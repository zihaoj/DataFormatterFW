

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jV08uKrM6FB79KkWQ/BXj6f14A+AEGYHCn1KCZ0VbNfDrIZcnPGuufHJK+Hv5nm3s6nRgyKiM9sc
4F7llsu1fg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mEgnJcfi/PWt6bgCaWhRPqwq5IjLbeR1jUx0MvpCJwM2ZaVfJri9hsTkatXmdNCcUA+lNz/aeW/F
sDcOGbKVVTg1yq+5snf97hZTBqSUNglBuzjNjNh5un2CSV8ttVXR1NNGfiSI48u+j4z+zgRCHR/z
6KlAJEcuLgnW8V7gP+w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gAWNd8trXwVN35ZXcQr9pZvhMTY8Fr2BewQ6CqyRY9m78MkTXCZV8O3jgNIOdO+CocqGe2s4kyvH
smrgW9IF2qrCszLKzkgc0ZEvJzHuATyAuaVMmaI8nwX2gS4L+3zO69yyD4B0lZrTuzCLd0Zrmf4v
y5BgkFIcSuXaWD6dy1JqXGmmj216DtACzcdp2QPhyp6wUg0bGBZyGE5sBbXw9J8FWjPxIpsSHV4Q
Vqzu41k9qYmSRywgNXJAIKQeMzc/FKVfjJz8u8Mlikz1SBoYSS5MQs1ZNvIJKZW/3NATqtg3O4uC
7XLepcL5FbU1FLplwJkGxjzuRwsscvZCMPf5lg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d07uexcfoDSmo0IeiZkVcW4bOu2jF1UYttWAexxKh/UquGZgKoVQ6QMvsl91Nr8PRoO1v07KRGwl
QHjbK6XSxBwkxQ/l+KVvOK+R4+WnUBOH7oSdoxkKL60fMkQBGcezriVNcTrE7CDAaKZ4ussIlkQ6
lhRmghszBT4Zf+kEzAg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
daZKqvXPzEDHQKunVq9aTX0TrtCWQzs5E1QGwhxofE7fJMfyTgGknuSxjT9Vc9jsSwDO4oPkvfpA
vEvC5eUK/VPZjFDJeIWJrYuoZzb15vXOGoDqlMkexDaM10RH9rmQA/WtuuATZUA4JAXe4UtIPDyC
sQaPdCzVIrKkBq6B4iuapu/PBi5ArFwmPdXWMmbf+emJqSYmx9L9aJmnIyTlgup8Y9CcNEG8gsG+
wAGtBTvupjVz0FBUDgxxwqHRcyOQ1FLt6zne5zpMaYrv9U2RYcnTLKV5/OtW+SKBTdf6DztEuM2l
jA9Uj/GJLi6W64bmvtYcsl6/gv5M7/95K61cNw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 77520)
`protect data_block
lwHsuZKyi/FxgPWtJJA2r55LVwEUXenJ4/uNgRVduTI+DJQHwSmE8R9pGYosDzPyV+w95qkI5D1O
3dx/TRY+HbRDxKy/dQpyrtIKfjbxlx8+vtffmYj/TscCAjc1zV+5WbaYFa/ilgGUqVkx/XXFSXyt
6kNZWGZk3Wupxp23M7fvFGlVsK1RaVgVyjWTKa4+hhH3e8pJQhGXKm+WAv+RI5b3l8zn877F397f
x3cg7HnWjwAc8REY4U4URN5aCGyclO7NvkWT6n66LgKuzTjfoDmOHDyvxbTm8GINWc+icuioMNpR
vPJuHqWGHGmcg+jqO3zyVPK/TSK5E16C6+nlLrR+b7kW29wMVYLhfg4frsiYmNyno1g6FqGOP/S8
9yabuysXNv00LY31W5SKQcb1qsSdZg5FJA5tViB850OfAKmsrKTbUO+NECT+aUzZHN6q5sl75o+h
Su1xW8f470bgIIj2QCDyuD+zYOn+CVrieHXgupH+aP3gZ8JZj1ZEhjiB1nV3CGYaK2/LfiGcR1UZ
X7ZFCKf+fE2coZzQQQtx3jr45XwVAjNdVs/K0mY3XQGsP6tPyre9Gfk7V4pSviwvZeISUBjfUsow
Jwky+OITujVRsHsQOM3IWF7ipx6wAUkktt2fFMdA0Str9jucp2dvsYJc3MwFx1yUBPIeGGx3x/83
dCWvQ+h2SrADtVuPgamsbtZ58/p0nBWJ4cAt/4WyBcyPY+D97yCpUmqQydJBVPVmjHZBVNWdKUaZ
/TknZzh0Rvi8Obqy9krO7Hzz22og2CXbjvpv8wf9W0RXRUkKTHVRPH1mdYoYVV8cvG06YK6bTZ8s
T6v+aSTsCi8uPL9amCxn0WLNTdcdvvVxb8KVoRVW37ae/NAma+AaC+rO7VDCYPcyNMfXRm8XkGS6
Bcko/MJClNprf1oI30LTXs63dzXPWKu8+TmYtciKz7MC1qRmJ/jFM8RBlX3pvIiR/XNcvo3gikA4
MZl/GtPQR5tUjG3IWd+OfmzuIvYtzBoWOjZM/6QLwh58rpxDTG5lO8J9vKX5dIFZBYu7rfquTSb1
sAUiKms4uAZ0dNXi/ThOeG0O1q8kAneHu/y5HBA3LWpMzENjpQLwvCVUox9+ZLWLCFakGoKsZt4O
59+c1CoieSBd4mukMnZmmj3g6dDTSN7MUuApQWURnIFnVyraHtYnoPmArlJIWB3tRdpIqqb5aPv2
MpHyOAO6mmRlPNMgm4gRdoRRuyIwpsicgd6w/heH+eKcQKSe5WmcTMX6CNmqzbpnmMwEMDiiXu2o
meH7NEtPYS+2jH+fcA3st86ZGvOdVHsCyqgCD8vdqA2jPrXq85he81WNUk3lB3gMWfW+NuRaEY8S
B+zLcVV92Aqv9libZGS34AZrlnGy4AiqxtiEw/N1VF/NVLUTw3Tf4AkLDCViE7txYnxQN4eS5OTm
iFxLgoPgwQ4ncTHLe7JXZNUfeNWCO2O6qi8vTrv2JIgG1HY/eB/fbLpruEXZPjgq/m/4ogSvbSd4
wFgf6tgOmXuSw4snYf86Yq4jqr7dYqeRGFLTJSxYE/+ouHaozxG//8wtUY+tkkqDL45OHy6qvwXb
g3oTobMk0k9EAJg3cIONOHDMnb8RZx7HX+6tlKiOd3o9uGp9IpxPzcu/s/KsnXKC5afkRl2AGOx1
O4aDijbjjV00dOgcPrEoILW7Qi/wVDchNuvcmfbzdooyNDV3CjQkaiTzYhAW6vBB4DMvWZ98iCqg
pYLnmYrWEtYI3U6pm9q2bOdbBGPHBigYfTEnnPqKOUgZOCyi3jxLZLNzW+SCRGoVtByFL6P/GjuR
GTpmBHL5YEt+dZPriaHWhJhxATOBQ42cQVx287fOe7mR6T1aBiStqinZWZGMnqASXvdIvK4q1EpM
eHZN5MMM9QXtFYggO5A6OHOEl00kOv7ZECjC0VWq8cmohLSiUGoYQ1EzM2miqutYue2W3sOIWwp8
zX3tNsXBCwkTk6Av4rNeqsj4BHW3NYV/4OtqCycePVYXg1tJKhQ481B83INz+n65NLfI0M00E+hu
1CGpdp7WJZpxmb3cXs0aVSjqJ6xDD7bwiTBqzj/xDqxaYm7gQDGNLLufW2ftaD8XV2dZjzmU/sAw
C5E6K5I684ThQCos3Gy4FANFSsQJpomPjwiJOPViP8Bw3iJyk+DFr64GjF38FuR3VQDy5gnokpYl
CpaF3W2Fg22dvMOKGqJ5Va+Q71i3hCge3rhCvPN/MAW68ZMHnLBFSG5Q4L6IJ9qvHPTD0m5YKO9T
ccsoOKhDY/JdrPcoo9tT4jP5oBURHFZ/D4U6T0p/9JPy+Btw+KTJWXLwnn+Y7pHphY+76cQ9dFYG
D6Mosc1xgJ+i401iAwq7Sz3nD3qQMcQQ/aXQQsxI5+JPj6705xHM3eVs89KOpSpKM4cIxeqPGcCi
5GRQ0LOCLIXqpvG+YJ3iC4LdEHlLvbzXcBA55F6d9URSxdmgBZ9l0ITx4i8jjr9u0zXq/deQjQJU
LnbFrYiQGOqXIZKEZzs/ROj+z0DejYkqUfNrO5FhhMichkrBZAwKlWGGTZBpEmYpnI4n5omL5z1k
UMRelUDjJZUfVTNRy7bZrs6UK9Sh1CDblfkh9QXWtDA2DZz4oN6A7/xGqtF0ZYCIjgjc96kcP4TW
fYeBT1ExnOQ9euqcZEC9EE2Wakp7QPX4VPOgSlvO88YvsBSjcj25D5Y+AtAnALucnjLyDNw0UlYw
TUh0s+MjFS/xK0TnE+nLT6XYZ+9pWI+zWGkCQ3b2X7kK4mwzUoA0NmDEtqzwAI5DpMmaWCL0+a93
/vFyua3Zjx7dBwkNi5rep5XdDlQo2pGgLwUhggX4q+6a7UdGe9t2cYp6DtotrLlg/HsOispLe2UT
O42MmvFZ17LKYF2eh/aPzfgQGj7IjZ7m/0GISfu9Y3ow6LnqnssO6EUW8UHENLnUISr/Y7X37JzG
3XOnGFLwFpGdUR7uqwlzBgJm/sC8lrtR2G/hQKCth6tp9EbZndPSFFtJnSX85FQwY/9VVQn5hLcw
KE+tX0AKe56GcDkYfCWoXxsacdDLfxkKQmZAsPJ5taWy4ccU//0JMOhUkyBiAWmex9V7dJYPHQOw
/bge3kNtHtz0LH2eG60cSmtHzJn68yvJg6Z7fcNyuW24c1bVG+gC8fo/DGNMwahn0gu7p3Yrm6SY
Qt0JdOxkPCy3673kacIbs/cVtpxWtI5fUv4UCxsuwI3nE4RuF8mADPdODB7IKV0mQx0w20MvJMc3
8+vmnfrXe0MIVgNS6N+LA9yhP5V7xfaTKgzTIHL6gv7nJh/qvSZlW96GgsqulO9ue9kRg2u7R/+K
h6EwZ3XIimQLap6/t6SvM44sZyyQGcnuD8ZjH92SHzJTfTMIaKLHNV7txYhH2zAuTf877jseixVE
jLellDTfrYqjMJ1NuJK0wpW6RfQZH4KTNQaKXV7/bsQoo97Lav5yMuFm1Tnzha2GZs12ErH52kP6
SLC0wZeDJa3GiiIs+vFMP7IwmrluE7emOqbUotwaak5IakyCYM7xcYZos7C61WyUzDsEv6C5tms+
W4xfXeb6NnqrkSXumvH4ppTd1RKljeR1MMEU5sT9eLfVDLKGw/MnQB1PRVmTFfjzvr74HSc4dbd+
BFXejs7leZaC8wnnFm64wId6vua0XlsG3ZmHtWKUOVj8nU6NGOXvuZR9+VZzree5IVkkEeirTDEE
L4B3VA0f1kCE6+nDZ9iBKHUuAEJpRbDxf/DZB5UkS0eeUTsF3sFsziwIvYFaszZNOkYlaYQRIVmd
68l4jy9QecG198OeC4qxaUB3mQ6gJmBJrXINDDqv+sTqNOWOjcAn5d/9ALJdanAT1tVqnEar4veA
Zj4tMh9HqZDNBuplJSPy63yV0Yz9TWPoXEkscUhoS2K7WOt/XLSontx2X2gi/gcLtNwSOjsv58oU
46yY1B2il78qH3POilOwbUIN9pLaNjHeLE5LoeawkK/ibbq6vYz4RJ6ipY+exicNvu+nksVmdbqg
vv/ieb7zdqv5yC3QTivSo2TjME7pWMU2T+l/+GN4Agk4wK/Qn6cM2Uus2kW03nVC9+Rw0e0Jav9E
DN5LkzdFpdy814A8YvAiOokzIjA/dLIYVw4qRJREmdx6BYoP3q8ooYt+Bc31oOmvidegS5VlePPX
M2UtybzIsO9WGHPFV/V87Cp49W/LYrFeEABY3H0MkQnkuy5hEhaYxX4HyjuyO2rt1msXW/DyXT+f
JK82KLs9YLIjFaXdSMLp+flfPixwAMzzdcpH3ew8A576LfHfdhSBOtCg3g2lBw5MB9wNIVrzEvAc
F1hI8VN08XpgHswer0SQk4VtKMuUbPKzqHkHyLqGyExKwnJlkbJzaNNpRqV1Z0Q0gso36LqdTmeH
nn+X6PYx8kMnc2ubppIzahpRrhf4trCVOFBlRKu7wOUe7X/0H9qv/8p8k+IMaA6f2NwFU1LAEp2w
55FfUjNBFg61p60orz2bh9lBh+PMbhZ94QsNoxges9rnf7okqJa+GuArxhYlSmNrhM1vrCZ3kpVw
FWQw+M7rv6R/0ObtyoZmgXaO0ZEyceqB/Uu6eNW8DOOb5dbeSJHyzUQq2hwFvhKbiLUod7iAS48j
ez3eEnrxr0MIrux2DthHTEo7mX0an+PcZUhXZ3FBYNciiSa7ZKVPOmupVFYrkl78h8bGudnUYgUk
fsERVyEoy/cuTZSYe62rMyapkuRCj96gDMzDym4t/LmJ7cUY4UwHzBd8hluKgvdrxfsTAt7NfCrH
/VAFdvTvWEB92orDupORcSu5z3AO/71sZEqelGg+AtbeyFx6dUCYbD+W99qGEhpsTn4bkh29iWO/
HfaTzfEOVdP6nC98SLzIcfkE7H2YcxfMW34NQYLvgSksVYoTQ+WOWMy0svyMlqkZ/+rlLdl0oOVN
4vHEj4IVTwWUIh71wlYsQUu5L4eizycqOz+pn8HxlGknQZx8giSqTbaDhczPpThy0lupdpx4fkrF
e020m5eng/EV9hn9LgmXpSi3facLWV2CMfj6tGp2Qdb0zf7IUl/K9Cq8xp44MbK/lr7CvjbFD5v9
9H/JaFCy2NrYaG7g/7yC7Xge/ks7p7WVCGBIXjgDjm0sD968kYtcKqROfJ1DRlhlRUFs15dkD2HK
k50JGLxRz91vM2SjR1cMyj5MMa+VjxKGxRmrKvGX5TZ1ULN601so3GzVpDlm+Vy8c5G9ph/nx+MT
+HhWub4qz5OnYN21GbH9r9lD42zpNyzGa+Tfygw/Qm1lyf4uT4sH/KxsC/lSQm5NbE6oG3o19VEy
Nb/eMvJKIU6DAO5Ib4ag3xFswoLauu/JJf42piVRhksqgKL36aKN0azD9KjIB2JaPdN9dwHH90rU
uWcMt6WmvtLMMOH3L61lsSrEAkO39k/SUytcy4chltlx0qzMHZqod4aHWm9ZqQvf1FendKLHXec8
bZRDuv13LVhB7+aIZtNIhyTDMkaZuCWOKkP+m0ORcttNCuGcJRTxYJYuhbuXeZDG98aTFjzOEynP
R0Z+c6NuDj0nXo0JITp+Jfx8wVWWKKDM1nSvbvtqI2JLOy+2w9aiByJioAT8uCr0h7v5zF6Hz2b5
qPNNJasFSUmLbNLTG66TFlam1GBFgRF4F7yfIuNYDDkvmC/JRWwMJoMitTRuYSuaJeK0W8iJf6V0
hU7knZdJVq1q84FPNzewdmtzC9XpbUFeYHDY+wN2YpJYFQUHOsT5eBaFrLWXc/1rjdWkhHCMIcKj
od8Z325PrdyoKZQeOFxjDKJw0zUH41UsW05exr5sbKNLu6lIqi1ZgDQ5gDSZ2rJJqjzUsO1RNILT
zlZ02gAWfSbYshz3q0/BRxSMspt96ecI7ngnqk8/KlAyJxcE7GtlZqIyer2V/7b2WfZ5HJVQwEyx
RdL2sG8OnDvrWxRqZMPBNa0VW4gFpZsgh7U8pq25O7DSHXWsy82OSQtGVH/lFlJQnYx3Ir8dWSnR
HKZYaAU0pPCWoTqC9xOKZ0LetMtWcYTcH7HYB2NFQs0ODehf5Fel5oi7PwgbB+uYjy4CLnh3K9WZ
5YQEp5QMp5s6jkCtiKaKw2J3I9BIM2FoVUcPwGKuzFfvn4zKgiL+Tq0T2KaR65MAqYLZXc5UJvge
vChf2kwW7Yckkt0DQ8dE7aUWfcvNc7G6KKIKFTjKcDqiAvXoeGnGjHH7e4/57j+OIEouPkR3746a
SM2BVZi7pSth2XGePnnKJMTIQMF8g2nD7W1PMSwxqmEv7ZylAnWmc23CHsw1gZCuew5JpGwXPPYW
BTJ1PWCs5v/CQadU6DpJ5aoezuv9G3mTYbDhZ/xm1a+SzCsfddRQO0YXAMHzzOqG2pWv7J9QPoEU
Es19rPyUosjLoEd2TmrD9JmOPDjAULNYNI2GVx9iJtEjNSiOcCwaCn7Frzkc5dJm+1Wq6Qn+sCog
wcVhj469wQn7wPCk4xW9jkTwoK6YCPVey3ueoovwI9BnycfyJqwxsHVkjJalo63kT6qktpzCBfTX
MY3F8Fq4j9NMQk5J3HQutqvGhixudIW8GlUXNe0mdY+vpWlOEDnjuLAVfixLcp6e5sHSqguvo6q9
ORqxDYwUeTYQYC/mEFXiocRHWviJ9BII01/bsNGTvsSnsADuAWKgcwFPQ3IGqM3EFQgfduj+O2Z6
78Q2vtp1Nml37dXE0+gIqH7IGamVefag4ASwOta436ghSREb6amW5r0NKHckQ+YUV+m1iaruV8xc
O59C5xlYXuR7KXyOWpIxH33N0lGTvNMvtgah0ASy7EYbGw+didRx6fXMvq74eB7Hm0gvffLSYHjD
DcpNgxaInLlw20Gs01z3p5U/BimQF9rlOyo0mhOpcooNrs1BWUfk1BiI9GalFfhzrId4czGBCsSw
t59jfldgAV45YnrH7w+U4q+iZLaiKLXLTnSpBcI5JZ2rWLVPUSkuonigxeNAiHMTcyLDmrYUdD/U
69jxdIdTMNNWhfaNiP23DIPEZQoGbBik0Xv9ERo2nEobq7lBtDm7YriXZuTz8b+hW6VPm/0M5hzM
heQn2yZ/dVGwcS18eX0l1Fq7YuwerrI0nYaINL630z4rm+u/6TCHdGfQl3nJcZyrS8bU7yytkFU2
ph9tZtc4YE3F0QWO+0OGHXu8ca9xNDss73ZVjSwHT5+PTkvRCKgucGAiViw3wplcFi5mJe50QZDr
On3Eurctdl/i3s7OjL4yI2B77AoWCZ4NoSbEweGXulEC+DpSDi2m7M+au2YxoAsQ/lm2VfG7HPpB
6mfkHSYSgq4HuuPNp+BuvpkCxfJG8+1bK31p6rH2ubaIYc+9KKNgMZAvEzoONTb9FOJLYHgTcT62
Fm/239XpSgseW+Nb7AAsYP6CedHoxNyzq5woU47FpgHurVGq335tCNOiY28zCNJYpXasfI5nK2oT
VG4Q1unHn+7vWkhYm2J3QX7Qk94BcNA4pfVRXqWxcOgl0uUaGuf+ST7lDozyHp16JFgmuaeLEvkt
XX9mhiOQJ/rXrdW6pQo839rwiVxY4ZRbmBIHVP7+namDy8Na8DPDP/sMJHw50KeNdOJKmIx6S7Ii
/4fhVzXlylWZ9Ktnc9yY6UCJFI1TBAENFK6f5eINOL1U83E14HXMNNbwNq+ffwikl3amtljBCR6i
3Mxev2g/oCl4h+Zabm0/mWN+qy4fhlkleccGa5KtqBQBUAuQbtOrd+R7Q2S1G7fHeySLbe71uM2T
IKtUZzF5mi4cwvRWiqeVRKquk3uIwmGm5vfW387eHBH5mD61SmBU/yWRiQioi3QCj1Z3dkcOwULQ
TNmi6oG5P5CjajtaVwdFIWp8mXzEfEn5EvjnSEyIXiyT0VwQKy7GFuQv5p7tVsAEE/Z+aQF3WvKj
wUxOhiyyHBqLRwa0hwDJiEjp60MGm6Ze+gh4urnjq2t4mKOaqtc9lGQKbKWsJtsI3CnDtWlY4RgR
jU3UT2FtPe4W/hTs+9aq6CGZQUiW6NOEqSwntYFx2+c8qk2k4ecTsUaSTV8gEpy5UVbix3kjwzL7
Arz//HR9GM7LjGmdXra9tjvAgJGKPNk/BXCzF4I9ygfcQ4cgiyJTQSaNiYTCsm1Kg4F0B7CPZdRP
zQG1bOQOnx/oqmZRGMHcxH6+kh/slcjkloGEgxSMcHI8GgH5DJL9gIXj+b21nf5GY/uJnB8/Wvfe
nZK1/UTfeJO8UrSaBvySX69pxseK3nA9qBuzExbpU87AgWBFhkRkc9GhJTv0YAXLh1YEwjIffg9P
qzU/wLR5jtqGoEJTEiTd+gwd0CtgwPBZCJCSThVZ8+heR3YPVYBYISeIVgPsArZQ//4bnX5zzV6F
H7QewmXf8LW7jIVfoVaZ1usM1CgTV3vQPVdQ29gfzB2JflSDwNH8XJm+S11Gw0trMEcZ3jznj5su
59YUqMMB5ICNfdTKNY9wJrq79P78utVrRfvuTeIgU2sjKghn2VJkbwEVR/xBQlued4HXRJBEWK/7
Glw+b6OOVxIxSRJfDmstAs0T9dzA5RqaGDP1OkZ/I8+IsSrhtCDG4hHLk+LUM1Ox9VMBrQp5XAhT
Lackj2Hz2qZiZ36pYiIgq/fxJMV5iyzFLc9gIomODxY3QAV4uywBBAsunlqqKxzpqrV+uAgkzWkT
JK7Lx+GEEqzEYN7QTJ5fYGeplYF+HsO/zsureK0pB/HB+h4lnQKWw/BWPef7JGU6rfakV9XeVwHZ
nJPR3I/6Cl7XMlukfi5uo+57PAM2EX/eClfA1dC8ZqwIlMnIhH/bn73vXI5YaX43Q9OCTh3L0qha
NAol2DNJ1nHUlEW9nhDtXZpIMpgL6Euf0Ac04SfGdpRsA6b76q46n61db53bUnJGpVfjkoF+X6wS
HuKzH+BxOpbKwJGsMtmW7NRyMwL8j+LcOQz8Bv1YJyyw9pjUhw6QwLAlDVRJMNlLNb9CDdmEg9+L
fGkw9ejxmtTMRJOwGAAqswBJ5d+fxFnFl/ROLit6obF+ZJcMm63Kqdyub8kaVvbHYkm/Ojr6OSi7
su+xfY14XSrBfDgXmESkewAYtXfBqTxR9dWkCZZl312SwZMMy37DQidALDEq5+7mozYlC1BiSxMW
M8ehjA8nP43/BpDxp9qsYlgVSvP39k9f7NX/bDHLxNW88NFqVzxe9jvGE3XVMTrzlgUQIF47R0XJ
ko5Vx+wVkVO/S1zc/iz9kr1fNnWnZ69z0Aa/kaiLt5+ts/E+5heGQiPJg+A2kqeelwI6rKGRzFeD
FRhsxs5FgNLYSHftFL0R4Fk8wMF/JOy5KAluHbn2vQCSb+KwDE6UUltrDBtQK0JRea1UV1VTTWMq
o6UE0T9VQNypDZ6Eh44kABrs3/ilZK2Tj4N5QfpBIZ6SI8/K5RFrcEMbG8N9yrDPKEGWVFHR/mVK
OPdEw6byg/XZhi1FxhYIcdQlR7R57pmQuIDJFFSn9AtFSw+/vw9+t0cJ8IIn/HSVI/beoWm5Yk4s
m9v8WilOLRoxWgF9fS/pYaJM+cpq2ZuckHOoHDGhzJCrBoik0PXe+6d0EFcfxOynAGXWQx6TjmUD
hpoftYCR+jdQeq6bXlCHWE062Bpx06pJFWoIUGWPgxleQ7Dh3VnhcO9K3EyMcLuexT3HNWnvEh/1
jXyPG8i3amu8sV9YTGFeQQUVX0L8Sdq0YZrWvP2mAebHVAllLu7+ZFZPHhDcChRZGjG5XzOZ1Hbs
gfRCdzWb75pac8Uphg0KhwVVQrCjE4e+v5pOtRwm4DiIWMhaqCRiqIRPKuBYIb4XrMznXJ0adorO
tl6pSDqF1unDnh+23eXHABmr/5Aso3Lez8WNK0h71sox1JE3fLLVBdCXbCMsJz0KnQrX1WX64rhu
nsDdeiUO0ZnEwWT1aY9vKDQRr5N5hH8rB4pNVx6DgYqjN328+YRFu3F3Vt/MTStZ95Qr/8r6ogP6
beZtrkAO91ZJeePk22zF0m1k1l9/GV+AStDm2aOW/zr4ao+t0gVN29czgBRhgBa+7QOpq+M8B2jv
c8FgoKVWZ3Lv0PCT3X6cJzDOWRIUFOdKmByGwTehHoSnR8/yz0qdgjzPIPIS0rtE4sIYsLgJli7S
lWTkM74Zdlixr+A9zJ9hqVEjTcHzO1vkG8aNUIY8PHuQt96uF5fgT/m1I3Y9X/aUslec7GFqHtp7
DyvCe2AGh8JV5whXQuNg7598ZgjiehYNwdtUEoUYNWl0mX8AZddzN9YlbPWaXzXsbG/+mWwwktpM
9d1Hd+J8NmRkMe/5oEY/uQ0e05Akq1uolzAMBxe07DP5OGauBwCT5Xib8BPsmM6npcXpJwzVIK+J
uPFcK+4NT9RP4xPIhCa4XDLU5AFi6GmdaapIFuq/0ZwBQeJ6tzD1883gRfMkU51PCcr0VyorObn3
faRf7vxyICFZld6LVVCquup+DSmd5cPNr4Joi+TmiRRbLeCWhS3NEI3cVD+Mo0LhYkKxZisaXIDx
R3SQ/of6BGKV30VBkf6pRurdRsT6599MiS0Lb1dVnW0SKvi5Z+PARV4sJVfjADN1X9XeX2rit3cG
PsPhMaqEcNJEdWr2o7dHfWPjvPrXemY/CmLhjcR8nbrbotKIX6C+EBDbHHtcDSymeqv8XHt/UGxW
cUjtmJ7rXu7a9u6TyrSBHcvekZGWI/e2aDt4cbxvXPMB/rX0pq/sWn12C4UVYezCL1ehZ8FcHV7X
2nefZU+8mM/NtZYusNVx0hSy6T//FGnCX7Txh364W8msH2FyPITwpdpgkU10GpDSiuNF7qQ19K1p
ToBHr1bGHhgCTcPbYkcu6OkxsZa8kGSF15QtWGBK1rewdsfFmlBpGVen6o4iw3LDgvLRyueeDn8N
XZaZpgjuPDHr754whtmGE4hqsCEG8+/84MUf4SjjP0rlthH2eHykBYCJhyda2rcC1igYFAQoAa6W
CVlf7Bl8O3cRmcd4HLGgipE5f7+VTv8rxU0cKx9Cgh7QuoNGPnnpkdQIEBenS8ZpLSAIk/g59tLY
e7UwTb0QKWAfYngU6YcNZyXCyYarRXTvr9XBPz5acTwDdtaNDmO+28L6B88eNdbtIXiGJnpGlbKk
XQ0TxyohLMRbNGmAG9EmJawaEW+0eal9nG1nOAR+5qeUInpSUaAf2eK68S2YqSpjxnRdyfz+9k+0
l1nTpgA2iZSSbNWpQN7zih5tIjf6g2OY/1IA87CkM479NlxV65uVBQfO68gKI0GVufy8b3ENMYMB
aB9zQPWkmR87ESDB8ZwIprDyX7VZQsscZVIdjrNQmOzZpQJAhTHzOSyaqTyNPn/clSGNVD0f5wkw
xuEB2nI/A2oPZ6GRijaH3N3/JlgP+FtIDLF3h7Rzsp40ppUImHOLbCeTtK4zDyOMafC9pZfu8TRw
J2Rs3Mf93aLZY8LqVtBHCRfZuTycdkfC8PBE28rND/OP5v+juOFu8Ccmc2Bs4Fo3tKVUHAgreJhp
Z3sDlojXxdprGAeMXncihj5Fr1s8edC1ZdzE8vZDaK5WKTAf21azMGynmBBObScV/W1NcrhmgdyP
CLAGa7g9kxOJVFs96rtENiQ42RopjNqTQ2EtmnX7Sx45A+eQr4IhZzghXPFEmxtMtKfGfd1ARgWT
nxnjcOSuB2UOmvAF9pTkHaFCrfrg5yAlVRjO2B7ngLgD4ZgLaftU91Jir4dbFKfBiKSgAoljMkB8
Hkh0asRhVwnEjXv26bcTQqt3i+rhfKxra4OJeMYtLq0hJsnDNvHzNOzzx9ac5RtUmVOpbgj+iexj
+l4KRKAcdidL307ZQEVYqv+n7NwKryAABdUqCy3sO5pd+ROISL01h4iQRabYQ2vhH4Nacwa3tmrL
e4abd9l8ISe+f1nI5OAUPJqcTF1Lt1csWnOK06geVjhQIPIPUDr4A4l/VJjXIOuNfAejqvHGtv1a
h9DqwI4euxn9dNLhQwpde2vBb0UsXOb6sjSScQNiuWVgNaPFl8jY8p27lCOPEoPbGktCmyzoLLqE
BRYPg9bO+GKgba+CP4bV0tKgZqnsGTf8CBXt6UIQU4450lG4unfrDpEX3D4QBd3TQce4eK/n+6zd
5854Yjzh1UESJVJ9MJvYrLefK7wXpLuz+1Zb8inRDMoVRo17TZNJqFqq5j45GAt1itasrlVwgM3O
3vkQfthPfqGg4K0dl2QmAQJo7ZtWYqhFfbcrZwdWXH8Ix6Tf/PPrZXgC4AQ521ifnKHlhY/3X5p9
/hLMgnO1YZffSmJ4JZJqfWy+5O1I28+jC810B7DoAhN3VNMgu3DFt7XjXk8C0GF73Rk1quvGKQS5
HFme0TTe6P/kQcGI3B3KxE24fna2J4nJxWvlgIdRupaoc8q/gaFsELh7CgSFJzT7ouoKR7SfTNQH
sGXmG2ZP5PuD2ZPcpCIXt+uSiz5actYcuo3ButlMvL0lahmFG6Tjiu4mNMIuM6UzngRbBSz0I2hZ
yM7avfw46nyxpQgid1spYK9H1xHpB04BC5Bp6TFYGZbbpZsDXRCJMKKEmNTXrNBl5j0dm2/CQojR
Snx5596YlU/Q4UbYLEKMwRoWVxy6PVAg/RKc1lUALu5wrNFBLZLNeotJkb66YIxe5kIcsVPcs0tu
YKdexWoJcv6YZq6Bo151AzPMV39dNMP42V4/1z7NyNjTZMBD3DlzSsm5cKaqCZFph81YhUrQyRDK
pKkgTx4uYcWBgyi08ywdctzX/YO2BHjeg625uyj86KdIWV+lCFl9/ep/kAe6ZFeI2161lahEPfps
xAfanLTDm9lqgKVGX9vlkjOE1/9JUN+35iT609WszQrGDkrTe5+LTTxhRqZgAFoa7Aqp6wH9xBcA
O4/n72UFI3vUUE2oJ4vcKqLaC5NQkeIphxGG+ASzXqlXC+ENk07EIW2i+jtY+W0LoxcjonOcsGQM
geZlpYGDIRpBlmirNU4qMfRVe0EoZwsAx5QpxzBQlehkp/p/jAWcKnW48ouwQ3lHqOeL7QHLUalU
fAGg+slq7cN6HkOblgEPHTKczC8mbWZ9oemg1y0pVWJ/x3Iq01IbMjACtfWiCEFmvPHqR5Y6t7TE
MT3NjrffsHUs53H2XhybqFSlAv95DRgQPn++9bh9k49vUNWKEjPXIn6C5gQGAjQzH0Qla7YCpdR5
ZHs2ALPjOhRqOWMXG8r/ykfPY8vBAEpLvn7hZfVdr5akz8LyqFyH1d3YkYsfmAczyzyDHdWHPUhi
T8eq4FV4aKuZ8ENbZz4UkA5HrXDIr2qC7Izef1svJJ1KUGKKIUD5x4O8Xrdh2Pk7YJH94H4B/vcr
EpXjenQ0dFAwbRbhRSk3LB1KtdSD2UkiLgjBBC1/Qd+k0shLo/q9MpzV3po/ZTEC7l/LUM7kFDCA
vflb6eSRhlg+CrOzllLVCY28PUU4yv2zT2LLnENwJD4GAl4HU2q2gUpvY+PnbrDfEAiDz9aXVmuq
zBLppqYl3ksyqktrJSRm/fWHxadLXXyvkwQuSE9tsolHayLS0guFJLSQlkbuqzNJtrjrXg9S0pPj
0D4ZsuLEjvyyHxnOlnNKz72EtS4tTKStZu38XwAFr8CeJWSvQcoytJSmY8EG+7fHA7P5Bs0YI3+9
WeYf+t8sIhoMN43gu9Ei4Zxw175UxKeElECiSfcRSkyMO2Q2q6K1So6+7x+jlwMUbJGvlOdcjxt+
ncqnFk7CP1P5vmB6o3c2vabMleRf53KNIDaTg7erB4MsL3S9cEATr0OTVTAJCSyA5TZ079mOozLD
5d1h6C2MUdu4ci72LZwxFLpbsjzPptCPSNARN705Ax4nBhrhq2EN+d48iW9hUAyG4jjJuPQp/0Y5
O8NGq9w6e/CpYxdHiiB+AHeixfPy+Rb+Ur9liP9qHTWhfc6Mz7xLmiimLiZ0lvQr5800Cae53cc+
+heryfp7ABctSD6Jacbj+L8M5j90VYA4+32q7r3OlTk/JqZV+jxsHQEwwVrdZP5x6o0cIhXjWNC4
WnMm4OpiKsldWfOSdCpWKXc3oa17bGKd4QLYqL23lIYj3LvNjyrF04HMX5NXV2Ol5VRraAq+eefh
O+AcDBnnUyiXgYLGGX4EExwhPVkQt8GIpShwvvLmWhYi1dkgCJFJHZz+oS0IclPGlkSJjU1SgvFD
dRg6rV1fhEWgOcqKLtsoGn1BLC+Henw/wmwqHql/1dzYsa7yADICN8i73qbYRCQQ5stotMvXGg7t
t67xFDA8VC/C3G9HYLBxli3Ar5BiGYFjenp1aY7F7g6aU/OR7Yc8RNHwSxOE6VZsdaRxT8v50wYL
2mVxCx6FR+Vw8p/MEW2OqLTdIpKh6N/gZRDAVVtatt9DGMDrvfMz9woU2NXUZ4+S0Z18E6l7M/Wz
1rBtEGagVynk+MwcmkJtbJ6V5zQcGeFvqon1r39aKt0rwP+NjBzRMjF0NVNtoarQopCgyNIn2flN
Zodyb6nB10RMnj38csiJHey106OvaYmrScnxJYz9L9CHgugwIVh3/JegcIulA83i7JfpOgSJKe2e
T+/oGZi7odrQVrT4e4ug1VigieRqyNNZkRRvwUpL0HXxzkRJ8/flr0zK1OniHwF2U+lDXtnwoCBd
Q4nkrIU+TJY/3mDEqf9qYEROZywx75QhBYQpOIwsad9KlJ+VKzlZoYJkIuF1nzW2aDeA2K/Ybnho
yTmVe4YxjYTwcJFDFPoUtBD2Q/z8X8q5Kp5wLS+aX/+oH5lqcokdo9BSjNow9TOWGEEH9R6E0APw
4LzB9s4gNEl7maKkIrt6Ym4e1nYfJ4H8eUKn8wJo6RhKQnc6Lhw4wmWO4LfMqsmvSmI71IeW7eHh
00sjdcKxqkvssS0JWHOyRLFpqjSEUdlFeqUkDPNJ7UDOscYU8hsmGF9PnMmSIdUi02uRf47vQIH5
z6Izxloq0gHZRhan/EryjU19xv8UdrdoCAaBMgX4+L46OfEdUpvflZYHRfDSNxmn1kpuS2nYjKtn
ZbTM/nkSl7ieLR8AI5Ofb9uyi8QSBmvyJwhHlqYw1ZZcXp5vEGxCRax+q/s7zrbveutdqWhvOAEP
eTBfJogHvkPhYPfWzigWRUQDgbYbksjnB2X2OMgJJsicxSc+K9supRTm9+oh9x+ZlCzMK90rAYWx
cWh1hIgRokkg0AJVr3d55Sxjga7+GiTON4gQ29SmwR6vBDHxcxSf2lLOX56UC/Osh3TMWgxVVzDC
pRI1J+PYsCQfonOgg/LlkhQ2Z7AaAc78idzgVSYTPgxOb7193yMx1wQt3SB/oJt7PxmP/T0gKSQC
sAiM8IIbiC5SjiBhWSLO1iLanskOfcVOnUOU1+ifu0zH92VUKGzrioZi//4cHXL7PVzPwYAPO42G
cX4uMNOpXR4JsSbDWOMcmnQod51CaQeJKJdwludTuSvoKdwC2g+1W+lUHZebaHtCDyn0ECkv9Trl
0FIkkYrBtVENzXCwqJt3yRKdwSVe6RBbGNm0Fwr1NperLTz48X9EEMVOc3QJxTHZnHIokBpgwyg9
omVssYUIJcxnhvlnTTDGlXE+qV9ulbmtxeCXjulOHUw78LlhTXL1Qt2+rGE+LPeflGYH5nZdpuNF
a7pix6MJYEl/nDGDlWUsSLI3uW4AA9U7IfwqLF6nKYgLna9jhAwRqrF0rsbkIH0AWHYkhV+8nZH1
jvOAA0N3GS+iSXCzuoREQAv5yYpSeWbmtUWrmhXFUxFsyQFZRDEXpuIPfOWxFMfyvnTMG+F+l8e0
ODv73VvFbAz980zLecxSW0QQp32ojELaH+tNxfDUHO6+li/3ezXxXafLsCs4sKQUstCWs+8PfJ/9
YMerwT2IVigRv3ExuJdBSZbkjeoJfxTmAun85lJ0WpAA3S93kV/8IJNFejn9q537BuUEUdo2gRF9
n7j/+242UIAcbeMLy0pu0krjJomjdqIAbT6cqiE8OzwEhEKyKvJSvTnrDBLGrtHv9sTKU6W4HAa8
utRsHGszp4WkqzTEB7T5G2FJC2KJXzDTc+20Sq3OYwKR7Wpv1hCq6s0WSR+KkyvWuMNK31V08v6T
8RGAelxyG/+Hl6iCdRHNpQZoEwDeQqjlf4VAyxE0JuwhCH8EowXxmpxZT8fdKkyfILlwCdqPRCW2
kSpee+VAU6+lSq9NqBUZsvMh8DRdEpkQj81hbAPqTOjJfmXwXEAOgH3oxBaSecPibUCi2nXxyR5m
+ZMyG92vFlzFfiRf+/b255FJkVF+Nzjjjd6KX677FiG0MiYU0ZkQxiJopN5oBZ/3vmh3OOxmJWIg
ZzvRYjIhcxPnuEQfPKLf8ct0QNrQd3xBbguceqsroJPBF5LEZDODJyRGUqlcXSrZiFn/b2oWZMzb
C6VTMx81lFWIWcA4ltqX8uVur31BZE7L6kb+0K+RzqGzRx1gFmM8M0wk2coYtbl0/9J39MVT4xZY
iwOYOks19T3lrUE1qcSDI1XR7wsh+oLHQDKoL94x4LP4h48Oez7dIz9ol6SsnFk2zgm6O6c4syWE
vagQ7HnMfO1maZxkvjvQXyKK0VoJEiO9Lr7zlmAr3I+JCyjNw47LnPhfECAH52K0LMMBh4lpdJDG
dAbl0dF41ktchWl6gIMgiiTPr1KR8anLIWU5wJ27bBeBENxaxPpsQkD8NKd2QrThQXxaWH0rLZBl
GDEUjXxjmQ8YU1mmN+FZjkdenqbOmxxuhVOc+kaP8O33CQZbiiY0lb6fNHmyv/iLK/OEODTCwseU
lm5sU0ZPoW1WGpC76DHKwCp7zesTdViQyfm0swSQc+wyw5+hiJ4fAOvspHE521VLjX5HbcTc3PoK
7GvsULSO+qQDxJ0UToTlPXBzzcZnCxfclKAvLkHq4MZbhFZwm+B+5iyVHiXhnR8T0fXdTygckhlz
q3Rjc/W1GQbO7dozlstL0xdi7JN+470EGhacytv58WbFzQ3Gz7SAz3dHn78n1PnD8JtcHX57YWbU
ps1YvWWm0gqhkHSwwCT8EtMl+BSTq5OHgv+V1cSO2QLdzIJZd4YIShx136cH6xVNghgi1inh4PhY
myYrvptHYQZbudWRHBcL1Iyy40Ylaacjl6GFTsqI3oPSUYLL74g7ThaN3MsptssDmvK+MogjXujt
8XCRWmCn1VJ/zOLhC4BDblUQCd0E0pdhzNodfFbhvFVmAz/km27cwh8Cgg6kkv7xtGIrGp7JUrjr
3Jkzn1usAOXwdwSUiM4JCHhWyAeg9xO2Xohmij9YkLTbNXMqW8ppBiKQ5nvxQ5e+JSijIdpPmmGN
vW87NhQ679qnBp8VS0Cb5YWOKQPpX4ETYyPD6dWz1smHKg2BCgBLQ41BOjIZ7VtSK+IbXL9NV6o2
kS8fzpaoMYwuVy5nbVrZbBaXJoXSaEQjoZdzBK61+T+uYAlVF+Dwklw2g3ANdU1xTVGFPXwTNHkq
1QqMyFEKeJalyOaIJ6BymT/psbtDCPR8eQQliTL/o08lTOf8XAMLgtuLKbpk9pqrw/KLVuIXYJKw
vgosCIoWvtch6ldDERySIIUbNyJVBbrlq842WWLOucSdRQnheEogZz2ZglCWH+DqR5aCt/8iIQ0a
6NI9wfkrRe8QA/ODyV1XkCOEgqaBtssPps2jxegMbexlbumz4fZe1XHRLAyRB2wv95GvW2Hy7VYw
b80WfCJSmhF8hcYcKCSAHSHAcKKyZbiMOd2B5wm1F8vW8qyc4TrVT999ryec3aLXfkVgCo78Lpky
O7XtunFOH68sq7BjjBwFpWI8c4NmwnQ60LNOf9uG/0lpayqaiJB8fjJWKyKYcMFzN3WAA88Ps5iN
kB0dW+W+kRuNOEudAv2ijihCBrPvlCl+BFM1ikBrdXtVAgyjDFvW69eVSQ1QUuF8ZHmXMaY/ymrU
2fnDM4ruO0ZldTjP7G5khAIhaHJu7Mc1LiWsf65prhb4CT9YypgwEVT4iwSFEkbVyys3FqsYdPum
VyEfOTXyBnIauMjsdcrb9xcdkmQrf8D1kZx+dSfn5D32RDiKnF6WTmyLGUdHf617w+1p64II/v5L
1293Fca0krqPqCtOvulV9POPbWF4F03DQkV3xuiwi9etxLlw9ZdCibPyCIhhULhdeaqnAEBbKhDq
x+w9PNq/IN2bkb3Z+T71NiP7xMyj/JbQOsHiTo2etRoFerXJYpq1EDUZKVK2Lqa2XubfIIJZX3a7
1fIyH6HedDY6MxsUHWR7/wW/jIpFxR+oi7urFQtyBl8lcy2v7rUSclDfLbuujpRn7EK4mU9I/A56
0AIKKpnyruXc6YvQXuj5s90/aX69j/ElJvoZNdqkgo+k4VE6ksOIVZrJi+wfngIVMdWGUuk2q1OT
DskGQVhjUel53teMqrT0uYfKcsF9qIZNADzdoUjoMYiWSRloKLUO5vJXOb1uBF1UrKj9C4dCmob/
b23yBbJZzcCsVcHEPh2vgoIlL8MF7dSq+53spnLB+ucy6zSMe67SyNFa6y5O4tVeVzPrZcWj+lgZ
BvTOPmTWxal3h/U4H3cxcR2yIRIx3Gf3dEgjRyoSDMFA0rxN6Ibcf87WfgIW42EV4aGUDXBacMWx
yRlwTXEKSelv/yiXF8Sy5nEFPqvfw2PZmT2ln9NeIhn0J6AczzXafQOKH7S/7oVur07xxz9j4k4M
9OKUS6i1zbHLixOAcAE+vIFMnbWUpRkCVEacnajzImi5r6KSnXTtmNXZJSPztOBPdafpZzR1U/Bd
j8+QkaA5ERKgxljfGr7cXDgIs5x/b0CEfTtfjkNK4zsH331sLI6+X05oGDctMdSUiTUZYsZz6VnC
9tMVjhdra4594qTUHC19Bhr12H/LUobG+8LYKBmvB2EuF2KncHzWLBOiksHFZUSOrbWw3F0qxinb
r5wZpNCYjIzbiWOewDcnyYqhO0HMEQeNGaTCsTBlsSQ6VH6FlWYG25w8OIVvZZ82KvHwvW1MeozU
SkckgtgpvhFoDbiXmwcWaBb2VZaDbX9TDYyXe4qeCELjznBf13NY3h8yKRudPgLriPE9VZMYRKLZ
PCwEqF58plgjfNe4I7i70UzYvj1osO+CPszlCYeauib5YX7C5UQHfF/CIf749u5AtpKsoZzm4wnS
IYTw9H9eDvF1dt3qru57JoyQI0819DCnotJE2YR9WvzHht8BIQ5nNbNnfnU+aPxQxo35LTQzCtUC
TeeIPXc0hjXHhnEIcQRfvhtb+zBGdk922FlsoCrL3Vx5eD73dphJvPltfCyMdEL9Ph9rz/z6Qbgn
VMPQLl8bYVqaRXtkqLl02SWmozisCL6ueyv0uhRFFexV/YRyfvsZkVZPS+TZqnACgsypppAmn7Vl
2yexQuoiHi/zreCzLMT1IFq19iykuw4DUxclppTrI559UlSxtHOuVgJhFyZ+atgxZAnBalmeyJgj
z9N8NVR/tyFTTq+lU+hwmAz+u/N6j0oB+U9HR4erYcVA9acgVGvR31m1D7zw0izMH5AX1SNOnDSP
REt2dQZJTQhmbO7KQ8vORl+Js7z7WaPA849M32MMoLSH+d4gxqEMIEVHkvbZ2uzaNk8z0sTm+Kwi
oAqTZkeCP2uhFbMV759W22/4c4CillAXTsjAIFg2OSLix3xCJuRw4P908MPU3r85puTqfFjev0Wj
MYrRMXxeGcIcnBhyK7p5qk5HOYL5FeqInChif/jrQ7ueNSdDoTiYh/3VPa8KAM75PzAapoLM8vRL
hLw8OfJx2RpodZFCn3SquAIq8817WsBSekQaEzE7YHLrEZ6kusv9DpFx6wPPaNegUi4gMo3em1VL
eYexdPaDiwqNcWKbcIvSs0aO3bsi1qUnOd3kG3WzmfVt2LZJ+5pbP8pBeEV4+JK12aueOt9RwKPp
FyiZDkgwxXPh9KQNREy1Z4eUE0HuTxug6FuRycei1/7kMUQrV9qeG1Z9Ek5q2KXW8g0jQ5bO5t2G
rSEc2khn9y0NpnMwZNfcgtUZ+ELVB/sFG0OeGAeipxClZjOhd2YeE3O4jm8CxOlqn++bTpCuyot8
kYzXyPz+psT9S09ihJW5HXZdjTwWZJ/8cUHyQJ0itU4+PHqnBfLjBHaKdJP+t8E4gRsmRox/rPbz
IL6C69sZtUyFQavQ+RXBZ/iLoVRBWOppppZuqByPzDyrolJd8tRwSZ5ZJhPwmBnbZzjxqqDAZ3WQ
kVYXwfJabWDhpdaRbA7mP7mtgbNjd5ZGZvNtrLqj077mi2pDkpozWd/lfz8nRmSbh4niqvOCxTOL
9z+qw+FIC6Eh8CooCzDrPr8422A+2vYVpV/FCqg/VRi/9hm6nCUSUpGvHe02dbJgX3z4yQ3t6kHm
/B0cLtxwRhqk0BnLyiNHZLMmEpWzK0zCLGZqCzWxlNT1YN/wKZm8IGNfXvKN/3A3rjmTD+klGy/F
9rwFteHiXFAnnMZSCx1evQ0mYtw+Pg37Qd8zGm5PpsQt743orHRvUFtj/hT576Cqe9P/VoMl6wsj
AMtAOF+Hbpr33QlaPuwnQ9B6ZlckpWP+njY+oXf/ie344fDY6vi3y7aR8/FqVTvVM57aIaSsB+Xy
SJI8PZX4pJMFLURsVWNsjIs7JIiVJU7FPK6HQipXAZDWfiiC+ynHaSkZom87DgVcWcUIshn+rgJa
8RhoEFU5CxNdeWPhd7b7KfajfNOHTzlqXzN1Mvcp5br+kzon/hPxXKYH2eu/2inI0wZCClswF0Ml
UWmHMo80U5ut6OgJLilrzkxJR5o9etGTXII0cCO+Gu9dtiz/M8q2YX8VffaJRGrVxqEUpS3YGoRu
ILjhfjrtFLefiYrXL2ja0c5k8aNii0bXVRtkZZCu/Ba616fhHGnz1J2a1BW7+RPBOYylRQPgP5ri
eJXgfqoW7WtiTXt6l1aIS8w3fB+neTP3yuV3hwMO+ErLJt6MbTBT3efQVyBtFxgu2Q5Ze56EUfDj
wZpWjhdlhlGgxQQPW4UMa1k2eW1rA+vCdaaKFC/KL9DNzDc0A9TO7ND776SduiqUNarl5dwgVt/k
v8k/Bh43gI0jy1CUiECariVmtJC/YPA7vWYHnckGYW3/z7fGmVPuEUMJr9rMqVpRuuhg7llzw2P5
9GkyoNn8qwDC5HlBKVAxMtyD3u+KuppEH4RDydqNZYhbQzJrRlM8q8TPY/VD0gvI7xFYBsxJiB5Z
F9kc6fB+0z0zDs/Kjc7myyq67C23vwsi/kS+47VKNosQaVZQMFkVxcD61VZ1zCq6OgEQIeYBjv40
62nYK7+8GDJzmoMBOVpdTXkPvtPOFSNUBNUMQWrxgVdC8cpIdPXqAESd1D/lMOJg1uq1PNWDcdKN
iTTBy16IdzOWIY7haZmMwY2fkC93rgAnb69OedOzK1pco+3BSFQ1gO2yMfiR8x2NViw5GsYKU495
qkoO6BtEMSK6FG+LvwLxZtJwdC8JBei1PTdgUkv+p4Pa+AsbBatWQ07Jw1VLah16TlwwJhJfnGc6
VBGQP06z+bGiMbzvUa6rQCC2X6VteeS4QT+cII/UZJvtumvEXvV2qUPXm83q2ycO+Zj7lPHR/eox
dJu+W6z6H0f1SZSwCUnOrZtO0ssHlFF6PlrwUQJ7tEheWnONcpLcEN1DuuVgGv9hgHUWrXzyvW/X
Axr9+Lu5mcOfVmsjxA10bQw57iwqdO7OB0NxZDXqkH/pKcXESkZKIPv2CzJOUjmZriwkOnFPTQba
kROa1afsHycNtPIyVCak55A7Av9weVCZFH6wMDcCpwFkNwscxS7U9Bu2GXa4yah3FG6cJOgFYPxr
3S0LjR9qNG0erqtzbCY1t0k9p6q7r7l4aBWShiQsKG7bboyKx4M4eqaVwPdEEouWtIk4Q1PLzbyR
ZBRBaCi6uww3tGhT6PRpaB9IBlWH1sTmku6qrPcoq49brvp3L6JPTPjJTWNEAkxf5EIn0B6ZBJJH
h5P15Ug+DpfSPJw/fcwyKTXhSZLVbAZPpltN0MtnYUWItJng29xYTdQYowwv07uQRjNlmn4hQtHn
vrCOfzVFacejQNjNWtn9TGvvLHo0f5YPfXbEcwS7vvYKQEszypU+uiBdpg8NXkosEkezA3NKkF8Z
vNovxBZPD0QR3pbqVNpuIpbqtAsx5Cse9H50qVEDiBsfjJPn1GDozULCKOjPuiueLIvtfQpQ+3XE
foEEXgDPVmveOIob7NT6jVj0fW/k9u62sYEiYdaZkMN+cRLzj1LCJGSHjqqK8u4xb4zQpZpjhbNK
JD+u7Nqsz8rdw9/6yY0sP+t4bGGixT+YKdy+xr38szXo35ESVrRpcxhfxG9ShW+cYk27ahhHmwWx
vpar82RILFkKm4ptXSDrOIs40qb9D2e+NIcPilRqYkKVOTBEh+lDmFEyRqDPgYfD48Lhwud11Qwa
8ByQoC3Hk6F8jEFeKpBUGQCHe2s0VSh4pjHH/FSosffvv8QwpIEDfJRtp2LMBmPBtGm5yGXd+lrG
ZmijfcxsFrOUutfZYrhpIKVo7YmuxCJsMzwSC+CHfHsgegP9irxDnaC/Da/wcE+aZLBys5YsOJiU
wB1vtuGRfoXLCPjkvjKdXhxdiZhrh4OIXT0QdYiWD3gIAJrVrQKvXUkmivinMJyQkP8nLudnvSPc
E5pJvGk7aOUcfF8qKZteS7mLWfgYxjuj1BFqqVaD8f5uteGaf9vR+7Tuztiw0vHMcylc1561nna6
BAq6mig6VBzLsHLaob7SHrBpVM82+WL64b8XTBhySUxjjR13I45BmCmNCMhAtPmp4WfkqEMZLaxk
tYVY1bcaOXB26c5M+nXCpMJUWHpqCEyZTHYyHPXWMGayafStLQfol75T3GAhFn7yc2WmU/vU0eIi
CT+MUUOHDKd273fYcp2iyT+TLRjOlplbZUUCzq2NzU0ZMRvkhbQcM9cDngqG5YQudPk3V7jYySZz
7oqJKi3nIkzPP0Rb+KKVWailEoWIiZu/Y/O2uwt/HEKN+5ed9uQfb9A9zKT1IKZUNlHfU3TSYO1W
pA2TuY6yh+CfvipU/1eZ7q1OCrkiR+PeaaWs6ND1p7D+/HAMwv8g3GJa9VC/44vZAR5lAvvQS1N2
EKnT/vK1j4yAiElMCcMI6ZzKouj4MTJY2IBr1pbT+5BHtr7qtHczyV9Qv+SeHoLu6pAnPrX4uQvr
aFicTg7cmxDumznC9ZfPzatQr00HlERuVXA/gE5/8HFfTk58izlVUNlI8G/iIPefrlYzv/EwWOVR
jLwMcuTFUff7mq6vV2qQ2/KXnvIOwUoIVQVT5RNm/GK3kYaeBWlAYehVWKZAnoiopp58NX+tE1J8
lmKT7FzWtCIAIUGQIP1h7xpgUf0BN4VuEIc70mwTkxftZOa3waWJirY259Wn5YBQeC6zycTxv8+A
f4hpLrxEtuazncRra5WkyR2xtWl+iltsaQEUYfnJQbaIO1ZBpS8YPifjPF4TUs5Y3tCXjtT17f9c
RbDyEBy9jiR9g40A44WSooKLtLQe70Wx3OJJVOvhRKJlZPXaMrIoRlh/EsouqSXVfFeA8JA9fXuF
N6h7ONPv7NGaAvSYdWwj/PW/hXFUOBUz/8XbVUzi6Kc1xJlBGf6bKyk++yJ552xixVpOGZRBnjT+
hQEJyrq8i8RB+1FRmWlXKP7n3vJJ/uNxBI6NHEXItWOtwW2foQm2JeB/34gvlMFwXfxRjOjhahq/
qF/mIyJzIZH8sv0yCLeC2VnPCddB5EjdIDR1YIwtYmkzOF4nU6tvgn3KDv/b+kalKAzqDhRAVlA5
J7B+KELG0c9gLq7Zal7mFpI4fqRDUoQu6BfLxLRa0CLmKXkwwnJeB8I353LaLdQzidG70al9TDZm
Vtw0/OY2Nv0Az5Sr7u5Xf+owdAUQ0Nk4MGFu7R4fIS15pvguYrTBm61kW2KOe5Ix0fx5TUG3VqPX
P9YjNX7knVGyG3PoKuavsJ5GMpWjaOBfz96fCKQYmAeF0/S9QdnTTASaXc32RLr1ktAByX5nKsFB
LEYNYkmYAowxDs30fYN6diQxzpyM7SSto/OmKFlS0eco56NBJC6UXEtaY5Ka/QrKdeMPy/t7leWs
V+EsI/GAS6sAwBTQVqjAMu+ERR750cFo4uFZ+CuYWArwh0PA3wQCC58a5qDKrLuLkbocWGCbmvea
xJlqST75jGtqQRqjK8bV3Ii8NiPaU3AWUqrHHzMcWe4eq+jsEWFMfmY3w4oBLlDbjxqOukACpE0+
wgasEV1vMKwP5rOps8dkDD+YTcOjLvp/GtfntESbVNfU2xr6CCdRdDQOicgLWJx0zxT2e6Thy3Oy
9VFFg3b6mx2zWtENDsauI8X6724n6qC7wGNlCGt3TKAkxu/FCevDKc0IOMf+K0b4MGXMAKJpf/10
n67pqMiY03SNfaPb6JYOSC11NorJ1L9+GFqZJGruP4Y7Ly4XODtd068cjaVVHbVPp8WQu+6nMrnf
011oLUGcpNAgcR4zP5tUxUV2U9dynYl0yP7/xDVHxHsfa+PqRtb5vQmNETET+dR4QY/U6P61v4Ph
A8LcBjFIjKEObnofXh1fHh839SiQ9oI0J/Hs8yoipdE8odWHTdm1hmEIck+jKEWfQ63RCjffNnrz
Y83WwQlIHcbUxSMg76D03pBxfZPizYhYrahF7/1okg4C+yxSbhd27/E/u5wwPjeyGpOBns83IX1r
u9Qs4USRcUix8UsppTz52XfS18O9O/LBzbZh+g0fh0mNr+zzdUCQJAIg/r5YaH5jS2JQcPeGBX7B
lcUy7awNEFjEql7awsEihczGbzVF8jo58H4E3Iehv3Lp5t+oXlU+vPX1rr/XiUrUPQhLys1dsD50
LeRzzz1A0bCKY75pR/iFFQyAcclQuZrstBY3MfMe1NQMNouIVjzWShtrlmQye9zsAnH+vs1UACk4
Byl/oR+Kb1OaDYmrzFanfKBXXy+z2TqOv/v6B2FuCdKcuCOGpBCG/9mymuzXiSyBXliZVsF2q2LX
kYH/agO83pqwV0AMZu0XATwEat6/Hgoa6ALQqL47tGlVAvemSITcRgO8vldeYwgqVh10yB9+/vE1
GvS5d9VBndgXVdjXhkMORvrTwROcv9cZgOKbp4LNGwAEVpVjHP5I8ArqIvvmkufKDJkkkh9Ypw7p
fFQ3CSsQmczDW9S5lm2F3gB3VfoIUSMf3cmFuFzsIX9poOKprWgNwsTDTovxTTrna+NxfBcH1uLM
TjZE1R1+B6m8vgsQrTxZkD435KhTpbU66PzRxPqeJnCHx4/wnXFGOS8obbOBu3ZeuEHEKoRa978l
GoVVuDR6sl5vlMrAZLH8lG88cjcGIPipxf6sG4HQpjkopzilhZiSn8xqiuD1ACCTjWeJAWZJZBj1
AtH6EgJcybPPh6n1pGgOMoh56QQShn4Ut15BjU6slr7fL307UvCZJRMYSD03HXUK/NqKydMNzxxI
TjBc3qHkxhOrvBkg9jWO4STbVWOXxFE5ECClfMUK5/rIeXDj4dJ85phHf6ct98PSI5lyZiMbsX+Z
g8LOCtteY+V0ZrrAzWRvcqyeKSQ4bNwVk5J9j5UMUi7uC9P+f/WbZPPmedOzhsp8rBeTuoaP4QD9
igratdgfQQoZyMU8OJzpV1ZkEPiMFE81MFZCAEEVF4XA4mK60eJHoFAUnPFwaipthHjPRY+Lm4su
3Bs5y0yrj/e6mXrHWco3W5QiZ1TEHB+fzSEXz3tLq7Q2Nx+hrCn3KwDB/16+bmAyGuaSFEokDqxf
sehjsPQGY0x3PYXTD4XqC8cs08mBiNWYBhvRI+hvbTJDFHChQzCn2g4QEEmTO0TKbCHtmL/45P+1
SPNbH2jP8cVwPE5ySqFqVvCjz38x97GkFiQ9cl9nS5pijBvPJqeNtpr8LjG5YDcEhfDdem8MglBT
MQVfeA3WmPaWPQ7KQg+ZYADMQERcs868ckr1fXETUuN0yKSE5VHR1eSohSWxK81bm3MVhw1PiFA4
wipIqCE2yYIMb7pXrhl31BkySAiUPfuyOsywkLfiwQ3Ssu08zsoUzN8Y71Gn+UWF1ubgWtKiO31p
zYb7P3o4iPz/cT5egyC/MlcsTFN0LxKLBYG7tjbWJDefOrCc/aEA2TNEYXeA+UjHrUzAO6QslYmG
xSMTMdQn7GB2stKPtoc9hNSLxnGtheG8UNTg4ezb6Tp2eIUMyU6/tedK91KHp23J7EZRH8ZSA3rj
P9BR9QJO1kEM4jUrrwSNV/wxImg8NBDbeIq8G6+ZZcBHr9amdF5Y+6N4dCeH+MtTIXZyYRsrgZfQ
sJWHtDmLHqKO3MZtY3kxt7CKGPnIl2sEB5PjMGZGvQQE7dkhER/fKrWf+3y5p4ylPWYCH1sex1gB
aDoEWmbOjkswxrrM5PNx8dnoo9/J6BcSOEqLPhN6D1Zg/L04ouXrfL6eQvjUw65HDlvyfMKipRLh
Qtb9FFtjP8u/ibyRdokqlV7ahiEc7Z/0x7QvHA2WoL5ja1w505vWiPZ9LDC34a7RGfJO0H5v5N+J
Dtumu1t+azFVsOsctRXjMioOHuOm3s4bXTnuh0baYe8nqbVBLaPPrf2yeW7Pu1IuauuZ5u3VjM1S
UsbwBevtVbwfIK7IgTCr8t+q41uszHGr1PSZ4X8M2vVkB8n3tA+OlKmJ+frUqweasoTQRZRWMn6o
EUtm2oieuUf01tnV3O+8M8oZQd1B81TnIn7/aRZ16nQYKCTDYE7dcZNjOSHQ29JsPpLwXknJoJVo
I53R7oNk9Dh9ZY0miTazRwHqeYTKgDgh5iVSzW/Gde18jP+h+l1V1ACRhc+qYrOzDrODI67KfIA/
VNVvvRHPNyiKpkkfd1Ade3jkYGOlgTSfJBFfJPdW5c9WgevimAEigxRF4NXCe1r7KUW6V0cKo5Z0
Ru2dPHVl7s05cMUp9prs13zfsPYZe2HjCWXvh2XeUz0CmyzvfWxM3TUmv03xHTbVOe1NsYM9TBI4
z6Y6uBT48IeWrFPmC6lqWZhKlykUyg9dnIsCkx34aVEQUfr6ImsOL2letLKWVCgo88rTjLz777dX
R/FimLCHv33nKNVaA963Osz7XR//LQGRf3m1D+e2TQYIQRLTjimHOozkZN0mMrzPkyFvEVrIAzDH
6UPBG5ge8NQ4zXFoUjNs13d0Cd0jjVHVcs0Rvodhyi7qzCK/AST15RkGRsrR9a596Y7Hi9oMCD+u
xDuWQy1yLq5RsJqBgNpAxD1Yb47gifoNtL32bPzdeIn/QBXclhCm4azP8MPH9w3l71C4/zUaGvd4
8oHziZrS6b3lE2ZnuDZ1lsV9rBOiAsdBQfxiFSIjH7sBQb5MtgviS/j6agwbBf1rMVE2Poefoo+u
lGY8LWwyn4QuOLzxHNzGff4E+UN4zj9bTiDInVWjtsd1L+A8xILBsKVzdx31PP0TX3ycVeo3yUBM
PceW4VwV9HtkeF5vsHZ4V4bvEAvOo7uJ96q45PkFu13/Em/F5HoIysJm4WWKMehPXvATNV+N1Dlc
zqEMeZVemzTLQZqIRR2ZBK/kpOgLJZno9HEzr3dZxG5mDEm1JF3HRFsf9SaAte+Kgq5db8qgFrx0
mvvVok/7GlrSfud3Jl6/dm0fQBu75ZrEprF/T0jYT0HHsMw9S0ZyBv6W4L/XNaDFRoeG8bF1x/K5
a/TvPxk3N9HLATvkzXeNAlrmsgJC2kA2vnSLSZyEmjvpwSfKdqKMKhEcir8Jt/AjekWK75lBUrrM
rQ6Hl2A4DhhrtWGYC4TomFOjSIoRlyVRM9kzKrL/orCc+FjvMfTb/zUQx+iW6KXOdDMD1my1QaBW
Ufrbn/iCMK1HhFaHOQaJXtmmVRBiNBs94b2de4ny7nq3sSutlEoJayPuWcPQIJr/SJvZK9up2c62
xnRzQfYQtzFRysoO3WEhGzHcNNC1b36YJ+LJ8jkk/GX1m4bngoCD36TgSaN+PGy1oMDDlb/LQGKo
Cv7uHtOXVNWGd+f9Cr6I0A3QnoKmvG6MTXgOOqH5WlOXwjWW5Qskmt6TU+EUXYQdI40Midt71gNa
D/QA8BkHyHgoGukN1dORY0ZrKCZVp5bah35V5uPtjic0snuOojr7xjRxS/3xQ58yllXtEtvmHMp0
HZGezzUlELIMEEsae6Cjt99gtozB/98/92QTLIzeoNfn+xl8ZYtYxLsj6XgH3uTe9lKQcnnPcWpw
AMEdTf1Wi2+eqScn0gd2l5QRna377RTpCTzMAUc8T7/sGQFi1DBwN8SDqGjgTYbl/VzWDQm+eWg1
xtfFMlyQPzVq6gA82yqyQsO0m/Zz/C5Y9R6m424MtJxcrznj7B7hYXjSbua51V5QkR77384kxoKm
E7zbLmzSSbI9GmMIaED38qoMEBcYQSZEs+2W6VPJ/X0hmj/2PbSQ/DZjczVny9qOY2LatLEK5GGt
qMVAxt3jG5RMouwQnL2UrK8LGaVy22W+yt+9bi73lj9poh0+dbdOsIIjYXjlcl3xKHQ3cK7V25Ba
9Mi1FmJK2Fw7zlCMqTOoeL0whrR5DiqjtE3LBlYFlGS+l9tGTHr3YYu5dOvZUG4lOT5ZAyHiWG2Y
YPpZ2gxFJSMbqKSnOxkH7T6Ls53s6DKlR1eYt10m4iDJMoJ9k8LF09BF2ineIQ3Os+DnzhDmpDZl
gsLZv+2H7mFB/5PPW6UejYNwXq7iT979WyCar7dpx6E29R9m6q7qNkOx3MOk5bcpeTlsAZuhQYu2
ABckqSf6CWuG7uExjzy+wMenuw0Xjk6qFvLj31eX5+c6hBczdqKGMyR7BPeJ18+TGY+Z8bvI7tTZ
2rC4JGISZNRbmtb2Y4iuXQkeaTumHQKXLHnqc/YUnsj0PQh8lNFfvL3tu0uRrBYVb5A95lnhQU51
QBHeSTyFodNo3YNQl8nlZzBXOT1MmDJIFZ0n36yogebLt8bYeNW0KKTXcdmrMK9iVdSz0v2e+9vT
mf0LxU+S3jcvQ8OxY2ghj/S2MMyMxvNNIwEm/TwJilf+9INaE3YY+QNLh8KcTTRCjX7BN3dMKgTX
iGMxLbey3JD+iat04Imo9NGUqcnrO52Ees0C4BrJuuasDPXsbaA3EMZmJdY6tViWcNMzLeh//xVz
KvB6mIV3VWciz3B2CfZvx75rRQkEs2j5sMhiZqgGSQY6MpKHwBfBC+4sIaQsYBo+m9+kmcbXOLAS
Pw6cSCDM0Mzm6KIiQmSBVfpilG7byiZtrKBEKcBaQqz/nnlOiwwqfq0TB7L32ldsm93Bgmo8884O
E/XQOcGeS8P+JHswjraGXHQ0xFkqOqOrKTgWfPCCyaX5GANLObQ/gsFU2FBzjcyf6FxOHx9uMPwt
gLareYD0FdAoeYevgom7vfgVamcZqjOQ5UgdHsi0Zf0UYJ/vU2d6q/t1M+EtfgEmbKgoP19ZpUfO
SE9MNUzEqLjPrULr9gEEnR6uPtikujm9eRNgDbJbAClKiiSa+6boxfc2W2+hCaP/o9dktKkCxOCN
Wu+eK7XnnYf82bLQvRFWxyYVdENggXkjBLHkHaFy5kkSrj6XTTYVnoq9ZbIA0B0/BugFFcyRr099
Es8iAY4PmFsHpFziTJYGYADu3b6jy6W5yPqgsciBw+eldqFIrD+x5E6nNmRGcPDp+/94BZbGt5AH
D6wkpeZTeFx0Oaj1EGQupkzWWtS5AJV5LoLiTUobk6XA7W+UVBoWMP8k0vBDodOz/87LflKXFiMX
zkwWnV1fQO7XEBVniXdZlmJukDKhTOdCQoQ0UG0ebj7nxHzgwuiyi2FDkqaxAHkMz7cCJ0Gi/7I2
ye3/g12qwmt76OcWH2mgRJ3l5rbKNE46YhSvfg7aXWuyWcKZgDTOAX4/fse5e2ImXM1F1QchSaaj
DNd/ecVjZQGb+vOtZuvkZpSXDlCy2twDyj7kDeMN0oSQHbiprScYn+F9gQremacf+/A7KC8moDEm
b6iOxe9eNFLJ6zxSIn4xSK9NKvJ296TAvpQ+jF2OyWdaf/Lvp5ZaHeDzMzaLhu4sNKf+v68FgL7B
t5MAW9tfcH32yfyAP9Tg5lr7q7/fWWwZXVGSTDkdhjW9skc0WsP0k9QiifbTie8gQdjVo+2K80cv
4GTKRq3fhyWYUMmaMQbMO30jU9AG89cVENEXgd9THBQgRw2xqe3EuFIdpi7GBPeYETxGSYbdSUI8
ItqK88+FvGImifqhpzUBP10EPz8hqTQxdU7WNu31cLuRmuNqdxH3/AkJa3uBYJy6JrAcmnXSkREN
uyPHZkC1P43tecXQP+Ic40zblo54MG5zvaRkmIhS9shAiOIJ1Br+AJgLLmLO5PhPCFTaEvXnTzT1
gDepkpJNu1ap/WfVefeYRCsMoGSgZRiTy+HlR+Y4PpvwrOW2QaKmxQ2T9hNFTAl7BocMQU4qEpfS
5yMaZXdV7Wp2Wx3Sa5Ze/aE+GBJVLjwhAQ7qPqPR2O4/kigZuBrsrB0r8UtJ0RzXic4mdiuMw3y8
Ni3nvyix+cqG5sNFEck4wIMTpHJMzGYRcn+61xDcqF6rZK4MpV91dhiJCYty3lK7k6Q2+4kQzjON
C2VWg+HV1rb5c3o+aOmxYGL3yngo06ceAFRtJ8ycllC3Y9Y2D/Bf1+JS3b1GgvZNBBdi9t5H/Zg8
se/7CuCh+ulqqm+0N6e9prfmlhxGo76W6brmfKKkNSvclj2c9Ufpn3xYE7LgdCRoTyfrMeP8poMF
Azw8VNwBnLBqzSQQBlPjNRHAEs6K8sB8Hu2xFpkLzXpeo5JleD1YyGZWcCeeXjF7Pcdg9FMHufJM
bJigyTHz5kMb4yW37go/HaMe4QfG+fcdCplpJJE8lGAv6RvaCQK/vzOrlPEAIb/AxGJv4xajKevj
AA3aab510RDf3VeH/VB6Mjg3O/QjOIhEqPS1Vz0kYH9AcRaT6UJWfYkTPX1MleTKYhnxKDXlmGmT
qTLbRKy6zPc6nOR9xMbbvGT8qDo1yUdxbURVvgo7kwTBN6+S9KNgtj44e6WPeGvJ1HK3FvP8wJAK
11zFRwE3chU253nC1BrWC2zpV3UmTe4op3wgdqVNbzl61i0cbgcj5Q0MICKhvAWEhyuEhff1A1ll
qDc8w6cQPnd5o7wVz4EOPH5M2Apjjzozb6mzqLBcngmSn6kPLOrJ+d53YJcHZTGpZtMneH9U5tZP
Ugg3M0Jfb8reJMYHzid2XqEeYaNEbe2sC9d4Ji2AODX7x4B4+BO9Bbd4xiVOhxAQO6cd61oph6Z+
zTXMRt+G4tx1+826EaPJcNdcIFcYUe8vuSQly4IkZoL9kplGIRDQ11jlSE/3soGmiqz8fu8WLZ/p
nc2WOQ5wECDtEWDyAcaHue2TSIfxixpo3yLuWwBp8p3vyC+DUVDPLNO94crmgaqAuZGiUnPUoXNV
hmTxihpCdUIc1DQvmWhnsdnZmBJ0bmpSP4N11x8N5iD0NMhvqM83yQyayQURI0LPIL7YGDPWp5wo
8z8cpDXCX1iSkObf7mJnmI3f+WiSdzEnlAKcizHYNl2SeNf8tPhhPa2pO9Fr1+wtsKtY3NDIrJp9
RoXJYY8jdH9P8z4hctmFDIGL09bgoyfyQ0LLXFXl/OkWydvntLMqo4wyXsVSK9ozvdnwSXuvrK1Y
sJo1aWvOA8RswCGu2Qw5sQ/errj6kGxissJpj6we30OoXIh+XKeN+bVcgz9K31lm2kx6mv5VZlvc
wtiN8KCXxBMNAsgL65WIX+LpnDlwqTJm/ssLc1suKieICQKGlN8Y9Fe0hzs1eMjBJ1xcgdQCqB5c
yBOwBFMs0L+dshX/UzaOIm0dJPlLzxP4ANNp6cDMKRJR9+ugA212SaFUOnpDR2fjTC4PKTZfcuGd
+JI95T8HteJrvbzaer3JOE0WKRt6GMrDpHLcPSVILPSaleYyxKaE1bZBoxMTD3yGYtoF9cpGNAip
fm8xJxK3ZY5uqxwy/RP27ul8DvkgmSqlCFjCZSJ0RqXFvzBW/EC5KUu3hcKTN593EDSikDAYv0xx
KhZl2hpVicUtT5IQ/fPxttz1XKZkROxWE6Ns/HLRCHxolXZ1W4Jiijd5usoRB5Jq7h8TN5QY5RZ+
uCOA2iwsEtthofr/vMsLyYNrFs19DOVHe+oR2bhAkWJxUTDDhWxfa/uVEm/8dPqA/tx+imJxpwNl
I8/X9qBxvs4ZXDS4BCIG7tluSCGiLGPxggkOvwMH/smT+XCEbqF5FXzM//OAArTLign9Fyq/Vr1Y
+Q1nth1VWEwRc/7+e6WJgq0vL+J/gK8GqiRFnoV9W19gvGnfCjyB3aGiWYXBnFlzR/KC++GRdLFP
1q7MAZorBqnJkNjEQc996tXQlknMunAn+dojh2WZAVGUV1+pU6XsDLiErX87TVC2CdjZXzfk2+n/
s0fZL/Mzm74b3HER/JGjcQuSf4Nk5aBO4VGJstODZJG0kLU8Y22w33SrwAphaCi7MvTKuHMsCtta
UUX2ENDWPQM6T+c5ob5pUmjPhF+msAt5qqgeegLx0qp8Cr0Ln0pBBPwvrTw0us2dbVeHzjF86HbX
j99T+GQQm6X2Hvr9dgkgenUG7nkWlhPoomsMbVxWi4Brl45+EI3+2gTubRFfpelI+IrTzVLBwFOl
k7dcE9VFxhPryudl1UBAAJWbIbs0HqUj2FE8R8Wbdynu4Rhhr81idUFuyeWZmml5uHOA6ufNpa4a
VNdnxiqiUO1nxQ3HKZX+SPV3bfIP4q2UaZ/IF8C58rtcS1avVdBGxPo0AoYqUXgGbFQnj5E/PrSS
a9UM3LFdxmWrUb2U+Dd2LFltcfoShRYH+hDupmEX+gsqy0UL4/zvO9JzturTAdGVvfahsU7dWSWQ
iSDRrEzA0ePZdwk/VNEMWoWlWEzBdEts6AISl8Q4KhC39U6imnnL2y88GSbxhQhnKHM1cWiEBHEL
hwmtKz7qRDl5ngZ8oX2lh+rTYoGjYAG5IHU6NUiLunmY1c05p94qXplmIjRPt1ODsmnS/WuFjtmc
O9S7YwQcAzNOy1UUfaT39XIjybAlr+graxBQJxiST9liV18J9UMPXtIP8uVbJ1xHMkDESIPTv4VG
KgP4yCTKzL/2G4WR8NrJH2bDaEexb1Bu2FgypUAV6oGBxslQDfSnUl9PAth8UeBKeaaCaIysqAmv
lGDm8uBe31N2XaZo7PATJP7Wd2OXqhWOMv09eEBbUSuKPvcU6dixQftOoRD6BOBm8vXp4FChdxYb
riV4HgyDcmqewkR30pa6spjxpRskv4qSvJHxMumlYa9oenbAfdeZTsPsEGns/5lNrilHVBn4aK/9
/eAa6j49MFygDSu/X/ZD3rdvlsgNwGvlUzJ5KDpccRgS30c4XImvsNOAoLH33Ilfd36m+r/I4NXR
U4Br9pVi6ybuiWMxjzM9ByHFY9QMW/8ZBfFBtcPRmc2eBr5pV/L3NWhejdomFfF041V4JU+R8Xm2
lcIPTLt2Gkg3ccVEdEW7SZTjynU4X4C/NWaj4n5+IrsNkXmLcAGSBRWz3KXKVthUqP2YS1aiIK63
lP9qooKynO9dovxy85bNOh6b1b1w0WD8nF/Xs1laGeHN25WYx/5zru0/OLvPTHOzQ+/W0FZqOoo+
JdwCJLrKE/3JaAF/qa23HgzN3UQngPBAMJKfFihtSQcEH/P8Yy3EsIYSPJwjrfmrcWNQ+fSOEx3v
YE0n8+0xyEAxC+8WDhrC382FXH5/KAH9W+VC+4P9LJds5uykI8KcnBw9nYGQ7YtKXvCPvYwUnu43
JUUFYCj/ti00tZ3u1nfT8DDk+UDeZJcE6sUawqefLQnTkFfy4W5wV3gyUnWfHG3GVnpIcU5WMoWz
TTa2LOwo8bNt88Fj6B+cEatoqhAdlZCJOjty7v9a+QEjTeQWLYjNh8jaITj+E6UkPipySLNUo06T
mNdZHtagypIoQbtsojEk+Wx/K+SCqYExASUlhxMVgp3l4gJvYVlb/Mh7apV5rtaZaU4PLe9SZsTC
GNws51zrhqUYulOmGEkx55VEmulclq4pzRoM+sTWvYS0oLJDgnulTxIjYVt4VLjoVJkSMGqyXGAF
JGb4OW89ObqN4TwuZhTEKhKCt/K1UsyoAimTQpJgpG/rhJlh1WZ7RbTDi67nnw9AQiVc6CxvfB9/
035KzmoORcyQZ2YO2w/WwZK/ZJL81dlaUm7bGIu85ExTvccP70Ji0X5+3OGFU5WQdKJZDx+LshfL
znlsXnHtI/NoCCJtjl1vECXRBchEwmBDGa99ErY+kZnZ6fcQYGJjhSpBmL/BIx3fFk5evE7HAbus
sJzTHn7+68GfSbFuxEw0jyrIc4Pd5AG3jgzAJD929a7DcIn8XDcPpXd0YqbvxkgM4z/iwqY0H7l8
Qslpsz65NoTZnGRhXuTK2xseYNFEN8ISR6XaGjqhGkDpZ99iVKnY/S1nlxVIxu46TCDZmZ6MFb2i
G/4bS34QGgqkUeDDn0b1PBwkoh9CdFsint/PdlfBgvRIi5wv16jaS7YLn/Td7KK5GU6hY4RqsSBw
ei6FCTFHbOb2FP+DAtcxxrreDnVfUmlqfuiuFe3aCOd66VEfYB9NS4LU2hK3EBCE4USKAx9GHmG0
QRbG88ZUv62EU7Uae/RUz054WBE5fNYcNp5vHsBgsThImHeQdPha7fszWInX6Jj87wbhuIH/r14q
99GWpVh8hTSkKpgOVqDP5GxV2UkvcRFm4T7NctTvQuHK+Q+s1KuLHAD0WUtUE7koDy/zkLH0CskQ
BR3PQ2FaIpYJHWzw40qqlH0R7JvLB5d7UYlBJvc53tPo8ae81tIeCtok+DccJ3lt9284oJjT0BA1
aEX1AOnz/adPVvgnqYZtTNjJHI6VEPBF7Sq/cHT+mG37u9Wbf5gyUYOYAIJPrI8yQCQFhaspxorG
XmEKiRTLA4oWSzmVtz4fXNyBQR83ORB4g34N94SvwzWWsOGRcCECpi5CcwxZdmCDUT+HcDksXTz5
GpQhqXCTwjlr/qKp6NgMJQMvyqEUZ36swLDs/Ew+A4B6ooTHre2YL30e4n019XmPxMDfHTBbQhzT
18kW9aaVQg1I4ZYL44eKdW6BJfusXxf57iyop5VrXI34QztaYVjhBVaFQrZ2vwjEvQ4STje+17+D
khQNsMKlHud4PbCfQNue+CdRqfRb9K4b8aD+4Hyx+CUX81TtDrIUkjIWHBfFKWoKifnh+6xAChhW
NgPCOXBwFb/AQ7YFeFVhuMNiYrxMGaGwkyl3IcnGGykEWSLDpBBRhtunVW3S8JqZ/zkJuly/C2WQ
L5L3JjtgdZUCWww2xavEd7dDyWcY0bpU6cl1VyZ24//k2X6ZhMOIb+sz1gzL3ngGJW1o5jArvNlP
emr2jI47L2mCIbomXo0xxeM9tPNWk621u40pC2h3uQplDLdr5RmXC0+PCrF96c9VSUzlnKs2nyJN
KEWYWHX2xI7rR8q1NwnPiLPdLUpCJWd3a1f0zK3s/cfRq/ZWPw1j+UxRySsUjyX2KgIAHaXtjyiE
TjNPl4Ew8r68Pd/A3dL8am/mI2N7SbOf1SsCyzJbAPiJLkaIpc73ittcUYjSmNazWGip18w18o82
ByzzJ0sULWZKHo7eD0xfUYcXDcqk5GmJEpI5/WiJYWJCpWZbuAg1uUyNvKTVQGOzJ41u/QjA4K3b
LzUsVXekVU8qVvtniWoey+SfziqiTJsk6VL0i6GeugW0Hed0cfGsZok8BSk5gULOp5ZGzbE0O3g5
5+e29rlAyRwLhv4NWWxRFVHAUGX6tE9C6xhKCdX71Pk4dRLN3lIF0JLo+/ftAdrk1X5UljGKXSzv
a9S9BoGd4Dk6X37UTprfL6LNEyb2oCwarwmB/qWKpQkQnlodnzi+4HmQosnY9tmTlVod1HWZX3ba
uv6Y5xWKW47wlfzR+M7Kd3AzPSIbu3ik7/8VYerMKbF1vZ3B6O3jxcYEwiiEtGB87FGS+NhP8bNy
NVXXAFYi8U5WmHSylibK0HBN5nL9y+tNS9srqY7dQbdlp9oh/WbggxybULN4WFyVDJIoZ5qjXjxr
U1RxHl+TF5445v6mMWCIvcUS1++bBnsVPIDiiTWvbCENJARcntOMYQRT3oaUJutO1NZJWNJqUQzs
2uHGQBmibi+R0s8QzAqFL6BUa5o8Y5OZcZ5PMfqg7Xhext6qlz6rQJY2h+RLNyutS17dWiJxpWeX
G4QMSaiBHMZewzNHRkdhQW+kOEH+qM2DC5mq/VwOLyZytFv9HetlZTX4NZAQVQBw3nylJVyT6OPy
19+aICmQ5LY8uuNkz4YKnrPkyzr/FfZWEIZht4sfAnk6ugB9FP0mYx1P5kg9hwQ2RzUlHU7OHYN9
ZNirN33nkkmtgx9nSxgsk+F2oDsQiz0NY9WnWsCRF6K40SvxjILRxz1EMQTdOVlMndBR6gszzF2u
vIYwRfH6xXGk42D9rpxGJ82WjXy1gvk9LTZAY4NoLOS9cqxPMV8Dgx1X+IAIbUjmCrx8Yn5fFtOQ
02K+S/IEMISv6vNPH5OXT2LJmTLI+uuFMU2/Z1AetQYVaehoMM1dBHN9E0mML89ZdUD5V/DMpY/V
h6HaVG1zqh6lMKXqEsjCYypjq3RGfrX6OJH+/IEYI0RcrP6CmqRShCN6BYzbiK8cJxX77fm3QYGU
TRONZ33Qru+6Oj/RgeGE0VfHfgERe1ZxpoqdWAnxK9+2jgyN5jsaRPiYp45pHzsus7AV0FyNAaO+
96k7G4WABqYcOunN2+0LhnBifQMPS5MJfdOywoi5WuIY0kCvQ9zgbHXXA9C7By6ly83rep5acVLP
t/fnweAKdq7HtAds8Jjw3QvyOJKcVs3zgi4Yo8P7hzVDalpkkBP8V+5584ASDJ1o4Zi70DpyOl+t
rBSA3juxJRHkQZRrCDLbYNfpfbRQezO1od5NkJNB1U9Fa4ms2hhu2x/aVBlqlpRkwqxws6pn9vj1
SJGWrT/NWzSmPBDvvGZPwTVjGKwq1wVvwkkJRcsO5nDmRdjJ2WZw7xY4Z15vFXzu7zb+ubaczPMK
M8py/i+pP3b9umh16dahlJIOovQWt4Pehpd0bAaeIS8W45eU0pQG6cO97mduEnKp8elVzbDHopwZ
P3RRjYy8uH4ajSdhbBMTnnBZmsaLNp9boPTq6gPFPGTcI4sj0fBnOTNKKSo15DOoNBBEgTOyR1tS
hXHtBX8KQCa5KX0KhnY9VN455K6RknPVTK269VDOzThumoVYEs15S2WrTrMzE0gWDYJ/AKf0f/G4
uQTKFGWHSY0ecCpwBGK+cRr5fGDv27vzlXR7dtC4sy2o+zwLwqfwZNNmhE5vnf6+81VCvSOwkZo0
/UbL1zSiyKKbkkrSd4sNulxz8knlsn0sPZmGdNSgE7bQOw7KMtBt2WRxDcsCh0VploOqv5oOoKBo
WqcY8ncyEeV3ZNKgiWq+o0ElRpxPZoIvppSB85F7Qgq2fIlrR3DJ+4wTWMOS7QJLVFRQUc+WHmQf
X0rYqzXDZ8pXRjF5DCuARwExLA6pJhoHrqXFYz/vvNPg9Areli01397/PQwfnuvNvLWr9T3+g670
NnK9YDwG4xIVWAOoCxGxXVyxNYOR/wrnNPjGR+ePUuebDO77BlvX/gOZ7iHHg4V9+hfa+lBFg1Fa
CGNu3R2QI+hlnI9qPHw26u7zp9xZkZNaGNPQxjPbhj3K9aTS6vgWMsR4rUNaImjzuyHpQJHqCq93
NW1iTcl7PVnqRBlxrcexnDweZXnC25Zhge8c9oBKVyNh4wWu/byQLUxdpsLj1B+SDE0ao969XpTA
fZezHpgwUqRkwh3/nq6XoCFZmXhaqmMEjfk+l8xolkUjmh1MkxdGNfHCq+IPwTvD83+rYC+t4uBK
4JDGpwUwOISeL4bg0qxGfM9yyHZy9dtObZGpzuw77uM0Hol8ngLGHqgLkN9uTqNZIvHJvj43/X+D
mslbB0LwY8kpZVilfuBZqEFfVyQ8G0qeUYvfiXCYw4G37i7+5UzGBaCiBPYPc5k9YKGptNr3mM0O
Ya1UTImPc860pzrRRDbm40CBGm/MLCahVATa8//plaP8hm1MQE9j4RrJq158+KGHG69CvtZONdC8
1Qz+0BePr6ZdTke7XFdfM4m/3K8eMOpyrvjBkq6zMdS6VADn0b/tJaICYrDEoRf/S4p9f4ufXGVw
wJNiOJeb3LFEL2xwKIVswu6BVKpMjPgZlv3Owx/EE8fSqueoveec2NvKcbRE7o3kqNQ21PI3voE+
8WKWwnYwhvsRL4OlzfcPMjDUtrGVLlvXhQqMuqftldNQz45VbQj+yPvHjqdQOf6UR4L+JoCvhdHI
hccQ61vTK3RVN4XUz/qMOQpJTGfQT5G+wopP7KZkIHbvFDpusLgzt8jHO+QMld6z0buyOw6LqQe8
JUYr0lMdTEC+wk1GSHJnu+ZYMMoP0E8fT5XeysXy5s8i/WDxi05054c9AAGbW1vXUjfYY2frMqYb
qekMZsTxjvPi1Kh9LM8rsf4FHLRXlc6yKxbJ2UBWOqhY1E1WMj2ohbt/OrDIRri1Zf1VuKhoIt88
Rc/GRd4U7q02uthpTFQRS0CozeEZYFLbYJiV6zeZipsyyvX37/+/+J4n3SFBppjmaUkyKo0NCiEE
O1NcFUWrtuNibpoLx58MUJI+yM4M3VQqyCo3UKHZfLAAAv4uT37n1F7XQWIj/YqrjTWD4ZyjNvVR
oG99a5lOY5keVONeUqpST7btd2e/NBSz+okGO23MKE1M5pz3JGHKSYOqvsKz7O81LtYRSgUzPFNG
x0U/q2ZDvp2I5ooCelgkfH5I7tviNBdwTgnKJtfQjMwrhwZnxC9bVmJOSZt6Pb3wuJsVJX7qbFmO
Ck/EhFsHfzg2v5zP2rCS8dfcfj6hbT+IPU4i/cWDjBY3e4jaKjCF0IB1fl86vrc+MTKfvp3GXVaG
ZCJ2sbTuT9aKDSqYeNqJMD59ip4ii/O/N+gTacTtMA/a6ybFhAyLJoxDonOlsBLweIQjNhlpQjCJ
KfY0/pCBOZTfQrIygroO9RGQxHBlNuVH39mORizimAhi624eWfFqpYvuJ/57RMwFHgihfKZS/+os
NkZ+FBnjMDHDpneAwz2F+qRULQKsTGVGlukFQ2n+LAhOJD9Lob4L3H2BC/p7lWUD9hYvZ6CDzSlb
N5/G9oX1UupFtOWqTx5h9WmXUcLaTFDSG1Ojffi696uVIEzbQBXAxZrsGWS8LEbw5oc8RYJe9hzU
+3jkrw3ECV56EMhn2g9DYeZFqfUPMr+vMmATXVAoowbdhNpDYGP6hJN6FFS0fLfQ5liAkzZpRIw7
N14fYln7Uyv8i8xoWOtnHvpRG6nsrTAw2c0P/W4thhoKDbUUEH43sNVDutltoN2YolH/aAjVYx7v
qaaMnyzCfKRYKzAWVwGlcG2d8ijHV7U3f1kLF2t7e13JnU8AffYniJBvfLD2t4VClXoon0tNxYVJ
LggVx8K1Wdevha4NndMKVwrcHRafL3fQdBhX8+3DrMUZehXJ1HrnqoBuumgxHcEDAboe411niRPf
7kEPmsFiZX+WzCQKHYLt8o/g4HAcksFGqnwSGxKYeQb703wzyg1Uekr0IKBoQ3BzLVFePTnpswfu
tfYhlDK1lEQ24vo74Q+y7/v04odj+WFi9C8BoJkcDPsP/6DrfNmZm7yq3F3R63DiCv2cf+95MGn2
0e7tqYscJDX799o6MLTSfH7JFvz0wqsdG7q+SCFHGm95mdUMunV6pR7SC/evuNX4zGXxKBpH7nyv
xIppqRBvQMfVYiwe1yExogm/inWvYbRQ9GImMBS7LBQQcHSwYJWnzDCtWDAk2a+YCloHi4wsioX7
ZczyQlCs2VdpyhvePy85nSxmHrMk7FffRqWnmvFEdCsyn4DZmgnfWvxt5+wRvZRuW1V/ZCJTW5km
qUPTaoCtEDNIwbgJvCKZvGxreSKZO3xBD0BPTFKNkSudgpLMhSfTGpYyBdwcq/yLRXzyI+95gx9h
9qdIDzfDZBIgJD+xV9TG9UKgTtNh8PnBybsitCk0iZt5cCZ3ZMMvTLFHYwp+ObOp1af6LoRRGj+u
wcMvCfzgTu4ngxzJ91gL62Bl1qWkasroh5dCGWSPbmUu4anClvZeO4SEcv4LV3UBLU/lRZobnkB9
0qPnAfmR39YIYwasSPXDfEJ57KYyZQ361Q366//BNwkpIzNHnJ5qsW24/epH9VsqrQ9zL2r/cWKq
NPjOiHzEgUEt2LpMiTzGt9RgKdVMWNsduPyaNGpHZoHBRXvQNuLWWXmm5ZWEk3ZisbZQbxfzyAu2
vpvbKtxSVVjYnShS3W+Qw9coR3Gt3kGAScdW3W9jUYZhfgzQqELGNw4Ad1d8eZE7wQjG9ZeHPgNa
S7kYbPYjdh7aTzLNrW7fr9ctct/fnqIexJVoNPys9fSTZQ9USZIu3x6aXUuo5PDDfCR+w3pXAD9J
q+iIVrVyZORdXUNppQLnUMWLYc38EcFBUda7fE44th68witbCFBu4svsbn7Z8DsobbOZatnsQm18
ipBik6FQxPFIqm36thmWj0y4C4D082ZmAq3Yu/tjE9BkLvNxvcVV8Ylb+m1CdfPTzXQeuLj9bVMB
ZaTzwpoq+BRKiwqKWKN+y8udEELgLRs5GlFHy0HfeNszqHpevKmW4zlVjpHCT87SS44wleYpAZOc
7f5jsXpzDTbpS75T9VDHjFsaYA5ka2nMxmrj2pAPPaOwC57PV0PFJZAegAFpHBqNraVF6SWPjeZz
3iCSIwp0e920LEb/c6ulakOQeHucO42EH51TDqnartN38JRrcqJD7CqtzfR5mnQCp2N3OmGkHRfO
mgWh40BVnIX1e6X6AY0qvkR0Hqgyh2/3cMhrys/d7qnt9SfmO8/XI6JwDVnloTTVy4dXqFNwXGhR
Y/etMl5nqwP36ql8/cRIwSNUfHiHKOZygvIbch2BmYe/u9qlhQ9S9C3LCkuIPcH/52mn5Ic+B7qs
XcTTFkZYx0A0QvnhMdNDSvzIgD2KLR3zrQOPEneYSvOciwnrrlP8YKZXEu7OdQtiJY7/xWruBlbp
IUOWmS5TlMBKHaxcIfyt75/o0+iEdaREUmISD5OMJhRuaffqyknYtHA1Lh7jdy/8I7NXcHaQVbLW
qoicPt9OqvhKj5LVtpF4IE/lO+uBQPEtDjQbIxBXWNQ29iL8IwH0su8OJ0/NzzRKD2o6vDnyBlVA
YWD4JXqzaubHfl/BMMscbE1/RrjA5mnAjVNkdbGwBhJ1Yqim7b1XJkeAlP2xXS/WwWvl9JIlC4tY
9iepssnG6ar48eR6ElJNAVakrMoItptooe3W4P7Yz0NSf0QOMy3sNBy7hlMGYATdlH4VjZ31QB5R
Jk7ZZOe0/f5jdkzN8vSoaCJv5Bo2LtLmu/UeKpq5ibVNh64cJIorcrelgQAJciRnHTqFCUuUzMx3
QmTEoeg7Q1akWVa9t0KBvvhTJ3jOS3prDBOOE3KVzoSjoOBab15DhRbp+pBL7TqJUgR4q2jne9uY
4jgu5rEuxuQx7KyL37B53YGJsawZ9oooyHCbqBNnW0K4LAIudFjkaxTSwvdfcA+6mw9/+YZx3z79
jsWehsC0McnuyKhXyKHL/Wb2/HsafXTlo1qpZ3pbYFs6nkwD6pORK9N2eMImUG/+cFsRYTDlAiat
zAATAC1zB0+QkyyF7hdGEErfM0rpuwd80sNdrIolRgRjWEqtpg1NtyPhICNfEao+uDH6DQ8cc/EW
4vr382AyDKHNOv/QtIygsANbrHVAXo8UpXlOndsFpVjXHteJBIBMAWKUiF9N3pjYLDlVyrVGQ57R
dzYtgWauzWhs4h6zwPogpu0hojvPPE/kjGfrZ1nDtoUh4dFiEX0x7/sNpOf16fBu3NXiruKh6nhA
PZG26pIPEdcqPNWM8CeMTpqDUlssMIz55EcqOs3yqfZWNCARjb3ysZt7O098OBkJ4sZKX2Rd4Yok
s/6LQXdumYuV61xx0xJlDHBSilVVSpjHU9RHdOWO3Ot1tJXfKo62a5mOyGxWEKisVyErFjWHXYaY
7l0/89NPOXy2TBotoHccuGKBzxVC5mfjoi6mMphXE0p4dU/kSY230b5i+I7BrKSG2D9nGiZxwmOi
6XEzJtcRIjr7Mi0CdlEKpzk2bnjbYLaBkqlWwH6Hvgy1g/bUhE45JgWiP3rVPN1ZG3Tx3uTkz+3h
qNvp6UWd0ZZQA5NOSJaP4xQu7WFD30F1qVqTTWEgNXalT1gQMM0EzfVM+BnU9L+lZKbJBdVo7g/d
vvgflZSlKqKzgBB4eCXr+/3RAxQmLR9xBTG1jwME05RsRhCoHrFenW5Qf/7T1OOB/tvjYokUBj8d
tmGac+zQSfaJNjCjSwrll1rxuHMVrODw8BLhbhGozcXvNS/9QQYkYd1Vd2ngqSTuDO/vcj6Ba1+8
ja+4kls3MNQULVDCmHNgKpQ4mT/B1YTDxgb738WNgarOby9ee8O3N0QHSM2cXqgWjyIJtn+pc+eE
ht6G/HSYzZ5NTX98l8fxVXdwOZb3MWcOGzDf5f+RrbdJ2w10Df1TU+/AlEyHXE9DMcBkb6QIxh4/
br79MNTe9DLbMp1HcgkwaL/H8LnYuV4vtSarf4jUfgFCj94k63tIh9fsr2PHVMTPo9x3TQ857qwP
fXtzCxyyhRG34xAvVevJYsNPn56fv/3zniqh4sAjrVMYIDZrstSemFhqUXX3IU5ma1YzaYtN4OST
Nd4xkJuDxeQY96i/V131jS5iXSKyuZ3eia4jCKltyDonf97vgTfQnVToYORxdH2BBOVuqcCHtPPV
zLx/amO6qECK9yK+pl3ZH9m5nJjIuDkcIJctfuCbhJCIwBQNIWCcBYZ5W/gFHoTa7tJLPdWbJlXK
tP6IPwt6Cl934CpUO5NMjeIhmXiW9JRt5hK5oCF5LS5nm8YhbC5gEipoBFnmnluIOzLv9y2GDXI/
hRRUVAnLONrj8FyPvnFypQskhYIVv/l0HaAfMY2mKYd+aooGNVKhKQ89NLjkXdQQDPmW3EDVYgY7
gpIWRo22Blu9gJnNFmGpF6Y0DlUOsKaZBD1jXRRLS26FlOz5maGcS+vsRLXXTwyd2gESQ3EPbikP
E6kTBvr/DxLdX3NHFichJQtVa2GKO74BMgE4LflE1ZNv1cfZXoGM87aJalbQaJt7RGd4zHoN5tWm
JL6B07qW0O+l6e64uuxh8vqaelWQ/M/cw7cAsNVvDpYhF0KVK+oLjwUkSkM/ipKchFF7F8+pYxx/
q+AlrS+vyQ/hY/JvQOSdevsZhA99coqqH/et0kZTIRJ2cncyczwY7TZyHLT8MlWT3ryG1DfwbJws
M6ChbbBanyqLsUiZzmHlmxPpXMXBQbo3jsGxIkI1XpAAZFv4b0PADNnpFHo+bDB1v2zP32pv8965
iL1R5DkeoGKbdMy46zuOlfn6dP9dvw/4UAMm2jyQct/FvUuHjdobu6tOBe3GBia47V95pwIWRc0n
iGl5IjPWh1I/S1T4lR1XTMSRfZrODQt9i2cWmsrfEB7fCqZeqFacAVOKpUCOGMpaWvfI6U7SkIOg
L/3iWF9Ecfz8vsnkk5zEcFt8lw9xOa/O+jp5Bap3/2hZzESLGOLK5Ar0W1ZDCp8TcYARb+9ztYtv
hBzAu9U/iljJecwDhmNXq6mqJAnh6KgJK8Vz7LQYL83O8a5CDEw8+ACxD2C26VOa3CldJB7rs/J8
3Rh1Pu0vT/tnc4H9Njc5HvLpm5K3shBkPCuocmxxFxVpDB4LTJkhwAb3e66g1iXLPTzlHJewBL9J
/cgkjnx26oJXYfWIu0rmGwOy+4M+iwZoXi+TycdV1voidaMf8YByvRhqXm+UL7TzAz2TLDR7McuA
/W2wlibYK55k3h3vsYsY41sXgOoTpoeba1G3RyHoKbYak+qAwssKb4b27XLB7p+8S35hXMJz05a2
6qbkSSZfgHaCDzrVbZwVy9BEr+3mUQkUb/sfeYAbcQ84tYBLVd993+ACmNfjH9Agmh5Nt5RWAR5n
5otFyOOybBN4GztFad8QhAZngAQdQ2pZtUFFDSDuCoe6lT90z+moELBbT1SweFpQf2U9twUAeNUv
IauSuAWMndWnBGa5j/MN/5A/txc/cV8Agj6v7v/xPr7zxxHic8TwEFwn3Wj7lJUQN8Sb5ob4i/EW
8qaPzYKCJbj7kozUtXbKw06fufaGpasA1J3+zPl+Qw6DgaObva13TE0IlmI5j5rYlv1S4Mf8DcGi
Ug0DyyX6SuR3HawLRfsjyHQ3VWpS3yZefbk/YfzvmP3Qm8+7JpbgGBN3HeX78T+Y0mGNmFz+YFIA
bjpgloLvIs1Yf22rqT557pBwkOB9uGn2jZXBEnjZZBYzeupjzXH7efDeSwSAedKP0Dt4mQOp9ysq
nqffBh8/LrjCfBoCxLYicFg9rI0RbywXHdtFdWrxhOVXG+jDqd877a1H0ceWI3hRwY1wTq1jbUDE
mNrJvsMxP/4kxTEtNIqIPYpexIbjK5hRCV0T5l1da/KhR6IYmE6h008aFHvPqEOw132Xx+w9cnyA
J9LQ1PRXRovcdKIIZG8dbVHm3/QvJAlGDmdLd2bNwcHJzNrrGjjIYaoc/GhzBO0vadXHwUZde1Ab
wggNlhjHVmqY1ZIDzZySh5zTP/IcgMbt2dFxZs+0euVjon7vL7Iil0UbiQH6nfMsM3IhlDRgqJjy
nuzUAFgZMscxnI+NA/1Ecx6qy41MF62U5jXtAhURc8RXy8Xvfm3Sjn3Q9VnpKjx1kSiQxQJb27PN
23iQyqOW642qvtuum9/pgU1xcjsWdg+Q8jCo+u3+Ga7suX9Bg33cu1wKs3foxXtasTMW+8bip2Is
1CltvO11RotlLL/p5BIfVoa38dwcRTP9MEIYJbShul84+De2KqzRDEmQ1EqOAU3Q8w6NSJRVqzU5
0dNKlFAmC+0hpHjMJTBGmIStBx/gBvIY0tfSMMmPxE0w85SEFxeoaUgl8kXp7603O8Glo9tAfXOg
aKmRdTVuArKUAVulICjpNWGA959yGFStxOiCZMuIRikSQ2Qtm7MiYiqWuTpDL5PMlbe8oVd4Noeh
LC8cX7w1Mp2WxlUJerXiY8G3eE0oZGh04Iz4yFd8lelm5+ajkEVwe3Q13K2bkzLmoHrLk1WCJxHw
ZAru2WHkQgQjRYCMYEsn3GxSCX8D8WarKne7uEZyD+DG42qYdJTQNxMVX0f3RNFjiM2/Hu7Ewndb
cou3M+lnhqgp/pa1jC2QQdFgD4OZAKgAhjcySRwxbHm/Cf0PPJ5TOD3i4nISrqxtqcVe8wMTqpDO
LUC2k+jdPSrWZwLElosTYTfQLtVv79mf4YR+p5VOhuT2HnIUqi75mm6bR8RUylDuayLL4yFvUt6y
4X/lPezaXGfnlI8aIhjL0z1nllspOTPoqMLPrqmkVh22mmMaQ6wP3yd9Nu4R8cz182mqtsLeP+sk
tgGunlaWLIgV3dUihWPhNQcZV75VTTnQTRGKHYzVWBo/ZhtAAveFBEHK/jd6UsAFKOD1uUMTmfUr
pwEvEDIGsXmUsy4wNK4qDpWwwZCJM4STzTxaOFCN4uiUsJgFHiIyK5F43NpraXyX1wV5A9tlSk3V
hIpSsdVSErj3WJSV4uGlW8jZITUBhabWH7rWyMt1/GR5z6Iw5zJtDSGDL+QXKxXFThZe17scLBTb
fg6I4bO8ljyezwVCb0f4ALCw3nzhbpu0JvFCyx+AC+TxNLF3/4ZqDl58XQjD8hqbW43pFiM6mt/A
aSEGj86RgmolINwOgSZn4Svn9BESdI5BRaB3ytGZxLLR1f7D8sYDqjzeDJE4f3cjyvfmgi/4l9+V
B/EFqODe8lk43w0qTL20snm5fxWLs6FN3x2ko/iZPZqccpU+eWysmej9IH55Z6R8Wp43R8ByEo33
3OXRSXnUcrgaxOZfZg6IfP/CJdu7lBb40ym1sHMfPjumEzDboxYuQ43AW1OJjd9QxTxrl0oe/iU/
G66XW8Bg5r8CZ3XjESciJpHQh/6PWU25+wyproYbs7eQHzoq8EnmMRLt1EzzybHLKlEFQ2PXvuys
a5bc7bIrcgEwCEu4FxrVrt2rYGHRSzGEvCvoPXqpOSE9+uwsjJ8oWstDS8DFuqQD+nI2qOkEhdzY
3XNcjp5RwqOjkverUOD8ejy7YU/YOxrl8clEQ9XvHVS3SFOCk3CqkglxG2G0YlY6XSv6F/7T0xdg
IwJ7rlTtfkzVye3+h3qfXsSw5u9juo0UfsSgBRhSMBARgyYh15vizlNNDzKiw/dwJsBepkzDGevw
jY2HjNJyPHS0r0w8ia8GUhzaXBr4Xwudjeox1NreKPns2lEVikvpWQzevpAfaxSSMTcOYcoic8Op
fa6wqLvrUKLJMuBXpZKrcPOpBLsDqEclsK5muYlpUXYgSm10Ex5vUxwd24+5j5M+5tpMIICCJIZF
+rYd65K7SnCXO/gZYAlR1vFZUvCeAhNL6KCV/MlJCKaPiJG7pbZAdTOjU0LYDPfJVF+I1Recoud5
AGE7UhWgJXhR+1oPqEBlMQ9ZX3igIdn8zao3vBMJAXWXAL8gf4yxewy/3yEIiFiAfUaEEjCBwolF
hD35nUAant/8Dj/PhgViqAQ5vV1OmFY0mSfqdwZlF8wsCfoak9ArnFPhxlwDHHXYdi+jIO7FlGfk
8KrdNug10LId9rdrQbDPYjvey/yvjBWQ+CJJxqbosHq3Ouv7BPIbj+dLSRZlcLm6d0ADf848+Kyc
u+lx7AijiNr3zd1c0iBSkPvda8dif5j3pNr56XSS3JaGCbCO9UNeONrxFOx+hfYGWsPM5gei1c+S
emFE2w5IDSq2cKCYOnnCSKvgaFPwl2UwSgi/bV56BSNylXo6wfvtg6PjVufiBf4Nfz4D9M4xr0rt
c/BVzj2NRn/Dhy+6EBRb8ajJLCYGzSYcSXdkJFrqsSonCumSME5DnGunmZrDh1RTD2iVPTM/PAmB
jAR+iOaC2lEJVASLDfdinFFIFdQ8jDnLcovlPQSkh/lIm/IIX2cTZ/WAiR7Cw+YhV/Dv4sjPdpbt
nlHXoi+Wh2HnZpyNuqzrzZnqWjXDynBUXLfsE4NiRq/1a+Y5VXOF3d7TJ1rK738zMOuPLxPK7Lid
cL3JLhMknSxE70wQ9SLvyAuYv8mh9/NqIPY5910sQ3sO7G2+GK4/aU1brSCf1palqm+mX9OMV8dm
pk9R2b9sM0jXgwaNxIQEttaupfuFuqr2XjXEBNPeBctEus45O3mY3jr4HB5iJ355Gwll6kjxDj+q
7iH6KeZK/DleK5/oQaYowcfZafuDxQ6O0qsKgWGCqlWWMJoHPE5nvJLVDkTz2B963xmy7FZTUOSr
xbUapI+XbbMUYfXWgiNyInsiGRXsDhOrlHi0Z1QCB+g27TJuWIZOTkuj19VXLWXw2wCFJGK1V6/S
oGWgnLZdfwcl/1y+Au9EMYAYti2ezAds1EQdetSFzaf2uDbfHOu+QWan5xbpCZnbEdXLDEIRzHYD
1X6Wq5a5p+j3qF1O5GHvoqEhNjyMBLlfwh2DuqDTpF8PGd7pDtDPyhMIie02oDP0B0Cj6cNrMorX
QS03n4YPLnobQdKMGI/RmfjkohuSEpjXOfQrfflTj8x48XA9/e4g7c7ELweZAiwRWCOfJd1j/YnZ
mzi+fk5yFVjJD2kfAIgvVR1XqdZWBaZvlU2Cfq7SSc73Rx0wuNmVWmwESnUbNm4ygt9n2Kqi/AAL
K+bb4+Qp5C9RJDfED/P8/DKfGP0iXaSZdRHZP8+bAFBVHHWjrw5Qz1PxbUl2ykh8fajr2j81oElj
zOd2gjePKL1CC/w0M9LF8Ncux94IdoAgOiW+ZBMUV0i915GfNSX1rUNuuPA65mvIWF2e6Ycfmeh6
kNy5iQAnDq8dw+OtKGV93MLVixRo/POeK8HOOWcPU1tuAfiauNcmtbJJvNziXygb1JDQbvoE0/ez
6Z2ZGsR5A8P56oWT3kycaq7QMKGrkOziAHDz03iur4WH9bVNjGEkVc8c84cHkuY+PMzePUBivaxW
reAnXfiKDrjHJKEpVUJhYVZZPs1KGnmM4HE0I6xTPJk7IHTDj/4rQ+vq06E/ZrnJYyf98HbsCY23
UrlLeq5UanvTy7bjvqnYCSAxTQlwfXfi3LRGUn9aNBzcWDGxoThR2qCanHDdCAsNm/gh5R2CLbtS
Sw8t/n0c69OG6CJroRGBalGSqBFPkkDD2ZlsvXGEvAJlLrKBJY8ruX0hANsrGR3HGchy0u//x9P/
V7CpevtQO60kT2Nbn7iL+Tr/UILJDPS8ZCbm1kPD6VyGVEZWoj2+hJoV0eP4fXUMSoqZNhRHJ8h4
oBV8IeqP84Ix3TGx0eL3izK0S9eFw7ByF4llXLY7Yablj0Jfv1I+E/bu4Lh/s9smIcMP4MHJH8Aw
6HO6oXMpAcPiSutNz1SP6XyncQtY88U+pmKn4tNKI9vd2WzKRzqg414YocRaNCCWjMGm1jiIEdGu
NMT6gGSRDYeSYh9Z+VDvGq2RAoGNJbiO5K/TZkmzFGIgKJetXPxWVp0UGag8D8JCw7crlOEQHRvl
K2HZfj4bDdP9tvDkTB5ECQsPMWOWCJTAIT8jFD0xpRIGCQ++mocyZvvaHcKM/N498UNFUrBFr/+K
tPc3aO9V5WmoE0z3KlhP2p3mqetBQqCjMtYSm5vYpkK8F5bwxD6tHTNffuVmhj387zU5EgBoPfNI
I+GUfLwN74FSJUYzbE8v8RnuqwG5lQg95hwyVJ2Ofe93p4lSwfkmOfuPOULdTGFYj4l2gMkswH6B
rKuSWolcYnzYjUXdBV2YKWzK2Pw5080+63SOat2IPr+HHEl7TOUAp5LyL5mqJRlXrEOJvXmTWaoJ
yaNuuJ2UcNsK2+9rwwTgxN49HXVSWXX6x6H7S0olb31M0zeMy3Fj9KubQI9vGJXoYW12h7yJtIsq
EuWKP2ZxRfOU+f9JjaMpE3h4TzgAksEcs4YkgUAA9AiYvNHSPEexP6JoqVYl1c7PsamhuFXRl4pJ
tZ5XFU5gnSHuzBlRx1cGP0GyxJr/zThqRXGem7W2m+rIfixBaOpAZoOgTLd7k0S/qyVuzCgM+1MD
MmJE1onEYVAZ4d43Z2VMYOs4g4OXa7X24oQtuuNcdbd+sJdArp5a18jWGinsRapqoR5/jOVBsLOn
gKxxrk1JftlW7vGWDZnoWMkAkaYagn42yQgwXYHNuMhbotY0Bd2qIoaidRcUhY464oP5XKOqters
4A3juWY4DopLBDR53EazX7NWxvqz9cRlwIazNPz1z6Izkd4I2fPe4MVwVcY81YJcUhT9xcY3XfBp
yTJPvEjW1Ujhn2OgCUUctPFxfkT7yX/xQvTDAKrQcKATuiugfW2tH2Bm3d8kifK+xqoD9jPV7uZf
vE9pvKGIoQbT8f/A8YGpTcf49vGOO4mcNT6gfDhuikEWWjuzdZsVtTuJ2Y2Tu2pobIwMe9QRn/fB
0agcBTsGxorDm0QYibaMEyRdCmUeQ0yMg7FufMClK40n3DlVReZ68mU2FO/w44RLmh49Dt0z3pet
ilo1UfdN2+2JdMVxpK5zBEGc73GINppm7zIFvFYRc1CHDnFN0utaAvxJTR+lPQPq0aoNBzhBrnEH
CLTfq+VtzZheypDMmoAKKTrnFhYYWEG7/Xe48qBwMZnoFDn/KkRDHVGgDkVoMKnykQUw1zCmjC1h
uqI28uxesqGrcSH6KxAmFmHCsitzk8apQrqCtdqo6l7XWZvMo8knkJCme8tGzmxmbjrJZGsGTBlK
J9dGD2auyVTpIhKvDOVmghf7cq4finrZWWMhx5vjsFoD8l6VCDWYQbEU7QwAUnq6pZrjSDQbVCQ7
i4k2FTiSfZJ8p2XHt2xL+yg3mGEiaHso6QxxJRHWpQzrE1w0kliHMq/F0c9WuFzoNvuOHPEon4z6
1opfTSECq0MN4caOhnFkawWyOO7GOpBigy3/5duLxx4TXlKGIHzCg9gFG7GqQJAfSBfANCIhZ6d6
fAFWFE3th12K5zNmlLpG47dcAQIPUNma2wTgq5/8D2DD54h7wMaZtB/8QVPgtLCx3IMEtvP9YCt0
GXGRGTcb7IR4QyPzoAa7m1FLioztHYNocKw1lQKZSaHoOO7EQ3A0J4IvV/4vveafAm3PAGlehgmd
/ZOZO+IOFzKy6XXd64e3d0CjVzl0WT2KkB04MdSwxSP+ye9rZl4crttv2SV3QlBC9vzVZbLeKRwC
ac0cDoWBc4UvLEOltBa9l1Ht0q/zerUjTr/zLLzRNtc9qBGBXiqkYdQVMGtbUbTn0jli+rrVrsrO
fmK8pwP/AkrMXR37uPRf+2pDXaUaCcQ7zM6wnwpsJQELz236ercYdVNo8To1uSZ6nvezXVGqtzHx
r2sFsfYd67SbsgUWBNS/zE65nQMirULRpm28tsjHZdnW8N6CtBdW97WgO9BYrTx9HVtePJ711Rkq
BhaLUsPQn4rPXmvq3h8xvc/nmv1/cnIQovdjELQpl/sn2UwLwXUhQuUtrG8h9na9ipSKod0Da02m
1p5RihKnodUU9rCPOtmJsohDYFL4b6nS8/HpFL0A0SbuGUYXoobzq5vCLIPjqAPig7fQshIiAoN8
spG1hIiFIcmdeOfrw3kt/plWSq7zL/nsZmbbnC9GosUEQ9GXjscoYqEPhMK3GC7WdOZfDSpvG5MX
LJEJHwPcJsOYz4FGf8UXlk9+qS/viePytmty8y27NzyRnJ4sAp5dDhfrdamSlixX43WDoUjZe+wC
wyN+pR8jM6JdqvvVMp++9TXEYgqRPKbdWXjQ/zs74gz+2M1F2ZZPnvsTPy4K7yGox8681Bjue43/
vRskXNuDfiED4TV76RMokqVrc3ORX0lQoLD6aSK+o94ejVigm/do2GLJjhYlDEO+SEb7eFfqdaGe
amkFua0A9VOCFVJTFgdTpZQYdOTemFM+gzwTl2IkiNtN5YGYHgzXUb7/gHfu8BFjFKAe8qfvM96Y
mrqBT3fLLYgVxIbU3ZbSQvy8WVcauJcLJ2uevYXszb14f0vI5yCQEnAya3mjV4486NG7lw1z54cN
Vgxd/Kn+0U5wVUh4lRwUtS5I+blVH6My/rQWlh0KZBiLzIbFNG0whUD7yZDbK2fYRs8t1nue6Su3
L8RWCz6FsSRYc0dnq1XkooxLUwJZw/pZogaK85QBedRP1pC32eV8zpHJmde3zbWCkpWPlHRsfmgA
lu1tyyXuuzlHiyzd9/3fup+/ddQ11MsHuK4h8XWjPB1UjAlY2rNh/rLQ1nDz1E8M01bN1YdHMXAR
fS2DVbfo7Gl5iYq/kC267cJ3P0WkiP+gEfmQIaM3CwmgGJmS+wYB/xLbE56cvbXHsokvVjU0MK3m
NarzE3EsNGCaZ3vVW/gLKavM/KzO2C8W2tjZCS0ZaWZY8MQ+mrkHnHI92Zq+I6scIT01F2tQoK2b
mAQ0uJlMRks6z3eAT1k5zQkNSmtEbahuBhx4KV/1HJspJbensSOZKdxVAdSiLoy9ZfAPddfMCrgC
W3pdUhaIHS0hx5pUgQKhdZuqYQzYZl4ecHoY/adGHpHMiUDzJw72Ok7kzIA5cZtxduzBk+D84bnW
kv0qh1XSGSqxJuvqdS08nvgWqgamm6f6iwBteU3EeZVG0R+c+I4ceAep3loxRnqqCKaB5/dSYpz6
5dWExiklFpOvMHzW2t0OV39RHimQs6p+Htwy4R/6+ehEAmXJ8dXv2FrMuHu1ErQ9fBFaNBOrUm3/
oC8IZnBMPAyZV7QRQ8PnAPiWlEkYXPq83sjcIeCEg4XtZr+kS6EqicrxcD3/iqWZYH7YYvTkv5h7
C3IbTAeZ8EYudM7zyBFtVAum7PYNIzCyVm1wuqjKGshNnDEq+AmqF6UuWIryDdg9R3aZyZSRtaSI
oMldRCoG4sWOZApj9yOA98SKX0zvp3kQdJOdv0pljATkrsNr1z4WusR7ZW/XFgJBLFDKBGalsOQq
Tpt7b6XsZ46lQXsnZXFWm1aaqTu6V+CkkMwvIOCM1s3DjTih2UoV+XKNK+QlkPjTwT+8+r8xuHgy
ZDxb81KOaa+GfODeA2f+lyiZEb3JIXxgURJ0RgtD3haxZ7gN8SagCNtPFQxmYophuuHRIIeHLAQ3
+Nq50rneOdxfXOJrH9c70ITByB8bPBfBWsLXdu+0mTpvvaK9nNP+O8uhgBksK6GEiaVvJCeYvrzJ
olY3wNvsFyBdF89hu5JJcIv/58kVqY4Vt0RuENoMPSndkj0RIAKGRdVfxC1zg67X72NtzkyWFNAw
TNCEdiNDHbZRFj6aRpPeyszxKt2p2Kazz6pA2y6sU+jT1NIY3TflC6qCM7IytpcDPalKsxRx+36+
Wc6DYnjo4bUNht5l89jWrdhiIQP+yinj6gEmmIt6CeCcqW0awkaQpcUmjZH9DXtegv4+ErsxTvEO
rnjUHxmQFNFiWbnfQCCD/lBHohtrdDfdpGCg5Jd+CwurAYLXVai+yMCw9w02FE7zT7ATQGVmUO59
++qY+ZrYLW4LN3D3AR1qyrPoYMp7i8yOysX1tzwvmLcRUU4UWza5QrbhOYJbEgyBWik3COO0RLyU
AYjA5AlKWGpRL4EZ/BFMubza26Tdq7rmzaQ6JqmItYTiEn1MKiPjYrnddXChBkfh0r0jKtWdjh/F
KODgJObUX1qDs5yigYUY6bDizzUWF/3S+z2+elOFy6pUi/UD+XjVNWoOpKWKbuWOTroqGKtGgG7j
OEAjwzBoiF/NYFwhoRwxG2SoUgJb+JhkVg2pGvhj+V9e5npGdKPKbU9LQvGB7FXagywlRB6xOInM
axecwpYAVW9aGmEZN4Me3S4K3YWZkt07wT6eobIWgjLKcDUggkW+4Jj9dKGuVXeLQxZ7kdDLzHBz
x65OpCXGtoK6We/urE43HJdPg+sCqjehyhcd3/PhHff7w0p1jSH5osyUtzK+rKlMlKQDGEHLPl5h
kFVQ2qyQJNJJbRftq2ulJ8jpt8cXVhoO4sNo+gLLOLZTjt3jHMLnvR2dB3IQ31G840cvkrxHjJrC
e8wiythpEKrqEHiju1HkpGEmTeGomEwb+8VWMOiVr17nL6QH99Loxi+wq92qMdHSkjdXWzG0Okro
/tF+ZSburXzQE3EH6wNoFBqTfsp2v9PvJNlGbDDpGnccgyJXRm291609a78hQSb3jdqMG00UdJOh
7d5yZxVfxiJGOk63l/AFYgLZjkDnaT6wLlRLHaaCKxqBjQSV6pXpZ7ePDCbUScR1s6hykELnPfiy
NqrSy1MnKtP7MqnNiidPU/RL2w+OrFehKB5UPP411efpvJee6LI1MQYbklYjVeIuPt/mnHnRwfxp
YfynAf1P6Gs8TGdFQF1Oj97EFG+YfF058mvDFBxd2dziGH5YRjNSX3beYszmV3h2AkyLyIerFyXP
IUJ4ELbneli172WA7JH105BvkGngUYT2K9gaeCSQvmqT7ILZ7TAPdkops85nPmYYSxQArWwo3HY5
kGRpwqF0WjqWLaJIJILgYrf+TJIqk4Hh6tted0n0BEWhA0HcY9B9RvPcr1oAhwSo/qYQgzH25/Se
/u5xAHd6C0GLiKWA9DS3uw64/7l1WHqUnQR9oUoU4z8ViowY9pgrZns5ZVtb2vHS9yOz5puINGXB
uGwvG4AH5yPHgGF+OEbYSmkFg4+VGuLsEiDy2unftEZF8fZieH9o9TGHf4BfeGOIW+9XpF378IfM
b7S1MCbfQbuqyOp9thbbAdnWLWlZprL8jMeVg4ZjXpDMBLtAxAKAyr37Bjdq8pyMxe2cizOX4c/k
dKtDwhLbgKiyoQfeoRK4uqNG8s+neOcRrKLs1N2zQfCZxcnc2neNFDt+MC1GG0TkRmQf3PorI07G
V8BG/uY4PnW8QlZGsdsG6HgPKJxlYNiLMLjj+NlGUb1m+SMVcKXO49m+Qxk5hPYH9JYK7hXAUck1
qdJORpdyktJQyKFjl0kYLtOWwaG+Sf7GvTXttMo4pErsMkil+tvsjSgEjkCQQIAcd0JcIobuuXUR
T9FW7wAsjhEDmt4z8kxiMI/77Mi1GudVrSVX05jz/L4VqaLMzYNZfI7sUMtS6qLD/CkURZQeAO9a
4UPJzUWY1zqcA5Z25D2Pix5zN5b/O3OL84xQaS+hdIsqgLkF65cEu77/AV2vic0H77FuWewbnSe4
M6pO63jPVQ+gCf9EBz1WdMFHwNeBDGYyEG/Yc/ubAL3jTTE0nR15al7THPNybvhDsAzE8n/v8Pb3
JMFpUFGfdC9UPz1ckDtCQj4E8c/FGFKkMzCaVQkJr8AOM3EXr+5XiKThhlH5U1TIjYp4nycWWAAe
4KRPfAAnYP7PDMgtZUjUeUbTnmOwuNbzXmkdGeO2ajgjCqBPUfl4DPFlQv7gIVL8EFB9Qc+A51wL
9c6HZZ7zHRoBUWA0u6qBtRNFdaHaj7xIEH0RJQFOelnpILEOSy2idNFBGzvZ2hd4JcHhMj+r5P2Y
V36vuqIjdM58I/RRZGfDx7GRU3tm/mYn4ebUrxY8V6WDqfT6anp0a1D+qrGloi48g9GIxExogkWN
bahbhQt0Z6fOvhTV8utgLwZPhltDxNT2dJUggjP4djwiTWVj26dLGtVr+QneTtpPJO+pxL+DtblR
NFUWQgJcRGJyexLRQnr0S1W+9OsN8PdDYxwxlFwmS6jJm3cEPg+bA5u+2ak4rX5MDZC8AJy6FshF
ZdIsg5WAvhUSO1pRnamhb314MsJjzw5nx5t8jqX9Rhg9FMdbLvE2NdJ1I1Hhe/9OGqi+KGjGqiF/
SdXmCioT2LkccchVl6S3DXZgEvFHmKQ5PYq61FaB0atmYJyg7Kp3q1DjBKXu5G4QCleDfhm9/EOS
oBfptRhO1EUwPpIHWDL+9CFahdPEqE8McaSq5AHzH0wDwtzBOz8SPLGHZ8kkcnCvYwTXo9J16Y7T
HHOQJSzGlWYgAB5p3lGF9uib/l0VYUaLe1ex02IX2WW4QKo5wNa+5//WhoYoOUTzZmkMY/hUfdNM
BVxo8+xIwOjSmhiB0me26ZdACxd285HuPCOIqq2sO5Ayk49xWf0tr+mespcQwQFs0stVrqmg1qhI
j2R21Nw1AidbTzEpR/ruArXfdAaf7xdc7oUqsAbztyY+jMrGgjC8TSV7GyL58eTnrUrJeeLR2y+g
Frk702BPDZpJ3/pxKdbubxmMJv7qj3J4ivbFKttQzJ7DhFPbMnLVrs6L+xMJwRPfx1foMyVXCS9Z
Om3Yd4mbL3d8VpIyxMicMAwttw2dQboC9BknJ4Q3DVM3LmfHygJ8y/wfof53xpWXA1fTPzzCircC
wnfdYFzNyY/UmX5FpdkiPBfhIgC6fOFJMQntUCx/NdKiPWyMimMRhUD5n/FtyoxRmfgvc/pchwqq
slJbo/LS+mHXCmSz610RvqXxLz5fVoGmQSMFhE8oLsr7IjLP4TAe8V6tDg73pzHx36F91uOlTUwg
eizLblfN/GXkJfoIy+nlzpk3CU9HYh8oEdsnYyakBDvcoLAC75K/xRz7fkVPxLzq5LFjhNdkBi6X
ff9NIXDDcSfJ07OQ/Hq/hMDm9JEwKqkgL7mo0sIGA6Ijz9poNYnufjiyfPD/GMwb2z1DiJoWxlsf
xmZ5QNAaSmTUJOGNKNvUHzk4t2tr1j4ME3BOHmmPQG1XNLl7hti+xMSLaRP3vbYZ/o3K7848hBKo
Jz/mpxLC3aexf8sKDOHaog4ghfmf/DDlwDsICKv8mI1LUPWGex8qnl6VlmlstymuPtK68HozbwtV
UTnRk6AEXNhOLaQbi73EmS2dHPZwx4/O7ZFj0fmmyVrQ3m0fkJ0jaa7avWotfqwUr4XusRPzO4yw
HgxDhhC2TyDyCQcwhN3TUZH6mLdZYSwRri+7HZo+QDXV7mh4Krdx3n4b64kfFRJBjoz+qzqnXqe/
6ErrP+QQN5XjI9U2BmH/rQusyBucV83f09s1Ya1ymhuPuHor0Y3SErUFE0nh+kzxVGiPG316ji5B
TCP/a5LOkayqsJCLpRppXZiu8LSdTy+eGdnzG74m68SRDtaumdBsaedtWR0xQRw+AObCvB0PT4ig
Fgi81E2ISo/g/yIqGr+4PtGw8+Hi++CDHLYPAcbLvVEqdoXTtNhj4ESD68J+LEEj3pSWHgIVBEKP
0g6S81ZpEHjooO0ePSKlh5sjal4Vhw5nlVLguMiBo9Y0+Mw7wsu+UFnSIrQ7n/mTiH8zTRgh9Ezj
3haz5kBnbf+dZmNflD1biF9ThZ7iohfx7FKUSR5ciR4Z5mtlycaneQl10XonA/8e5mzwCm23ueRV
8iOhMoMdANxD9/IuX+y8CIB+m7h/v3ErzW13KXvrdT2gsLUfr/eHWekYk3OxXEOtfCGjQecQW0MN
3RHlxKkQyl8nYz7HjQq7PDpoiR3JJBZJTI967QM69y/Z2rrX1Ux6XEclnjkzebILandlgDL/G95Q
zmZy8p3Ns5MFHA9sG4X7YGarM5015vZXV7hlam2BRgkgAeiHaCQe8OlHo1SaRw9eBg212rDObGet
5CftspfPgjl5VrubizNcW69W3JtrDpIK1Idz51WOUKh5qP3Ki0kqeHv3B5SfE8kNBbHRW2Xvyvu1
+ALhHc3BOrtiowrJOH0WLEVFb07lY7JCrcuS8gdGrxKZFqn6wHTBEDM1VIwmFGeO0eZRQ4FA1QP0
LcjgWpF5/ANDfUDOwS8SbtsaQo8zy1HEFnMG4ocBzttUzSTns+ZvJtG3MlM9KeA51c/zuLeoAzK5
V+wA2xIwB0ASpompWn04Fm6yL9XhUptWFm3YsBZu2ln13+dWvruQg7Jj6LcY+trYlWBXxQ7+tOpu
kWn0p3I+UpBkWrKlsaTbNoTl6oYN22qkFXWT9odfNtzTWnpqcuTiuI9uKbzcQUdrjOBq1j4W5z4r
e8nkAEJ3P5eDj59SedBOaQy4Js2A2iehW9CT9CQsQfkI7UpBI5Q3TRMTLPtPh+wvYfdpPCwLST+t
ooDqpmXCzUKRuGnzI5D5fp8nMehyrS2h7d5/ZzuOuj2ibuxXKJtWUS5zSDs8bls0n+o8iXUsNaZ/
PcZKFxYYH22/4crXwC7HlxGiYchozdWkuryk8htpRqB2uDRabd8NUOj+lX+P6MTvm1weJPgXUaes
tt/H9QOMGI3blGzkbB7CfMstTDw/HRaBTC+SWNcucAid1KyhAYG+Q7G3GTzzWY11AUPLd+su8dYJ
Z7cV3p+RrrZZevnMcOM5YAdJVA/F6d3DaT09I+cyflDVWJIwSiszt5oPoRaQGgN+SYgc+1dr0k4r
tLG68yIoKMErtWf+ueP8AQari8p2NI8NR9BcFgGCLgZxfoVz6qFfgunalufiqBjQz1aK9G4yHyC6
PoMqy8pc0nm4TKkuypAUQ5mteJdJC85wDhxy9sl/W4TVeXuWTbUl5OqHYyR13n0/o6GDSCA7VMGQ
JPi5/qN+B+xcdZ4EaK3ztJfI2g0UflWSq8wJm9BBZFp//mjM8fg+Ny7v2kErnYBooLbKP7NJAbPX
JVSxpFbJxEKiR+S2VfjlHYuBtw8kLP97Bi7JfxulHfpLx9R43QT1fReX582dRZBvGAcPxrx/20WO
331WYqMwDJ+ZwdKEWpQYc5MkQXQyl9mN1kCg1ZpVOIFLIQqg33LIR1Gk1WXUuR/XgMWXk2qEQ6L/
xzGgXlBPFibeJIbDRWkHR/nurIHFz/JbpwGL1oaBFvJeGUziWSTW1ONrvQEesFfRIUi1C12lOdK8
1tSNvfp6kqsVg3Cz1l3027MHr4mih5nifLfwACo6hwZNOyKCxMgxPFk7WrQx/3psExuIQCB1OXpD
PlzzDm0Sq/vsJV8lVwSi8BXMP/jCwJ+YKZo9ycwFWLQqy+YPMJnxVaYibcgfKS0ph2fYd7gWmZNQ
pKlmWdfrARfHugEWGJTWqy4kw2OI8XMGkGGzVU5odVHDZ42IiFCkgk+QFvu3urxleM2W1YD0wIxZ
GmUvZQZLvFB4/9kx7SColSITuQCspDv+GOjtC7LyCvothMdJ+hAfxU3cGhT2y2KTD7CHlzABgYZg
ISklEaeSqm1j7CJNZhBZ6H2zi3Odoq+Mjd/ukjHHSW62qBnsZPxxKNoZSzM92kyn+LSY/utlfnRV
IRtaYndVtZaqRnC3DrL/DgFKP0gMbYr29i+o1T4Hepb75FggYF05qBLBNGDzyfH4x+T3d+1PEMDi
8M/EIV3twnuzdp3X0+g6jjGQBTa5bPb+4pODyfjN1HTgA8DgPCoDlmoErKIDPW3SBXgm5Y7HxlIL
x+taX0+IjxyBryT853X/kR3J8b4n6CLoilH+s0ZDpj4RG2wp9MnHq0ZykKYxJCKX8X3akzo9Rb/a
vnd/L6O6/TbtlamE+BQ23GBmyxWpm+6xsHzvr7MwMqeXmWXQCJyREVd02JQKIMiQPan9w7pG2YAH
SIdUYHlcb+zLq9vClNM5urqsgHioCGHceCGlaU8TSynMs+KpuWuM+n2WYxD+yDGlzkOQ3hrjveMa
YUytYCImDNg/foeFv/0gZrCtlSYd8aIryAdzBxh0YD/wskLgM8NItdf8kSs52R2QG9zlCdmkxUWX
T1WkF3M87i2CEoSOmRF/PuZgBO0XxW6CNJCKRd2PtJBkDmGDTF7Gx1sy/L8Cs5V1lHsrM0CpjIWs
1kRmSw7sFS/VHH69yCv36zgJ7dldkP2YRp9rKgDSOD2CcVN3fbgs8xWAoAZrp3FUksE3pwlwjBbl
SMhz6qD6q2mt8baLnKu1L+O2xQJheC0e+PTZBOpGHa63m1YTB9N+wOt4Phayj7LjZWpBG3M4StGh
aA8j4srl08C1/t8zKF2JjODpZPSQDlisu1yLMqPHO0iW2wCw/k4JmOqvKBXO7BwF3ZawlEIpmC+v
iaaxUdmoQSKTcwhsaDY2RlX5ttLIhehc52JLZ7sO6JWC9TCHPRDjoOCjQqdkjZiRvxwsDBeK2UmQ
lVwgNDYWRtCVRRokRjGu1bW5tELDF/gmVk/0a0rMBODzgGvTXf3oIvIa7SuX65Eodr4+jP55vp/Y
ClDifIb+0XIBGAWM+UGDFKG8eZ1m8lANTsFvw0MookYY2helMIlH5eeqqfEAlzG/DXKU7dVwp4Lg
PN5Vvr7V0F2gPqXo0egWLCzBD4Iq5n4xOqlZ4Rh+6rZbgxmdnl2oqH2JwCNWJI00YwR7H6jDu6dZ
KTzmkk+/zKNtTNXuOcC2MaOqoex09mKh6cgAvkz676G4o7E/Zf3tCKTwGPiBkdZiHAxjlRMZYuN9
QfWHGwJsN1t8Po6X9epXJLjPNmuXfvLoyzrJ0ZkDYtuhRQqjpOQ/bp7sfcnIgUOPNxAJT4o/n2/b
n9dH4anOyFqRMtJg8kFvzAHOPZ0GGTNjwXOA5JhqVI5G1cj5R6zG0X4XhYWZZc+acmDwSV+hexZq
Fp4OhyyDaLYQM35xiQj9YrzzEU7KWNeIaF1Lh6QVKb/L6vnseyP14FWKC7hK36HP7+G9Lioh6W2m
EbbrjHEzbBgfn0ks5LBV6P8KMfLI29+qTNVg+FTiJuFL9Qj9vLqcxdWiiTEs18gruXO6Wd6WowMI
tet4ZIPDR5GCeCwdbKgqBrRMOZQE9FrA6jFUA4tOfNNamL98a7d5X012gJz+NuE12DFnRYvA5C0x
EJYFv4hv8CclSe38HPF5Nx1izB/u5hxhbjNJG3jN9rbbS3ZSqAczYihDTvN5zDri/tbtRZ28MAXO
v/UIE7WcqU7QLUFkKS5hA+vBtSqedam3hLpkSxtczagNBcE+kaR7gEJOVge6zLXclmegdfRCFkhj
2wB5vtUpAr0pjw3dbis4qCimxfwqT86qx5fk9sWrNSbzQwB8BTRuoB3uWQeOoV4yQ5txN60Cc0Iu
eOpzlfk9zmyjeBDxb/OrAvHhNM/Cm3VigWYJLCnGXS419rwMyMkHmO0dmp3uHsWoMyo3RTl2zvE2
qx2ePfD2fK56rMgJD73be4OaVWmudSTrl41x0zyAAuTUu8j/ivo91dlTXMxmchgb/SsbZOuL43Sv
NU22951qI5YA+5ZqzqjfWzFHmXPtoA7nzxGgBC1TslJBROywElIcfhaMOVCGYlek2V6DbcBKX9He
fZQCjhG0RQDXMw/o4XAI7Ceu6/iEcVgMrw2z9Lobf1B+n+HvkaApd1XAu7ZZkAIHVAJlQw2d9Ov5
9qr98FAK83KTVMAQn4fuTox0AM0Op8hJFpn5D9k9Ll39ZwabjVUVBombeZGk9yCfnO0jsp3ZrDsN
UvYH6oPO2FeDpWKP3mE+OuPJYPD2bjnikOxU3v0fhLIrp5dt8O/ThQFG5ud0GLvY5j0PnOpHXLhs
RR4GGzlkn9aHvaXmUNH3nGAVM3q/rov3zVd3nCk9Ra6T8wV1N/hiMhP1v8t4jaMKe2LwRaOnTVnN
/snl0NLP1cXUKZEREG6VvFm6lORSAhPVO2VfCp1Xr+Dz+p7ssvkgskJ9AOs1kM+50ltwRSct2kld
6G1X8s214s0gdnU2YbUvcySyfPfmVSjqMZDW4r7kBaqjM/g/n5mQ5nlFbe7C6LahKY6LpZW0i0sQ
RiLwknmI4uLv2SFpUaATHQSyoqtqALUapLOhczEgiCDM26oebL2S+H9AjEiskOnh5eUQMAPvofzd
qIY2wLzSyL6T073rh8CTQHYKl6+a+1Lmac+MfuhFsg1lZbLXIJRKBWGwPv/lPFZAGgKPvMs0ywnk
mIBdiP3C0zLVjv8JCo4fpB6TcfzqxuuZ6XF06MB0KjxCNNo8CToEA/vSO23CkN0KJDCzwnpZIfkN
ogh7+QgpAWr+AT29WAOF1rLs6v3Jk5N0FOi4malats6cCUuSZCjfZOVwd7iGvst24sofvGecTMvM
Ztek64ylxnfzsgygWskjUdteGxA9JvzwBfylFyl8wgeW1AYg1ULo+qT2xyY2I82mYzhUAdq8BTOq
kJi2jT6w6uMoQdWoka3VW+eGpT8tEAysZiXe+e+AtEjxMuSfCCIDr9Sm9skF0jvLOLtGAUtY5G7z
DlC3zkgHHsKrGZeL80FluXXCpucqkw/m8N9yBicPcZaHCn918Dl+Jmr3WeVtvHhgKURke87DP3gC
9HENa1Dy365FTLZh4EqoeqUdlhOPRj3bk3mp/aci7TGDBMfIur7owYiBk9+WwPd7UOanaMLnaijh
T6oFEe6bdbJ3dYf3HK/777Qr6Nr/SAy8cGNThq9hBh3KBZPPycaJXWTdnmsVeaNWR0Lw/Zsa7nbG
khdJqwpSpEpViSmZJ5okMt3aO5KKsL2Q1t5fohv7hd5ZnBE8EAl9eIWqsl5bRuf+UouunEXamLhR
oo1sf2CrSLF2ktvO7ME9l4RNEXp+bT6LtD1X72V2RNcdMlr87covrqLvhtuGz78NRQA9Sqgm5Ku5
HRyCV4nZUeYhdJ9nILxZqawgnRbROq2UoYkrGdADjPBa04YSLefZYl5vq0K+VAxpzdXrvxYJdtHi
1roUUvlhlsjb84P9RpX65YzRel7kCcMsm8mJh5QQZCLuYZybYZ26YP+NDj0fqvMbMs7nhsZ2jB4B
5DLUJNQQyBmTWw1daqDdNXHKG3tPlzH0rm7zLfpdCPfyTrvLml4B4CCtF8YSsqK2oESQYsBbqAx1
g2a4w2hI276/URYLxO3i5l2mZRN5Q2cOrwnY9/hAKdqKSt2UFCopvPusYnHMCFRFwiNldJ35zGyT
p8UD2a82W7dSF8RhwjMe9Yf8tLP7mrmt7g+Ezr3ycKuOgS1n0E5Aho0uq0O5l73Wtyql+Gg9jv0W
eqFTYT0is2CesEIi8ebE9JwgJhfcGXVaJifiHbfzP0O+Aa+vJRK5bmDKHtRDMLGQbuglgR/Ty+8h
8wrgrOiKV2vTwKp4ImlL4cD49u2DvytJaaVu7tJ4LUnLAUAG2R/+ZPkiIvaTj5kxkCSUsw1B6Qcu
uv5/jWdrgJmbk6+SYSEQh3wpxpDDZdPIoKXautPxX403oq3/MT7KL7DkZrIlmr5FXS7ahWbAjqQa
aPVfBhv0P7uXq/sACpoo3DNC30WivlNogkx4Tln94bmKw7QPmOQGPbITW3rYXc7ONmY6RXGOFlMQ
PEBWBB+kR+IfLwJNThu7iunlDiy58W1zpgfQU81MbJowSto1IRsBdF7QQD9BlvNJTqymUV0T7JDb
JSQ9V0g6d0PLlnRiNgN58TWs7edTFjVgJoClugq1fX7heZW/OkXC1Z2KlCp4d0gmckSMCAFGsxka
UnH5amDNwQVZi2NkOFjsnoWKxda5pRkUKv4198fvcF6B9Ja6xVEQB9AtWUc5i0jwvOWPZ3N9wSOp
Mmxdz5LxGz3Tw+HCre+50dEN7K7lRXkvkTKMvlonczpKl8dWkOH4yEbaincJp6zq78n4NWQ5onSh
63Tr/IYNcjrATIrAUxXgAIHhFkxgRimZzFYZo08gA0hXnpbPCjS9tsa3wl/N21yU3/oHWvHQYt4W
vmdwymI4wKZs6jq5P86bG+wKv8GR6YuzB3qfaFvkyl1R+8gFgjRFJQXr8Q79JKXsBMEf4PU8sZ9P
RmaSD+NAVKMzpQYFPwa2XUkVzy6hqvLUR73GyeSNgy/8GGeGPUUj5gyy8gsS9UqrwakXn98DQABu
plOxISzS7+iyPs67aXdJ+UoO27IhTy2pm646Ot0D/RG4jE+v9MsFxYUIzyQ5cXDmtO6xhq2T1szE
8dRN7UOJU/fMcYoG3Ahck8ywlbx6n+NwJM+foOFtEm+1qqRESgh10wowkvc06CSNTdXs5/GZYy7g
S7S5A1ujNJZl2ee38+UzTxapRSqoX2RtkPdwos5qQJmhJWidAvHPWIQo4+/1WHTHDNFLyx1wUIfF
lUh1Jt+U9ExiGLgIQVRlb+0OXS2aLpOU5m6JhWJz68JCFeX8cVOC/inzDddRie0LMzku5loqirn5
ZSseuxaudwtEAt11ysRqXXXEgI3n7JtyI8ocgXPH9HpTSgruTQFTcT6t0N7rmmMTrTyiElF7JxQx
yzSDtnoYwgt+WaIVUGTjuym5Qtv3iY8IV+CcNi9uGu9fHzpI6MoWOqAlVCwisSZJRyDCvLfMurSH
OCLmVgyQH42nVwxJWFnY1hAK59lTXlhhWxnR77K9mWJH5vPGkJ1JFvq3Etn/NXOl7zVvWDNklxFz
uk98MTZQuh79ihbV5fCVFtfVlZLooOY28GLOWvZYpZeXRsnAVAT7emgXz3cEJN8JDMrqrSfuD3OE
0T/y/pKF2A+KPmLy1MZyadMJKZr4R9r1t/v0HENrNG/tbytdE96DLfcTOVa80s8ajueND9tW15aK
uQKCuyrAJT6e3mssXLtfO70aflUaAGy+iMYiN+hxkuJbyKnPgeF0XBLKu8uDsZ2S4LchfnnIP6fo
p/z3sd3JcKq87qNvApQouVrMDKPNFZ647qtGXD+YJKGgkCH30pZK7H7TyvBSLaOkyDTlGPZFByx5
6zuX+UH/Dlp0PIMYUmNn3WVPjbcipY0EeqQGrRtI9vho+r51tp+NJn7iOPxVUtK4AIH9yMMW49jf
OLJSL0a8YrnggnstXiuDjkgleQkjXGTgJdXM0T50Pp3d5c6SLEZNiJuy9A+VXg8KOgYVnCZeB6bQ
8CSZMj6Vq2mB7DvWH3+V+O8tq/4wRTtPNXVvs4ZKrBkZqxKlZcGcTizfO20JeD2buE2w2iQjUgkH
an5ujY7Z5TLXzk8+BTdnIv2gb/57jpIdCK87t+EyHmL/h2YDtmk8T+ifgVO3ic1BJZYQhhgm6dBm
m8KNRJsDo4NZ1DtIq/3+Xggf7oTYVfhwepiMZYdAyK9dB50OP533rTnVsULraOYE0Z72P9rkVK+l
CypcgLGr63Ktu2HX6Rs3Y4Ys0vT3hV9xFHj0+kkJfD+FV+kjReT69l/AE6Nun0RXojaFtht1fbgH
5mfbteiLheHRFbgXsmdt6OgZe/x1VuvU6fVPYfnsS8L3gu5A18/ESkCdCczN2blcCutG1aXk+ZVj
r+Rb3U3ktIrWp7qPBf6qTjG8x4FvyiUl8yIgUR/adOAR3ZsiEbaILRRWMZ+4GbA1YMPdN1cbXQLx
P+kdL9KPrpoga//wthtfmGBIdEOBaQ5sjD5usEVfa+QvywJvx2aokTEDz99W0IUrxxGgMQngvdNa
RnobV80SloR5L1k6mYNlH8XpS8e/P2PIKBSV34UIO8DFSqBK7S8G/UMdCvb32Vq2dH2kNkal13gG
0RMZuiYEua9QWbV3YlNkxdablKUJ+3zJA8UawGsmuagmPnk2H8ZaRXq8+zlkIgAiR6VraKfw3Cb5
VlsbxtY4ayO+z2P63Y2g6Taou3eJbuaHGt4ydVIEa3/VOm0c3GQeRwDE0DRbc4GBxLzNSrAY3d+i
tP7zOKfbmGsOYauf15wbvRblLhyfl7dLGilW9skguuMFiVPikg35c3Itg4nSEsD1QyBvOm9OS5Ip
lehGfvcBpTCfzMuuiOl6NnrkPWHyw+N4hTXetBHj3oa4AABEbeqUcyMS0mjYPsoIPb+EH6PdQr6Q
Oo/lhArgtiKUQTFHqEFkl/1QDwQcXYss/2I+sUEjQKjwgtq7xeeOyueZt+5YfGKHp8cWt9ImKvWn
ZO43pkpCKh0tCWF+1dP2rvmc0/tEB6zIugMyHXvo+wvlSOFD5EL0xwVIFrYz49cV6WSx0EMD9HCl
sI/kQ569QKO/doCgKmZojx15e86tCv0h7k/BGQ5c6i3R8XpD5UMqYDqsToSKGMYwk9YUCQ9i54uZ
yR4A+7EjhafhWoMv4frJJC4M4NkHJqIXKXY5BdwknNXVToLoJaYY07qRnfGE71/pq09r7+x6lXD1
muis+mOPLA5g5endi4ty8ooZx7x08+jFDB5clYo19fLI3sqJPClNE/8Knv5UoZ4dPfAnuun+6V0g
qQULNBwIM8pGjn2AgODOwroJR4ZoK1zC4rbP3IIFRYtqj97EM8SUY+fJiIgB3L6Y4XCSfU6Ubu+S
9OLFMgGAkVs2Vqh13YBwWmfCJN1tIFZPIkPQ/AmjC2h0Wwo69dug+L0CE/JY7HiztqlbcBYF70Ol
YKbUGktv49SPmBJ/riqB9JzI2DlQu3G7dq5q7aeJh7NZQXgS91Vfi/o+JjlokKzMVZTdXcG9etBS
fEX1xCeuY/reTYPusGAn2DFY4hCwyZmrPjFHOK+iKMbyxzmT5UjOzFqQQTwofyqiM90A1ym8PTDN
ddXrmARHKT480q1g5kjGGFPnuEc5EEuO6RfPGZjMXzXDsZ2nxXMiJ84MvqJZwZHwZvHOTehfnQaa
S9FKiJr7gWTTBUC3DkrphL2ACuIkHSnWANEW8X9iAvJtJqR4ciN4QR8XncPNk8RsUgHgevn3/pUH
A8GraP/RYLzeYruXtWsE2zr2PIjvm//S3kboKGOo4Lf3qK0t+GUW1t70Fvp+GkVgeSXw6A0jdTHh
O92dQy4TtL7OH/POD3LFc2jXXNLjllJ8s70BRMmyTqQkCdDZ9I3uA5e1x1GQF5NjilsF3RYrD3wk
BssT6Z798jZAdnpU5pcDnePozHmxg88AZ2YieREMJCMwdgp7sbyLfQacf12CxVh3n5s+cIrFHwuG
5bsmYrMnjTfluqxHY0DaOBXDqZegdmokduokvM6DfICPqFnZzbAMvheZqaR0oFXbCO/o3AH0M/wn
agt3d72w3f+4QQhbrF7N8OjV3rEBj7fC8SelAoH7gysJPpUCavbhJAjedr6oKXARgWoNpSqnzZXV
yU1VL/Ew43/xCe9Ap9tchjMR9wm3NC8n2s6jlE3HESyDagZq4RABuBEtRK4s68yvtK+GgSw6AO3s
b1sb4bw3EvnK7LL9NVVaVafhQqzIBTyICOFoZftIlRzZdSu+o0S6/V8fPmaVilZdMPe+6uv10m6F
H9kz8cK1x1FFhMD8XCxjCFfNiLmJg52no/mmn79O8TLApM9nnaNv14WnbIMGpl3m0zveU6UnIWCy
UShvwMQaNJ3Up6qsPd6Jg6t0dIDPDHcNtdBQDyMQGg/5Ht4mx8Y2h3YLyINDpq10IxCCEOGdn9qw
o6m6W4GR+wteHoK5Wk0lmEOGMxRHSx9owqHo5T7lhVKsTZ0k3Ytddxu5sS+Ed1E2WFPS3v2YoP1Y
4U1NHSbg7lFsb5Nbgt+LZgKZ3ciliYTldwLiLSCzyLPQPee3MyuWVsEDugVfAo3SjhpNBGVCKAmo
6eu4dzujlvnZbzzaAAAl2WgvPDIo+BZVuQzMgJstjmdrXbcbGz6PD5l9cnbB+y7JReClVSpZZvWQ
lMiMLVjPDQBlvrOpadXkpO2PF6wbxcCALkfc8prjui4tjC/Zj4VutfuHM93iAF/EzUO79+zkJD30
arj+uZURHtiNQPWQlKv5UCbFi7qzNA4dM9VIx2CzMrN2rsyw+zJhzLDzzFCKpqpJKykJJTmiI4OA
jNFFkh5/JLFFo/k7EMNC8KlIR1N4nMfjstW5L/AL/heuWDj5vVjvEY6AMN31fvBGZOV7PMukIviF
gM9Sj94UrOQdpMvsIv7cA9Fu1Bh/LWlC60CdD60BOUOHRqYxj64jMlRKOp114+2H1RTxhIPclBHw
YC/QmciKWgxGHXog3YUYB16+aq8N5eefQhS/X1dnxF7VzSXTq4fzcEk+ZTaTE50Ky0Et7Iazb9p0
eyzzQZTttrHvoBI5bqk9lj120Z73STLUSIM9RTC6K6P/z1F5BcR46bWRpi77eGuI8KRlutfAB5AD
oY4LG7eWhB+dd/r4iOZPpMXVaTePL1b94XncAmKiBNy+ofkbLpepczQYo/Kgoz8sUv4DC4FcKB4K
J8LfuwZo8Cuq68zC06DrfgK9pIe9VRmRDHEbvb0L2zHRkaKFK0oYT6DQB5OX8+mzwzwstQVUcPYd
4c4j5AX9JAjJZhISB9pwyHWS3Oq8hiUmGGuxYFkSal3+99m/clIW48cUtTWAou7JtTmWhWd/0PZo
y6BXvP05bTMk6BrgCB7Q8WQh06nOsrlAsp6OMxASA27Tt8CAqSWuyVp5C7Yf//qlQCdG8Pi7p7O0
/blcT866uYwxFpjKbmZjAH1YCAwbsrP+wlSTTiNz70Xt/DLJPPS/BOg4rZDNBpBq0en6FymzjnS6
FCMqogQeHk+c0TfOtHDxciKPWaiSZtQUpNIel9gqzlV8LGIY0O4WC3aRneQFqWLET0dwZqmPQmNh
1LCBw+g6tiU8x3yWkz0uCY2l62yzpS7Mi4XkOg5qEcqfDjLGoq5NdTgHcBtFYrp2ufBz6WuX43za
wbUWgvv5OetRsfJGyNbyIh010Fm5aoz0NPc96DEna+pygiJnmVN8K4/1Vi9zUnAnB5p0s8G5HnUX
WSwqMIbdQk0qnoIOHQ9oa9FHd16IzAJWmCAWujZeZ/NSt0miSNCxRZIzXMBc8FamnJmnw5fmrxpX
1FFqbnI1Bzh7LGQuMpaltzGySwvl/OTk4ae8jhjHl2pWUJ7RWlDrjv3v7TQYa/cRuftgsTYJ5ZaH
qXMH7PDqaAZgzEhUxzWRn5nkbir0/yO+y1NrDHXfGoGmXMxWP45s3miHkXHRZ4LdahVunvRNvgJc
tmrLzT5qSkEj1FVAc+dMaOPeNdCKW10g6lP6qp7TiusTRrRamF95KnmG4JCpdPSqIWqMzJfXsq9T
ZNrnS/C4V9fIpH2SIcy94Y9xNqVxMSz5p6AaxFqwSPKKLW1Km/QTA+wSbp1js2cGXdHlsFig72QZ
aqb589KR8DSNTM/ULC6ESbUlQECjXh7BPP6jn9MayuT7SyiEQt/R9L4JZja/bURPnwhGkOpQopz9
MCHFiIUjc9zG6cOcBesTkTG/6GpQgiTmc+nKsEki73zqY8wi1+Gar/GPU7PiTtylPquG+WQfgjCG
ViUj3ra+Qdz4V2WZL68B2fX6C7wt1mEXb0p2dCCCd4Ib+YhcG91DAal1cgsFHo7F0t9fnffO+E87
y/RvFLCJF+CNB5QERkigy0zY3t+Xk5FZZUGQWTbhmRJCzPy5hhQomCS+nS61qf5TAoYsu4h/ir/N
FdP/MnhzYx0mj9uyUJwnBFViHhtueR9vViI/JSHk3WMm2M0Hv0WXOGYfbxLRmpH1ulcXhx+tNdsW
a7+0pdJy5DoHbQz7HuaWpevLiPJers9ot+oDWcOuEVp74LmL5xHIs/PsISZ15KRdw5aMcvOhuDdr
nf60KhZhVDBgC48aNgMkYim8j3/0HJHQ9od2kheOVRESNU82oYnX6csdkMKs900OptEDRbt5Ogyo
VI9V7qOtTavUbYbnRmlo20bMDJkGgqpYrchSfdsOf01DbtrKznITQvIRQdTmIpO3sbbdokGveAHJ
iOiX1IM0H1v6udJc01zA/SVCE1MOMdkJpaXIAZqWHwiEctknUBygK8j5Py017vIwDoNwPSbi9FSL
B3KlHNKMJmqXOunJjChgt9R0okrfeMILkqFOkmE5S8UWUzIjPpOgekfASbtrihgqh8N9pIZytiE3
2Viw9y1di5l6w9uWRDrw57gF7yLUSnqJq6dEpSkqPKJtmlG/c4KfwccUswkaFBgiL+MTBVqrXSox
HWOLpJDz767GiQW+sIwEaDC4NcsKYY6rdzc6mQemCcPcvNZyU1gEuoMKj7WHHhl7mzmp3RUZRLDL
vOvdnY02LIrOZePhrCuMNCdqg6MZW1Och7thhQekvBZREMySLt1CDHJWpuT8g8/KBwhz3t+MC5BC
9hpkbSQH5erdK0SAthJe+tfvMrr4KBymyZMKypN9+HTRzYn359uaf84dAdgf0CE3twQwpbT3hAi0
QXXGX5+AexH9lMDN3OGjA86nnARdt99kGBF8pA0p7ME8NYBLNzIH+a2RrpoKgiQ5N/7dYhftkY2N
Zv+t/Ab8aQviRTB4Rk8sLO0a3I/a7uBhEG53DK637H8EWPp/mYNnR9nVNU464eLpbJ0GLUhc7Xlr
Tjqi0Ez/LuCZ2BaO6h7NiX7bNgo9JzMBcWaHfoJ9RK1M7DX/Aa3dO/6EyQftDiNelo/Mr/kfzaBJ
jG+CrcKGcnVUjjdNbOkR7HShvKKfIsybX33ap2l7rq4p2EgacUBPRYq4IwL2bplrWS+WTSyjpokf
nvuIugjf/6Y5gRhOZWchtm0WlVKyVWYNTo5I1Cdcbi/FZp7Imw5vIYEUKEomQdsm8UhwHgwuQigs
TxYINTvxAVO/GXmBvP/ab7f71ItGD+F5L7kHNKk4RPXe5tczJKpeCQSs0QmCY9D5RWNk8jY/L8wm
LGAv7jgze6Ogqo6YX/YFPFflqMqFTUIhxTx2dqOZS+LMAdDcX0KwsUE+5RaIQuxOdL6knVN1NEPg
n4bTHKzgRS5J59jxfJGjGiHvzQBJ3rDewxaNDjFy+zkfbfbD/lB2Vk/27OmOxMPwUqU/SE3wPaqV
0RBM7KBPw4f0W64EjfqxayyTIrj0D3nMKfyrPjwxM3BRTpcQLUnx3hkXExTWzrBhCljYJR6JC7Ql
9SiZwpZVIhw7jMVQvUmB6OG9vhOFklZjxs3vyKsbY1oJGSzQuv/OPdt+WwzRLxH65+3pQRfbEf0v
1uU61tokrxFNk3aAQBCmQX2JRUbUpcjhiQw272OoqRjhS66FUlaRXqiBxWUekYVqDP0/3ZK26g2C
Jna5pj5+q7Xtk8XKSjWi/JzS7995SAkAr1F+bCPFTTxuGzAlu9W5yPaZlarjpg4SAwmhVuk/AdtR
bfRGKb8jG/fXBRqpLPSscdG6ApiGd1VG8mVzqCvXVf82X7+y5es7Ce/RXOG9puSUTYNe/622fv9X
/QirbEp+m3Nx8kijLOli0weyCGLxVPZWNlrHQ/SKajUu9VCUMYz8gTbx0JmsglXj82UyJ8fEaFLC
okJjc6PedDf2eWh4OZFLihk/oLkyqzir2j7EutRNZS6VznDn4xcAWF5OHH6HsnH54GNEfoq+hLsL
Yr5gUEvWGG9lYdM9Wpl7SgiFEolZAtcV2NPn9/4HbogMq1ldtn7bEaKuvlLyn/PaUynXkLRnRtyQ
ndtHQIrMEm/IkDvVRQ/VG2D98XU6hIABiJ74FVOJHtBRKgsTSC+3PawMjmZwhiCnoTzLRUzxBUJe
cLaUvDPEis8Xv0cQHVTKxPskSDq/0x6ngC1ADJiMjdg45WHrhvrou/Lii9r3BYkVa+V+4kez/c5t
wNIZZ4GiBq1mIzVJ3ldjvEoFFCthVrQynpnH2Pdac+dKMntR7FaX7aOsUMdCYLfJzDv3k2T0jo3W
tfdVfWrXd3snK8fbH/xdUc9KaepdLUk2FyoN4V3C6/Wm8O/Dn1abeTnoBrzHtKMePYSLQwnNYF2O
llhvQIIuxILvzS/0onzAm5n1RuAP8euOgZvxwwoHR9qxRuhf/lLBKMKi7pz6l9kZZpDJKetS2jPa
LTm8tc/77sGQKEC9pguI0Ax88XA4EG5ny44o6v/twUZe+UZCTQ7NSpwXMHSIgbn0WKf8VE0c8iAs
OAeanZksK7JU2A9i7U3gBX7zdOL3gVrsWp4Vxkevu/fzBCqWukoiT5VcPuiIec67jtry/LPXJWvt
qQtq78u2MZ4lpx1fCr9dHLjTRX1jEizNq0J7gXjjBHWbdUDAqAeuB9IJQyX06JvID4vgoXnOfYxj
3G5QbGiCKBMBzzowd0lHG1o1Ej6VYiimU/v60F75Sx+Gkge/FwsRG0SoWU0iKHpdlFeadXwSJCer
une20JZK9xPP5uLG5jHw687mk8EIp9tIFmXo14OOL8YqBFo8zzK3YBMpKAIP7snYc1POf7wXxJi3
IZUOvChCqGV4VNpNABqO2POY4Hh0IqR/O0vM7JwXAOMqM0W5BYNj/cTTGO6Uc7mcfbmLLvfpc9cL
f9lQ4LYz6vMtGf8UXBKK+PzUzUS9CCniHwGqbf7M33NdYGGozah7yU5WTbcwRps3rICx6alCoVkq
xKO5MSrZ3tYZIhtiw73GyDbs1+dNBBPYbqN+gWYywAjGeS+/TZPiR26vCzaYDU6h6DKQf2Yz5vAl
Zz9XqpkHADpSz3xcBV7cwIetgFLQ3uoUt0uNh+aiXV8mkiktMLkAcYnoiOPb4OB9OVqtm0j7ACQ9
938CEuFL4kja+k7U1eCh0qmMujg5UjWVJwWIRVHmNKk+WIrbYTvEZTi9xDyUrQ1kWpvmmBmYBhTr
3yl+55hEUjkwnVUcU20KVKWTnbFj0uorCpqLlsjyWiEMm3RszigW8nmkZ0UG1AZ385NfAyl/6lVe
j9n8UKKrMpmFk1pEFvG9nJ4S+blKguGXR6ZqbMMwSj/rE49wveFaFceMlAFnNVHKSk3Kqbr1Utqu
bbAdciX9rj2RmzGOfqUnQcEaFA2ztvpA6IJGAWWSdEUekZhjRbrktDPHQ9uEAAU5T/Z7FelQTG++
yFujxoBpUJ1dU304OUXDDi2uDwpgFsWwg3+K9xZ4MxzqGSkYw4nQ8jLaAK83e+fuk0UBZ9GellbO
hQlNP0PTDQqGN6HPoTFjqcJunVqPfvvsPNfLOEB7eTLtGUdWtTUonUe95J7BnsciSzbAD0zfTxKo
VhtD3ENWdLWpkb7W+HX2IcnZSysg+1ohyQPmra1fscIjeatCehLlgV8CgkOkUkLDYYQaD+3HYrhq
nAGWLV7i9HGH7KiRqkn5T/7aSrOAxbJQep3eYXPBH3eYWfxRU7EUZXRCjGBe1jXKUuvUHL7f53tR
0Ff0U8D7TxA//a6lOKf+97TftGNUf8SFdaM9zycXT9rLFIWxPT2Ftfo/4tyhe+lOyBr0OMG3FXlz
AEQSziGYxoMxO8B3jG0F4v+OMHFOuef+1aBYlZPB5nW1VhPrrWR3VYa57vgAQbMAuJi81rFVtFnT
7spEOtOmiexNM240tP1D45YvftPzY4p7pxvL/jiLoCehRzYnutP8mAC/7LwHo0qPZ8IUe+OWJXr9
7fhNAoyb+q+9GcEXc/fBwcrcsRlS9aanNW9fkGIP8EtV1MDO7MP+P02h6+TTlx8jE7U33BSgbf0s
VzbdWEQWH4SPItRavPZr0bGZeU0x3G9fG4BpYzpwlnLaLGwgxORGELTr9jDOAN9czlm1t882xmEQ
iXrxQPrDBWB3eii0NVz+APGF48kmSXsLwIMLBb4Xz1ac7wW+xPo31dF0AP+EZpJY9e/9gjGudh6g
g5RMtKlRsNQXOXCnv14yzDIr9eqdB5XVEKRJE+am4rQEJAqLs156mV8kv5sXu5p53FvqFTC+j0Y1
YzhGnF9UJwR2bv9rvWq/NsJGmGF7OAmBfBCC8A9lq3AB3F1VYF5EumLnU8tSjsdRpAGfkhNPmnu+
oO5Rh3QbzGGI4KQE0vY+/7r1vu6UiYYGDa61FKr4YEg0il7jTSfbSt0grwpOv9Jq80rhDC21Ja3W
IYpm2Ib36SwQ990282ijr/V+foVjX3dn5edHehoSLPAZVR18K1eNXDAcXH9N9fllDJtJg5pCrBlj
rD3+IGa3sIY8lJoMmxL/ABrGkuRbHvP3T48HZ1h6yuUXtfgG3Rp7f14pQhXlSYS6AX9bV9O9z8qn
/Uzii5ih9U0BhoBU69B4YRmx8LWqzcn9oH244fAjaL9IUpQv/0kdJktb5J08sw0451FRI+4U+8bn
meSj/96GZQP7YOsfXE7TpXwDFjiefTxbW9vx8bQJNGLTg21rXVUIcxPFg6m2d/gY4lGXDeLp113+
znAu2uxv5zs5eSjrpS4W/CDhqsVV0ahAZkhwsjeHP6GTLP1TgP3+CCJyHTVEc/YWvH6nP7LoElVz
oiE+9n7RqKyWg8KHRBbczpUY29gLv4bzoO1LZgQg+fT81KPUWOpY0J7yzOILUYbHGssh/m/X/5qZ
gCsb26lKI7xS46TelWXkgVupp4uW4juGMD++DRH7bkAFLbm/X4nAdWFRhpYH1oSeSojS6dmYYfIZ
f0cXvS+vofvhxraV0ZMZODY/xw16kSLcWGq6NxdHszx1m0/wbnVIWiFXmdv0BeHUk0rLr8F3YmxY
l8bNQsnvTs6Dm3vkFKKxE4YxQUl6WA6rZIjNC9EwA1zIdh63WeY6lw2cC3QJ80t8/N9Di7GyRVN0
qtwsqCnTSjLWIZTZQeC7VN36M/zJtTHlJ8bi7jA4jWNjvI0hWhvwGF0tbmSynQvkxneAMpXQSaSr
7C5+E/Bsrseiv1nsSDq/f0h2COvrdNrAnKefodVegYgbTQFFAEsvuO/ACFqE5+y7BSKevTuejup7
d/sQm6ardILzJxKgYxSidMQJEIlnjAz4Jz00tK2gmyi428TYMivaeQQcjFnfqUPGpFXVNuQowmhd
OhV3c4LLVEY2IcXWm5N+C2HRFU4LJP4pOjm9dCQ4vC7a7HcoTbi4Gs7yjGjLyzzshMnpZrvwTFog
xHfsaDBUPoEmxWDpXZZfEY5BU/QzlEvTitjZfJKTGSlrivYaea5749M/wc3YJZYNsQpoRXguhRAj
JQ5Ajs2iJHoY6B+baX+nhvy2Ipy/BiQtPHHrflNLs1OQ+jFocUcOExp6Fqt7KQ7khjQ1saNO9Lnk
/dhAHamUStxhtWPdMlEmZ6D0E/kOMlntN0yq931uq9SoC1qfFKo3Xpcahb/PNmz4PovKXdWkJfAc
TA0GXYbKMEuUKJZpDah/W/AiwTlnD2iGIaGi7YINbzKBSrPFPX28RK4GG2ZrLUdqZ8pGUY727j0r
Tou99Q7AB2VuEE1mT8/JJZvK5QppaCmomcHDMMEIcV0gtPFSbwpixRNKTzfao/7s9vt3LXpbSDme
/IR4/vAkbQmNByggrXHzPLJwAY6oNtoly7soqlpEGqj4vwPgnxcLOdbSQqKIF2bpA68CQsA99tGo
GUxPm0PSam2YU+fIzWVBlPaUjopYXH6eLQA62uw/kBvh9mbqT1Ne7fhM4oB/KSbfKu5T6iXf0AlU
xbMAiwWvbqHQ/3+utIJCokPaNSsqKuB1kbJdLPs3/J48e4+A3+CxWoi3ePIOtYD6EoD4OzTgyx8Q
IaKATlboKVjXI81yA1ibcgv5HPngSDMi6EIThWlRTS1s6TdzX9Qq+3v1wRZp27mq94ACbZIGRKYg
UsE6FQmoyHnP+cHW9bRujXx5+rR9wSLN0T3P3HGM7AxQqRVoAjUHqEApQXwYdnVDG4p1KIjTwKWH
c6sW1w9nsC1cVlV7XN5Gta8Kb0+HfsKwc6oXek1Cko57T213Ydrp6Vym9iXtZYs+JwXw2r4mbq9p
n7H7vXgxG5oY5d00m8s9bhiUCUNQySXzG2qsWq3KpmMPl4wyqviaRGh7ACUA8uoqfno82lkm8xOU
wiXJXpNTe090T+3wOjkHSN3PR6curkvObqcskzTllLOMTuG+LN4ii7BQ06Hw1jTE7x6o8nY/nKwF
+pbGymOmZMl+E8a6T+8kBjXLMdwIBjkLloJaKiINor9oRFPh+7ps1ni/zi/fTtBZ2k6oRiMCAHNL
ds30iqaQybbP4ep3NLNMlALfeVtqI9V1VuBtB80/VD7MYYSoa3eFO3gnlUVVHs239x9HwcOd3OnE
WWyYcnak1bvJC0NeeGg+hE1O+sIR13dQ7KpPDTfsvTrJSzAYM7cw3stmN2F9xtmDCNvgp+KI0ZCO
MDYT36XxzclBh1Ej4GbLl35cT27QqeUIoJoRivRGp5KszjdBgXonlC8McwwoYsmh4p7cl+GC0ixZ
AZyq0Pl8rI+gbfdf93Fr7Hv2vMUo1NNzse0Sqs0TxE5jmAaVnsh6Nu+OkaHoV4vVCMt0ij6yO9+q
oySTgieR+dvZ9IF4xIed58DEFq+gG4rb+TdjM+NGRg9m68iDuY09MONnh4O/HggUs4G2lNxV+jO2
qmzCYTkTDnHCzGAB936soJMj07FqCEgAs4be0J1yIR9NOLq9b+EboDxBTM8aIFFQlrQ6LRMkuwPu
hj80vZCYZ2EvG7OHiFk4hKSa8QDI7lEc01VJOSalJ0lz4YFXlO255DuppFPYDozoKkcrsZ963GBx
Uj93RJxVl8k4oW+pmlhLbvnA814FN7eLxuL9kHPDClfILBC2Q99KtpJ2geM/4U0T39MQJ3bbQIiq
DDCMmMWIlU1km7vXZOlBfPfjPsEAanOTl3/39vhsw/PXIILNKTWsoTcjQYSUUlyn+oLL2YsTrQp7
XKK9qIcM8daGfbvNJHUHNPatoNETVpISlqreUt19s8WrZDj/aiMSocvPWMMA1Lr5RwBOTXbUWRnX
dZ5RM2j9PWgjwXb9IdvCpuaG97SR+lJ0c6yg/7qTKxWE9sZE3nnwZJgdAzeO0fO/9TVaW0jEa2Jx
CkoXxgHvsOl3H6MJlZYW6VLdyAabkI/OS2SWAfiCNzNyVTiGU8gmlLQWxrAf1hEfH4UJbRxVzfrI
nRLHR/kHr7bHoVPvlNpyHxL357Jrocfx/3xwCQYa9eOigrOPNqybseXaSpZmgxl2L5HKuxLD6PJx
ZwgPDkmkHSHdeIPsMgnQtZZ2uAaWB4TObyTcelq/JC54GXYoEQq2E/O1PZV69LUZ2zfMa5oN+4bO
nsaK4QJMFHhlkOdsBckY3GugCliiuM4gOgm4naVlkRjJl+QZCBWfEJ4DYbu0DgHipGe50bPvMMUl
tdPfZA0YTp9MQbhlLgfIoMriWHvhP1ITRf5A7Z72u8nW7FBfdpRtyUSoMhdSnqFeD8eLFQmZIQlS
H69G5AwqL3v9cw/yjCwWY3Y5V2+jjHH6v+zisQunPYEDjZCqT9J41hCMT8DIumx/Hsp82eErvM0r
r4w4vz36XidEfoVXf4NQWguGDY61Cfj5dOOK2jOBTlV16C+8F3jA4VYuBRTWmo6TezI+5XASDjtw
QrYGViP08CgUjPEl6jTkNjL9Cyd6ycYwqT1IO194ASjeNelSyR54Jv/JTzWheSnUxu/0e8lD9bav
6tLVKKTSJXOF1KO/a9HL0uQoDi1N9fhNhLYHQvFloJtLRqsBp8cpdS1uYFma5QAEeyJe9Gowbrxq
PqUXbmEnzIrg7CUAooUvzziOqi6NsBzf5YYTbD5GCnfD1saTvO3X5hoftdzQV9sw/+vWFKxgmGsM
STukpZM3X2lG+7k4NxLMe9m4JnOhMDcFGKXVk67Z9G6OoFBanJo2pTfQ4DSUJwQbeeIr+Cs0T5AK
a2UfrTRT/kDflfKZzicFO49vbTjUGMqwZwa+JgRY4dtxZOrML+KOSjL8P7B97HyjEe65bLTFwhMf
6uaTpJ4eNIsSMxDExnoHLXWx5M6FMVkzbut7OZajnxlIxNJYhXnuMi/4ikgnX8DpimJS3AvcyZNb
l558IkVaxh5fG3gMqUaizFo7LD/H8TZOv3CPZiYVzFWBTcY8XglAq13ivqGZ2VFbAJ80m7NP0PGA
TwD9ABHSoDSWixWuyqtUGdcJDGjt1vqoy/cRBY05lffST2QGqhZ7EcGR+00tBXj9iiMSHarZqYRs
Nncj6SYq/5qvQCGnrVWKu+X77Mj/M/69Z3FfHI8rJtVm50YM8zmSl7XJ5SHOOkc87p3HUvrmSHvW
X66X65LlV4mVmvmEVIazMgHREwVzjtzKnxbYqrIHK60wNfgZzNylVsC/prd8KdHkuhWXvMK32VUr
p7XovZDb6rR8W1YGSjBPdayqVyhpZkGUSUgkp1Af6PQ9bsa1T6y0pYWpPXicW/DQVDal/QzRQCXS
SNKVG39Ha0oPzVoHqV28cgeqlR7JMGhMVS5G/HbXs4C6sWa4ABWyFAopLSldInDS74ST44tiWZ0r
oR7bMbSztGJvQNx14ix+xkZXsm6boNCkbyy8wz1nZ3bGjJU+VuobB3j4oq3Lr9ooPrlpf6/UyslF
GGmxEh/i1QbkZReqs7r26jk2/0mJfPdQUjCu9Q3lSWaLlnF3iGkBAx5luNbo7qoTL2xHnXmXN2z8
cJnPSXWOBGHyUso90+Xo1KrzgPZ8rVkc7u2aQsMrFB1MJM6PzRSI1DlCnTgFzGcwbT45Ho6YLanp
1plAw9O6CDjGT7wCWxTnjwrm/eK3l9Z9BxrVU7fSxX/WPVYB4Ke1WQ4uZftLr/Ji/9VuAht/4LTO
S9qAnBI5Cv0zIbexIvhq5bWvhlWhQQXWFCpx5mPOvmgrGVmdPh6/WnFdcLQPDkoPmHzEfvGjIRrJ
GNgboZ4ed31smrB0yNrecfBzUDelEq5whE5zanBRRZh7SQH+pae3Yil9yrjt7EIy7r5UVODulSsW
gY44iHwnV396zoDG+s03rS5hEdJEq04tFM0Mqn5zKBm72si6gL/TDbWjG3oo6Z3BksLZEC7o+VtQ
IgLDjQ0gxAlnlmwuRsfK1NdKfjhZF0p2yAj05TM754KU12YbCqM796Hd7I8KP5+hBFZAiO11khzt
LvrvJ5a/CsVDgYD/PGV2zCZ+NVJXID+/6d6EiKqG8wDcSgUdt+YDSrI2vACttmsTqECwQ6vl1WGw
HjDNUDlvoAPzGgJE+MKMxxsEiXK/iVX8jLG+wy41HcYNSlCxYI+ZPqwsL3S5y2pqgSow00EqldTm
lfxxp0uEUIPIk2zhrNDbOibiuaLmEKyIVHBRRmt6O5ut+Tmshy6zWKLdeizd3R2fdV0tE3L+jgUl
jl9jRP5sMEI7xI5MijngHEUS0SlmwN4Kc4nYlZT+3w+5UxCZnt73Yt5T5fDJr8xrjuUWQg8SSl+a
sP20+saL1wD4fQOP3k7GHSJd6QqTBWSTq+F37C072c2bbd1Ow33LJQf/AWJHRv6Pczdx6sZcWICd
kb0M2zWY9GxcPv/Gr9Nd+RtdqJNt3NmFOVjS5UPtmPbHn3eKI3fOAZP0c0+Fqe8vTPfmkBgwXeTI
/uP8pwuN0/wjL8geNQkvZoS7ervb+wUJTlb8DbXqyAQ7ZHIwXlXrkeP444IGq+Yhp1E3vBcVdBYP
MQsviTtRDCedBmwSL4UYUjacq6ExeU7dX+RlSbYtstQD2Clmmlh6cYSSYl5maqG1ZO2khK1hvfO1
Lg2vfzkB87V8JrzhmD0cNZ56EHF+aVXYQl6ne3oYK50eGEmYmib1o3x0LiPlIetxkkABNa79Ri14
44I6fXfRjSWK3hBI9ieYc3T4WQcxrymySHg8CttcOdOV+15dhVbB0sHp4Glzj83xjzMmctSmr1A3
EbHHOhlsvhbaSlWOLCAMZMUEuJLnVzV9J4m2EeeCEQEqjF1oTO5AkCuqQp+t+C/wFs4MnusN8UZy
jsHzuG/5F0LqqDWcIf4QZbD1oXopHwHsLbzhC/DbETS76awth5lqUZ1r8vOnCHyVAIGfIwOqz3DJ
IEBtADuVtKQsrxhbBASDjOLfdsaxDtphnnBG5YlEOMCvE1KG73T+4f8iRvba77SbP4BYQ3aNricY
NUlMGlZcLzDjs/dO820TQ1ntw0ghT7b3rdV1nCzliwQrxy9x2NXENRHHLERsj3jV0UfHGT+ttHlQ
Xim0ArNmt/TGykC2WAKIoSjCybqh+KHdX8EUxAEPnrpTwnho51VfvNhnmsCz053NPK/0rvm22uSt
HnuC4UOTMN5XI1p3Wg3Tl26KGZ8/0eCjUCN3wg+eHSPz99mCcWVDEr7NQ0XJFbYn18BwKViBbcdE
YcwmOHf/DRq5Ke+DwTflsj/hbKjYmpD77+WZyux070/3WhUxc/fqZ7wIFKteBtJN6yjNdFUB7BRi
pMLAy9qsnE0sonN2BUvy9CyTUGWWvX+z9d3Py4PZC64GlgtO8QP+us5CK1dOPqgNS4g/2hLtIIci
vgaiFzEul3Hr9dF5Z6y6wfV4KzlsFCTtMZSA27TLOkg/gRjOg2bWBw541+YwFkCtl6SFK/OR8x5l
fPtIZFglpREqBD6hEeYyk4yJSUMA8lC32X3CCokLHmi9DreZB76xtGMervN5y3oe0iD0z7eFngpM
Xnu+OhXQrSRWNo2H7BfOHOEO5amDLXjSaj9VgmN/3gRC2ZRTw4BS+IGIVy742ICxaoG8uPxcg6jo
6SwmE86ZgCVJPoz9TdTxKT085dYFbINP7aTP8xWWCf5lDF+iLkG1gE7ANGtQNQKdArxwermbZT0f
SkPV53OgVzzlaFwWZNN2Mqz2+cB5r6gWX4Cs6FYUaCvL+afokePHfjm+5HPpOEpBI999zndZcTob
8RtkNaulEIHb5bjqSjftPuh4ReoBUkxRhXuQma6Rp3RljEqSNk1qvPcVhhsxPFBUrzgE/B5qO/tY
yTHd1Eo3irORP65xejVK7QWSiuvkic/UdJV3Qr4qsgOa+Vk8PHShDmt1uJNRXHNG59RMNfKAJIoE
qxp3QJjfvOlwrXJvbFo64blv8kAqCfRH9LL1V2jUSlCngyVvXrGUewU/T99dZeJ0brZe8yz3LTmB
2Hk7iX3KGQ4vXxJVhwT0nARya420xCOO/aGvx3jI1PBbEwwRfey2RTlSbqnJ7FFhZ3Vs1GNn4NjS
OC/RDYJGymdBa6OP555eTn7g+OtGPsuWoOod/Hxx5ViyEFyBoup1IjTW27SnZRM9MA6tZhi94czC
WTub6hmjWw2VbaPZq7qomLHpEnN7X59NmCSbqcmM10dVn5Yv/ffhMVkjCbRBtd9L9nJZAprmq5iZ
Ii5BtPX0YNKdTZ9Wa2KBzWLzVZu6Mh/2dEyFr5t/zZalfzzR35qsdjH619cKSnDAYwKm4rOeE+C2
2VfD9RfPjSz6tnZQyF7Mgx41HxolyJH03XLV8m7Oh4nJj3zDdUwFD4TOswVpBddqNH9e1Bp3sNmR
RwP/CX2HniiwsAslySc+agohCoajUyAaSHJoJgem6NwfgLHpIMYDJXw4xvNFVxWaio+o3ZSjiF9/
RhjmRylnfOmnK9L1P85DoREVC/X4b+Nl/rxtfmuN+dXutWWKl68+kacYYgqnHxw7i26YUHWCCk9r
1aW727/ywzCCQZNOllWNweG1V8TCt9Nf1U/dmaChq8sq54XCQL9xtD4FpA/baQmyC/XBhUwoPeYc
1rxli1xLZoKfSr78CModEyZq9MswmVAPo/djvQM0oMJw4ILT5s5VyHHWC65oJLTjOp+P6fDoGy6r
WJxe8f+EAIchcc3RsiILbOuXPrbwAeW+Xl7FpXMYxFqLpUjIUeVvYV/aSudCxX9vM23KquZEhpXK
ah42SJH0O+cIW3pDmmNtoZfwXEng6QiLNKEUI/tQ2/sAb22Ze5JyALrcrnieqDzPbLeLDvE2dMcG
3GziOKx256hpK3slg7em6DwxqibaKs7uz1msMmklgwrnhFaGaiL5iltTT4qm4KjykLLeAJQlhUdu
oGhSsc/0cf3gUnzB3BeLab48aPKlD2+CDaS34NRJPDp3NmqaPqe8Hm90qelOMDIMnYUpFfCTGhJS
5+Br1zWop5vxiz6ZSQcbd1P7LSXOpIwu51VT0EF6dr3AKgrOACU3P1ttWxkI8BepnFlDdyqdOcwd
QwVAvXQ0cLWkkx+U/4DfbT34hwK3oYF3RsNjg/zpZ4N4UIq3tN1n90CNrF6zsSp3jc7sPCW7+qSb
7RbbvQtzC2BNNU45eX9wEoKrSklJ4pjboF3g3ctVpW7IzPvGx2uqa7dYZk+bto28dL6HXsdOxuFi
HbOz1oS0Yl3XqJRkHUAY7nYPPO5bMZfLdGMLP+t5GIJA6AxZ4H7S2X9pQ+FXxsv5bs2KSMgw75hG
lsmg520KPlPth04TUgwY5Syxf8veTFe4OZ7YGqXF7qHfSODNMCTZK7oygHGx2jLRPs5m6DlqgvRI
cWLlv5Ita4eXY5fLWO2aiv92iTWK/PRtMVqGWMI3ebaq82NdDcCxg3PuA4wbZv/gh5dRNw013mdx
xcV0EwyG4DI0Ihqv0EYDJfNJgJEYgfxV3CVo+xNgoLzUadK/V+Da/bKz0CizMmen7lpStCmdJKwW
QH3Y3MPzPhiZcjCPBsrrXpx0JIyEppX22bnoAqFLbemBrqXLB1f0H3qK3ZlYbfgDoempI5vkRgWJ
aogkdab6U4IZcYq8D4tDJ0/O0gKZFFzXVYJgDhbY9Y7dtL75lp29uxVK3w2+hwpOqeob/G8VPlpl
QrE/sHzIfsAk+VzBlp7rkeT3vcN+KIA5DtZOg1MH1MBZCL2XWX+h6hI8+8KStviqqUdWlGXVRG3o
WysxPjeoceqx9dkpkpifRXqgFxBGFWpUNtAvhhOLRENQacOwzqpPYZKemYJ4+ZCb1xtLzd68AFtz
8MeqP9mMJfX4pT3VRP3IaiiDxt/9wiaHGsVykKzcB5XtBpUmiNhKOV6v3qDZ+PNwpcG+Ab9W9CXj
CzVscXEndoVKqDtrWyVB3/7QYolOBAf5JEOuUhhUqGpXfbjttrM3D+u07Y81qqsBAxtGNs91Iozs
4uNMSeRSpgGYJPjOIq6zX8hcQuXeq1EBgYoAjXD7H489WQt+TmmHem7GOc4fZc7pQtHlTpwZpEps
jTXxi1tuSCZ56PLTpDg6zGFYhknaI0A5Kq5zTYUSZXRJOwArP4/+xGtL9y9W9Ef6nRX7lMcauhIK
DxbKuBH2ZEdBDQJR45g9iybUNjHBJmdBnUMeAOP60VC0I0jIwZTExmX2hzHC7um5ZqjfCUeWlKQ5
igASU/hR0yUn7yYxsjDQdhxX3n5cuZhgI13RzRBZKM177oSLLmWcTFsls9cEtLdHzkyE3WiHlGii
DFSPJtmu97EBLJsX3i7jvz1yUKXcpy4LO7LsWE8aFeyKyZrRCz5xQPQk8yIdncJnzsGUaGBs+Yg0
OYHGXcZz0p3UmoW9xSgb76GMWR8zm9jtfy6BmB+ZEs9M3timtwtMfq7INVDznNXlp5F2vuSPE+Sl
XSw63T0I7xdvy1H6GbhOnwrNtZEQYOXWGFzBjKmBr5cSlbLB68vvad0frk8vABBmbKjh2jCUFyWC
33BxLRpeVBgYg1gf+IBV20qzmBSGIybiVoXfunkyMYcLANjf+e759jsM+kCPIw0sT7+n2kooGERc
J+eMgw9egxg5iv1zlQJ6v2JYgxWNB/NXQCPYuRn3bIq+e9IBaJ3EAlcIxMS24LHUX4cBnKhjVETO
RMI9LiQG5ROk6vLaCrwuRfC5H1gtz30ele9QRelsfoCA8W2OO8qKdUwS/+6Viv7xxNKFfonBpfJK
wzGmniwO2o37NDBrDOdUYjYRl59zAecTGJ84+mPzGh3mZ9Ho/DXwR0tw3ziaK9yNQPX+HgryDBWg
9a4bgpDCtA+lADnUmzkleCB7UdbcqYtQNzgncuKoO6Eyaj+TzWTLqq0RyGqJP7ot9wTbQ8PprUYY
VSVxWGDQBnE6EQGlRkYwuTegaZ1QtjYEnlCYcb+WMvkRLIUQ3BURCxZqV8DK2WeZdscCx1WaUDJb
55itTviIIxU/lo2pjmSI1hS7iQZECrHA3Bwfgkw1POAwKw9ydLajfbOn+8buu9jJrDKe8ZhbJjsv
C8aEs5xbROsDj+S0FCWhjUID0rN+yUvxcvXNS8OJ5P6aso9QmrAM/jN+6RaUhpc6YybgnfrcQzEc
bU2IcMAjW2LqvVSN2RgGzFcmKD0HN3dIposaP6azpcWwt4EgffJ/fun0MgREwQCKBQLTaMmbpCpR
Ngn598TGDvr/eSa3yFDM2ZvfJuxacRYquEBP4KZloKxlXokMThy20HNJYhH+VTjhbcGmxrS4rAkF
yxtEmkIUyUa5KV1ZHuxQkJ/gY/cxWmzDDZuqkB/IMZFWDYVAeRl10+0YdkVdOcXu8Ra0EkimRTO0
t9XhkcmEyZI9JLA0g/TjNAMM14Z8q2D7wQoZeu9W7Yp/zFuN170aS5wbcyT8YHdf7qqXkRDG3x76
3XG5VI50HvupJZ0D7+692lHYhV8XfFHCkoeMqUhNCgTuicCPcUY1hBvucXhVCpBv9npl5zC/Ayyb
fph0xJT8GSWOE1yRbXqFasa4faKak4AiipzJs9Yrt10prS1w7H+f+THpa3TYX6TotDGwSYO1dO3a
tkoU93NaV4gPPVYLdsgHB282eEd0UDjHdis4ARrnMvHAFapzySV/J1txlTzSE24Ssv6zDE+HxncJ
l6OhnnppDSrMOxcpU+2++srYaDDIuZMJWwe/Nz6Z2a7TsxvZM6QYRo6DxYODOti98podHjY/irFj
ocx16t1cUp5mfKyj07+YDF+mZS5lWS+0/mNqvzGe9J1njRMZsmGgDtoQ/aALaVVyp92wwd+UIT3z
jOYJc9WU4hC84wzNBuCJkD3bv8OjcvLvBmaWMJ+Hdc8a5NSffAQBa4+hdgUu2AOEJ2Z1A+0w3kwj
mhQXMK1jbW178b5qNJpZuMcJZzwb40MrjkwpD66AOnhx6V+JbcFpEPjD/Cbm9mpBAfURAFcgcuEQ
bLpvi/IHnUZPfToq07tr7xaWRio8tVbWry72MTdKHMsDSHMNiYp1Wdr3zQZ0SL+H4fgTm6q2E9Ax
oGiDK17S1yE5hnvrldBwFRUDg1oEeOd0ADYudSTo/Rss2Y7exKf9qnc9yo3Ski/nVCitZElubPPQ
FEgELCXXQyhs1aGbcBWKOKcBIo20en7Hg2zfzunNJ99MahCRVP8v4f/fKU6on+r5Qk072k6LgQrj
s+ItnCmIKAZfseBK/UJO0rYa+UmRUWiRj0rC3nBU+dLpzYYde2ghawjYw9zKnQQS+Pbzz/vKd6sb
fuuON0+4pRUQ39ha3gaVMaEw/dO9SZkoZvsgw5jqH2WTlLtCpg/Dx7KqPZN6bizaCdYluYAIaGYX
qSJdfK+4O9uKFKC5iXeFl02Dj8tOvcraJozkhJB+UtqCO2f18aSVOLPOiBnfpRb2j+hI54qQeg1R
TeTe3fAqPZoxTjGvDDpMctKVXgWl6lnULKHqze6+HoIs5miQ5dDDutM1OcFYpq42rH7SDrXTx2+K
oB80T+qHQobE5H0LBioQKVnfykc9p5nIe9SqZkEq33QpWkmM2DQHXgcUViqBxnNqHrUvTBitRlKp
AhgCBJrzFCyhIui0T6vGU89UfsAxjG49r+A3dzx1+mFFcKkB/JlpvKP6cy0hFZd88m5sNeXy91Xt
Wx1w1g3EUjaCXV2sB8o4PfdEtySh4jJTILr8L50uSYyCWbdtRfKUd2gKTWn7MUzXmgr9KbYNfljC
UlvUEGW5IWTEEqe72JzLhgs4AoVE5rmGj8smaAQwUR5qxO9iVYTwRpZ7JLvz8dIvGcsTOVdZH1nv
nSTfvxa9uw5JQMfK+fyQ3I6qgNelHf/JJH0xJBSooMPyaE/M2+8gOhEden5v4ahhbY3uiSRezE8V
N15UecCvyACmf4AeneGt4mp8Uf5HvjkmH5Xa0GfrzXzBQDsdOgZC+JlEqLMt5aIf/6MazozH2Cw7
45pZDEPClUqFhYdV8oDahyGgUhhXRuZapw4SOh++P1vouFS/9Rg1SzoHQd1zSbUKkU0dv5J7Stbx
zXto8XmifxVz8FNodvIoq1E2SbrcaQqCZr1cekJx4KZjuBNAOLKziy/ETZTHTV5/+s5ovSc48nYg
af+6EreWimsXdRWeS6aNpXYF3+39d/BO2SL52Nhabi40oetg7qyp+QC+KL0ph7mIslJdU+zVOFdu
3TaX68hXKmIVB6naX7rIEOZiQEKM0tnF5mb2R3f36PjD6gtiLmBO+3OxqzglRknOUACl18fo1yl7
4H28o+L/0ebVLS0ch3A5RY1MCqmMPbqZ2P6QC+v/bfgUc+zNepNh9LDvfZda90g4F6V8wNcQJScA
et4SxjaaGRfXpeKkMs/0Py0T0grwbtB1DuHCq7hX0NLVqPbFKHURQXmZqLW4phr3Qd4hXywfoz9y
Sd5ZxtKctLZ30YY8WkK9THNHnRDiOquK4x9UwguPHGIUH4ZS6EPIijoyMZYxDd5g+y1nJlVMxkgx
eyOShAi1I6MTMlaeqbzH6FWukD+NTmqRh0fqFvIaPTXd3GrN7MgsWzT5Zcnt/3wiFUV7hpFRPwQx
hqOswuXWv6GzAPMdcG29HO+9LfiBicsNUXjv9k2agyjiNol0qwIJT2vMJb3HPgAIVzkBPOUPmBo+
XBfF3xtxNXkpKNhOsz8IJBQ8MYyhG8+iMsGvmV0I9mizl3p/DZd7aJeSGO6bNsn8ZTWVd+EQ+4wu
5eWHPngkZOIASTdv0jChnAI7vTX9VEyQLM3fdcd3J9WxHvA1A9cr9F7ovWzyHy0Gv+3EBhLmKVoc
nb3t6hWS1jlYbqiBry3i4wWyq2/0xJ1rSF5jbqMECofa7nXJo3FFBNDldOadOdpKdET8HFsj/duc
fLgn0a2Uwz8q4Os6aeD+pdcYn/uNOkT8iEchZz+AsOj2qWIQ3mJh7sR0a6zyOevufwO9puYMHrf/
kccGSr12BLxNP95z93AUJDkHRYOn2qeKnjvSINAtR7+VD6j5Ha/uYhTiA650Jo3q7EPQluSiR4hq
X87eLlcqkRoagiTZ/iRnHdFyquA4wjjvhox91DyEE0ivYss8OoluCb0aS853lMq/zb+9f6af57vg
Oncqp5tUH7zL2FKjfweN5F0/50WKwhsakK3whSiG208lHXs5rlJ0msF5Eq9JWR7IidB12KeETDoP
gYAnrWv/S0VJBE2I8Y+h4rlj0000z4V5+dgTgTt2dOpJD00oFqAkIaQ8M7kDevsEoYoJOQ22oF9t
YzSrrBBmcyflo8f3fAreTL17dITQicczoYCmeDl6Jt3SeRJRqOMebI+5zq8yCk0YYjCW5hbv8Bze
I+a866XGAPEhQn46XBrZy5kbeImg42BTFPyiQsFbQ1O4cv9RQVyuLHnMJOkYLJEx7NUFiMR1xt8Q
G6a7vhjZMwYwerL9zfQxRZCm7NqzH37Zk1Wdk8Q7TYiZYg9MicGlO29vjJEJLZOar6KW+zkmbH7w
EApj87BhJxTPdnoz6PnLWDJzvxnebRukSpkk21h/C7svUHDOMfb+Diyhtuy+i3YPdI2LhFL9MfmU
tlHL0Naprh8RP+fsoZiWtBO8qpEbGtdvf5zaNZed9f+Jt0zlnzmT62rkEkZMB4nAUXUlziPdozeR
p+oM1tEMOYxx1KnzIOmNQHDAVGqGmR1nv6SxpwGoiN+BDkTWDZwdr7EtZqXHkRrGzsLien8Uom6o
zv9UoeKpnQ0K36nLASGZFMlS+pteT/Hw0LlDAMxeFS1KYue24Q9ozQWxP6Bdv0ocGjZgIpI9abEW
LsddyPWH5V2srblTSD7b5oEqKoFsf/WMRQ38J3akCjnZzRHZYfi541INdXWdoDCW7N6EMi2ib3ln
WiGySfcFnDWuhtnZzqx/epUxazbxN1Hcb/CYePJTqyhxsUeQMik5XttL7+e6z50S75B5FUYyr1wE
5bwcCwMGyoBXPUqIEU+aV3uA9KlSfMW1EF2NggQeehvXU2g/0Ke3ob5rAa4rMbwgxV5x2qQEhQ9W
Nj47a+6sdolSJV2hz1ZeZ0vRJVmR5KLOYTXmwLoZ+F/cV0GrcAjQxovkC9taZAB60PE0pUAA+mu+
6Q8ObuZAH5b+V3wHiGIkbAUHkkbSYl7PHrfUbZLvwectyfPtbe4UkSgoIuXENgBlOJ7F1XPbFH9W
LNgKA0YUIY96tceYUNe0PPur31XomAWrie+72Z7f1MqS9MMBDgSzDmap6tdSCHnlVnT2YzlkE4+l
3Kdmm9ocumnQfzgmekT6AryCMNmd0a0IJHZOdB/+kKPobNektTG0fzAREEFJPdaYVOsWBEkJF07x
/HKFj5lGreOo0alJASJ+t3EBLn6KUY2v8bmbW5l+pjqxnkbqbsw70q52oT/6uu66pbbq4ev5ibaf
Ir6LrKDAh7meCJMF4Uk/EQXZKkas2EkYlFXl+Fh7HzeEZn+aP1hXU2ofUulQzUGrC9CySRqdrzQ8
tveVYxbGo37Qi3L3p9MEFP3Hgc3bqJc+Fjhqne8i9A0UOOBMOYNj/BVmCFKv8Rp2M06k5dh8Y6s1
Qr0WxQDrYDIzngIoiFSzcWHrcCDFzLvW1dc1Cdyy1G/kqDUi7rGzoMi8BRafGCeUrI6n6Ndi1Pqw
XMxAvLkkuCv2WHGOEhVZI6LSjzxLSRPgNyz9zyHBIh+sOVGTxkvvkVMQ8z/K9LHRd2W3mwTFOxtV
rrbbC/xlgQFZk76vFHuZSjshYkQ8kQnWqzIxF3SreN3en8dEzRPyl+50IGfV5OxW25/2CP7TD+gV
avKTm8/6bMo4DXJs3uDmtOMtxlfc0SSHfWHlCnC/VAobF9jIj1Ycy7/nyHTINec0B99EhoCzbB+Y
t8Dfj/8UJTJS8sUgnVziv/1fzjd5fwJRLng1qYOPkojpnAeZTlVm7HRr7exa7GWa6SWPfZOldEz5
MCjr2EV9quJBjauX0aZaggjg5HeGOPQacfwauEU+4WnEhM03KcHbb2cR4awVLgArxGvznKOYFOhF
S3fMB5sc0SwJlFdoXx3rXNqTkZPeJmqUMFf2eYIlexTg8h9mHUgy6HUXSF8Z/LovO8DgGNePBq/0
d1EwccVH57GHNpr9G3SEswsNEUBQLvcTegaXdjg5pd5RXgGz09vKdReyDShmfGe58+2+0k8Oad1n
eRe5n2Qzkd6/4HS5K4Jsx3JDqsEhj42+U5nvfTtWOzdcGXz3Rz2xwoueIBt3gNe464Gs8CenBFon
hS8Viu5WW2hl5s2G7Q5mouDZDmwR8VeFWulFMfTxsJ35RTv39bOVWoe9d6hV00/NIMEydaAzHGxY
SzOU2bYOlTHGTBv5tXmiTGaZLZkx+CsuSVik6jUYiPROJIQmdVuRF4TmUoV/ImnyKW61+L3kqPA4
sBOxpM1nGS6aNuidjQe7XEdsvupm4RHlU6n6rBuj+YA4WUMbe+4mt3qEfy+BAvJ7ElEajvzIrA8n
BSbKR6j/mTx9hQ81GD2mERSW9OsJb2asLqBuoJ7tdAlyfUSGI4BzVJf6AJIgSommEZ+/FCx3SEqv
n+UTZvfHofyk4EYpSDGpuyumGXapms0ZQwdkiPABSVC6dRSNSL6E1TYyCsiMDqirsZkXT9isJh1S
DLaEL23+QIfG2rLvT66qJY7g2xzJHxBmth7Qm7qvFLJnv9TGlS8bE2sDlDzk/Wt0a+z2a+nS7jwx
cFs0C5KdKo3xmEF21BbMAKb7XZ5RupusyPhA41bJmieUw+1AzJSO1HEy8ozoX7taW9JYXu/qmhOo
pxn+b6E7CH8DucmCe3hMZJXwoPagW7xw3EnSPkHHi3cvEPGGlh1Cjua/zrnhfpGV1vLSlQ1nHZh6
MmLS5Frk7y6uUZbN9vEviygHV/mVquQlzwqwEfsPhbq+SIoNQujoyAy2lVg9VAVnRWElh/egR13j
XMaGcaH/cmygyU7eRpk0yT8FNnmgIHht+7tU17wHpqE5r+QHq3CBpM4LNIW8fnW8KufkyHZMQUO0
2xRaIn8bkLfKo6GMb8uVC0vZ8k+UgutH8OyuMXKg/N9J0iXimb3bbqStS8nQM+ydXDnc7qwsDcBy
oUu1eZKNSI1zNQv4YpJ/9jOpWgNlqAL9/CA40t4px0Bcm+EjiMrVeRpqvSOkWa/whE1dPJLbVA9g
FHK3y/XXZPJ1/WjYTJhaEmJXXVm2+Vk2fmF5yGCgB/ogR8tGbax8rWNmBR24wqxvLcxHCj8ue3wK
HSvpw8zIPjIGiDCDML4/0/JvaTzbVo18L+RMeZlbkBwFGdl0GBYHc1kf6B5i69XgiVTO4nyOGlh/
nkr/kE2P2q83oE/f7ff/fbk0YDG5L1frIY/eIo3NR0eA9v+g4H06RqJqtTCuJOlAlG9xHeFT6GPf
vFoqfCoF4tk/ynC2hccY7UmykJtJWYds83v8VzD/d6ciMUwvIhVbnIBBiXocH69yQoOoBgX8lsm/
YIQl/MAl3WsexlB982BJ6KJ4Lk+hdAOihCkZytd4m/r2hpqXS2HMhQ1IluoAJDlb2oh5lQwQd2lE
HQBOkr1P3JYToyg6fK0r6Vd9rCmBrsYw8TzBaJK8dKD84AMxOFhMkStdZdgqFHJWQo0MR8OO22NO
EGP/8KbulgYuR/jkVpAXNKGPjo/w2KfDOzGXa64aOmBJUryXvagRwY8VA//9hf6SHUqZglxIkbo5
epRBOp3nXBjzQOxu+2PXysIwTmzgVNrZ7j+QJjiYrRrsFYK7L16MgvUzCJrBlBYkOO47t3jcdzXV
W6K+mjV7zUfbbEg4HO0u+tfUKcNexJ4dvvDIK9X0VBUEFc+L0SSRs4LU9yTUN0lozSADvcipjFZ3
DOQOMgKMKXg1Y4oCSN9W2tcrmBhnxOaFSlBQjvU91KtLr6rSaU/ZMzVp7N8imS9W/zbYhUouswdR
fyrjEkheqY3Cew8Mth6XGW7/3Nf4kj5dcSX4xQ6NopoZJnJnUlUcPqYHOKC328UvCXv1PXund78+
aR/8yXXuPNB/pDE6Rx8e3hU6hjvjvuN+MC+7DLvHjGycNM6aa2le7a9FC2X3S6bDP2PDybsiSUdw
TaQ/Lr2/IVKrVNoCA0KY39BbBTURxRLeZZFk+lfUgzCcM87hHmG+2FFBjL+VD/Abvb9AKQ1C2aoJ
NvKD2TvRsVomIi2zhAIdehI7PDhJX0w5NLaaDkmUy6OKpwEGnuTmU9d4goMEnPRhn0O0ky7faE08
LUFX18YlfcgwkgGWkQtJXVqU1PA3rEROtQr3KOa1t9GkmLs7KxRFuoRkoqwgv9pAIjXtFx2I1SH6
DC0zVD1cGJGgOitT3VgtUGmcodkU7ymGtfJBy6C6SGKSLCKBu92zI4+xEtE64wF8a5v8cUAOKr3t
RgW/jKWBlZVZE/lWnxGjsOJw6cTO1BoT8+v1nNz2g/4oqmLe69EQDQrQpwtJSSCDpF0X/bjUuffy
yOfftfpMkxa0Ux4PourIAkNuOcINYJSFlD2Q2ahnxO3mqKlWs401Pamo3IcS/Di0GiCX0B0qlNAX
KMM59zMwsezf9jiJzSu32REwR87raV5yxgSGwLz+XlymhvT4aWJe1cOHQjnqJo5i962KN4aI5wGp
EpmDzb3AbnlBJDOzIW3WOdnvgI9Yukr0BiXZ1ARz2RE6NxW7P0eUqFMwe55dZ9gOTzKEzUdsw0Xm
jJiMG70HdQL8O9sSk+RUEWfTw0bGnqvA+e+LV5R7df5jmyUBb7CnPayIDJoEiTnXOpQWN+a3JWuN
0V4x3L+frS1mMo5I8UjSobGZDzTFZgZw+He4yogNSa9bpujcyZQ8fVAt2OtpBPqIX1Pc8WR5YsVp
tspV++TxVsoaJPxgLbrzeCDKUYGW8Gidpm5UJEvDTs7g0WvQ8l5YqY7EcDvm5mrbvmy5pi1e1aT1
+xkijNuXUceF81CjF6JOsIYfrp0/Z+grKDglZrAQzNoEzV0EiopRx635mXnaQErGZQ3wFPESRxLF
OnhfVujdTrccssuqCi26i0HTye+8kadbQgsLFBy8eGlwDVeBnYOJoeoO2J1TksI0EA/s1L764dyM
JPiAQfXJaehxwkqfO0g+jjvZvO3Fo2t3uLbeOt3MFKDrjq0/+fqvoWgoIKEb1f/gM96FkNZPzVOj
m1Fsq9dIYb/OrQ7xHLD5H03tWbdT2kmCCi/xXejnGeK3EhZptssKoqmnVQ66EY2vNqeVMpyT4QBJ
GArPnIjpRoEh5NRaJwo/EEjyF0tnKVbbR5VWOjvpSOyzArsNVnurgt+xQv59Jug207FcNg1NcWjW
yGs1yg2f/3kLn7+VSR8tdUf6J1okyrVdZqRHrtZvXKfYnRyqqe8haDtlTU8YG0D47i505Q+Wu2Gb
M4XQQvS0C4YkkLP8gt8wXYqSYeT++3g51xHIn+iK2IBhR+VpeJ4Bw34sFz9U+WMJtIzy3ffySnBN
XDt/iPVn5VTtL8ZEeMQMX6XetEMvocjwGys6sFxLpgkxuITtaJadCN+KGTUTxOllHuM0MUJv1HGH
wXH7DuLXrXjgLDN7swzWRXS57YEzd+ivEHannF+KDBq+5EuiAygzIPwayKVIoxIhySEFUNkq9b8D
wujBjo7yeghDmulzuXEZYJnkWWk8EGhh50/inFbtmTrgrxZ7G7dN1CbykwiQt6EMXDskCmMN6HVB
rZ8nkGDeilSuh2byRCBRNMGgXTn6t4zPCD5D8MmUAuOSP26B4KgZoHuROOB4c2rWog9R5ala1ShA
NamBADy1ryPwE7ygaPUFYrluNFftkxKiOAmjGXJQpmpzpUWnqmkKA45LZigGfUFQohPClunHsfEB
F5VbskqL3oR6GkL+j/+FQZp2K8HKLYfjT1hEtABqhmTp/sNSmnJtVa3d4hen1sJEkDUqGF+x942w
2NwajiEJU+oMClBLuMWetW9eMXbXLuGEeHUUbcFVRXx/4/pfxzQqhLRpB7AsAelPQ2wwS/qy8wDd
Wdxo+fsaPxGkeoQ+EZig3z1QsfE/BmDt2c2QQMV6PYjDlKAjRcbNRWyF+mkWGMivtT+21/c+qtie
iPYrz43b2ev2VNFS6m7ZNWU+ttuicJ0g2BpJ/P5fFFdVBG6RrX1gbwmtfO2kTE+4D73b4YhmrjdS
+LdxtdKnXIBfuTF1bwxgUlFNJ0mCAEGZK5rud9YbZV5QHa0SKkGQVjcRfy2nwJi4uweNc3QOpImL
R+Bl3qhdvrbywBQdJzY4rel6TLe1Zzo1bA0DvH887CRXXSE/68HLvo9FQPJYfBDj0dRh/KkMs1+6
ywvq+p8JqyO/TzAFnH/Q6pIIPCwE58PGK86oj9H3hO3PWdoT4JkD/UIxeEg9BB4pLISaPxMQpj01
qcnKDGYOlpjMO+7FDb9iMwyhCpWfIlJDEVCOIPiOFEfEEGvk10nmOt/dzWsvquoBBCdm+k8CxiFx
wNvbyFD0owDvvVo7wZM3jX6RD4nbZoQLaq11hF3A3lT/lftVxHUiBogg04tkuud9vB/y5qEP8PRx
KNTOrEWJn7hdXd3pXXonqCUgDztTzTP1Mc/w+DUsqY/x9Y/s1SFFdLQCjaZzOCVZe9sgRLvC1EDH
ZPaERn/+4xvzW9VqGOQovswrEjba9kDL65EXL+oIVUg87MXd3MEKQM6WSZWh7JKahdNCspmFMyOQ
SWJ0XzRWaRPItwHQo8QPgdwnfpOPrM4oPkN8H9rFszVfodcKfk3nCNvGvqsDmcxVSwfhvcLL9BCr
YCtSRPUjnj3U+6aECvwDYghHKvQhs0fwXK2SRln7Rtl6Jkxq3a8KBeSXbzoH72P73D6iAk+kksko
AJS4sjuPxbagPqZ799tjSntLLgk+FaMJsHrB2gn/mnRtM3ZsaF84g0UJ39laUhk6F45BzbWKNA/7
UNV9+E3OeUQkIeRbxHkU/A1zGFdQnk5Rcg87Ey2gY7O8Pa+1W1pdVavdwUTyZXPkTGlffpDo9Ek1
ekpDi3CJo1X4/lp+Sopj+XNHeoGWNGw5l/hPyht/0Y8sygqGTn9b4l6ChsrspYaqt+oSE5iIUaTk
YqBAh0JecLTs4GPke4prlQS83rw6oFAs0rsEanhsKZ74Q/64ALinzZyU5corvaZFlUhQBuoVbgrq
s67PQxmB3Mu37oi9pFJFcMY/FOSBDaADpgpCegyNygDP9WgGulj2IbrvPDdh6IzNQvY2GVvGjHNy
riQkJNSy+5IHgVtq2OWK1FCJP4fFCHRzp01CjYDYSgEc8RxXkCf+ks9KWdVlTMUOw8ccFSxd1Byz
KxcDQyV0Zm5K5C4AFO5SgtoQGUSAVZOBBgN3lZuDLG1Zg9snRicnGd9OUjWdzAKbPGrGTo9XlLkI
RNAf2DzqxeVPS3dVxnRg3PEljkpDqYlVHdkm6abr3gGANV2JC6zuu9zrczWT8a/mXDxYA0KkX/Eb
iNZUdNmE+riSf4m27OnK+Lx0NxJO62DeihcqQW6O/Y4T/ZbPteyIa5p8xLCTiLkF1Wb2UnwAXCbn
SBY0YhLP/knN1RuzAlz0K0WyZRQO2MqB4Dil8o/Dj6mhCMPI6oAG6nmg92dAeZ7iUueB0VBV5rZ/
RCtW5Mj+IJojO3Ist+reZ4hqiqWBMQlZnAHOzGYjyN8ra0j4eIOwvns245nB7XuQP02buhJxGS+3
zXHvs+yw7C4un9beGhGuITXXw4BBllmMgr0AUwFKVBLfW1Jur9j1fe3BzSxmtDSlGmVL5Oc4v+KB
IaLTlPtZuKOEaKhh6MRfB9j2RrbtqqUSRkYm/1BEx4L6HrTXS9K0H85hiUIwEeG/s2PNJt4V9zUS
OBZhLWCJwbDgPdWeakE9zVmGSEquHV4s/eqdMA9GzM6mnk/ZxpBoYiA8KKrfXzKhPA5/tUmEnxRh
LGQr3pT340grJg8AVQeppI+hIGH+tOj09UJfZstPNsWniLKD6QZk0ItVi9dPuKNToVBlVz7o0uKz
/vZLqz5KE07d3M1vOiRwR1+E7Ficor3jYNd47eSzUjm1JNOgRd4S2t927gqrk0J3jbiD5OBmFIRL
Q61LhQ0K+LY3aPoxAknSWzjwpJ5GY07Ubh/Qa3DPYumTZz41vW1LflE/KjQoPo9lmfvqH2Z78lBL
Bz0Ntfo9Ni9uhDpT96rwxgRiBalqucV4P5zd3Y478ZaqlAd/e/kXKCp2MV6b3/qIhRVZCuKNEAGZ
BN5p0Hs2zWP6mXycK6SR9asqvBKTy5vUJXJZFAzDwyHdtKhbMzNGhmzuCNtpoKPFh8H2Cglc27JO
w91NunG/7gEl7sy0lDihoUmEBrmszXsvq0XkZ27/Ux4LCwfQF6Vagj6oyUTPiq59GTkxULe3HJyq
RmCRVxiCU8SrI2FNXuWAiaXiNhQ8kot9Z/FNbfvESbypH1Ex3Fpbxq1s8PRwYsL3qeWx1cVSwEnx
pegoNpLLA0YjfcZsYmYPDQeeactfVYY1kBMKzH3AEcNm92qIKPWuipaCZQCmr0cb0M8SXRE7SHq5
qPfrgLo7gbx9GsfENW6kf73K4kyFMKDgbEwG9tRRT6hcRf6tglwGXwXLrptf+sKwGGCFEq/dmFHu
Kw0fsE/ymJ5iola8FqQsqDb5WHJmTSjc/eYfv7W6wqgpTnXuilSmaXNsQmuyM1nB+f4/6s7cFP+W
1KuWVAy0Nlera94/oCORtaYDoXU1YF9T31dRABGVSGbi/nvzfs1w//T/nZK+14nAHaQbLrqwO47N
zcGzARnp0tg5Fq2xq4kJqVSXtcNhAHYuo9qJp5XxYzmzyiq9eyM83SaCpObiJ3vU8oDqoWzx9fY5
37XADjXGFg4fA4RRYQnoGkYOZr/JJee2k8/UxXeXhc2SO1neL/LfR7dUZziK6t3HvfKnR/pwoVZ2
FXmvTixtCVEy/iL8xlOBl1YLQcsbpnvh1CXM9PP6ZnRZOilxmyGQyQTbDfXF0H4FgjrY2sGSQBKx
kdk8qdTO4f0zfYeZUKTtRHC5kP5I9EmwmnPqeMtRoCQNAgWKS11hUZX3Y0ojvdH/V2A2wOY5nWgR
KECAQp89UH0yqM1Wlf95GaGK/qh58gTy8sYO2nOwm4x4SrdoN5Aqp5boq48KkjNZcyNAMzWTvsGX
iLGf7JSR/ePegopcpV8EIPsIbe5ekt3OStFpVTLBImrdueTPCMK1rFBJNf5Ee8rwHMhtcYQhSHVg
Hna5HW/jhTpvBJMYUgXRPhs+DvVIjBnXHbStcnRB9DcxDoYGwQz8kXNwp4RJNBKfPnLXgt5Fh0Oi
Yy00NaYWI7YPEygIM8ayNtbSSAXEelcQ3fg7icolJDoQDzamD0I4Cn1L0eIa6N8/FABgsYyoSB8e
zFgvWgBZMkJl9V7mH3XeXIHZUYz6nevleh7J8v9l73XAUKQgev6T9bR3x9bmBNlyMpo+mqblcxvz
YH+C9hyYDcel+2/wRPbLMi/H6Gr6eQioww7OtZNDBbVf8Ug2YHWclZia3ssjI9CdakfzYF5V1+oX
q6BUeHZdgJxTZnvYeOIwBWYQU2i2OYbuhWcosBZ9LB4dM+y6/SpKCNzZ/R3DqGvn5drShxPMe1kG
hqiNthI0Wu+ne4IOIhTJe5swQaxlavzVVYU2cGS+JrGvovJr8VURhm0ZrMWCU3mMiiGYqpbVADUF
3fAYKxLrVNowoKyuYqxpdA0Leg57n4eBmhZVbuQ8501ce04c+iLvkjQmaB+YCi7NUvZq9jo1Z0b6
JDX0H03ru/josAqKM+PzYavjQFV9waqVTtP4cscSICLolSTXiEbC/73JKtrnjRccTPZYvvApMXP5
14NDA4bRPoKWZEUwUonfQQPgKTU20tJoBropwioWZ/Oc/yd3Ch5KqggQHIN5Q9J4Ckkqg25hOvWK
t7Vt9LDwpdg6AIe7ACs3l/OCbiZuRG3h/24AfsVIQ4PAMt5KbwC4nrDSxAc7ln+W+qAZW6OJc1/G
ne037xEn5jCEje+pQTXX0Z0pArEqHt67lOl1cRYeb7tX7l4ACdk+Ae2e38pHWgOW8Q2xhyBRAvjQ
Hn6Tsbub3bbaXfecJt6j/nUmXLUbuOzEOhpmskhiroQFG49X4c7jqBAEuW8Jjct1zRaY/telhkAz
gqkqht5aEMt4HEufsWJjNZd2z3xxRJghkGEnr1G/R0KlB2UPH5/Av49y5H7Q4xrwYpnPEK/Zm/Ry
EY6aOpM+9C7tP+sGEQ+PJPO6Ozjy+juGKEds6YFTv5gE272u8NojOwC8hbkzNl1vzphmRxwSSG8u
vePlbG2OtNMDRlhuB9EuHZVgvsjS741LIR+EbhkyiyW1DG86mvHOv3rGFPaKr8ZAZZcs/rqh5aZd
58EHheX1+3xhu8S/xT0rs/M2jUY++06yzYdsnjaR+/z86CmKdMORP/2izj7tkS8vzQXx+5qRhqPK
ARS8l6F1zM0fmaN7KvArYFBaKncqGqL6nQTJJsra38yE1jh+MgmBSsgsofxUc1lyOJKJ5GZlJbH0
oGkJjoMeszfR83G19VcaW5ZGmsIccxc+UjE+MISgDtrF1lMTUttiNL9FTlg+TuvlwMbtX5cYZqr4
rBw7q9/xSZyHiYctdgsN1jbIvsG9bawF39dYsX0skzwi+w8LpLKBKttPiwiRcm8PQDwDbMsCFg2C
ekfvQRSYhM9V5/QiQ7vpkzpMvPFcv9lyaQsoRBTUkfuqHUliGfxumekMKsjF89KDElRvpZKqAzGZ
deBGNyhp/bNOCjT0y9/U7+1e0QkRkqA64RcOpaDkjlmk0WAPBj5crDDS7CoFYbtARQDque6t3S3t
gD3jOfWJ02DqGDS1CAAVHUyp60p0pUt2BSXlkUhCyso0Uvd2uK/e/qowGjMpJa4y1Dfd/Zs1UPKn
zwJJXO7n7so6b3C/bzSJjyYAHds6HwiFzOH1rlzbpUfO9yP/OwgOUN+cnjJrRCfamL+t1A6wtccl
kFp/jteRbyJbXQq7N6phUqsMf2QgtM6t3NoKIrqzqkcxNBKb+Lx6eVHGJwwDdxCdsStpD4PUlPdc
/QShqJttm819W7ERIW+38k7v4GF9N+goBnwMzS/0nFTIUYEAOuuEDYQCYK6GfGXCYc02RPFQ+4cL
cXoEopf4gPibDUpUw8YCJe+6Hy0VT6CLfLvfFYDLyQAQHZ1s4JnovHl/HeRYPfHgR5HKuC1Jcj3j
5q4z4lnZyQDeS+D8ruFsTsKzsPlEglFj2kclli2VrwYWWp+D/BaYiuucbXW/VGJVbXZoz0qs+EKS
9a/+9L3mY8JyXpDJrrxj77PLeeZOHveHZlPgK0y19YhR/XX+mvWcXS3CvZzeWScoIGY3XEF2FXdZ
fE6kmkoyD/c72fd9DCoA7FMVbmOgatmXf8sDAwnJXVnRiQYu3FiD4VCbWJpcq8Fx00BZEQBI+J6z
amd1p2KhIkhKXiKNV6ounCZ6m+igKKnf4dLycaowUHIHAYCs32lnjWH/CmEu/osXikZ/gI7rgBFP
IeM7rkmFbirqKYColEoUrVa+KOli7OF0D4lIp+uP3NgBokfGlHuRQkLnvwqPnADhryl5COW46ivp
CJRiM6NtV7veIH27aer7ZU5VhK1AEY/4uBTP9fpw71fgroP08txFc/9wGLs2VZXlrq7B0x2qD0MP
g+XHmTsTLfF61z6VoSuEbOKej+34hoXGn7mfnW0L/a41rggshTSxwEYpewMjlNUx4yP1Vfrp01yt
BvSTMo47ixxu0CYVIIX7MmMe1/6bPRnuYKOwlh1Y5wywbiU3ZKXsIkMi0+esEnurah6qqpRI1Ny2
w9JN3ICIONYqvMVeiTVWVD5CxHAGUqr1PpKAuJ1Ug5zraWB1xk5aHuCF25IwvMkR/NUfokv2oYre
ZFhqzn+zKPtEKKU3jeRFp7vYZx+Kmr42OjWWdDYMNiV5HQEZVfk/CFRRwpv7PhSTnW426bT2vtv7
vNRFvKc/0WRvRUkB7kIlmy6fNls1RWG4nBs850+7UUpkZUCWPONXl6rzAwcW8/5oevZmYkoRnoWC
xA3kAN7Z0E/dQtG9jJ2Fx+OlcX+ZWtCn6Cz7/quLrvW0yN/j+520pMVIZmOhTq34CNlJyfWKDhbF
yyXDG4Ooy580ZCdZ0CPLWcxQEQaaGlOBtJNv4mUfnYgNm/WBTu7e2yYX536wzEWY5g8eLiH73guq
HT9QD/bmyaRxuR9Khp6ZaipdbyYUO/WPfCVAk1rxHVDlU5DlVQ1tOlL2Opt+faMNIZYWSyvVvqk2
JCH0UUVOuuNaTYNdCrV+P4/BQuYceN21rzvPnBN/zR0yzWR2hd5sQXdM5zY+PxOqcOIHRk4E5YAN
99j0sVV3cQ2tgYUq2dD6GFLwt7Q6ej8II8lSnAcJGWgGpM5WjSijVAvKNWwiJadxbW8eN0r1AzcQ
/IWNVFrpkgsfDSCVNfmylv9JEBTHMczhabEx6sXpB0I3zidreB5K85O3HVKI4ToxFaxku2q+a2BL
4w8MDWu4G005El7JMDtvhQPSreycG4FP3CP9HmjsKA78DFbf9AdFty/8U2wxYL2bXXMayxKUXPlD
mAXsw3eqOQe3pc2zF8SpDQA9Le3hYZF/x6u2I6n36k6JfqqFWkLXFqDqT9r3MZ1+BqMEfk08+SRs
s60pd4hBZQd30w5tuDlcQYXu9tKW/Nwv6k0tnQzeIbZMdInHBNcwJ5JvV7VCAZ8obYkjxkwA8Z3C
5/lwHOw3OYpmbu9AHoBE3ie721IS6hXXXf1ucEWGs2hQRWO7vdWtHkymkyOO8hDK5GLg6rcRu6J2
kxdUhHmowtxQaSCXKTsuAYjZEpe2PqGuNR8e++Eaix42TDdLMdERp6qPkmayjytMZ7Xr93bF6/Dp
tSzZx9uS+jGc9ZS6uWffcatzkVfLi5NtjBV0fMhWlHx9S3l2IZ0O7ZBnodHEk76jHGVBwzj7eLEP
jlF62Pz5kmE74VXp6Dw1u5NcQ8d3KmuzvtiO/MtX1ubl8nPHi/HasRMHl4FP0UwEJav1VkU/Xq9e
DOFei3wg1hWW9TxaTH/NenCERXo1lAFrKWtWQ6H3JTxX9VHAB8pGy4llNTXvRAQYRa4gcUsJilR8
uimeAtMMDdd963GXs+WcsfJQX62iNJg16Lu1X66AOpfrmcWkiVs57w1TUBvY+iuk6BQFRUhy4Zdh
jC/QEaGi0wJPr0kTEiI7tbY1ycTEt8YwEXQPGrn40RBzHbaKBSEfl2ywvo5pq/tmqtK7DHuANORN
RsLScST0Q68AMFn9+0Hj0BGtElwkjz1rNXusi7z+KEdhCClIIQM8H4ZI6IpI8IaOTLDT/HPiXNxl
bBBE2NWDnWdrwlPUNP0I8QViEEzo7V/+aiT/K/jlhFXENWnISq//H+JJVGFvMg9Yo5jLNQA6u0TJ
tJbg2a5zIZQlBhNNwnqJ680+5DZtdOoujOYVyVstgnD8tVlZj3V7jXdHeUez7bahkFNTde5JHLVs
dtUWs4fPQ5IEAG5DRTXnQx52HPpZBh2NPGh4/2/nei4KLuXSCrAqAN8sFcjkA8eebRVXF/7YZmVn
TnMo9AGDkbDz9a7BT4AXu9uPQd1nEb/UALINHlYTbJShCjtS+yu1IpJaqWndNBw5wVB78/+4iRbx
FYTx8gDU8z8oA0+YNUMX1UGZietpb8NcdEyTCfAPewYCKLbprgXDmTXDJThoFOArgeDDwA5hseRI
T+vENAiOoOamyiPP3H4jCQP1bBYkLGLVlu5d1pQv39A6Ri3uvR1oiZLyk+5dH700Hd3WqCjYZMsA
NMZYvzjuVUThH2RDx4V/LoulUoU3p8OkI5It/3U9Qsr/P5zTeBH1g3AhOKNtIlGDDWIZ3/c88J8a
3OKouevUG6PZG+QqUyVEppiW0XASdK20zsA0qA4+mo1Ga4XL5ZrJfZQ/6bLmuoB3bRO5HMghWtRC
DWcY/7fcRJorg0K9OUaJSh4xtceK8HtxQucoikSL1IuWxSilpOuOr4iQ5vY8tWCw7qheJ0EnlBHZ
bgqLz6BrtycYoxUwZ3hOkEmViKajDj3n4F+9Cmwb543lh7l6yN/7x+pnpqWgzBUMudzwl1q/XvHd
eHJNSzkzUl6TQDyG+lgtnpOQ8FZrdLjmkb54Kt/1uw5oTmgeTBxvouIpF+IBjU49TNUAevOfEp5k
oDeG3NH7lm6K+aohg/a1L2RM2vUuBVeYaRlPC7tkpDzs2TYPTRzSqwiKeGvdcPCxdPomXaLObWpD
vONKYuqN7y37eDR7sM/wxdFMaxOSRHdlpvuLq5diC2ko09Kn4UYmLboZdK/5g6MIi8QOn3TtmLke
EjM3UHNZA7+h1yeVVpTOgKF1YlQt1MfSP8X0reMR0KTXSfSyrbjwQzLiophPl9Yg7UwXCJ3CXmqA
DUmr5DJzEGnolZb3dgPoEHoiHi6lLp4MK/aZmMywJfV01Xi1sehi3qr4F+ZLjT5VfWu7OfbpFiRH
zGqvSWukzWvAe+HNHkPjmOrG2HEuP+oD0R4T44v7w+wxLExBfFgSYHdhOogtuoIZ/5Z3DTxU/ZNN
MC785UD8zZSp5nhD4vvPvZknwZfEFnMttjwIiAvIZwqxGyaO8X9P984JCr87XsWy5WqxyD/HZ0f9
D8VF2MxWGx5V7QQAeYjLMEbIQHX5s7MPjf7IB1dKM3N5bSGR1haPcKbvzz3ad8/CJ/y/qOWE7ZC6
4dykVzFfJxdNEKyiVvuNYKTLbIwZ3RrQh7DzmebA7A2WT+WEwStNqK1LiJkY5bg6YesL4FJncgx3
p3MF8mbTka0fMVSBCI8gyPlaM76z5yXnK0rBFInEbVQmAmpfQBRX9FP9oFqMb5rinx7tnoXa3/GI
OYN07djQy4oRE+GgGnEavA0K0HGA6kFQRfpNb9fDN5D6X1IqbWf8ERpYETiNdJcHVu2qVPzDCcdb
6PA7sP1gMm1tq6qOn4vjMwCAFBCeRbcIVXQCRwG/VZXqNtZXreMEJFCDeC0feAP2guO+/OiA6zTq
sDUvpZKDSjaplM4D2hbstzNgmd8JYlwIRwH7uPuLckh1+HEfnRD9PQ0OLrw4Xqj89O2S7Pbs6g0H
SrPz0e9kF7Kz2cUIZ+XDOB068O+FYg0nINnLVwFVkXdN+mEXTymltY9mR0pJ7eBHMQddx5YUZj6i
aNTaP0ryd6hxPf54bZjwiNK3cZOVRntMq+aWMWVRSROkfZ0C9TLJSbBFfiKVsXvOSvLazsjptGka
s0UaVrSruQFegrB66Ww95Ijx7KfmIIt9GkvjWcBOuegBILtUD6x5vFuP2lKnGR+wbmJpSYNA9GsR
uyEk3mdnZjGZceKuI5Wphj8auOcQ10tl2ArSnYhk7CxNCofufA+XULC0PArLmN/HYHp8O7AxQV2X
+u2vOcKi5jNpylUeRWUZImBQIJhHigighWTEy7q6SuLm4WgE0jhy6BQyjMr/Gbm5Dvh9dkPtNEOp
72kLZrUxrbl7xO6mQiPZiEY5wXMH2vFryD3/4Cd9Vy9y/bQYFicbQFgmB1XGHkljT+59r6Sl8/l5
eiUgVZNRR67q1j+EO9QHtLWI8wT8PBZctBUwIP/qxQWqCOe+jFm5EOkVSRwcq/llhc/+bXur7cWB
Nu7XgEycmsvHst48oV6rSGRyZZtkjyr+1kY0Zj5J4D1q/bnZW6Pr4YdVWEuY27QFTrCJh6QflS1o
VPH13pfbVnO1Ask7xQ/rWNB91UO61aQE1uTrC1e4TkHFnNczbwd3FhFSY8m2+dwmiVYYnK/g+fQU
ELUtC1rSJ13H/cDxTdPRR0Iv2sEGfc/Lj08Y7hAimpxq2B1kyyvHBgeoJZbXHjKyDJNNCPu96KTQ
NTg+ejA7Cf0UmhShduqCr5VDmIhT6jIHKa++7l0oND4LbmycMaYp2HpOnmKoDCWpsJH1bfVsr2fA
w/cKopukKRwKInNlbq3Lr2A32dnfuxG8CKcHDa9/IhOIh6Sma4tORzFUopjc7poQySOdzSC+4ex4
Hv4TvW40MQelDCVQjWuQwFoiCfD4ZcnsAS5L+Ez7vw/Znyualb0UjHG2KAnnPMgsVwyu+f8ou0ET
wgOPphuSuNSLIJPcvMQamwAiccpR+Oiwjq/nHOI/XOlHvMHSHhggwO9pN0TUsgcU3IbewgYT+ESn
XEpE2wEyYmv88476teEyqHXvYvfxTnXx7+fQiSSVC2P4BMB9NSkBXL2h5oxLuNAgFJg7DnpgITFR
9AXb2s/nCcxf8F/2CYNyYIwfd3kiKlI00K2RjWEldCO9MXVmCZpU5SA/3y9EY+irJhGFP+GxVep5
ZZMX1QyCuI21M/QnRmSpd4989Wjn+HyjcJ5l+YTVbSiPOD8G0uZcFwrLpNaKU6CAKx1+qXlKAaB6
Tgzj5sSf2y44IPiQbjYwLVvCtDOIoRAJREwrsyDr6LqVHffikgg6G2X0yZ7rCW5dzzxPjNoJFbMK
dKHs62u5jxrXy7m1kRBKH/CUOTCqbbiRuRvcqrHvivSWEb/Eem6daZeaN8cqHksaZG3wZuV4iDdv
ew4ppqtHYqPPB5RbYjJTOeFtq8z2BdqE7UO1gyNqmMoEktuPb3FBlLxZKhJ1gL4shBtkf7KQl/k+
HnEZDiPEc2Uz1NfBO2tqFJfLN5Cvx0LXtG7n7Dx7bgzBVg+FxXaj+xXas3tJQVJ1lEq/yTl0v2T3
MOdzBLU0vTQf2ZyjHP7OMTJR8Oimpl2E8yWcPRPDdwhQIHMl442Qgq+Gb67m7bQl4bXNwaRHO7it
anEkq+wScTIVGYUUDHi86pQciMMPrjO4Q/4Sc+xuQR6S1iENktFSmBFrovGgXzbAaYvxr+X4GNcg
QXsrJD7v2upVV01/PWjK6AIVmTFXcosR8/DGGgiq2eD5l44PF3gZJca1b9HAKnTU9QOPJBC9Qty6
A1eACa2/iWDr6qlfcaE1IO0lLW7+Mhx6q5Wks6QxQ2YgG9eQJNKzMf7Fayh02DvdLShimNdnzgUd
qlUWDZ+mDkaHBToeLoHwhPGXTAjhLBIaVo7FV1VkzOCBqrdPOqa2VSGrURZz/pAWjvB64UBI310O
8xjl9Vz+KmXziXavE1N+ifnkAT+DDsBHtyzVHzy7FAKLTGDyiZBM4G7eA2kmqTM2Xyw091xzc5Wo
MHsC/kRFTFW7P8+63ISwC8CYXA2lqtV1Fe95IKKVe+3kkjpEclicvV8k34kcrFljliK/ktq8G86G
8dG6Wrfsxl1O8vnuzeHqfbVydRc2aNV9lU75sSB73zS5xrveq3+hvJs7MSZ/ScciFiCItq6i3MTL
+sxfEWxaJOZLKQKRQfqiVR+/Fx0w1sEf5TqJJRyjZeC/hpxDDNoBwOLmx+6LAQtDwjczeRw2m7Dk
K9GHShysV3YV4xA1gVHLqdSNn8vhnKF5AKm3VTMYs3jQOJM7Nmkf4qyr4TXJPTv/hT7EhMIw76Rh
EJEITmE2Y/WnhlPL0SyfBiNwFb1ruI8Xn4fgSaQCwwl6E8N+oki9+e7Awg5AYBPutPUa/EfiIKoQ
OHv333MhpyAbax+Jo2ezK8skEUTWFw77HqPuFjYg8N25qVUCb4KP+9cuOFKDMtx4I32b2FsFUOEd
xleaz74eH+gtvgPn8EWymZKC696tucCu8X0zmR7iYRom6c3ZpVCV3anrNRfWrY+nd7IviA9MO1kC
XR7/U+WrVsCe8TlUrnsFMlvuZiNhnXDIBYFbRilT8ftHd0MRW8/w8iSFR7xeOuLL/AKonlV4PEsd
K2TXhj1DlyBNOLkjpt7qDd6FnUUssZmYx/Y96Wt9s7PQOkentfqQ6wgQiDjx5of1qyP95rFkqz1E
AuIzurAxtjI8Fk95wL3RYo7Y0RfznjWLD5xygx30x5B43sYn1yxCoiUJpn50HO5GtR5P8O/msLpQ
itIpY/MB++1RNjbTgkvLvoKZOthZRpSCmPzR5fxOE66ARwu3s637kX2HYhZ16lMSlIIvDySYElUG
O2D0mnGRACsrGjQ01EdcgYKIlrUwaAlEjHcOS/D3z3hw4hQB6RhVv+2NNx/o+rkc7b9+vgGg5YWa
tyCdZMEU8KchVH0CmajTGwYaL5gYTVmET6CZNJx8R7sh6TXenkHKCdW+lzEQrNkNqkXLPGm2/MaQ
QhuSm7RWLuL6BmQYd80KvDtimLQby6VcDzleJtv6OWOz357LW+SMNU2o+PJRP7juD7XHjLsOvreL
1rZpAgZi0F6lHg9VS9d3dJkd5TlmCa4DoP6UuQ4PmezxhzpdHVbgTRxKwGRotvN8mJ7sHOt0sA7U
`protect end_protected

