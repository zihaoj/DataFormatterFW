

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
h6CvGMJe9ltbgvSvdNvxr+xWElLeWWQogLzLu5SuldOpiRNjs0cZqmvdfyH3mn272uSJ+pqX0ncH
zgfSG+Xgbw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P/ZbEjSY4ib3C94+peyonjWBNh7YUkpPFze1WlXDyDK129FfSDjL6KVm3ZgQhqVSkEBubIIbqeU9
+Hs/qG6Sdyxo1pGfCc7QGLjOkCs0EwIOIRnRPrhbqAYoO2HkPf0q0q4YBU1AQNFgcY/IFPAo0RUk
FXJmSS9UWYiWjffzneY=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fbnuJsiiuYCvY1EZKJuO1r4G2rdEap+7MI72jtAYyXeUfg9+dCvXpvo050i8uj7T98AtzHE9ODva
x4Jdztaj9UVTDy6KWYiJ2VMGMoI8Bhyhb1wWgQftG2VCYIKqM6ac9+yO9Ax2oBcjxLrVToDoYr3d
rtkxCKh8U+dzxUCH29Hu8IYb8rzNZMCNAPXGL7cvUOot/NUpsklQR1NitFWS/DQkM9HdAlU4WZyA
l/EH63k27KfI27RvYKodYxFUKt+5eb42EGAA1pz1nx+ZWftnxKQHxCcIpatLCh4BohXh/Lf6m3lU
rt+FR1MnER+W+tZiU0qF2miaPqE9pSCbGWdMgw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mA9ctEkpntDb/h4byoy8xKqUG2kY51sDSIZENRkAkDW9ELlCoFEN52ijlYWikAoAmSeEkemViFUW
sJE0N6SWKlmE/846mpyavlVJIk5+1nM7aU1NtRauoDOAFSbO2YIBQAgHgwTajfMNISGMsCDTBeQw
u6xCwDcxE+h4t2oiXuo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Iu5xymwO3DvP5tF5nZqupqUHRLTA5JgP50bco68vv8zRTYF40vPWMmLORwGgDE2elxhN/mN//O8k
W+eMdPtoeegP42sc7Jntj0BUC+3J0BpLCzExs27LCl8xaFftnO5ouqUGBTjrckAtlShtp70vRv1S
lfIhfZdVOqYbvqJGRSy2CnargjSoAGerwsaPCQ+nG6+smjblKDdD30pB2G90mCzKuAjDhJQDULN2
qFeKZS7gD0L/tk3t/t6v246R8UYakPTFOyc0CvEO8CyDqPLA90YIz/4UrGsL3jRVh6Fvj7zaUjJA
rA5JgP85Nb1Uab/vKFP9/pa1ecO4q9MhoN9jGA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5024)
`protect data_block
8Om9Znm94n8pnk1ODuAfJ7zazH4IygH2dhHNMN9UkP6bgJBg84CYnbTCSJiCQPVWSGUJV3ZyiURQ
T9IliWPYfcbAe+odW5p/mDkFPQlTEqykkcQCUCDQy5mtRF+gJvRlcu0HQGgkpc9EjgZsT93z8I3D
8DLcSXP9Jry1FHneM9onIAPZQftC6QJV96tEUzNclV9iU5odvd4mRGnK6es5MoUVPvtWMMAV1GDl
bq1Yc+JH1cti7c9odcibSWYenDJJRirNU6/40+IdNvKaXh/jeAR2y4sUVagQZgkF5tVpGALOFRpl
qiDLz2j56/MySDbYNaTAtNn3abMcrLT+IG2ck5mPKP7PHj97oApHaYKCNj/lcYWI7C31cQDCx5qh
oEMER61r1zY+TwnrAP9/Zmr8C3Qvfpl5uK0mKcyTfn5Dbc1BvgaN1N83+9Qkg1gMf3fNuPYy8Sq2
PM078/Lgf+yMJ3l63xY9dXnO0SkcGzdk3sdwPl5e/jCWinjzijWZyOECEsqCu8uDpQGjOmi57TTH
9JUEP/0BVCUaoVMpZmuIO4Yo8quhAnchvoFAqlKUSg6ayqY9ICIPVjDUyE8tef3p8V5TKJG3FIrz
lHW2h6EXvUVGT0mHDY6r3ZVDYYI9zSsT7IeWhUpBUNh6axQeMLPEOEntZTXQdMrx71vXCIee7sjO
b1Mvid9ywoWHvMwQnxFwOiJTHi0yMY31Ds4MuLnliR9ba8DtptHaq72a6+7o7eDX6Yqc3BeDplX5
pX1pnZXSvGqYXpSalFKi4n8+z5alfCAOi0YB1Z/4eM0bEFvsWpysgn/qWzKV7+BqmtflZLwn6VhU
QggPP4RdXrBjw26wmUqeubprKs3nr4d6YBkJ1P6TkddPRdv4A9WqxISVP4AfLj6gAp433EgsQeof
l+6TnfmhSKrvJl9UfL2GGG9Urum2dpX6v1Hp8BoVKLxmsTt6I+N9Hl7FCOcm4ghhTFFNR2H91lVo
aHNWgT+aUa5hTo+5yL2JpV+s7r1BLPoU0dnD+vyuHTVnntvyvDD1cZ5NPl8+Ngo8V/nsQZE9vlgo
thrhXago/Fi2KG1ojzYa2V3PdjxbZWn+oKwaq+U6qi0fXwGTaMfGB5axp3KQByeog80fBgIxSkIp
26jOiysNtnMTmY8qCWljRx1ib2DP+MZv9M0OSor6giqxPMS6rWkfrGAcK32dwFe5/na8F8ieVVIF
ZPkVzqd8mOq3IhwccZ//7ULLJE/AgV3FLzB9LzrP8vrtPG62u5rFH93W495vPHf93FN5i458sh7h
telqgpHlyECGEKvALhvabKmAeyyZi+EuDrSh+9Olz5mCsiIlxv3CVGfXY+2AjdDnUcrz0ZNqfP74
G5c1gB8910I36/42XArTys7UErni5FFNwArvxCBP07dP3DkT8PiAXHlKtRArz/F5x5mw7gdIYuC2
ldK8SL3NzPw+SBaMNyv45g09D0ksdX8WrN18m9GbnFQFaXm51jouvd3gTWHS0eYwn6DEfGYRyTr7
2lKJvdvCZRWcicEQPvXPCrxAGauyBkuy6E4lGJTi9qCtiCOzS/7lq3pVqonwNU8nzMjBrvhm+CMr
FssePIgD25M5MaykOxEcvKZjitS7ieHyhoNMztyhr0DcfhcQVKZ2AddQOdFSixlKrWmksqNiD0Xn
3DZ7UfxyPESADv6w5epZN4HavqlmtAYUzZF7Lj2vJ1S1M72x1dpWOxC5b4beMGnnZCk9GjHf2KLz
12BVkMEX//OQEvPodZUzFU/lAP0AgTcy1qpcUFL0pjEFIuxoAl4pF9b1+Z3ZCVZmluKtBbCUpAxM
FXsKz3k3gK3vpNsmIPlS6atRuzlJpgBW6dXUocx3hlr9v5yhgNBs8i/kl6AThLy6wy5tBvOpfJ5O
hDMKiigygBa74T5gYpEpIgXhbw0FaqUmbuejSj3KM/T0O3m9q3fUupgjk3WwOrLzvkwFFpXuOGGr
X2VVqaii4qu6LT0inankMCz8viunDZeVuxS7Bf4/3vGWcJzYRkKwpueDRxYlqo9VvBUTQjbMM7In
38bTpFo4X3wgtpgIcA2XjHPEUX1CZI7PV9GfYfyHPpBj3ap6X/OM43eOyyh4k8thYF6c4ZBLq9aA
BAWv+MzXW1uBcgsmh96FSK6OYV4WLCKTILkLfNzAnls+l0VL5ZOecyKo5CDJ5SC9JnPI7D+inajj
f5AtDb64QYXxybnEnP9rmcnljTYFOKFN6JZ2M02L7c9AneasjwNbLoB9KHfFiEtfrCqerSwoBHHZ
Yr95NRM2SX3vjJ0Kb34IcFIRurkN6/2NCkeBdFnAQtj3LJxcfvXCqpCDMIghAZY+3UAlxOEP9zNp
XdP76VWyx4w9UsTEn6nVEmTgrbKD1+r1NUk1SxAHLJSIHn+yoHnsw+PyAFvx2tTVz2dfw5vlILUc
umdewHiCqUJSIsOz9yUyVRuf5uHX3TuauOuriVj4V6EjPT722d+b2JlabaV40Js2cC0NikTJ3uAm
M7SwEBepr+f9mvx3CRGpmH6tmMi5l4dxnZu9WwFkpBRxasgK2eVadW/xKJWLxYs4ffYMc53+CmDr
1EFuN8aJObDDqZuQOABT/4eFRy6fkEhzbSJQpxjBfrkrGWhTWN4oWtJ/vrwVGOdzgPx0aIJne9GP
MFLwkkS5vnDzoKkwULCDzgQihx/sIsjSkJ838Svu33aSNlf45RTsKQdq1n7ozlOWsGl4j+1fM/1a
O2/TmpwmeN3UzeCaACszeqGEanF4Sbphfx8FtAv9bNUuVLVLaeRjARpoLULDq4f1TQYRntMgD1e9
k9IG6jArJ1wjICs833ux75UHmVs/tVuEs6zMPs2sxdTRsrwJJOfBathQqgbW/sFHVSfgjqHAC8ww
YCyfSIxOM2xUwg1NfNB0MB/UyWK+iZuSqMwxtFAUMkweABbwowqKSInhXw2IDlJudi0LBE2xaSrO
5mYwfreOqsg0lNQ80xngK9ZVTvZbm8T2XJOt7npyYzO4sGtZVjGiYNMXDCSXjD26EPY/c2j5XdZN
1D24igJsWzauRFrIKeop2i6Yqws02q65J7PevGBbqgks/doc73KkVBQsZllyee6mzdEgzRALJYVR
dqYsG2Q4yAFfpsHNpKP0UWSWruDYqhZ49iv09FpabyY/BTu1Fbq69xDbzreKd37VtFYM42UpuOvk
rUOWP92EvSmNIymZ7zebkwjg0mo83AdCvcmenNr1geqWnX933ZEEBmGzl+uG1gcVrY/Gs8Uc2Ozj
YFQAfCmdUmd9mY+EoEy1dB5gTb0Rbbvmu2UNMtFp00+lWVe69Kndu0gimeoTgtTdivo5k5h2qjGh
6zxOFq4Y2+aXWaFEh1HPhuHYYhCeUxcD3NfOKHW//WSlNZQK0DTF0ikpu5uqCW1I+S+tjPar6vZu
lOc2wojm3ZpqjvdMCb/WMscox0Ez77aLokt5yY/WEtJ1KU24rMSJPYO9PQFZZx87ppGGzCHG0oZ1
iCz0JDNe8D70hxTkTRHR9Pcndqrz2WT07Mc4rTHI9Mgub1IPgfN0+4ABH4iEIS85OHqYlj9qZT2D
G3N0NekW7c+R7O7QklbEPe0yCNuAQpZo2OtNOvk+arZf0Im1FQsQ+9nNGSYJmYVhqQ8dxX80M57D
sumq0xWXWUvLaEZXOUu60hbqrBjtGxxu0O0t+ZP8WdiCC+konEbswWPb1pvvqlwyB9lKIDg+4itn
1kG/FJ9VdVe4EntmV9aO14LYKo8mmjYaHgK7SbUBodzOpIv5uyOhn3rUQfrsIyFWQWlKCFdEy07Z
6Sc44DI/h0NfeelgZ1tk9XT4UMh0vtbJP4LfTwnQv7+PX2DpRPc5jp/Dj8kOOTpAobNkJr3AZZVZ
1jkJtpkM/WrxFA1TJtiIN5KBluRDlQR4PuQ90l57l8yFPFbW+RN3vSuWb4jpG6z0eUtkeGkHlyOR
ThFbltHfgQiyqeD4hZL4HdH0dWx7Uaumbz3K9BDKbzapIZML/l/zNZIU5qrxlSnZfZLAvcthm5eW
J88ejvJSLsSCNy/QKPXbytLm7yjOUhwDOqdkRf5p+n8kpr546BXgQYZocz4CWb6LKo/sBMZjpfLg
dtALj10tm3tKQ8iy79R3odECDbztz2nctD6oNilz/5Ivpzwx8NGqnREdHAZekPZqXrxLGJtfnJCe
NyESZ8vzNIj4RL6T4Dc61LJbE9obWCvxbHn7CkRgA7d+UATxAroTYRiBmFImEqnwf5Pl/uPeXF2N
fmbxtCGlAhFeVawixmdcTir6qmwLObMpwBcFAGaK442k1uI5sOsPg1Ewubw+LiNOs1q+sf6bYTZR
RgKffl5s6J5dlpy7OXEZ68mCio3OKMopM98KiyIYIDs/zmNpNGmzGKlNnQoRgk36J36zSkeijee/
yfMY/80P7NvXNSjoAyiGV/+MIbV1RNMiDk4dMIMxjIOi5pNXE/E70DUJxC2y+jkm4R6OJaKchk8z
97QoTLb/+yN40C2hUP0R4SfMRDUUoAYjP6rBrhgUWsjSTQ6BWEJkZD3/2xD9OBFVkauTsnWyA7bc
lD7afBgFuxoNniqYFNiHCZsGf632b4OCJiHjeWqeALAmLMoC50RGzstbNgx29mPG04Lbm/u7iBSv
VFjwOAqlUQMd7iuspXx0lxOx4tlWjmvYm1d8q1JuQnyXsNjuYMYuIvt2PX/Rs9HPAB8SDlZQjnxc
KDZqy5FJ7nwVyKMq4r7rIvhT2HDvfU2K0fzF3EaFJOH1I9dratWU2ygPCkeVN/iQJay13wbCHH36
I0gANnI32+GUWF738/P62WI/og6P+QGAVadAlhyohpXu61dULVO8ZHBLSAbGL995Pc8Tn+tLcabh
BNLi69gtLd/eCZdUI8vXmHeNtvXxKx3uVMTBqz7SBj1prq8PpWMRWDei04yPEY7iz27W8g80Czcn
xAJPcu2cxU56XSL4Ti654Y8nVXd5AashjN23XAy/2g3ylU7rCgL9WYwUu51/BqEd5oUlWiehLOJY
MePJksW4C1QbGUbgtSMxqGVhUa69Wq3bYTgoaB9h0tntZ2pjmD+qyEZpNr0DzApOQVgQ8Zt49cyK
VBftX0T4QTU0CTRJgmsXQgKqHcc//TC6nTbTRpmzNq0IxrNL6UtOzbbUvotcUKWOLjuU7NZ8FMEB
3kD3SLd1FvqEbmQKLmfh9l8lJRivDsBBm/EEB78Vqrza82w55o2spFlkQKAZoyQrWJsI4h6BCqkH
9TIvU7L0BPA3x5/uT885vWIrxZnkFmN76I9PzRbJ9rgs1tjz/seLJPshBqQy2L4zECHtyETvJLgJ
3wuWSA3t7bb9md4tCl70NR1GKQ2Cj7b5Ws/YDqJAM3t9BOVo/0mnh3s0V7igqYKnFJ89wl2Ff7CK
bDWzVR6FihcrfX0Gx/K5zrmKo0qgtw8yhaz/kce0NFD2snEp6TvNtM8d+A/7iAMjZ3hVEaG9BGaC
6p57B248RLxmuxN49JgJKOyKzJxQ4UPJqNgNmJmZpmASEuhnWCPotgsiOfqQGm1Vu8hJQQhIPNE4
QFFD3iw9MpuX+4rC3JbIp31mU2U04YhEMBsZcgIeJbikoSK9FJaO4sL68z6OyUdzKlwUQAf9Mchn
iw/hWmKmWH7OYhdA/KYnIIHaIL0KcOj5b24RyGLomyKsikCKVBWJApfigEGBxz8iRU9OVvIixne8
ASIwPUmfUsaWJx7dl3Q9YnV+FHjHzd0RXa5lHp2IIYlqxsvryDvIUV3WLzWW9JQBBhDVrrwT6pwY
k6AXAG4U4CbxgfVx15Nov2vigPRYKq8Mjs9flPQRejuughtBmvvjnsuCaElIgSd5/jn/GQugIkey
OZ2Ljh2r96U3qfR4UzPo8vViFcx4PuCPRAjS7S8hM44rqrT6bqisQtYAHWXAW7GylKog8Li+xm0j
UOrQCjg9dI1oqaNUgwOwBkrBL/LqPTLZ4vQQwnpp5CevhR1W0+rvllzAMbL5EtsozaiJPKeoE2J/
K2cirqApqfogq1w3x7KP4kfxoSb+b4Glppc2n40FCmNxxBb8S2p/Lyzq7JaBlYOUVdEZ57YvS5bS
Y07nfPE5VzC6oLFXLbTLyQqiBaZ522+JkTxabaEUyu2fLaZ/Ylp85prnWqj1WV8xeTdWCWC1lzHd
yUZBh19bWmsAnJoi24uaYFgWTFVBgrKrQixjFswmiWiJ9PhOjNDLvifwPblHPpQscfKFCAr6UiwU
TU0S4l4CANFygskWMgeMvT+GHFE23z5zZQUVIkIw393Zmda0wCGPjChTFXzxPsAC/1fsNJFaTxIS
Vu8x40qJoeNkKpF+pBTCvweej4LK78Usjj94iJaUn/vmtIamII0JpxBM/qhyf0wt8sGtFOShhIvP
nV++EmothTYmVnfjf5FbAEx3Zzl2garV1nLsss2MWeaE3Rz5Z4NxnZZ+tn0Wad1OgEQ7BU2Nc1Ds
v+4IpZrx4q908fIh94E4snAa/xD2nCIgkwIXplkevHitFvN+JbYFYz3gH2YdvbzmJpnVExKZ+mii
z6JDZhAKiMRsY3s4UuvO+DoLIDeWoqliX51MZ6kiDlHZ70ob8vnp6RSBLUazgKmJJUaRuaJpn57J
UQTYkPyWns/1Pvneft7PrgDrDEauI8/lQyBnbbuzTNQaIgzsitU10ATGJ411KteeBYAdhr4j2MKU
QN6BZyT9GXE=
`protect end_protected

