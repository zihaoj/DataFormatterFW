

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mqShA3L0xrr1CXM+0YZvvtaaRUJ1WqHYA1RkCJOxptKHHEZLZ2TgJlJnf3C7aYSPmzwHBPgrEZ4t
59sA5Y98ig==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MsiAoOXS03LU5j+lvMIHiTAH/76YLmtmAHMzaEvrbpLRgWJdLPDvkZ2G4KrBYwycx6q0zyT9xham
NLNIS222OnRpye8y97Z4zPgF/k+fzoe9+Vs8CWpRHz8nk6+f6b0uArY2VEg5b7PPDlTlt6PsmkCi
T6ruBr09P7+uMq+TDm4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cdLiP/b6Cg3Rbajvmj8COjloYcjaYIzGNU4tOjn5Nj2i+hqW0uuYV/wb62Ban3cr1mK+DUGNcziO
81eRRbw0ZDX5lmoiIv25wRLqUlqPVQPhdS189inchZozOdz85xbDNO5FRT2jRyGIAgQI9vBlr6Iy
61XxNTzzT8zAGz7vaSrYNcmgmFfTuNhDKxvvi7Ayc6I1vRu7P4gbScFBa0WMMOrcLvYpnO/9nfiR
plrYmMPadMOYBckYY9NhM9TfVEfCFxm+qLVjb50vORqJwd6EIeub2L4WUJpFO4KRrkst0TJ5mqZL
Cpnlckg6l0srLlRyRThWFvuWbiMgAcHezzck6A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e9jlbS1OWz0ZIS4Verkx7Cp/oqMwNUuBPenxtOPRz7MMFBJZ7J0clStLHI1GtMjq25gVt6Y1lDPH
spzV//m1IH5JReHCGtvCxl9uUegxewzheDdOOL6yJEPGaCFIk9lHGqWBnF5uteUuswXTaUSnX9cD
1CtwOmmGvUOA7Dy5B1I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YkT+wIHcljuI62r4ou0SHGK4tNN4pTAPncGz+/uG9RXJkJJkOwAy0QMgF998sE3bQskkqRitfALy
TGocAiE62Y/7v/NTKuWndGS8MGKgIi30t8b4B/pbdK0pyac2VMdGsZI40Jk5PPbMZMerhyLP8RnP
wNdCEZiEPw7IWzoYzJwMoE2oczEkviBY1Qx4AHm++6e/BXfpQdYo73RMqp9ybDmrX9k/xrDfe9hW
ydn8D+u1UetmVzbFjtSnGhOOyByAXmsM2T2WvDoiIodFPLVgpIVT3/MlHhFWWLxbJcdBitX7zcmm
jF/FfyufENdqG+S6cqog3/Ey8LLxEYRqY8vBvQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15200)
`protect data_block
9KhdriTyr5AOskrxWVZLjy+9Duc81mrjEE2tCpDlq6RS8DcWAxt2O3TDn8oN2vVyIG+Jbsn3TKPx
2KqiboM2yrIAbZUG7vVq1lWgGZPyYzyMkDpQaMXjEojRJ1bgKda+G4QoM24u44zC2b+S2sTADJS9
R5bdFRIdAEeimzXRKYWx6DlYauXaQozm1jyqKYJwVjaa+MgagbJ7uiVLuZlWXSXxrkpwxZzwe2U7
FBpxG44NEpDRzUYGUoeIiHgF5hbwc+LokwDxBa7DvoZOlEaniVUA1bcN2EIwzZjCaHvvhScIrh9l
/yhbGO+7R/KPURAoZHdp/BKPvLA2zcG+SHscp83g7uA565XNm+2Apt7G1Gh+wGrEXEzbTQSN3zGz
jwBYCQqwzIJfOSz2LVxLnqpV2Xunev9RukvarYui9ShnpebUb8Bx7t4tb3iKcZTu+bwh8JKZAuRf
lKWuGMthgROnKLgKB+BXSNzgvxeMrfRBZyciKutLvHMAmDNg3Zbpq/xGU66o0t5CqTfWJRLssXDp
B9JhCc+HGtpG59Lw6WH6liBjE/MmlV2dMDBFPv+LROZ1dmgEjWsR0ddwDEVjt9GLYelPC1fYFJ1L
1Igqkvd3puRG/+qFZH/c5NsmzFOInEUgDjXb0cczhIdbCXIO80gFq1QKIsVdgRaacA155zOsj/iX
hjAL2Wjgrbg1Hn9Mwu0MJ01luRxywLkSw/YtFiGxbm+UC9qleYqrn7ZsRFDpghUgHitMjGnNxzQd
xceZwzRnKwvIrnvn/emDa+yctKkOhU/Id6JJTRPhu+TkjlYxmbt0HPqyGu2o8DYiFIx1Fhc7jdB1
w2yEbp9nd/lywWfAtUR1TjF4gCvIzUeF+Ac+orXwpuQz4PgIF0a2q0tMc6mkl8+JnVvwSb8v6eRx
6oMpM5c9UckssDZhLQ22k/0bQrST0RAlN37Ht6vB6d/6PhxKAx4DgHfak2diTM+HxAQJYuZldHoo
Sr02v6aNoESczHQXKBDm9YnsIunqYePneDoGeZTIvddgtFD9A4KLZ03JUuMNla53BgFSPFM++9BN
xMmnUMmQiw1VoSE7pvEoqkafNKM42Y52wwJ5ml1SRwP2PIIMB7al6GUeXCqwylsHV3CDR+YDJntm
sFk80Zuthl7e/pE9ABvaxRltu8D56XWTx6vJg79j5z6h7Ry7Nh0HeERKpg6E3lE0Pl+h6lIDvdmF
rh6rpnHQnHfNJn04522WefLF3OWrud8CW7ZQuuGQevO8xLSSoj96Ao5o9jE5riJ2aBdPEMovY9Vr
h6CF9ciDY/fvF9D4HmQM3hpFvPPCpn/kst9UFvRmj2k8CUng2Q1Y2qilnzQmNS4riXMWaJYUK/cp
OU5NAJDXf0f+59HLj+EAFL9YuLe7B2neg5Xp0e2la7fmxkx8rNpjiJmDU9KyyF9hXTQBTklTW+Ua
c4huyn/VELbqowpLMgFObKH4dn276SdiHj1u79xEx79pp/Mogh014vmQQUOQ4LSqEOnybKjYcp5Q
92gVi9j4esunseAl4FWex04U9u5P5fabcaW1u134/jI+/CknUcFQukHeq9HSv7Mn5WluLCifWMd8
tbbwTC+iUHAXsg/s7/mm1rY3iZxxa2fUUrNt45szOA5fkoWghAtPUf0J2+tyMVf4t5ujOx2HRF4j
Yc5G3whb2gFrsNXO1BAFbgn+4EtNc4p9VOXKl6474gtcBqaYDkvtr3JQIbc+O8O6lYod/tuui4ww
HWxBkSAsoHhNYowtVCOMGYgiF5VYf4ow5lL6BYJcG5yg36wy9bpNi/Ryb7I9PhPqm1Q6qh0fCtK8
Nog9iW3XTl9nqJyC/Wk5XrhP9BC04DjOHJk6avIwnwIPzlREH5bbtKgNMXKiv9Pp6WbEOT7yJvey
57Vj3DmasMEAEk9BVgHpYXnfLu65JEq9dYvv6DgqSCvt4oypDt/s6SyBwvhsIHcoZxDsBorZ2lZt
2LnIi4FjG+wLqjpinHGGccTwW3+OqlgQ2BA6PC8N9zb2EEt3pWOW85uLZzZF5qYd1tAPMD8+jesN
nX0AOEoRsAcH1VLS2qOO6XMaKeYeSENbYgcodd4HLsj10l2H8GCMsaQcwv/r5JNhHnY+ODOz0UZS
VwrvJ4GcqXJCHVzC881lHHSKJBnETBrCe+vaz6m202suVbtH45Y9L2k+aW2wJU0ZI9BykBE21Xqq
I5pFtqNJZli+Y0zKHEaUmxw+o/42/Uy08tCslKtuh8T3H0d8vJ4GAQQXVmK9nlLBrdJEVnb5MxyW
lHN1nGs9JqpH/GA8qQUfghJW+i9s/g/xV9mHI9FKbKIaZuO/TdxdJhbh62AYrD/iI24aBQKMIAPp
4ksKcDX90s3zBTegaRGSv7cQqVs8NISfslTqZEIjBUjbWswc1lW9P/ZpXshW5hZBkl3Zo+I3T1n5
2cqLM5q4gxH6jrH99G59+19WsGUfmwI/pgyW3WQU8awV9SMqse3VlHXrwdz+R/oSp/+C1r1RbFsz
7CwSwDwuOSW4oHCxA2k802o4Vi9ztKRpSVNq/BhozCZr60eYq1wk01sBiKQQqcNm3S2YlCI1URBz
Y8Yo0vdlYnSxoMtIz2bnfJjyGgHvTUUQ0yXKtsLx01yJ9jY7tnGcUB8HNbK++oehogVgHAhFGMHJ
hx4lz3p11br6ZiZ9ETdmWavADEcXRcSqdWbe/a05Sy8oy9LGHrqLyA0OGRqKayOTy1MUI1cFnGLx
4Wnq47UVKvgHAZA5bQxg1aDDm6OyPuLPevSADM3VDGBpDmS/oWunTupEXK5OzXGjyNcvv9b0gm2k
cWhQLs2b5Bcq+59PugpnHAuxATn/7EJnSmiq/vLDZElVa++vOMiT/62kcGKL5+ONXv6rqB4y8SpN
URc3yb3Z5SxcaHfHyaPI6hldESWW1f2R6C1rRJ3ELuFlTja3BS8xCIFBK+m/1sl/BOKJE1WJEbb2
rLpuFcE6u9sT3Wngw2DCkaEJVSnfisSjrZZUo2SkJcq1stdGFfzr6Gk3u+8ZoKn32+OwIXEbxuJc
zpqGnSQGCirg12XAriXwcYaUDWbGOGNu7WWROJBrfpEDWX1xKm233iA8A6CHFewZET2OGPyn6gIf
62C0qByVjNSfxG0OnZZe7WdzHRyxcTJ0eWPqPDPb91Y+yJST8bXFvEKkz0/LeYd+E4JurraXe07v
jlC1b08m30peaevNt08xtkBkTvnXYwF0Pe3zdU2c1MjCVV1J+gOt+xDpF/5wfky/mtlnsS6kayd/
gn4KjUI/o1zbUPGsbnn1N9u9QlUvqCasIARkaTRQfwNFwUm6pRmgs7wQSA6l58TK1tSedwsP+CsZ
yPTC9EsoAMFpI4SLZyiTlTdRBfyOTwj/avXtcmuyLL1A+1SeUAyiB+Advr9ZJE66xSfMDAmxCVcM
hs3zLsjlUQqSJZXWOUnIXxlg6culTVjLPxBxrDqQKXXZ7Q8E8XmTHYIvDsQb9qGX13alBu7PK4UI
4iBToKGwg3+81vCs1qM3Yvl1b5oAT+vihJmzPIjkwotWUrqLR+x0dIx9AH13Xg4zaOIEU2xYi5eA
0c8tRfxf6SZFOvennkLnfz/OSPsQyYTzzn/fcY/HWbf6YH4yf6yaOud8POJWnS7wPQEa2i63vdOS
oAD6dwoDnuwfzLqEvn2kbLs4JitEGKxwrL3F7k3/kfP4/PsyJ3OhopgkbZDUnNEJqmRVua8FGtLn
NZUueGrcNtoaLcH8kwSy8O+rwCF6VZSuTF8j38ZVHEFSx+yFA+5uJGYVWPtwJ3hCm0occ6HUDT15
G+tnXZot4rfvWifvLz53xOn0kRkHUWqNxQ3AXkYZiqwN35wYctd2FTNeKuuyxmjncCPPmeV5LH/W
5mhCsGIHAp5Gg/3RVT9K94Tvj9f0uWtyYw96Tgd5lyZDONCp9B3Rlg95QGfhcCE5qiafsCob0ug/
GgVK/gln45MBF3YkdyiNzr6m69gtSqbO5mwHsF1mQke5NVdtt3kbBPjS84Ba3Wu2DFNrTm5yeIDM
llgG4oyzBorw5NEDbUBSCRtO4KAdIIZ+DsDJTCOSiQrt2NsPk2iJdSu6p2V1UHfiRUxaqn/WKCMA
uHrOxZM6VM3439OMqZ9HdabWoUXBzYOL1N9GOcJM8GzfrTDiHc7dGM2zMzaCyjPB8q02ksA95NMp
mtI1T+nn+xcXiWW+yh8Vsd+FFrnwVT/G9d6iuthE6suNm3wGX9SSpP2yAhadUzcv+r3Sh5mOHofn
7rdV3Aq6xg/lRYR+K8xo/39GeRq661OSuVIc8Tqx6iYYXQepgQXg2prjP9J4Jey30ShxfAaEe3hX
iIkizikiJ/aEMo3blrAl7z6zkwLlhctvFgNBiEI+tC6QTrkpweEyjC/m4cOAd3iP/AsaAtb9DJRg
/YqqSqHUiAWLYxRS+PKfedaItRzJpG4EB4nu8xrr1pDjEwZoZ/y3kfkAmMjKXsFEf2sYaywkieQF
RQECCFGRQOAME9LeBPuydjIXzNm9ljSXF43WVV4tH5aGmDaBJurp/p+Wvr9KY+kvUWyPSoJVeO1F
cp/2tXAGvIlfSkd9xCB2uasYPjxZrVeNvQX7JyxxZsyX7bnkxGpVTMz0twGemMqUmo9e6PL+Hm0O
5gTD6BUaMo/QfmaN/HOMNbPAhOVVE4kFxwQfwj0fVHU0opUBd2n6BuiKiIZFr5G/N+FBvg1J8duB
bYp60mbX97NsgE7cZqoqMDHynoffKJmpdTkwuovI1ZEqtWhneczFnjJ1JHbzy7EZSk1C2wT/HsPh
ymTz35mZc0Y5pk3yEKF723MSPny/cNx+NPvkMeETYq0dendEBsaO9l6DR76GdFXItdjnX6nJTijX
8l81BcSuKGug9P0YjRQ6TLO2ao/D3sUGh64lKq+Qo8mwcaNm1T9bYWeeRVqLXdXfj6NdkXqktOEk
bcN/x1AS3pSSwXuqa1/P1dbfZJv9FYZR6y532ph/6Sjirccr6aF/gKyeDNtFTTZ4InKSpWi3TmM7
2qrfOjPK46LF1yH50DNxJWC7yYjT7oqRtPMG4hxozc6DkuGeIaeBc1h9xA3ZyskH2kz+vZYWfp49
baOHv5JIt+xC7Rqh+s8UvqbLxqDoa2mApE0elAF9lZm0c+u9FDO3S4aQYjWRNsPGq8zH1F7uziGy
BSLMMBmCiJrdFl9XtrWJTK0nvgI9yLAkkuum9iibdKcC5vsdsXWwTC33lIXS2V6xEhCsnRhPyHbM
+if1iHf11ZYWKl87t7qbEWimM/ctkryivMd+KesuBhhTby23iiNg6l6618JRd53ncJs067v2Rypf
33mxwOufuo2FjkwBs7UgotuK5Q2WO6dahNqCKkJQhA/g3qA2kabHX+Q5U1zixItAxsZpDGYi/qDQ
EReD95HeuSllwxZz4OZga9dd8P6Xj9zWzG9UPvjw+WWBH+inUn1MwntoybJbgPrODq9hnoC+9yhj
q9QfXSpGJaf8IXlYDrzZIkznfqH1qZJQkMW5uQOcI1GmC8ljYq0erEv5YEdwuKT2x+ok1JP3B7Yq
s4tR56Un4SVRN1CAiKgKuu33hdi5SBeiJjwedHaFHiTo2bUheykxscFn+oet9Qs5lC4eU/4br/NF
ZnIeX6/Lz2cmOkuZdPOj+bH2P3AwKSjoOVBH1kAeAFQ3EoZ+yyrDn8MS7/kclBuXXJWnxka5xeBR
O2GlbxjhuqUYqsJKew0xGZc/sGnr827rQKRIKdCjQagA47AD7wdmHaMKCkxi4uj+51Sd3ovmAJQi
/MDtWYxE6jM99gw8eFO3R141bQUQgfnxoCLk/QiXNpVi/hY3x+Dp5t9ZudoE+0w+m60Ps2eTjV3M
si0E3/abMpn+lx0LqRu6pzbeyTO+4QGfQOR2P01ndzEeJ3BTAp2EphIGjufBz4TF+odyMA3xMJyh
MAv750fzuGfZHKWlW/R98pWbKg/yeY//rIJbLvu1Ndu7OifzGR810NYAy0dpGmU4hW+Jye+CE8No
/UcwPxn44eVPmYiXjYmDxgSgir3LVP24jdn3w6UQoyBLD4YJ6nU4pPZQivl4gp0DdmndutK+Ifl3
WfoaGz6t5/t/gsH4diQbHhK14US8zrjUPICNvjbfWfRMzPkkhoWpJF06+4GDJNL0tD0tPvhyk0Ve
kOOr3s+CIe0mmLwcrZXHpFixabclp5ySM7VJX2vV9vZsWWobu40qr1/qDo2LVoVzDdEZYgMzYczQ
5155CicDaNajzrYmHp/CH3Hue093WEUEUt1wLUjcGk3bFcoBJd+DTbcYvsLnqOREgf9P4MIOBVT4
0VgOubYtnYvB1lcdRAzCVzQ1PEx1xpmTDq7VRDcb4hrbNs4WBtGQHK8T11z0TstlttsDu2nG6u0D
AYZu0MGZ+ew33skPTvMXuvubD/JB9ck7v3qG3+jQDgxqA4HF9Le/I8kAwTRllqQhNLSVOzGk38Lg
VhRw9r6YE7uOQnkWkleLPqr6eobgnU9IrVJy6jm7UaxZ9qxoxP1m6ZZKRyVtEcXTvf8XXQd/0k5q
j6+tZ7+pmJs+YKkmpFmL5MBurLWiUrjnwgAT6bvZX6yrhm7rO4E5+x1RsNb6MjWH2zsAIZ66uNUp
0IjflzS7/S6q3/VDRBGZ8kvuZRzj6U2G2HgH9mf/V1wo+sB3Ov4+mZnsV3oJyR5iOdVwgZp7B60y
MUpLfz3etF2zku4ToUN9jYshR9FS5QwR41FYo789QKXv1WohkB/DH01RuWo8tFAsUjEIap90fN7x
GMLqeI8VrZ7fAc5IiEVU6IXcTsRoCeSLxBlywHM0OIsmf56gQ6CDmHg2ARmuEn6Nto7pUlhT1nig
DNoZ6r7AZOrBD9j8YeCOVUW6R9nEsOcftNF6NnGdEHyGUS1h4J9KQLlX3PJRE+kCiTTsgDkIWGiJ
Oed2c6oAMQ7BivnbAxzYUyysDGi0CfvBN+/wW2emIWvA4q8MjukEyFqa2BJ3KJ3QitWFWHpxD62L
85T5jHcstk7zRZcsZGycKrxE7vSBO01cpe1F1VBYFUyIuRJXIwtWIeEh5lTl8vhikETxSsRLdCt5
c+9tPQuT0nAutnNrN7PW0Wxes+86jNRPQZUTukUxzJbgPtK6jsw2kJkxts8t8mj/1bsGxWtR9znW
g2QdQJKGUtOK/EPum95xT7wleKtUom5ex4i4a32WN6qt2G12hmfCmpY1JcgjlDXkvNCH4D1ms7Nt
wZ9OZ50uN46LH0dPch70oSByMYf48Q9t3lfBX4MLtS1o8hcZWJEePKH9cp1/ovfoVzW5nmM/9iY+
xQo8yPO+LBioai78ZZxJNUDusg6NBKLSSbYICPevZ0viLiAegtB7+wZppy5XcfNkC6BXR9Fb9lMJ
dOH67MC198xQuCUkwucjZSMGVI/weOeVReectjvt5rCLOSAjWhoIGCS010c5iVt6NDBTJsapgmT0
1dyjnCj5//r3fm+Kob9uu7zskHeEr8ti8InbWqR4FO0CDAlmpUQG5odug/3mYndewBsqOGlZYrgP
U8a2GMOAonx2S6gb7ERwEV6swHS/+srPoSFqfryEbzh8Ae//IdXZCJSahGEzUXEvmxAY/Y33+85P
KnahcVCE4j3QjU4USpvux9Umvs6W9pMHz3d7duN2yVOJVgF7254e/S/J7utVB+aLv4xs/jvhK8vI
7sCOkhHKKA9rrVxsNvOpB505rhNH3J1b3fThfdZvwySBWokj2TFy2hHGs/bkM8n+ShloWOz5lAXU
C7Cn2+92Gpi0cLXmbvmGww/gEi+2kYEapQiZr0q0sRUZ+cJPrJacbMLlrqgTY8HDJZT1+RBhmiDw
drYVDEHMzlI4NyNPkQygfX9MU7UDti9vt7frQDNxcnAUVZXHJLN0LANDSbQGksPqyOX+P5hBUDf1
oN8w/G/9bsdnVSzb6+GCk4krT3wqLRomx06iFN0oNjcAgLO2ZteXLuviMOdtO8K8vKvQLW7LrIe8
zkSMHtu93ww8tPn1v3qlvRwyi/qrKP53geahHAHWbnRc21TDUSv30OJTSCS3lfUURILRwee/La3Z
XFBX1SH04OfM2EikTea4BON3iRy+QEO1AZFMz2L1m33R5CiRWb8vR5ha/Q6cMIwwyb8dkIHCZr+S
r3Rx3vc/9eLabhLCf3OS03N2SHDrhPbcu7am3IxrtSE9cc2fvlJQtSyPnAGF2UPSL8j3sDeiqWtr
YKiD+CzrkmNJBEHSWkMg4i0Go9XWnfgMYqad54Ijv1QKojE0vXSKdDu5+FLHFvmF5fU5lcoLnXN9
HP96UFe9yaGdEYwyawNk2Qmdl7UxECJqmybsxvI3PzYWTUp4fc8s+2E6JWj4Y9Aq8huqBTFZXSBw
ZP5V9S2PfUctHsj420jVdgVUTHxuBSLEs5+hWLcwMJmAQAWHgZcDYrLQU33gj/yoOf7ekZuFtwXD
+5RsQHsInpLYAKbDkHQxwastnPQlM310N0gheTZFpXVtboW767zuWcO+U2M87l6YJVpSEXYMTOnh
o2yL+jRW6K5gv3BqQF2807USe8n4hjJHdm22CoUuNEEy1tCb1WGjSY9Ho2E485kAZ8E4Z03jueMT
A7IgtS2wPNpJa2UC/vjg93eoQZFbYnMtObkl1+c4/uX8UkostjF5ub0Asw7b0aY+ubk4GAf0fMua
hNp6bP/4rpx6xAIdqFQLanLQDcX97Udjev992eWmbDdDoJi3KkM5shfWbwggp1GT4KQEPE63UfVx
XkjMnPptm2u7Wi7jvPjYJPB8O/M+X4TEyCTuBwP3DpAjOS4LuAVzI8KGtdNAzEgdsNrcHeGW1l/2
/CiCuQBFPfRF97KecHaFnY+KA2RPPc51ryji5YIUtQN8kreWic1VTpT+0shIf76CfdYmmKNKixF4
x9MU+zpHHZcBjsnFes+DJgflMgnvUNMVekU35eOJQtWx/e9W8ot3C6gld6vkIA4qc/oAlhiFns3J
0Bk2Gm4tG0ET03Ot6E80b/G9Y7NSG0/jEc5MqWKiWzzLDwxFdHuL8LQy29RkcxpzJd3r1A7PxAay
ZwWL0kFPFBOFUiZWJCCI4Vd7jBSeQQlhlQZXtdpofWmpq47uVGpTRdb4OKQ6eqF2+jK9QLef9TLL
Y2dSTYsZcLNTBtczTr8BvZ2gH7wDo4sKcHkTwTjsQ2s8ezM58Byfg5Hms0LoD9ohw495YvEYTICa
byIwQH8R1mX0S5J+1u0NTymDiBWzE5oxGY0Hm1xA5v+UAe9b1vr2mzdq1QonL9XDAA1aspfsjel6
GQKpCseuLxivg4+EytugcDS2emA4w7UoVepmp+QMVT+dPLJdaQCgpyBHAHK66S8X9FHvJG+Ho6nT
QN0HMtkZ1Q6TwMY9dqpYKEMhKDEnmkNjrIcfDi/iQuQUeRd7WFVNzRJf1TTIzLv8J8Gx9mgxBCz1
vbQGOEvc7DImcHVqShtFk4cTI3F9bXQgtzdClns8v+z0iBJaQgihcB3aNxl3SW6RVlXxUJm7JyyJ
AoK5Jap7cw9zrYXjiQVG7YKiwtg/WYitiOgNJv+j+EStbUz8gqrMQ1Ro0T0D8qwVsd/fF+xmBMzK
46SP9h3ZIc6Lcvd2tblghpjtryEfilDGO6rSIejGo9UP60b91oJRIq9s5RTGy/5JovgJw1YBYk4v
5Cm/b3vjY+UnnX/kujCR4Tk2ho8JC/9KOMpUnSiyyortQLuAfUgn1KDhZXRGUNYOOY6OV2/XHLBA
KA6+E9E8W0S9XyiP49jNEDleml3YUyZmOWx4kGW4xsEqv15JbeBEjmgkdoE9DvFYvFIl1D9E0jQK
ddwDxu7Ly6WSIYlDlaScUON6JHUNTc1pZHD7AEtknumDTKTm3KdJrd20UL8xapEqGnNZr4ID+lol
+xFG7czNwNmcsGoNNbJIyT8F00mElKtAEun9s4+E9WDU6eGw3o64RgsMy/Hs8OZgmXDAhsVQdnT+
RdsBwIIayKmjuYWg0QomPenJUeb6pIhp6C/UH4qPbx5jgGAe7+CW9Fd1yzhXhus5Y1S9huunoJ4y
drBZUYugLx2ATFmg2WpLnI4E4tVQj+FK1KU3Q+9JyfPGktwdRZeX4Y+c+5vxq2lbPLZPHU4tQewo
eczMFhGKGDxfjnTivkBRxW3ClS8MCfFsnqaCkBzzXi4oHXN+qXJrBBa9VgjSAjOhvk7y4flL+0au
E0kodLisKoSHtko6VqsVMsuktYvnKqEUquPOyFdf8b44CWKnJdbZR7WJNXxf9g8e96mHWmCfP3KV
lcUr3EyAI4tgYSgqC9b23zKqHRgrcIyocDMwKMOwRCH1KugXuoFfrNc08eiBtUCujw9n05g9DnUq
zKlE0t97G82Syyg3DVkGuYOIw5qSrDmGhYt26anaM2+L0apDjprhyE8tUXEUKFCJ91VTzF/qrGuO
YDTi0Rv5gPD70owjqMLp6adqLuBwyGA4mVdKpvvf5UctK9hrRcB8WXFtzXZOX/T9VRMYBL7499I7
ANHEkfM+kCxCKI4bSyCOYA2jZbropCCtwxH3Vl0HChOcSW+GpgASIZgUsd1Nwn8qrI+DHTinjcu1
zW+a+cc6DIpNplZihtrst6bSECtKN7nr5QYqDnEOVw3sVqpxeOZEDBAWMYzAxvpJz/5hNu7FPBWQ
F8dctvyBfhb7OIBaX34jcTYXJ8BqIFNO8KTbgtDWSlqd5/wNrOVllHL8bpHaBlzmkyAa9BQaGQQk
jGQjQ8qMetISPiLEHpYACMw73yWDTLskrYf+XBR639nVJ2mgaaX5zWXj0P+hKItjBFAEq6/h+1NZ
E0ztqTuGwdzjPQ1o04/yaaLXXbgOqY21AJ+h1go/TQvjzoM50g9cicWS+neNcRvzCQ6I2l3OIKRw
nV55/9zRTKmZwav2My1yQPQL45Oe3of+tOJcjqQXfdGT3cNVhwvIT7MmZ3k+0Sx6qEwRKo3qr2bX
bDWe36Q7qzvqZ9LO3Y/4Zh0RijX9T96C6JsVPtWn/kbVlyHS5zxf7c5N8VEGgbtotNBv5Fmumurh
HKiEEoDcaQFZLiQFoYo6kr/QSSIFJlFmx9Fgwm3/SI9GyFzzcBJ62U/NlrfkTv8lHeAsxzjNbV4l
lZpYUhHYDfkGW4AyuIHEO7P7G9DbvlNqf7LYvnyLv1OvyVZwc9UwiNl5JoA/JuDjLdW0Ozd2opcq
0yyV7nu3uOgpQ9y78vQpKNblO+vy2A8qJoC0DT+hcX0tLTinPTlpyVWAimzn0Vu9XDIiWSYXZD2F
h1rWMcqNL2QmzIAsm65C8Zt9OcMdxJyorS3RweUh1xpYlGMsk0EJDtglB5q6eYgNiF5wbJkz/EQK
+AfaK0/QPnl6fxSMDpxn1W5mQyPbND3Ao3IdzOAakCan+tofa4pkm7czpeYUtBgXuC+bcGTZeWNX
WDFrNF/dbfrkQqHh9ecl/+EzJ2ud7krSoFYSP4LzMc/rIMUDa32PhsrExVco/HRqW+6f2aqNujDg
tNSM8SyzwWb00STY2f5q3bESnr87oDRHyt3VSr5aKeg+4t0evBTTjJ1K/X6yZHFzNeOHdDV1CNGZ
Bzu/lTiWIyoPIQM1JehSr7SCffZk2nbwiGg2nXPcRM7DxNzUMy6MPjbzMJ2xOvp5XgW4A5f8b5En
GkEOOs15eYrVYyRD1aG5VvmAOqY4diqYiuoiM2bfPkS4xP55ydzpjLJmKU/NQkb9Hv40OekTP6rT
wmTaeAmAMgoFjquk6gbIjzIFJtEDLI8iEqBwhCRg/Zo3zyu0daha+0AUid3MrzX4oCoaD4NMlL5I
/nydfxJAmolrd0CLHP00Dutv/6d9b3QlueyODdRcX67lfqbG9wSYIZ2nlsUF0b4ZeNgeLZtaPk9r
BYydCv/e/OI69/0Qe6FlnowQam+OvXBA/jS96D8Ld6ewPFUWBcoWMbOCSysR+/X2IkWKVBGcetbe
eHp2+wxlsW16Qurl9bVT4bK5Q9cUt+NFEeTynGMpx3m5rteO8luqoL1MppKIRgYfYsjDOGlQ7WWA
HT4H5Jxd5jlmPdAQpd6xC7pxa4+lD47dfH6vHuuLk6vmMTF+gZD/u5JPT90sTbV1MIwdjfVLyg2A
fkGgVpIv3EP34/krx6UE51/ZZ92tKOqoLHNt93coRHoxXEWB/GwpEwV9LbfxRILmEnXWNVgp/giG
4/sUdD7XG+nN/sttqtrSh6JfHI6+V3E+HmUcdMLIxzFNhoG7g+LmJXMzfBqA61FAS00h5uxJYFs+
/+fz3R+q2tfL+D4XuPlhtwu3R1R7RUIPzuUH61XcglRQAe8wi1kOntm+ahsKwHWNE/deYg6ba5yI
FGgs6stR26mlbDHUbQKUP4fcpcg7O2/SXKNlqFNKclApKJHyk/oQNZrLXOz67WZ4mD30XezO+98Z
EnBs55YUmPfibGOKueiTXHXGLnQyUwUWXggdHKUFrUAW3k15Xs/vWGUXDFrN3b7N5a+SGwdlquwh
QbyU/j950XeXyO6SUxPm9MmihBZHDk2Z8G6ZRQq2c1CFcvT8JeZrkjgdQ8oNi9GRSHtgCdAWwjoQ
KAULDza6jKaXPleG1q7bFT/VKXKCVjYtn2MELkcDzIw2ZyXiRQXR7DODeatO4tjgQlA3ZjHR3uMO
wSak+J8mguK7yjW4AmMQiDnVEJvuYPmO423kvKox8K9slwLIDewJHTxqX3JrRfvAeKWl8GVDCt2S
J75SbIs+TK6RyH5fabJtx4m7mMJv4gR4HHl/tat9Wm5m31ou2McgUmuWqBzwhoHiBK8EHXwsY6ua
5grz2TcvLtbgsLLwlV5b08BMTNUjKO5KZFcmUwHAylOAkTPgpbX0WEnjYwpbtTHHAXLh5qXSZ/u2
LVsEQcnuH19ZTnvCdVoR8PcqeiTc89WmRZ581ZwiiwEhzr+F4ltyoH83XoUhiEldZTHkn7RpzWpx
hiallob2+um4tHSnyvtP3/gWrkCvA5UEg2FW0a2apOLMHe7bxH4kyf06RpCgxWkZNfEoLDOsczy/
5xRjRUj1c24DzUb/RcagXfeysI/U4A6q/iOINxLRAQmjMolbk9huXy8KqyncMXcvG00ENwNJONKE
ndOl8Z5l2c8WHpteHCzejox+xUx+s5cRk40flOhueEO6MROYjx3uE5EKZmbmjWM6xIGG0rSlSQB1
ubOSpb3qwSu43RmBdJcv+EztTwKajlcslfJ8d+bYji6x/3mpVrc3qrGoNFJgvpErp21QXBrnD0CP
fFJNxxbaSsaFEV8cNw3yMhN1N5X8D7Lf8KQb8NFjfS0sq4VSQKwKrqiQUULSSrdUAmDFUOM95y7R
B44Pf1denlwalMO1Hrfh73xgziUyImDIP62AXfYXs6uX7QQk7KduYCacpYvauxhcpfH/D96v8Kn1
0rEQ0s+hVqhW1gJ4mrLQBjmGtuK71Tt145XTJQt4L4MJ+RHaocNO/NsyCOdvGdhLsbY7vdmL2TTq
4ph965M/v/OpW8mJM5Tx2G1Qft+daEdD3+qaUo9BvI/7w8EB7UIaIjIgzQHNX2HJRHrPR0aiRXQv
HorLwS1SH0LAEwvfBswj0WDa5H4Sz74+bQUmWGDEuGBkKN7eCRJDmsIuLbs8okpUSlDjbg/g6KH7
INx6w1grn7kk4OkNlM5lJghFTQzQEX9/Q+n+2QhLAnRxMJqgVpqVHdreiAxWiGQTJtZpd8FTo2JT
Ud0P6NOFbqF6lOG9n5R7assoqe9dOLoru1E4TnZwLoQAjTnSWuv+xTzXCLz2cjC7UzQuQAU0PLnG
0OVYaTuJRBhqsFVr1Au7EWaKGYMuePpRKGTytcwqL29qtUz42omWSL8cfhjkChvBfTvBcqeNr/XA
RAseOsKY7+1tFTUnt48Nc/YSpjtWgvtaigka1GpJszsfQ7i83JMFe79AO9q0VybEsbRGoXRPEWcQ
IMpLCD0Vmf7hEbDPNncKao7BoBO2Mmlg6zXpLcdG+AZeuYHVCuWkPrXgGBVPECPTDEiOXrpWxryr
0RL4E0tzaWhKt8QmK6ythdx0ozYg7zrrbL/imN94OjlXfCnJAwqc4GUpescIewhPOYRrTfub9E3H
q3c+2fXGLRBzHXRj8XzTuSZRuM3S1EuYU2Zw0XZsbgUeRK/ISe+I5+beb7RVtzs2QeQKinoNFODd
efefa8Ty9h9npCefi581ecGtu2pt2XHzKmyuGPnIOlaj324BWmT+jlR8KrF3X3KbkALcL7XcB97r
9vk6p0CyU1/zA5rHYnFfcF+9EA+UeitAeHlycUfIRN2kGRspmlkfDTHSmX0Nja7+GIDU5Dy8UwcI
UDZTg5s7wXCnDw+I2B8r4UEJE2+iA74DnGV3hD2MeSPXHfgqzN4jkQzBfLpMWlFQ4E4gbp+qo1Jo
uE/6qJj76ALCAI+RZaZetZfMAzt3G/GZPj52H0Oem5NNNto3NHCQGLdxE/B0iGjC5n749u2UbWB9
9ItTewk4M1dldv57nlp2M/e7g7IzO7DLmgzcYc1RS4d2Ku7MZwaaFzA1S625DDFXJkw0Bx+oci2G
WhFkI4BI1UBpMaPlqyqzSfU5WVPbbjwQmnDF9kIua6lqxEhLMl8uDtx9LMxpfPaAek4SZ25mo07a
pahWkTrBFIqc1rCeaeM3IPrSAAWZkYCL5w3eUzl9Rbnrdd8pBcFmV27IYcsYSmlLLr7MRuYzt7Sf
U2LQI6GAruuOWM0xW2mk9BmG+S+T4tmR7qAZzi4iQ4sniezZFasrMVAeVAw4aeE+y/Wt0V0VhqY8
sy4f5flbAjych/L7magcvKiVm+M9I8hDEK9rrIpHceUDq1s0c4fPZ1ry6oVfGj8FwyMSdppUN9VK
F9DLC3vkv3NjTUYogdxGQUwVJpLJQ1GwoGvpaGaeH6NccMMimMFMVbpaQpdGLIrCluvquNlMxiog
z52fIaj/OYvg8tLBb+na50KMe3IATtkt5hrZIMcyB5w5mrgkrM2DNpTcnu6pDr2PX/D9Oy0nutxc
XyoUt9CuAG4fQ7rSmuPcFFzKE7ujXI6nIbHhcXeVz1J72kAB2t6HFGI19L0Ifb5GHGJpiKDYiyEX
fVCKZgEGW+D9ues0DrZ6YLyf9cgGm4zjeFbdBXlTV9s13HV+cr+UGMTU5rEJ+KXv4ugxykEF7SGg
0CxOhgrdBdISqfP/5HwjT+W4NtHlv3zzge7KEMRUvKCuhuIjdGjr9gDujb2gpH+fUrb+26Aak9Ys
L40Tk8bdbEVRbhE1Sl3VytY16M6wNDkotiktk/Q5VtIcuFu5kTo+xJaUUgLmR5M0MinDtIICwJrW
Qy/sMVa8X5pSG0w8afRbAPu4ROHCQaduHHbbg/ynUFdM+qRMsaev0WqUUvSkQ7F0VO3VCyjXVZDf
mGdePvNVV+REWM4kneGhv/2Cujb0m5JacTVpm/KbVMPA8Lda9X0PhncQcvUIBgZVkRDL9fNb8IL4
XDj7aRlUtLRHck4xbLIVFPsravCF6XcHG1yyfI9k05ON8yLCE1IlXhwUU3apieLlB9fKLiTp6CPi
Nl/EnujSXWnY7HBC6wfMvtT8CSSm5dRUNyxJUtdYiFwet74GKdjm10NBfTNCYJXfwBBzfOls8ek0
QC5LPi8qlq33/WcVI6LX1LZifCnetP/prS9b8WDaPrUziZYWamP4KuzC3vp93rsD3mH++esI59QS
VN/5iK9CuiODifvY7+evcLNvxAVQEzzkZy8MoYuOYpTO28Ah98Vhk8UNIhQfXxeGkTade2osBZfQ
mhXbk1xYnpMtTRrIG2Z6u2DmI+okkf65CbyveEsV53dGORtZ6O0BWNRHIlfvh3L81qRLyBAIicY5
Tn+a7qCXVoN7ECGTVkZrEoJJOkIOZTJ6VNTQjSUKGFKrX9GIzUhbPHZwcNnu4ittN4fOYyJx5iLo
tom/Y9oC32suj3IBcKqYrlPN16HnAwzBrC6Zx1IwLjCyAbv/qfLTa4BZutVUpgsWlbaL7PvfOlai
EgCB5SMGF+A5wlNVdehw1223G5zbGHkyr4KzZ9uNzMAj47JlF0cIJDjPjD7/5R6wqcZt67YvpMiP
fBHq5LecXqEfmBYUlV7/rQHpAIyqCRL4uQraNKBLdltxA7W+49PqbKQlNLtbP8wDHhiXIig84dXM
anqOzWVkmIW3ukNv6PvlEOhEjFVRDd5xSM184hYPwNKYyazrJmCuvYvF/8S/+3UVikKb5N0XjAVO
fBzyIR5oaP0N4uhp1VrzlMJaE+ytGTTbJWP5VAzjHuD0kEp3MifvCrvNu/OvRHWnt2QySz3LQ6P5
MYO/7SMmlZ/bXTK/FxO6JjH78wXIcXqGH1hxmgIIkMw126GwZnkQh5f7+2LLu63XIgL+FQ1amMBA
kmAa+4yNMUZi+1v33TlgUlhNVjPIgN8iXpVzwwsonZbsSN/gyfGIx191Zce5LcsVJv3Xzs49VMa6
IpegfXifIGE9L/XrnP+l/VWeErM2cXZMngqM6LLyxfzeyz9+gRG0G+yrgke6QpElM9OWuUK/Jaht
yDAbGoKidw5cmDYfpGeKdhfetxaQY3jQvepj9SvnIXArGwJiwCZ5i0qY3fwwHN6UYw8jfHSmbfJZ
HbQ3yfVQ8P5x4avGSuTbNhUGpIN/r3CJJ38vV6qNnOfAiEI1PLeeoNcmI1BEG1HoQahLaIysxp05
AlQlNH1rRuxlZ7Guzu2p+g2kcU37tdJPRgKKZHGPT51olYvvAResX/2yCNq1yzSsharnLWv0VJT2
rK046U7Sb2vxoQsf/LSQV9bbuCfFldcZ+ZslsppwdKMoctqrXMYdgFTO2eJCVB4wbaVmJGo6u6Tw
Yn1ZkSXVn7sT2aO3r4M7EscJeTcmBU7MgQUMRz5UdZDSfbB532wYNJhMoG7viqPJ2qEjh5htr3fu
BSc1fBhogW6Cyh8RORZSeRNYMHH3fkXRI5GJSjmX3Gz5RLmffbOkw+5BM27hMzeRKb4xz4OyXlrs
mUNRf9dQcDf74VjAt/LYY6MqHrAD+2esP9KNHfxvupcQHdACI4uplBEyWniwhZX2Zob+FltGKIs5
hpAjoGJ3qBNmLE5Tnhmv2RlSyTsCRtK5PhZq0zOIOb8D0hzmYYYS4NLYwA0ZMgDmEJjjHwxtdpuH
01AaK4azHpQ43CTkgZ/xk9geWJcp9qrkwePtXsb3QZNNNVEfOs1/hSVsgUX19g2ZWhuS38TgluWH
V0wJVCFDbwcZ1YH+J33xlzrUpz0GZODwP2MCEXjMf4YYqsjgwKeQpDz17pfcgZug68dkwqSOPh3Y
OBT9siZJxqUOddqWRztILc5uWu4nGfAHJuVjl3mn1z3oOooSauiyEzP+iMW+9Wc0rOviFYtz99Qf
XoeSh+32Pi99qhZQwx+jlDTSi19obG/3/1DBYy2lHIuISRhRmkC4df4+KKXKMbnMS/tZIIb/XA9+
VCqqz04TEc5RBIZmWYeviyazuU9BtVZrPi/+YcgJ8r4NAa2RMFpM3m4j09GjrOtxQKGgv5K0iu+n
wXKEmBiJRVLTlLJu9Rlfh5bF/39hPcA3zp6Z7wak4xi+4Ry/aB1CAV8Jvv8w+uHGamr8FriLKGTk
680+v8NyNf2a0GUUZ9z2gjoYj2NNdpBrsLIfii7io6hy06/ZfsAmkfZdU4jszciTY+OlsRmZOU0Z
yPt1LyzJrTkj8X9KZ8Vst/Mz+v+4wNlWUZJzP4KXusbCjD6pbFO/wNRFi5ncP8sWDa28XX8a20J3
H7ZcMyyCY++PIlG1q6TqzmtSfiAaXkacgS+h7bug7EkMk3ColFtQBIGO7cRaA9Lc5ft1Zs4+RlDk
me5HAleO4jX3dnAZBImzAJ7OhJ9Az9LOzOV4gRBqe/c/mG3GPElG63VqTD9BpMwask5fNA7uZr/Y
I3RrsGWfgdoRn9HYmgArsEJ7o/TUxoPESw1/NdA3srcT572I+WRkeVC9U1vsZ6DiDw0OLFhl0Yfc
DsBRlsvd+d7UfTc3Jeq/qRRnXFE+RIZdRgG6/8+H0L8k9CdCllqI0JOZdf2WBuNkIhThMAumrxMh
VYGEOkXSIMmtZHRfqP8JWuYNHrVGvRmIY1CVtYGVkd2q269BkPHzUX3vZuyCYqoJPYp/wG5xeBrY
fJzfh+EL4xXg0AGEKCmg8aBsn3z94o6EXjRb5bfG3oxzgKCjSz4IhXiCh1/Q1DXXaCm10sMgkeRv
P3xAmCYezJVrHCjK8qdqlWkYAsAEKmYLaUTv4LWubQuQ66YArgUfNBCcPJfMstJr5ruOnZZW08uF
teT+yJtwEkTmaClziBlv6+fdPzdh7tpnApYv5wTF2gfKmD++IYmitLb6FpPMW5XgcnO6OeDeZRRt
l412oMIK0E5n0P6zafB+Oa253s7lZmKcIF6R0XjH8x++l9zYguZCn3Hk+JzkctAeWLhxT9HqllSH
nbFRQbS4is7kO4fz4dL020AV8x3BOK0TU6x+nbeIRaFw2YY/BTAmZyIdZELnTfE5OZyKmhk59Jnu
USXIuE/olqsZyeQ/712ZSpLgz503IggCIvRbq2UlHwFdZwtRU8+xzp6knSYnPkeRA0uXWBkljMao
RybACQ29VqstgcswohT3x3Cdr80ojU45+zzNRLekdv946F5lfNaqaFyYkKji96aLy5MFV4rKkoee
Y+XthTgdPtqlzRMbKwpuRNXMKRMrSAKipn7f3/erkPdH1A2Z1qm1RL5+JrP/EzhkRIWfWWUWKHz1
el+I/u/gnjT+axJkxlQbOgfBnbuvp3MX6TtzNLQvm+MM8nASRCbWjTy/MknuZ6AF3RCBwqj9h/O7
HMvpo8q9jbXYy7VYJ5U5rY0Pm2NEN/d9N7OyP8KGMT4APpHXfNU3eN/MNsICyf67Id+/hUVO5BNT
y4AzkuHl11gs/6VhvDPHYACatRLFdzGJEggNIO9ujbsarGB+kXhDntjhuc6dKGlOGxMwx36Tl4lq
2ceovBn2u3dSNaTJlDDEhMvTBcwc+dd8O6Ro9v61kR7qUAVaFSKQIYoLhKWtAuEgecFpwnhnC8w4
KTNJgdcS/ypxubTgulgupe0YMaRt3ch70541NTINiZPMRosq1vqVw/r71FjLaFGAKsmxvGTMZh53
AClLO+qSXEf5IOtMTvSDwR2N2Xy1FIGeq3bN42KKRv1ZhPQxaXZstxKWqyFQnUPOY5Ix3t6tTKlE
3vBj7B4bnMNjjr2KkVx9YJbQn8T/jpscZOAuYn3ZSt0CIzdKCYljJqGaldUonaDeBAsrl8NWGf6o
tYyA1Jj0DYJYr/LXwuX1OvzUPmraBz9ruFEvpyaq9id7gu60V0eojKS8beowh9OZJ9/Fi6l/MHmX
vBsrUmKPUV9XEoKT5qLIL/kmRFz3h46hSNFJNwLK1ru259gTDTezJuGpBG182Rtkc9mXFC20azFq
1evs8b8dg9DsLLHJHK2Ry0p9KYyVF5Itgd5wMONvz1IqaTSWau5nUgakBL8MQvbYwuERoqSTAnCb
LvbIMIup/K9Hj2hhNZ2nf9lbjozoEGNqH2S+b25fqcQ2q94A3yLJh7UAvDk7D44Q/RFAJ+qlBibV
pJiVTLrJ2Opt1GwLYVmgdhvs36iSIS91gct8qXGEZafYnIB0u2hpi9uXnOye6b3K2Nq3SKHSB2W6
nGVfGcjg4mSQNl3sLH9vvc4L9JFup6sMpbvoeXBLKo/7OwLW5lIuPRmBLxSgL/E92nW2EfXpeUYp
8x/RLRtWNP8xUEIp+vzRXHw9IUy7bvax/XiWauQJityKrFdgRFZdBLso5bbgXaDaelgRil8BLb7t
WqtVPc9spnQtjpSC00h03U+5SCBDbZuv/SRL3uSXB4hcdxsqqbgtvC2/Tuv0Ws7nE7WnLEUMNEZD
VMVm6stBjogjbaK4fGXT/cfYZAN2GJMxPJhGIajJ8E3h0XedIxt2Ba1UfV/OoHQwpOPR11/Bx99f
jqqr3a2MERUPiSTXjJehY9Vi4etDRYA1sty0DJP0e5JO1ozJoz86wBNr8Hu1NJnuJoadf/s8SOK0
sir64Oas7DHFGthHvAXKgggwP5yvXuJtgzPZ8LZIddyJyCkHKH6adxJNc7/uMT4qorGnr6Ss8qo1
4fNBAldtSSRr0NhzNQLxW5xvN/8mZG5SdMXYnS4VJ5TRS0ni8Rh6aHgdW9doDPypwOD9N2GoGtj3
9nU/6H4I8e1ALW17vzBFV4Tdpdt6SjWFySEDx0WH8lTx+/pwo3KATa+zsJVW/MwqpQR2fCm7G2Uw
fGRNxBSXXG6IDa49QozPlUH6FuMPOpkYr7yrAdS1iTATERP6Irk=
`protect end_protected

