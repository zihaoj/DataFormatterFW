

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
igspxRBvZTl/586mNdrH4BQX+itgOCeZ1xOzm9aZbUvP0UoMU5TvTDXkimIeEenF+LD0DgFrCICq
OyRbSMJ7JQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YRQhrmSAroOiD1bgLLadPnYM04gJV4uAj+82+Xbog+8blLhXTxB3/UTJk8MmcIYY+btdA2Mkcr4W
vOZ+b/TBUytWrSyGdj8/SUu4yCdpwBDZ0YEJXp9vZU0zfysPYTQO1RtloeHeOljj/nxzfU8JO+Db
qpN6CPtIH+ilgYQ6gDw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
N2BeVmmjyQ/CsQIE4JZ/yf8177W/13UJcP7zdeLaTDJri1seNWBmKCyWCyq18RPFjQfO0/txaT35
bdyW6sQRFxRssWbwWh4Y6YEhtQ/q6OP4ZAFAVv0r007J/OA8jdphubQQQm1eh5B/XPtFvUv++cTE
KoEIuebQXW6fyrLDhj7Yp5dP65WkU3tcUEhz8uWaA3xrs7vfI/4Crr8suNQattesIPJ2JthlzmSO
Xneb0NLqYo3RuKOD8o2Ihf5fg2UZo0rCS9si754eyanQ6L+9Zd4JvSAvXdqAASvkbV/gHP7/3I/s
1R7KAdadkd9Dx84J6YS6lZchMA770COqUFFzlw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sAn7OmpbNaLGVe3KSsDOYCI1YxIuh1s83IP3Je5Wm4JFkRSwsgP9UCFROmwCdcvkDDnFuq8ysvfR
9j6WvsgNhxE9ciKJnL+R8zmgPjxOzQ8U/BHS5f9y44rdX2MmdwTijgqaWkbE9fMEmn/MxvG3H3dX
fN2OWLeFpOulkej1TV0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NUQUiunqpt4DSM9cFCfu3SaZP7zUQxovsQqbP/L87McvkmjHlaqmgcLM8LwgY3+bovOQ8ifV3wPZ
VbFoh18SQNmbCCpwtdCEgauh7i3rOjM56Gar2P8O0c/bs1hx0wHagO1XbXdyic3a4Wjr9ph7+hja
Vmnb8Oh3ootlsg46NA3ZsMiCPanLiaUd47D0ujs7ZqQhcCtDS4wuN97QhDxcmc5PIXSc8BAXPLOy
ECyR20WFQ382HJW2V7WyKnRRIuJzb5QI9bfRoxKRmNJY5phbr1npTBGzFUDdQEieanhUaXupH0Be
uttrMyA7VuFJZINdLEhfDKM6bw0ZQcBF7Ihfqg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6336)
`protect data_block
IGgSlau9R88LlFKk0c7E0hS1NWdMHRZcY26IlIKIBLomceWfL3UdJFG7J9F5i8E6YU9IWOtzt/pt
SX321iUOlt4pK1e3Gt2AHYj9GH+/7Scyz9yQJRdDPBJVoVxGn08+WixUfuiHHmMNa1SdmuNfO0gy
1ZuIO82AcWrBH2mfZjziFvy1fDLl1BluNK7xOTCTedkDgpeHkJjGsfooWNUcGJFbd2xSovXEUDDE
7vsRwGhjWT2xWQWs048taylMjO9NQ6KhJGd4vkUHcq36DzhRoPTP88u+Uw7/fnWTUCvAqPFJ8vqC
bGDciA7t1ATuBdC3mp2T2ygm7c5NSMTT3TmMMuYM5sZHHj+dRG+Bh6Kzrl/RlMko8y7ZNEkqs128
8xx9pPUawTgt3StCj3N/1DQwRQYx+ZdE5e2lfQKdrWLCMcXFE57aQSHx0pbW4+bu2TexA5BuAmJh
AnxwiVxmbpIeOM9v8cubZtAfXlmXyhQb/TEhKEzniFLOP3xBDjcyzvflHMF5JgOPdrwvu+mix9HW
7miZVOHlmRfnXGKV2BRTMC6uaPTq9JZ4IjRMWrh2CvCP1GMLQNSchzxoZeV4Jmc1isuOagcU0NhI
GHmh8krX1sAbo3F0PFIWAZEISjLW9143EG7DqQf752RNxvjtTpqw5LN+OS/eCUJpLBhD8yWECyim
1AZfbNHpglizVrDapnxpOHqNMCKF5bv53YMYFOT2AGXi8nMCI/VQs1qg54sQDlkzmVDBnQ14nN0r
avqRzPqunrj+LP3w7pKDo+9rQ7poIf79U9M+xE1WjveG6c8C5nGgsBQlZ7MNNa/25utVvAq7EIsm
4gyFFtVgnUThgmBgR6vOo4J9lRwaCOid0eQdnvcUyhoRaLhdenXai6wG0ggLdLJm+hwttFnXmZxV
gyxSG3GuIUPNe1WHjB67V9MOa/dVo0a5C4AZgFAVBACbphTMNRDIXpd4dTyJNAQC3pyWRWCmMV5/
QQsAbb5cXcSZh/1c07lM7ajpoygN+yLTBnwt4vgbwepxlZgvgkNEphdJZjH++tGxJ+9J/m1jqL+/
x0PdOuyU/7uMIsFKEDOe9NHt1T3xohEguJ5eI3a2rEz6cCMs62bHAzcYMskzE27qZ7V+2friTkxz
wO+7Ba9Z+R4m4z1Koj7kVVuA+CAuO+BOV2gN1jT2nAMBhY71slR+YgweZqd73YIJWPNlDWp5EFhK
NqqsGKKdcYfL63umTwcDtW4OwyCbE3PMkIas3VJBkOCix6QJWI+EkLRS7k7jdVG7OVEf0HlQdkcX
yxD/NiqvNnA8S8WydQBZhVJy4UdsPjgKImsPRsH1i/dE/GSbz+QWdFOM8GeIdYWTPhxj0lCCe1Gi
gvFTWv2uDkv932ZciMdUK7A2g1PPLJCJmiLSi3H4NeZjiReI+jfdoSQzguQ6YgUYxuqLVphIR8Re
eaJiOjlJRWjd6uB4CIaWigKp+Ku0qCiL7Gi1eRaGOt5gMsj8wNNkfjBAefZZC+t5PCTjClhdF89p
6sVfyAB6UiMmTrWxPjrackqKEiphoL1f9KPe2aa2Od5ju0kLADRIA9PJ0GinLVZVtpLZ63CrUK/q
6MIUzyYXN4VKWU055vtbjjpknz+KmRdybVNqLYHYitERGcHqNIbAP6vHEebtdNjs0/M50eUYhL/W
1JwLRI1A+hiATP0m48S5w313/Xc6v7QO5DrUxCR6s8n5ogjSiRLbuw9HRYphB8M+jeQAaILxqpvS
mpAfiPy9td4tzRhANqyA66otJ8oDr+5oYJefQlPDHwYX+CkQzbBwPGM+JpFF7MP779mCmLY13L8i
DuMaermJRqCqOujetYad/H/v5ZfmnIKgmQdOhno9B8kiRLteear7NIcCHtzgjeZPK8S2LfC20b/9
Dxu7ClNy2t2mV8NBb3vZu2ogqVFPcoQsvw6jphELJWoufZDhlv5Pp18Ia0PIlQ+2qRvB3vCWf3Uw
g4hyNTqyk657LgKHymRSgafjGGK6bvsCz3WUCPWFmsDS3D3LVug0lJNxwtbVrKnd4UAaAYEHWYZp
Q2c/QMkH/gaHG50f0qzP6rWRi1vIZH2n+FMT36k7rw3zmuG6yRvDH1MHW/wlbMXMroCiUHLkdl5V
9seseFyZIQK+QCo9jUIaToWTAYFRj/edAfq1Z6qX2sjXmSEmJkqpF/Giu/xB+mZjFnDkZd+JkEVd
ZJjE5lAT0QToiGoIqrMrKa0yZTSFz15eTSIJuMMewQYecT2s6ZbO/DCPI2FzsPecmtymxdUAHjNu
lEq1PSnJuT1HGsMYJqsUfRN0ENjQ/+tU3QNM6UWn7mGsdzP9EnTzAHqtwjiE/c8CnvgUGzfwNVlC
jFj8wcRSYkJf3BKy2qjjiadTbjWDd1YcyxpKuivJKWZw9/sGmkL8v4qa27TF1viiptB7GgD32C67
7MDg4MEnbGgse60bKSO3aNlg7fHmmDw6h8j/UfsVLrUPHgV0bm4QHPGhnY1oEKQgDz3eFaXBtIvY
2qOdCK4Sal1BESyp40krtyGynfaq+lSGuRt4jsoBvJzSd1FbQzLKQUgEe8zbVnk99iVDjaj9EkB2
cH9kvtVFjtl0oGvjJSSGQo850o4bTVPcBs/p79jdH7gTcNzVP/PwAWT7z22p+mCH0I+feft6VgMQ
ydoqtZ1n0hP0IEXqjmB3Juh+19t5zpwl07AldPC9QH4TH/Mb0GxZBPemyZ3evkF9ZdYwI+Jf8zbf
GSMDKQZlV34ysgpP22iID6zGAZ/s2OOK0yw2at56SO/X+wA1FXkPPCejmNmWLjv/s7OtBvyKF5Ow
6DoAds0GJWRNVzcj4QeRKRqIZmhT1HUR6nGctGQYZdj/Vookvc5bTbzMtzKrsYKcvVVK20R6utEH
0AcuTcSG+sR8iQBoYfc9oiqRVgwL4h6XZNxlOR3jNVou9v3mBEjMbMaHYVCy94MWLSTSZcHuQVOs
3Mwv58tFDWbWMKPEqBNNsOgwEapbtlXA3Rjl7H8AZrzBeZDh99fY5AQBNhX6MDrGkzhJSwjy1m/o
bdPJEyVCCsKClweoSUJj3bMifmMkHGRuG5V6mTT2OmvrrGNRd+rJSaUN2q0M/VNAVDz0DhC3iAfm
GgreH56XEWQOGC0Xlj+xom1H5rXVnXIh8r8IAw3SgS6wTj3q7D++Abb9qfhTz49NqXLKfYScX/8/
itChWeAzkxg1WwUYkZ0sp0bdOS11MzzOWlxjnBdGnkFwhoadtCC1fsglMxRPditcqZ2m2TEa3aGe
LxfvotFN5bClMfzKgof/SvrePzHWHyvw4thg5ach/9I4ebnkr4SfweqKIUWcR26OpVv0FPwGucOk
p3l/XZP4GQsSYeT6sMFq1ZZzTLcrJXX6LVPpLX0OGZFLqSCrLTopua2nlS52UHhkZmWbNhWVSUFW
gzzeeNoPybzGeHY2GcGsOHHRoDh38qOTz/fiuTURRcd+6OtWnqutRx0rP+vd3MKWXnd2Q8nEx+N5
VFRvsvMtBPYaRdNEV6W8qMuhSOArCVuQ1FYOAseAupMqdy42zt2kD/C7m0dGnDAZKkcFTdkBiDC5
ew7JrqFiXrwQtH/LdhL73ZOWZkWdSnKTqEYj608P0YO9Y6CoeBs7Xpk/Uowewwn2h0DvqgJ8ck4P
tL/sSJZ9ES1/cIfQWQmg7w9eNsR9i+lc1hBDeag0B8N/GzElgbmqlKM+prfLgVhPjnFgLduz+LYl
+rbRQfMqyOtIQznSrHSd1vwBbkf/hixiiC2hHHHYONqXhNJquAxoX7MksJqOpJinVYSKh5FqAwXF
ko9SstJxVNrJg1Uo2h4svf4dcJQBBoL7t0zdkDeV//SWW66EwuK9ja3FtzRURspsfV3JNgfdmY4i
1rOTBAvzXeAGDGdDRS/4nzzm5kwA/vJjHYsmH4tUYcttv2AbErbMm5VkNmgh2VxcLB3xiUteIZRt
0t9CcuY7+sTAdPDbIHrPt4Ul3ZkJs/Cqr7dX+48d/U9GfsKQqsSRWxF9367Rf/7x3Jc43svqm4oT
Pex7yqKL8qNWGFKxYsWIFL9ZFP4oIQpcruPZs+X2oggC7426iEKuZxRbV8pF/OWOC6cOyzuU5SRP
nqiWTO5+syy8GwYEv3BfwjSLtAZawisREjTi+xZ2vK0nxdHt6IVz3aQz417HFx4Ckocx60QYwZIy
v6QIu0DzCnBGfDvKs99yauhkZI6qGLad6pTcVthkfOOzt8wJG3G+6bspQd22Cj9S2prfmPggBLOk
T0BtVLyCqKnN7HBUEgbsX9KSZj4WlpfFplZikIKWhfjMBuaRpKYcAgV9zuVoMTbJ2neIzqQC5TqC
4h3D0pKO3qr2FO1iLdif0Z1+Nm/ZIAoKy2MpHS+JpFmqYA2pk8xjp2SiuafA4iNpcmQEpxkXZ52N
7APkNcaLru0wrzZjGs1fzEtD1lYmD5tC/xVM16Kn1t/PPma1cagc0hCD/FN+59xxBGB1G54NWJaf
t93DrRDRhNOC6/leUNFXh9+k8rvq9vyAVrwC/4Wg+jEKzHqi97gjo8yL09zt4xSbo1Bjd0Q5SyU3
xEoKq325xDyYyVYdTZoMdCrezrGjc2xp85DjHJabVRDCdQIofCG7pwkHH86/oZdFXRcNgH+cCD0B
2xld+b0xDr7zvbo6vy2WHWI8xHPrBL8j8n8yHYasRdVJQea/5ak7m4g7Y8dSfWXFiHrvbFQq6fyN
V9qGAKV7aF/YyfSqwHDNTtxkBU2OIaMHGauFviqzDwXvOaKOWTrq07o1+FvPmVHTzZbtMrvKEHIX
v4OrPA/3TJ76HJQ7aJqyIP09d4XuqohgYBjqlylxTU2qR3k3J5LYmunqJjS9SAvGg+J/GACdW9Z4
pucM0qRpHcYCO2Kxk1KEIY2VhRYhVCNujXSvy29VNj32Y7HO7n+ZkA+hJ/a3uUkTfb8NP1uip/mh
w3oLFJP8hdaSjFmifclW+VFqd/vq0uiOjl0VAt45CCAAJ/8Ul/8FffV5gSrqZPHzeNMchHoFBRnN
85Fardve3iG1xIq3sTlnQqSwUMLrDupNncsas6VCMNow1wEQcx952lpKxsHKS6Eam6VqNxAVtNan
l6iJQ+NEXno9K1RSuIFT4YXjfrWeFCAaKJ+Q+pOplxzv52mN2rwr+U2dLKcnNz9eiUv4rg80ziJV
OsDajoT3slU1JpUKWchdbi81yEyVT/LUkZhym3uMMxmDCscizlwadZDtYC5Lhtdz6yc2d+iRyY6L
fJ5T8eQfUzNs93shwj4jm3R+gsRqhlUEsQkIe+iuIpPrXjcG0DYCNMhsybOa+OisC5rgXGmaNbqi
3LG2795j0NqiG1+fKKg7vlRMTdNQw1LGWrmakx1NSWFjEyDvEbHJNVJbrwpT/rhFHD9z2TuraT9A
uLt07yrFmNzoPtFccgWWGKDE1oqutyPy4esvYEz710wIW8VojQx9mY0xR1mdwImx0fcnvDm+0g71
lHFy3e/Kdx1xxOIpse206FKEZlUqQe0cinrktHp2G1tq70YMbC6xrDwxjcQAW/30JIXbZr1/A7Da
+cy3WzDmL2VZ9Rf8QVC5r3yv4MwFZDqPcUeKOTdB8xR4nSf+NTklI9MP3uQqR54mhG6f16o6Ms6e
IFfJd2gOBRBnyrBLoUKelmyu5gpqtmLiG86Xa02gurQrFlJa6PcfSQreqbCojsHO7qXj0biAaKaX
1yo3dDtnFs6fShcDh1CAFw9E1G4R32e+JKZ3bIqBnH7UrQbfJxgG/tjWtV3kmbAloF758bhhOI7v
Hz77Ze2u/DnbbIN7yON73BRRG6MmRnWGJoQ/IPWSZDl+eFDy9SQSKgrYjJCEF5olo10IScfw586e
cqi2lx8r8jKrsIM05lMTR88044CaLMjvoHME7vLCZmmTZXE/wmJVZoZw96TTWLqVXguxntolsVpw
OI1rFRKJbtS5oqHx4YOdGn6xVygWzK5pLH6Tfgv8sV0v2QL5F7uE+pfBdswaPOJgQR9YCJgOHa0w
P+Qaybo2BOnsrQR8jZXmp2ahaPjpZoKT9jo1xuiglR0E3mD6fiZOaBkH3hv+JR/GtR3Ttrdd2ZFn
EX9Rrkq7p4Q7DVCcCmmv7Vm07PdgVD+Aw/JYwxKAeUBa5lK2HmtgyRxWrKisBFSOEekzUj+/jFg8
mXPXPqO+laaF/m4ClTIavRH/AEI6thv0RdqKgrIS2AXb0ly0y6lkvxqpboTFNgwg9XFzbPcfQK7R
yee+TcJpUlk1rTrkJTEo7TyrPeUbfPWLnxsYr1eXFjrJ+NHdYL4YaZki7MgTEcPmFO+HlJ8DImC0
eG9S+Z2zCMaklAjIB4gbDWJrlxGs68o0vOYVpXN8uyGWum5Mbr0NdoAzqfgDuOXIrUIa5oLO2yeA
ULQpT4kd2otq3IDszF0/2t2XBE8GWB32QOZLmvgxC4O49FZCrOpg7iHtwn3qdwuxWHb53RvaFxKw
sD3215EyU4HMlMHM007lfTbJvVK2ZxEvUzTGMjp/A1mCWZsNfK7CmZBeM4oeJEWyn8D8sxwqY9lT
7a8/WO2GNiuDw1fcSkhaY8H0lI8AIbb8zzNSnr66PISdX16dbnv8ngn5Rx5OOV6pROv8HdLaBt4j
Fn3w3VX1jtYcci4GuTkrdozS2zhol4aH9xJqSbHrqqbatM5713F4VJ7LWerttRPhLGQ+UqxsQQm2
kjebnh9LMNUuC0ShA2/fM/EcCoMRgMEa9KHAO9bpc2jFvZCKik1CXpwbG+9P5CsKZszb4Cd4l06X
+fhOPfH4Yb3SkCmkiw5L8fzzciMYMvqkIGwqk6uQGKmciEt7dSXxX5Qez1QV4nRFG9BmpWYCGXBj
4j0VA2GbMBdPQfjB0m47ynWf7qEKrNoGJiA5bOTqWYoaGrnuJKpFhlXV2GJRt2lujVqp1T8br+Wo
Umaq8c4OtVyendAXQpFl/UOsrwnFL7O4jyLKGEy5kPrKNEPbw3ZGpt6+gtMJ6bCXCAkI6vKQoju2
0dzcEuZtCuEt081cXYXUajsBa+IaisOFLz86naPUyeqzdrINop7wUMNBp5KjuM/rJYSz1uQLWwcD
KV6JKFk6v72fKCBb/sQMY0936u2iL1pfBpgXwU4oH+/z1IRIeKMRlpSDNWjy+djGYj+1FU0R8pOs
MQihqbo7BagOy3+2BZbkmKg2Z05E/z5FSPGSWIgRxFtPLpOYX81/LjVT6dSnHb3HSAsCJkh8muw/
epBn/Fg37TbWyh3mvDdlyib4Cvhio7n1BJt4xNfzoDSbkwDg9xiF5vC04Kc+yIc0ZKd7gr+E/HI7
LBMntmPmyWRT7xIYjozltEz0YH2QbS3KsxPCOVDTJh1HaPUpDxrojYvv6HMSCwAXQEWJodvXwXR0
JF/78yGlcqB9uLde+nTu3lxkJAWgptZt5XcoTjdH84tsJEKVdjcD8XdnyAZBHjWilOBHyeje5GST
veO0CUuTUviM79lZ5JCXqQ2QFqeRLIxoBGBxc8U0vrRRBITEpGPqMyR/Gii3XE6E7H9JK3/H3j1D
MerLMdiM8XYGSVh5HCJvLKielcI+zFYitEhc7pA1LHk49gosdcM6WoiYm2mnKcLZCOrJLVv4ULtG
fJYMFrIhsits6OghIQGiTmvR7nHg8QytxowlbZgmxh3IiYs3PSW6UstnGdAe4FJpb4PG+Ik+uM6a
o5GdJxCT+o3jCaJwFLd8UzZmqrOdfysde+e4Wnblp7H2T/gM8jLxxc1xjP3IFVA0AtCIlFUxhJCu
4kwOiQuY4O3A1tUttXQJfPaZSB8coAdrv6peHWQWII8DpdwDBsPAw0d9RU7Thf/6fv8RjjBK29Xv
3nvod2pzbcI5cJhpe8VR5t0MJl6m88y+FaZDgpum69pirPF1dNOGTDu8apGyJ5pYnAy3x8CXkukn
M0WiU3F0Lw6uV0jNLATm/o/Okj/+y0S5+YXFHHc5F3u2uD4vVGyl2TzF8ZCejdAfo5UdcjobsGvO
xpjhliWznzs59kuC0PJj36pwkk5jY7KPIyOM9Opf/HS2JOMF7gqFiFu7oUF8rxswGvniGnC9r3vW
3uQHrR6Q/9HbhkmbYMhQqtcF/ym9YYxbIxARFryJPLFUnGtu05I/ElsQpa88WhNMB0D5XjFEx0Y7
HlMVwgzJldfCuW6EoenmDnMP/GdGg9fzAW6u0FzXgTIvCo4z/VlLf/8lWTGsRGyPPygBpWxJWIkI
NSk8mYmSbe5tOlTz2McYUQhMeD00BMkJJ2MbRC8Jf17Tyc9jx/INs2LHyYimqRMBgGFsVH+QJd2V
CsLL7hPBzxKf1maMIoc/c7XWzJTsQXkNoCGP2nsQH81xGCcnocnJ+pic9bNYP4ewZDvYt6Sjl62N
hl45orFf3Vk1GP2ZmYmnYmRlnIRIt0wuHV+6iUfSA3CUxbQvb9DkFtOs9r9KG0Lmzi7UL3wzNOkA
lj8bVi0nHRQN
`protect end_protected

