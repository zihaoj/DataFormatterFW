

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kOs6tXJzQbaly6q1YmMa5yYN9ESbbI4TG7psRElo+D3cUANPdAkUaP11Rtv6aQHEb2T1YtO9U+cF
QayzFykWaQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kpFYo8t+C5u1/YR4XqHEKItFVPkWlU8IwR+gPeKPSzKkec37IKe9K18s1a5/cEFm7diJTPXL7HF0
VohSaTQD/umF1kygcF2dRUpCZFxiW+tRJV/6A5p15sfIau6KYPTJ99Qood+MhSdY8SDBgJltxPv+
mPAUHnNV6iJTo40YZTA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nuHtvxJNEzsHpCj0HTDVYIIPhkVs3FpqR86RYOR+Lgls4vDSETQdcjLkJffsedVITnrjzagoC6OU
ZYtqIhFE+nAuFdTu+Nfeq0/XsIyypKDERqipYVA5oKT4O6e0B5f7WDKVLUdIXmxqGlNYI3n7xunu
KlmuCo/9Vx1SdRi2srcsPh7NAch5XDhhsoudnD3wThbSF8G6K9fDtg4OHGtZ1p0A9+kCEFOp6J3j
SDkl9VMjNadLGP8mDeN3Fxx3Q4QwBQclUhLnMg0EtEcKXjDtNvVjIRk9z41mT0ZkvwYpgMo0iEvl
2bB9KT6yQTFz8UeN2E2CGOaQRVi37eKhp+oVbA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BU698lf6zciIHkn7xp8lnUJyUCWQ0HaTNdk1/2z1r0hZZ2nF2bvMM7ti+v39w6AcGQwSTYVLbJgJ
MTQ3HSB+aKIwEwGoSPoWpUt78ixT6W8zYoLF9wlMTaeLUNOZ3MOViMI4RSZfgmfGn1xP8cG6lJWc
Ss0/U0d6OievndqJWLQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LIY0j2vauyVeQj3uiBvFvvm8E16QcWzsNq85IRlylxI6WJVeAqbjJ5OQYvJCBd0ynHfPWSkWL8Pu
cLuATqKC5J618+iWZIZpqlH3QDcCQT/k6zYzz0TWv7i0LLV+EftpiWlSVXka5RewWs0n5z0s0vmT
PPVkUjb1doz4k/HgJ1s81qAUT3zd+t38rGj7pUDz7LL8tzGsO2VhuAcS4TTIjIiRLaPZlyIBSrNU
RRDEgRXOXwNJqdKCAQ4/By1550ciPmC71ZUGFRTVnx2IqYfaKhJjEoNX+pHMIsNx034TrzeTz78k
EDcVF3CuWM+LXcdtLj3VkbgGr8yVX5oMz2u+aA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4256)
`protect data_block
reUeTIWVTh5m9fA2x6v/0sEzPKQdEvf436eCI5QX1WaaFa2okt8lGnKsNAZztLeXILTOM71F7Os2
/1tBs+NcgnEPtwYbZLT146P0P7dbRAM18+o0uS6T1qXX9tEXyoGznu7QET7XvLcbUllwigorffwc
4wLi7dANFJV1vFbBAJUe6kqw/5rmbBXFITDM45JsIYonDgLdBUW4+ECeokFwEarMroLZFCY+AcB6
EP5AbWOn5vXbPxW76/+kRHTCiJ8naQKDYFYK2ur0FsOoEJxAI/N0MzNECjXQNcThO+7SKhQKBQ/b
ZHfhZ4jREqRizr1hEfO3zY9tc+m2UxunRRKTLIYNp+2mvjY5JUwTiWhCCmxlr39o/W6QB4t6d/8t
y5dwKUXFsUT8nI41bbXUw52ubp2G6r9wry1ioHZWHWPkpwnglWDq9zqoSQfRdNS8bOiTYMDQMaIl
ls8Ufvw61aoP4cUwFFV41tZi9GEWz4eBJ1x1m5OBoojm7WZO3azUUl01s9MLxU8N/9ZtQCgV+wC5
RbYcSI7eayFN5Qyl+iSdQ+08QXfdWWwTWCvStufguc/+Ati2AT/VpOhuR+C9ol73qPhUebdBHMtV
/yIMgk7+MaqdlKAlUrUjghKu90qsz+ByKT01jCOLlcIu8VycI+n3r6cgG7TO6U1bXrlvjpmaCAae
m1yirFFeWFMnqLEa2ZYQxYspj9qYccU39BnarIznnKXDqyZl3ajRV+IOXZ6vUSKyXAk6D/WUuOOc
kWCmoHsVF9i6ZtYsV1nqwRuQ0ykZxW0SK0NHWv4D8Nw8oBsj+k2w8XVoiWiRNJEP1EKlweRfNHew
qYEfWJq0Xbn7YOPVRMm+aENZYhOD3OLa0vwIFO3f18ktvAkihywwW/axwxACPuEiEO3LYd4LeMZP
FA4/wD53ShH+Xt51EIBmEXyD3dWT8MBHdWj0qrv0CR8AWzG9f2tBALLSq1Ogn4iAbfC4D0ik5cnv
TlvJpH/PoFNA5RrF/uLoustRViTpw2Cdwi9awus814idJO987MclpNZjDngBDsFRMkD6A/cNmrtj
eJXOGKZnj6dc9WzP77XyHc97Pw0HMbEuH8WioyEda9UeYalTpusMV2awVYPRc4pYED2yZ8KWUYRS
Ph3JcTujad5qtgx4tCmp7TORe+uIdY80MPYUl/cNCYmJiNFRirP9HGVefaxuGS/CzQ4AJ+hdO7YE
5f/W11euc75CHi3A/kAqvJF/UhycfYBhrF0751fNduuTLDi/roP+zK7VFRvcUoIzgRSmQrc4Gke8
cGgCisZs6Ff04MbiWP5/3ry0qW/tJYjdEr5zIvbH2SElpfomrFAu1hd1MPlUcYdPGEyljE7gfd4H
riD2WAB9PFRsxmpGVd/PWItgL12+5A1e5mb0QotIdJqKfUhzxxz3oY/1Nitxmj3V3m3Likox0oyD
ASVrZfP0lwHHZS5qXYhAJ92iTjxd4mEeX4fIPNy3XXTYyxjB73LKO2ckdinstL3lENxtrU6hJPE2
5N0GGKmIcyrNhSCFKvwgzHiKPSrojo+JVt56weJHVYTHFhRT5uIDCpbnPFzWtkxyH/dfUPTOYIUu
PF5T0UdAqDvmx2lKie+61DDf2kU2jz6EL2WvIp7DSg6X9THwMAq59kcDxUIrBlfeCa1l4O28qsKx
cWAjaa+loO9XCyYftGTGIGLADLPqQ3Gm6708L62o2NQqK48a8c65LA2TXO9Yyj5eXaL75yT7uh6w
CsJo0sKxOQSPCjqlkXymoFvbMUdNVvEOLWQveZsF0KyY80NzoniZpv5JmNVY6/e+v3YG/PyGFyc3
zl/HcCaoKLFnS++OKi8hbG2f2jXgO49M7VSyCSSgMEEqeq6jODUqh8Ig/wQhzwvI7vTvJuYURBY5
ZPwR+TfkkV7R2nZLzuKQnzLOi0EnhvYW/Rg6RSz/uN0mXSmPxE8FfHccjwWtSvvLWKmd4XmaRUkM
mDOJ7mMV0k+jHrxa0eHWao9583p0z10V5YHTgChbanLzcHWn0mWQxVfTX/KYTGEywKoQLsc/AqmE
/FwDBKXcA7K3W0VoUiYamTHbn5jgynTzYP8FSEQZ9NsteHEE74aBn4Cxrjeb8QMAzCr1W4b7Dtg+
lut1ADanGvLKqU7XLyZb/Kr+y5dQrE2ZAgt3Fk7auXjRgWygSltug/7paawBrdaS0jxvtICZyaqy
w8xcYZkhFaF9gbWoDC5izKeyWj7CJWrzoj+44L9+z0CfnnMFYihjteJmNBWyvUwI2HiQTdxgiYv4
AzhgRmzEfLVxtU+sz/sQcYsQUYYrA53e00D7/7HgnUw30Jj3LVdgMvgtusiMg8XNZONKOlt6wQrs
g6YlBHiB5Q4HBoHaHSyw908EUuH6Cd6f/8SYCXu2J3q49imbpyeGDRuYJsG1gyAT0hX/cGKGCvDC
W/zYdFaQwpQ85fZc/f+mbOjn6l8v3JGBtcdfIRpXKO/wE367Jv9vVvYwVtBXdXApSy6moy24Z98u
CN43Pc8q79LRgqPt9qUeMFIIKPQ5VYmoCkDlRgrpPZs0GQX7nGbPNhrP5dAsCXAZFiuCUCLCd6Wv
cAxCovL7XaMMtFouwYQW2mcJ84f0gf4aA1T+23MGl1Mrxqv0OqAprEnqefrNHHWBMjGzfgmDebSU
2jVkLwjZVZ5wZE3upXPxFbhkZGHWCrHuIihu/bbho8ONIUif746p8X4NSdmgrpcgJ432ZTzp30JJ
rhYa8RqDEZ826YCFItZBV3gTHGgp66Gp6xZlqtvXw/tt9xZHYI/Hds06HXcan8jajLsufC2+HGIf
+db5RmKEiIBz+J0Lrq6N2ovMpzWnFN1SDIBj7RvfPNeC5zNkyjbm8Oo5cgiwpq7aEvCfgn1STgG2
HFRvq9hM1HCKXo2p+xCcQx1JFGLUmbN4hOM5A/VMIhmVcTsZHgIJUqvMn0li05CckW3/xgAu54rr
Vs8iRqPA0udmKPa5A0PyDQYQNannfdUAZLAT97g6c7a6YpDC57RiTT4FylfCUo38mMp7UUKmJi2B
yAp5IV/V8YxSn8SIr/Arp8co4lagX68QOkKJ7k/AtCAK4PZxW2JT5fHS8NuuQDlFZpFT0olanhRF
J4R9Xsfhn+soXJCl1c9K1Q4ieo/roamqxz0NOOD1cHlhAWlj/1mgZdEyv5M+YACiMvQ+YtgM8oJH
geRXnCNXSxkIV0I+hJ3PW3FZ1/bqg83ANqpglUME3M6zClqV8X0Q3ySP3n+MDLk7McJgeQYZHe5f
lfBfCqF4+tkOORP2yTBCC8iclOoK79mgRslb00b8iOoz36VIUS6+ZWf+xPs5ifXGA5UpSqO5SCas
q/BobuUp+0RxZZDRdjE0eyggzPEkUxRwgqi0DyeFgI0CG194HcvqmGucc0VZ0I3tIMd91Yroq2/c
41yorHFqEr5mfwNgVo4NcW3NnooPcwZtM+e3IXmKqCFXM+EEw+h9UfR4YzPaVnth+DobH1j985S1
vz/FFP8m0UL+hSGd7tqOE2Al5lQthG2lnoKdMJKGCdJuqhcV8BVXhzpbSXA+OLpUB8n4uqXe733K
0WznEQUmyaFYqcJ1ZHDi0Z3+4p/kjd9ueNGSBhFsn0ZX7GhIuydVXqLV2i7KG6nVJvbVzhVKw145
UVvs6dLDxnEKynTGb26EoujH1IsvDzIk1itxNh3Xbuyqa6JaaFy0ZFyS72wxzWaFEde5yBWqqBzA
eVwrcO7HAt2LdYnl1tyNjLLm7ceUfANkwQJ3Z5hI8X7LwR4Ce/OEJscE06sZFDu24YMRyfF4z5GB
neO6FCEZBF0fPiGWk8GLCCYFY6/jUjhPqc0IUqkNs1RU2OJziT5AxxH0A0IiB089SPFx3NPSx89J
YV45vNSPc73CbVxUUn4gS6iRQw2OgFMqTEjnsDvdAtoYQ94OE1Fvp45ryGQZzKhui+Yd81b9uWv5
xoBYtwkwfGcPCc0DYaoshUOVAJBeKht97SsBMeVNv2y9G4ji25d9vzGIZMien2wtN8wyYtE84frN
N7KsS5hoYf4Xlr5WTTnETEBxP39qNYToipJFMQvAQkxd3D8M1EYxlDkALTcvi+mBAOjipoYCdLSW
WaJ/E2XOR2Mj9q9Ctt8Xpu0rS6i+ackm68pWroxQ8iZ9FvjkwLvTLrSoGKpLthBdsw6zPqbadiDd
Kd4enY1sON+amwVOxiX22nu40grcAFz8MttPnz2BA+P6/B4jAjRfX3VOCXQIFyO3heKmNQKBEESH
x+hrhyJz64aU4bdncMlUcGwaC86dYRN1R1aI5g1skCJMh81YKxqviXp3h03nVw8xub20q7hLqjLg
+7ipDQFhK1dEHmZi4x+PUsgT4padnxTzGReP9c+YtzlQ5HPyKhfTNQX1kcCszYfp6svEH35za7nL
SKwfVj3JAiSSSWAlwrpVPnJliKo5aHDurTJMitDieG8isxrnzhLJQvgDmIFhqjlbU0XAR0lj/ShP
cKnx3YPJD+rUTMO/+YN03xhhbY/t3EZBR1KyP/rMVLuxVvzfL4keLrRR5FIlUoXpV3duV/FIc1/8
e84taroDiaOv67sgSOkLIcs2Ja3JZpMHYnKLocycT3dYYk8ZIZ9R1H/t5zaw+xdkO/mh9aoPVqvW
l4xrydv2JdpoRSNgCs1gWqJz3l5mK1fk0+Ag7f89CUvwz2cLeSbJYdEDKbiRnSnyk5DkF0o1elAX
BLnNrORAOqmd49FKSTdvy0VZ8j3w1Q9DMe4BPkzLqpMH15O5vQu954OGK+0EcF2qh4awK+BMJeKr
jRQWdAAMqFLHLM8LU+4wOYshTKIkdjszvnKjQx9X1UW7AyT93vHHA9irUaU5XkC0UKpPvyvjd/s0
R2/mykq5dtArh7V4F9veRauOvJI+dEcPYC7V6W3bFexx/EVpyHLwwZSojfczOHpMMny+USreIzgV
ZUYZdgPE4V6HUr8YNRTSUu2qe5foEeazeMjQeiUgfk/sDTUNiTamwm1o4FVBb7dlsptnMvyOvXbm
zr/w2oIg4jRHb6RyfXIVnQhXfJwlWmTJtjthPegM61CSOl4wECs+TTSA3syMBqEkHzAJYtByyL62
uMaiULh+tM9OEdO2Vx/bfQbVuFYQgAg239oIJdBim1QV8eTmYo6OYZeTMn18bqyRwHYk9vGtrRjB
xHtzyo8BT/LCWrYhMtCkqIssRalc2TZYWBo7E/rE5zjnr+Wwg2530uk3R1o0iVn4hP3e/NddHdSz
5TXPr2lgRuq6OsjCQWQTPdHAm7qFyypqveEc/8zrTEuUOG8WNFrySnaeU7cR2QryVtumQrnbDTSS
vk6qqxI5fR6DYAv/hejKTmqdHfGx9F/NkpZyQ61qG20YT9k5vR9fZTT6h9sLZsAJgPneHpDEiFJ2
dOrFIxmO6vnrq9oJnI8bE5UOp9b83SJrnSNYI/hsJ7GdBK0P3dHXpGUoxmk17BenbGkt2c4jZEpk
V3FrDzC5I7wOkoBzYD7JIgrbouXIlERdT1OQQ3NXEELRpruh9xDzzl2BWxwM38btiJv5L58uRQ2m
8I4raAlf6QiqbnnAy2UTqQVTkxi5/yGvHmHOAFtR+9FEehwj5MDF5NOFKAZ9P0Zw8285td1K7rRZ
mRcNfaC5aMAa25wYaCP5IJ92R31vR4KxFQzGeyCDqLZSAwWbikc=
`protect end_protected

