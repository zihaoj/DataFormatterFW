

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DndfBI7K3jXgN7GHRcECwyAER1W1Qh1PMsFelxk+HDT/ClV9Zo8izeECQIpMvK29OdY6SSkvB4qZ
+AYx/myMTw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CdiSOlcZSDfE8CurfVdELYArX3+TnREZq8E2Yz6CqivQQWiw5RGxv4Gl7Au5kxChzGyLzNLvpmhT
ppQfKBpf+XrJYAfKx28pTmAx8X2waXhIlI0DeX8Ov4RDfCu2fd87Q/1t9q5AVlYHTpz7Pm37oQMC
BonWIfylGOa+liG14eQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gt7F+PGAaFvQvayxMkye/PdntejydD0eqxluJporKL/eE7tO3gqhoJWrHr6EJ2JeFopjz8ez1QhZ
7fAYU5KG/SEWjH1mXWJASfakqz5iOx3/i4t+1xPIK6IS2CWsRDWrz7qcp4f25fwEKkNTRTb0kA3S
z037QRb6Gcl9T23pQbGxiebbA2gHBh4zigT1WwGjqx80nEVyADg7jOuLU2FeqX8nsBo4aya1AaGy
GqejeJaJ5IQ7EY9/zBAWE+DzyhN4Gv8mYP8lGSxa3Sth13PiRU0xsOZGac9yKFHDFVMpCjhoYAJR
tGl0wUk3TSBcSnsYqPGgP97x9w0OHGuDh5JvkA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iuUGkiCJWqD6S+Ivv2+2YU4CYQvzOyv4L6Khf5yoSOlP+8rsrITJxR/snSS95M2cb2SYmzGxjaxu
2TAok7Q+ox5BAM9XQweWOfuwovlgJjHrloEcnxbtYORZwicYwSa91IutF7z8AhDo36QmuOnZx1Z9
NZoQDVYrfJs8Kz0Yenw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
a8x2Lj9mmpL4v+zPKabbpGXEXECaXjvwa8IWoZyGK6gZzcKlusapcFQp2jYobjGuXoqhkYYp4ANR
/7TGF2cuIszd4V+i1ZZL4M5UXTQh9kLT8emsG5cwnR+Nehucye0a/SdOcbn6Pcg7yMce/+zpuuV0
ex4jlZMAsXf6i1il2ddPdtWT3k2AbR+Am3/f8ushp2fsmcGMgRVNtOOYROsCDX4KlRdas9YXlkq5
9d+ubkYzakIVQa0PQ0jQJQPW2/C1fKNsLisKy4kJNaDNwiXo2Ve5N6Qxb5irFP8wZ6iapscbnarw
DNy84LnVZiSVsU3OP8/S7YHAsdW5lukpeuJb8g==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oHWnYLE0J5rZZEnXMuTAQxu9NgUolVXZM5hq9TvCFq0x5b12/jzoW51moxTIzUBj2smQ/sB1QlS7
m2fDrJuFXKoj/HCk0KONHoXlaXmLeXQqL6HYfKw/j2F2fFIBmmAhAJ5qyyPkPnlXCvkE7fsc67s3
qz8a+KKsHGqGWBdeF3lAT6y/10HKSeR6oGugaujjA2CDnjVv5Me6lAzz5C8lRfbolqR+3RNm4o5P
Ra7RJtGQz1ANkLxMLrxpjcw7kXNTLrC08BCVAukRWzPhr9a9wfHitoK0WlXx9s/o5jOgg3Z6WSqF
sJxU74LBWwstEEO17Re4mT3AJPySE6IUwgXMTw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 961680)
`protect data_block
m/K66vQYu9QA1BLl/gcAAFfMcny+9uNb+4fAhl4D0gOczOxS35KAJpMLCe9W5beGdDVT6/Bme1U9
1QTAVziLvfG073VdceUFW7v4x62FN98GsFAOYb3NQBws5PJlHOxrqytAvHLjefs5dDwnYJ0m1M0z
jYVlWa6w8OaSSogKZjp38wg5tCstVJXpGYCnQuws5TpG4XlycavHFtWQt/sbHUZmdU1KIZuvWAyV
HuBQLjr7lFTd+daVetVsViWJ4HEUcnvHfgFys27TQtqBeL4XitfT6IP7vK4yE1yw6RuO0NFRq02c
5hkruW1O8pc/kGFvnqvbpGtIRay+/HWQYi8AYyEK6o6a/kLQzByZcjjeY6KsHwSkLFf8d9OaRehp
zN2SvqXqPVFClcGl8sYgQalaZu8ecBeHcAHokHET1R3JR1omlBrzkK+QmOLsrH7ZWYjRzYDn/Om2
/B00X4hJR/YG0K3kE2DGxyMHgaR4LD8gYqep+TxepGW/nccU/+FRshxMYQJ8FQh4+A4oJdKxRtev
BT4/fcwszOl7luSNqfBArRPvL/vyHmuVREysJdurE+6F1uowqaLi1QS5a1uvliP3OE5ONe1FsO8V
bsLJnCcsv0JjJPtM2qvLAFtosYPrQRzKtWVXBT1YxuXDwi+HqRGgMF6oq0fqVU68lKhprYRS70rC
xeosXQx5709DKO8HIxJjt2m16VAI+OP0csVyX8oTBpdgUnx7CtbHB8I2BZPhM5qd5SGjdsP4XkIJ
u+QCa+jqKui4wcmaD8sSSC8AuaVT/e92IiSFIwx7GYIRD9GK2dzW9cQIeIkMUZlV6LFe0aaWAg6V
YLsjJbWTVRQSlbB3LJB5nqsigRWPS/Thddenecf7MY9dxsFYMqimuyd+FOuO7oMKKVkm+lFMSZhB
wGw8gQ8/+j5J1e9aEyOfmabZKuzuF+VbBKTGvLtJq+e1ZEyyJZYiZ6dGhezgn4A6eYyVLsEGQp0J
xeMXIiXXDC1r5yo3c1o3Mul6K5qMNyP+q6Os84JvleBAUyi+TTgXX6OSNuLBK+s9olAB/BnXJz1c
M0101JpIU/K5y3YBSifSp90jyphnz77XkpoLgXV8utq8RPyELM/AptZt2/UMu0YyHgU3P1/6uiPA
zvXRzkoX71DB4BvrgIXVVqw/KfWT0VTp000T0yMfgznPh6+9BIl9YugN8gBYO9za4hvD015iR480
7IjW8zhS4Rx0bvqu38dqoLpIi9MskGZuW3qsI+W4bJTR8h/mLLeJeImT+Dg52mpF/TAqmAohO1Ye
lp2PghmGkQteaW6d5UeEuP7WskPTDDaYbDZh+ZpFe2U2zmabYnBLk9+g2q7dxcTXLIJJ1yG867gs
HXFF4BoMLXR2+hD9T3y22JS/9+3+B6FnuP7FkfVvLMz9ppC2DzGow1v19FHxxcd8YKUmnDdoyQOa
gu7dfr5bFHmSUBUVHEdFBh5HPNq2KfHrfLmEABI8ldTDHUCoShwuFd/5Egq7NItYdQIUc4OzPcAl
NGrxj9q5k+G55gsISqkAcG/UYz9cnjROwxme5CgzcrRWzMJikRXoaHkYpZPhaAsg+CCKnYRksMGU
VSzOP+d4G/Z+0y5fKEHfDnHJyhKeYaOinEMY0YfCXAdAWxUf5/bgAr1uO0HnCDktlc4MfhrjAe74
0oi4xN7COyrZQr1qCMQWWSgAZw/FDc8fq6k0HU9LkvZJoU3v/Cgtc+gcX9YRWfheLArTOSqV8xiu
Q4WHmVcnvTkRQCAlplXHrvNQLDPZTaIcai1lOglSvQeeMqa7NjhFZDmEi3YXGHwWDdA3ML4ZnAXD
YJUkGRNbWcjByQoN1v742NUWeax9ZR+rGLA1TM6kjUKMATA0ThX4A0WtpGaC8HrLXc6NlSb1GPaq
brzg6er6kHWtJRu7bgJB4UsucYGqCyJKRjBbDlykUy8iNLcgPYw/ddms5TkfOnlVoJDtysbNDxYj
PyA74c2wUa0Wx8bqjCK/4MzTCOOGsI4J6MWyq7TgEDsZTZjH6F4JjiAB3vOUeQ0VJGlPfSdZVprC
Rxig867BVqO83DCYHat0oO59yFFQrbLDyYTJTAO0d3BgqOyx3K0QZfQ053GUw45+A1/WYvHprTL1
m4BynhUWQ+vxwuh98iRYKHXOy8lO3l8VURbjRjAYy0ToXmM9EDOkIXtRoWs5MYmeh5J9qo7Pqvcd
cOi/oo4N+rG3v68fG1FavTcH9U292ng0xcyNH2OIdJ4bJkY/wNoatgz9siohI+2/g4wgUMh/dU+Y
BflvfiQr/mMHHcPSFQQ+2Cs29FGqNSWyGBDrlX93YhujhFtXRPTQq4oIplX3PldyW3rHd8DMjwXU
AspyRdAQWjJoHXkqursUSVqv5RFBYAfrV+UrphVurkah6uEst+s9Q72TN6m80My45VTmAufpEFKT
Gy1/7MlCP/7uc4UGqz1cpq6pcfkUpGVdncjKZvW44RZ9dMKW85mh7Fa9bLz0+ElWNJcRcrELXxxD
1UNiMSZPz5AYy3ui4DQdMl29H3UV7ldB2W2w2N2ansTutEB4BXCmQIOO/8EX5zb5dCMG0yxkEdlG
pa6WHu9Id0/y4KAf2hqikOcnMeSkH2sDCfE2Z3Uma6YHI2dRWKFrj45PyQfuEx0lhDs2nSOl4ZGY
yur3IETiFFTCrjjyLpJXczOGvpuNUbMrbYbmehTCFZTIwtmMqXaVJTzM6wabrwRO8Yig4rOLxdKV
cV9feQ80LvGBlTcjUHqd+4MG3CaEcj81VMqRj8Xe5P21pRLAdn5Nj8198mpFs3H6p6VGYFHEq1nC
YkVvZtCk7bPayZIfi0evF0vzbSWYNZi0lCnjW8JmHRRbYSvzPQtaIm7c2sSlh2Ny8mrN1sqH1E8+
0hbnsnGhX7ytpHVVKLMnNO8My6ghYpeFpSLFQT0ktWUZV85mi8gVMiyFqc8coT7nl1xq6CyVHcb5
ttGtmNICZsRme0gv+x9J/lGInjxlc7NKaxWi9KHNtvJ2UO7Ho2KQ9rVlgzsM4cl+Pe9ox2fVSMab
nI20HpCp/jv/6v0vkoIP3lV9r4WJBCNYk1sCZY8KTyfOYwOFIJ5cT4A8ocVDY8gngPGckShkgl1s
0IYD+N7N+mIN2a3fLO/wjsI3a00OR5n/WMZH3CNE2+3kGWE891geESk2Ml6v3V1VZteKi5BzgFwv
vVA0VgBP1euwd3pjT7Pg29F9KYM1gCSsKSXyqHRLjkfY7gMLpnqoo10xSP5z7DKp+YTWalKz21Rb
tpbISra213xbp/qHup3O/Bj6DnAR+JFOcRdcdSi+NBmQYN3dKgULlt5QFWEWiytjtXnsiH6TkeVe
zEIfXuIAXeSGOmGrzOZm0d8+D+kmceo59OVCsFAwufuX6o9/Ad7JU3EExQYQ/fsIB3Ev/xW6ddQa
lYHP0Y+5MDMFjjzJoXjK6VZR49lqq8OzZLRIl/njaQHjN12rllBWF4WrVHNTYCivMEDHsLokkp55
xDqvSkggkkQykd/puO/QuWImUJ10nZIlLupEPwWMXMZzDRcRviOR7WITKf3on9Vr4x6dYFJbhvNx
/1uZdYOA514GVZ2xMfsiGxVZN7q8dyjoiMfCoB9z/dlVAZZLI2UtuyS8qdlxHFr2GD9fQk4Q+Xwa
E2tygc8OMWwx1+y+Z8VdU+WsGP/r0jgW35nedwv+uuPyscGh0vjM1h8GeKnSCc+rFV142KVMLMzl
AWEd1+GePU/czbT6o39er7/KgNDfOj3U8fnhH30WBArzt5QhHTmXgxotKF478waNmzxDl0Luxgj4
Pe6co+MldYPYh09MlqDuJ9E7kd8MCjUauE/9vDs7R1/I1wdi0HuCHVD//6aHFBKzsQOsxwT761zc
rI6wlsBBpl6cQ0y8iO57KacWbXGrnbrk2TojlgEuccEREHvfB3abMaOR2+5RVo+i9+pyXw6TWMuS
b8oISgPOqgtnTglGmgjnuX8dLSJ0Bc9fx/EmPr7piM6KL8XRgN5pp6h3FowGtIDsehjjDwF0Z2t6
n4yGXrzIadzpX1FFOdlzDeyTDlaoSkEEAZx9Vf4gko/NqBNCj3bt1uTiU80PqzFjDbXFstnpgkEe
tSOsFuIO0qx/4mGrkW4Ib46ZYbehScHhw5oWcCyRR+Mw2J/jFD2INMVnDTm0Q1Oe2xK6n7Accrbm
2/KlwMAUKFVnH32YPcfwz4vTlSo+pFSc2D5tQB//f56SUGHzSGmz3KCmSF8YvPadnB9vijl0wwka
q+pOd3ByjK3/57INQrrE0xhDg6y+xvR+GyUk11azAL3mOqCAndYaUN983H7clndDxir/wevUxYTx
yYTU+I7Vng+2zKH1oko4Fp/8+E6i82HliGy1/Hgv0crzU8jX+uYWCQt/YrdaSHfzY5HgFAIipvS1
VznqS1iUfN5Y4oGoxstBCkFzIuHniuT3J0uS0ENWePJTA7pNNppu26ozES1G41HBZVKEWC939J75
TdiPoArtCGSmbH08HsI8ZDtOBPzPtXG2y5EdPyEKy1C3BQ7DrZyZXV71cOiC/al4w0d6C5FNmfDL
J8jiAulwXPZBmnSA+BWS+falX0Uh5LrKRxg91mWvTBVFq+4cMUxkkHmMmXhC33zhQsx2vwKdzvIK
vDoNEy2Pndatvnzp1vzAXCkofTkgIjv9QZ/BOn5tA99gSE2nwz2Hx1nO0UsGDywgwBgpgq6JnpJS
s/qm+WejnhzNE/6qD39O/Stu/TTAl3ABFhTxq5uPmYCmFMAMrLbSbl+HSG4xbm/e8keCvZgprJ4/
NZUIbVITvisMRzv0X/1Vix7F6okm0fJGBYdTOwmXrby8f1dfoJ+MnqpXENNh1fsm6EmPS+wBF2hX
pIkV/0eA5dJfue1PBJoTj+ppXxXeea0fweqwkqrd98MQ75qg8p/RiT+duTzjub+N8sljGCnDyhjt
pc8b+On+qYR7d6xAb0jfFApOHnrsl76GgZ4fx0tcTsWIu7vaxVhDwSvP8TsMlWRm1UET6FnuG14s
HdCwQTa572Nu/8UXlHT1exSqx5KvmZONf7zGLw0KrsN90dT7kPmPOGCtaObVgQE1Tfxy7f1Wy8V6
xlJFN8fh/rOgNhnzk8PeotUHtgZ0sjC36ZE+YNWb+L0p7CdLFR3CpUYDK1b6umflboEuSXRF8NoG
ckm5GeyOTlWQDoGSu17HOyi8R9iPBDLLjnnRff+mGHHrb7bjmTwtD2/Y9GYGo7f5TdouuUDz/Buw
PEycftzc5romG4hGb1Z6gKXyWewEAMP4YTMGQ9++MKNWHDlBDYwdS6OPcQVHMYukD7IEv0Lu7bjh
K0HhosEq0LKXPKZyqCS40bVHsDsKpz1LlR/r0iNhT82t074Uqx7mUYLpzj4NRXD0r9gzAuD+S1xp
gHwX3HyubZUNV3mSuEDF89UiySSo22wmpyaFhmpOsChEj4vyIWcDbRtg63VyNhYJ73clHV/iDc+X
OrVORg+xJ/dvDjYV4twheaT55sOyrvS42qeqM3T669sHcJtuQkrxDHzi783ESCtmuJHYZ0F7zkUg
GM0epo0vIzznGadGsOl6ZnGyV1M90TRXaVedW/m+2u8vDlMZtkVJTyFRtnSOJR+hnJQOHivsIhsx
VfFi2ikOQtj2ad5ZcOdacFLnulHk+H23ufNAMs4jPSJ7IP/LKZHKm6llYmiZv8mnBqSsB58pMJc+
BSoxR8kOF1N+b9vcAgAtYAKYU1FOlV81Ez7UGawVqmsl0UYPapp3eNEnEcaQp6et0hNkk9CpKkbw
SDSUW18VVPRy/aR79wHXOILPOrWiR/XcdpCmBRfzZVzFbbv2KIFRqUQUfuywOMxBm5L6CUh/OMVn
Zx8pdt+xYSsGIFC0FFz7rAtz8v8tYteddaSwXq7OeyztuY29IZIVeoCwtzrgOZ5Vr2f3QIjoDzVY
n0tOvS0rmnS4j77R8rX/ZjdXdah/KjqRGaB+PVCL/VVbJwx8Cf2QMCwFa9va6ugonuC0xrZfpWeX
dtSIFV3QxeFvh2nyr9qbayNPDnypDzTaI90bgM3SIbwSI6YP3NPYwOZmxWwprmFeN8f3BrJtMJ8N
mpOVL3005rx0EDrfWd0IhbRgNACxOF2aIZkM/LHA5hpX0qiskOkxWyZLTLt93Vzx8b86w2rpgpGB
SOwXq1K3v+YcVkdyU3c28L1itz0vRRoSGxaIAzA/vaXWw24g7gqMXyNAbB7pyoM4nB7ybmpsgiOE
c6i0yX0/gsDh/DG15XEVSPGU67ZH6z0EuZYhgU6QTtYp7MVnmFJ4+bSQYu29KcpMOsn8DU0INgCB
yGfYVrkN95ofo0MLbThaV/2klojSyEjYdXSnJ8e+d+traJyTYjpTlvmBkH+Jxda7pf6ZQWNCBKVp
29mb6QCIko0VvqlsHXtUbz5gkAzYxISIU1Pt1atNlVRhe+KSfCPZeefE8Rgm6XYGkmhNRVkQ7QmR
8b/9ONHTpyJdVMfiJax2OecD1zetT49qADv26X1z3beZ93Fvz49eX72tw7ySUQhC0MenZz8vN8KY
O7UMohmR2wv6s92PG6GPgIxqrkJxBjS4DQ97tZgv+qv2rLM0v50LsKOplL7OaNMHuLbGyc7MKojH
TLaybSBF7l6hHPsL93wzDD7QvMM09J79PzZhZPukZwZ+e6ElNvhdabND8wqEVCqKAcXNPdWjpjq6
YH+8L3VZFWVBlt48kVuwCARRIsqZmkj6CNlJiyTuCNryG6ZuXUvmVVMpevymGrGRmtFfhv3nD1iS
EF0K2qkK6174Ky+ppsORGZpzhYYC7XomH0N+lBsm5jc4leyz77a203mQFmW2cLCz7n3GflV2ikVV
lKfpK/rpCOeJWXAcWhyqw801jZi/xcHtAFzQhYApSKyGdwH7Gcyf2Lb9AtQjsx+N6w6iMaS4+fZ3
+ZA5gxehjAqZWNmB3z+805fzhk4G8g9V1ctYNRpBxwzFOsKERIzbhu9PNPR2mIp6S3pf5RuEMpDa
svwnp5K1N6q1DhF3eYkJ6sXgvNrHw5mEKZJHAogzJO5eHZ3o9vagwAljOXBqt7zQvDZVRt76SWS9
YDSOGEX4tW888NfQmnU6ctrx9MXJ94h7NXfv1UYBI4VQVnJ8t0MpnWMSQ8k7UEhBWHGOHbeIw3B5
Tj9Im38VxUNs3UXLSdvfFPU/jxS9cK5Cohofm7LRSGozfSE3Gnk8eFJ0VR4ziOaljAqpwZgFJL8k
IPRzx97d6jed/REMgig7xDkj1LqvTp3JpXkyqvtY2bP0CB9OP9U+YaYGGCxOYHEYErMFar0WMTVa
5UWhQ1FM0W0KLmaUQsEmKKOrJwEpGLUtOciszJrjBAM1VwwvSuZPQRV5K7YsMZKQ8VbCjMe/EJha
buNFWPoVi/FmrhJoQgocu1TctYfnZMtx+S/HGlkqnz1f9BTaTpnxKvJx0oAIZL/Am3ir+vzE0edT
kvCJJ4AKH0bS03DHOy43EBUhF/kPo0CgYGnlx5IVgTmyMjJnTIUd7jTgj0j46mWI9FUBH0nQF+5k
C0pWf0VqEXWO7IZ1LUuM1AxuXegzD6uSMg8Ep+NzANnXgl685C9Qg9XUb7QCkBDrId0IsGcD/S+r
JHC74iwUucg8CRUvnYJwIZ+15Ebk707ljhoN8qaUnLfXqHtyjCmJbcSe6KkRnDn7X5GPvMgWsOVh
jn5GCdChScqYHvEtrbGkofmdsuI7TwBDDoi/5o+MZWE9Tuc/tgdhf6+UPVyWEGWi9G7Xgda/B5Oe
7kKPFL564EFIpFhxUzrcPiogA9d7j2VEky6CWQSE5JEBRnTR0Erozb8O4X82/g2IIj1Ej7eApqZ9
fbGeRBolVOt6C1NGUCcJHXYb63qwmDTEieeHWyM+NwZT8qamdDmMQQwkFI4DolqiD2MML+j+Y2/U
oR5KfDCIZQrXVV7sa+MHhveOMoePBjYa5ekzyaVlAgx4pkTUYyDu5rCPl1is/b2z8jBatuk8IPVP
399S4j3hj6vJ6ffiDVAa5vWVw6VIljIcigfHAyTkXb4tMsClhRAwwobgYn0JlB+cBe+zkdrKxLEs
WGp5tuOQFmzY2X3TrbUz9XsrGCbc9qRxFgbEDtt/bHLspowYVY2IJg+aaO034Xlifg+SY0Cf3uQo
+Y4qDNdBXqhXgxAsYnOn9UF0bFM+yqQ6zD/gLBSQdvMryDoIfBpXzY2hJMraDrRbPirJZKsCpr6Z
WbTI1TrVX9sIpNSRyno0oLwNutq+9QNv9pvrMc4unpBSJdaW4ePTxWMC7wMiRZVMIM2z9z99U3M9
giABG2+TawOTNyo/2E24eV4zORjLXMtckieElXxKoKgpRBh025099uPFvIFkOjNyArh9gS7ffo2Y
KqmeBj3wayQDGCLjZ2dEGM8hY0iCeGIN8eOxK+MVFznkwegOU39JJKQOSxqFjkwouumVyDIDmnCq
HW75sBFYWycwV05c+HOcMZBSqTb/Nw6gLxmxOY8Ha4cBt6BR/BSNe6d5W7v8YGB9BWS8VD6jPqR+
Y/JZxVkl0ypMyE9dApcVWz+ymbk8Ru+TmKBPMzJx5mQBGORaOwHK02QPlS9Z/Blc6f1XVJOf26AG
YPIHKT2UNv7TPvwx8LDQtWyFXM/kwWFzvtlCieUS/rZXluw2D+42VN6sqGPa2v51H0YX92RKahzy
tx65h2dWA06qPlwghdGkTfarKzAi2ejsKgKdSqeanlj3dTgOkepk0m/+hhcWidqTLIXeuNFpW/KO
uqcGhjvxWLdJMY+9Nv5n1m+MtlcrR5QjqnvKzTBAZezlflqfqrtTRexspUdmcg0SQ6rOK6aXwfSD
DGPqRaC2sOucCHjNTe0ePtqocpoBliSZciSs7mh++2X5ylCsfDVf0Jj51fhRlPXlfUqV962uFY9S
zh1gJn8Y8Z36Yd+AOZnLVfzsk/Ty5wE5fpCjwyYCOsUf+tjFVDNRHGAcxGu3AXX65mfLvzB+pb45
t/7/qoglzoBmaq9/jALNtjelftRMK0KW9fHfwpDdnJD5TjNiQVpLQTP/PUFWi6eo2busYJC1lHm+
dZt0nqbw/nBZX1vvaqPHTBbs7Ib4GtJZRLpCBH5ouRoZrjFv8QRn05CpmRhNzTRir6nK8GFQw40U
3Eo7QHbRvX03r1cBxPGGNl4kKig4SmpjZ5NpcfCQuvmSaqS54mLjbQqkILzoNfd1qkRL2uz9d5J3
XpWU2AjMeLGqgAk70a/2iMPuSSF35iWIXFYV1kCoKlrggz19TDI2BVfWo70QW2eQ7VIQqtJjp30W
tKka1xDTr2HZYq7EBD9l4lFGEsOGO2vzAet953a1EaG5uWDZocNoOZ5G/zr9FxDnSmJl8KLZFR+Q
ZkFphACG0tgOd8vs/mVLOjagh4r+PJMdBxouWAJgKEi5/LMOGxfuoUciG+6L0FKSqNkr48VKpkjG
OJ65svN3G6X4UaeIVetLbDqARlLcDxoztJH5WLMyz3BA22t0Ry1h3dB2e+9aZ7cizOimXlyOdYlx
tMxkx6do5NdWlw+7yB0Lju2idow0V9K6cxRsz5juHQCpYhWyx8Ic0q5g2SZJXq7MAkFl5I8Exz/8
Bpb9BIDQ864224wN6QIwjcM1Ocf7aSjPZSw8M1nHQjM9zUuXeEWVeX2DmEfE8EGX0uGgWm4q/W1x
4suwQ2bELLhS+RLJ49QAnwkkCSmsZN974Hauw0qYg/lpTWQdTzzmd82Tk2yeITumLGcObs7EiYx9
07trNs1LtSQUVOb+1Hzc1j1HTDtWzyQ9RirtN2sJjOBzxtYPoI75md7Kb+dw8JqW4Eb6OdDgX51X
PoxHOKg8hFl47panDbzS6w8UMmj3e6LTjo+R0Ij+UAFysfDEeSyoDg8lYONX6zRI/gSJ3m/IqhTT
RlHC435y2eQXwuOM9XTyqgVfYt0TOSSJ5MzCPEEOg6tQBOtlGjqjy4DvZPg+LZ32McQ8+9RDZ691
zbGy9uFgkQlXqshR75seXfcMl/+HFcbfH3FpTnbPC74UHvIMN1aJFNRvqKBdy3z4yIArpj87ln0y
4pswglBGDtc+i6l46BE/o7k5rS7K8qr+yf15Gh64cV4p2p2KsQxXMfZConFbv7V8ogy4OS7QEUqM
RZMpnPuZjDQiM5K88j28SFmczheN/6AWEnU69gYt3vIOxhg5w1bS1K6noMpjHufbUNWpQIUPQio5
EBJaJgfh86yDJEoj8iYGWO2NV/4EpdHoDKUGUWvdqTHapJ2SdfReBAspxDzx6zAj1FigAZmAx+Ao
ncnrNMaXqXzl+0IeCkq9EcxkBPIXjFs+puGzCed4+Hxhjn5N6hx/TPk8TaekmNI10LKohL+WWQs/
goYBhUPiU80q/j0UoQlSMz1iRYzVaz41V6dRAtDUtN7E03SB0H4Gaeb6KyFpNIvHVZIgY2sH1ewm
Zrdpm+0H4iZR91yGlVLArGBXjBtyYWlUSTwWi4Qiw26rBu5yvwI8ff58cxzHoNL3lM9gORcHro29
W11/ZmEz0OXGmO/0/BQ40Dz8bZz/uDIltVTcK8JJG9dgKqxQRWUYsLxSpwa8In7qeRq1Ehem+r8s
wX0k0qrI4+6t2WZfUZjVOXv8WgTBzFaOPFb1cyP73/4k5gAs9nde10WG6aoynQ6eTkFt/wgi8ArE
e8jlub79wryfLh3r1bYl54pL3JxkmFe+D4KD7D3DrVZ6gIlkbh04sTkVpS5VtdGp47UJkI2cbkuZ
+141FPX53uf0AImib+jj7Nkz+sI55qEN5nbDzymIqDnLPtXG5MmgBclm7ESDBwezOFSt7ragbUDZ
QxeZuUqnEAYL9VcWx2ww5oOT+IIRwp3IINgKTuuVONQh7RQAfaaurRO/AE+MYcG7WmEiaUyNOIFs
XjyXsxNpQHiQosYbilHqMV6wdfRCXSE3eb+XMIoP9bvGcRhwTxZkNa/ex/1omb8/ZEBsWKQ3IIJx
V4YZ9NuTHO1PpPXBY1DCPK66+d6k3MK/l7xnU8JWmTNwk+JJUAQjLiN4JdDQbPl7TegCqasCrorS
dkntmkIDKTO3i0YmCAPqUYjp5I6hTaVUhDhLB4BZLM/YUZtp1YdNYEQTUR18TFNP9HsC68WidP7h
Cu2/zdFhZCBe5LnISD0QPV7igWwjHwl9G1uPGJpgkt3lglQeEDO5J8YwyFWVgOTF6ervzBDT7C9h
fWlM5QQeJed3rHQPuE7WWnGAQDl7F6sqAnsQTb43e6L1cw9WKObuw3urdVzMN9UsigWUos3anKfC
JxbydlcrD+2q+MVgdj1tHB1PPAlKSXMLmnE5mBxxnatDyVy9ZZl0lI1h7d84uSmiiMIlv/TPW4YB
GNw5tIB6gF4gObStFodLsgpE53BGtvSaZcOw83RyvA8fLtXYJVVpVMGjVk0oeqgWGE9/iYczDzwY
s3rdPdYsB7pibc4uA8mP699iEi/TNxyHR3WO2IKHCPmBEk5PUc+5AVbxVe8LuESAIpozHyuQd7bG
xLFx297DLNK1OXwoSPGIKJ8/SDAqzaXrAUMKbgRi7lgjo9ySM+5FZzF6PeIlatuKN9+gnj48Wws/
DqcYzwR1ZIUzEMQGFVYeRcy4vlTdImJYje9TDh5+E/CNWznI1PJyb3LS9uJyKXjnBTBrxiw33ufz
ND5ZST8JveLD1t3k3wzCHoUtWL0RlvMlD6wflCmvpBbcV6KO3h6smA9GnlNKMTB8wFXTWeZ6u8T8
vWsKcbRsZv6d6UrWIr7tC6r0XBeemFOR+08MNjpiGngBq5xlAkBBX4ahkzZUsLMYCqbq1OpJ4E4x
Ea9eAFyOhlSL0Vy21ljbEp6ZhvrzCUU06e/HVKUCEsg+VaLEgBbsmyYMBykBV8TFjHLJWTzp5Oqm
BnVy+dQSY4JadmIQcR4FDV+rediP/9i0Ia+KCV9SeLBny+SJaZgXqig8rLF0OGXN90QY51ADzOZV
fzy3/DdZnQ24QA8F2M82mjNMKmm/+U02wljczSYWNJut/HN/d8BJ3eUI9QT98k6viEYHV5nERKQ+
QJHXvpciR9aqpqlidlKZ77hWAv3R/tf0d0qTbsb99VtRfJ+0l48DpYsEsDfTAQfo3aBkj2al6Hlw
Vz9l6k4mWhajQSvwgrgUOcXVJ7aV8DKfqCFEHyQK37M4cxm4E9FwEzOKkKmUQajPebtYMocEiV3M
/yxs+6Ke9oUd6Bz9SVmcQwVf1dNzm7U868bgi7d/MJdm4CstEDsLrjK6YyBCoDM6Yhi8WevuXL5v
4E3rlf25am4hGuKSFsBqahYM0EKr1Sn7ZtW9D8D1R6geX5WS3UUEOL29ChwhfnWObJshDP7qHOiX
VdihQ9WsSlFLwRzpf37KIKUhOZPxEVGaW2ySHD3IIDaLzv5ux0wFyWYugyXuiUkGma3UaYRHBcJh
2VphU+WdmFZlGrTSaQOMZV3n6tD/YCHXzyjK8Id6Tf1OK7XMfPJk4T/XuV2nKguTC4j/HqlovYTG
iQxZYEOSStEOp99k2tO5vGVbW7WqSNN3JOErxSm09Y9dGQyvdlmG4HXetLMMm/Avmv+kwazSfduI
XoIvDRBWklDQ3JaQAbJpjUaKIsc/i9WQXJC91eUEByQyqFMEyfm/iePgJrutV8vCdNyxs/HatciF
UhPbsxKBVqAztez4vjkg4DDBsVOfbZzmnJC1gUBM8qreFF+Sy+wkI4ZrMAyZRuK4I+UNlpcqJtaN
tu00CRwcCcHz05EB++GWaF9o7A3vGlJtrVlv7vLJFEB5E48SHuwNNW8vMLLduQyShhbr5DJQBmVc
xPEfnXwSp9V7LrZDp2OjeX0VjNfarQjLCB8X4NdznTfKJ8lGMrfWSKeu9BaPIck95xTXqNA0hl7w
F+ZOtX/TcOPvuPLjkBsxTyA++tYcdfjzWvSiODsW0WLWQK68GFtKtLq0mJYjq6oel0Sf9uWXR81Y
/iB3zfMwaQ88S69Pc67IhSPVt9VAPEPVDfMyQHJFhis9sq5hmM5Yw//Ams5JkyKEW/rPU++YHwpj
WxuUmrCdyFdu3R8Srq1EMLp+oXf02pW3hhKjf6MMlhMpqL2gBJf1wfRcIT/WOTVIk0c64daiNe0u
7UDUEThUkWgrxF2scmy41Kn3gcoXOIltZ0M9XmQdo/AllxbydTZvtGsGXyr1SKnjqerVch/3Kj1E
gs6MBYDREjkKmlql/8AWf6Vzy3FuLybENQU2kY81IY7DCkOrTQsL7NO4J4ngLdnVjwB2pYXI2XEP
3+03MghSUv9SniTTxVSpZqPUrQemHIF1QAgy7X7EJUJFYBHvxMWqtx6hYADQkvQb8kE0JlXopiww
z7W3nVTpuwJE5aUNNYE3VBBkn9tbpDbx2V12myzZ/zCETDZmW660/7dYWWJxmer7CI/J98T66vs5
icBAFU6/zTNQQmLCczBaMF4FIBZ3+Zn/aIlnEEnzsO3gnEgdnjdgoAv3RK2LllkfUo7DMzOl6S38
FLd74phUI/Knl9DA22AC0+qxza8De3NSjLxHjTouAL8MjHrPdGsrQ+ohHZYoMSMbbchX9VaBLU6t
hFew+llLjc5RYadrrVt3g9ot3a23dBdgtFHF72KU32ZOZVq3CaMkNwSiaApGpoK/sii9W8TR5wQd
KzITJMbNFQLevPJ9hUdLMazKtDfMGM805OKB0WzZ2iZ+OrcM629W02YxcgTQdAdwRkQNfEE9Lqak
CCGsE9OHp+1PljcQDkOaLHCZrvIsXflSAmS0axPqKyzSli7bKsimDTXU/ptqjD7FlV6eDCCBS7py
Afk7bDKWNOYP0D/c3laGbD+2zH+gJqTjDTC5DY1ijJU+Y7Uck+XXRxO311GhWLOfLqlCu5banzUK
zSQKXCdV2Txrr23IDAK1DdwBplkd335pmvmjsrS013uHLQRSv7fiJOshMrWIXZT0zu14sbT2Bobn
09scoOGGe+dew2Ks7ULRvqFwpSx+9uOCpc7heqBUYubfYTD1kQ5Br8m6KqmiThBwxzjjQUIg5tbY
BXuqFMgzovmGFHzz8fduoM0eAIeIAE7CiE6FCd2o4CAuJwqOIA4B+qVXcl31j+XNWdVX8AwkPcvr
FdeaeEzmLDmEjIBOBIiQVEelGBym2z3GONCruptvxjKlRK3sgyzVtFjvDxew5q+98ec0izC1MsCs
D8UrPGb/zR1mODOUqjH92bWfs5vasQpzams5IeKgVROjHKmd/EJ2jh1VpWYiT5z5UK/5mWG4/jc6
W1hSuE9HmLiVBwzHULGGeIWPzxmkCjf/QOfw6EIJuirlKBMCan/1t0TYKLlO+URBmbwozzmeFpLz
60XaNFSHqB8U9MS4U5RjjaKUo3OwCqBXi0hHwF9/v7EK1otNmY+rnU7aCz5D4T00OiU507/ZQrQX
EE1vhU3oeKhihRDyaBvf1TonzZwx8tZXJ0ua8R+M44WIqM2vRmMgZdXWO02QYvN+/DIRbu/zHjue
lS6BvLllLL5ESsWexrN8QX4pjCVXTsGdU9RscFtBP3qcJZBlHZHhw+ByhWJE474wIvTX3UU3ND0R
rDRTVbb8ExdB+KAwiuYdRZXz2zKLYIXqYWfBBgmr8KkM1b6Ug4X+YOR3UF9ux+TF4nTSTzplqHj9
cVhOlvLSjQqIuX4wvjPSE5EljjZpub5dCZWizqTY2RvsS7uxbcx1Nr/UA/dxeiC0DPK/5ypy5faY
O/OQPDz5tCsF3KzhwHIQkoMHtXbwqAseL62mXN73DWMCpWLVIaL/dfkTWGjIhGKf8TKp+mMIBQcw
YBU/df0rFudDzHA+3jl5GSNnQ5kmVTk+si7WzFz+ZIwQ5qnNIMAhIvzPLvDAhs5vuqI+4hfkdXaH
j2yaC1wCJhF+xVgNH98HNiCtcv4jW2ppL+fTSw3nS2rx7OdHSb0A7QHuo6LTCxPyzFg79XsKyVo7
vEt23A7/6RW44EomYWwxu4HqDIYfmgJyrKN2p+RtZo+H6VTkPZ5EduSo5R8biT9xc8/sAZquL9Ce
Sg16v+j6be1P+yFbO51CGhSN6V5n+LlNNWUCbeAeo2usp52yaUPRh/0ZYa28WmU/bumLu/Im36kS
wWb2UX+ZvWU0BlRzhn4yd5ST5IMDBHshxLDXcib5sTMyQDJT2wjT5F0HuM/C1mLK+WLnYH+f4bze
4JZq4TGASVuCE5Es5DC9grbb9sEy/eIqCzgYPD4rtn7ZF2wsIYoDYbSUO9yc+v5TE9oX0gWLhfR5
jfAIJlaZ3SGI1Ie5OPK+gjGtUTqRWYnachh7/VMUlIFsLdGF/177wWGrxMUsxYiBm1sbHoGvLUcd
G18GJnN5vp61JRIoTjGAT+CjSZGaS5G+Iq+KGu521tNSV3DfUXWl/IzilXcVHGqhoKf7cXPOjQ8E
Ml71xGKHeoYaJesmLzRnrX7/yLNr576vFN1N8yqewYy0JZzxHvFIi7SfvVKoOqu/ojPGQEdaIhjc
QmGhPbjjYBxa/NdZYAw/GWrGNIJ9zCUSWxIK8abAElW1db0hzcLQJw58+vNhqTZlHzhzfcHizmUv
YiuXB7q+SC8Rv3TkHtF57KHySCvBZ4NQ+zQ3lA4gMlgT6T/U+eEuRwzCgIkbMYbZStJYv5L+7H/W
Es7kV1LZ1f711wi9R+v3gDK5UqhBhn+FdNXn/iG24qQqpy/YwWEnwZg1m/yvBgYFZnQiNMFnL7RH
pwrghXImTxO1W3PzxjplrTChwr8PmHUAY0g9lco284hjNV0zgRwcm6mpmbEGegencPAZcKJcwGsr
JRBLI30/7xUTZqshA6bjYRuwZpVssxSgngCvvZ7s16UiJD7w/zxwmP3tIlQWziv4xUSeM1mkWB0/
+SkaHK/tgxuxWXebg944epk0uQIrYlkP4UY8vhJJsBW7ui50V0BHPCU8kEb8W5JErf7maTG/BOCm
YPTEoO68Gu/UodCqOFY6CXP2YcgMzc5TC02VEztnpeEV96G5CmqBZpZioTb89tPESkxaEML+bb5D
Zjvcyu/+psvFUdo7p7mhthAT2x/cIZCpPmDgX8wDQAAlhC1yFHAxjcMfD8BKpp9/erJviqEC+rBi
UdBAvek3aCkLrm28OjuUT52bvwUbDRoW78rHelxWPz2hem8Vsb4L2aFf1Jurq9sXGRBb98xm28RM
4qMR+aq2OYr5wyqBT/vS6aOxalblqqqxRAKgvGrkfYT5Rjf63YO+KilD+AWKMT0WpHeHMU78p1jW
4hQAlBqoGmDx4QwXlZ/4+uhVoazgDb2hmxg0mPOmyRxzQn6pyZUZJUpIc++qlkQj2UYt/htHn4Eb
Big/PXBqROvSfOpSUvliqMZiJrRHG2JRJq4/+WCRnmlu4h9YmNJqPWNpzMGiVv8yZ9McMwZfE/7M
ntEHuFIX2c72RKJuYHwnAO3cejGfMl5+uNjyyEPRsvj1F5zxCjaiVwVxHYbKO21TVMRj4jU0eMUI
YlqHeewjr1Twvv6WefIl5cT5X2/si1gOfvAEJpWrN1NVFQ2XZq6VyRVLuytzU7HYYnt8DsBs6H9N
Iv8dpUjw2l0sieR1FrGA3HlAQIakCNBarPdwLRydxamWiPbCgysLRCKKj6YKVz4mLRqCApk47wEc
sUS1lXf+sPo0IDtHVI5vJOMi3wFNanomfYU5Ng1SHuliZpr8/Wi1EUn+wnh/yVlnKFLnWmT1Qn9c
HjCUX7Z5Z2/gvlbeILhTyFyK4X69o1RKlk9Zad6vNFuHdWGYxzinvhUdmxaDxpGRcEoBl3DQhuJp
NQD3xkdayJl/efbeLgSADfhXcs32g+NdTbYh34p/Bw1Bh2/vBBnTbqAJzKBsnPEjQWMJRm+yJ7Az
NXMYgwulMq251lYYFUjsz8FM40G1Zq+efdC7qgyA7LUvj3F9o3GCXaY50dCLaM97J/hWreMj73yX
dx6tkkjxiEeOYRYfowXxtZ+bJmvWJFshafJ1f2kLaBhVU0GOkCceYc/Xy3Wuk5GEmKCde65TWeTA
YZGZpfRTPoElCTRkGrTbS+OvowmOrNS6Hw3SuvRyAJRPFb8HRQ+fKqNhqKv3KefkQStem2/4Ozip
4cbg53hRCxnv/S50bQxtHevi/7x4Gn8dl6OYUeC31iBqLuMxJiBcyLAko45h+4Va/+SR20Tq0a2B
5B8HOIEqUofWjBuCJBtBuYdZU/5fgP4IBsrsm2XR+N39OJXBLNf66ivnsVXoK1RKz52myjK6fbfl
7Un6lJROkbJAINT4rE1bR1re+VuQ+KmzI06O5we0amA95NfqTZ5Iwb/ZzfUg/vbwMzPEM0DD6Bsl
taggQqak5HCX/UUHeB9ipkPbMfyEmLnJ74Td5urbIIsQ+vy9kTBuY54XSI1TDmVanCEMok2v1N2Y
Xae/SYVoMUrAkoAGDmVmbgzYZbTCWy4FcyH+/Fcg8yIQt2caeF/TuN5CrcaKc6Jkz+Of8InBKdaO
szDIqEI6c/0MqBF0uMBc5Fm0Sg1BQF4Zund/84zp1yMGu54bSQqqYJWeWp/0mOjliF/bMskxjE3Q
8u2RAarZa0gT1rTdXRFxZrxlZaKrmXX/bQPD0WIJETbJGpkHmMK/WBIy64VCe+1W82i+sfYrOa60
zoeVJjBNGaERqFhtX1wc7twQosE4FMfMAcOQ+PvmAVcjYA2Xs1bE2CIAH2S/fab/GCYOFa1opGEL
Gp0mZnjQ+Erb1zZwp/uot8pG32aj55Cte31bpc/GHp+ZyX7ODxogI4cWL42SEtuoFhAxSP+wL/3V
E/wVJchw6ZHaSxwyW/RGD2Mi5oNtH/5e2mmWG6PHj6vw7yL90WoUsjNQkMYbQMX1lrZCB4fTxWd+
cE4SDM8gy1HF1h2fqQ5i17aMOsM8tKCgjUcduJCwaOcspZoKrEbxuw0b1p08y7lKrEzBaHgodY5V
Xrije6K9iEc572cPe6XzdGb3UvVcEdM70pZr2vivsO1lbar9s7mpjc+W9SgwoeGe80q9SoKBmBhS
Yva62GG8/WMv4KDTIpjQFAqofg/Hh+RTl3fEIhU7LCIbxkw1lkKHlmyLdRlYAnj3hTAzt/sfqY7U
RkgPWFC3Ij56XLOYLE0byFy8dAQY4HhLUBjiWuWBdiDAvMdujLqfs6vqJeABtVAlsaVYIjlUDwfY
H8DNrZe94ElFo6YpBAHXP53C8T4DoH+ACC9J9zg0TLXf8FCo/ZOTmY6lzWlhHGCYGT9Jq8MnYCxn
g2IAsHGwyfJ8iipTF3a3RZRCJXtyc7R613b8ksTgs9iXuFaBqu7Y7w9wpi/wkTtvfaseOvVVqtVI
sxcnx4RMP2N2pUiEiwsbaWOUFfZ1OS96i2YBp1M+++tgmc4N+zJ7Si8GC0xAnqdFDlKOA+CceIXv
eU1ijK3X1psWgQRS35+2t3HC2OE1jAVw2Lt4Yqd4289auRfT/K/bfHI43r/LLiYIhBgAi59daIHa
fWVMxq9DSXpDR5nMCmJTjshCAZej+JODSDRumWj0GQlJfHawunYUB1fiEtZeMm9+xeQv18dTSd6n
E3Vacs2ggDyMkiRykXKgny5/Z850hOfh/I6f19JBpEfLKAwmycJiDEwglMfhBe8DKDmBYqbd4btI
aFuzaHCbXdKqRv1BvNkR+kNdL5I5mwifb+79IVlJPYTB1IoWeWH/L1CbLGmG5DSwoP0q7bgg25nc
nnXMIMya9mZ1gErAcyNaejJ5dCPn8en/LaFFz4qgH8h2BhVNeT6UotkLCHA1W9kLHe4BqFqF1nEK
QzC0VkXZoXVAFFhy7RPdlFcJ6p9mVo+8YHGdr2c4rpEeURQykhcTPTiWv2SwX0DGdlp3nH3MwgVJ
B0H842yOXg8DJxtkvRkySg5yhEUCpmP2YDhanJN7FsyvYo+2uC9wiubfsx6PV7H5gaNNIT+rmPYl
lVSo2ZsjQpgDW4nE4qam8ST24E4i3sfipWYJ9jFyHIv8t8ukutV3NyCE6D/sCJBapPhT8Yn6TJKg
eXkc00AZG1dXllPc1Y7cINlUxCaMFJotF8+JsHf5KdK2O+cgnKvue/jmnL5rtXy6xUQ3akCRbwUn
UY9erILPTScnBeI1AFbQxkBUQF4OgDsi6Dg+WC/UybqW1BbzWflS6ZbCPovwfOrg2zSDnr4YVSGx
tv/fSJsyE3Yydb7LX4lnKPQ8WzZIRgTKrzzHCWBoixAd9uX+GsK+Me0YOb7gyo5eWOOxOp15fmls
H7vYHrdWKOw8R1zOLE2Us8gVSL70Qu+vZZnrAKzJmJAb13lAY3Hfufig5dJhBuCPEbGIU0SBwnee
6ZvdO6ZZVaoUYma7nKBbWA0siDPDWDWSzuMg8IYIy1oxVShUCk5mDiPzKF66QrUIjFH/Kck6U0Mr
jMwCOHtAZZ9cko1hoTH+PVHMWB9u6giil4eADfTxN6FiAUxivtABzC43EZJxUSoU4s9i4ohOw0qV
/Y3i/80c0cbRguicFSf4l4yr7UkPeB/hjErwUB3vFkGodtjGxuUYpRUb8X46wfXCl+Tp3cKMJtf5
YtFYObTRU5U6GcWFekFGwL8p0wk4I3+3HpYfatcRiHjeZbvOCgCWOjd8nmwPYGUcCV4tpqlavcKt
ND0iKeuCVZ5goHIMLhoLL0vvKx4J5zUOvjrCWnLNmeA/J/qvv+l5+PyI6wfFdY08BD+zpq6Dpy8/
yOj605DdvaFBqtCmG+UaaSFnVQCSOdaOFT9Iu7IhVEQ/VXlYiSMG1c/DlYO0wMuiajV55BuFLN8B
5fK6eyzuskN9BEuFYYLdAOOcZMveRKjvgg+TLtoS+Isj1/KyCGqgah4rL0HN9D0yi1usZcfzTs+M
npePfJij1CMUUqquNxhsnQM7FZh7s4zE3rPVi5GUDO/2EIJI/MtbhmYSpmAhQbSW2ZbnbRs8A9/3
91NRJ1CwNgYPMSJhbXCZro9L66Al346NynndCwvZDqIITM2Pxv6CjvnNCrIukyYO9AmwUi9aqulr
kqKpX35lloVk2pER4QBg/S9VvXlGfEEWxM8OqpnFRX4dPb4BwWJjr6b8+CvcARdPvUfXroUw2Zho
Lhy3JJr3DFCuVdQwGgtT3avt1kDJDtCtdKSn2QNMM33wFffBkbB47gLVtbDFWD9TMMfSb1Ffa2yN
E7mPWeqFMrEmdCTkTYmmj/RGUoc73hrRgj7jqk2DSVzYhtGCqYxnrNUNUF+o5OXlEh2Kw6Nve9p/
iYyFQGj7gS7gGH05WdH6b52VSGSDEe8YZmSU4Ot7OlCCXCaI7knhtYhOZf0WAuOKLhrJlYkoWYyF
9vvN45HxEv6xKaw2XGdMZJPZPBr2dk9YrLsQB6B5bcH857TRKekk7A1J017thltxHfRpOtmLKrFg
x25e4KtiDIpJzO6qCDSgRte8Gk7MCgDgLSc85OyfSQKpz6CkWcBX7fy4N/YnG7pVs5QWKibG79/i
F7VMs/JNLLJ1BnYgMP3nQsqVzZR4OIBbDhk1HU8IEng5mhJkuFeVbDOl9y9qAd6UeTAYf4x67A7w
vDldrdiadsKnBtRx8aOIeV6EPJTor+nqveo2DTR33MIJ28VltU3PqPZ/chdwbmkRr4ZFVobA0o15
29AhvNUkwzs3ekopnXSk78Ezofv3cXTxXfJUPPYGFakkFQY2vYB9/ngWJmODySPG6tCTpzd6YVtx
QEVEiO0A8scHZiFopRn1X0PhQyoxEQHr/dOfKn8efTwGSGxiTC0ucFvdoZQMqPSuGA7RDWoErX4b
6Y+Bd+r5U25B5JGX1KJ4Vq/7pX1ThjdtH5A4RK+xP8FajK+OHU+OysUVYB+hAIL2bwGaGJmetrIz
aFm53YxysjsXdlx48DrT6E5tUCHBrdbPHTCFGMIdBIvRNkaE7HLix8rQko5dOweW95LnG3BhVHio
BwdEZatbf/O2Z4tuwp/Jj7r+vxIo9i4dyrHVBc0/rQ3uJf4IFAyUPk4FJbu3IGfJC+tfcCAEl4rU
dr6ZVZuQEXi6nka+WI3NfHROVl2f86h8zqCiPCbh7GIthJLpkc3W+4oDSsThKr5bHZhMznyQgMae
fbaSwyL2OFrTeUyoNFNsYnpeJXsIx63vESAU4ze4RwLPUZM1rCWT4mVQ4aIjsP7Z3KmMWNOSHCbL
khZ9eX2EZJfQimSjixu4ebIgFFg7AZ1FrNUJz+xZbZZLZFvY6Iu4haUg+le23rd/Obj4ThHZxXrB
S3AujNIyTK/1Y2pYmETAweEkqJPJ1IobzkG2zg+5287H9P0b8DN40PMqzFtsP3ZE102NnlqvamSN
Jv4NdxMEu0j+uIch8hBHrhPXlTF5vIGeXGDQ+bX6ptZJVmI/p8cJ/AfJxebuLTHZnZwdyhT9Uznm
XJ2Ijq66Q7HuK+AI/qzNg+D5fzwv75OrRjhBnfFW5H/HkMhcVqRFm7ZK2kTMipHU4vpSoBB1aPkx
MeTsKzBfRxkp+TLFAWwLPXsVCnToair7cGlbMECfs6IgjXcPLdWQONRwVYNGwDvejoUTyYY4GI0R
F6daQrFSD0xHbb+3DE4D9bHT6drN5W4jR6QS/k4tp8Vmn2yWMOWngd4jshwsXpNG4A1gGVjeNQWF
MtmoDbNpybrAQ2/kFhPR7N/E5gmsgKSLDV+oG4UamudVOZmUp2Y3QXqL4rJC/2BFtxKLHIv1Mme3
Cd+B2l1xTc6oDnmOk3KQ3QGiZ8u7e2leN+lxvVkprsv6ZF6ZAKixa1MXrmflG3SZp1iKCNGAV73l
4qbQVa4ypedVl3xYdu+Nc9amQDCqPtXcD60Nf2T7gzWAk0kvigvZVnBJ4UDgRfsBPudF8fcVGoVY
l62PXx0xWdnNJxl7TgXn5cAMxfNAYsySr/ndgK56ItkmXTNw8BwEUoe0biAJa6zMt0lG8SLZM/jB
zeLrnRdearBuF28Lcxrdy4hTVqeLHN4kqzGSltdEV9DEh//0PiwErNO3y+k2+dXUIl4K5yESNWHT
F+JwF1s6Fp+C6jg2bCaGcI/rY6p9ubCaUU3g8VmnftrUtaDdbq+pK2qdq3S7q6bNbtOV6cejena/
iyZftnA1KDCrHB1+T5Uklv52aDX6zR51dW9jWUNRwXdkPDihMrGR+pzXA4MzdAIQ2gGcIAuucBLK
vEHJqzA5xyFwrj/ypTCn/CIo1Uto8KGfTY/BDkTYICKUfeHQP7d865cJ2nyKQTCjDhob2diro2F2
jnsjNcDc7A54yhvlVTsWbgT7Fxc3NDfMPYJdaKnNqEfJYVqly/YWINHIRUMSYY34DWD0YbH6emBA
ZxqKqsHWaw3dwY+SpHqOVDG62YUwixEbLJz6ZHoYrvzBBsZRUFVGnVFkdoQHjBBClyxHk5MWv0YO
5oh68EdSHYZyaN5OKJCc6dubwX4CkwBY/ZE8j4hsrdj3R8Wl4Aa2cSsGVigmWsB7Q6N3Cl05JCoU
sVwhiEmi0wps+CfNEwga4mte9yd7Q6XU7NkFCI3cXlq/tIIpg95Ok1SwAHUUbrIH7i5U+JEYJ7Wf
i+RMCxuCax6EW4qBQ7yr9Xqms3Ah5JRJ+BOiZi8Xe7No0watwTcvF0QvSE4tyPQ5hB7r/HGYflQQ
4gkzZz0e3nOb83noGIl3DUT2V74KWbGkEi3uoDBUxnfdF6T5vZ0fsqEp3c91PMkypVM5DlsMFRjt
Ba5URErx6hJYujw/X2ecGW4rV4/Lp96NS4mw0RDosTiTZQzi4oaZ3ude8daAomWzCWcUn7Et63RK
2OGfp9BMk3+r4B3DS+o/c/cQube+1rLIdAu1XElZuGBeRphe1viQ/CFfXSu5B6jt8RgdWYfzLLjP
euQBr+YQn7vCTyTTOozKPrdhkF6MrgCvNHIl/EyU595GWCeY0PAyZJ95yvWXBwNRW/T50YCtbMiJ
t7pHeTK1YUksQZ5ClErsCYt9FufsHB4QvM1iF9hPeKrjJCUGQ0B5zEMqub7w1+BjUn+kmV8fIcSl
ASLp4tnl4ZK5Si6yqdxBG4vn3fKN88obux+OsKkjE04K891UXJdXhTADUlU1HqIDHp6yAkmNQyah
YHQL4Rr+uEB3gLpAqYbNis/PGOkVAGNmHdNAa72fNLBEmKaEgMy/mgqbQ6FGIpCUaoBanuVKNoA0
Dw6gMUa7OGecC9o5I7aIFr7eM3HlDQVFVeu6X/LAJ+NN2O+8wMwVto2xwb2K2ANPmxqqzsnrrEGH
di/MtGx1N6o47a5+lju0hCPeSwTHY7nXaWKyI6muuwKS13haEa1TEclryBp1gEGjQwzDpNrVEWhg
t89mC3pybydLETkGnL57CazWdwHqbrbj+6e7nuHTPvF+9l9tqfTJ/pFaMmSGLogPnPW4yrPVmAJo
I3cBq87VFyj9iY0Ooyyr0RnHoWUN/tTKVdO+47xeGR3oSN6/dXSHezHdUMqUebpsGDXvStOVmhhi
V1o0uHN8wqT0sapNWAue627Elqjvnan2y65OlywEr4RrG+NqVDobJuPIAcC0AdXUupbOfqF1xv32
FnmsXuk3iL1mY4V+fN9PkZgQTA87hG0y4gsDdFe/hCdhUU2TFSL/WO3Djmch9B4U8Ea5gooMZlx4
oc+xdc6Pk/r9AdXGKGAwsLilPnGQ7jFmHCAGVn0/2smgnOY7d6QlOJQq8hmWSYySIM/689lg7L4K
3v5ccGi34q97VClrbFz53v8u7A8ecZ3NVlrkWi3vaoFy+BKQNGkkfeydtLd2A7qlMH6YNasP4VVR
XvpH6PwPK9HYVd4kXtIpGf6bsl422+C6mgwSdUM9Sg45aMPLToOhEvGmF6z8nphYGCB6/WLcuME2
lOq/pmKDCpZwaRh4U5t5K/UHG3zEWFmtf+mRB8wnDErxU1M+bpSGyGBSTPLKQnsvQUeHnn2IRZyG
YXmltmbSuuyH5Ozo14eQ8b0WenTv5abKJSnZhSjXUonscZwcddvZ7gQpCE+Bz/DSJJlZZpIJ5KJL
OtNYmW2uRB+Cyh83tcf7K5iA+xIxpugm3K4tzugxVyqc7G7+m2ZVI/QKi7nx4/AxIC33lgdmtWLn
I+6fr1BGYx9WwfohvCzdV3wyBZ7aQ2eLapaqLjFPvktuL9DDp8+E02RLRO3B7lMcgH9PBg4JkTtl
qPo2DmljnYVi6GZ5MnDWRKHy5oYNWnsj4yZw1cdoEfo4AY2GoRmOLF8ra54LDoe32Th6dqdevJzm
rwq8Jt2twMGj5CAbiH1SAuknhmgBxu+06q4jwkTk2rZa4FqsMdpXV1vtq6y9Z8z3ALaoNipaxGSy
a9i4VRtyYWhkyYOTusIT41eiiKD7fDTtzEPawipfOVze5QZDiI1spZEuWx+PMZbwY8wtcU7kqjI9
twMUV+eK1+bUo4Vx80771vT7f+G2LibjIP5ZOD/0snjjsoKSUlpDTUaJSPiwCv3ZdNHu8T4YdJVf
imBX7CkFXsbp26S70XEDkNx6U9fcqa7WAAe7UyPAgq8+clgP3FJSao9IJ2sexkgM2Aqh9gZW6gxo
5PHinPsUEDzu8mIVAKhjiLq0/+Np8wNJnMSeiKMOdJb7GJBepSBDW/NP347Cv5P2SAqj5QYLCQA5
XM25KkQEZWquZvOeD6Adtg/vXhSAtLQtRz7xLRUt9E0ivRjv2lZopo/x5x4ejgHHaCgHgWVgqGWl
pVphAi0cSSGw8SRUN9+d8u0nPUxZStjQUjvOd+GAjF0LMV2qKUaKWx32BbFk7PI138fP5BUtGghE
uiLPYdCEO0+cwQcNs1v8BfLWcoY/rlicoi3CoZ9nOPJuSqB92+/DA3o9uOGkyJWn4vm+lGNCJ+ft
VyKxKmbVOeZPn83dc3elSDEVI3L/aZB7Ob9GCbth7IfDKhDY4BDW0q5hNrzumT+Ks+dZNvzjlwLj
6CIB0gr+LJ2V9lQE8uNnx7wMyyRTIHnIfDi6auSWW7PWHSjT9xsV0sxIq/wYVyYIrBKr+OG6rhQ+
zJyvZbAWF0esYbqgxWXZqkwg8e3m24oxbjdlZcrnSGHt9BNRj+NKvh3kVa1aNK+7EgiYLORSlpbD
jrpOGqRiFt1fY8H5q1Cum+dEVu3AtMh7hVtPNlJw/6oAq6Fj/3qER9F1f73f+QIzKADiSyl2kTVO
px1riRmjpSdbZzVlyy5ot+Acm21U69LZHGT1wZn1ZsbS5D7pDB0I/IYam/GwvFAzppZJRQwZ+xd+
uWJuHzOJHaqkeJHpz4/s+s2mMubYdI90GOaroPk8azOMlZQ+2Gn4TjMRXtpXGyp4IBaghRLNs6Mc
8GWgjToTLK04gkuf91sAModV2JtfFPikrzYumtEb3kMjETWLs7NhsjPQQqqON+M0AScbNoojYEum
iv9UmfAG25PmcOFCSWnvH015qAb0EvOf8yzthC9TA3j0bkxr8rSDUJbjhv9epQQ+jFhVhsJDY6A9
bjzC+tBRO8xwE+ka0LLnAcn06D9CTouG+U4YDcML3u++EMsB1/l4JeD5AQ+wZlBKOhAcTOWgn0eI
4xZxO+OgGDd09egjuhP3wgyd55H/vGqWYefTRhsDlin+D3gvLaxJTvq39Qzx8RT1dnRpJ2v+uPMC
p3jX+ybG0UTcdVoTOeOWtrVuAjkVBvypIUJfEAQ5m3do7T/KoDBtRgZ5eaHAahdNs3bMDPxN5OOH
5rqSqyBPbjtJskdB6bU+a48I5u9MkimVlQ/+HFiK8c7A0U4Pyb2PknZtHIcrBeWm4rOWenbTjjZ1
vfJAeBjX0UkCwZHXxVn62bQj5WAyjBDRHU99C1SsxDNXOvGBBIhDNYwZpMvixC7TKHgzLxs4soNa
R+Eu+4TYr5TqHAXoNyiDQvYRYbm2xbVG7st5LrVEmiMXVLNWFOJtoruKZijpg0+GH9mfkjASlaUs
QG3OZZKKQgr61CIn3yl9lkvcTkKQs/NMnphFQCcgYqozGTWjwyMmelw7WLVzA+aDHpXbqIpT7YrS
AkZT+TSpOu6Ds9xXWat69JhmXSL1mZp8N/Ng8YSDBUw54KQzFqEjNanb/2xccG/Zz9HTQ2BSJAAY
e5/dCcC8h+U2XSQkcY8GG/nhtoXVGd8hUBnDzSScCypB9hwRQkZ1wqkUQ9GvhTtxbWvzJ6srsel8
c3XnPTYYJof2JA2RnnI8qwQsaooLrWDqT8BImZDY8tKoZyNKlJphg7+fZw/2YVVGB+ppmxPDPtf3
yNbA4MJntgLuCJaU12jjvOKFDutswpFhw+g7FKpsqHWwWnU7MDI9FY3Kzs7VTdxV/nWfz8Ce4C4U
BfrrvyrX2cy+LmN5hwpwGpRCIdUsdikQpxxN2I8YsKEuOVGW3ub6RLz+qRNJF5KbMC+NHKY7D1Ks
jawdQ2GQ47U891F32GjxHkxTFiAq5O/llObRuQKrcXqU2gkxH40YKj7Sn6O8XAwxhsQWaSxF53mP
/klpSr+6n0L8t2WFLbitsgchzLNyneTuiepsDsyBrkRCd6QmzrMfns/6shycwdDijH9C7nde+QRi
bjOWKCbpgadT5fXfaPr/3tRJ2UjIuHBTAj22qAR99o/M8lJX8uA+GnZYmntge+yYniVC/h3WlMCy
cnepl8fwmaGVPqQKtF9pJMc5mfMjWel+Pao/8o6MgeuNW4iAVeA5jIYyuy8M30hxVHkgKWR4KAB9
EcLJC3q0P+dpCyLCIYB3b/Hpfja8S+9sB9ED1A3LLinBNEhn2E9QAWV/XsxDdhaIZU9BXyYVyKhA
R3GeNLJsLEPsCPxZT0wPLjQIlXD5hPmH0vda/ITpBdaXFqn0r9AZP8xgu+GUirmiXzBio3edTqj8
V6Z4RtJ3KE38Z9DRSfP7WYU1XEM8qqaF4A5uVRAWhkdDBxMqNiVsskPkOszVbyXTs2dRb0gUU4x7
BAXIOZVTfDvV1iYq+fJ1R+AstvNPL55ELPhDq4Nv02rJVwW9QBE2MYwXun1nqN9cfPYR9Cd8oOLz
EwJzoL1CH3expXMuQlBLkENFvvFMsN+Gh4PLEcl3UFieKzKxy3U3MmXew0r8No3xl1ywjfsI+RQC
LSGSmIF9BEO3EnGd/zl2M8saZXCczhZX8igQrEvCflbA116bawcEiaahlE9BS0UJ/WKn6Z+kWvQY
nwZ+UQfQp/KbQN7HUJzNYYWaWYr2zCDvN0dOFXnMkaJa8tHg0EBwp3lz31eviJulXdz/ZlSk0zxt
gQ0l5dUFe1JnGjdPqr8V6Ox/e9cRUZAGRREBsr6JrE9Y7eB9oHkH9se/n3zAdL67uPmHro4xGGOC
xWz9WCYt5SXkSlkVue0wFLL6eeORIkBQvmEkiG9r/6ahuTDPiMOW7lQBrahQqRoOu8j7uMO/iL+O
Qdw+5IWQsUV1nxknLgxhTljIPkoc9vwk7auONsb5xs02VA9NlhhrKyzCsxyasHIjALHEk7C29zsP
Fos4lSE0ZpKY5k5fh5p4qg6AAUnxJ9KeZm7pBH42Gmpr7dUKfPyuij+5bh+b732r2/Qn3oBmlCPc
WE+yvWXB0XwcBHhxxxtekODSMfHihymBD07i+8JRFPf4ZMh49xz8cEC5FJGSL2p5knVoDd90SdtR
l/FunmSdza97VB12PP8SGkJwj44RPPqM+DbGdqgPyfv79BB/Gi9M2bvaSus5fMtIb0yP6GCkiFag
8+/qWIvINevFZ/oBXWD5r7VOZJwiJYVHDv/vda0InswzBJyN2M6LuMVEeQ0wCG1OiTLXV/zKDVBv
3wiRS2M5ey/BmIxg/eQpw8Vt/nycqpB5f8wrYEgTi85eHaRZbVrqFMXkvoGlk/mZ/fkJA5moD6sO
QhhEAuTAZ33X6iWD+oBrIShfLbqGTYPPdggepqcvZUClTyKI8p65/xkuTvboBQu5tcFai1s7DXdn
uKmfu8uEenGi27cBtiiPIEGcsnQTQGh0uagHcpUNM1Gve0W9n6lxpI7r2HOQACWtcaz/EMbPyQAh
JtevYWt+fXn67YRmo5uC7TXBH/Fn7wJXbGQtbwvZKuR9pV3hMqS/mCxihBsBHkROFfEFt2jxdlXk
BmSP2lZQu3b/i7ZSecQG89YPAYA795YppxQIxkss2hdXBOXdd61CkpsE7wPpUsx/h9ecFnYj2Dx7
8o8KZkARehpVAOyvsUpFioSuaTCWQd1a7ptMUSeOKf0ykZ4LGjaESZdG4iRKbIC4GQYWP80lYzBC
GvBNYb2oyVkTzjcHDwA3mpIoWvck0IKgfNvxadA2bQ+zF+gx8S/L6QKE+xDR3gtkMt+9BzOsFvGP
q+fSKDODRBKaTpBb6OREAfHGduz9rz6FEy5kaZ5/WUYT1i4X43Cd11UJjih8Na44ceCqDRYMRe19
/z77VswLZF9q3S0d8iZZdvYVLGsmyHVgmOkVJ3pQQ/XoydiUnU5q5lphj04czbNSZ9vjZFWvpCHB
mgBf4YYmH1wjLnq7Qux5IxEhihJgh+Vu7RlrKbBzpRlkjS+Px+k1/+VGecu8Ghz0P8hGkJs6M7nO
QdnpfmvcxKC60EqCl3xJWnlAf99Ikx3cAYEtz0vcTmn3rAVSEipJROp/rmrPGDxOUiPNyh4rrtsc
2A2xgenhudqKuDZZ5lOGraPLgDcMvwhyYR26wwlCj8VyuhLAkrOqNZnFK3qm268DEtsxAz+z7PLI
7jb8sVSLkntBVRM7nrJMg4ANWHzEbRWGH0rnQJnqIkiozohMt5cCR51cH+WDBnIG39RLZCUvkLZ9
fUG5vw5h65I78fCCUrseY1rNRCvmZ8sI8VWy4RzUZzlBm3X7iCnUuE3xHWgmyZzBNyr7p1cvzDO7
4f8+bP6EGkep29UqNPVH6OxDCXvP6Ah5IIWy19n3mckxqyu+3mfxuuOCv6fsOuMDlznd/GJ60bbo
Uvjc1UhdT8WZ9FM+oAr8eVRc5VsWTxVL/a37BFQvxSCjDXf43xTtmakDxiaAW0toPwDyHCt9EY1o
i4Nf+Bs8fQKxTNsoQhqEeVRW2hqMf3ju0H+aJZWFdHNrNKvfRqlG69Osq3QCUbrEH16CPBRwzDLH
p/X/6PWPlrcln9PxYx2t+hxOd4TZe1r529LcQH+e3Yym0Tcc8YA9zrNbsviSliPecL5yDeadNKE3
nbdjtuDKWvuj2N0U/Brw92VPNwkDXFiKhEurQsbM1AeWGsFl7kWozyo9P2tlNBjVIBKV87UgHB69
XK3/eQtCUqgEcMDIwBKGoTr33dMNOxGtX44U8VDa2yQseFEeb46W1cTlAHMt6glOE6QyARN7H9Fd
QSRvZLzTObdPH3bU88kGOoCBv73fftqEEQ1fsxPbR1uQy9KNPCEQDjbZEZ5X/RajJj9DgHdUaYdC
Q3wkzPcUDu+lZpGvxLVnBNMApOWDZJByYiHjJlNmr8dbdh4xlMXvzR1XoHVFp1bctl/ifm3d6D4o
fUOjBDqrJ4HfB8hvSzW2Q/ROrbDmIHXLpMXKJdmJ7m8esSH/D6t9TgeE9d4Nj4DGkChIqW7FdV9Z
UPFcjD6EiUC12fvfAfsZNSj0gK75moHzqe2cQcz6PsetxEtKXg+MESaG3Aghx8Vm5Sh5d7iCx/jG
ZOAyK4mUIBtBwAF0WJ05jUZSxkJknqANVQTrnAdaWG/oeIkRhT+SfrLQ68c5mNT7zRBamkl/e0fg
tNvp+Kh9EfZTjLICKiH/n0inmzpQjjzDFKYHZBF8MwEu3vxWPMFFGpRNNUo1Cvl3vGInH5zmbe3M
YrujK0Kan35rPLSy2M2BTD+pyRYsupEWNhH4Ssgy1c7Gt8/G5scM3ImfloS7xH6ua7XVK59UylmM
6LgyoqbqEwMIlekxYXpx0bs4SyhwtSre8j5ALF8zJNXAL2XVpaAosD0XiKu9mx5QayogcZuyj0+/
xMPUXPSsAnW3qen9hOwJDvdYmCsMsxtZcqHVThO8xsCWJP4aXwphmTLLz/9oZPSbu0J2UbPAF2sZ
ApCX1vCZ3B1zsE9dpa/+lX2YAVdn0AaEZEIqzqWG89QwezLCGPEPLBwgeavX7o0h6B9w3AqpqBvq
1OvTJv0TxahftruQFXCx9B650WQsR74oUlMWgDH+LXrbRQoH35TXACJXnhSO9HMpodhGJzBz5kWm
bJIXqLodkrbbJTETZiZYJj/vauFFk2D5Sm2HrZ/W2dUVWSvMV2DFXQ9+fSa6m1MfuGmpS/oTVS6v
reL8SWiUEjOEccwH2HZJuOyAGzIs+dfIZIa7Yw98MzC3gY9jNXDGj6Cc3/+qyu4MtwuClI6MkVMO
IGQiJfMmWqNOKkresrSEqx0r53x4bTWnkkYbO6N3/Z2wKszCe8JwJw5z4d62BbOuBX+vCDg1PZy5
IJk9J9McmgJvHN46fDfh0oaPfEwPmx1R2K4gFlarhBq+8AHOGCp2Xtny9GkENEMEFGhOTImsAS9r
U5T5gNvB/67qsQiZXZ7pgTt+CoKSGhxNlwPv6IAwDe/rYbAG5IpNeaZY4TMbWxzdipvUXpuCQKck
MGvSDC+xqo8Q7QXiKLZeGI/crn0G5nTBYHe693rXjzSOpA5rRvbdmp1RAXfEyedUVmnxtdWeY6RX
sxvYavetlekCuPE7S/yL8tvwG2GKmKYCpKO3nVjej96i3DZ2rL/+25C8HA/749hmyQceYbFBX2lv
FIA87UtsjDZptayZBPQ8OVRbiHt/KFbIZFWvpdoMC9Qszsq2A/blgKcUqBEW7a6+5Nkwn1RvRfqD
JrcK5dnavMxyPwf5sO1/vEhasuGcBx9qsJyaBlx5BhePigoTnq/MJ/R6s6GxTzILsYmzegxkkxzH
KmIdxtP/12BYjKxCdJ5XnfmBR9QG/Kyn8faGbvZDmLn9fbZ2eJN06433eu7hoNBvMu3TFYUbCnxS
1jwE1MkJnYqZQfOLNS21KJbP23zOqpEunqrLmZgJ3v3RGxH2er1dZ2aYOhP6gkmlJ42xhvtqz6SV
hryrNk/hQAQGdF+0vOuiDcjbFe5a0Gfc92Xsj8/uWqf8RjXUnZmGUE/IuJveYUYFP/rYvqfcylRJ
r8+GinPdVOJp9oqN+faFrleyFx/AUSQhqkxFBc1RWjpo5lCe/OPmm2AAlbiSEFTP7XmW2j7sJJHG
7mHpa2GuEh9D/GWdWnD8XiFSDLZF24vBrq/63M1Wgyo/hR3g4weGg90SHqLCBwHp+wZ+ysnxpEps
qDcYE3H/cRVxVVnU4S+j0RxGKiyCexNGGvJ3o4c34zq3OmobCTH7C4Jhgf8ac9rLWiSpvP9GJ2I8
/X+JngzpLtH4ck4/g2b/LFddVcmcB/Yu6Ix58RL6B+/wkzmkFQiHT3OIOTslXO+6GQGdbAFtab9l
/jUwWcHex2tjk1JV2Fhl0FA0BRFvov4VcSVOEa9yOp8F449r9A61jOTO516gDZv/Xg3xdBOTlbki
9OjwxuRsQLxeJgkjcQw24IV740PIdHx7JxCLehua9/Fp2v4BItzkHrxp5ZDGVUZ0/QqB+iL1Ubs3
b58s9zlOPjMn168RvchY/W0BwmwBpVI5IK5Nwo8Mbu8D6bO65nICVgl8Vo9eu7HUSHFMnnIsOWX+
3XvKSAf+0kICq3KbeTND+eKn3olustCGivstn1GvjjpCs3xbEK63PEAyICQ3F6RP1CaTohXPMLur
BRB6yR51LIhqNuas85EWXC88AEUcnSVf6lt1STbCLincnumbcFzUNgId8kH1ipcsqPdwSYab3GE5
YlaimJqfKWDx79DTQ6EhXsneaKw2m6A3UufJstuOPL9yt+0X+j1goYjVbMRVwi3vKnFkkHNZEGKG
gHke2EvJO4abLr1CuPdePxVlt1sjjHi/LTFMxUuRN0rAIE++QbduhFmUKc4Rv8RQwF2XoszqUxp7
KHM4+tZ+89TIiHJgmmeGKjGeqyUoru2PlojIz3Hw2RhwblBKTjBtULUVkZSK9jufc/E3KXR9xeXy
8CnIL4aqXjfJBZlb5yOkJttg6ZEckN6fV40H0jelsR2GjPhvLTsCboVOQEgDENwA2vey9gJj/zNV
FoaVptl2BQjEtRNBd9vTQadWg/h9vDe7PTiDWB7ZJ6qrDz4z0fDttJOuuet9KEa7A8nqK9qmvVoP
DGhexDYRfZc+QF/Fasz4KymE2ZR4ZfWeY0kDPPbHZsYb3dncxVgTqtpYeSX8Me/tvk8dhv6bg87g
mnnLB+Qy7Ok2Qqb7xt4i1L071SM/Nhjyman+8lHSjNFOn7UqCtPLBnB6ya42t5NkcYg/+Nhv78sk
zZdwB0E/xsMLYKDwhO6r9OHtqDLG5wQPwhSYLN7dfXbD2T/8bJ2T/+fs/92QDqZ9Ct9j1C5ta6Hd
fZaU9DP0cjW4rCwQM7g+r+pkL8RHt4I40qc71cGU1nI4jL8OL+xJhZxb6DdP0AxjQbBgwpqsB97r
gsnh24SlmupjMaoP+WpqY86+5Wsie8WnBfc8VEfvoA9HJL2+c//bzwmvfG7bVyrGui177Uwn8Kbc
UYkn3pdNl1Fc8k7BDJ7DVE3F5Ut81k64h/epWUja+qeZUwt/hSZ2sW6+8SWEJMHwO10uyLM5sPXO
eA9EtME7klQAuGQNIpR/BQn8eL1qWUtSkahmUIZEbYq0WKMLyjGfI25HRnpPyLNxPPTBQthy50kc
FzRWzNP3nL9kMrBF3d/HXbt1VdnDBvHxPeYSoZnrPM87y/Ww6iwFGpfhfF0ukhtU1cVzB6xzJpFF
09/8XAAUOf7A7rsRaQIih9PSL33IeuOAyaaYY0kbkuuUNCGzSly+una54+U2y5RfhP1ObLV3dXka
UOLjbq5+QqWDCZ7990xYOEPVq18VpDCDLHoJYScIdXuU+BYQJNCSonuVjPx28sua2Pe0AJ9kxnHn
2ws39ZEnSY2VntCVJQVnakIInOn97agd04XUtbUP1cEM0/KwVtN91dgjRWepm9pyfiSLNjc0vkHa
caSs8Hg/5W5RzLuenCYrvLpOaNPnjqfVdHiP3unIUOLGoJnefL0qHFBOmrixTvH5Vh56OueR50A2
rG50uDQWBoK/V9zC4XhdrMdaYXer7OWMWHLDp6XvtQNFmNwR3Trc/av6CXaPYBSC5Rcf4KXtYCo9
7To2QYSfQqQnc2TrNdTrAinsmbkTzD9DYt+y48RUIRItZjU5rpKOT8LK/QJz+9DwUjoyb9lEU1HB
qIdVdj9fGSweln+Za97E3uSWp5Vrn7/0PfIMo9z835poCn6qLIQBtNn2pjg7+7lU1StpTQR86mcK
exlkd6TB3P7bd6jth5QEaf6hXXo8PHhw7MbpWMnKpx6CwIRhM+s3Nrgx+Y3a/QGYcI9G0I/ldysT
uFn+ekcmUc/g1yeLByvwD25frNh/c6r0vFtZSMwduWbNF7oqF7JO4w2wvpHyTElLD89DJ6wp97rZ
GQfPc4NJBfBvbeKg2XitDQ/KF/KaiRgREGxCtUqvEdMOSPx/yXdAC6WI79ehCZi7MnBuh3q+VVT3
VVV3aGWXSU5MQ/H57DF233hNk8UbdFaURlKHfAJBWAC6DZNhtA4U2FuxQsv4VvWPYi4FwsCCKY8+
alQivX9V+NEGsqnsycFaI7UxnFlu3mIpbF2CMQwgjHeyCvy5/atLdWnbgAEUjvyaQJ3PiK78VHX/
+C/rM60E+P5H+EchoHUklej+BYAoh//WsKbYNUxuy/o6ibvrhH89sn/cjpPglcpq4eREFoybMlvB
uqRRBkElYIE54pNJmbWx2I5IBpfAHE2bYwfwyQ561d/YBjU7AzoZ0IE9Y+/1r45Jyfx8noNl2ZT2
If6vC0Z5u1LIel8SgE1ATLUGWmxfUIi9WBpTVvx62S7fGK97+barwFNPnlsfNbWmtePw/Na7QGCx
VNmH1FwSGXLWmHkohK8EwOjJtVda7fMXeTk1OsHUmaGOpjl+q13ABAFwlxfFjAo5yiWc3shajil0
MqxV5NkSRIY4HskWq/imIW5HSRwEgBtFERhgSUfoD3REWPCk9sUh3Xu4M9Rtd9QSE0wh8383geVL
WEL83rIjB/U3LW3unROCHJkxBDzfNFktofNxhdOmWc39PgQhlJiWl49kattv4PwZeAZFe6T7Tu9z
h0x7+DNJACdGGitJvsYLs+rUhmXHNcY5jg3H5cEmtcq6BQajEzLTMuvCpZo45M169RQzNl9TV6sF
WTL+YO1GVvYkaJtq4S9BT8XbJLlUkMtGEq3vfPF73ShF4fY0HJazVNPyfPChLH87SWoCyjwFZTAy
TiN1FYowmdN6SWgvzSWNIY0I0oAruV2jpr9XsS7uxOplXGlSR/rhpdIe5OhxblSbGVDTjkCzlXPR
syLWTWUD5xhO7KQcTxhF7uw/rnXqOzmHfXtfAudzkCJQ0ztYd0wXbZJf6T0VQvVNvuX2bsv4cxE/
0NXWI3NOxWfjPHddX4eUYjMEipo1lOTZ5eeFDVe8CeSkimg95/h5RSsBLZ8C1g0f0VqNXVruUN2C
v8yayyT33j0JOCJsGa2ZPIHLyn5O5F6Jkd1HFvclX7uvlWYFw32E2UYnsD7xwKp77HjYK49Vrhxh
GXgaJKH2AiFYOw6Ph1/t8ajUfIeAo5+8AsU3aVgjJ3fa03l/OZxfXfjjMTnKUGgNQx8ZTIqJjUze
xMTSXB26WIsfv8IltqjauT4FdI3EXcQAITMLwkKRwNG29Yte7niakZuO8vKfLVUQwozY544+q3hq
3H0jdfwQvb3SgjBUW8CKojNGAf5cZ+NFXrtXYY2VglNL66mZJWEgYbQIMpGFZYEUJ8RhFYGu/TYm
mX1IOUGw0UpsuBEQXwZxit7p77OVPwKoB2pJ1a0Mz2i3a29Wop8X9oskift4rSUC1IsukD7gcpZV
ghD/urSHCz2t2t3DfMfON42KgKBDWOpVirToqxkktIf79dwxzXvMNFbqN6+yLH/cKMjhhkBo5+56
wmL57sGbPlBFIS+6UaL5SA1Lj6AKtcLzHeZIfRpyEtcMgnIr1Z1x0Z2zNSAnpmg8THMzXaAhzi7L
/h9KfVmxKOgd30lkjaCKLqTILdYWTv37m+O/Wd+hfqjShqFitE3P6yRNUQ5R70IppGVzLKCh3lvN
rwJwHKXc6SYbfagI6bs7xDhK6YMg49g63cde9+hB4Xz5yc7C99cJ5MHFNmX5svrBNuU7pND5jZPj
0Ynoddrd6cTiqptqmpE/fJSmUot4gxmMlGvR24LvA2DZdbAPVlOHKxJA66ku+tkkIqXhlNOL93yA
hVx14Rz3jB9FG3b+WE9W/qVq6erGrcSNGaVBNRYc8xQ+g5l35+BO83Rdt0XmkJK2erjS0MTnVQ5m
BzVQhBy8ejd85iplZ6I6oIK5oOPAdpRKjiqIur/7n5HKGGfcdFdkJ5DYml2aJyB6FeUo4CWkkdPv
JWTBdG0+NLzuLAyVlFqUhXsTGm/HPbHevvrVX6a9DcYWWkLwG1nCFyE4+B86MpYZnWUjp28j1RCG
17QRipvshZzdZK+T1Kv4bxe9cCstKqKrsaKslkVIU0Q3lHvp/nWIYuI4P/WYkahfeWcCobyVR5vf
lLAGvP16UqM2chhWAOU0p/jk1FWcOdfjfZ+Zy9WTqs/TcTo/y1K844r6HyRn5JwDLC5gqhnMCgfx
A033ILEdv/hZ1GCRV2kLifW5hd+hxNR/+8GBz9t0sVuL49ZiHZGqPRQiGdQ4kKuOXGxm7eHO8hLc
YceTHXO9XZ0y87Z54pXd1PrYiZ4whG86c9mVUSLQ7RMK7veOb2PVeUWArVEJfObRav1cxm5/Mw3e
MLLecTNZxk3HhEnim+IylFhQGToAb8YiJE3rT+rf9oOwnSi4M8fCTWZB6I3l8mFHNTdG+n6a/FyK
qdbkQ9UwYyZf/pE+NShW1soMo83rxbP0Muxu/VyzbECtbWvqudefEozSg77uR0CaNqRq8h4Dp1Yz
IuWe5qCdln9Ot6tnmq0ImJkcxhiozILunM8CMyISlZhtYMGsvKkC01nDodI2Mp671tF5XJcbz9eb
+ne3cRyEbNA25944r9zieObuQTqNnnAZ/RKIAEK/xtnTfTxVgxE5JLqzb2LYxGm9Gv2IsWSmj9mx
25ePRArF8iN+lM0dqi7AwYAy8xRsLuTsGr+uHJ8zDQHs4iwtwyZxCzY0irHq7FHpuL1fRfssxy+z
sxS8HiR+2gga5oCYPjfWLOHsc/DzlU6t77ravAPCYk29Oilm2aoBNSdtLIFi6XKfzrglqX9Z5Mk9
b8QSnDORJdbWyzx4Lkc2aT1m5QdNbCvjNw/qds/epiRegSM1w8jPkUtTsFbNaDm5wQrlSz0+B+s1
veXkDyvj7iSKV8TOosXRT58KWsaChLBS+2RhOqChSNh+o+0GNeZwQqTKfvzn7MpkVazmio32Mpwz
o3lQ3XYA7k0vlEYVBjszE0gDAYaf5H9Ys/yB1te6AzwOq+Fe9ZAauLJ+lIhdlKoMJlobfeybmP+B
9NME1v55TXiI0WIqDmKgm5T/Ro78fDhZA3QF6Kery9ud4pU/evdxAgCHCY4BHVBXyJxQG7giEc7L
brVsINkH3uEQY4X1GlYGbd5/UhtpXXDGAqQWcDlFeIDK+P3I6WOsC2a/oRCR3dGWEtSgOhzEcdUm
3i3fAYXvoQPStmYxy/b+DlLMDZDXe9yE3FOzDGWGyNB/4ND2pCoUKfPkwAV1WCqdie+DARbAftEz
km6gq2+BMk18h71xORwAqVxarG2hCITmXyd0Gw0KbWYzpyrcks1UBmQhFAVJVhvK53hPbgog58gd
CKnZlqDX4oeVOt6s544uyESuVrg+U1g3JNRAQVxvaxUXiJxRDZJRi4RHevHe0XsGvppc49ny18+w
bLJtRhMMIHlmqqref0v+OgnhahPrFrtTeSkXU8MvaVQsMhr1xqHZGowvoAro5QIgoO2Y2kKXTfOb
N6dlPAEdKGa6ztZ4IULM8vy7uua1EGNl++DTfdD0aj3Dzv8Dsr0HFLfdolvTrzeKtRH5Iq0FlZfq
qbhTcOf3Sx/wIzAeKXpFEUO6kn6PYlHBWuhZDQBV8zApNqZNnVVqGCSgxl6QpqrNjOHsftBndQ+1
kZIUwEiMDzp0i7ojM6V/exVFjSVbQ5MJ8XwfstprQfdIP3TmT0665vLogBv2ajzQwx1zhdBfIF6K
bEyIAr93LZM42WoHyhqPG3BGKl7tuvhKxahRQOjU8hPbHumr7xpxvU8KpaygBbjmE6FFLhahABoK
qQfuXfHktkofbIM75lAQQUb6Gk42ader2ywQlkDjGNsTRMTgVCHJ0wHCHdYaMQJ8vGg2wyA3ECbj
itszgew/fi/xsSwlO9ZKv8uzf9TWlGDD9u3F/1geBU7PgspmNkH7IExhELr/+kTDMQHwYzAsQQHB
8HpC1bMXJRnK0ztV2JETK5CUB40c3E/eI6LMTRiU8SvOzPdRoL/aXefYj7o1r/VUm73j4jNeGQ1q
yN/G6cxj47sanDHjVEpThtymqIBk9RMJFegXWC3vkfi/b8+aA9ScAi5+4QYHlTxjpGIGEvV9nJQQ
qSKHDX7hKImECyEjne8Z7rpcH8eYMbb08YjRdtaElHQx4z4vK30tT3MsMOMgQCUPUz/lVaB6fun+
edo54StJgFJSPuGgDaC7HqYQSRZBIWHQMMEjal5YgCE9eF72SSRFtoxw1V++y53Xdqi3SiAHk9o5
vvIl2lIF2EepvSGIXmnHNVfdGH1fUx23Bgz7H/Ow7pGZmvJK91OPVt4AmQAlxo9X9IqXYdxzLYBW
Ol3TksvYUaUczFj+IssLq2eJNQV1Efj++717Hok9CCl1PO5sC3YLzqP5pBHX50GTMvb756Hp1kyZ
YZORJCuCZHniXR2VdvC/ZxM2NgCj2AAXAH1957DrHP7Stqin4AERPkmCQFq0bz5czGxly+5+oNdw
PfdK22TKnkGb0Rf2ZcE2acjIGC/KgGKK1Mv6he6sQttby+UmwplubBvL4AxVkULuhaZa5MHlsDB0
WLrcEDGA2UuVY4XIei6jUdA4rvCn3pSt/6B2UVmKo92BP7xLv+SZfpRJL9zy0dLBt4bXEdjqDqn7
qBZ+Dfvm/FBpOirSxWg/wzEqqfoHs7EPcMsNpOOulDNEwwKFfr/6ABLj9fjyvDRaTINJNsf9z21I
z7o4TyItDqZVirayC6QgmbVFkjVJovxXB6zKCzF/OQNTyb689y8vfJQqQro4GvXHvygxDGDiCFj5
A5XFW0nJtxLc6PP3Mpf3G3VedioxhxAbT01J8U4KyTC9L3yRRbTpG0n8QBfb5n64KQ6vS/YJ0LYF
5G8Fg0Ri3XlHft6knx1vT/x0EXAMEOUyar4zrGm/OKT9hjsL9+M5EcnJ4YFRe+wSMIFmmjDsYzWU
beVPaya2wtFOsJ7okaHx0HgxoQ8KcB9vUtUAKPWz138mr1m0QO6gTvLnLKK9mKgn4diJsp8SGB8m
553lpOtgUIzHWgHjdfhO7YxIIhlGKiFAcCuk8hAHOfHlaIJ6Wb0me+2EAzjehpJiLSmIKPMdOTds
vHeBi2IpoXG0hQyYO4AR8loKzi7dIC1niejwQgURJaeJYQe5Q1ExC+tK92HpvRTGAoNcBLG8h4DF
a4/WkhZ85lWMMkUCOCR+CakwP+cyWhXLr+eowschva5EafGyw6bXNBH84tjZyT0SFS75uS233KD3
gU9A7GYWkSwSeKtTQkGV7uzUrNJR876yOlJLe4NsEEqLcPldeIr2twFJZbi6CmDadUs9wYv1SSB5
TUUAdHSydCGY0aDpY1Nfy6YYEkovpaR6Xq8e1XslaMVihBb37ipO6o0svwNc8OpqAX/W/NKIlQPB
ZHfKhuzVTNKy4yhjcsK0Cwox3ONXPhou16ott+VC3zuKjeG0fVnkz0PpC2rAkSopxweeR6HIvDs6
mwy7l+N08klFAB7JcErlAjJV5yc0p2KnHQjGHSzHgG1fLmR12rcviuWStsle8sSleiB707sTimWi
EcYI8j1eE2JwLpMxfKrDQKUBB24RjnmCKEneOi9TbMdxGxFyVdb/hBaZJitDordr7QkHKIyzE3vA
rhABpk8lDDryTGjJ1REf0kd0SPp8wKtema098gfmSc257ZF1t+iRx560hwu/ltY/dtS4RqZdryiB
GOpqvdoqxfDDFvUNZyftQmQPjZ7BeAa508lJQEfOrrWoXSoZQtKKy3uX+kfG76VVz80GROO8vfDa
5T2ov889h7r84oiyFnPECPJNXLHwnx3CEqsgT7uFuvZgfDjxUlpQRMBBJDGTI9rJmW2e4KIHyihv
X8YZA3AirFo0Y+Kyw/cFGllw4ss7t8tl4MLCuHCFXdJHzci9B4dJ17tdUlBObTs1WjUQ3hDM8FB4
fsFSyUAPUPodeT90OVYlgycNFlLCnvRy0jo2+ULJDIrKanA4fYACchNYIfc0uQcUdtIua+L/e+BY
876+pent9Wv5K9y2Y+ES5DRxRtokRe7qANbNdHFPgv2d2woX9jS9/xo7BaFa64ZlIesTPJEXROMJ
CwOJFanUuZQVCx1c05bDkP3YC6aMYvUqoI9EX9213pWHoKhqnStuT/Y/tVqtyTOZ6KeoiGfFnnhl
b/5qDsKJ2c6OhFstNyTbjdS28DqHF6LSzsCdE+qIil4BnngHZ7AGjMHJWwocMJBgDvVNl60WPwfs
Ug01ClfWsUC1COzoEBKoIPdepmdoCtm2ZDzjjiYI6K6z/OMazb3p03B82hPl5FOlmOTnTxG0EVy1
uZzPL7ymtCThs4Cd51JmMrmYrVrHEgY4bOtUQqxo9n1mD8mTrBPhl129TPGcXfQhKgI6b9ZWjcJZ
qYfD/Z7Pi+SGrAN+WADNRE+wxMjYb+buH+al9ONRoayjNo+pDhxVqL+5KvtXQMx7+b6y9YYpTcEB
F24ky3S6xjCaDxDk0SPrFGpVLPsKhY6etA9KUzourLsTAvV3cnXTl+MaYNdoImR7VZe0Dynx+W8c
VuH6vxs6cwkJjthB+QWZrc1klQpxzLlFySvZppm6pE1xxanrOQ1EPMy7Hv9J+BXsSAx2LQRXDyOB
xW48jrGhxLQTmAhIR4o1HLpnWOlSheFBJN9zDiSnSqcq0/jj1UuerS7dA7TjsNZX6mS4jstXez6g
wLqAlqaNOzKaCIVnXKBcxCJWQwkfZXGPPDtCdU6nzb3w6ayNyX2bGIbb1FeuO8qVy8gNeKCAVJew
1flHLAy9C9A2+M+tFPBGR1/0jmQaKeA8mjeJBAwx/xc+Ht3hRp3aiHmLKD1xssbiyWqfBwUAVqqI
BrnjcT9KUJgM9r1AtJ0Xyq4UybHSQvcIbQErrjWMPpZnioUC92c2+fKpoHEAKP9TPJnOykSiXlHn
YUFrpFX1cUoS398xBR3UJlPpknilJ3gBgagezanQE9E5Z2g8kVboV6qq5bEMlKeI/Wj9VrEChdp2
V5QeU0CE+0P+vk6ac/BMn0aYKDoadf5hdOI4zHgj097bq267VJ7ZwM6KbeK56M9PQW7Xe1It3kT/
l/L9SrVC476QAX1dUIdeXgTdKgOAO8PMSCYibskvZ5FfXTsobVhZdpDRM9b2tbljDveuGBKPd30F
++csJSrA4J1Hqa5Vu+qrQIP50BPdh+LFk+Pa1CTepvAADHJQxB9O0a16c17GVS8g38z7ihMHBALa
L2QPLELPb4T/4HR45/rnkpVtRf7J4cSYe0OtSPrH/qps8/EdSaHQfIiwQqPbQvd4/ELgUJZ8baUs
xnYM+TczgzhXeOOtbcdbx/Sqkf2FGOjTY3yjTZMEnWcFFXlKMpX0Ga247QfX+mmVkCIZQ1xos2GI
KmlU8GOmiwufN/S3MDXaOWMVKvb23PMTrTL1a98L4+An1Xu5RVE+RC3I34T0+KSYeH/DSkisGPFN
Rr7GX65m1M48Wy7WIg09zRKTj8bok4DTmi6o/16QcZcFmDdY3MzKKlfo2xuaTGbU7hoq6rU2SbZq
w40jh2zmklHyxsZiD2y2MB/yfRI6pgQcloL89/ZEYgfpN4FD7jCakbWlZ/FS3R4vU/2jEGKBxcTA
tiXOcEQdSY55TjukITuofl3TiYUGwh/+IosPPu5AxhkO08SiPCG3zif4Z1zPUEAk+7gI+EQeqlOS
yGHwlev+SoL5/ptkdcNufMsALGM3LbVBcSuJMZs1QR2CL5mMCCFCDdhqdM5VwhZhX7NC1BYGM0Be
iR58HT0svCOEB11J34IJPpUzUprA6qFDy+9ojy/r0NIbJ5+uySfKm5y9Pxrrf/CCpB2mEig2KZxx
Z6KQUv+44y45fbirJ+7si+tQ7MkBM9RTf+dDj74myxHV8avJGC1tyIoZl6xlZ3rXCEHhsKRklJ5k
Hex+moTmc7aZXH6qLZy9DTSRO2HVXqLyzM86p8xoDzQn1PjzVeW+XjK7pe5D2Kvxk9T6YhjZnQjP
h+P7fyBK9eqxpE+dLPRw6gSOwQj337Asw5A4XWuacgtc6o8seFdmXMiJLNhnmzI9REeqXS118D3u
yDOAzYpqgW25Vopsu8gmTBtshshwVb0os+NaYjsfDr1S4C6XZ+5uDI3ViMRj5pNRzT7EIc+IfoBW
5sEGrlht4GimmMg9F94ggFp/VicJ1XQESmb6w1OZ+UEME357C1ys4YJ/f5y374D260XiOYvIf9+K
E/2ofslzlbgvYeSQvWOQ7xJu32dgnstGR0sV56llNg5oQFHCn6YkYOL/Eial9QXZA8j9b3iscRRF
JtXtYe4RKcf2wNC/tTypwgSuM7pW3AmJ1+viPWLA62u5gz72KM5sVfmy2ry3cG5W51EH5LQo7OP1
yVlGCN3mfIrVEauqb/SQFxjtBp7Zz8psq092hGn2u79T+luLV/XERGP9HbNYBASRcqije8qsq6tX
YjdA6YrqgAYFu3uDmbJlrrTmQJyNm2tSQJ4Re/s39cHpJwScTbpGtwrz35xVoTN87uK0pv/Wrq4S
h4o4n7EL5HyG86yQpQpoSLejV3sqD3T94RqA+OSW1yufYCTN69RR6GAJgvZgY4v9sr/Ew4dmMgpS
oCYiZxqRX06Y5hNNGFS0QM0wNDYO6iwITDStvmf5vC3l1TWgdRn39rS/gHlSDf81uIYkQqJxKkcc
CqOymEMTT/vO4rMjffAI7QDdnjac3gsaqlZkxt0OXuTkzuwcGaCshglHFdrotbhyQC3itTMa9p/e
+ImSh+65vCfSY32ac8dOebkj6B+4VwxeCtivsx2uH219XQuEEZ/LQARPGjIuuf7+vR5fthfiLbkW
tBu3Yg1Lq0MyBRuEbg4jbWTx9ozVGoVwlZnOEWZXKLmydlPDEgdL6IrhBJXUKOxCHAe3XvbCYaCK
+xXyA3nRpgQSbYoknKGQaOJGXWYJ6eCSFnyAFLn8hj7EhTdD/sO2U+ZRTRDTyM0uDwr4n0UQr1U2
wD6diC/1xJCXM09AWZoGGO7XeujH+TxfV63fqhMMNPLBVib0RcXNT37wW9Lu2Rdo4IgzxgTwK71P
qq4Zamz9aFXGmZkfcN9ibPFtDqg9ee1G1gMMPRBsp30qGh/r1Cy2ow4IBFszm63UKVxDK/FXR3Qq
7tjDY60MXXiM7SfbrsEACjHkEROSGqpy23BTUZjQC6A1ya6qmjLKQuT3aTTvcoNO5Ru0wmklZE1B
b//BAeiTx4nVme+n6booMB7AOr80LQr6RGl/27s6IbeA2p0OHrSB0hKkFLNcRIwcLYlkDBlDZ2dw
+khiDisyVIwuw2/wtD98uB86eLAXhuLq/BZ/mpcTCcl49Js0yO9VcX9cMuop0hb4TFoizUX8TFEI
rTJkdPen+wWhfkecY0QFIh12rMxYBldZPbqvbxW4lCL08kUsV61iNKyXFicBifMibiisYGURo5L0
irpk91OJCcF0//bRnFPQhc20DTdkFyiNChQGt9nQRMl09aMhlMxIG8AMQkKcvii/e9vIdgTj3vie
BLFKMqGUfnXmjG45fTJ/IuH4nTjzc2usNl89QdeT2+sWA64yJdvDcpOvEqfgyPPvO36+SSeXVUrZ
beW7AnB4QMzL9L3ox80Dego/RzICZF4LW3U4sqn/6y+uFJysi+y9HwDM5JFqiNmOhRmBstN4yD3G
bVUveuAjKrKYaLn82pdF+EEvjS9lGwTxPzG6UOvg3+U2Tdl2PoyUnZuRE3w6tv+v36q3Qq4BQqOy
zMJ3DP3wMRUuqB33BZZlWQopXbhVBUx2uL91wfkeKN3DCvuJqrufira52DHIApPlNSFnKmXWymPQ
C4ZbgIAZTQolKirO3AQiSXbAIMgsyqADYrKktqjMMSIFfS+2PL/+hwMldtydtcaBXYvXXZYpZyiC
gtsYXh3mipV7R76vGPpORdPE6MJ1bUt17C/J+XBUmICfnPv0FvdmXUfrYH1E9Nw2bKxj1rroCFwK
XPMACcPp3F1FeiCsMaa6r5inLK/EFCNoamlzzCQfea+0y17w7/NPqqqvkuvB+kNhesJXd3qGWs7L
oupJJ0m9AgmjCw8YM/EfxIOjJEEJVDBgoZdRNzw6h+dn4S5lVUUjytBz6f2f3OEZaEfOp+X3xhi2
dsUY+QRX7UrrOsCOHycAAuO298CgfLT+xclugRRBgf5rRG72ebqlwPL2O4y3+sy4eL4KBrTlKqhA
/zQczveyS43HeWrIBMNvEyUn4FODw1uRoojVErVa+dQaGn5pCDeCh7NqrMPKPiLFUkZRoh4fbq7G
g19G1aY1bSNjvj/d2Gvt5TmhwI02q0sgpiMHIl7gfRPmgg64mSJgBLtdZXcuFucPLnXXWIDI5cRZ
JKE/eo/C5mG6bBOIQx/a3dXKFS2GxLhZoApQzRVxD4jDDGN2gQv/jw5oQeIninxtFj5C1ogfnV30
Nuof2uQq0WC4EPBXedMLOFZRCcxNb+XpT0JDWFE/Nfwz8/pll/D7nR174PUbbUkPCG6OTimA0xMk
39CdmhNxGpoWqSvUiQrLApJAsjALjQLpucL7dH9BQd7m1OWI3BeL+9peMVnXT73QNXNVVVe5lYOL
lhIhONs1lIzGmhbk4KPmQlBROoDWbKbZgiQH5b2Wtq/PIVxSjrzTXlxiPQgsO0VFXrPwbmQiCHE/
r+lT7lTwI6JCmo0vhh7iPZXFwSnNv+1oTWUynmPjWJr+OXmVL1fSNDShyombJdDIcXWK+rvTT5PS
6233gf5BxAsk7/h+PaqhL74ZpPoB7d+lYzN/RnJky7fHMfuFI+WWtL3tbQDPpm42uXPrHZVhTgga
7rj6QT871jWbp1ybOtCO2/KHETJ4wV/3AyQ/qVOXd4rL30Q0NxnJRmEeqXG5n74iny20S1c22fq7
pXhcYJJw+mpcw2sSfv6Wlmdj6hL9y4NA6uv4tHSkMHZZ12+vaGOcVysR2lDwYGFX0phZphNRLz+C
Ku+XhjKnFIIoIrnsDxbTm4TM2FeMni6snW49BzCNwKvkqWo3ZSq09qrOaTisJsgkTiDe7r7//JOR
haw0WWSN3w3fif3nuauaxnuVicHBHfQyTZ5WUiS7aIA/kfzQ9gMaVIFZ+7ZcbpfigC6geXF9lSdi
hP7mjoqQsCtqctOPmn5JbKjefYCBkPrqw3UIOwPrLM7DAahUHEM4859Zh6Xj/2cenY1cvE6qrbac
+3oL6h5j4Fv85WFGKrVR4s0jw1sLhDMtbaRItZ1bHCAwyMyxI0qk1LxQUkcJF1+9aVzlcG5Jzl2o
99xnBmshCIKetncWfq5/KZdIWbE4SfRdZjmY0keuIi1Cy3aQoPrly8Tf/x5WTBfVib/UDrH3mRix
nJNrvn7xJ6kTJ2lFFhNxg4h+uD8eOqNQrRNwv4ACdx8NgZ2twfQOseDCOCNjWTSMZwWmqjpfmqBK
ADuLo1En30fxfJA44tW6jqjR7Gao+BaVigmw6yBV9MhMbhlv7H9Dn/mrVm1TZD5o2Wdb+jgAq1tM
Ge1QopPhPKwtnBMfEfu5fyRKjLrlqa1LTIj09zlAC1wIEyleaBvbeIuuw5KBBJBs6LPTw/f7CZ5H
ore54FQrwmAbbFfFjfQ8KMHm2uXy5oGnXzNBLV88ZRwGRiVnDuCBoRDk0IMuQk0j5jxjvGFsMwa3
+pi2kGxuhc/WRIJx+ny/bdW+gSZclrjxd5mHNrgGJiSX60z68oCCiH8yey1Du+wlHLLgZCAWRM1j
1qUHtQF4KqVEiOXkBuEtMb7TVgjeBBpSLqLrqawInngZN7kSY26MFwOyAc4YN8AmkDqEZwJK59Iu
4KGEfhsxUneLehQA1PT3taNgCZCCXAZp9+gS6sd/EkcQO11KALMjeSCqZs3EKiv0nszROfFQp3HS
bVFwIUMKsVJiebcruedjU6xcCGj5MVuzmf0y+7h7LCtD+Z1FRtVsqwppgxAmRXAImL5Q6qzlLhYn
CJ59QLDxIf3yAJh93M0OcMsH6rBn7N7Ad+QrA3IcYzwLxLwSF0otgj2EKzilC5b1RTMbgPnzePbO
NhNaiZgMNG7+GM3aHHgK0W4I3zX2cNJTDlb8h7mLCYj7P0lLdiMBYjQ5ogd8QW9ZY3JchrVl0Amj
lhhmEe2cVgwVLMnWUWtloLCNVt7TcAMxEm9g3EkozJJ6eDO8gXLUCHnzWkegQR6gQlmpNqvqu8AW
NpAJzDBBSLMIAp/rEi19e2hWieyv0r87MBSLMWh82PP3bd5aIE+IlFg9Lk+Y/BtiYezo0Vy/oIj4
wraodoGJ+a/r5kvAp0eBU47pg3jjqZkaF6Wxl7M95HQF/v2Zm1dUerIrP0efq0vlCdqz9kRrJ8rC
sA9MSQ6wFDBGpgJD3VpE2QiF8NiFqa2vanz0jYg9rbf0GEfeCIt+hf/gACRxHll7Y3bJ8xkGIzNv
zgpoNokZddx1k0N/Wg10GONuF7YIJQ/KvEBzKl0eGM+cgLMDW2Z2aQgxJz820WjieMnb/rY+Yzef
vnAiPg2vfwPoSfZ5SQ3UNh6h+sULJPA5MvunnFiMVKWKH/mEJlXCqaqs/1apIyMXQXzKgOz1dOPH
pTyXOucwjHPHZPmH63Tya703Ui0nHolm85uYrwZGlFBqRKN+STRd9goMfSFVvF13C3E7/Xn+3fF3
CutLgnzofoeQvN7103g4uhioYN/5RPLUkNWljDFrnoMtYrsyGV12zpNFcvN3RneBmHaaYwFRljes
6Sf0YukIj4U2leKfUj3BnUztlxY7oaRPCu1ImnBI9nC64ocV3m1/GwEJztX2jzOT/F3RcFOiY6Tz
IIZjuztDOXitWOsRSEpIwNObXUejLbKI2MoUpjdCdRB2Dy0KYpG6FagICXZdXEOcUrByXGCFTC4A
FadVMgahnIbe023P2T54NQAv2acOuUksaNBpIVKzDjU2XvSw0a+s1NnG9A+C89FklXv8RnygK87/
LxU68oJQX30iEhNji6dyyY268p4kfhoFOT/PP9f7a75I1GbMSxF6P48GjrYRYiI59zQrJs9W073m
AtX0E3EebNwL2EnbQXrwy+Ybv8UD9qiPt4Lgim2tpjSF3j+RkWTmA7+iEWjF6vtj/XqLn84WsX0w
Cp8cDpxtYyI9isJQtSZSRTkkguIIux6+4lDZrTstgOx1mzHSBTzNC9UPWrSB+BMG2E742dUexJ10
yqATEVLWpqPWf9tXwWze4SD5Q/04WVIzvatE2AbIPOAHZ77pv7Xhq8fhYXR5HVyl6v6RgDQEd40I
MfyExNsZvwP3unOvQb5/qSTOfcFH61TxT9EUqX4VNzIFlpp89DF3Gpqg09l1z5dUSevVH9zH7Hsy
QQx2fxEGb+j+8liYunGPZ0YX1tvRJ+2jP9aD3BqRUy4Iyw3oraG6lhXeM1h9HGirox8zUTxuEcGU
iiZYNLwMI80A8kKEbqI8KphUij1iQXrb7SlAmmGTYU0X8BtHiNtVqOWcE5TFvTkAMj20o4y2CQOR
W/08BKPSMAOoQmf6+FSb9xEJ7STEVyEOLzqLS1f4DcN9V6rlgK5Q503XReHvGJfh9dg5whDrSc5/
oO3iApENLgz7RZGjZuNbwhO3fKSaPhGRiTkRS2B9poOobYbcCcK0u40RuCAm7bFMu9CgEnOhd5Wg
nYQwnWj3O9c2R1bEUV7IvHEatzeZaIyitO5w7a8d24q+cBDhvDZTdrVHaPFdUxjmkAHLPPCSlZ5t
8BGwtyYmuPCn0vgFkO5qUAm6dnwbgst9ESslfFYyv8z52J1zQb8VZx7xAqelbq3uhYo3NmYeZTKl
CqUJqk/0EYGqlwcQtrksnvdo1wBBET8wppyJULEtf1OBnlHMcfdz6Ea0iUhXJY0wBWgQ7fYGN0vU
/Upg0Hb/Il6QREs0yyqKw6maxCdtojSCHVrAeCm8keKAtmR5xRo8teHNzN6Kei4ONFiBSTQXIq6h
tqoepIkj6cFIBw2YvN70UXTDMP6kLebPhCf1+0tQbVpN18sqbHOS3XkfoILhz8r1nd/bdA3oN2x+
8msENScnO9yoOiD5troMO9SG4G2fpyrFDZxN9sDfMz0T+hfYq7S0anIrT0kzAIrrVAjSS8pr2dZT
g0aMxqaifkB+xKpcpKP9Jhw9NNVvAkB4DQ+B9GCaQqEvBsvbt4aE+2R6pIP8t1itVJQjxhF3L+ot
p3/GtP0V5oBprWtdUb0iF1dfRKeGZ34ecbixiPGw1PEoZD/4L/Nl5OxHEYkL3Ni220+hOkrohrwp
ZQXn0bBa/vxYOPWyHylO3DLvzr1iS76sUwhM2a8Ki9yxCSMD6d74gBt0kmqccsQdufgCNCDeE9Xz
OxwYSwxNxMEiHzV9OWIQj4iqPHPir8We3S5kNCDRDjtnV7+JKiMx3kbE02nwkNGSJ1OzEerVczn+
sOsFudX/WT9Q547sckdA6kftnyH43WlifJgE9V3CWnlSQqMdWTEL26GKIcOBAbGlSGZQVlDr2NxD
GVHijRksY4rR4/rWLwGSSnO9G6RhG9+ls7Jsbp/84ti4UwxB9MVMRcLrfMJXwtteMSkDiLq83Ltw
8jobNuZDlGzkLVWlFusDfyrWjWJ2tSzoqeVf3pea7SA+1wmsXWGTcJfppXrt3UJ+9sN6mP+7+ECt
iEEhho+mI+DlveSKFAIWKxrHHmT8uPQrtAKvhvBuNoUzarzss7v51jpA0kXW2sIcIGJKsRvcjaTs
e4etWB3MJOc7VWAIH66kdSxlR60jmGFDwOcWg/HzV5cDrt6NpprvGa2tTqLvJ+L0YvjuF4mBoQcG
++VbPLXCci31+eoPfBpWDHLsYgvUr4YLeT9J06U1lDIY34LFFpI8PRySbZv1CY2Cibe/WtHC5EWn
m1q/wQkg/5X7guCKl3izAmB0OfjBs093SxL0mbNPhq5LUfFYZDOKg0DD6gxHEv5rmBHOGtEXNXSg
OSOPqA+I9arq+dW2SSw5zqH1D5BdOcvhgm3MNjcdsOzPutdgmkeUThX1Cfn0DXn4v47pToZs8sae
EVWDzVKFg6AbSbERkLxJNYjtbq0O7Bb9n6Bu7aiZPSI/lgm0dfZaV4TL5/6g0yexZjR9pYzXqlFF
CvEGeY0AsCV6h5xJmtb/A00DtaNp3/OTr9nuoKEBN6Ag90uyQgLFF9hSkMbP3wUVuz6of6UhjA+D
dOo6QoiFju936hSdIAnMIZWMUtU+AUFFzcEkKczUDdwImIyWKRsUU8eSGj7lkT5f92KBvSWVjQOY
mtsBCheF6PRBWojeP+MmiDsxEWdv2BFUWVDB3p8MGAJ7QOdG31h2QwRbdoGJRf+KNTOUiPPu2YCW
+0oSrls6LmrQfa+CEDhRDll7R/C2gd5SM9nlBrh4O1JV0z98lhhgJtihi+pKV/NVGTz9w+0Pe+CB
vZziILludBVxLt4j/YDIY7qePY0ktFMWVritsHmdw5dPbwmvnAerPhloC2X2YDYcFvRiQ2uidjz7
WMqAerr76WGdW/ZfJ3I4gKzTLNoRJTe3TF1+Q2USXPVhteUz1cMYKXVqR8dTATMApHLPr8Vc7/00
Z0SHlMTzkFDoTVh05WraghUIhP5HhCT04d/B18YU1UV8aHtKpXPOntQ6FDL5Nnc+O7PUBC0ZbZ8L
y5fF3Rvbr1LFxnkpPxfw4x4V9AX84p6w5N/zY0BVkhViK2nIF/w0sdhV4Cedzw3u1ngD9+DKJjwO
FyDDzhaSnFMAesFmmIh3QWqwr4S8yLM10JXSYpwYEx2WgZLqrhJbEIDNhyx/59HLv4bG3GoeTvnr
3AQQ8vDNUlNo0hrzx6J/mKcC+xKJWZOUeUkn8J+W6qEXKZ9SiPcy0YO4Ub/Ev1K1dSD8qo6KtGdq
UU0YgsAjyOgj6wNGMZdwe/6Ha8r+Snpmgk34vNOeoFBU3KbR6D+8TIWJiQ/UzDMWqydybKSEVR+A
TBGdRHP7an7OpRZlvardB94cvnDAH41c6WyUEItRa3Alj5EF9hyowu24FW531DfXoW9qvfk0cBSA
Myo0YHOEDEIglmwrHQSF3+7LIN1a7IYd/miMmFkOJSO8ijCko02BEgQibGHsfehUJ/zy1v9GPaOM
UTHKKiEgHY5Q+OWybdDocARyYxyneTcWEbV7SteFXuIDtN5VVU5tgVz5Z5wZwOqp2kGAXhm1L3Pt
SxzxwKwWmA9CbWyhwUpml2l1nPqbk7rEbl/vIrkTnNysoktk+7UITrPE9unRcOJxNNEbAYqiuejf
iZEmUIiNjEO7dW4UgNMFoh8Pmsi1LGXR+r7xwERiIEzYFCRg6B0jM2iS9qtyJkxeObCruuloav9B
ydBxH0zEWCp8x0XjBdf7pQzII3RgqHAx1Dbzv86N3rRYs4mEA1R+6rEzLHRVbCR10bzB1n8JwN5/
+IVxXji/SLQLbkp8eUBn+pXp5bMrrYDhYN4nWeimPs3+GM85etR+4WJQ6oHVubno7hZR+FKKdMNC
gFUcf9owHDwWEfF1L54sgyLDptBdZxiCEGWmva/tPaEoPF/xfyFM8z0bF8ztxWadyk/XFnpMYGZD
UEgKoh74WMah8eF6cdH0w1D9Zsw4fq2vNBFn/TORgqzROL88kkBDhHoiLkhqEiUxHYe23gP4PuUL
AXD7vCQ8hlBjgUq61403WphLmWFJZTB+OOTAY3Id7xW1pMPEAvfR7WLyKorldIMQHSMOzv/AlLli
uNz26NLFJNz3Dq+reMop9KXXDwkrpC9BCeEUSDhcQg+R6I3syFn4u2bxwIdzl1tpGtT6qycvOSHM
vsnKIo6J1VriF7o5ZvfW48uKgM/ePUJ2RNNmhiKd0p9Ku/Sg94nZm4Ri1iOQ4gnvpR5hNdWDTuGB
rVPt+5mQ9Q6IAc6CnshFV04dJgY9ZjzcuG3U+/FRtSGpL24Fq/aAywagGxHQdSsbaxw2PyxB29X9
4vfpuEI9nQNG4V5g82OFAFynZg7E1XhKe5mm+axG6mc8nCFZ29oAcSf06jy3TJWAXSBMeWLCpU2Y
PbAxrhHoI/fDykjCHzhYl9HaGuUzS2NTXI09wq3TbQz4YkbQxXJJJs3azbhtNtO+Hv8D1UnPyfhd
jDcxV8xhK3bvp89hqmA+jALPALPCFyUFlxF+Z1MW9KI+Ct7iYHGrOPPEltX7LzD7/42yRPZCI90P
dsh2FzE2zr4xLMDq0Q10FF5X1Pld4BvCDE0XoZwhsiE/yQ5Gb9cJJqFsOYW8sb9FPE0mu/2NexrY
oMVxz4H2/zXTBs7qBEmyn6sN3v7oIlX9gVOwr9iHftz7iQcSCUjlbf457BgDRFS5SpZaejYzG4lf
epcjddbGSmeGvpAdJHr1ARB3jz0lq9pI74UNZNNdd+TXsIAESZ0WoCaQto0A9/gqWIgl4MHJgt0f
NZEZq8t36/NFB9Ec9WxX54ZmzGNmjFAbctJEg/NoJa9C8Vh7OgHgff8pWASioa6Yj/AiJX62YMlZ
T6Nlt/pjzQxZwH+gbP/xLH4Z3qo3rJlLRY9qAdWr1tRFrFeYdaix3x7m7uV9fInkT+58M4LdnkXL
JW5Ahkg52HBtM1mLDv0+AcuOWw5auPgZT6/etQwZUfcgbL00a9dXGgKx48PevUM9CXn8WmbesS2I
HW+IU8droRanrNmj8OTjDH0T8xOieB+l0q7HxrIWeQ/5lEkt6SDTKUUpMtYy8rzIh18JEHmZwRU1
ZMNGKTgF+KxvpWmvjhzLa6YqDrumINOfUsmJqArWo6WbcRuF1iwRbUAwRhW/fVVy854s8COVZFoD
5BjBwh6YWDAQQPjjXQxNZkdO455GxG5t6BkTbXrJjiu9Kk7VxBX5VVuabON5QfnUnOVvwd2r+uiX
okqQm3mQr5LltpNk5hp7+qmIBYBc4MrOXda21N/mq74CTyuOlqTtD5hVaC9nFUvEV0iYtSpKoBgy
x8Lc6MgxEUUhW+TlAy8GLd4isIrsSuXbAI3ayTv8jWlQIDMn8AXcQjunIOQJOqKh1TG2ybqoO0fw
2f0Dheca7SB2f8UuOu2l+1/dxZkUTzlGMVPdVgLz2aB+RnzSM6lqO+OUuQCUl8swEtBH1TjpSFEW
xRvLiLW/AS/tjkC0Wn0l9kA6dY6r9R7Ec3JPJ6EsP+7D3X8/p3Y+xEdMl9V/zDEghsxtyutlLtuN
ztD3RPk/MbTl44x0r9gnAy/tZrWIqY2DJ6R35+nUMpCXPHpI57pEy78ig/FUYqFbWsYgRFPBWMN7
1bdGTqXewflSsOxnq99fdU7Bqe6zMFGi8GWusSx0jwQN/ikw4p7ntxrk0+WIiJGl+cKEj0AzBse5
YCS6TBzHwEL45IysgMjSGyTlHwe0WWsQ25iNZm3c92mv+sUZrKnfBRWz9gAhlPLqLVdGzfrG1v10
TqNO9kDN3jhfkuLQas5PJF5I8ho8Po/fJ6GMDahM6ezw+ddHrQ/vU65kIwGa4J5VM7op7fK9ifB7
j2rvt0GCWEFpHS5jx+jbiw0EDQaWOUoJX+KHtZxd4V3vQTGQdk5fmt0bncOVHyHKNxWK1oUHOWTA
ZpfdtoVDbovxFfDjU8DlJNl0y7beq/vVKLrLKb1z50brlFHO7xa/hjkHhqnnbdz8V5fzugT1PiQg
2W7kVPjMMVJ+J7lIIH984Cn1fyhK9dp6BQrGxkwKDU6B6PPGCB/GfAS2FxHjmPJ7SpRLK64WQw4g
Tx/fFFDuG7xfX13rQECuHquMZMBerZXuoEHAeKucBax5xZwxUqb3VTCbjXudSr/ZcnDUPLsSHuVG
wYf4gvstKCPuFYsWfYszyiMs1nqirAsLh4pxsRuG8iHftCLVdZlantNeGfti573TN8BHqYEoJcNt
dQMWLDxSIvdIWj+QMHVH5mRn+6Z0HqB6ScoExkZXZC3SRIK1IK3EAEy7/btqAI2WkIEQaM7ThUmy
HBHoai0SJYvUbz+COdyQ49lni78M1TUjv7IyN+hi2IVXPbKQ/QvwPZEf60tqadkrKSs/a/uvel4s
1SMJNxgxwpgdBHPWPMzrMsng5Uf4wEUjF081TPX3riJeb5kaXKjF0IAc93crH4YkTTYag/K0jexL
PMBZHSu4PYfqw61K6gqDnwHIgKBY625BeBC0WvsayFw/ZIKf4NbIfO6aK3eQDNVRSGoYoiEpaBQ6
aOxP4GLIMLc3zWsGp12GLTjhJoz8IjSokpUGz2EQxWbiygsUaz2CF2vYLnOr1WY6hjOj446995YJ
fCYzqKCEdKGVlH5etSf349FDJKtOeMEc1N2jZGQK0T8/8RltXA6HhEOforTpbagzHiR1gsRnjo0Y
iXMo/1i/vkO8A5ufaMMtA3ysrp5q3dVaK9EhYqw/AZpPZmhAHUsIWocNxFC9UGrti2t5prONQtte
6MW0G0NV18CsaxIUVMHd7WlQN2Mcawm48+SVlc7meoqWpQT5Di9vhjKVk7BbvzwbCQ2jEvMlDSA+
BlfE5/LZRFcKOaSe4/xQoDzXGdcxsSialSQe+HLhSGuWmhl37vtGnGNLvopnesn5DNUUNoyRjkFc
IO6lDtoslnztSQruBYu34h6SDUCqaxwkWxvSNMeFNP0NeB3KZ/h/zio0AL1PSdk5A6MNg5T/MWDG
LZauL8hCw+f7UErEqWcgYl3tgIky2tnWLVaGjWFBVtDw14Gr0zK8FDg5uS07My4RxqvkFOQNlBdV
wXcGMnzIEAKXj+Pfs48pIFOGmbMnjQSJCWoq8wNqChdUF30dOGOnCjbC3ahlYRFfjPM5Jif9NWPy
ZA4QafaQEzV3VKcl8g+IcDaJNE5KlcFT5zSh2GrN9er/1g8TRavdcgnFq+wXrLl4pQEQzET1eVgg
OAZIotu7y2jpviPeGZ5AfPpXnnlxnsA4Bh+4TYYWd/bq0vH0nnFz+kgalbxR9BcTml1vnnebOitl
v9vKSQx3hTDg4YzI5Sm4IQUw16iyJ6jFUTU9/e3dQvYKhxTZKLJUfxVa10Y1zXeQ6sz0KkO72cpJ
UyevVJo4BGgIeola5eGjtEYaQJCbyvVt4ioQpv59bpfI7GXNaYF1U5JLR5BpmuePd9VC4l3Hk6K1
1lOrIOS/oycToLDnVe9yFme9y3M+TNFyEk0QG3U5TWG1ScGrmsjwW8uDrvZ+zh1o/CoEjrUBuJ6U
ONYXxCyhDEKjiI2ZM65MixE1C8rDow5re9elMJ10ph3IjjxEkQR90pmmrXuDF/+RzsUGmcEEN0vr
O2vCuyw8KClgaMlgKmvge0S0tP27FQ1P8T1sKIWoVFkufRtZGdxlxCU+75tnhRcvma9NgnsQ2k9x
42ULuX6KmTSJwv8mZlCW5THcOQynD04pqbXH9K9BG3Rd3ft/OmJM8spqPJGbXPf+DU9z1XtsOAxd
Ul8VmZTeF+pzJPCbW8lgWqmqMGFcXGmj12mZN5U6p+drdj0mWM5a/EGUafM5igOezRLzZL6hZyoO
S8v6fj42AbEs35BqXMmmLHOlJXUBm7SWBDVLI8kwxjmSxS2SWOR8LwcbCRiVzgXTC/feB4AN1MvF
EaUq4Q5zXBiaeg1Fv8ZieWo3eOkmF8j1sWGPpTdRrJx/VFSyLDSXL+SbBxjOD/4QR9kqSp7BMdiA
THhSzIi6qXhgzpT2Qua33qa5uTF0+58CktUWD0Jjw11hz6oxagy8USp23xjOuEdjR3opQ/jL7BK7
i7lKDvctDIu22PvIpndjPqIjZfxzvXUCTdv6/PAggu7rtQPw1O/yyzncVFpP6K+A8cXngNqayP/Q
9ocXP75LkkGt6GkCR+K7btLD04Z0I2ccUyahNnv5aefxMpHuNkoNX2omhSJLn2h2Vr2/yMPm+AxD
PcTi0SAaIoB4N87gjfR3+SUBzn5wb94NAyX+YINdBP41WIN4FeVBJVr+TGFGaQ7ckmdG1YnW9vv/
hx7fn0ah8AfYeE03Ic/GRp76awT/5NySnMH2iCjw6oImcJ0Jj71TB6KiH+AdYaHsneDATev67eav
a3SAJ/Z6pl2QwViJYt8ja94Dq4f4eUPSbrUO43LVKEUaqVX5X9IchYH3nz+OTdlL9THH4oah870n
j+Q6iCw0yovug7S98tIOHM+G0ZQI2ihwOHp3jUf1VkHZpYybANS1V4kQ5ORKYxAsILlE+hmwgrjk
tw/BsItQ71px3XhjV/AW61XUga5QKmJrEqVfKCRKvCa+nVAc18kVzc5sQgIF32HC6M/BXVkg5P5w
WizpmKN242CI0A+TdV75MSQPFYhuLGsG7maANVaG18InRCN946ZwEahl31MzulgJS7+vEmEtGzG3
/3jC7mz69wgT3+RerjKqIqugUR9N9dUyxx7zPt942OfgDj+Np/8KIS6A1KkJ9C01ZmzlYm3BC1K9
SUJOQfIu9dLRmjk3icgI2ZtFpYzVBa6C59fPYgSrEUyCsChuXl1mm4GBUqgTH2e+lAsvH6ND6SXd
YYXcYuVCidiYSlVfm5bMj8oPNy3kEH+CcsBHfgqLVN5myHYFlIdxLoXI3F6jcEGMKnNpzz5pJZFN
F4kpRbNZW1jc6PcgTgslTzW5KzOGGlYlxL093b7cxhAfCTuuvVrawdGT7C/hxwMFDYJGj7XXtCZD
AapFUKrlQ2xrjrVBZfyhY40d+hnP063wY7sOv3yYW7dQO+BfpHN0h+wOhx/labC1Y+jKduUEzhGM
2F8Ejppe9BOvBfujsY3W63P5mSwm2Epir+mBBlfVdh4gMiODpdirDXUjdo6XmpCBaEKPI8Db0s58
G3YNblv+T/uz7WYeEOHS7vD9r4QDYt7LIyu3ry7d891p9Fd+RuNECtYdAa+297U7WKWcZgJFbuNx
mX/r4XlO7r4KCmsowGajfnnbrZCtZ6j0nm2mYo1z0qUCOLQSe0kTH9Oug4ySi9CDRTxWOFlkyHoC
NLq1CE0jOnSw8CIvk0HyOluZmcM4QxiPByX2YkY066MbrONQM9Ifwp17Qgup8DJ9G28gnHozHH+G
3wHV3I3zahZ44LTDGSr2xlGg2N9KC8PiKblUvx1bE9kNqtId3/N+zUaWtCDaa+a6LsqRv/LIaD5j
svwciFvUsPwgY/DxJeRsDd8y6upHqH2qx+V3iKPGy9lohhP7FjrLTWAdnIXenGjjxurfghUUknna
Y15hyeUuXNfDB2n5nKq5yKnMyYE6YkVlCEO4V2BESE2XP6u5u36RXrDVbHNvHWPW9PBdvC5CMgKe
SozIn9wkVfXlGpnldOcrr+lyyW7itPSVb4xOYvHVRlpQbayitaTdN8MB1GxQBSqm1YehBNuUPpjD
D4+K+8JCW3QvIxIzVtD9syEWWn/NYZuL6xKvF0r4po4WR0qy12y25t/SlZ1aCD5Lkow/QaHB5ost
LmXyH5ZZObgPnHtgz3hzEs1iAPIH6V0ZQJSapKpZ4OoDfY884eunHCzKRYoExB+f+U/tWzgz9ryq
52ace0o2J/Bxiqr8X6XWhva6kkXKnjKThxBo+SisOUfuTOPFbEo92W0UJW+fpAHVYOf1ELl/PkoX
IItyCOgWcwkhBQEXbEJfcr/UFZnbLLRHVn4u7KxsWP+wURz6bJe6W44YBbA9Id6NG7ZcFt0JPvNh
3X9iB2q3fG3OUZzis9DJu2MDcz+nH+uKaOS/vuqm0XvyE7klZolSO7e4JCApQYIh7lsTKDNU1j24
P89Ssz5V3NUkgUbHdtVn3FhZha9H+qiG9H/eRwoWdoHw7Ej7uZKuFZHmarBGEEfccYvwawX1IdhN
AzjNB1755FxjxoB6FXZIsAUrWBRgTziPumedNy1U7y9+Dyp28RDy7HJpBKFNA6eDHO2bfXCfYD/k
+dTOTh/F0fYA6yGSo55QRb13JyV3d+ZUQPA5Xw0Api46z9ukFGgWWxpuE8nmfpnG+ZzQhfralgcB
1xcIJ+o7PVkJH92oOGbMMsW1RN3ZHkX1OqnORU6yDzwlObxiKpCQX5NqAWWmWM1Gp3klgV2NHf9E
U55Dozp+pLhUJMm4oNb+0f9HAjddBew2hYApbcq/TGhYLyR8T6qLrPQVKzR1yxq4yFG7kdZvYsrS
Fq5xRNGmQFY9Nmup5bDUqy/QoBSeFklGIAv3vlGaJsIBCAqPzOyz+4CgS98UtdDjUgflREh+laei
nL1N/Xr8iorqvPYYuRgFU7U9Sw9hDTwzxkUdeUO5MrXVWgY9qfuSVCU8my/9aZdXEfmwydF3AVr2
cKsNlqxPh1TFfZ6vD5KYcY81oEfQwZkke0lHG/fqcH/HwEBpuM35vofuArneo/yXOw54ZZgFsBcD
7+3r9+X3G9RGpddKwDZf/zxvDlMTXAmVSKF9QzPxMY9CS1bcP4Gpzpfy4e07AUgbYdIbLr2kcZZF
DSODtXHIKBcq4zwxEKXXFEmiPT61y9DmHrlh1+ubK1sa/BSQdaK+uoMXfvG4HYDwFvMO5/Uii9t4
GJO6G/vHAmT8htwCaxsyALiSPJXGnZd260ES3PBLFP/3C9MH7vCP0twS6vObGyHIEtz/cgA2i0rT
IuN44LL2sc5+u7I0Mb8nQ6bvPBEZaE8RPoUQGVtXp1yjyqIc/VrSOsrwIJQJ+PLVjP/YZpdlYy+E
P4EqW7DjBXDazhwetoH/H5ITACn4PmQ16DqxI5t68k7BkD48ac+pLQCVUc3PBZAJhcg0WIpRx6Ua
cjwtp9LrK12i1yXCcSuYFYA6LVa8in9rWs5DNYher54X+wok2oMTXDNy/rngQQfUoYcB+2EKLPiQ
CMmoJLWhFnyJbWDXTn4/fu9bTyuHZV/arBdu0RirjACOJ3AFVaDq/E+A9hySfaB2BAuhPc6PzL4W
lTq8Wfbt6i/dR0SelcTxkdrf/JYgcbfxtBUeoutootV2aHbFQ2XxTyYqwEFscSVdHMLPyPrAsNpr
zY/cnRil+2OXnRey4nM5q/HSg/I7xQxONSXkZlnpKXa7DDtYw0ojrk1+gtGUuZmpCZd6PFcm+KrD
PhoALS39PZYZnYCfk0VtWUfM84ZZr6AaCyCusbXJVgDfxSmbi6BZBzKF1D07QG7HBtXMV0np51RV
jfmJs1fdexNg1PtRakk6yh0byCA0bZ/HKORAl3xCYKrUEoRGOLmSyNsDx8BhvX757Uyk0j4EYha9
KMKCWa45NTslIr995GyYh1haGW9AFJiSiRLNmDl0ApKhMzcyeBj5rBVT6Vim+5nDfjtY0bqnCWs6
wXd76eSl4rircvPgZ+I0g19m4JMNRPd+IBw74RzTK8He9l2N7Io37UmW5dVxrj20BiizY4QL0Ezn
Txc5v1Cj7Tev3H2nTXufuDzehpTXO9Dqdv+unm8W3CyKpW/oyTqkYqGZb/kU3m5SEnaxcgIUNmtY
bcb25as47bDutVPy4slNGJk1PF3XKTt69Zop0S4iRzVe+/mXym4BFrkz5xym255zKvZeNtFcUwbD
Q4k0+ZmHl63+RcbAmcJZaks0Iw15on/gvTVizHfY+hMdE7dEOn33XXTNOLm4glr3oZwAhP1+5di3
fU4GC7gBESim4CtHl6LT9TvRpvgP3VZoAUYvkXpyxL2vW/5llboPB6l5Vyhyh2H+Klixhuf5ulY1
wTe6+OzhrNK1F6h1e53NgaQ7qIuTcAQUwW5jRn+3uvKHn106DVYCfjEIfu6ggmKhmSYEuI3dXwwz
TaT+ZUqduYH7McuOOPyB4+0npJcOWEFiqXQ9tkRLMruF2TEIz6w1aAdDFVUVPbnl/UqBMercmHHN
A3sIAooq7CixNLG65nqZR98pWa+PODeUJYFkmL3sL4GwNaHgp45EwnALMcl/BHLcoeVWPs5Dfi6H
04NuWgLpH9Dan2dJPiRdLwh+UsgB1rLykD9tzesZMXSEWwpTBkadiIxm3eJXSTYpxmJAL1K3N4ZH
heDKHT1EfWyN5+6gvmslqMgUP20Hm959kq9TBi469Zoi05bcrL38VZZTtUtIVmDUCOjHYFBZl9xA
1Oc74t0I0jjPuAuVlI2oPZqDKBlMwivXL7AxWmz35KUIrBlcgzxfweNSYiLaGqM4Y6GYGnIZIwfC
JGtrUZjo8D5+n2uU6eM9CVFgos14Vf1QU9RGrqGNkjGA4ul8wC3bqOn5hxElDy0zdqs7+i07pFAz
6j1TL/R4Cq7lV9VdrPmhVC1ZcMRx/AGEL7yh8VOII3ct1XH7dhcsn1Di4FEqTd6XvpP0+CqpF9Xz
nZNj+qyRx57x1prT4USmOgT20ghRzB1Lose3dTTi5Cgc+Y9xH7hsRFVXC9DE/4H5Dg4RMJ7t/jyI
xSHwLlwZiyge8sqkbpTsAPZy/mu7BfMi1zTWKTIvV1iXaQnBRz3PO+AwqhvJptUrG4Tsh6oNMGZJ
PEWDL2bJqU/sydcM4YfZiwi9u8+VQ4W2bh9+Uv9BA2yXD4ZT/F2bC5xnkuf3PerUzsSWQtrCiwH4
gnxP6IGDecXqBl8x3xxxnvIFvCOtxUmD/AHgQ/VcfPijyX2XewxAImn0ouiKmBKeIdDeUy75Csx9
CeFFVjABA2smc0ThDV8bbuI1U0LoiF/QoVY5a4wLgnPZr8hqAMLHwaK2SqCZysUbEAseUNAmImLB
Ky+1A/Re79sOb8QR2BMib/XRnShAUtLODoeYdvjPuhkyxc82Wjqi9rwBk+kAR3zxY5Ri+I4YUXHm
QK9QEYOxe1A9MZs3FSB1EOAfa1+Xf8RurqXMidzv1algCN1ZTf9g4fCiMMfgWiWTcEhqHutVrb11
TqT7r9hUFFPfTwSx0WxGRM4rmyUIzATYBRxLJDWHilxcXjHO708qV/V7GiCQVlTv2t3Vo8wIEUQU
eX4oiPQfmMY3UlrkLAoVR3pBWrZPzJ42TTHIUXhyk3r6sHXiOETgh+7yyRpLvW5IJgDpXb3iW//M
/xC4ctiqOGHKRQYhAf2Iky6rGf+wdAOLwYOribUMCOJOpdweMG9Azu2Fi3C55GTZ0MqicF2+ZsZT
ITKyQk2XOfVt/OGgHaIMV2PJRHUt7aJ8IKnurn4EqkIOHT1r6dk3OLz6sguFcNMvEnxcApbGFUda
4o9j/0krswxrefquqGwXUmuz9ROtDH/F8DoiBatcfyPVa8zxG1KXrc1TCIJ1OtdMTvrVli45nTDf
dkEzPWYHc+8uBq9uiCbKe3/jVp9cTZ1iBcv1HvzdW32HmPqQcjWXUXMS8K85HwDSfOSiOtsIGV/R
QBCThkgZfoylgFYDoWO6j3VXp3zjANSBprB+nc27VkBwEHCcuzOGOhJxeL28rNij02zWsOs5u5Hy
y3i4Rb3Srd/rLlwabH6upH8WlMLDQGaCITCU2rUFKncG0UDrsRDubh7QaDaumnbcJU2LzGITqjZ7
0QULXwwrKVO5RDhhm50NmeQ+JU7TPeo/s328TaSpUDsbUXfWtBA+eUQcId3Dv3CyqzcsnHjluV6z
jibM0I30UOKmJ3qb3JOYmIia7QbipweH86fPv0PneHHjGUYIRxd3xskIVrnAteOXu0XtAlaH3c1T
Zpp9TCnU95ug7Zqb+D3rQOIa0Xh3yRAZGxdTfdq60TnUjSUWlcpDpSeWNgo+1gIHfclA9C1BH6D4
ds2Kg+484CC8r5JUM3/ox/7iMIw/xgZbvFHl5fpdFALj7BZdeYK/ueNNpMQdCjxlL8P0NQ9yj+y3
8x/IZ/5YWSn6krP1hrq6za8ioqnAKy/rPUOVS58oCwVxdzlbMqqsaWYQFJWOOlUWSkdCSWh3UORa
bzC7FXiUdUUYpKpWzCxUgbWVgLRrChleBUXVp/x/brCK9xsMOEGunmvp0okPjx5SQFVtzqyjmcjw
3WToEaSPJNsLYrs32fKexPyQNInAsN/osC9iB0sBOpYszqaFWbGxuNSYLXaNPf/qE1/ZzG5ikpZB
Os2THOWHymEnWEWHKwpoZbxMe51fF9f1CPKJ1yDftACiImz0rpwfFxsOrpGC70VCJFZUlR5+mktG
gl0SvGi6KcYSMJmcqp1rVhOniS94HXPxRHlul5lUeaS+kAXMoL4CqnWcyVGRnCpyk6SUYdc75MI2
1KiGPLvITlaQswKbTKXK1yNG9UKTGXpkSu8ha+Nk2mLyHcLrEY9pU1nU4xVm8R/bG/nsk6/zzVlV
NTyQYLe+q0CEh34vF+HUKcdywihnodS0h1xbJLQzpxrptLc6xDiwPsXQeDBz2Cg+lycpe+f7W9ar
tbjAP4PxUF6wdlvY+6ri+aojr07Xe6hnRF4FUnuyLYXq8uAWd5B4uzC5wr7z1ap4fHl2EgU1BLcm
ukPunatrkUrLo6Y0DeErUofcOESMJi00sv5UMI1meha3VGK+dVetxtsRrTh8r2FSdJYdx3RTY0hZ
5DVaXTH6s2phDZrfGFC8A+JK//mHk2SgV+/y1OjTZYHyt4oscIjp6YM8nOHO8JfVcfvMg+Wg8zCz
Lt3yjNK9YT4DFsJroTkXYAox1cHyjS/Bg21R4vLyMngM+xp/SP3/vDuJW5T33YADxBsyJ6SkAjmj
JKnb5PpAYpKinC51Z50B7UAz9/P5REAPqkQY8AEnEm8fFi5WVU1R7wcuApWX+b/wy2WrHXWxGAK8
Wh9XVQdJhQ6h9xPWn+zizey5g7/GXMbmsKTWPzbDZk5RFp19QtEZAo/oElQ1yRVV4eqKZLNdHD24
C5sWnWI5FPnyT1WSxTX5CBD4LossUcDIoDhcA/OI7KeNfEfpMJzd9y32gchgnSOsc/VKx5W5wBk+
E7lUYZS7038dxevBg+f/xBZcjpr5Z4vCHCuAw6e086ZEpmGF2n11PnQg82mYr9D4MbN3DXl99lID
+CN5JPjCCGmgCd14PbA1+GfU/2rpr92skEqliEAVO1yGe3zET7MVfUDEtJaIhcrsw2YCoc0BNVBr
jVzVAT+nOFymHBKh8356EKDH4dObnC6jTiIqivZobHqaCqMNpoU10LcIYpUGngrCbp4CS6+yUlmp
ox2PO2Y9x8vR6lmZaeXZ8y2tDfssnXEJhU4PsQNqW0EIV1enuF0a+It1W0yKq61T7N+xWeKLAxj2
8k0UtCJN/Q0ON+lE4ZxeNyi6QJTCLdnK39jH1mhAqHJDravX+T+EmG1og0D0k3oC0hG9gWUoF/Fr
oY33FoH+0WkytTKe5vn0kcc55ApWHTtggGtv0aXlpVy+1VQiqOE8lnlq3veQniBOmni0CjQTosrO
654O03svahTbNJDyEaP5w4I4c1HUevYq8SFxFRexYT19cP1g/w7YeL7tj3nIeJWVlLhHr8Hj2EIO
7l0h7VWmzLu61jLJaNzJuTbXEWb+9FGWPpTr23PykWKPF5I2UGeCpczjGI2ZJS1k5bNahtxgscpI
PRsu/sch4DY1gaPynFMx9Iie5j3X2wEoEn7PLMJHFgb/E5gK29obszKU73+IXVZVnKdiVNSFnoGo
JkPITwtN6W3uPU2qquP3xWUPO6RO84PbW8G8XIwziEn70hq8pwu+iAF8Cy5GrH+AEnor3qKrPpUt
J8YTQVOAeq8zG5C6eqmDrmfAUxLyPFG3ZfMZ7iihLNS8L/MhuMAOfqyWbbUzW7jTm8mcMEqRlXsr
4zyb93paZqUsQZgraqFcJFzAmWxvUqqpyGQviWGXdR7E1mgEoRP2A4GsqiapXmsWZzO0aP8LoDqZ
6lACUHUxVasFblsU/96odQFZoG0+NvfZt+Qb85cxnGIZ7zt5RFtagcdYEejj6xQ/0hQVvJ9wxnWY
nBF3of9hBmSZ0dHv/ND1t6u6HRbIEFB0hYphbwhowXshQjeTAvZREl/GQHmuZK9pgUZU2jKFnj5N
TcQlwqjPEw/wQIr3KcfwtyjgWVxNvfPfVD4ZXs8zZmW3330huoV7Vm02oYEetD2LgylpVqcO9MiH
HHJCmsZScUtQPFTjx/cOZaKd6XAxw4w8u+T79w4lyQAN6zqUnpS0z4su2RTKWVLDGe8pwZ6pWiqX
NMWDn1HeEuGxblOq23HD8n25SHuhMTRss88I18crCoRTVNy4UKY6Fi5tKlEIyOnfEFtORXk1T5yF
p4V2g2ukNvkyd/r4jBbVzYAZ1bYoODPZ3M05OhhpjZ3B62kzBgVLfIPXhKR4K+jhPaPISmCDwAWL
TdiidKWKQExG8i1S5m6YTh7LVsqQLBhIdimZbg/ckOgPQOgwNM45rLL1G2bWcDEJRamX+93hFqyF
raw3gsgw7CnWioi9Q4VbgGVefdCw16GW8Rb1bB/rxw3JbyrNRMm2C+Sh7saE6JDHecJ4HUjYhw+k
eHPgx9KiC0iXkBUU99EM4yOxayUyi4ZAU9SMO+oikfuS5jaEhoyokpahYboEVrJZHSaQhuTkKqJ5
0pjsd9BWjIkbgcoKDuspQI/6JiHoq7zYNcV2qGLkFB+UChaPqL/BuD3fQXPT+nkJTCdyHJ7H1XAL
MjA844rUOAKvDKwVBhTVQ6KVOCj1Ln9YIg3QC2nAseE3jXa/mNLkdtYNlZXJu+TIP+gOTn1vPqbt
M6IoewwBuLDtoNfiqgEIuS6vFF1daz4gDRfRePqDec1Kaz4MAzSim9Gv3oahIk/jtm39ZSGaVDN3
bw6Ukb4gZ/KF5O7t0UldAKaM0XOpkB0+8P3BmPqiYZmeCyNEbXcJ9wN1apMu2SIcbeLCGOfHdjF8
vG0NRMu/zP9aMhooJHhIoHWotxFSJ5ZNTXpt5Gaqtf3dmi0Kc/NgruUYgarQ9KG0gtIffl2Jz33o
5wwN8G5m9mzOr9AhxHw/UsTb6d2JXWXrU/kGmH3JBjrQmrNjkpGmjhz/b/GLr5Rs7/6kY8u7yzZo
D1GJ+ummBxEFXftiMwlqsWHQAYo7RwBy6Kvxd7/yWNvUjI1xXevGtp7UPiQbnymfyeV2lCrWUfKm
UB9VRe2EoKBD6M18l5ZOB8ImVTF9CNqsM1tAPEZC81Ekug72mtk98pOYcZEkuUpBW530rBjoDrGD
Nn8eUn9cs9xng0UsTiWdUDF2TgKWP8t8Tr+2wD7GXfY7hJ0NZsPYSgiXe504WwKp5NnSwQsJoPTi
qslos82GLE91g/BVh6vo/gWzPK2mKo1fxy6bARR4I66qemxl1i1rIJUdYDxX4/sGcn7FGvmN7rOu
0h1iLFxDXoKC7KFX4QT7ROdF3Mm38V2k6qAn0/vM1CluRrnFCZhJA+/Dm99r7WUGp91bH2KyM8J8
LYORvj049MpxdUuDt1zAltHZ1LFbUdvIQLhWgfVEQAALG4dLxr+Oz9V284+Ry+RUh/FYUWuFm5M7
Z5MQEyafovolSXupBB19gi501nYgKyIG6PXAKAfhuAWWWLow4q1BlDY6DsUwtIYLsxuvoKO/+6u5
4gvYQf0kSJkuXtu253ONgirV9jjxvezavVafncalj4J/PkqakfGjwgls0xchp7Si406u3kahUOeS
XbxCn5X5JvmSe7gLqP1jmuSkcXkUdAGhFXWpyLcWh+hk1lpr3OSe7SEfyVOl47+nMrFs73lHFeTX
Zox1S9CF66qsxNUf50r5MgP+p0bGEEN4aN86vG3goZZzezlQN/4xP6fE+RB5mnk+xHh1lL34FwKG
GmFBfxmI/44BJwlReOrDfZF6zO2sh8f9BIsAn2GJ5ua38DSFT07K2bE0EYk85coXk5jS37ZLd+uC
dukATYjSLUMcR4vra/kqukI+0rHFNMo6omdXgpWTduH4dx0S5pWhKQ0QfLM2M5vSWEWfkKwPugkO
RZDtqu486cAnThk+teIppRTEW+ZLTM10deA0n03EhQfSHhkeduZbQ902OhZSVVBkGrnlflWme9w9
S12Y5TcJzGDNwK+SFvo3T/XSx3PEaUECyV92h1LDwlLFGKxpRgMpXpZFCLbEzlbNXgqyEYe0pbQl
lIMegn5XMJzEHV/bCHMN/fjntYAqtbFnLwxkLJA7Rc39v1gdT8EecjjTQF40vzQpVogu1yAl6pNm
dFo95toA7R3fqxac7QG6cTbjgsZrSWyZi9dKuI/GTDsV8CIaiM4+Ezb1SUbqIaP4ABP7c4Nxrgc7
OlHqKNw9tppaBmU4xUFSShhrJlumlOYwVVm18CY9mVG3uVK3ADa8M/DWnh6ixPvDb0P8a06ka0lN
zA9piQovgiyEXCr8oOrAWYbXrAGSvJGZExgC8eQoH7INlgxrgyOequUbVeOBOf9E2pFjHA5L6Eb/
OV1frR82o8KoTGrOBWbLa1kqXzoiNZSmBrwNJPEyH289Ug5A1BTOHkuwCViovJB0yNyeHTe0am5d
FE63K+BFPJqKHUcSIEc6dxD1LmPdjggP0y4N3ys2PsBI9sURb2v7y5w93CW5FMDEHu0tUA1KMHUb
xZuTQhbcy6ZIrXzaNLogzFWkG3CvbUZb3KB0iz4/7f4nwvs0HPM3Q0yj/6TqojyK5b0SxIn1sA5S
mdBlB0dbnVf22Bya7I1QovspQ5IN3ATaD6QooLxaVU+rIjfrtV/CrJcisnPBTxvpvBhD3VA1/2AG
XAY9H1HG+JY21isgSWAuiU+fVTdlshkTN+MRmCXMlz5fap4PSYb+wamkyrKzC8J5lAWZ+6Qv7g1/
wpJFANGSwMP5OLaSeWdnJNmmsT64/CoQ4/qI0q+sZFy9cv9rqVsFBKs89/W2MjXmXR2AVZH++jWJ
V50NoLdkxB/QBaL7bE+fWwBBVYXH4VUtUf5YOavgUCbuEOiK2LXuxRpcTtpCl9S/j/HFePR+l+Ra
W3NVX+wsd2wZp9qRyonFN3qcMJ4VP+I2xAyyZLlI6ArDZDSm5jnWjQxW3LJ1li8vXyaODkYwyg+/
rvBeKihOJ2+arBmgkPjFSlPbQFscy66Wmbmyxn/lrM5Sjd0yuI9ZRi/D1KXJkJ6LAwQ8pt7R5z9T
a4DomyjF7dUDJnvAp1/Dk62U6KqH01q6tK4nUJsxn1ULV555LlpIfL8EUulUvKC8BID4chU6rkMG
O+TU1whjqyqIgbgo9mEJHJMZtQZ7+Dy9st6TraVpN/kbhjXdeAPtqfjiuDbZykJBDJ4bBJ3mfDkv
wogtWHywv1cDap7Z6dJz8SzjXedADCUH46BZIm6Vdc+LGkqSJpfpN5ojcPbgu0L10D8cn/M4rJY4
/SSVdfNbzL22eUDHzSNXbXALg9iGCVALvNYtJerc7XlUqNlHhhA6AT/RTn6Cv2GD7cIv+Q2PT4ol
zNDBTpMZ9gtsXoFMoVvbdkNa3h5VrfuD9psSrq5LlnxQNdj2/5bTVTUHGu9L3ujWd1HuS7TzXgXe
xvhWABi5ijh/KLHMdma7TV1Bs2bvXKGF2lzCnlq0mIfixCdo7HngJXKZt5ohFeDeoIgr55eGnVjc
vOyOxg40AE1YjcZ/Y/yt44vE0eK+SmoO+Q50JZuFAg8g5a3TPfiqLE1lXgdJz7/e8C7r7Xo93djr
ZcCdu2W24uUltnmtErVHLkAFb5CgE2ln80xkBIdpVnyon3rzMqIlMJ6MCSKIBVGf+byOxI2LDYHt
S40jAc9BufmDF88d35J9rWe/7yhINYnB5JYWm64rUJzOtRPFjbtu7fBr9sEVUAd5CVoqGlQNtS9C
MK5zvqHRUm85UPcK9XSRPJ1Cfzka/TYiohxR7k8GGMJxgdLVOGzvWa6PccguJuk/i8LWQW0Aadha
F4k+NxYLnJ1FN8SkNNFeXYAoRFTBVhflTcVrlly8xDwwIw4IjTpnwGBWQR6/uJsoBWPRWgg0yf1A
JiUTW5e23gMPOg/8jDgGq4Cr+2Gk8JuovVHLeJ6R79zpFD0byTBgrEh23nRzNlrJuq0iD1LVrB+7
777JtG6LsBQ+nZY77gKnnHG6aARg1zLjNDJO+4sZZTx6W4mK4cc7g399aM3xb+80qsgiEdaSTSM3
pFLERHdfZN2JNBVe0q3nKOBDkQzN9UD2fdB0AoDpD/AUDqIBOVfSGSvRIYN5oABM+QjH0d3ihcJ8
Ux6eN1+UMzgG2Gman/tl8xYzXb/XOsYpUxsacX2r+GBnt7Ai//4oFVsayt5iTTjH6mg64+zEGaJO
ih+iqcTtpyMVUKZwZVVdoFqWrGt0LWQuLipTuJN89JEaqMrDyY+pmhhrWSXx6jQhFgjhhBAyyfuB
J/EukdIibCocE7QtXPwYR6tii/WSPqRpsLqTxTGnr8TbJuD+r566hBnDqQO2IGeQfBStFexyVhmO
RAGvOZL1ZIX3HsZV+HaRcJeUMbTGA+xMV1v9El7tJ9+Dsc71FaSOpAg+qeJJhv0zQYDcrtvGD1+A
Nd13Zp7qQF+2sQzxPvfv2wNbMr4yXWVPeIonKso70Ih9iccZaioDUPClxrJXUY4pAdXWFX/E51de
AIVZMADRl7lsn/nBE9jnByxZ4dMJhWbYdG4icD7g/ljJvKCR9UZTsGIDbg51E0dQYbd3JCjfMTx5
y/PhjoMw7mdI0Sb7SfSrWzVQbJpjmvrD871MNtKq85Th49OTVM+r0QZuHVjBbzpZz2gwtexqnHDU
uqunnCwnRAnId2SMs5q5N3RDA5rtDBqSAVHu5aT/3C9agPLoMRlYpqTF56GK8NUCuQIDFX7psmNI
2Q0n3xIbpA3IHn5pE04ZQVccLvGy0nSwMJ3w2Jopn4Xu1qTWRdA9OyDRsUz+sQXRUs0XBzqDkzcM
7/MS+ilwvBw7iAA1UlQlIsWr6dbc3BRCxTHT64RLXNMRPWxB7rI30rLuRyk79qXKm0xKPrY8+CM7
H8vaUPMp3m9C7dh9LeMT2AmTZKt4iLPvbQU6a75/Z8h70FqTX/uf79Vr0CLCoqqOW0/Gu1uih0wY
Ybdx1ZBaIr6R8DgZQbuiIMY0Ey6oXfRP9MwFGmTS/SErc0XrxPxorsO9nJ3ZiRm5QJC90TXtNaQC
niyeQeD7tyXp0GIU2rdRDnnPFH7dea8bKCaIEAagkmCsugHWTPFc2DlF/Hw1s1dX7+BHXAqF5yLa
hAgHwdSoDmZtJolpg6PoyJNKMKyEo61nVjaqsOW89TDrKQmeGNvoMtSYhr+g6Pqua/qglXNDYbwZ
nibwBSnWw3sK9869BaaB4ckCtIb6dVQ8RVYMRqiCtYlkW1ultG42DDd5bSY9eDLPBiomkzW+NYKR
VVG+NleZXxM6dwGmznbYBaJAXYs6k6Isv6CCGdtPW/Egl7UfAgqdsW+xsX0PA43i3DXoIrzjwwvP
uqU2m03pXjO4b7pNAYEzyQXJWPz+BhMmfjZXTGO77rN6tW1tf3yO97AAOiADWHxBn0E89atUHCgX
7+7xyDkEpVQnSneAeu79+WVjRQrXckQ7jOd0bKyypZPshSX79GjQGRTvi3ZVmfc4nGstpRu19t5p
rCR6dgg4P3nT6k5d8Mg8wvH/U1vMcXPWuRQCLPrgsgPTH1ZoDWJSNtanVF1MaFnfyuPbpurXr0e/
cxSvNZSM9Le9+LVyXvHnnNlMLpnP0OXsg1LTzlJkxWYc9SciH9vRJq9bqKDdja4wllPg8eRr6w5X
mDShwnZv9hJMG32hD8EyITrtFuc2iskknvJ2N/o09XqpyhbzlHNrcPmhLI1802iGsJF3KrlClg+D
2AHXC97xaW4FeVTiCznUh2Q0th4tXqco3pOLgwhK3MB7YwNmI9alFXNKN0fFRnkxc/RJgHeUJjSn
LYJMSdMHDsJIxtqWHAQC0xwWt1zzboM0fNtS45Zq8KwxY1lEkNuK75MQzVWosHwMvCZtMlTi582S
D2Djei/axuOFHl/Fa/ZTe3Fj/6zLRbooofgta6Cx1eQklZqzSKdAB1fn67q0j17RyJEoje1xRtmr
fZenZEIQ15e+nzJV8zbNUuhzFgr0Eo3M78FONb/k3qvsJ3ogh4DduAJthomWzK/LFztmiClPuLON
FTyXcCYU0mFY3gIE9oTvLOMLK5ScC487qnKnJAOctqfjwnBJIvUW0d8X5zfB10MAoqvwuaHJHj32
x7CL6Viv1Tz/kNgRs0CffzHcOd61VyHEMPti5QACQ0SQRs5te0DXHa//+7O15tEOXviRznjlY/dg
2WULDAuucz0LIgoJunhlS5SNmZievn7gjw1ZJ2bRhoc7Rx21kDTy0b3TmfrAeOLxvpEsYNoN0B//
Zn98gxdtIJFijWKambnVX0bomQve5r8DoWztjzhnRz2jBf01RhdJPkNNgaw+PFdBljyVZD6u9u4j
Ra5PlkkFw8LBKh6DGscamloWd4+Hw61Io1fCfRK6cgxJggreN2qD8bEtK+17to8kYzIUjDXsJTZ7
7m8qkEIlWuW80gkfIEYaWdAlCGVHgSOaiWv9tooAhNcJs7BVMMgcKC2n/TaeyM/zd+SzsDbgcTAv
7nOuCwzNXfFqGZhFLmqGUwyHZbuCVianqZJNMjyDIeU2M0BvRYm0al85LR2MSk0QlwIo7Getxjx3
bnnzG4pABqGVmWluInnC/f/eqdPr/+ncZ733FqP7g5sod9cHCCzsV2R7mMNywpkAFzsh9yn0R2xV
PY+WYLUTsLBT9mGYJFD2C9zeDY/D+bWVhzKh/QaHCuY9yvMvtkaC2sgZSXagEafQWSioES5YPSTn
MBudyFxnRqc0Razuil1O8Ll5xNy212cq4vsHpS6MIQ1kWV8yzgZsqivoPcSuG/b8kc+2ZjprCLTl
9QUxtqrAFGzTnGYP9u37BZsRP3VB+O8A+0Jr5GHjjnsCK3Dq/MH1dB8K/bspF/AZshH0rtoTgkeQ
rLMTVTH+MZoK2mUeKONz3vkWHfs7TajjHyQ0eAGhKcyOQAVxNMtSEGzlQRMBWx2WFGDBrtisOTvB
p5qOQ38zqW0SlcOnBgZalHQRWpXHnCYWUzfvewq9nfjSLjrPdtPRv3SF7vu6eh8JqTz2Ci3s+doe
glXk0Gt+qsV7pbnIi19hM9f/y/K7dR3kxr5sBV0JqHLGifrsc2QvWJm4sdc9kAZ+BZq97GZ9VisJ
ZmTpdwQE3iH5qY15AJUPUdeiEaNbJ+zEBKdPYPPCgAvMm1kHy0WZC7S5dGOU6E0AnsGdD4OD0Rm8
iapnVGfWJtKOv9awYEviwfp7n9KNYC7IYAt02rrOcDCz35l4ezvh8e4uyvTWGRCsfnPS0x+2PF7Y
egONLoCFzhSdk2PTBNN9PDk2um4TwFQC/loo7qyrF0ylB+e8YnA57kzPmRV0ZkGmwvBcjoojdbck
pvnP4NxZ9z24n4bLHp6N520K6q98uVACtBUFR/VakOHiM8RnXziFv1KUivSOcJCXmpZz1DpVELWi
hy4MGbRHC7OK3ifUITn6Bl8T2V/OlrQvZoEFFkxSp1MxnLjBcRyaD+t9IPPjBBEWrGIyGNfi9CL+
HOaDQgAbAQm36RL7sH+hybHPOmKmkcyA/yzHWB4dEhhOhm2ZV5GHBYS+iH5x1ugjKb2f8bRurFB0
L54tSzcJz8gVSs2xDr5SToWJ12uOBW6c6VGZS+lpetJLTxkd9s3zkptmGUa3li65VP9sq2dt3gPj
7QMtSRVFIIyx5k5cC0UELcVMpggawDcZIv46VdiW6hAfGRRaadiAEI12sEGIyRTz/fKmDqhg0aj8
/zB0m6YpQ9XwSjHs4eusPEP0haZw0VRIbUH8xM9vffpVvkNOCdcIYsXguv/eLrM3Gi5AKUaVVvBm
MHgG+LngZzOVOBKRKB5EM8AXbUIyrZZ8T3jOmb1zAmbtDfispxMNMkcpfVZYAvc68YgwqUV5oTRZ
dyUYC7tuCh2DUcSEbuKRfqSUovRfeYeJFb7XrYjYnEESbJ3mBErRR2eiR6o9dlBL3FmRq7bwvD2O
tNeYBTmJfD32KtY44iFVrkOvYVFDxVJaLhEKpWV5vWQx+wNKyNWpi9gIWCcnTPTwPkf4QkYEGlTG
fwC/QdatXwUTq1Axmp54QXwcCFQqJqf5OmBc6YtCdpcpIfrcS2s9ciAIDGAdnz8zymBeq/w2dnmb
jLJmne4vvbO6OK8u0natvLLRuv+MoCJkuhe5la3FKFZiD2bVnBRufOrAC/TSX2XbfGTXogttiIoB
Y/FhSxQOHSoCI479PXLEAKzPtfV1qUoChIttpmxPSnvJd36SU9T2F8a/VHR+cjAZAZ/DTP7Rrv26
YTBYRD6dCDLHtnAZZLDhrWryLqcNah9yFIEW78ECYwt6bhyeXxUye/2bNrzQzo+ajVqV3YMOxOwC
/x8aSpYZZrgn0KDipdlyOpuG9Vb6AH67wgYLu6lj0lTDl17KKN0Hqh9OnCE51O6M/7meYEqOwAli
kUsIaRnbvamFMYUtcY7EaV+zNAMvJ3vrzqoFNXv/14piXQWna7JV9sUcoMmqXsDXlFtQaGa7qW2U
gXMJ4eUmOwccCDBo21isk6mqlslROzFHlW8z0oxztwIDLj9m/Bev6jqdu2GTwv38e+zubH8H5S7F
9z5fo8uSlkTuPFJ3QUMV/2Nl7F2RLb79KCaran3QDR3xxGs02ZGxGMEGHSfs14Nkk5YHc9R4xjEH
gWu2P9Vx4lsImUh0aisYsxkqDUhANA0nhdpAiZYlSZZdXPtAiCGFLktQw5gkzu7lL2UqEavvuAmP
tbUPbniuT1/3ZIm+WlUErspJKieIckN5e4mH3wSjhUvCHkwLOW5PzJ+rcjTyY1QRjSpptcl6gSuM
pe2M3p0ULaaPbrohh/0XVRXLq6dVlJ2fHbQf4DXY87kSW4Jn4XK9hzZZMSJsWzoiS95pyH56CXt+
FS73SecWpLvKlO/kPQ6pod7wyq4I4WiKv/KqudHHRdTcjWli89EbetizJdWGZXdsimQF4vmJtuO2
g0GJwM7TPCxIpSVnWhzB9Sj7Sof+xQyNazrfYoKbb1FH1Fd05/KAjA5vkMbwegSEJzBkXnhDUZy0
SKHDYsDSbtkDEAVD2kiD0IwfhCt4/HUw5jUoOP/9SwwudKdNPWnJYavLzmZb7kiH8+yCOCGwI/g9
FB8UKqusN+RMWJegjXLHz5WUaMk1f4lO4afEdOQbBlQ7kGJ4Gg7n/9r/MGPwwJaI0oGQ3l2QlZMX
m4T2sLy/OXgGGph96Tu90Zivilm/lnQBJ1U8rjZBVIHglPp/ekYMZI2YQshVAH58q7KSQ8R4H1bQ
pzE7OzoLHPuQtF54+rLhV9rghaQcMKa8Iz6Ijpqrk3EJe3xudiUji4bML3h45mCnw+XsuFS5bS2L
ZFaXZajTCoLlxhZJyHrxXm8PFCGlaFi5l/hI5XnO0UOeJJ7R+DTnTcEEuO8w6kjnsQaXhHWLBja3
oQSvHEz3ZNNWLZTTuWXzx7Y68UFUvXYrY2sRWJH370Lyk4Ntf9FjON018zKFOEYdpYywgzfL6Pve
T9UdbvILq7Ht5A9nW8l4gkUNXE21Sv24zsj/XR5WYkb5TF490sjb8ycM9ET3jMuBYlI8XEXfv9E9
xUMVuFfg2VEqEGUOmJmRchMyBNNOjt7QsR3QI32vCIo+TlkCjtNerRQyg73cLB1JuqGNiCqeosHu
//LVuDxo+eV12WQ/FEGgEckMMIQpFm0uT7aRP0QKEKwG80UVTrIMPtFpVXTgesVPDlClm1KluSAw
wMtM+LrUE5LbQ3bC+yTHRd/0jpHdNYME70Pm1qjYH/YApqLxcsU22xRwWCQvYk9BHa1PeiO3oZKF
OQZPbZh20vAHmBFDVOKyARRkBbBRSWAA+NpFCafIpEQ1rmPixApElr7XGInHm+PlhQBr2Fcjyq4f
NFdl8pEH9P6f8XeHU1/7bYMsU/8fjGFerKHHeelX0QBQwFHK1vYJVPJFcMUSEnuKpJBlQHQQOm+H
Ny+XuoxuD/Y1+5e35+lQctVreJvJ/P75Ioei5OSetagMb+Di+RpnqnicV4vc4/xRVXQoocN1TAft
damQ4kAfpg/yYR7I3kLTFezryQ48nlH2H8ogDUEmO5/zVzncZoqGgNqWTyxjtnBY9fZB1NZ24f6I
XgZ4vodpOszg2iHPzA3R1m7s2dlmzEqBcv+IJB5E90mD0fFUpVfwwB+9ej5nSxnBVdA2S+QXv1Xy
apBCEuo6DMbg8mEFft+WRDsLRLEvpmgYTTm5U1ZekZA6RYTVjx+nqfMK5F57BjJ5YMOtmjQT7x8y
CZdi89uAoVvcrT5GsfSQlR9tv7sq6FH8gVX7YpqC+Tsyuyrca7pwhFgoNI+98K1B2V6Cc6z682nx
+Dl5eJihhLuazQ7dLDHN/1UF4kaD2IGfriCgeiY16jMCRhyuV9UbZJh2UpXiGOuEGLPYI+0gIJ0Z
LQsa1mpfozNdnegYiX9YYwzOgfrgCzbPQsLPYgtdLUhB1SmFKWVhH3JpMU/nQMHR5PiTxcbM+U4L
rnDyGgy296xH0ZwQDlqH9kh56Pydwv38OQ/bbWKhHMTAHWLeJqQXhdCR6/ep7tOz00UkbH/UXxQy
XJGdTZVK+M1E8K94dX4K0z+wnRVnvqH+QPlYTLmKetgnmuL1ZkmItStJ8NGhzpY39TGIotdpTtPC
e6LpT7qvyqLp8clVXnvQpo/A42XkosOcZ0T+FePiUgGdoO0dxRkvf1iEnmEgguWaOtLS7HVJ1J9a
7oIfaQILh5BcoMQTMFsFRvUY0buyHUzcKFce+cZy6krtURS7sU/TpAIfzHzQMnwNPMa77kLgrC/A
2IcSsNwNZMrEZqAQJIBkmp19t4Pe6w4CrWUn4tfLy2WKu6A9wwMoAn7OkMecPU3fRNpPeZREAmzI
vAKF4AZdR1u3/Fznp1TSYSqoe5nWw1dVyE2wv2NksTCk6xWfRqhmVdufkdrXVDWuW34JR37rWvpM
p2WNej1v/1IXcxs2zh6Te8nUUU9BEHGps+tECr5T77y6H/7FEtdLIRfTW8c29Dp8rYiJpjua7c6y
RP2MqTwpKWr6oCC1OvqN49sxRku/HF0FraxLclcPn9tNDG8gf4E7zZBeZ9QApj/10pAE1G0f7859
ALXMxxZ7OP42tV22IPxPIyXXi9kPK69fLdCaUKKc0lyB/K1j9X3B+2ddflXnpA1Hj+E0qXB1jdCO
B7J3KA7rc3jbVVkFYc/pleKTH4nk714XwL3jiYUzNJ1wutzgEm7Rm3aPdirKtKOZt0iidb6GNuLU
xr3HgNazsPtZSE76GuGsNCvVKmPREjanGKnQn0bWJY8aVeH9tJP1OjOxOd0G8agHIlxYDKLgUVQS
bQ5RmcunHrHhj3t4vbtm7XvzjU0RQ7bnTknae5bfgbrv0odhgIUkNEHoF0Tz8FoLQw6Yrq4muf0I
mpyw1E0Xz9UHW0KFhhJQqDIOM2oN9sNhQnxsBnR6Zv8NwWFLqQxKe8GYULCdLSBuELmcomz8dgug
yfc5GobNOEtmERWWBloOSLaVBegxeuG4FNAgRaHjG8CyNKU6NM02jYJj9dPwtITYjmj/sNO3dw6U
tQnGcRFxZhV6kZllf4xIeOPIGWAC4q6x0lun465oI9wEBmowNVc1xWAjgc6aW1q7Wryn1mgPZy8V
/V2Y9oxv5Mjew9fz5I1V+2gP5vCNHRd8VZF4Y8Z7a4dSbzv02L3pqvMXyOYM3kRcJPedJJaUCGdS
STZf7RagaQvflradG137COAOwavj6UvYu1PUYigjfJIVrWINmfpAYseBeePayLPnpd+DvhmuHp6I
NsykCF4t6BhDjiP4PZ/1nD+Pin8gHWWk75ntOD6ljgVfdCXX0WpUTea+VfL6PoHV4z1GCvE7uxk2
jw4h5TUNPzbQyMBv4M5lC4kmPDYgX5Dvt1oyaRFBcXtP85jLs6YlqAb48CWU2YOFEpTDjWdfEn58
QNEV20L8ajXCMX6h0Ur7JhgvHRGxVDsWQLp7pwZ0uIRthi90OvRgCp2z3V1D+95Cmv+sUsnXn2yZ
I8KTKgN3SevfznoPuf+zeW3ontmsribXojnL5dz6GRCHmVzY57zfdkq44K/CW/hpD+ZukoqMnUNh
uH/npuKR588G+qo8sQcKK1wJ0gfrqNQlUXIsdAEdlXvFZcJeg1EYuPd57J6L/ssNp1S6VD0t8fhX
RISkO883aOx4WJbJxvLavQ07jCDt0Uu0PTDsWEpZE4pazgbm1IwYMHL7Kuiy2AlLEKMZfgR6Vv8E
gVIUZNYn4tBudVumqf3Ov2VMfSGjiu6151bi7Y1Sp1I89XN37USa2Qanhbg4ugE7nTKieO8ABxpu
BS50kezf0DnL//xEsosWIvutp5pQflLxTnE3TQrYSpF8UY7g3JlJgt7leLf/ZY1xBG4zmVE9HOie
G3TlUlGeBIZJj+mVMen9ToPtfGZItML9SjtaqEREIodDlo5qBkTx5n7QFYzswBgifcyEInKQEPBN
87khGYEWye2EzNhq0/VURv7jGp/DjaOoXsDGqeUCyECZE3AwVEg2oNoQWADtgEXi+WcNH9BB9NPu
sfiPuGl632r1uiP+LGOo1+BW2FxzJstppp2mppY1hqL9Ztxf7F3MLzVOQood42s75wKkA+pkExSm
hUq7hC31fg3Lv3atr/WRRBt6cl3UpfrfH/wRvpsXIEWoANpv0Jat9R043Bvm9RkQ8bPXlbqMX3wi
X5pbbYBz7r/S3LWd8tCUPBK5FkPOzP9z6FbNIKmtOx1pWB4SH+pCOt4Me//MKr9uDLeYoLsyt2RI
a2uhte27JmxBkjZJZ5BMBF80Nh/tracairD7svNvrXqU8Erg+Dd1qKcM8DgHRiTD/6vGsrupTSoE
tONYGNb9T/fLIeIQkkEjl23qjl/CHU3xmSnCrrtrTmhI1MzxZZmCd5mjdZSA5g1Kw4hto6VZWCWW
61x8TXnj4rA9CAaUocQAfezc/our0fTUQP+xpC1Qfw+yfgWNjpUzrUsnsOen/1wNBOoaItup12HR
RWHQNSp3dwv8US5fSy35kMFZCBNjEa6fJSLHbKz9P23OOIthTft97MdTwPWeOkxH7RdVnZT09mgd
1Xwg+RGnhRF9ps0Y3sArCNXBR0SML3YB2UWpGhuwfebIT9tcy/V85WjGXgq+6kyiJUAHZw+jgYiT
HJjAUQc8Rl6NePCGoqm6yl/ruS/U22DBVkiPME9nM5bphGcVC4aXPOso6L43AlY6T3lddeaZi8jK
Mdg9rbAr3P0UBpBXrwZ4Hxupmrb9wRkfIFvrkoZpCBIVOAj0Qd46HY6G5zVUTYMhc8Add70lb7jP
ABdkXC8zEJw7GtPVI38WqWjmHOtxc9QGJWeLpppn7yTWmihYmJik/thc0jlImp+ZHrBF2GImwpXL
Iffnmu8+8RHbXBkKBWh+381s8dTRbPUxPMhaUCOdmTS8TWt3aCRnUmi9XZ/eq4Huio+FYSTPbAB3
SGvXVGMYkPF1z+Sw+qvL03ffrRQkhvBsUVDxSrwpM8uPNG9ogTk5kljLYx1HOO3taRFRCmMPv5En
WLDwHgsi9cKP/KU7/2uuYOFvqCg69LqRIHHAluxam1coMaGg+OYA/69/lra89eBfHr6HYNO2ztkl
96iGiPBidmvUWhXhTW1wpzIGgHlZoroL/4qjsvE81BLK+4nvKxSwLFt4fI39QP/EMcKRw1eHba9E
7kQinGYAdUcQUgaQ4vt9wLhjiZ/O9+FSi34tj8559RprJ5NkUslU9icQpEOlxBvZukQlmJPH3DAT
42tmnEkWamfxi+JkUPsDzMM5lIsUEdSjUe5YgQ+lsrOGWYBKipDu9Fvisaals1/tTV3VYmdfGaz0
IOB8Zjhuzx+OOlFYdw1hMrGBH4nuP5Dx2y/4dOJEuMETcEEWMSW2Wsx84QxDHy+DjAuVKwyvDMsy
MHRwi0sYnPizURdsfJJ2zlf/8+Kw29CHo8ImybzHmRHbkDGwHA+AE3KOU/ednXY1ZvOpPENNzLfA
DRAIuZkN7wOGAtjrdkju8eZWeC6MGUpzgzHp7rxcB98omu7q+ZyO58IdfS5IqQXshpU856Le0GNo
H9dTJ35rWa5W1ul7X81oR40Y5Yx/p/ADo6+NaHl0z002u/EG+wr/eeQvhG0CwA1UNApqOEBu6GXz
toMzjxUyZxZCpLtgoo1qP9nj3WcHTyX0Ad51LsjVLPn2lhu+uusN/mFlsD7IN0EifhokiqdEwXOS
A+GP1oHacyfmLRDEE5NAU9yinnIluw73nLY6IfxC5u4W4KyJd9TcHpZCxzBL4V1I0/cKtR7iv3th
Ag1OOTh0SuB9bzkUsiwRdx1u7n9cn462Qx5KgSLZwrlU+CSJNGeuYHMl91kPwzQ90QG9fSbwQYB5
cDMJ0TEOccyi4qYzZDB5e3/4W4zugI3ij57/IgsfhX2zvU6gLhzZwjE5OtDTpM6edBEPbhuRnt86
tJjv6KaAgAwRcLZEKogLpHg9glkwU1Ilv2yjbqDAQXMlMDOTYK4+uCmh3Sfazt86IXVmX3yIvW41
Zsm8r7CLaxXpG28hgHsh+PdKzcphECP5Rwi/oTSa1tGKnQLVIsQKkwpDHXHDlcwTfP04EAo46hpB
QF4ClAFE+ViJ4+ZkkWx/n8EmE/Z2CIRD2CepTWCFUk47OMgjwSA53IZNMNSbOxETHSXa9kMUhSAK
xrZQK3IGPjIa+wrperCE/3cRe1gmF6XpBRjxSe52+jP1rCJ55WYwu6s4MmpstbJZ9qahpL2vnscW
lJ5ouQgyOLL3Sb6PjBvtjDamBh3tqDmRiQQNjemqHoRQ0hUK3XG3S9Dvo7i0PRrM6+o9/4t2L/Dv
azEYovKvHMn4Bi9iv+cfxxHRYE933Ve0xX/fFy5mhMOsekafXycZ81EkJCHHhRkDa2sZIkjcGWYO
3gt2IByX+GqSltZBK8vXZmcFeO4kiXUbl3+VDL0eskF69R9FNa7eH5WdAEmtLkrTQMfIK0GmryjM
YLbU+y9cOwqNNNMx96mrqhAMbN5E7I490Z6f9148ptd+x1vqfC2JdVBtlQ3QiXUvF5fLb9j0gMqm
8p60gvrNfvrK7jQNleod4QSEozjfkouhkyWoFY6wOfcHelIa0yq1fVx01sI3pQ876/QyNM5286K8
DyKqJb1V1AJiU4HLvApNVf4HRvCzwGokne6K0EOZABGkEvqc6j/mmj3x5Tzn0eLFbZmOtBLvRwW5
6hvEFfTO21nsO921XbnxC8aVtSHbSnTrhQHNALBeP53KjOndR6buSAwPpvHs7/TtDM7WtKk4xUMD
IEQUns+EubRX/3og2ln1mpUsoSr5OM74MHGz9D+J1rCw5DTDzGHtCqIhtYGugk4daYK2tkc3q96r
dYJgju5/bP8uWBKImx4gspgVVomKQFh1LXeEfVr6b/wXgw1jtpE8p2AVhl3wuoXt4pRpk3grpCpS
sq05mGw3jre/nJQjcNad2cufJ14HX5f13WcHVVVrix/qGdDJql+EoiFZyfqZ+k72z4pjOXlW/13f
81FGECbrCgz1q72cH9tH8sB/xxVi7se0sPzxrUSPlp3H93oT5hSy1DIx/1ZJwP3g+1klmPF8SQKU
r6LZLFem3bEIdeilchFdShmR5ehdpoU057raU0tWkWCopDofmP2sz8oB7pldALQCttA+CsTwz/Iz
km/yYsSI0yFPGffEbDAX9woSihAavw2WIxO8AtLHkT7J4QZAjzgoZ8Ei3gjV84ajH1oNOwDx0Y+8
VuKKn/KSkRLAB19Y1NQJNJkDtb0CJ3zW7sdy3J6n7fdW8H8q2bKJGe/drHWHQLZYLJnJZ+PJbu97
pBco13mMIclTdhsLpRXiMJk5gEDh658YjgCDY3Jtke0qGk+pxy/o8iNo9AJ7AdfNhy2sub1n28To
Yc3SCSn71uu9kO9ilpd3Cz0idPy+bWZSoizH2GEeh6yOjCYqgT2BjoWdnje0eo3f7W73arBinrIj
6/Cl0zIQmYtXuOD0pvBtEmc5zlTjOqbKwlVIfMjc+54U6D30tUO70nMBYMWE1xDJKuwc6/w6BUdw
ZivuJQPbrjc20Gf+F0mX6qh6x00k0tiVn/WOH9omOj0ytU9xEwPpRnLBelLbqdtkzm8iii96Kr3K
3iKkQdIIkRdu2tSXdUzWV9uWsBW3dONdsAAa/gDmY7KPitYohmjCGQ2Yzh49FxnN6iZJqlPH9SKH
BV1Gir9CNMQwhnc6jincj2qEyQUn/Gdr0KpngHvJmocdFgmMFKliktF8EIQkb/Ew7ld1yw33BMPj
kiMwKGeJqq47c83DKCXgqSh8ZG2KpW0ODKB9pc9l0ACJLUOUA9OH5Lh7zV07zCD7G8teWxn7bC1P
uIOftSeblcVXMhRxxb7WgEpd/ME6nwWLTiNIvjwMpl8s98v3MJRWIhJTQ67qLreQJckPV1cBjC/K
4JzB+KkU2+3QiIb2sIyEQX85Xjf8qswjhueP8Sug52rYe0crZMQd2lAnLt7AVW3bxZTcWyh2whWd
EijBX3Q/oMLZqrKpT3+fxeAodl+TyoZsFqGYh0FPqmDo/FUDILX8PGn/nlQ7QmCDcnQ0rzSDZOdX
WrTN42hhP7j0FhgPxhMFo2UFqk5AvNVHR/GshwPtm7PYCF9a78SxiPA0iMLnyLQYJf7clXetWLei
wrfFhF0mncuKoJ1ivQ6b4ExUq1l+kmqH79x7t1zmj97r1ZAOq6DiFHeYCk/lTx8nrKtRx4CMiYGa
+XFwI6wBwvA4HKmdU3C0AAO6W5KgrKSjiE4GT7F6u4yypVPiDkhu1w550gNvstQydgX6Cxwu2G7p
0B4QmqpDIIcbDJg2NcXnZbUtNBE1NBQnmWNlu8C8UeysVeRAkFqnufyjYduTIrI+zmzYKDerWSIM
1sD49zl4Z09OWYncgs5NEWcU/cUc52r0r7HkX+TG1MSG0BmcyhvlWMudmFVg2teDkdZ/b67cqNqV
n7rRuFsFsAINcTfUdCUyaEZkwy6C9tA/yN6x1g6z5tUimHm39kk0q5s2xKg73nm4dXBM9UoazVEo
Kq0QAu1+s3RKCkHQSRelC24MPpZBoUcOsu6lgzmLOlG6hkSUg8O7ErOqqgIBLmBRdEVYK1Vumwih
wW0+thC5Lhr4Zpsbtt/ezzohF9wu6IHVOcTR0erqUcQxYGGGOBEZb6lRq7pFpFYyn0D1MIdZ+dNu
ky4dPm3iTyvZ2NPDYV33bIyTZSCUPhsZ62y3sH5dXKRaHX4Jz8qWDmyrZINskyeBnje3k85QO5Z3
bRLirjwwlmx9PaWVAsvDjHwSZP9ikFWw/aRSZdhyRaDKIFDl6wlathyJs21Qv0bOjNI2JLWkHrTu
IepHs1y5dHWob4DGXQ8UfMW2P4fFFCnYsmXGx3yj5XDuinUsIApGqDJx4XpkEal/iJyczA/iY9mv
DIS70BxZWwVGd195PtJdT70mbJhvcoJsVOaWD4A+4TLssoiutzNnpOzQniEONDnaM23YgAZMdA7A
xfJ8+jYp4G3ymqkRojTnxnLtg/vd4Cw67/E2CbciWIP8TE4LeldSsTNlGKegnrG2rnWtojHWyJgc
LJCQsaKjBo5DxjrKvBMjnL9I693C9D5MCSASgoNhN/A1KTPO9g0AE5ACpQDRreOxwxZWprZfOTaE
99O919eK1y92mECnOs3PLIFAPxtJMqStfDBOBr6muEKse2a6dBj5H/o6OqfiEovQIxscNXndSbyz
/ijin7BuU0u7ZSIMwhpW0Drpw1+/0ag7GNLJJPt+i9X2HMB/YkXaIk5AMnWhDz63YBZc1lkzWwPT
PALpQKTJGbLqS7hMz/QdQebmGK9P4EuHmFC9CIDnfSt3iOIzFZGLjxpybyzGmgpOpsPQOi8D1DM1
EXBw1da+zkSfEi0pjaZMEBPsGADguXIkwKEHaA1144wesFFQbNrS2qY9tS5991v1PF9zr/iCENJE
yG8+/uXNqVrWHK29aGXn/eXakw50SIkiXIsqUyUmoJkC7RCFdOmaA/QubaXKvptLi9eeLl+bUmdr
NuJsub1h0vC9hPg8R8OPyxOu5WlwlGmMv7TRlQ8pE2KRZ0AnHYNaOMRlewSWtobwJtYoHpvfka/m
yaXZszSb3KDmWbnk4q2X/zI/3gONqhZLl87uQ5u+h8QUQcSE5q/6OOCy/6bVu1xk9zLAZSTrcM6b
UMPLajZoRgWa2LJCzhbBsKfpGfPKbefl+1eK0Ra50pOuktL5q1pZRDjFQwyPHnskmhen1Z9NzqW2
7ANxmpIBFobynPBed8EQz/cJESN8Jrnv6X6fpqYizn5nd79nI0CLsE8qrrN6i88uNUgr/Ohc9Tky
y07Rka0wIYXY1TL6O7gU+KMRS806vNyd3UL6SyUuCjCDPABtqhvPpOdkZ9fcTx1WI4Kwju4VYOWr
w1mNEi5HYxDAZetWdPTN7iusaCmw9CW4yfH56CU2vZjFBhaZyTt4c9LPMz3vZ1VUsLQnJnxG42zX
z/2PWdBIr8zrVtvKWG8d0eMfsgOMtnVWpL56NKgdxZFLrayFd0XJ+cg/MIGadO34wantRX3btO0d
tk6SClYc6eQIy2Eo1cxsmQiXVwj8piBaDWV7wZ7gEN8YfbNjntDGboTL9NEFsoybiUsEraBO0wJz
0+ZpxsZJcQZZZDAxNxP9W+CMuWPqtlJzJ5ZjMWasSVgfvDbA6zrf+PiR4q44+xFR9+VrCTZkPJsl
u4p3zmh9De1libqAHng7bW9B8WCGdcQ1Xaar5dOMZr4ZAVEG3oj6vFe+0QD5L9fAK/Dr/eNSwAOP
jqefXNWs0FisJTbu26ChmP1tDMkgoVxKTnd4ZcfaFfd/JFSohJNXIfNF/UDpi2pcA3f+thAMaq7w
8VemD7XhweGTB9RRJhY0y7L6dzUxe0sRLyYabgk+TKlI/qIURVLn4gRH65tK+Pj8unguGDv2+f0O
dj+7nsoQ/k3oY0G1g+l7xaAC/3EJXZMgQ2RxUSlm0/9K6A8sAi1iyDgkTMWoggVm+UzrtefDIKuu
eSvuXnUuQX0qShcwbDDL+rO+KXiQPdkRKiCIjjrIXvbDWGjq+0skqdFQht3vkUMk/pVRTSsF+mbp
erA9as28HFRepxv+aEap+MimAH5vuWFELQmbrOJGxEjSAbXCF7q2QFuH4i+RKrWozgFHw9tDwmuP
Ufs+wmyNo19pjuYC6fIwHHk/nniw8zsS0SX1mM9IJbiZXiLN9GwHxFM4vY9PxsG1r+rr/bgTy4eI
UcZ7yauVB4DpHZvDn5o74PyToeS1ex7bFXOOxKG1q3apGf6aB+HAbn0Fwjg67FgsGvfxrZV+Al3Q
hDYn/XhAx/M+LBarV9kMGAL119+cBbCBgzgzlKbBgHS6GtEZXg11fnmBhG4pROrmoo1IZqCXnNHK
bf52v2DTmwKN96NUgeyumv6IKRabkpkOQGomb+GzQeJolhSKLEpHRNCs9iec0em6tNCu6bmGJO57
D7wwmWFoJFz/cEmK9mgIXN0jjKtHg24zwdUszX+7sTLaso0ABVw5l1fapk9F7WnDwlB20F6V8MeK
cHG7WNXfWXlFbBkkYwlBUf2QXn5irkhuGfee37vTQoK4l3hZqQcWoXQahR2aeTqg3JvcliZjI0nh
U+N4WqIT7YlUujkuuHZVKaoVnrbMBFtot08D743Fvxy8vhTeeRTAZkJuPZOOUihkMK0yefUe18bf
Ztg7rmTgRrPP8nTV1JExxUZY9jn8PBraN5uiZunspaskBVbVWRySbT/N8pCCq8nVzSthQdcmAY5w
cCLa3fLASd3Pb9AHBwiEhc7rZVMs+z75+YI4CuIfZ++q2qRveLiapIJOUeY8QMHhDjBkIpVp7S8U
L6BBGURSPG8nq+K0JE6wDjuQkHqw3iFy6maRzqZatFOPpUIqhIK36wT9DCPszaFVYJFb5+AjhmDb
K/jUsMwV1mWjJiFfh0u/RU9Pnaemy4p3m8RJPFXeuwQSfdga0vBdADhz5AFdXD2vHtpEFzDGj7Kh
F9c1/OJz/EFXhrJEXLo69FvpseMaZ7AkUIduKPyCwUy6zk4uBFK64G0RsUSSqThWQVtkVPzl1Byi
VDIGi7j3U0+vxGSI4AhWG7UpKs4AlRR+hJRmTdYXMLNEAZKZCND/iAhO9BoBOmGyuGRhNDPzzUA0
GYK89+UGoXH9I/Cf7tMDsoaM8NrraEtCWrlFdXNBAFqmL8c6hiw2LIsrMC3KguN6FDfFbZ4RWDQZ
pIwz3i3hqiE5Jq11x9JgQ8HDj/Ay35fQyb00e5LSo0t/m5bykr/yy5s2qUNloaHe0pcHZkI1yuxc
KkvLIo4gnOnUifqZcVtmxo0olZ9NBW8Iq3SujUwlPt5wFdCNH2YCtambwtQtCERQvmoVl6ubsNbh
VtaEuSTgptqr3Vmikn+doulMTmMrJu4NPXivQmKMg6NFGvXGnG3MiBt3pgW8MH/MXODkD5yEJL1H
HKSYob6ouShcHWMAzYW5EqULTGJWaOEBVQdstEtGbFRxGXmpXrEBSQ6sE4NOdVPi6saTSnQsqnVw
WPm3RZiw7N8wKae/9MH5WX8icDj4Gta+jQGuk7VCAaGAdStO8V06pIdn0LgCOYDkPjTcr2nVynil
e5v9nT9ordveQYOWQ/Gi3II9JLAFwhiQGLYA9n8Rw7hGrT5wOqsFESrTWJF5HL+0hoBk7cG2PCCg
8ciOUNM6z6SOdeU1DLyB84ftgx9jirE0ogDUXrrq0f5/e/URh4yHfJz7mMIafdmsDt93dUBdOr47
kq6HEzEsCqqeuJlqAGH8UA0dqn6+c8vPGSFEpnfNd7+U8cGa9ClQz6McpPX3+dOxPJbk5P3DgMWX
NooNMVmtUtB9Bl2/sVhiCFLx52FxbB+qjFH5yMgAaKtsuKIXs+oZgz4Edj7TFiIGu0dB/SRaxoKU
Ch+o+9GJQK5Iy+gvd6vVOJ3iIvo7Bs95y0OC03lzWjJ3yCsqqC8Xw0R2IDR7JfoVNeuaGK3F2KwT
m+N/e+oF6J5qjfltjma047b14G9gEzmDIdxA6rPvJA067nrHR4SJ21yXM102e9S+erZJbFEQIi6K
Vs9TkeOf5MsJu5NYt/9ZvQgE92lLnBX4/V3uxWxhMfjNoRA4d0kbiZqYbXZ9wwgdH5I0WVdoJ+el
TZj3H9mlqMNCX21ttOxITS9QDIiqaXHGFtgMJd6vqNddvIPzHET5kI2JYk8ji3gtRZc+da9MTzp3
lZX1PT5FI4kIT4EEWBvp+NmMRVHHorDc3+4DPkzzMgooAFjdwV7b75SDyouN9fMw7KHLfbZ5ca/3
JhL05m0BysTMm81nY6nbja+BEKQNIfzAmI9w4eoy+Qfx/yNWZOoaX4pnEh4U19eGa4KoCDh64kpe
Xy2yN/SWBAAI9kUHvZSJdprsQ4S42rR9RM+rab4IPpKs+l6kc7vywR6L2h6ajUZ13p3vdaJOiR+z
Y3pOPbNLRE0JyjElIayxf9frVvPs7KOzTQcfe9VKupzHWDIPFacBPoUyYfrQL7zWgsW+WfVeeuRL
uywnUbDf9w/v84/6S6XjydnKcL8/hajM7Gtjwh6bXAFc+tw0SPDBukAN9ts32uW3x76VJu97zJha
Fw4BoOeSZ+CY6zNCKulxuY6qVVH36rgQv8t4VxcOVrtzClT2uTIkHizpa6/xXJmeM0Nh3gVNgiyU
OsJ7QSx1QosPXIVl2bc9EawfyQ89A1DCQ1oKIGSkzEYsAp22bJY9Tf/9Va7D32FDPDMKtUwpsgme
2Q/4elNPuJGwFuLpCC9fY46N+CGESnm8amvQbSOzQoe1VCog5h6pfbLxASkWtq4UQLrcJCwTZ/7R
OgaMYvW031nO995X6qtcvjlXXMWjIABB9eY6UQ87cp85Uqw5iVK2/2c1HkdtafOhouCjlZr6z2j9
vWKjhxnqfhWd4fm+ExXjh3+Cty7TDbtvNOygHWgtd+XC82YfjFnY1SYDV0TrpaSi9x3cubgIRbAM
Sh/1Nh3oFdpVrluAX3kJNr/HFrNc9TF9DQSlV5+7X2SzVKsSW9YcDOs6mQ2PH+KJS/gWfs9cHUe6
q0KdKg6xHkrbsxge4IVyST2mPu52xT1UVJotE8J9DEUEy6YirlrzKL0pTDkAA7ODpHSdxgIAvEYy
2lFPGXAZ8aRrADgEl0QVTxMdKccPv9+3e8Zpw4CZpBjo+mMLJWlFvt8gBy3ptF5dCO7TTwcebEc3
e//Z0Vj6xoB+CoqpFXalfzUc2ti8sjxHUZ+wnCF2xxGNr8A7QSuqhrZ6JScd8C2lJoqRvVzc7uY1
YySqd5En2qAqM5tzPeSZHh7ZbXn1ALhGm4W+omkKvydi/KEbtJkxXazT7nV8BS8FhQj8dar38b/8
YFWroxaKkivZZuVMokjBQXhR7MfR9p8FXT3aGuZEScmP6cQV18oPSfUs6gRRgmW7qiY5U8DrhWPi
SAfJwr/N23SGCw1iWQ4IEGQyqZEd9o1pJrhRepUFaKzAxu9kYV/1H5Fm2zt+TM7lqnLOs4tL11md
so4lQkKcShSJBAv+tA4VdWEDqGh2zDeMPdrNFPMZZmkF2eJWKFRNIMXUodfiyBKWN5vK6RzlhZDg
k53X3J8z7wY6i3wmU7vymPKZNP8Fy6k7RjOq0W/LbIct6o5O8tnEIt9ncQ+nlbD4gMcwL8G/ZN0a
ArB8GBRXV49Z7kq0id/1yXyqkuDjlcUf21cPAySQq6nT20hdzaBJsil0THbTgtHcItzvIx+JkR8w
OplVXlJwyYtrnRCOCj+zNA9FtPj3TXkQyLsr24zVSX39Qpsq2HIH4wvwe4GeLZzFX/aK4jzPE0ue
1vgbOFa/XtsaqiPF5MHLia4PVkfeRiDNh5Zv9uRIkSuRpUFF3EEgMVuj8XvTaHA7C6HQm0gX8apQ
cV8LwpHpO9VOihhEXMPDzq4+pH6i9ds3PUEE3zUAlg3gE0Zhy6iKzsSH8YOT/BaPms7cY9N3RI7d
eXRIrgWgw7MQFrGejL/2cTc1FwBPY9wkUv9hBbtk0mYzwza90M7HkHjryFneFSTPtPEZf72CoiSX
00T2imQnJDnM0DVil1/aieu2DK3fyesEpqmRqKlng45DRjaxJW/835Yb7DWgLqkIobldCiL7l5hS
gM+5vAcOgx+w0BZkS2LBG5h2WsI1vLB/8+A9+uWD/X0pNGlCDJ2pj5vA4MWjlc2OtPNnJD03rwZC
zARg71bXB68VfS8BoQ+Cv4AQ9Dob8rPu/Wu9+yhiGOMAU3zbz4YPO4wJJXdXXakyVtEI5iYLrHZg
9/u3xFfb21P2IT/pyPLVD6nBWut5dYb3v+zz+occJD2TPoDj6v+5r1RyYMqGAWcN+WTP5G5i4XrJ
o9sZJ/OCNsSXP2f5KHJDtB9U0q+V1uoRtu8UWj8lCsEG0/QxOPlMOK5uLbI/tCXEv1gytnNqaGIY
UvzJwtn9OWCNLjwE8snr/jPSwiDg7EkeeL1pspQCkLB2ITWrhSdBFzjz8aDtGvtQ2eToxY71ful9
0R+Bxv8i67zbZC1XvJMCUm2cpUxBhXtAvepWoLRzJvSx+TDxrVGVkEynR2XBD6l7obN4JQoZY1jD
8KiMrbz0YRDjv1vzuz0O9mc0T6mCR6RFWNAhJ0ShE7WXbcWaFxqFAKrtgX+Ng+l5JdoN/IX6JAVn
5ChTmnwyERk6FG3FiaJQceqTkK9rL3dAd1J1xtPOHjPpbXEgmLjC7h8efi07JRbAya60mJaoHRwx
b6P8f7DSkYzW9T0zrkzdl8ujF1NpaIjwSxquNRcxP3+VNhd4tHnz6fEVHUlVvNtMp0UiLDS9GmSl
tTYVOTKgdhljqslWxN4TGSiBy33iwqOJhA5PPj7z/K195325118LB9csJQDTJyDfqhUXeVFmdYjv
KfSzLXcnkMoXtqprvtA0AYKnvBIvoB+WEndShdcKu/3FbS0SAccyg//l4rJgUQyoVQHs6W+eGafb
VRks5L0VTnCX4tKeXB3uyHLFtR5/288fahzPIUghFP7opmL9qXz4f/5PO4HAivYjuQPNlf3JJwve
GhdgWBGr0FXaJcTdAIZH5mLqmXwWDXR0oj1dRMN1Sp44PXyObUdg2MiNcFw6WKVTORcCsYq0ZQL+
gOXI34sKTd5wrl1RcJ8XDH9Fsbr2efLfDZrjO9xxMOk8G03dl+L8CjzELSf/ixgJmOLoWgFVnxec
nqilMv7quHbOxCRt43XoyqDhATzeZWsjrP5xl5G24hN96aFwbjN7Jtdi/uljcM5ju6PQBv6CV56z
G5BP4j1MTmwR77+Va6mIgkcvcFoyImIgd0eRZFZGuU0JsrZEjg+mMPFQ5bM6T0S8A5HJEexe0TfL
oEgGURUnnkDvbQLxntk3LOOp0r5DLtGExt8yKFn4RzXIDhrQ9TJQKE+XeqcaOVq1xGqWnOlLv+kf
ik+WAyPb9JVi7zXTMdtrI/FDKeXwnKgOjn+mwaNyqL4ANwGhYRCxwxZAMHijJHHtt8yxMPMAA/44
fhIkW4KM4tsFHJ//jBBaViyCGPymK5QUBJ1BvsWEqP3MPTrR0n90hOpqZr1smt2MkvBeBosahXQH
oMHsg3qvxNElJWig+pGGT+ZmR0N+upkSZgspzTaL6xmZVFHIrAZOHABOF3IbBY/g8VZLii3b2Lrt
bWojwX4hLYK3MdpAY2dDkrgkQeg5gIbSRCT8giW4PQ3UFsEEXAIw7WXtSTDTobLJc3mAPUo1nr6r
NIgfv82j7F4kd3UVs+mb9AMA+C7k0CbQETtnF57Q8VD4hf/nWD0t+9DuJY0luBNInWzbH41f1JYi
hKErNrsHlnXaEiU4xms9apYVMylE9JGv6U11P9kHLVSEEQVJG6l01i2Azx0YlRuRKLbej6mgf2o4
MG9sU/AQpTfr4weoTRXlTriBiZ1wgwJQkSY+71AnTwwxXlM1JWU9Gsdv6Rtmeg1KgScJ2vAg5wL+
QVtuSwRtn9PSrxf+2sn6pfAdPPFoQGViDQqajIL0MvUDTbf2HhRit+ddxYxaMe/WMBMVZUeCagk7
Icy7rKI4I0Y+wTEA2inzkAph4kBFMSqX3tqC35qucdPVsbD2Y+sNpwJ3hLYrU3L06fqBmFFL8b4V
iFmh7fvNY6XpoDWRUoqs1lyh31gpL51WPIsweiBQQ2zLF9SU4AkbPca9B1/9Qk+UqNcJHV89SFQS
4NBXZBjBDcCuoFVguR9CnkKuF5iCkBgAGuQ9zF+Y8YlnEkK8GhsHih2FMbWgTlQ9AgB2VvX/5PMv
6ly2u+HMPj8MsmXcv2wj0W1PrDCBl6956bzzOMDZejL+ov9buTz/Vdl/rABK+MDibKjyVxRSP3w9
eVNRDVu/nyV3Hj8c7K1/9KXMAEI4nTeK7ukHLCSwlQiFNIplNuA9oAkOalGfKOxKLIXH7CLhp/z7
7b4mQ3AdZu+EjCe854kFFYjyzLss4jl8jwggaF4SNPT0YLGnMByVnCDy8Hi8bDOdRS1YCKB8qAv6
bydrz3yjiVxsLyI/l29HR588bFN+VagyWyTIoUYbEheAF87eOrHlA7ntEK2JFj3wdmn/tEc+XCyX
o6fK5Tr/pmY90aB1GftmGzKqjWPX2YVZ2PXP64S40P+rhuj4Z8H54SuYwH8AhWYnYGvzgPoIvWYX
le+TLOaogkE5gFyIOwLs3MLIkwyG/LZfCz4F/s7jDZ/CDS5OHAztIIaIlvGaMeHTcPv6FSt6logG
1t4wJducKh1x9Q7vhxfNGhTrFUEjAhF58nWjcC0j4wM26u5w1nxXcHWdarPdd6hiWuEINEFJsJl1
RWVG30ko0bzSa1NPTG+yznvU2OdVSMUopT4L+KpRxkXKuwTLXRHxQCiZbhpsT4BNQiwilTm0a2yC
uRdERYhSPFtGoAJifwAWOXf90QnbdWY9xf4BwAJcY6ABiiOooB6/0TO2L4Wud4nuROuHaP0CLzER
127EPw1wSgO9HBD2WSDI1l/4qqJophVSH9JczFSwthXC9qJWtwYVvrrsJNwXzMnWJP9WL9Jd3Mbh
2YYFAKcEuEAbb94VVu6r+Q9J3e5+zLNf8oUZyHraim9jF88oLx6CJfHyEQ2KmvPQX9sI+YS6CmXo
bzYdZnVzW27n/IjEQoewDapqk8ApiaDjc6PWTqHuvxCo0S2b5PA3auP0aDJmVISp2Hzab7jX5lVm
K815lonKBCSUa5ANFsXKIjVkDNx/APK3LEHvMydWn3/aL+qju4KVDGujt1JIhy4lDFzFvSpckBx+
lCyrqp73bWGXlOnVrfvWhwi9xFpQZwWYC4wVnto4qC5GQW26WFINrrfIDAwU1CHW3tZ8aSal0cVe
jGNeBRpoIzbrkwbLnX8JjBGZqi0cn0vcg5nH9HE4RklQl4KIF6W8dMzthq0dWsg0maj/tsr/2sFW
CUzFxLdPG0cVFEn82xQiLOcOR1CeYKxpxfnLoS9cXIPL+Cvd4+Zwryi7PkwFpWFm/iAQlUDpm9kN
MPvY74elNWUK2AKneFFDz+419OsEKUmrfSAJA5n/SMv4HfFVOaiNjrf6X4ruy/aJCtz1CcIs9G0+
6sIa5RwX5Cy0aXygk+Q4XdzHkVRMNRl8mgEOifKf1DNz1Zhw7ApPMde/e9cLFwZslbg7r63e5Id1
mbsiHV1hDNsMZO82BMk+67Khx21nmleM32NlLfcwLGv+FmRCwrWr4McRqcIuaL0PCJwK67H6RMFA
fk+9qMBtMa16rmutI4lt0a6J1jA6gsi59ncbMaCcth4iB50G7GN8W8AJt1tpIBwmBnNHAtmwT2UR
HxNf9kTwiBVVtWB/TTrqi7/Dsoz2npGN+k0ok6nMyPjt0Z++Afn19lCe4oiqI2oqXkt0hF48J/yP
3/jiho1+qa/53nykMv1Citgem/7OXzyRtD1dU83Xg4sy+23lGjJpiudSHi+l4PcpM2shaXyqpAuL
4v6yhQgc7OpvAa5Fpq0KtZBna/IcZvbJLW4/YTeypxBmEHTfQNZ1APnSAWm/Qw7P8VG7G9aBY4Qk
u7IUGAF2oiyQEZcNn402au7jIKI5mqhuTai7Qb0Kcf3ylmVIFs5FWGMS7asUXRVNCBKFxAo0k6pL
e+N4hrwXsFfwCaazw/UK5VIUZN5JoONyR1iHF4rbgAX62L4KUQDMm/SubPQAAuSWqDZTe+mh3P9/
kQdHVzNBwolaODAjGHCsUflf4uppvdU7m8lfLV58O3SGuvoVHF6WhyVb4alavkwstTn2285UcVQf
Jtm/2VCHtLw8Sd6Qg5fzmVfEk40ggFpuuMJjp35tQIsZv2vm1DAq0vog2IRwVskZb0TXw+55ASMl
ODQUEf7llxsh7NreIsIgxaL/T+JRy8LnRMugfhQ+107+nz2K46vPPdMCzcGTWOETzVnvVMycxXfP
hNtHQPfeMekQQrFE9njyeGyzpaWQ9Dg/OFrAmBel9i0HUaQ5+VMfkUpQBljoidO21Pm/1kLKjA3L
/Z+ZvwMtJPcssvnjYDDau1MOLOZ9yMVvQb8s8xTzfkavcELwEWJ10XkLP2v2oNiEgEtrdsW5c9zC
cOfkdLbSGjohAHym5jR6h274cG0NuGFovMjXaESiggIwjUmEIdv3D+c3t1MMBRkE+Pk/RJqb3NBN
vIijNAr2eRobr8BhTtxseh+j4AYAY/Sa0w2+4ZrkS5Y2xuEyB3MYMJrH5XjFhwzgPjw18BSFEwLY
O2kLlr+TTMZNYTxnrjE8uNkjmr7caRWeqDzRPpn08Fe7nzObJgTNnxt/CfqD5lOj7gV1WjMnZzuw
FInvCg0HqFuZC6c8NQtg7QEie3zVEHsGZnfEMAABiJ1fwzHkZOLoiPGVchAQhvhRtDB464qvuSzD
Jg/aSoWMcC3zeNFvTJIDXyBdVZ3K/f/hfHOf97dD9MC8ZNQXoLOvZ/zvzOAwDOpEw5temyvXEXLi
FKGwSYlqS8LaR7/x3NO8/RB2dvdET/ybsoyftyoTKi8dzxcMKd3x4z+BC0bjxKNdb1RxKxaLklG6
mDIV/lohMSYTmhC9nu3o/OnWS54bddmjPSUAK86GRr3NtsJ3sPvELTGzXBz8hVsIi5NMwJYirvph
UD8l/NgWZB7natmSqwGPF/HxuiNNpaqCi8I8uwpWCs1RJqY/qoSCltb3WgYfMInZb6mK0tbWq5i/
IXhnyPOfezbp99CTDiNE6a0Rmaq3V2BB/H84TTyA3BDsL5yd8/esWQHFqgu4bO+TTTmRuTgZx29d
e4IHOBrvk+vdAsL6GTIPHkktuYxQ0pYMyGUXUnj3rwNBuEOQsSLaPXEk2P6nRHs0HkCuH1OxDWek
A+uxE1D9KgHL3N0xHiRy/iuztjxtT7OIZV1A9Ix7hGS0TKl29dNMKkjMiJ3KxQhYy42BZUdOOoO1
7Lc5w616CKgvuLONUfwqFPW3AU3e/44vg2cDJYmxqXDGbItAkTowqBAGp4Y6V060VNvJMbt6nfKN
CmBz/BsGGYp6xgwP8dYHrouk6TjHNn7VxYO8W0eHIRGFmKEKRYRQ2B92qcqXc4Db7IOEgE5m8OiY
xB2VLlh2gounfGKNocknQxpqLii6wCxILe2AeBosoP1TO4E1IflESFiZqP8y+YVkXOSMGRcdMmgt
A18VbZT5g0eYv41N4DSPdLQ5drP8JCEijikHiT2tr0mlE5GTf/OQwa+IbZCHtMP8WmSbWFReWvwK
vUiSA/5lToJYz8K9xO24PSdWBmpNTlzWeIYg8GA/O1EdBwXaJLxYRZjE4QB+aXKAxGVWRYDKnKEa
XJ6T0ngweKdDWpLiA8aFit1aEQpLl7IM1YqlFrp7niUuOhmKd54h4UQFiLZf4gZVtj1oIiJcLmmt
OwnhXCg6AGqH0GVC2FEkvgiQ7EXetmSsH94Zh6wZH3uKh8YRVZQ/nq3K//T6XeGwfK4l5V+yKBtZ
nZNG0PefDsa9yvVnwvRci3OaKyEfcH+ObL76J7Ua+VwLl7yKNP7byQG30WxMprgl6+JaLLMNr2pV
5vAgBurdNHqc4rp6i3hdXHA69zncWSR1KMH8Sc19d+Hoq1BEk8zqWMAEY+qmsNf+x+NkwgYa9QYI
0tLI+OAUSAbo3GJr5BcZOL9vOot7tDDCwXu/lqjT1Hq3FKit5TzmWdPI7e3fabqKcUR3UPRIyG+D
wdKldDEiaNBQLMat9PyGRJhGpVx18gn1SXgK3BaLjvyq/UetJ+k7Ri1qv9bGMnKeLq/840kWaYSY
4MVXwO0NHm9A02WdkIv7KVkvKAMJa8ZYW5gYfnxNLqnbUT/1pdxR9ldquLl06eBFW4BgL6GcZrpq
yi1RMv/r1zCJ0no27rzKiwlr778qOzyK0Kqy2/EpNTixfYNqWlmQpz4+QAkN6bAuAsw7bT+Kcsj/
jRgBOEw6cWnsUFlVXXisdKqqPB27oyECwZbscZ9GDAvpYB0Hc65OsL2dKYZp6l9gBhKNkCmI7iV3
LRLtbNFSR4Z0mLx115Y+ZptSpGvkVFoknAz5Bt7ALuf5dWXKdERAMG+KJ4Az7ZdkpDgdwcvgkYZD
CMIWYolss6wsuYzGeBxSi9hWWWA77aDaFHuuH5RzlAD4joEL6uqqtY/0cLcWwPMy/FNIup2Y3RV8
gfhlWK2GsZTNbshEwtXCZMik8mSTdLkPrAy8HAxomzjk1NjgMR9Ivndb37+iI+lYzhO3qDiFJJTB
gaf9DGiMgMSsS9EIibhm5MEe6GTRuy+WtedYNWoizqAlEwFONeIoR7JptENhF53VI0keqDhdnU8L
9czIwE9ypp6pjW24J+kOkVbqqBRcZO9qjYxeP2oMzLN5FufjPGp3xbxncmEPWcwN0g6muwVcepTX
JBfpA8n7YD3rlEo0RteChSX0roteyHW20+E3y7F4hm28y6Dd27caOVGWinbzzv/EPIcLJtT3v6rf
VWHNMh+JqE08UzunIvaTT3WtZiTRbTSbQ4CR/1IJhjB0aD1XPKj5w6gj59zZAvsCO6BO+RXBksaj
Iaj4eqYFOCZnT7GG6fYSL6YiL/FedOQ2JNr2cE8A9WYUQIDRD0fv+YlE+T40SHWUHFvvpJPIa344
RwhYuwBgUIvwgBrZXeRt+aaIEQSA20wdWzP43KRa/9hgMRprR2Khtzex1bbYt5Sm+wWI8pTH3AnM
TRhsVZY+J5Qit43Ofud6V17sAY61FxKpG5YAdmZkEl1+WwV4NknhCtZBZ3SJBZT07lNXIktc7clK
BGq9fzR9F7z0RzdhxFMFSexzsHMSfkpPASh7goTntpKxQnRH6TkeFk8mbdYT5+Bk19nfqw1jpdeg
GQ/Qg/PKukwucXSCTfQ3or7dbVU3+DDyVMQV18eO7zmm2s46GyPQLv9kPY52jL2nFlkkJ4/LuCB9
GY3PSZ6n2FIFUGFrE+0RqTm2JU5uwdLwkXgJ5xtaY4BBRSwrUj/A9/iATw8Pee5a+8wYA7kL327m
JHrM/EQDGT4c7a2E2Mh5lLtXQgtXcIVKUT6JhhFF9TikDFcMPyma0dlNWOY6o1u7R/qeOvZd/5pi
doYLqOqKE8yuFEXuIaxbDzWIyCjd/0ZojkgfCUhiF/aD2MCmGcBobc2sbVsveVLUXE+aVTt/1E7Z
68OUFljSqlOtNGN0/8GDUeB3yiq/aFYKtHIxBllLjk8agIwe702XaV7qa8paZwGAsICMvTpVAPVe
mtEAlZ/RBgcyigKmcGRkrRSAv3Sc15UOuILn3MwVtMHtFuAO3qchuUolTRV73IBBL9/mP1EuXpmw
OSLsaCuIHd4BXKaMSp0hEum4MxhQXK2EoTAren+49zA88W8D1oJVeCXeSuKZf0SnMt31A65ZHaeL
uSM9obJLb7WbHe3G/tuEgV8lfpyeHpT0WXnpDrDWemlN4y7Qhw6GnDpLuBscNssft/M5cqi8e0fi
hvBozxbkrNjuOoPhgPuY/bU+WmEKrQmAg4/GKR4tYylsO1G/oCgUaPMo9oYR89TMD7E7LuQ39+A6
oS/SqbMA+I/BNryXj/q/02ZQklLwlnQBopC7bM7KuEhatJZ5J6h/WQoEO9wKGLosxy1lPwEtGC/q
D4QyG1Pdo/IbCs8qS8j8xI83hDt7zfC00ly5PO/11a8jKySiNNVPnvIi6oBFajAJfhCamdl7ndd7
izqlfeA5OSvGCSFVkd2G7HEU3ZI9giz4kCaG+lrHgcpYi08Eq4kSAZeDNzZ3UtehuZCeYfIpEaNC
J6Bk8UB9MzMO20cTO213DwOuUFQEayy77NodcbXiCPsM4cx2e3XU1Q6xqfCFTBmahwWjL1FFgqOx
DlU6ivIClnmsEbjcnZHaMO5x7SN1Hkx6lzhQvHs9CCj9F7ugK4WT6ePB5alGPKWPE3KOXauVCpSt
Er4YHsexHuYX2Jwsq9Wqj2NFeaf4bfxCbHD5lzgD/+qFmVeor8he/g/zUTELQJuKbDNs0cgeTh3T
z8RsX2GdOSjx4QgwSOrNxB0/AK7+q92NbJ5jVB0SJEJ/UvwCpdCYURU3HYR167MOmw59KjkCbzjc
YeTIBEN37wYg7TXABsA2V0RigteFCbELtCbn5pcawJ+UjV3bgFQZ6/IS+AlOqYLvtEQkEAKMQ/t3
Y2MAa9dxchQJVrWbMP4NgxeKkVtzTxoSKXW1oesv0URZQpFY/9fFL6SgX+pl/WZucLUVvxV4p/A8
NG5nKObXqtHlb3pGmCbfSRIlSRcqI72DW0ZGMGBmkKO8/LrdjzD+5hXN5T3N+aOLu/Du/FjqUVWa
sioMAC1DTSRz4YaYYIEA7i69mLDFN4lANlC9MK0K9aDRuALv+hhMO+G8sI2wsfXnUDiDbPlNfoSf
2Z7+ckiawK8nWl5hj9vszRs+VrFClNoVEDLUcs13GHtTz/hBIoz2LfAwwBgW9gJehNa0HJHNKXDp
XLnahIrME5z4eKcnbjjokgmgr4HbIyVA0cWW9uv9GqanrvIOwk5nWu++Ay1cgCMPe1yIZNvtmlgd
5DRb2OQQB5IHXKgQ84K5tcPOn9Op9F1YIP40XrGlgxc1W9xrvn1848Zit403QeJinqfOYZVOFqRh
RLw6vDF8Sug/q9XuPhHg68FXqrLM/L2thN3pYo3A7veCXO5pMbNm9lVfp+LxIuuYG2UaP6LwAUAy
t0IZOzvoMtPgbeU4GJcsdrxxXxk80znpm1lser13wWo35zi2HT3NtbTZNEwe9QeVWaV209bd3Eoa
PGwoca3sPFtInwTUrUrDU70BNaDa/My9yTcgBu2eN25cApYyx4gog7mNSDRGGbaRFXtqLxQ9CToW
Ya+AfFxepf0gFAYeLKgZvCfsFIzXYWKPBzeDi4+eCTxAZDVGhMl6BmTQC0yBqwCCoe9GORvgNfWU
GXO9em71XiBrV5hL6QcPr645CbUuc+uUGAoLrW9VR6dRUrXO8tYLufEdap5NNIL+ZO52Si2jBUvq
CFiGms/zvA/xx/qHLHU8dsnUIAdRJ++HztLHuwlSrypmI+LcAIBeCSnOB6ONoanOVqk1ay49vmtD
iLq2OG1dT/s90utn7RhtwI0ElSrBqH0Ocb8mebIS+EwijkUaq+4GbL8uQ3mr6SjsJevrILY/27+5
saNPsVpwSQkltBPAFuwgMtxABDTDds59XQNTw8cBfaMbFQX3oa/7rIHLMWCtDI2+tqBB+j12oEdp
f2MM3e3wC956Vl12K6k4RWmU29KHbT6E37nBoKPq4ZKSnUnfMiH4Kk43cY8nNBYkEpyKbYYkkYAa
IZfTRtKMHLxtc5pA/cVLtxJZZ1v4YOks6uuSsfGHAya2BYA1zEsSBvMQ6W74MF0l6zJnAwpWUdlx
+c0jbW/xKKXw4JdwPdEy346zsoXqWefHnkoPqkEXqMyGC8O7ZjH5MoyoHK/Lz7a/l1WZ/eVPlJme
2IJf6HjJP2tRGVPGk4v71PAwqE6fCN2tEXdVYzjmRb2UjhFN+/BpdsNsIpsDHKBLiHQYI3YsoB5W
v7MIJYCjk/csawDX2aqKSnvmoK5taru5VKzsndxSFLGQ8LdtgywfeRHmriXScpYGdPyeCqMPY1qw
AAFDQaoeyw8dkZFj5RfB3M49GOw7IkpXpSaNzcWVM+w4XxM4DYgNnlbTvg1APzq3h2aFZf/5cdj6
P9z1faVphXjvvNp8GRod8tn2WxkalrIy+SNviLZrH4jLe7Ut7qlxNChMUVFAMErjbqoXVs0Knck6
wNGuyXi0KhD16A2p0y++9yghrVZchv9PTDM7WzTGY7avVfdF2ndhV/LptD59qqJ5JG/yfrzRP+2b
TV1Moj+DZQLU512L3VJ5lLCcNG9WQ/rMgXhCLgibDnz0rduAATDEwVCaj83ykv4H6SQBu7tm3la1
DnnlpzKC8rx8f4WVDE51e22i9h/ICwhdd7dMj9EXUjYbUjzHR+MQWI2J8b27mKlq54LUXFZM+crq
mWnP/ssPQYp3mLYFg9HB+7IvPapPyunEJPRyiRrpkBAI95iIV4x1yMMepuu8LxFUc8bsLFx+JJaC
KdsHj7CwyMf0vMGokSgunnYLwks0aByWB3UNwncD3pq9KJG2JFWx7YNBK8US0X9C46AnDEdCuab+
Jp4204Sz5Ljv50YsSWt824UNChAAZjc7Mb6DIGGVFZ081pk1EPI2sqFRpUQhgQjETY5/WwHSMPWE
ZNsyXbHJVvxPDnDejmRqAjs9Lmj54edmBF6FcJPywp+zafjpp8d9Zq4IrADPnZYAAx0xfXXJwsqe
dRyD5Gtiy+LpvXSvTlF9QMle4BVWHqfwfv1U7dmvpI1rQMQfU2UeY2nRSREM7zkyK0w6Kr973MPl
gttupPUx7+D4sY3DwRVYHt4OvRCRsSFBNcOdzCWQ4TPAYOsxjpvHbQ+o67gnxBYyVLKoaNoD8XyR
UKLW8zj8siiORC9jJofFVadzVQ1HawHGa25GogWCm/F26XM4TG822lgGUYlknncSsqB9575oWVmO
BWXaElF5k6xHnUD44HdeMBvL6dw2BLVoEftgp8RK8/NACsSut3aXRDOoEt4w3U62X/3rYJSWAZCf
Y7iboj0c2N6uApi98T07oGvF/3TpQqAyhi8C670ler5DFmMUKFdiTmLPrV8Mkb18jR1ah1jQSRl0
+9hetpSrc79ejJixAd4LvetTq5RUDas+kdG2r4QrAjOvyjzGiBYL4xl6rgPzRb5sIK54REBYDCFW
089c76mQa9L1p7sKriWS32HDfW0BzK/hD+2scOyAtPGvFEYfMd014VCcxL3c+OR74XdtbyXnlctC
hoDXx++o7FLP77cUWsKqBjN28QNhLYO+O61X4LPSd8nkEHCrGFTzfMNmyANF1VBUGLgIIxO8uSIX
zyikwIPSgF0BpId0mtUY1R1uXo0gw/KVaeIoma4FuxwPJFGfgBed2JLZvgVaSuptza76gBcpJ2OX
aEs7f94bRRzXLjOkvfHck0lTrbRCcUqhyl9DyO8l0fSu3x/jmZleOxTSw3qyTNCV4c8SU06gfyif
DDE98y9vD23eqHL9FbCAq2MvSw65Bjb9Ewr+Sc/6RTtbk9EFTOjHe3PnpBou326iKsKW2NFzHKsI
xqocnrKXPlhoKXSrCl/z4NT6O2apMBlnSa0zDVixUKj4mimnCbixc2kFrikUeTHOpmx3s5RQ669i
cgcEaEU1m8+c8a0ufa/209zfhSyLSJNALw4h5f7Y6EFcEzUz0Dmfzo9vROMz7CsYAnv4SAZyorS5
L3HLW+DSVvrLq1Y92X+q1lgoEupDpRp+0Z76MSSdQk/HgX+O2cKBeQXok4BmH3pZJZowfGCS/ZZ1
e9O3nxDJdvKY2Vw6nvX5Rj8hjobTHvNfh7BHuozlKl6OLFHlvlibyJ7fEgCMGJ9vZXHD4LgCZMWm
qQWikmOa9FD39BzXTFZPBBharCfX7c7fZOksqmakUP61ugcCyKjXBWQoNWI+XBIGH3R8f11jK/Tz
wMBgM+tQIZ7LBK0wULGNh6nEDPfaUF2oMH0ffx0EjmehByckmVBt0URNeESApZ78PYzFBiUD1ald
TCo0Y7ZIGBVjQ1lTiHcOU31TO/Uds8aXrCYczuL1c6apxDzTMadvpfC0MirlvHaH8DhElssYHPTQ
FV5gRT1IG3JOudlsGTkv/Wy0pOIq4kDlfoEbAt6NAJkkoMITjsR5IVHGqje8HChhEEzt19B15va9
ui8FGhaJ3oNuALLY+AHatqYMHnV7YQa7wJ2qXV20fXkbgX/y6+GqnDkudMtm9bQ5pIQ9Gmaw7m4k
Vvme/h+v/S5mHArCrMba4ohkVQUOBISZmWuhgcmjUcoshc5nRii16E41Spfiwa/9+p+pkN3JILJB
aEKqQOUzC5eI5H0SxGIRgUKiuZNF0Y/fRtlPyof4tOVk2PQ9y42hN9uVulBceqykiYFoIM3qRBBb
jpGk43QSh4iqHXLG66ODWX3cS1ZkRPLLL0NeBN4Fuklgnb6q3L8USr4QC3K5nc56AE2RBPtpXjWo
b0hIBdvqfZIA2rAhUdoLYSGylnxffbX7Y8+oLLT8E0fg812xhelv4CLINNKJNigW+HbW2V5WUsyi
ipgNyTUr36LQ5Tf1w9o7wxLcf47gPlre7vkhSi6RisMv+Hvrz8D08Y9S6AVrNpY8iY6h2msp5GYk
UzpS9Afzg1zJaDMRQIv4VqzuTN0teW9vqogxau6SIHqxO0RRQbie8hAFBIMjAPSNa8RFXVJLWW8E
m9CaLL/bPJ1KabzmC0k8KLUi/v0h3E/fBAGjQ0l6GQLpYQsOy7Go2ZCzVjnzaly9UeuqoF9IvSd6
cw+tkYGbRLsHm8Q/NP0byFHOb9ZhK09F/otnb6B1cAS3jKkOJKT6sDI79dxfkJmq1dBNig2/5q0g
HFMDDcTG1eTgUohT4zfI1fwtUdPG16eaKTPC0M+G56Oz7eB0d/s/exF0QjhmVNZMB0vcE7Nluypp
RbFEtfREdZbQfan7oeSqNDy9E7iF02ziy0q2NIi/hqtN+AtDqa54WUb8I2WM/2E/Gzhnm8yPH6qG
n/qATi4vyWmvVaruLWiyMmfXCBcx4JrNHSqv870RieLQlokcE/PA+CV7hvbrON4+BSSvgCg5gCj+
D5S7hIxe4gHCj4ZKAsADJ1VJTZf2Nnvmzvyq5GqYb0qSfkHKw/AtyhWruyYt4pUZtQoRR8pSQNwN
F2kylubcVocqVC7rrg7FAloH7bkXEK6wHIpKSOXorZ6rgt387JYBb75ERNCRgMo4+GhLz3ioHn4c
/TbrtGg+zvuOBLh3Zsxi9PCwVDutetHshPYXKu6yVX4/P74Ni5O5lObWqVD63Du3dMNDR/6TewxJ
q870GBA35tvW+bmymAEhhhhYW2j5pcYX8to1GImBAa5zqTdP+rurbxy7Tf4PtKNfyr/QrTcyqcZN
9hXEcCnxWli14ASjHMR6RDctlaYqr0KN34HCUfQDb7Zf5z8dCGAAb1VWNWaV2DO9cSwQsE/y6VE6
Aa8BUqLy1JpLG9NCboq6aNc6qP0I4vJVTdbUHq7xRsmFhBz9REfEZdKDKixvbVsT/Ix5DFEE8p7i
maddx9O3M1iufr67QJA9JFFVN4aCuPNDPsK46XB0g1Zym+qVfvc1dNM+c4pQMdRUx64K/9TKGD/e
3HzDbE8iDMs/ICNb76IFsQqq2t7kpQlTu9EopkJijQu53qpU4oShUXCSV/2Hsf3rhRfB+xa5ON+F
mAtd6Yi0qf0Mffxk2KKsX+C5ZX/X5L0Jz5odsKlLJloSCaW+ql5dZP4Oirgj/XvbDxDQgLXf+F6Y
JIX3+olHbEoPwhyCeWt54g7h8uQV79ghF/R77garr75Y4ValP4c5zVfw5BcG7T9OFbyDLEhNxIb8
f25sLBxbgTVOBzNLwXbzCu2Sdgos9NoCu/WtZ5FFocsQZWaXCJsFXm8QTV76WqNHkNPR1DSuDPQ5
z8qnf4AHzBQxixId+hfCtgUI1qW2TKzOpVE9y+vW+7k1c2fXdNhRkOq8Yqele6EdPIe4QE89m+Gz
nMW9kszTShAyMb8eSA9pMWHes0mM5pde+bY724xT6fV4n/e49zEhu6Q874BVQNj7G1MK4RUllgx1
Gdg1tFUsIkB20fun0rQtY2n/Rz+Pt8eOFRp4JFDdfdQTvMd7Z0TpVZRJc4iwHZroLPyJo2DBlTyz
mdzafHLCCh7aGRt5BSIVL56EzHhOsIp/ArYpYG7d6cRr4DtAZBjTL5JUAKd0L/bxybkG8KzwTwCF
zWQC19m0WNERRT+mnZ6Om4e4EVB5BDxffoD9wIK3nBoOp6CuU8iLbh+lscmz87BUkMarD+yMETKE
BP2datQtWIBwxsY+UxqI9XSVWY3/ACk4mtebgOUn1wvGZmB8BpbodQxJyWh2gIIFTBCDPk6IdT9Z
dcHZAK5G/oml8JLFSXM8A7n09UISMn+jq5zbrX4MbWrn9QXzGySJyYlTeLQise2wqcsVMPwMENjg
23x4CcHxlz23EwHAzMgXCjqVWsHuHDnXXTzIA6hlAlqUdRSbJIPEaAa+0y8/lguzHOstke7QuECf
VEC0O+U4OGazyZmrd2S8pNwuMdUvLe3iwEqJvPBYrLUf2kMgl5ejiGVXPHh6exbx2PAp2bJ9h72x
jZLVOMfu2kV4iKdD/1bu0rvDcgpRQAAhH4ESP2pghUFuQClHlK9Uuv1XJpteLK3hDVIzjYzy2xPF
0ZSHjmEUMv+ns44/dizsFs8RuevzWl6xGbdaXkNmcVMwMrpLbdJs+j5NqEkrHF4CB7oasbjH0jN8
VBz6vXhnaUdFvuxdq7ptVrZdBOI1s52QbyAxjuO0/RqpmkkZFlzt7sjCPDWaP1bH6MAbUcJBsTJ+
H8UlMoz5tJTRZWK3Ubt4IcpnT/uiyAfFFk3+Olj4UHODjNY5ZcDOUPhQaIfiOHpJaZXBGS30BwrU
H1YuSDZl9gb/SKWwarZQwO2SJD4o5B7OrppGGXJJOR4AGoVTy+2IX6MCxEynwFWN6L5stalTGKEo
FqHrfNcLJ2TrLODOX0cE1ZNKF1ASgqLQd/XTccS6rXY3377/LRsURnqj8/+LZVpeF6CtlbKq9VRc
WNBsyedGpRxcl1vcVBoOlqn9F5muUuK0NMTdx8myrj1MwlzgoncwjdlIKgLRUswREm8wRCx8RBWU
zMjaFS/7aNNe+CFluUcreJfYPUCJiWkw66G8/F/8s6Wr4Wxmp5rVu/o2BnbBKxewhP+To8OIh7Q/
wtxPycDkfzM5m1WstUha67ymBNMuysfC4OpFz1tboKQotji72KXbF8q9luAyiAcknQe8FJmzQaxO
Cf2g9DZInpv6yUbwDyX7b893BrPUp928nXtpVosx56aOujvkI7/5O7EgsgMMqFMUZJQumcWZglR9
zflKMNC9a5pJL86X8BLYBhmKS4HpMzLRCUbCmSUXv+fzopGaGpvKHysJi98f0sTXy/Cj+DpV/s9a
FgA9Jnb2sXLmLUx4/aoVfSXThZVJoy+Ef2fMOhX456OqPyOUMgJhkw7HqIxCWlXA/Ur/lNQa0wQR
zTNXx4q3N94WQnwoAucJfFfyxOKNpQ23WHuM8f99c6mdRtTGhsfIZEAds0hFSgHENJtr8vulvh+5
OjP/28m9PzheUjHRAlIZcJ8Qe3jL4tmVJZAZflyjLjU1K+UFzvJmiUftbW2M9esJ85i5Ec+e7kRL
4M8aXBbGE1EZ0xFOQZfEfZmtg/VR/3M0e4rth6dqurZgyDUZvvkn1UNaz79nwv+yAZwX7jUwBa6a
seb/aC5g9m8lKA4dvU9FOnX/2U22GaSyZ8bh0Qy+NAU5XxuyVl1ExS/+k62UDTAelA3A0xXaKqYV
+rK+cqMCLMTwVLWOTt3JydxL2b/0znRefH3bFVWEESBKtdTBvn6+OvH2hhN5q380usyRmeXdeC5w
cP5UwTDH+gZC3pEAireqbgwkEROMjibEAD5j+XjKCPncBWs9H8AVerSUWcaCUDEtkdfIj52mED4u
UNFCugsdTIxuFEHu7zXsf+quHBanliPuX3q6In+NDfsfFcKnh300oVdHfyrmQcrmnfIapGJr7vGf
o8A4B22IuVJKXC8l0p/OlWCJasWG9Tc8Emya9JSV67OWVaQgS6x/cvREae7vPTmkhRcQVNB5u7lJ
ZIaNHfXWRW6lVOZ/0xmVcqF9ybZC9ioUxAw+uFaEdVL58Lclw5YOdWDPvpnvDRZE6EuIig/GvyMi
K3Ks5GVhVStghvf0zXFshRz+/j8IlEij35inos/HhjnKQHoagxwScahLDQRKHcxztemrtrLvz3JR
xJfGeO32S2DxTSy7u9WMPQHdgV3i/0AI5gsx4atMNj12bp6WKk7PQ3swq2wrWIV5JfV/xDWKYYmJ
jvkcU8QlQByYKW9MLRvDE6KXl103DNo3IT43PhkFgRNZC9BrTff0fGfU20B4r98ct58ZqfyGSX7a
xI25pHq7om4j1duR3UBfBnxkvbft2ye3H8Ht9Ca0xUUDyumYeZM5QpBamZi5e37WiCcgxBJ2jC9K
WxA6HCr2yv7j/CcfKdxFtLn3eOLBhMIL1wI+fCbrSl7hgx2C3X0KabhBL4eGVcYb3Nq0KDuUWyRu
+xsOjKV2W6CtXrAYF82uX7YHnC+05w+fGGrmGV1kJrdgGe9uWjGogqLwfxI8t+aX4xBaJwC++M9/
wTB2M+R4H5dBeODQoChIQwA/rgVVm2XHJaLYSmznPSievGtrIsRaP3+VtyBv75mRkLyrtEfAxiJ9
rNGmsvu1wVv/6znBdsdunZfReakOkLUQuyQGJssyoEIx5V9hyqN8CPdaFKfhFUjOvXxx9+qaqeY/
EbopILCXQB+Q6RrUiZAGbv5TPmvbhA2PIh7mFcaUMeE+B/bkprGAvaVXZdEJikCtO92/1t+W+0n1
nK/uzY2GeDdb+wslQv6s/oqPmE54O1dc3Q+C/geOJlVW0qTwPTscRCvSKapE95dgywMZvflTpTdb
Ayg3+pIgurP41TAXDDMSK9BDPX+aPKp39vm099mgjKYo/UfqMNt0iMjq6m1juYCsg2fS/CFzgooq
3oXoqy0Umqw7Q2dWRfaZfUG0Hm+o7feHwDu5JJSXsZkd8+DpXacwRt1Hf1iSRnllhRopMEBaFWei
DXxNvVPHpse1vZSEnTxktm2Qtu/2pweBws9jOzHOp9v3BuWhHUC7zj3xvnpwCLjEP3lxTXInJE33
ce/Lp/1hDv9qxtHw6EpSEAi0V8sOp/JVwshuWtyCnkIO2BdkFYfYlGEu+RAeZkUotZTsiEXDJYzy
29GUcq4RXJD4WaB/JXetr4MaLzQm8ry+EXIeq900XuhYcQy80LWYBaglaJhr0cIgLMm5pyM8sJDS
AU1WDo+QJH2QRyP5w4QOaA9o/B8Nq78RLkjRm6Iz10Th+rxvK7G0gAAOcOdAtvx8057XI7Nqvl3/
mnq95lFWhBY1ocNJ35fLZmfok0iQZSNOYlpy/UYUxfOCOHXA7oWqgBxGSAEQm9bTs0W5IoYdR8OD
DvlNmWqKCzar+/KuJ86LgiwPbqwGydMRCRXlXXJ2prlrFKrtOd3P1KCBoXhTCFRYcRNeOMiJf62t
ASJRNvIB9Sv09opmvTFuPm2yGmQSwVqYPJRvW/BgJF+mGngpLPbW1eqoGZTgVyTVvp3uPPCkpfQ+
ati9RwUHbcIS0N2fDw/k1R88zC0vm9JcKgU47VJenu3aXsPm/VSjrX28mKvM7bUPCoNePKkqeyfn
tizcEGfPfnZxP3sxEfeWo1lV3u4EKGCpptoqhz2GcyaKAG51uNO522AN7E0IRwSPiGhnfSHv4I/3
A0hNGsLNYUwLIRYtuesdzsUqT4wyvF2UrS4VhYDP7QSSeo5EQgz4pmeLVYFB0wMKNOoCsIrdZ9fu
dfcJmrctdAVFnKVNlTyQT4OpylytL6hQYEiF0Xu+7m0WJaX9ZO3y9+NBwzul8zS2AVga9YubzGHj
C53muvN5jVZBXbLrioWZQWagBib2a9nGM2fIsCAyyPdzn7VwirCZFf45J2VNFyHMjB5Pq0+u0AhB
JCOFCEEgVZZzyQR7aLVDSF9ljEQH3DlbRTIDs8jIAXhMWBWoFMhL3ogd55FM07LFxjfCDQMEplCP
NPMd3JdoyooumfBS58dFfVVkPbZTBeKpoY6DKRjKFvaH7qydbuuc5cwCAeEpbYMoY0GiQAli7uy0
h6hQS8l6kASPKoMRQraGVZXKe4Z5SBZoddmKMHLIKDCK8M3HudsmE5CeYSd7ZVaMW9QHikETj/3l
An7xHpdICr8CZOLrjULdnLPWoabTwYdczaBvnn8etK5qLr4wTzo2nVD0D27t2yVB00BuvrCDalVd
7PEgu+m/Zr5mTerXnvMd5o9T1oXkvn32GUd6cENGH5DzAsyhtoycJnbW1vUTRtXTD5yQluzhZbU8
haelj0Tmqt9BX8A3+3V+znBilvL4A2x1w7DUzIabbv2tl4JNAEaj3RUb7vjUC+bcu7knSDOLQsKq
iTmPmKvi7HMxPfhPVWE8GTHGHX4FFVh2ZGikS/2fVFBS48j9ksRv6oA/3upgTCD24t3OdcC+mRzz
/ZCMRJ2BTPT81oIecywl71txekdGl+YobZiw+Ml2L/0pToTUyDnBzWXW1Ff0TgnDZuUcE+97Td/z
MSwEzVcxqrqZjB3yswgVn8pcjwYqWuXeJTEblZpSejUpNMkw5VfqB8jjasFA3JiUvVvgt5zLTs1k
kYWtFTvqxOX+NCi4EZ8Hg16hzyYwLcvpI+gyoW7YFtrpuWQy3cM3xqhmhN8XNqd1EdOcI1YPyaxk
2Dd65o8Et7V6krSNBvhz51aM5+z57+Xiy5IQQQVb0wcp3U1i3JulyP5QQ3u2pJbKuRtSb8gl3hZA
1sk+4jnNpuDIFRv2t1EdbJtn+n2cIt2QvGoofOn9oEr2SaAQlHIXCUNJ0ini+c5k0U6s9CxZ88QJ
ZiKVt6mYCy8XaXfCDpRZblWn16ncGcCHYdSEL2hFgF1fXP94fjT6egTBHevrI0gcElqCFbXkpXid
uHkbYE7dc59+dMFm/bStzXpwBd0aZ+MPJYObjSyutdMOJFV6Nk4nioSO9Q2Rh/LtmmnxFz9EFB3L
UeXD8iv/O8X/f2aP24U3vBAthmyvPJedDTcq+UF2hl2rebTh2NIhOIVkwKvS+BFmdk2yvSJ2qza6
CJdbKbVLqintnaR+6mG/r0jkFRKMoRzRtXMQ7Yqrk0GmkwkJESXn0vdArnrpOhCvLXgJ3lhEurDw
mpBA3wu42qwvGS3h2PCeZ/hVkFccBBjf29KTPzqGEdfXXG0ItrUrRgVxD2mnTLsDRRc1naEHQ5Bz
bQm/ZwMWusG6pbOWflM4lAEr/sbHJPyHSI13fBQ/VfPF4hnlwYdqdIkh1cJZSE2vfJpBPZzCZkOn
ON1RHBniNUbMPht9L2kGrQqQ5LBbHUDbwS9wOhaA/Qbojdb0L75MKJup0DWBY+OYz5uukOY1ghnC
UYP67fBf0T0cM0QpnhKuKBs0FJBKzIRZvtqxEYxUn4+7Io7vpQ8ERMYgbxSqzNhQvHtJ1CsvcNkP
o90h5gplBY9RMUEXxjJrU3HzXjjA/d05vFtX0PY/ut53Kh9UC57fag+OgDfzyzq3/SEQMsDGYOiH
GFMa6bIA91rVv2fLZf+h3UR3yRcJGaw2jIbPfhf0TsQjkjZCh3iAdSBJAnwIoFYsnU7P6BxWY491
WFUzDipT7NBt2IXLWFjjP1ZwKMt2Y3n1R4j3FQBSzDQw1h7VHP2OHA4I4XFoTTf+lZzMRv0v2Ate
lIPwWLcDHvdfiiAORtmzukCpUpVv28UbyLUEHbHXfDjnXklyf7rewA6mSKwEwJOoMcFHPxtlpEO7
9D6xHea+u63oLF482c64uukKop4AUUOYVKIpjNfxjYmjz0pqbpzYmZNhgNeX7RfKk0a40bh00CQN
cv5JkpH4ABPYJZwKNvkDZwcgoKPYJUBBB9mczz+mISf8Caxyyd+eRf13Jv1OGqcBlum30LGsUnTR
60Z3dT5eCfLUUjY9o6PLG8i0WZy/haMlx/MNUjapWCd8+hKMAwQC9REZRAwh4HlIC2fMYdK7zCNB
9LvgbFQUuesWETsthVUO0PIfpZ0VQDspmkTgNfWbFVL9rQrh5GyY9xs5/Dv97ejZALgCXjNlI7wr
q1+zqN098ThMvyjpGZE+2zDAIzQqmyzGvn4slm7J2jDlKYWXnmdU70Z2y2Evo8rbdPmrHINub/np
eSXZHuxZwK+cfLxzx/pyxBLG5vCfmimczy2oVnua6S3mvAuRXVTqEdQAEp0fQkH6IjuiEKeXJzEp
W24HKjfB6P/367cl+MVdjJC3nZq2uhDMG6xxz1mfI6P3/rMnGKsnvHxnq7NqvTMUknxitbKTwPXJ
33ibCj8q55WGbUBnLRy6GXXJzTtXdNi236a3A9y8gb5AdhGVP+j4HIilnjgnMNlDx4GIkKs/qaHE
6N2Is84yYvnazerj3Qxq2cRDMuwt04PHc6qDymczBmNI1iI65sMe/6TEqoy6Gj+0XXbF4hHDhV17
oh9s2wvjeFvT7WOq3BkaATnFWE7bTYdfZDwDRHlk5hiQxPmTWvwwRDtTcokq+ZLYv/tWP4+lnJR0
1iiwopfOrBY4K2+AoIMqZtxboJ53Bqy+Pelwv/iKRQ4tpUyqTEtogNASAekO/BgyF6I+E3UPBNRy
HF5j70DaK8g734bejBqrfCW+IT4H+yRVJXoyfmENWzie0Qu9rihKMk8QgW5FFXh1JZIw/aOxLwaW
N/Re08y/bkWkYUVsv1TDjkizFq4SHtCSv1KatLY8seihSjPsE10nJVEagSZ4WplgIQ9JMQsLNT8d
HJ91Zkh9Zk308j5dpo9KYQgfYxboRCn2QuwAQt2wtcaDS5AyMml+2YENSykIMKYluYxJZFCO/KO9
TnyGrGQSylqmg4wd8fwH/6I/xNBPDjJQRSzo4/53wctJrT0mqqaNFc+wEXx/PkEJzlf94R4inZeo
QjD1ASAMxaQ0dTPu0CJXHO+6CVkURmaOIEqAovF71zjyxvSGaJaiDHpBYL03k/l2oguqkdm9+0Gu
S6HzmD5P2nLiELmvms5MeueGXF+5gfbmScnz58joPMdq0tzhr9874Wg6yp3HqGopc9DDxj81NQOf
0Q443+KjeNFeorkwRVOCKy+xt/KGe/mHG38LaQ76nj+5diypjLigdx3ZfjPYxvVCK3+WPUAWBDWV
a+IVKaY8WVzzv2rgWwT3GOhUItSjUXRyk0x3VnrDzksYx9FobKlESt2Q6pOgaTLexGgGtoLMvYtx
XcObQEioHq8/r47wg8yYRgdQAkrj737WyAcR+aWzjVQBkuchE523r3NLG1dYgGZpRPcSwxiKxU1i
XtsU2iSc5z0FLrAiXL+BC5s2GMJ9Yn6TUkcN6LJaWIO83IPFkyIhllpFxQZ8XxL9KvdgTYPxFg1s
rqqFI0Eo2TzG+di030uZdMOcSUwSatHdsEkbwL1yrzYFjUFWbHpx3+wLrni8d899oJ0GteVZiW72
VubzjTyWZN86YIax1HSsqGO5Aq+S9RZLacs3y/QZ4tplTNzDRtssK+mjKj/zwalaT8HyahOKuS82
8tGsRM4jfeLwz2ChzAbKtotRXYI5rYsdum+Z4OdIlVLLhvKijak3RBpHqAoSPlOeitv+4B51HyCL
MWTj7LQnyr0J4FO8DCOqFbgXrnzt9xeNEJRxGfbpeegLWbgxXGwuDXmR4tV3gLWhR4dL8bSe8K67
cP0evBvhWbsP6RK6nvGJzLzHbJtL2rapFTk7b4LAotuSaWPw1Oz173rQg5jL52PzBTWvJKn2ZyjG
IgaErx75xPey3L7ySX23ByZpVPMHYNAqPHlidnrr3td6NxmJfoKkNBV2QoGSytI6hbbi7T5fqh1q
/dWcFDif+Z5ImJpXFX6NBlKUWA1v6ab8iCM25DKa9PfdhDyMeWtmgXqJlvQ+yQdERDTiQq/Vt7N5
4S1MowKISu49LZWNdGORbg7UDPTxzkPyK8doKj/4KyCuD9yauWMkMarQCb9NZBEHnYUIrmM83X88
avCpdhMnp9pXXTBDJhj8o3qlUSt+2CTLTMydXw+CT7z0+wwJ5DbxOf6P5Bp+s4c3XLtSekjFtuzD
f6DU3vK+UW8uYdyEVBsNLYW4EymAW2qfXo6Ha9gFuLORXWzitLUVNi/XRB56XIWX71GrkYdS1PPM
1IXruXksTSx9iS5xSjXcOMB7FstrbWG+jaF3gtgl3u+w/HyIANQJxsxE1ynQQepOWa0o8ERjecBb
lLmVyuDpjPWVXfpAjRJ7ziZK4NqE2utJRzXXJAiSI+38oclkOvB/n8c0PKhDl63cOrLuFSFbFykk
Wr+OLfKW7n9PODAwCltaa3HCnr0CaXtl93CPAl2LG4lMyBY7MquJa8jLSBdR4MqCHh4w74bPDDP2
z2FeToxVS8TTasNWGYF5ExCX0Vi1PQx6BPcoYu5yoFSaBkyvinh/j3ipzNKCRVI/z6aaWj6R4uc0
kfpJRnjkv6y+1vR4WDf6rlSuKDvExJh75BpoyifciS/gumHgoMZqiEw+yMBpxjER+9nPO2v7jy1p
DDnUJl2HoBYegMA4Cack6VUnz9IhMS8IGuOPRXHhGRv98lNbWs5teCXv5JNoI7GyJHH3fznVhJVD
uh2eO0q7GsaBqEABMRzsGsQBHIXsAX27vEymAlcJqFkaiSqUi/MgbwbWsw/60XB12/oindLBTWzc
Kccf8EhKYoSar10ooCOYjvZZGepocpVQ333Rjd5UB5yHBIS6k+vECTfzcAgVAmGXsdyZMmMua8MQ
+akJZfiDbSwCLGrOmrcAi4C44+r28Jmn7CIvnsAQHm4mB/NEcLsmCsI8fQMn/bj+lFLuo7nteayW
nBWPQXZjN/bL8+LZhBoGk7Ze0mlcsEFlfpCk4NP3KavaxduWj7zQOygbpadIQKC9/qZfHxBbMPk8
KD+ZfdMoXTj2dzQZHZgA03CR4cgEVThSpakYRLXlHttYLEIajIQS58KF9DUYlfapp/Ltt9I/5/dc
4PzjQhFLOpNcg9pG9WAyWcBkpFgtlJIQv3LF0PWjiHMvWlQjIHrOuOL35FdGtkVIz0wqmw1H2WGx
ypKIb8YnB9limLNZpby8ffIrA2XkTLWV04+p6XSt8exVLzEUa3+xf/tmmfj4OezXZnlEQhzEDzq9
EHyqVe196F6vY375LgTfcyLjzSRG/2Xn1BGGVCzjIZx6yqZbWevhpmDTU60PoUVX6zXmHykLuwoF
fLTrtqwoM2XTMbo0CV1p2T2A3F/UFawGm0XpwqiKDVqFjYYzbFxfv671ML58C4g0XW6hSbevndfm
LCRjuaSOB179F2PQKgNjlUydBxHBYTeOWFZ82uz9CGP0x2M1FcgZ2v8+mil/P9PsH5tKH9iyZ4Fs
lfmycSzBdm0yMC77z1boWOQwtRVwpGU8pqRT1V3LDVNUBlyBKfhpBCQ9KNzl1itCndDshM9Wzh4y
lw80152lZ5tezWR+MwE811Go/Fm0sfRntgiDCd5bAv22h7zuOv9QjGso+AnOv4RYQNK+I7Xt0OI1
fAGsVNk8ZPNSxOz33QmIFJdMUhhYi+BWGzTOUYlyt2H7ttdLI/A9JiI+3w0YQOt03Q+LGIWkFx6W
gUPLQHfNxrmTwdA4LDODwIDUGX6OqNCFbKNYkcjGLiLTbDGevtoeMFjkZloFX8tqiqpbvTt7zcLC
Z8ehNTdfhTck0g+frMvM15iQWsvOI5yCYaNvTDIwvU1CSAmRnFkTP/lwd7+UYv+xMRMSt0FqhQCb
/tZmKUB1qYoTmZ1Yca8J037stsCk9JqAPgfkGNiQnHytJeGKXL9tPFeoekKA2jeyyqRJD0gFTTH6
BrHYAwesIWb9c9JQrtR05/kbUXY/5KEr2X95MwbZtYFdzX3iwzIkk/w105fA8Csdwt5EwTTZ1VTd
Gk3ygsvunLtF3EU36EJltx4y38nAwqX1GOIhpGTuY/JiFvbsDvp19ekWrJIlhgvbmLr91BC/blsX
zxHtkw7FqBn5meimKwE/drVvr/A04Jiwulb3fLJwMP0pYts2spySFRwWzPIdG9FFgoQo7E04nV1x
wI3JSQS97yI/B05GqwUoNMiFynvKdcOQnogbmSIa2t3CZmvDrkDhZ8ouqsu3qG7nN01sjlLRI2IP
g3773v6WCDF+tRIh6pXaIe24MvwK+qGNvIUv8vH/JH0OWyJQvTRIeDDrjA6DyjtpbjdoQYTT42X5
fpJP+tZyE54leM9wDVBiogaAJATADrCHkulOrqHVdCbB9mbQ5GR54FayPLBkeizzaLAgFRsLDtoN
fWz+Qkrp4RLY+LdoOXFDBlkd7n5SJkBq8n7NBlfN8tTpGMJmz3ingsZ6xHr+1QHyGJiR52Ws9miG
nT7atjLOSmh2HfTprorGF3cGR6yyn1q+c41Q7Pud6/NSkbPtod0O8D3Sxd15YA9Kb5ZVQTvYzWlQ
C9LcCPnaKMnJKfnUAitrCTygOdAdg6TvgoBzXw1NDcWe8M0GQ3r/pxVF4qJQPF853JygOV/Zxk7Q
QJggNQqcd5VB0OMcp9R576i8aHhvHMix6Ce/Gk1Eq1MNAl2jrEFGCqhprWptEbUx5XOMmcZVBxiB
RKBP8bEOGjXF/DHT+zW9dschz0ZObjvkMoL62Jn9x1u2tUY+QfFK9xQazfSsAFPY5Wy4+ftYb7ys
kzGh0ZnrDqUBC8gWiPMZN5PCU7YOY2ze5YtzKH/Awg1tATIqspmv429GIypYDyG7rnqSmE8wpO9U
4ktXDMHmsXzyN/0X3zg+dzHMaFQmpXiEAdPQXTv9tPrGs/D0t1KpD9Q+fMswNjK1U5I26LJWQf6/
0KhiGiXQR/TbIZhTi1fvpteObCKe3eva+WbZZNgKvQI+jlOXhCkxEutSx17GewSAU3N45nizuSHR
B2QcG9g58OqSVA9vFIUQhBxhhskf1sOZqKPEo9pmpx+/jzOfd7hdApaphw0NSljskT273dvogasQ
ycnTW1DfUFugERaCAHaJfMoWcm7ptLfbYq16WjW/Q0IIUzLaK+T30NaNZv1Dx7QWGkeNyACSbbFF
SXRXU1s2QfGE8MP9VNlxdMBKISjw0hskdnYAHQPx0o4aOxsuRDXF1MuCLgFGCU0QhGwzeSIMhdIl
j5gLF44tvY0HacKPWisJP00GNn5IVndS2o9bQEj31QR9R0i3UXG8K70ZLJ0zRasRid7ahCIj6jXN
G94k79NNqH21qPWWtF3ysbLWAN3Vw3p3Vs4aQxeI/VeRbRS/RwbidPNln/my/+WJcoEZGtXokNSX
VZjvypQO96MjgcLeRpnaFDT4m0AR9x71xYUGlcej/1kTBQ7nwdXO+8MTNESY7oEN9TNuy1n53L3o
GvBS5V7BH6gsINtASHmaUZGpIhSuuO7bogIJ70e99IAGe+WVDIpqu1216tjbvOZIstCCfK5w2FeP
L+R66YMC8HQDvxSTyk4l7T3AuSwfn9sxFO2YjiVhXWnZ0PiuiVxE+cL5BBBjZKW7AJ1cLLr0HjV5
R2F2IrgTvQvh3huz7O/y/GCJn+YZXMKQsCQsQ+6PgMCeRZfN/g8xa57BiOWXd7cMnrVlhElEt3qc
OUt66fDaJYitSqEqachWCHxyBce0Kn3yenHXtUzgebYCkFKpEVyPUQ1B6vC4UvjR6PZk5hvYRzIS
VT2pgAfF/8bXYkeBTEEwgqayq72x+ccxTxlETOzCP2RWbfWSk2wNLXryAWaYC5HmdlTeyU3w/IWc
cX8xp9KHt7w4pTC9VNBmDBrd4jpU5eCTB2Xcvz5q7bWEZRlGSEp2VF7KZ7YK+sq5D/l24/8Rx+uy
O/q5WlbsOyP9sgx68h44IRVkoM7kSfBm0gDw+J0YcvER/0H1ORASaBL+TDwoAE/8gTVZZr9hY1Ab
GT+SlwZIcoxYWNZUg//Y3tknCKv+j0IbcQT3Ullw1XgjTBff2HbOzS+PYQgLKQHtW9OI5EOtthMN
40RSySUrsgh1KMTTCf9lYV+IeM7Kre3RvYUpxW21JqoJmcSTo1qKnfoTA7pWUuJL8kmvS8vls/NF
DjGqGdDDvDjfW+DjaOxcCtzwCvi6j3s0NROptNteiCpEptAqLaIiPAvMZ6g63dmadYPnPqBapsvI
OuASURgLyG3Il784nPASYLo8WUIIYVMm8+paoasxy9EUDiE85DVbBhmq6DY3enVGGX+pjrTPeFPG
ikD/x0r5cOsZH5CXYLtX+76u4ix42fVSRuXsNYtKiIsuwgC9Qa2ousnsqKkc2nwounMQ7jkBGo2o
MKFYVGNhSQuh34ifeERDv+ONOmKLXgRzH3R6NYxAgln/mvUCKf0i6Ar5IE30lYJQrnfJ8Uy1P+Ao
bmlj7rBj/jLKVmsQqcPaQBGCH/w93zDzb5C2FqYKx5vtsCAfAHLx0nvYVijnYI6/CrneO3XkLWBI
194riyOVQyCvmz3IBLdY/9L0rragWfc0iUj1Qietx+EU3c2XfteH/PzAb8xQls1H1Ih/NousxkSc
GKtM7mkBfO42P93sQrz8Ta18TtbjGRDKkJIIF/v6xoHXAxLTGJrB/aWdvya4Tcry4J0m328in8di
kGR+2qvFFuLOo0bDRIembLe0FFzi53eTOrqiWNfhqpGaKI7MCn8qpMBifrOWoJmtjp7gc2bcVhSm
bXnQTn6klbXckEY37jC2uCwbXE1qBQni7f8bUdJ1iYk/JZS3kxTcjlXF0BMCqkbcO6KAcANdH6Oy
AXXdrAlOPxaw8DgIXIjpI8KBBMDj/kq71MQFiWrt07Tzb1HAqcadx6wVilKt+NCUignTgb44lIgy
tUP5FxbpmebSVakWClsNi7xUgDtlJ1BzD0ws/oahejct2rWXwDOskUhJ8HVYGo1ZD0ZOYMyeO0vj
5j3SvS1gNVA/UYiqL4Dd37Hxco5OUbwBti7kEorCNEbJxYwsQ+/KGylOuqzRfSYnfjXvSGpY568V
pF3J/yKN8+VTwBFqSGj6fVm7gbv0kAQ7FnU5AG8qUfEBcAXg30DdIJk0jQ381PFKq1eBIl7Ys8nH
FvTb9RyiIkHev7Lxb37VwslmgTTz0xCJSY+mEqF2BwCAfvWAa37UOihY2RlrMqETrZzvZrKcWvCS
ExpdVEZuxnEymuy/os4fpLaGaCzqv0p1xI2LXhLjj//q9DutHbp+K3vbYWqF/bnKpKtuuEXaV8O6
k4V6l6kMG+yx30zY5gqyPPKeDEnJOtuPcNPpTnlvnubFwZ9vnxgC4Uj2Gv/FKt65kkhpANazYdN2
x5JsW/XhpLPT696c64LiANRTUeEJXklz2zrlrowb+5+HsuCedZ7YDnAqtfg358p2a8CZZubntNdk
mWiPRIj8WEXGzu4CCSoOzN0U23Xz44A6rIQIuUEk60DdRaWMoj/7oWao8gfkNbkIWJeo18Osrdy7
P3rqjkwA8+tXguFDnmC0mE+jpBeIhBg7zHRSuyOw5R9W90E+tWgiuUBaURLIa70Zp9Mc+F7tlm2Z
Lv7FAPbIzLos9EO3K5pIpseOBg5Fs0iFcs3IH1qs0ak1HAT8SrMlZyNw/6wbjxlccsV+XdzVH2qm
V65ZL9DWbWRz2eLjeA4LhIfCm8UfsEOqtBUkYjYgMIhkFA9iFoAYkWRQFb/mdYGlXFXArostu7vo
gft2ROIKL3n9tmVy4qMfXW8vZRG9PQ8bUzL6R4bmR1X9Sy2qJoqCyajEf08CXzmflyzYROLCdaSc
/cE94uSUimDrrRsNUZPdLafy0qpK8rYmx/dzGhk25AzU+7UO0/eMw0lkc8SWwv2HcjJgPcKmm4Bj
r/iFWu9mfY92Zq0nEeG4r829K0zbsmz9oKmn59SXPBKUJRUXd22F50pCk3cFHtXZ0a0h2ujqjTaC
MfWP+Tvm70uH8QHwyVIfbSxK5k4mkQGRAyQS8pB6bdcrus12sG1HGaSEKz9xIpSs8VVN6Vn0ePmO
NlKwoEvHbsUvBg953w1PW4WLzcVhDnnA/DddyASB9qCtluSPLHVzkxWXsDdxE7/SS4fL4D/dNpoW
mmL1vhi9njCywWvXOrtyEwLtgwRAHgB9z+/Bbpj+vZxvvU5Dxg/lhQ+TbVIDT98S1yaL5QHb7xyZ
YM4023SO/teitXhglheXeU9HprWIk6XjEptoSmmtLiysgXh5FLZnHhayoukI9o9jSzOUnehQ9iEp
gkDf7fYrDviJUlO5kYK7aF5mfd+oSBHXxLyLzkLrI78shu8SzqDJsvHi51fKuAyHO9llFzZJfUh1
VQEAbjyAY4fFKJXdMZ2dUj0b6RcBeokEA510JlZxH0TSogr8l+LaFkse+FYqGiRmYEKecjsc1sDt
Rw3jwiPeQkeJyr+6S/++KIzLeqjEZFC+Z3i38G5DcAEYbtbOCf/v2aqicI0jyjjDSj9Vf1dPOu4o
eNuQEzMWAgrbeFQeAx+qjUls/S19yyJdUcyngC+3wJ3N4ah99XLi+sBG+wW8J0PXHA/2WqWOiBLq
tV55lyE5LHrmEZ5w5LxFpebmDJ8KrbrQ4uWjcMkUzs0bG74kda/mSg3epTB8HGx1wabuw9Io2ivf
16Ea0zasTMlBn2TzdsmzQhxigLHKlE/9bzg476ayveF23mIGZdriZvW1DkzbLriT80RD+D2suT0S
X8yRXSSDhnt9OWSGkv/9iqzIAiXH9EzfSTONaiYUxFxZUh8aeNNTGyjho1dHW4QAL2ZnUVsTvXuY
NfKb2FmqumK07SkKzkIv1mQS59XbnimCJU8RRbIk2tguJmInrQaY6R9r61prE4nsxfENZj0VgKei
qb9UmEeQ9Wl2cD4Rhd29Dj6VuZwKuzSpI7p6QvJdulVQL4P0b2CPNoMtIaB83DUiTkekhbRUoa6d
cjTiBnczIFMkCwp+FadoNjqkjrlCHCt0exieXQ3v/WvpOogjXtNxKuWayEL8+004DOxZa4vLMfaq
dlQ0ZaQPJi3HQlLFJMYmz7jkzWf+/swCH1gyhq/s03mQFGOCAPRiwHiE6OIoa7IzqMIvqv3EJUfX
9Qup9Aa7jSJfGEkTrrgRyO3EM+KRgSM23qBXGDZmsKYcYtN9uBBcK9Jj3LHdL/uQJVQ25wC3lK7Q
v4aTjPbA8d7vq3M3J5QItWOJRXXDHYRwatJI1CH28sxZOQVyIdCV5ejmQXKXdw/OZTSf5E6NBWev
Sh6uVK5AmprqdRHBvM2We7IBzp7qhZo+VLzzlC56WocoK4dnwBtETzzFjjfoKqVG6Ui/dMI9tVGX
X2AHTQtR3sJVPVmCb5QPPA837KKazJqf56woVrA91UMSINun2BzTEYzbiq1+YPbW8Ta+L0XvFTuT
HCRNjzmthdDkyJ5eDZtekxwe+BJ0MUS+Zjq9MpH6SvRJZTVH6nqRRYOQVc3F9S7UpjaUBADhWaLh
BBCMqwnvUkxCyTQLfcE+eecByhkw5N8yC/1SGm8jkftbJPWCS+8p2vZwoSUHg+lEfoC7LcoqkXh6
3DT3mJFkOQDQ3cUMI+YlHTGHEbI6e3w2eehPMK4+EWRLyPuuzJyMkMlKTgjFQ2IZKT2wT1JuEdPm
q/xFzhvJ3ZbFeuf3sp4pT9JMboxnz7AVTYQPcynT+ffnrInp3gnBJZh9WjcB+jqOe1iH1Y2jLhQM
kGqEjobmFYRUu8T6LdgchZT0yUCxFc0HXSL3eohEH8MUUB7jkRJcZY7b7hrAOnd26vZo/Cag4Fqt
j0yiStpycp//tYOxvapHc3dTb7n+Ct/O0aYsr9pZeeYtVJml/A/Nc1E3zcppAXR4zkx6dIflrHDc
HN3SceIRKI3x3BNOkwegQPftHPmOpMno15lzkO/vUV47cMJeAQl7q5MzbtpKW5/nv44QOaySbOy2
vJYADBAMTfZa6l7PdRTTPZYyKsn6IVf6VMpW3ZhUJp56yp3UO6r+tZcs/kiBTAs+c4y2stb8/Hek
l9IgDgMEXkxglB08A5JtSf+w7K/7I2rGp/u8RlVMZ1ZjhfBvUawZZh8K3VBqB/xZbekdpBYKtSVj
DxqIHgh/EnROX2okiZclTuRfemwYuVEbd1jCtmltON/VV4e7pnOphHYC5I9Dpu7Gzwx882xvoQTQ
lDGRbmsaFnUGsR2Wzg9sFTM4AuYO/mGTour8h7h9qTZeT5+85SjUYju70Ns4MsTTdy6EzXIkyRZe
rIj+Az+Ria/DRT90+IhHdimlV5SJkvu5JaANIWr74Y3tZ1MIRLipv4bLFiEpXJAmXev/9yw6vDdt
UGjcKzWrjvOH5Y6DJHpdpuiif+xp69qxGrOJQyfIOBlR0M6gbVg7bx6a5VGzT18BOmZJWwougI8N
F4chnQIqsBpoLkYAidgAxxGnIqhsXfaZTlyYriR3flo9S1CNVyDuFRMPYwVLHwYIKT4HUZKE3KLr
WrtMAY4uzKBg/zIuazA2jpRjsXESkLWVgQ43u/f3eO0OYlZT2yBpAutLrLFqA+PuYHfeVag+CCDA
FMQbQzaI+wUTSqAc2/uYnzd5gdXRncwTiYXVEz2Ag+jt/fvWbSM8Sc4YIZ4o5N17AvReVVxe1mTB
WK9Q88dpEeoe9j4+dY4NpcrkPKfnPQVPMaqIOUjRhixZwAkbeHslWislCcC5kbY+twY3LnCJyAnY
CnaETxO873jCiuVZvTXTqLthTDywZdfYXKsh4nkOQ7u4gTQCXDDhSFrWKupn8PdI0fyXTgSPdyRo
ZMkurflv7R6+p9IG/OTmM5f6vainPK+oW2KnbE7/Et0QwZWeRaB12khCPI9vZPMB8pLYhlulmSKy
uB2jyk5vtiPhX/aWCn9VHWV7gIbgQud4U7fbO5iv9pOn/D7XcKh1g1Tj5TynsNHJ27ndahYcKuEb
5ozQlNrPKEZGbWr2A4hFjqP0+yuCma3DiaFibM/7L78pEbrjCMKqihPMH1+pxRtFsLYMIZUhqp7S
9pDU8FMz6E7gURE4MvfwTsqTeMtFolOIPOLcCwxTfoBCj6kJJKtKxhsLOhRSUcn8+77FLes9iDX/
ArGXIPEH4P8k92KJd+7xtZ5k+Ekaik2psPuYVeIO9vJILtW755pbU9crmSECigHVAximz6xHYwz3
PRoyVdy0NA8eNNJlzYQDuiVQt2GV40PLFEpZGPZEaca+cgn8KWbXNc2yvnq2SYclaSHZdMxbxg++
XlraM9Sra8V7y6C40Vo1ORToM1QNejYVJ8RifmNA6Ybg8yDLRNy0HsUpSZlMwXzIsPq2je/0fJHj
3KhDSEIc7wlkl++xM239Pu0db3G9vXbfzza2HiLfaLpZf8vqUXc0chhQkOnAxMttitMRr+Rerk+0
78k2LAebQst9KmRp9zMc1e5zthlg5YWsOSu4CAR9cbYOyY0W/NOnEK8sYegMeyXSSc0kGX/wH2Hk
teVyglLG2o2FX58XOvSlttkHOlEE9QrG6AJV41XccDOk7v7ag2rfqF3/DYiZ12ZFEpGaf5pdeT18
g2drE1Cd+VqxwZzZshtaTZy4ooX5vNm75rqeXdfaRuGOO3jcz6P6fjL5hkK2ByAiPhZ/Dd1hDMqv
ZPYaKpbvb70Wk19cLomTQdTBpeYBZCca4yWu99TaQPnQnjXJVyh2K23mEdgV4aBskEtvJDdu5yYo
DA1cfV/w9zVbSQ8ugHYxlHPMazQuyZzdw+BdbKujW8rGegifo3fGN09Cibdwd+7g7ULGo/qlsHJY
WPBRMvp4tKMZlFvN0HCDaMv1TRB7/xsaXd5s7QXqaD2exBi7MPi4FDhvhlF60RCNXvWAVjQ03FPI
L/CtF8we9Ai7M+yufpK5iyh4slnbw3uZlAJWxQFeFJb+qjSmpFMp51h8Q2MPv5X/jP3GPuk0NU9M
wmUDBMY1IMQxWOgJ3+bJVQHxClGPD4lH7geQnxAZDUbkTu66MUG9NMZ/vQiKYckDVdesL7QE9btJ
GdsLgYk+n9chZz3L/uvjqR0A4Po5uLF2BwG31hN3Z7KLaRVLZWBKLF05UnNZ34U6q174qHqPtp4L
miiW2hsPBmFSULv3JIwjeU2X3LLUeWlsSjWh7gN129EQyYaQQloM/0oUXt5UVJphvWFPIQglUy8S
nzgFjuOFVE/TWYStPMRh0N4tOJi351Aac7ZWYYJoaaHLBvgUDdopGDpB39Pb+P18YzFmOqmjtqRm
Lo6W5RC0SkfSS6E6R46r/MtYuFHz+/PzCGIOtLhdfoGUUxllftr6mHnRW4R0/xkZ/yMJKpKLhFJh
XiBld0Gng/itLw9zIjM8AwJxzniiES1krxstA6hk5+QMzkDaL9ffnqDlgBei37cfkGHtJKOFkc9M
HF+z+IrM50dT5V7NuIBseqDoE1VC9FN4Wk2rxFJfPCDtGgCHtRrhsYtq+5es+y/Njl8xDdrEmtX0
DrrwEGMKJRh94Q6WiXusYABf5h8HsFYzm99NxEzJZuaDxTVGpQmxm0J/DVYI49nxeCg4piZRN4JL
pXLnOqN+3lMb6z+mR3Em30QAJ7ZXvVIxJCaU4RZ1N87FOag5bWPYtXrGwFBGqIF+g3sHVP219sX6
USkueCLQHN17DlMN6Z4bZ5DW+ZpquZYdR5KxsCg1iovr77/H+4ssQCP3lDfTjzX0T5LHa344FbUm
VeVSEGcuVoilVIbok7/rbNL0+EUBUc2sS567Yf+2AXf46T/8dv4KsB/ciexajvwIWCALmLQz+OGQ
fBIzVTbHXI6ThVenZjvLixNBEnufc4yEu0aewrkDmYqKCpz+pUJBfjjnLdVyJudgkqTU1jYTiuEW
grws7E+nGzpq2aW2qoZMclggC2t42ESrNOzpuUw6+ZBWKxJ9owGz04ue6mpZyhv+ikVnqdIrPGWT
rqNiAa5dHPATmN90iry7DSN0IwXbnY8Esn3rfCqQPkyzufkDD4ypO8pv+1yvLpL8ZNdanbMgttFb
blxXwcRxomJzTCthqX7gXBGwStv48tgC6u78ygJ9cBwLWdl2AP5I4NvLfRawS4CSwArNXQcc5pjL
X1lcZL2KBGsxqyuhUjKk3fB9fA4twjVH36mS2dXoeqF1VPNjj0866RQwVUoNdweXYi/LLr+9Ydj2
Q1LcRPzsS0OZZnZ0hWlZC4blvdg76YAEaYU9zIFKqaT7w5GNnfZ8rQx8i10Mz3QfMJTOks8EQ9Ko
J0/4L0aY2gaFEufTDzqwBPpH1LBqBV+xfgQxaE0q5GNXg/RBiqQhUBQRkMlRh99cajgxrZTLHmSa
9WxWEOcJ7zmyRuuAsHxvnQrmuTHIPlWqtOjH8S5s5HUbwQ1YfCeKgQgP3U0EikFxWejd6Ug1aIJR
m3SKe1Vz2LcJNDnZNrVlxb5M/+cvEMwQS0pFztTDHpTAx16JfNkxlDBDp0hTHBqRQCrH9BldGvW3
0eb0cKlU5AtbQJZUra3Fvnp41fwnRi0naE6OHcXAqhVVMh59HukiMTZwIaZNLNN36tlXgdHXe9W6
vCvVBvM/JT8jg+/z8a9ytxMy0Rn222gnj3I6M0h917LPSnTQwIJfR+2OR/bxIg88lNJ0h6kLlFDj
owBCZ50lhSs9Dhx38aNAkYcJJxWvzg9Cu9NWgjR9AEphw+1ZwXISGMqWboJt/m8nI2lN8T8ceWut
ZFRDrmR6cieZCUlpKNPomH68UzDqhhVuZOFWS4til7uxiB92DnVQiIvbbW/MnKCc3hckiWzHmIKQ
CLvXWg84X8D+j7VASMlKSYfkcoOuXm+2CuT7L43KKpbl/aqf13qmWqtt+Bx7Se5sSsBDAFUlGyMt
M/GOu0ZUx1XfufyIOrkO2poCQ/Wc/iulw7b94K+ga8zdKBc7Mzf5CG0Vu7hNQh1wzdP47dh8mFwx
0KpYOym7Acl3r2Y7vv0PQjYHjoeR0uhu2IVr9wiDCWDd89zZ3hXo4gr7ftA4ZHBxCP25B20+cy2Z
vDxrGhIFhC8qMA/CUX3JEao3LKgllqorIPgydOibU6g5hB8yVTDbu6fc2RZYe45rkRm2+ncsd4ht
wbvBDB1FExTxpcvLJrk+Pj3BbYfiWZwJelTP3D0EWTDe7dFBzIxtCKa+XbqLpkCaw2uW9q/ILvNy
na3J3hqWxZPQ/0BAjO53pp4Brg+J02oFJlLFY4LCDT/J9thHRzFC52UiqwhBbOK4pxsUGW0mrRaI
hNpL1mgU7kE/T4E9+wF3sjTQDCp00e+PLrQyyolUnh3R1uqEZGTVmquegu0A2urqJEppGEQWsbPU
EmJ6gtpoY8/IZ4vmaNsFR7wpwuXUlmLF8GAXI6ufsxSyv1/g9rIFkvretQs+JY0kcnjOZ1/BR03L
bXMQeno1+XV9+vh+09R23yPPTTt85ObMFQRDICTv6/FBB3m2YXpIuDInU2cvhiu3sXSXNpyUT3Gi
GkN7p5bvRToOStbFhA1oTNv4SP3KSiCXfYS9MEaWOvZdo//w7TJ4WZHoTHiFYRvQhpihOFbkNP0Z
rqa6WOUW8C2e0ZUiHROfewyZEKL4c01LIq7SEv/LQccEOomNxQwvns3yG4x6tnTpS4j4rSYnIP0t
gA2+BP+SbjIcPSlRxNGUq4hWIJ8PIqIuCaj8qnNAI57RYguM3uhp4vO4O7Hj0ZbMRdjZmnqerlap
fl0pYDZb/34mS5xgKCDoWoN67qDt5yeGTqBHXnn01Jjc+8qQfvF5Reyyf4UdKfdVqqi8VQkITMdy
gds2/DwvswyGVRxPuuKYpXUTHzqmmOauaCgajp6MGlm/fzHaiU60XzciVU6oFVJamFJLpE278twx
s0E9HQ882olH+1ZTFc22E14oycTKNxyEQAJnpEHW/GNsHKlbC69baQTGe2WeesBgKMCBjxlhsoPR
E2tduCgb701FWynHaTDx27H0Efe1LEiKdNHYZUzWeAfYBPqJKWahctkzr3GowtCM6Aj+U4E41jYs
mpfNUdJdFrPHnh3yFdERphG0S2cpOGU5nmhSBGWElpEcYGLqeZlVSp93EVdj3RYMznOyHHMH7BR2
tEMi/EGhEcly8jhAT0V0jjS2PslERx+YK7fBJ+EZoA2FVQksJARKW/bnQG8I58TGpp5NpXn8oigs
ME4CKcTfpJhzhdFolHCPobN4A1l2m+vtGJKkoPWzL+pZ0jJX//SJgQq6CMtuWI36v3mo9YRhcgbe
Nw++IO3KbIuEa5tJXcAmwUzIHIGkRmVHAQYxOVbiYU9iCwsyDYKe7cynUkK6GtXVIcJbcpMcfpA2
Ss63irfOXJtQaAD+ezYSBOhzT66s0sJYPu1VIG5Ix26vJNIg/a6c+md1W/UF1UhdXZ0RqKE8WC9l
POTm8kUFcvYeh3AveZ2VW0BN499YPI42H7CDh5eT/fH5UDYYxP/OFGb4HNH6sV6dwOdsxCHrDYRk
uDj0i/OnI4AVoKgKRZfT6m2uQGIwPRVF2Zo+dDyQUG2aO61f/gUkD3ZFyc7XxV4oxvwUOb9o+buh
VEIPf0XtAEztqDx9qh2uCzZErS8AhmVaBDWP4Sn3g9OjaorCWqtw0ASN0dgP406Twax26yiGboT3
yfA3KOoYiM940jWg5kqkc1xDm5PxQoHBooVViC51kK4DD0cOXA/mnIJs8rnLS4STXIflojKC2GmK
uXjaVwg3V3jBU4vcKqCPVs5b719RgzYvi8cDAyyHtZ11YmX+lvSRWuiCR7+cTPkDRNocMF0piQVp
CMZs9nEM2Iw/DDySZRnSmkCYms3pnmxHO/cMsXlYssgchZGBH+Ufb1te6+/hX1DCd/Ms/8GfI83b
LPyNxaaTQE2tfkjiAWECFm2tcxSXVoh01PwmLVW8iwNZWk0i07e1y3cGN6JWsigYaNhw4WLH1WKh
Ck2f3j4x9O90Td5Gv0nEt+auVn9Yc0PeCxX/v91CRmogPjKO1iRlyUo6ryffpvGYODHynI/RoVV5
yoB8j22i0nfYyXYjieX7dw8+L+tQqZwq/HOqCFSoQfu86tpbUjej2firdrtIkNcwxJbVG0qXl5Hg
dPmC5VZjm7/wqMat1XGGXlyrDUoVczFI+Ghzq6GL6PeQzx62k3hxTILKhgX5xcYzQ4bt7Rs/7yzk
G+4QKqWfeeSTnAq5gQPQCXPcPg4trm8y1xwrquYrN6P8mL4RQBFpbPsmCVRgQanrU4gPoD6fc1iL
8YTbJpB1gxp0G2A+LwL4qEf92s/VZKtS8Zwc4k3nxBdBS7+T37vgfMuZaHd+FSngEdfNE8gZGq6h
mfVfDRne/TZvMxK4bMybZecZKWhGz4y8G3gSGZb22+YJ7Q6BFFPd6e+6sKa3pAopXtKuBzu3cW96
26iLb/SAlVW01wA8LV8ql5/maR/T/KRGeitXmZC+q0WtfNx2WS8WdaN9+Fx3MNumnKIPklQrIlI0
HkOGMLLDZLpkhu0JtL1grHHw84DdF7OQrcyoNLel2zcgMpx1iGPwElFFzBN2hrCtE5oF2r8sO1Kg
nvQyChPvWiGIETmC5/tF7aA7ie9P+sFgWxzN8pP8AsxixCcndD+dMO2Nm15Xm0u+pQeNXzT24FZ4
J38mUOXwq/NYxxQr21rhBqfAXChmf8D8k0JTT5tqpfu78/08wS2AY6D83Lto6hAKa9gbc3Oob3ug
nhoTbE+cMhgHhJE0dgwNZEHXSgFfoXFGYOhkTcxEWcfryTxBzSBONE37dXQeYScOvD6t88dQjeOs
7njN3B5puB+IOz3V2rPXtWUjxky3X5frui4tHhr7FyFDwzPXOFP9BCWIsQ1qPtNglJddgg4b8YRC
uwUrf+NGNWyaMXmISmy17NVx+1oo1FYvQ8WX+RPB3AEEAxjUlXZ5PHq8omS8pxZEDnXcisWvONrD
TlsHkfTMfkcuT9q1HmBXXy0qrvRTqLjN+Bt0j9MoGASHv1hbPNRaiBJjKWJHwsp2a57rwFJVETPJ
QdQ5Iwcoj33F0OQCVTdU8dHkrcac3FMjpcN2GkW7pYz7CtUKXytjkoYEDlctmYCwrPJa8zJo1w17
mBJVh5hwzZqz1h8By40HsQu08NjNVqIc8PMbhcqCLm0kvrK+4ZudMjfjN1NZhYfYIlahtCGqsU1r
guog9qeliX+lvabAQKoWjmnXh6EZumCoojppB8KeFMGTmp3z1xVuz7o/+MILUdH2fR3N/Y5UVPq1
+k5mLSUC7Fu6I9lEwXOEdXZAMXa4sTeXK/sbD64Qev+lg6YDL/Yarj1HavsgAWsZc9lAqb4UHtyV
HE4q2MYh/I21JawHlmzvx3yBtBAKgj+0y+rzcL2oXFF/uh7ZlLAOlqZyZtzIlEraXyZPMW0MG0/N
fDiwIjzjKiQa1MU9ZzrOKv/+6dT3OPI4AzI1PkTZYGtGcNXxrbx0jdPXDEJGgBy/hp29/6Ol/fCp
+zZ5D7g6iglm3E0x0G0i0lYUl5qtctmMRD/3zRC2ByGohYxt/h5Bycy2Y/XMS3/nNkl9yHPcpD+B
FuomCEsEGnn9EmGMY5ZcOcx71T/f5dWkYxAItbs2KcQg2yhZBBQz0jzt7fS+K2jY3MPH4aSzlBnt
R0b1fuP+q31B1lUBksDC/FwSaPUMEMoDXXg9jIkorNYJ9MlC0Ai6ZQniHrKRdJQ8p8IcBRhpCnkJ
27Xe0b13jcAnhXILEoAjzKKEveGd5jClUgOaxt/W0XIRUM0zr95yb7p3mSSK8CYsiqqjTdodHWUN
Nlmu2x/jsnl6minbbIxCBIjvPJaGFXDyZSTNhhfXfiOYG92cWSuUgAstvh+2wCMdrnnLL50UT4j2
vDHzdZeS0eSNXSAv1xAF5SLurbAHQbKkphM0S10zbEkfRQ62cPYhqFMjfMkfcVfGQ5z4je9y2rEp
mlVMHeotHZ0gRfi2FMq7Qqs8hn+ZQS8thWKVC5A4iLWX6s9+/r08efnKTmak7mmsKqpckw39EP/y
KSEJ+v4axL48XS29kMVAhncGycb7GlfyHkuYNAU1LpHGfnxAge91igEugptz1OnqdoasM45jmRwL
fiSmtKp0srIQ55JZQQVGQXcp65lYAWP9HFBz1g6y8h9gGX0uLHcbYOUJx0MmIflvJRqBLybcfOKR
CsdhnfdrqbbinouSFrE4s/hHqbmnqLOQi09v8SCnA6Zn2OXiyV5bSPAAOLZH90yNNzCTkWyUtdgK
jTxJn/zVR19R23rWvIkr6PfxDa81WAwUK2r/ZHY4jpFu/0GukdS1BHYBGaShkH84rNcZFzTnLtl2
F5ogx9VbEjdn2DYziJ5XeCAsdRaYGg01AINus/RHTtstVkv80PLg5+ew8CNkU7lM5mG26vaFSotF
qEW4sGp1bjHwLd8q2P/PM4Vq4uNZFYEIa/fpBQV0VI7P/bp70rWm1Uphbxj4a4RqQuYDz1QmwRt6
6nZEpo1XVRHdaMZqc9+xgLET4jeuQrEng1rzOJ9i5NoXrViyaw8FO49qVtdOYZUlFFWt3jB1VOPB
ligKuyw+h8zy39FIbgXAc+uIc33ZyxXyUI/LxxV1qayxF9Z3ln4uel0NbmS9oZqgEz1crsPrr1KW
pzAqP6409BzdPsgCb1Q3bDFCOFcApktrD12MbqT4YOrBvyhvuo8sht8GZ8cpSlcTCu6MNr3lZYje
cIG7V2V8iqVzswxFbbY9KgMIDr1KVUsAKzPe58e7Yna6044aTS+4FwwyRl098UbpU8TZionsf/RN
2US2VPIDRzVaZtYy5+ot2QF6dI4A2FJFHj+jnc9jcRERe73C7iwAhoQEazl9XFkeVemAeKPMWvSq
7pinOYKHk2kXkJ+oMq4q4kpzAxZGXfb6ty9PwYID1T+Fbd1aBLW+g6tkBL/ZbtFk+B3+oM8mny/h
qyXhUAWmaRPEa21fxXhKj5alC4V84h2ZTVtKMV8BRmYAz8kgpTr8wEVneVEzBmJeHRCIxPNTROVo
5Ik3W3ElcP+3ZrCYh8hiA/KGGICgGcfbHMEkwxyuDEdLNyP9PqhqRATT+6n+K4BxSTBRXDpReRwy
AsvqUGxFMZSZh8EDeFSRtBeK5/HjvJYDcSNy0iTXCSHJ6Z4daXChI20WyY0xdy2W2TNdpDLbwWqj
yhh5HCEqXlBLHrDSk9oUjClN58RMDgAe0m8zbaGPN9unjh0p7wDy7XZKT59qeRCiqqK8nJ4/NIrr
qVS+Ic3oN0JJ7Ozo/ievMl12h6zdQcl7FpiDowytvzBjR4HPsH2UT5XZkXkDsc2qMnowBJIqg8CR
KQWSlGb9YZe9F8PwT/ybPivAlx0MMkQLYa0fgMGg0/oGKbvUsNQ3pQMWF4nGi2qt7MLmZHZMLqZ/
1KdB45G9jhGqOOviDSs8aDGUexSSgltDQAqJTxeSUM6DJf++bKCKlDHE4fgBYMeAwDemr7sVjFEW
uesEgNSBBl3/ca17eUET8wcPBwWWncp5uWnQtgmgbIy9dO9JF3iC5QHuYD/4rlTTblGlEQkXDwfl
FF9xa2aShsFEdXFY0NXtnyfbrLWz8E3GAxMsn2lRsMTdeVGTUmR8hd81ZE+SUIxkH1qzj/rIZnJV
iCVtW6cKMqQNTbqJ81+pNChqBpL6CSjwsl/k50pJnJ47v9dnQlVuE6nraAmvj3eJGHzm0SOwZRT0
NdLOjnxTZVXh2ViNqt3heB2EPKQJ7/hNua0GBnfrQdS9xTUBbl7Zact9LaZ1CwePs6ed/TqZDLzG
WOPj6VlQmj77IPe/NkZWS7ERH2sxSFWKLbVMvgoi0x4Lj3DEaHND3oQk3MKHTzyu08qdBVQR61Ui
YuO8I4O9B7zCLBynOHMcF3uRBQYzK1LX4O5x9FHtbrd+CZfbFrEz86FbqbVZ6a8zHa6CofTht+Eb
FsYgVpaNQ+3ZJrjYPpCfuIA2Bz3YaAF+r2e4byF61utDJlZcY4DkEuKbNmIpWu39U/LskZTBR8Rr
vtfYewNGUk7L9mBDJMHv4aoeIqUjNNzI7wL1V8sEU8BTHAZ3Jdh0+Swu+jxfl2TGMlbXEmOs5gSz
/+0CKJ14sXhjA7Tdpi7yvrSoiCQRQa+5loYLvASEZWe4J/nnWWKikxNmH3FiHcXbDvzxTlClRw4E
OF/KvUnOhK3vzOEhLQUjnj7NaCTCN53RHZqM4WqP2NMBuKgG9juYVmytlW/6/EOdXJYIFcxPBNib
zianUU6yMFQv5nNhcwJARvgAOxn4ayV7BCNOJl+2MhUJhq+s0rFK2vfYKjs47frI5ij0NvkHti+V
cw9uCxVUkT0xmTEeQv2cjGfSi4nO7wN7C3/Rn0Gj4EvuVrxFeaVq5jo3ecvzsiLrP+eYsTckQUZd
Kzv/62p2mBSqK/87mdVg2wVR8PmiJkfxdbsxDmJvw+z2VIrS+217484D3QGUNrz/L3HIteXCbS1d
qSja2Dx7vlqqo2/vyS6E31nLxNNr9CpATJuKrzXAl4LGFaqWAQJWHbVBOi6bEALHwPmI1mQjQKfB
2MtHPMfCvAYbq5G+h53ZIfm2iKxVChf+RBSfzy5Jgmt8AS7L5nvBEb4HLDuMN7248SUf+WT8k8k9
aScvoaxbTwU1MXdgYQoVVWyNGwJxkOTRqUvGZjBYo5RS8yL7S0Dq/kmmUR0yvurDL/N9RAnrSGq6
YuRRIZYP9LSBz5wmVKX3nplzBHcjXikSfxYjhJpEsH3rKWKIXbV/3lWyUXmOwGCdvBaWo2iRIlJm
CVJonqzeaApM/Tj3wiWYj1XnZndo5qDeb0xmtbVK45OZDGp29nGbo71yztIDNIPd/taCW7+hzwLu
MndzQog/zB+gYgStrOBhLs3o1SjVGF6iqCyWuB5hl7vy53+sA6ukCt9a+6o6Idepr6z88sJTRq3x
YvBTIQ5WQLz7grBn8VGIrXk3n/laKpZrwgAOldolsEl32JGENEoJMmO426fkvPCUB4Qk8FAfCox8
ZsEgaDPYabjE49eivROhPyklumHSPb9a8b608v/HwoJTnVov7ZiyBDfRRlW0I9d1bSlz/aRbRrEO
WU7fp2I2PiVYqAcYKQmLkjll3De5mPnl+eRskEHdoiGCUEnwYJaMDekTHUoKbuDQByDwhVS/pQux
kTvnKZtvSShbV/5dnRt20hw+nb8RRvtAcszaQbnMt1cxUZ/ItBKgsL26dnb+RClD+mhRviQ809rb
2fCCQ7duGKzE1dTEQt0cJ4OGq6b3Q8FvFOW0B7ajVpn6H2uzD9CNYWijYHyFU51+wSdx5NYRtdbs
4+gS629XFGbzDBeyZ2nF8vQsTA6r8EQoygZ4Ke+eTziJhZc868Y1PdJNiL+LiWP1s8xpJgnwx9cS
vt8riXr+0LWndTQwY3E0dA6h1imZjGJ1pOx/mgGRRwOX56fjNRkKjUfvoTITEguJvDxjxXr5VL2d
2IdjWQ4pWNtifHVZRYopjJTs2RXHEiOIp6zoq9znDReZoMarQCC8xz+lUrqL0j0aMyl/GUuP9t1m
PuKVbEs7/0Twb79cRxeIjCrl++J85eyG6bMrbDeWhCLcrciB0IzV+qTe7btBMeQKk6vymWtPTdw7
rW0fTdH2i4WU/XDlASmSK9bkAiso5MnJxFTy0KyK2EKtuELkBBHLCtI435IVHbFZj6w84epCOM90
qlPRdJJt675hMR1ZRh/2jrElapP3yEenuElJWHMOReyxknpOo8eJlEvnSnNf7yAXa6Tz/TleQHXj
oSIe99Ixm3J8R+kEHik1H1CyaHGmYPegJcAKtF8okmWL3fJ96fJC+J5MQP6ecViSYLJXObpnhqyI
OOtUGoXKF5PWKMOEwITubgBPhdPJ/+WT0GH/Bp2CrpWCIZIdt3gkoenzjtUMyieRAkBXQcLBytWw
rPj/9HyZ9my/HeZraYN1RTjvyyfud5XgC10uLy+eaCmSNVOs5nn1KSsB4TDbe6NWiYhtz1bStxVa
b20uTl3OAyaET2uvjHgvxvSfGGJ52u0mjxj7mePDPDMRo3Csn2vcsDltAZSb+CP+ShNhNp4XaKde
DOzexfdxhIyyu7m2NEUzuq6NAqr0dppzyyNljBB33ieiQsA7+NTnjG+l1M6F8ZzG6dl9zROP8DfR
NwzPHOU9ExOwWx38durFAiCvHbYbyB0L3XhVPhcZQZ37lSLnwliuIsFjSkDwyrU+P4R12VmzNIxU
Qf3c53N/94MJxFs1BA4vFhVTduC5Y8qUQAsrwmj0HHBa3S9EKgwusHABuS/vMzEhq7Kf10AMcunC
Ug/dl1V6IPVnyw+jdjn4i/6Nuq4oZXJCizQw/NFg0OH+LgUGpQHomIn7H8HuWqOrjIPjhz5/4mDy
34nPNPXliwFVXEWbCJgzHvan0DeyvAWgUJr0YZMnoOck6nfDPuxEL8R6DpNYdSdiFQfgbnHNvc8h
tM2jiVI66xLxI/9YSdAt+gO/hRJ3hTlVdgTXNkqvLo9BuaNrGfVXgkPeY7xNCpamkfwmzFpKMToI
etckN7i7XbYYRIov/+yNHrByk78qnUCrngEHgGU7Vq+d4htu/BqqWkKLpqYe3vmLpeQAmmJohaf0
H4Y+sr3m36wg50eSrUG/1av2MEjxT4T8puObZ+shYUmMSO9j5k5+02lGDSdKbeafulfEBxEay0jv
a5iwt1Fv5TeTNwPpZb8Pxm2NB5bqQMzVEPmPxwx6lD3K8VQLQNhFFT47FmEtYAm3G9keiEWJZSLW
s0t9iak3fClXgpOS+hNAMzZvY2QwmLN2Sj/hDnhwvdFsboGH69drCwrqhdjsLIoDtnTGj/aihgNc
dYhgpm9IfbDDs8THNcJui/SR4eGVuNVPkR7V97ltJ61gBKnQWtfpZwOq8qUmiWpAOMaMgNc+f7e5
ZBXmwyNhtN1hqZUSHpVUbX6Zyb3fZS9epqhhMv0VKDBLr2b5/Ep6nu6sTbC6spqhHyXHicGJw3Bh
O8ZkUjbfSkgdZoCM8uv2icm6tDg7ZZx53KGHH6sWE86tV6n9D8FyHtOAhjGlv1bm+rdDfmvIw2NA
iE8EWC5YekaJhnsGeRJv8jR96dOnus9BxkaJ8mfLhqkzZ5dWb+1zDrbnJPxVTvpd27OuandUQQ04
+qxyDSZLqjbPw6Jdt37vu1xxKQ836CFtOmcSijsLA7XN1P89yjJzDtgNtwj2aErcdsTM9L0NYkN5
OjuLb0HjWVBY41wCo+nefYcPCxDf067SyBX2krXtY7JO5HeBgBoBnvzYRxyuAqo0/ZAbcxiWIzj7
feUsdwH8XpQ1jPaY1wtY97aagF0w10rf3LJLmMzBuNfUnACoFAiPoxKt7ABah0AxKThuXmAbFhki
XAMOVm9nd8sKJe3V0a2sYXQ1asUSlpknJDg1eteHpaVCJhZcy3vLvhnfU+UzFd5Ryp/0jkMOALIf
k9yLnOnqMcyA8gkUnUYEhAoab3MrcY0E6PRHENXhCPDjmcJYy02oIcesulrX8gbwf+dIsCTHbSP2
ixUahYrDr1ELgrXh/3+xrugFrc96ZVMTJVintBsOZsfFWYiTa+dh1M4txnHk3Coozh4XZ0IYTc8s
ehxOSNX7RcbP5EntVS4k6o1NDwglOFyFCu65Lmbpw8cGdNpkJNrLEpVOGpOi95g2i4J2KG7MUicl
nTz5B2tGv6ROPZWQMfvHJVkDRmFSxtv76gY07GWwvpBVWMNYjvswPg+616Tygw8x4ekPQ+4xUr5m
70dNXTbkVoef1uRmKLwkXC1esVckml7sISDsNRv/icf+fxQdvr9Yp5TVlLoXZKS6GWxb5iRhsUqn
VdcBf6bXff8BzqN2h+TMIn6EDA+EJ6bWLhIxuirKaVi0TPE7A19TYV4XHbnbuGOdmGd1Ry9AvVn6
SAPxtBA7XmQ85gc1ItIbRMGd2/LsNGm2tB8bz7IiV7kv+PGwY9Y2/jYDRGbOirivWP4NIqrxVRn0
Wgr6A8oMNkwWpuetWzPC8sCoqvg2vyirPif0WAbJjJAnfvs8cydW6tNmWE2erARIFCf+Z69oITGJ
AIDxhui280BHzUdid3XeF1hNdGVDYIAWvqRm+ead6tLqWNvH9dtDPT5kYsCseoQ9LU0Drhx/3DlC
VSU+YAD0U+IMzMYS01IrmTsa5oGrmz5dr6YtzAZAVV8yfNszGzKQ+FW38nurrdGpZJcGo8E6+29u
WWroLXFLdy40bjAvYVYAwwCvyFKeM5IP9ThcZ3JI/Kx0tgvE6lIAenlsfgFiCONCyaalZXkn5lNf
mYHWx1icWY7XI5sDovPhgCaZrw+w/bZoQhedIis2kuak/2ic2xFQUXqvQI5wP205nvoB6NKhPOJC
UGn5mvmIpOq0ALnhujQ48M9WPztqjKAe+wSKKDUBLNTlLrrQzrVNzp1R8TrCbqyDLpXAA6VY+w8K
GLJfOXreaVI3/X71HDpQrdh7GcsMSmEX8wlr2It//eotkvFMN+jfXjDyKQpjNrsRWQjZjoG/PdnV
KKXm+fFHK8KXqF9kclQ7+TBvhKpkZ+v7ls6mNkNpRmZxnY0ejN/7Hm9e/EUo+UBASHOe1L+IRjSs
h3P2TgORAU/NMfJyAgeU13cZoo6mLCX92rpxPkoC+8MVR7vfcgw7HvgUzFKtZc4SN6Odx0kRyU7t
nep6knnHBfT0Vp4tHgEDhpldz8HbgwWqZiese84sVLwITgg0m+5g3LbXxVMjL1EwLjT3KzwcXVNE
N498XzpOe518XXBJhtXaXD+G4Ku+RxoWnkXs+a+Re7iL3bt+onoTIdRRW09LVrStBnQvDmFxawkw
NgkUejrL3bDqd6W8+1p4Y24t2pY/W7ELGz5kyCyfemmOGlFcaxP9+esT/K+MShW0f+x2DwmOlcFk
9rb68RCpgO4hlorQwXKSC+kprqLz0GqYoVYce00wvyTrPCRpP7easu9lCwAsCNVlPhy7iMns7puW
gyolpk/mv9EOGe2hf8hBe2Sg+Yt4RclTVGVjXUJoeSUmsFSq5okjZ84D7jtofsrEcm+3Of2I+DKy
QaM/MVwzHliWamKOdN8j2WaLzkNnCBspFXrNyUy5wsfD3iLTEJ7kEO893nDZFUa0dle5B/YifCYF
1mRcq06SqzVstB+sVMmq91IJuWHHfyqvAM6/wjsj03ZE5lsDdNiYwtEQgZG+VnFOummCbAsqgE/o
O2iXA8u6nkBE9Sz7XXeD3B0V48VEmX+0QtHlfmNrVxOenVrCbbJ9z6pKcRThMQ3SRDmpX+7fvM6K
njqPoGKDCZ9fYTX0cKEUBNdwF2GktJdmZ6gt/wavaUFTxpyvWSrf2R8wvkdRdzbII2gkuVmxQn3r
BbBvhbk74T15BPqMPEic9lvQJrbRaT7GoWuz0c5L5VczEkJDroW5j81bDiHR6iKaGiC3KWLGJ0Dl
n9DlArvKcPQjun7/0JyLmWGb3lXGXu3EvRlMKjh9gv0r33xwK4+XqF00JRelKcU+uSdYXLujDbLm
mT85Pp+FlVxwKg7i/3bBWBehk2cxqLVyY9XsCiS35ipEEXsr8XtBSgsrhFVnhK19o8ey4Ad6iK3I
uP4f2GclClB559VBgtBWh93Rhp6RKXdy1L5OdYIpBTZN2kx5kaUbvmj7TZaKIUBWNg0m6Vw+jIuC
tNI0Gpibj0XeT41ILTvFFIWZz3FzzV1+cmfe2AZ6RPM9Db+JHDGi5GpWcue/AhJjvUr6YVCW7fmR
oimNXK0qTF9Z0j+zAV0yvywgNtADeQu4qZIxu3tgbjoVJDwEviB65M+bxqWFCpUikm/wd9eacysh
jxu2l0ra4Jq6YLwwRfMn6oIXAkZwVJ/wAAzQDlifSSQHFNWdtkkQJ32Rzb3GcApBj6MEtChKnNgz
PKI8+5KeWna/jIG981Odn+io+1xDs2mKPOqeS72cgzzr1w68zBdGujvcQGK48Zdvl5Ytux3nr4G/
7OpTJKJjIpVnVTDcBNfUnba4e5CHQhBzEC4QUJjD8F1VIHB2jaP96pBIlAefVGGf7A98x/Upib60
RvAG9xndlo1FZnbD8SZwqZsJqoyhUxV1fUBttacinYhrl5EYI75FtG6sVDgfwfGkVTMogqkSxYQz
57c+K4o4i7yuMaeTDh6vJ8renThKWV8nrWGarwEJYSmJf1Qa+qUB6ryYJHdx7AIl4sEx1HEX1s+P
ZiwBDjZfr2A0arV+dJUM4fS+nhAMypZA7KsEwXEmjQt83m1H4Fo8ke8mPU6/cB5YuP1I6t9BoS/Q
CpBQeODpkeQFEKdS5sSjuHfpht4XR1fFkEUEfiLemnoRl/AbGozme6Tts7bDBta+Z0SBQTeQXRK5
IApm1SHaxdwJ68laW2C9mvrHjjCYjZWNjAnqDUViZ/C+gHuIE4COe3XvLOx5yWaUM2WbzdS819mE
M1PZ188ywdOL3KCU0vp51XTlEYWs73q3B11+rlRneEhiV1erYMeB79Pyy7QV3tUeEc1ZvZUEq89e
FFJz3SMZdDm/kE9wiRbcwfLiQEoTCFLU/w2AjGKx8i3o7k813GvZb4mC23vCvpb6y5v0bnqTldJ0
Vi21io1HvTxnM6UgXSklCSW3rg+F+ABNi13ifL6Qz2E3/zWy8bBwdxCqdWrH5YuLen1LOx+NGT23
HAneo1bVodsgCcQ4nLhaIjaeCrl7X1am5vIYdW3WHs52Fe3YSPKqi9ndrbKgoBEiQL25oleE2/yb
o1DGnxwy3dioxTZrvQI4cDC7TNLd4LobOJjHMupbZodb+YVcokrn4bEjnvU6iskTwZG8IhC9+6O2
USrKWt+YqhHehV50l20zfNhD4haLU8vOyTjj7faOQfO8oqWn4OanwCcY3YynYf3fAwh5pNx3eOfo
IRcywNxiPj4J+7zaG0tnlAEvrMaQJdUZGdmLPoyeJ9iJsvOGzuSoh+AUssYG4VHEoUEjIu509iKh
FDwcscatD+lR0BEXQznSyDFBJ5VZih2d5Wvn0lXKcJ8zj5o/Q75LuqL0ixaQUwmD2kIaaycAjtnm
wgcOw/92zdmlMfjMX9Fi6x2fW7iV0VECoviReo6f00/A1g4ST2gwNiJ6e5LOE4+yReeqnSRXc4PI
Z0NoPrn/cZb7RSTqSpB5jUBp+MTzJl9eeMAZX3fxZRNZ5nb5RYLFeybuoHwaUVeXh5faGAT3CfcA
AF4jwcu7Wr09AtTwgYxrG6AxYHasaqtOfmV0/Z+GBzsnDDqOmbMcwd3VVA44zriA4ILvK530QUCJ
s6pjTXaG2e5vM5f9GLdxc/p9zU5o1sC1OuKJ+bdRBRrZNz4nfjJpLT/KivFeUMuxmnP10CwRSDAb
8OpVLzfDNF/rQOXgy9l2IJ6Gklxi0GlraqRlo+iNkwJjfKqwGpoDYyFlo6HufmNXGIHNSkRl8cK5
CPSFE3KizlSJDa3OGPoAhcvNZJlTIV/z8f4oKH062EfMmORQHCCbPBAa79LBSXonJjuX+BlCVdwG
IdjuOfGh2JXYTD6dSQRPvTaT/cVK03Ss01GXZw1kMk95bJSwyKalw9LXIPDqFRFgpLOHqCaezNQG
pXYoNYYpFQhw3X4klXqRvsDin88SRe4IFjngwzoszyb9fCtbHQQrA0PoGVFZSMaZNqAi7Q6K4BEs
82te6YWazSFRkHel7C/ka4oV7oS5hBzCiNTuTMLJ0u/vFir9KpQ7T3/J6fh95Io6VWehjEedRDXy
dwqnDhizZnxHnL7DozU7WNM6uEpDETCap8sm3zp6z0576Sz8NdYTLgcJednepBm0mlBsWkBD58+8
Pfgd1T2Ab+Zb0bMDsrxaJl4JpVp8MB/1f3XaPwZc96V6N0MSzI9/+hmeIETD9chHDFZfnWFYk2zB
SxmyomHvX5SHhA5JaYIGL49KGlOA7RZWgrEEcUPgak7QTrk4mSqgGTBqhlwMz/dz+F61Udc2Jcls
O5fgczQeZ07T8//42OzxZES/9cuWrHtxlH/7x7zWtFRgjaMp1/JlATvyoQKGbBL9L21AmbPPxHY/
OCpfkSQe3ZOwBDbPB292D3/sqensB2bThWV3AxQEUtk/2ZRChM4fh9OFDN2VvWK9Q3xnsJy0Pv98
jkJwLjcZ4f18w8KfJ6Sqdrd/yo5N/Tv3SJbQYigXXcRzWDAu7uEiZ5ZsOdf5NAwR0xrNF2LJ+IDM
J4oUzj1+70X/mJxaZ1VkgFcF5iRDQEG+KSTzqk5UkXoiQchptJS6tMJLRle08upnLZNowr0Fzkf2
sQSl24uefNaztjw0jo7IhO7WxlrMC0FMRdQ9UHBdXD+wKXY8PWs6Ep8ux2tUj92yi/oTDdAWpcyV
a82eXkFBdPsbZeAZeQdWFLo+deGNR908fNnCF+KnepKfTTK9zrovQpuGz1HwVGX58qxC7gbZ3n7N
q++5ib4d4K8WcmUFZa0yYnzeViZRHTQ1WlQfVokUmmK43VtcIaTLKbZO6YcVXiOHODE5HnJpkN3A
XBhUmWhuaCO0U/VB6CuXfnfr1Fbipj+fffDHLcq+UoSFXJ/+6V9JQ+WlBbAqo6p7fknIrv6Dbn8h
dF8FOwLjxMD9cZcQZUj8Z8QiKNgAxLEQ6iHE7tGef+ZMq/+XwQRe6MbRQh/XejDMwDkV1VPUgj3k
9z83sxIIU60h+5dlk8AfRR2ovUnSTFZBRZzPMbeGOV+t8Bbji7gRlQ53fZbOkIGaCH1mVsoptK3x
exMvJv+Sp61ldnTgNIITwOfg3FKQYA6k35fIMZrgWoOE7Tw/WlEFmF6opdsKCgf0LXcl4kViRevM
TMDury+3CAu4gTgrRqHuzEow9oT2Aj+DlNQN+OdGkmXFGLjU3waWc74fdnzFwE6m5qVj1mmDvpmZ
+D5ePyy8ySwkbDu8O39HKyajHFN8MEO+CjI4beuhh4Y8dAUc1YPRlNQYPVVbSce2mRVX+jpxE6xW
r8+ZpomuZbg0LLif4oUTfcGg0bmtc+Z4KNoMgUOh7gNcfzWM7v4VoDk9zW472o/umXSKRlJ0eu4y
bOvcpxxjXPaxM+qj3xQitE3SBMkEXl5aiDkT/KSABxgTnC3jpf+/WCykImo/zW9wxMstX/OPGxN4
R1o7FAz7LWZFb/eS3HOtfc98Xn2yDnBjw427m602kuKIQRwPJfYOtobwYn/BppJYQl+nezoBbV9f
iWp6G2TIOOu0wNP9x/MtGV5HsYV0VHLwkVDeJ6GMXlWMXShMQct9iUjBdJ/E/ROHvBifJI5iEgtd
LrvU/HLYtAF+Rw35rcBei2jzS0xLYUcEP+5/WJ4HEd7tlWogDLbltWn9ui7DiAHjjPt92Ndlp43t
cGb4F2PNIebv/E3p4Cs3odVstlcu9MvC09b2YrXj6PgaTaiwJpZrfRwThn2vDkq9iyG+0TtsOTnE
Lvj/j1DhtM8e2VfFWOsVRwXpUjFSwe22yKrpxJnfRGJmgGME+o118zRF/XXG3PWf44rqinsnz6Ht
LzU0V6ABv6Eqoh2TbCyl8RaI8M+7qttxXFYu+yH1adF4HiiSLcxlaTHZbj2fRktwRmvkFEYhEOzS
K0NiwrtrN+M1A/9mRtewsj7A2yJoqtIGYPg/SeaJI8JIfbEGeuRM6HtsHS6uVU8u7iGQxLF+xHwd
7rPMwLtUam+6htkaPGbM4obqnUdtUkYfZwigBg57P5DU1+IhDGNN9CofBVbpJZwt7DGGprlxTgoR
U9o06jsrxmYUMVVXe4cZHczOk3Rt9vHmoxPZ48Nx6BlzATodAtD27QVjJ4nxEelGlF/Q7Bm2pLTY
zCXCDOQhPL0Z/JD/hRGze7QCPHMrMtqDfZYIuqo8SE5dacrxebyEGAKKwz1RqB0uRBUVANtGhKIp
UNiE5xJnB1YaE9F02/V+EF4NTwbQDIR0jEbgJ4AxSE/kKgios5P3Lw+jSxmh0/uDemTR9xxKCN9/
LU6Bcs0tPZ4SE4u0VqL+74Ymxup/wFjrtFjk3iYp0vRHv7mkP5ABwEudMyhc8LNxBDNW2Ovl+LAu
cTQSQwG7FjzLkGWhNev23zZDK/zpj85s+i9UftFc0ewD6NlCPLHw3XdTAQSGyTX1Ou8rxOf1xPjD
PGPEOHfZNfVV9Ij7cmPaPpZ5egbkebO21+nTWD7VcQyR6zb2w6aMAxDM9j0RQrA3hxpGhQlF6ZOH
8TelS0MB+sEhiEoEbYsPqQZZ6l+QXsn/1BziGAWS9ENO2EGwUjS//blC3Ap/j6i+8Tgc6EbAxdD4
62O/IL2S7ZqTVuoc0ictxhFh1OQdkTz4i6aY0W68CzJ+PviDlkoz2pmFuWk+OK6egYbsGIMDRiq/
CKxGdTnab7Eo+oPXj/qWR/STgAzEiQNUpnwPXRdVjwyD6ve+k09c12sfrH0cXs84x04pMBIACBkX
bfM8cuYt0VKrMdJxJz5Bcf8ZJGfiLPsXS9nngqt9N+RfPaZejh8/2uZbUmc78/fIWZvOg3TDQ594
fKDfzoL4SMDUfW85GRl6tFLTj4YOdjnMEbrApAqgx2rtET4RP6ZzKSqiCJoAdFiYy25Ut/RgxbOU
EOjbrBkC66OaKIvVFCl4bPaIOxLOb40iljQUGvMDNYIpj5Q6GskAFBz7oSV1s6rAWvCAKoKws8gm
ubFxzJKlEp2r33oT4zlYpZ9WeU/aXygZ0jReq+PnhWsG3TkD6Ee4voA/vYmzgtqYpnW7jTrcXEBF
nDW+UXhACPREaiAybUo3wdKHyGf59soxKzvQCacz8plqcNX+IuXZ8xjuiovRMbw7WayrEbak99Fy
74YfUWapdsM3nTpMQazI4ELX8Hx9iQHcaa79zGfxxdX+BE6gzEPvjjQfHYjiXi9aR6LZJWEYVNhy
ZhG84i9Pf1pg6wgzgeEd7XDaNC6OqaYI9Z9YNqdWQ3Z7cPl9ubwM1YEZjhVNAQonGwSyfjFd8vpN
qzZ50jMb968yCqOM01JwBIAJNgQaSSO0izlxcQWl++IqeX6ZJnp19aGKhpjNHTtdOMuFI1tNRZuR
NPzP+Xq25obf2t/ZLW0KWkUbhIJ98rSxSo1x+G9p80nTTIuWcgv7z5aiEHUHP64JV7W99EaZ06An
PNF1zYjO3Rhw9ydeQAOb6uNAg6N+GoPDgq6hSMgCDjaUr48XHg481Fou6U6Gw+e56gnXRTfRCccd
fhnKJiTnZ3cUt8g5vnzbrEeMXtSq+CoKqSd1ukPr1begXbawYWmhmKLN//0+88CM6vO6GNpDnz9N
BvioeVAy1awGcv7oUC30YVRTOGSHg3eSxzPQlPnNeRCZDSPZ9luZVnt6qfsfS/h31VgoLnIM7H6X
kQqUU3h/WounRqVpIJ5Bl6hmroqSQRpD2Q8ckm5EZfzbQJfcuGGcyR+AbRk+zhIanjXSmFtxFQ0U
WtTcRQA0j7WhpoBSx7eIL4upolW0hqpas4jLtyUFzZ2L4dbs4aORIvHa9i/ynL51gGMQhhvlZ27Q
ThlD8JkKxK6BlIfriz2xeJ2zks6MfrSJNzG3euovVUk061vkSBFjCC4Fp2bawyr8XHnj7etkjVUe
+1UQMvKN1cVAmsEpwepfBWpIQ+bwASB/H9VFlh75TKPM1AkekyheUkfR7FlWk377eJMkApDGpUZh
hT6mYZCP8Rq/6uj90SJ6F1eFWmE74KCFFp7Zh9yyvQWHaw5V/7vXgkfkg7tjgqDKS2/WjsYSA2an
jfJeTweoCoL8I0e0vq+Es+xTyGoZLS2qvfP+Ju/K5ReQtgutZ9hLocqD9MByr/+xNFSnelc//34H
sYKjKNnMRbJAdi7CWgu+fQZvH9msa1Du6LzsFOOrS97uZo+Lrthiv0dR3UWHR+we5aEdSn4YmiA+
Pka6XBEOsoPbu8HAAKbW1bivNFGt6RWJ7nSHFka3hinAuhK07xFPghojXuThtZx1tpLPpYG9BxLT
1U3APJMA7Pmtx5Y2DYJPmrgdFiMHJbJ8FLP0tnhrDe4SivDOGJ5qlEAhPpxAn5SK7zbaukzy/8aO
CijJ9XgUyFzoSpW1QkQR3tAZjtwWtr7PN7QUX8wrvTsK6NK9pkyy4XdG7Vr+9xcIedo2WBmNPy9W
M5w6S8jp1/W4VewyLNmB7vQmQB49EjvZx9ic3uzVdf1VF00UL4RFWh2Mym1wsA0DpmpEDpflOhK5
zIQNnfge1y2j6ZLzLaWOlO+pLnb9PUDGdERMCsZCR91231G3/uBxWVexD+A3/A/i6A2qWIXqC9Rr
jzNQlSTyWa8dAvUVllHbDAEAJbPH5sK0ulSLE7HdUdY64vqcm0c8Ybo88RNjxm/SJMhgt2wrHMUi
q7uer+ZlQ/2rjgqnE6ohYLE8g+lRuZXgTr6XcIEZuHezRBFWn6cDR+gz3nJNRu4OmPHEf0KvOeZL
PPlUrZ8BwFJiSFKuE6zQuOSBFR2DiYI3u+OTkZM+Mpuh7Gi0GGZ4l4Gtfy4tPEXlyA+DoqL7ANsF
Rn70eGN8MUx7oDHCBdN+8sfzr0zANNjGVAMQrILSleYKkL4Nc26MewkXz0qVU3Np/MQl4tSktR/Y
Tpi40B9yOzHBOeEybNKOgH7hlC1yDkXiIlCJ4B9yf+8fnYwkLIUkr+2UbaPu5IHG1/DyvWn+rqKS
3NkXz/hZUiieiQ/GcmHduUc8DhXijP/QuV19C1UcD8LMi2qGtsQI+52h181M+8+ijGkkC22Xothn
LNzkHbQheusDzNWb0WgeKzRfG/hlDWoNBlHmTIHKzlGJ9jgh4Xgimu7uVEKxRep0pMJDudH3KI/8
21e//Lg7IticCgZBxkWBJqO+uqJdBIT2eLbx9BTGzcf6IIzwpQnLv0q4Dhb50OGQt9q/D8N635iO
amPWAhL3BUhDhh2Xq0Vg7oGpN9jsMR6xQddnN2EFOp1mckPunqrUROTkuynPeFu4J2izDWfbIgz8
GqQyILbHPPcggwOX5pFHVsXpIYGdaVakgZZ3idQFqJJVI6YbWSnea1661bER+at/I/FlNfcaPPpg
iBPTJf0l01gmDdE28oXtLJsPJeURQ7yEXs2+KAZlpkPn2DjDadYgSW0z0lvtm8wGQqO9fnG0vA1P
ZO5igcHBThbxJo62nd4zfIehA8t7nrZwFWlUNwxc1zW1pGGxNXRC6viPQKHUmF6UeHtxqmQe39dx
UGJKBvviDA27jdMLYMh+WlDxlCucLGThbR6w4Nd1igQOORq2MnNHCTbqhL5rt17truRX+jNIgNQL
IZHJF90aifdtBGAXj2ndPReMuqX252F9tLy4Yglb+Lygkg7MtAo2tDNiGLOQm1gWH0WCuObDfCdl
As5Wx3lG3HIM/DL3qQXsA8L4HoEQfKmadz+tHzUqYE7ai3nh8H1lLhh+/5Ds0cqPvCTH9rpGJb/5
p+e9mii563oJahSa7hq3VaTeBnb4KdrbsURGXxM1ymBbQAH7xID5QagaK6DsPj5ZBGLtN93g73n/
1PQBpZ2+5DTbG5ImoYie5V1vzo24IPHdOuiyoEVlU9q7bJvXT/oGgoikbT48BpbFv3UcKrBsRVZ7
henHv0mhT3ZyXQ9cWE/nRwFwYH224wMCrGf1mCJmSRLLJEdMXLJBRJQJo3oVfHrv5trzAByROKJj
C5ynWewG8SLnJa3AoJUbRoLqmACsveyCanFRGkoZbfvCoQ4G9IcgdfpbJAMeFKb1sL/sPK2xKWQE
bwOsCHiXZ01I6hv2Fy+8c8N8QJhLGUuAjdvxU5nzEUAkVIaj6GQIXZFoCGc757f1/gbSQhOByhBR
17c5rlQVKbBRoHvgit+mwsSYJT5ZboJoToYo+XQplPVm7WZVCpSzgwxO8KZ9y+3S8Aaknbg/ef1F
0+Xlg/FAm4eJyIRjbMygLtkLd3jjFPvTRYsMejfvUBVAJu9pJjy4uOl69q+YtJSwh2fdgY0DtQwm
CZGgY1KQfJ5qB5fe+ABzwjEhNp+GRYzCxvyG8Nh8v9UsWUR28kKnxpHDnxgQlSW1mOOxnSjlK5gq
TJ4YNFcaHT+Qhvw5TSQ3c9tNKIamOMiYTHIB5msj96Ci1OmnOXLGMkbfAcmRSISvHdDM07aLMH66
QEUXkzmFrLxNGCtcSvNumoBgMW2y5Ug5dEs3PdpOr1cN2bSfZnImInPSa77DfeVQLSr6/wdjKOMk
0CzLsKEAWiH0OyMihF3GenFwnivgz8ZD2SYEWEwmNExAHWTYTOfzIgwJ9nR3EWa2sWgq4F7NMfQd
ErjesLEt3gar76gdbXb8+ucR0WjhggLQinMZCAw1coDwbu6jkrn2ZCqXQsExfHAmlj2t1qc3cV23
le2JrAzg8w2orB1kwFRgbQ+uQjQ9/Dl9eIhYM+dShEFm7/qa+oklwK1oAr4Lhy5DyUGrnlqNX1Ce
E9xLSdQ4HwTd9fHigAact8wGA6m0bdgQpApq2TO7MU29WOKQ1qjSI36ruqa8nLIOfqS9c0SGiRYz
ofT6vN8BdpcgYphs/NU7m5r7Qd8bcLcB/gETta6xONVgIccHVxtvZ2YQCaxboYFTDOTbncudsIOO
DjWZ+aqP7dACVZ/kD4b3v4MakjuMjzVK/O5/zghRVUjVjDZ+2G48B3MMY45o4PMjIt5oKOkvIs6l
P+Q4jrt2tl94yzk6VA41/cHErDcQGlSN+0Yz0v91yjI+DME0ri3+rpgs0m4pbVK7K0s6UHslYgev
2n2QwzOtBmnaWvYalaz1Zv1Vw/9rYnr5whLpyBk1nSPm/tMiZbU1zfuQWr+EsVSXIcmh+cS5CGFV
LTXuIMIX7QZKBA5AdJXQ4nq8YeuQMhOCslPJ1kpc0slBbtfOzB4ofIAbAWG9nLN2vtxR6TEORZyQ
98KwHi+VUGyePnmOtkkZiUmke31et+oNPFAyzQ8eXMysnOHzMC/RTlhTygOzGmIiCSyH2h8TpXF8
qZbGr9gnAs+35Js52XtTxaILlD1xZ7dq/7jp0z7d6EhCARDKt01fR9tGK0WPQeKGtUE81pKFSlek
T+DeSDqUYlTJq96X7u5l83QbsrmTkSH+JUQvjzmeyFbPd4lIdjp0tJaaOU2WLlhiJuMjiQSoThgg
jscalmOP+hNGgwmG/KFaFyynqmwCIUoonH/oENR78B2V8LuZyEwuhS4lRIEHft+cZ9amjQdT1ZJZ
NI3PqcY7elNfHAo6exMhK1CMv43x6YBn6HR1GfvHuqej6iFmsMIPKrNOoOumuRAE7K1gmGSLhB1P
YdJDWSXCTNvofa0pqnmsQzdnlvbK1SOcX46fF44a60sZD+OhaXPDBOdIe1czKOU8oLLyIEpHliIp
62Q3TeBFqBOOv+XOsPQTGGhE24VYeLmVx/eslAncRUBJjue3/7f0sGOWMZRURI3lhdyW+o2YwTbo
pPimQG7kzzXN4AG0uSPqHELm5wQ5ne8obduv0QvoPmE9sumFDuB1BkJyW/5nxr/n79KRIuPxlNwl
ADCBiYDp+4ZRf7qClCClVNEvmS7NL0GrUlETtbpCpNrDLj4eTGiNVkIqB0+kADzlqChZ9hj0m/2+
taeefxn28R6XEsfeDF1ngfbrpgnAYYi2DweUTBw+aUAAFzQkGR4KnzDfem0y4YWQ88FMRrGmoh+8
r4+MWjq1It/ANh42IKUO69G/NTBmKCyUstnlDKUMzMJ4xE3HmFe7AAZto/JBGtUT/HPS96YlM8z0
Poq8/q6V9yEeiyt82Xs+lxki1hvJfz8iQkrV5oggj2jRZSpfKGvRpj5ub8GdbcOVrjieO+4G62nn
NvBNYIlGdXFvzVeahltnthCe622KAQRO5OVSP1E0QbFgO2toIitkJzEC6L8a3U6qs2mGbCHAZNxC
imRcB3c9A1VUS6ds7qqTTjxyfXY2qiOB3BxIhEGphyMMoHjH+1seqVK+rkJ6/NHnv8Wy3zLfGM+A
2lj20JPswBKvg5aARukoszWY9bUHJN3WWx+XPbqdsOjAGgPmGno8tQTW7kDPoXhCjrYDzcE+ZLh+
sAO0G/+bmrwx+BbAuaMZUKgtRZxnPzW+aIAeZJyFSbuc4Sz++cRP94uNpfngILRtT2iBodiRs1UP
l7Wzea/NWUAdcQr+45Tt7i3DJfmbqZ/zUCuv2P+iHBEEz0X4N2tQSYxhz1NANlsftL93bjdYJBCc
T8WOxg01AA9uX2Tyzkqt+vSCvIe7tuPnRMd47LTyMgVImoP/kspx0rRAa6oNgKd1eA9GQjiwKdGN
HuH9GNUm6tjkRjXzbJD6CFzaHHtmMx+eAxr7YcH/PfMWWTKtvEggqHGaY9YaPc2ZrNzxRZM2AYLr
4SUgnQA393+7fgntUWvs4NBjhx/BruKcPQG6004aYRDyPhZbCEkUJ+Mfo65riZBc43mBWmKFp11I
5bii4Rwzdkr8MMrljfsinCUyrZzODzqNQQE+hWGqURE7jCDL19Jff6AB83as8W+3leycbcF4jHZY
JRpZ4K+BNy/0tAyYdgDlNNKD+IgmDjaj8OgXWwj5Av1FzWKXt/kbkH2Q57ELbPtBQ6zfvCbnv4E6
Ge+fp0P3AQDTfW0edTQ2I1UrqrC/YxhnnBrkEcVJh+bhX82sm9+zZYkMDyO4htncZJBdwwbxq5lr
yx07Y0MsXnilEElQUX7BlsehVgK9xvReu56yQGzPKGqmDuhQJmWP3gQqCkGT1GMEAc3whve2/P8k
V5TJ5LJggi3rIZDgGRCU6MPgRntkL4wHEiMe0bA0DIJsQyXgQUsd21vL1KgUDjUvs6hWZHSIqowr
zLJBZwnd0yfRvGyBNcjTxYnBLctem6NN0ikJlBq1m94K12uYJRMV9s5dzMhC7PhKBkBMpC7fWD8t
Vi/phpSLyyZwnny/Q7dzFLZ9ej1IYxCX5uDHUJStnZzOCLPRg2r23VBsfylY3WsCjtc8eph5e8M7
DgsovuAY9a2j/NlmVnhdh9QDxndzWpctC5POMcTHcF+IgzVFJfakPi05rHKuS9R9CbHs8Y5zgDL2
T5nAJaCIN67dBBaDLZmaTymwh0Tm2dOog8fwGrcF8C3MO7bcO4DCklRbuVceaJkaknlmRJjjDRbW
N3s0u3uebW7MFlQLMnldcftlONiQ9u5KQeV3hV1I1qC5qy6Vn3D8Jxecczmkx4gR90/vgNRFej/I
N6t51Hj9dfPqNhNVgRjdvGC2/9C7is38zKbCB+VGtDjQkshSXbn+vFeOsKZ2JDv/qbpPlpMxSsft
q6DSWoDO9nITriKhUzji3AOBFCqtOCTg7RaJ5/e/L5XD3rTGBqo9gUphFoZjSW2HTxvIkynT9yKs
qqOXw46XLd+MpyIk8a5lkR6uD6v0cK7Nt4wpbJyel1qx0wq+cdvVgdQ31T5j0ejUqZjRp4gdGEpm
+MZZq8iY2b92nE3mPP366OG1loV3B+jzgwWcGEzxzEHjTyV1Slk/4dH9VeA0n/CYMws6f+6YwX9A
twQvoX0+4iy42pboGrBJ8xCe3a4BvOcXnqxCOyfxHwOyoxZDGw3492Ql27wBgeIw3vvCDzy74vdu
xzgw0wngKjAg8i0qjNCGqJwsjSq6oz5CjCcrylTIOb5C1v1q39a/EAWPB9ohRP5aIncrLAs7JGkc
lxFDlcXWTglRUsgrOpp5IEpx+SEYUzxXQWBCaCKCTEJ78Ql6hO2OsU8+GB3pRG0L9DPPsDNAUvFW
sYpLpN7jc//zpEFqs1NKZQRrNRl74mK3I8aZDmP544jMBdx17E6VYV+JPbqU3ichTvoR6NOh7mG/
elEordsbPc7wFdcSX6f1ZMIHgpVB5JXEtX7NTQczNa2O71rJFCTOWZQuhChD3r53C4xt0NBZPAqH
anC8XUKFIz0Q9jABPNEY4IjrIuyQPy6cRWYnu6dH1sQ/MvcJqC/DN6jVpWa49nUAs7Vq1IqfDWrG
C6TshUomnElyXQXjEZLjp0qQtvefzJ6cYCsxkkIbcp+zxoIkpBO3QLsm5Y97TonFiVBCugHkrH8Q
4TCTjkLMyak/CtXFZJHnRiUf+B+p5md4cGJOWnHCQs7et+qroAjr7eFBS2gjCkY2igeMOedz8C55
R9p2OUbAODgnhTzbhH/ZjAcHH8Y8wpzVNsTlgFV/quMjAnbrtcXUYxbOTmMROH3n2NgN20ya4o5+
zIipF35WoxvJ+2SPlcG2korOC0Q3aq4rpEcn+ar/zQ0yU5Rjp4PKUnBaPw3gv7pdfQssHvWb6DM7
mqFWcU1tGJFX/vJd/AT3UWtUXQMOzskUTMe9BsZa7L0WM18fcD9f7iTBQa8n0vqGU8doBaF+E3gi
gduV/LtFPZY7kivBePvgJnyDX+cQ1v4xuYcKv3jnB6rQFAc7mit3VsF/bsnlJm0Ic0bta7h9lSsU
qjS6UngS4sUa1OP31De+hqAWUTIDGbTCQEOVmGayGLSNRs5WXVHkIKOt/IcR2iaatE0Hz4rKndZO
yPSOxYTqN4rMqrsRPZ1Eyj1B7+TZVjvoia79yzeOfSY3Qe6eUpz0drnYrJvhaXJuhXYGXfQhWThq
D4tHinwpjIgzXMGI5RWPlLTqUIFmISzLVCY5TPpPfUswcwHqw+x+QOB/8prS5wmi8fNJeuR9r7UF
EMEnd+pcAa6WKkWrOFf2GQl+LMgjLF3bJC2WZWo4NuOFZLhLz3d+MAfItBimssjha4KgU1tbGTSc
hgDFKbjmckRiX7Dl/3YcjJpH4E5IjF+zRbZ/EBCUWXHY0k/0oNzhVzaghiCDt59XaGPdyBHm4Ny+
RZGc86p5jYesZCXEyGQULHDY2Fmnk7zwf0zQOykioykDybN56K2NutHuJ3MAwTTzUcwl8DL6G6JO
y8T3G2Q/vNaIPMrg2n+spNEsUjRMy+7rZBlNfZ3S14JrSMc98PUUc7F1gwCS0pu/eXRHBxUB7rrC
lt46lspHE2F+5Vxw35roEkGFlNdeD5WhJgn2ttaNYVJaFvTwv3ZW89SP2h1UqHRbL9dPoSyP3dKi
ZExc56hnPFPkw87OOcli6f9WoZhTHS5eEKs+s6zcgI4BDKmzpiYnazE5dVNS82pQpEwbKdpSNkyN
gwbAfwUTnQJPvJUfo5RHu/DnxZRoIDlObFadVkYY+671L0vUoVi5Zgt4h45RJaB0/ZSCQKNLDbOt
CCXpo3et4Tw9C2/uNpOp/UAW5nbq19vzTWGMiCn2qg68TjSQDCdZLBWSeeLSQBApEeMvZKkocgOx
tCmymqb8crcdnG+0AXtJcVcl1PRXHb8Q8EwsNrcbdN2HIENVwfFfjH590t+4+8UsVs7IoZhEsYR+
9Pg1XaCHj2gMkHjLll8vBDycoaI91PvMOPxM41xqrq1kDrqmugIkndE9RnnW7ABSI/P3tfWFkI6j
Jv2gS2eqgloRN8douNysvJRP9aY8Yn+1GuS1BVqXhyIJE2B8Ox0F0aI3/uPxpeDwhdksS+AfHehR
ML/olEm1VYuC+UsVICFNA81gOgs/p4+ygXcoui1Oqtjeefaw9zYD6YWx4rl5GfVzfyMM6ZNa/vMO
AF4mOVZodLEFt8bwxIS5LZwFLSUufX28zSuAzIlvWEbION1n9v7c2aXjHbRUkPP7AGv2yfmUETP/
pEKTrPLPAvvni0XOk/PuILc2Y1tVufmtS+cjI7s+rK2yDRVPIrckrwEv/ACx2jC8zMA2kP0rvQF6
LxjmBiyChd436lUpjcT8Gei+xguxg/HD66n2bxgCzqPxGGKeup8UW6W7zvpzRO2ZFcw8xd88bBFv
Ivys2Kd/xwL0hiOXcg0i0GYDeRKZelH6JPmnbjvn7TdtlEFuOLl/X5tZyo32q9vyETejNJzunQDB
LdwxlubuRmbzN6d9HdVsfkDvkH3T3bavZzxqU7UZ/E7YMK3EZrp8fm4YZrT4n1sVTbCfD/o8nmKB
IDIIpe6lkP4RZsBJshAJYogIR8ku9POSkmc741SxbXih34hf2DiMyxx9/Tp4Vj5zg1Gc8Nqj11ip
Gj/pQQbPfys9MFq6odQB0Bqv4XJrjcYpgo9E6216I6kTztZbI45wX3L3HGzBa/y6xI5rPvMKRmX0
V3g7C/VBHwcCbINbeZNXjKzTeo3yF+U/Z+Fdk6NSaaBnL0v8Jt0MqHv34L0qAj4RbtEXHXBvMmH+
QmoWtuzorMAOaTTYFoc7y3H8ktpM6+Fk4wnP6Grg/05Xmf8OJfxZcrZkavKioPMOUkydPz5gBTP6
7cklNRQpJeG8ULg578U33+5xyNmep+b8IgpYXAG0FIzPKjO0hvxkH/FVjcIBno1PwQPYUfq396eJ
dLkdIWADgY1vgjCWTb99uh7R5P39lch4L465WBST+r1XA5MX6AGb2Cfw1GjyKHxNWg5nhu97gHNI
+fs3v0TfVcQKomdu+GNF45y9hTbq+tHBfjaiSpNcurVzKWaTcoVNINvhgvDDqFg58K9ZZyx16FJ4
LogfWTw5XO57Uu8r0445gLt8tRVBCG97uEj+SdCb1bGLhaxfuRHeGlhDxFNZIFnXOq3UvdUC8c0O
/MZtIGIl41t0n6LNlCJQbTzjIpmPsYuxiU7BoCyZOGpEqQ2g6CUri860mmmis7R2w8s0WpL4T9cu
yndmc3jYiaSLIcFZiNcf6dPIYMTHFSUzHokpGrHx8iFcUK8M9yEmm9448RWAxSu7UXJuhPC756wd
Z1U3bJbYFcqxNh9ee7BnU9oDceUMKMQbnfXl5as24EDwvs0dt33deYKaUXPqGZbKpsQ7gqvh4LUS
v/DoFXgyIZA2JkaJ9S/8Df07HK+lZeTaozLKAjWbNn/zrqxKUGSzdqQzW7boKhqFE5/Z334ZriIY
6EbJgkdZ6b+f+zo5/4SHBYL9CS1qNgOy9ef8RGc+NQ32XmdtIX63lBKv+BHC+z1beAAU1dq1t4yP
Zg/+jmmNVeHT062Y7VW8I7+QIWEM/CCT26l2AevYuN6vHErw70CLrFkGxELgoMEW5EF+mRBQSIls
AYhA9qHEwxLJZk0p176K+UWBjpy0kAUugF2TfiZSXCe1NvHugyHR3PNrk1cbbJJfqNgDqKhIWNAU
H92ZNFxFMvvOBmy/uwvBA9x+Bm0y7UhigW2+trdrLfrOPH8I06Ts+hy5LwWS70TeC3/6x+yUTmtK
uEIFNgxRRE1XMIzcjClokQ9OvwlLtPbayMmeSDD3VgaWjHfOv2uozT52Afxa5y86eYvnoLp+342W
Zw4rGcHlIkjh+IDKQ3eq3G5tQh+0fDWyosM/vGjVisyizbkQJ/FXd6jsWVIud+jYMhhR7ezizoyK
2aZDU5I2HNcIdtfJQy3BdNij6JjMNdIluYsmjRJWhamMscJv7DbhRpCvXKrVJUVBFhtbC2aehxPi
gM6QttiYSEpp6gEXT8y53ZV2VVoafG/3at5fK6/FuT2aRnw7rXxlJwYr6OK7vf0Ocz+aiB3FwuqY
9hzFsbljuSDSwqJYNdxhOC2Vy/39EbPOvb3cqU4XfjyAXY/b09Tj605lm/6p2+DG7fZgMDTvcA/L
hsgyX2e1+B9FM3D8SMuKeFad44m5lh9ssSWDHNLQOR8BRdOn6JQRzJ7gLmLYGWM8r4TFwbEuqYMg
m3TMw41hSwsKltzv/JL/ADUfYOF6B5tZCq6dAnpn1K7v5o2EFYpWHa1psfD2PEpIISq3Tlo6SP7U
ZjD4gQP+KICnWIV7cISk1K04TRnB5XgFhJH9mOCuENVmjl9ovUzqNkFTL3mN4urUG1uiYHrUgoAQ
e05rzVWzpd37eIYXZG/n+HAGEPI22Z2RwlvpWwXAa2N+Y+AHJBmIPTmJU3XP9ivOaQQCNefxOX3G
u+tVH1MOcNI4Q2gilflJUjeIPX1my8PBhdE2WWs7g/v55wDXzao0BjAt4wSksAj17mIGPr62lzEp
ZDE2b+WX2R+58I5mh6pT4+afQpcEZeJ/uoj+LI5an3v8NI2Ggi89FN8B7/nEN1mqSbunBWyYJ7Ak
M989J2w807Ix1c3D0CMCF1450Sm7NZofgKJTLjGrhxl/PueX4evTacWIIHintUqeu/QiBJNhBtzN
tNphXueGSl3CfStV9hJCMY6CIrVfeA8OIVC1+J6Z3ObGVkUEK+QaQgU5DvWJp7mK0J+ubp0qTLbP
zmNA+EklGdEYhzb7l0i9VHGwNiS7VzJXpKQCAbAxvEudVubqdS26R1tzDVhlpeJhun3+8tpdkDuY
hetneDzqY18arYHZUsrdz45J+5nJyEnGbwBhdEa/++pFRuWo5ogOC7HTOwaiMymPPr4lbKX5MNPH
ENU547+KMk8L6AILCxExmSfF8iBevSUeFfJk/UOOGhJlHgkCkeKp0lITx0IgwppRo313NheIb8QH
QpxkUaCtR1VYzwmk+MJwtgP5G00TZQmIZIpg6mEJlZl7RHY5CHeDgQaaVfiGInsmUaFo0rBfTDWO
dXx1npsdUiwwlXGSHpRi7HFLvmm7WZip5BwYlSVOgrwuykPOXDaHdHydQ7IX8qbebsGNfKO0FTPN
g3YWuLRQ0Fj1zUucz5ErU5QR6iGNnVBAwtBdiiUCHU+yi8iAKmoFxJ2MhnnPjO1p3L/xq8p3LtkH
d/K0xa81RAakVu+jLIELVLXbyrS2Wev+9eesCvR45Bx+UXex6Dfr86fp+ttXhkZwcWvXg/3gn6ES
vNNcypkl6hNInJ2T9Kh4JWD4KGdkhCNGb04J1fYm4CqzVViMUmBHcCvTqDiY4PhJqDr53GNZvj9m
/sT65GSBYRNSf66tioDRJ3McIb9KY21EFu4W3oo2fmjTahoASi6lcBd70Ibl2/8FkJRfFxhVj0VU
12Dqf4sPW5Es5yvOlkdUs7WWJR3VegayVqIFs0kzoWJ/yuc2wlWater8zE9YoR9UaARMMGyVdWnl
fKPOZaNw9g0zVJuEarIfEJ78yhHiC4Horcjv2v/ysbXoV/Edn37/Ufky+KFLHY/JvkugrSTSDADr
T1UZd2yFW5MGqHSMbSHVWlddHpyTHnc1e+oDLruJ7r9m3egfqR0hksvFfk5nbK3kzsHThvH+MyRn
Bmye94XrS8LMGz7+ROSxT7pj6oxdYjUX/Jcqxr4B9ApxAzXWcy/6E7e52bJajKtt9Jq4B8vRz340
8U9HFYDnQuBBknsY+SjxJ6CY2ibGWgnrEQvzIp9BZJ0kDAi+x0OOcQkEzUzXmVqvLibP/MqO0Df8
2DJeikg0n7y0wKjV/hOeXN1EneQalxm3JE3jJXutE09gYUNexN2rD8/gf1muVhrEMCFx0VlYSNea
LqgQNPufGYk93d2SavYMSqMOvdgcw9dI5qtYAU/TUoK4mdRK8xTS7Igwmfda3qNhvZE28uSLd/zk
vuDpoSYxeExyAwveLxfnBXRz/FNudn1NTWd6UxCc91s8iQDO2YJZG/Ke7ETry79laOpqiMb8ZJWt
EGHMqHJ4GGqxP/5vDluGILWaOR5gNayGUgMV3zHH2QwLR3T7zLcHRCTItdoLv+RQRHp40WIYaLwM
x8Oyu2m20dXY1pwQ5L+95RhtVvjOeoVfSzX1TUDAgSm5gALzQPBTGFUD+J11aCDQFB6QJ/bH2ClE
gSnoaYUJqfam2xwk0n1e8RgBFr5lIJf+54HCiKZ5Bt+qBpMY6btvsSpiYmsEJ56QUrTZLjHOT4gR
b+t7mtoAH3AIgXZo2tvvJeE/eGJKNlrCz/yKYsvrztHT/L7GhOtqkcn9tAk9uqCp2qh335mcPd68
7uXH1TMWGyVK3PEatSKDvj0HbGV/F1kKuPIWjPbQHpkfzu1zNmbwyQ3STGsji7mns/z0eRP2t9B4
hsxqd0J5ZArI/ZF22xTH1hCHK4QtNLZl52UbF0EypKEA2tRvE3YqU0NCK355Y4yP11zuIhQaHsMM
syFQUGYJIInHWtzg52hG52NQ6RFB0CrKruHu5vBDzzhvW4u44x1vo9vZ91Hi/+P6Gn6mJ2H94Jh6
XMvz6dGv6nbluHv7mUp5KrPD3VzHoBa9vKkLd/9QZ44vN9TkdDXiDXNdWFH0QMoACx1MpRCQzATU
W61kGLShW4kQTtmkl3kmVmzlpELy1eF2d/RuuBxleN953ffcxlFln2pBXrXw6B15BxL1nMjuuYiZ
m7buaFN3WJ3+mBOhZgBQm8d8e49MIPgbUsV9Yr2LMk1K2c3CTNiy1oo3/Cz7U56WGyBmHmiC1u8r
yj5jBHdkYiUd+TTMrWeEat5iCHKKmwJSmJkKStsPVNFNDg+Bihf8AXC6g/mduWMme+BWHfuHoQsh
JGEDEX5pBoVbhjhfd54yMpJdLKUNKT/oWYSs5I/wV78Y/7e2xlJfsFU6zGDWkA5yHGRST6ZBlgLe
cWoOh+dJWCNzKwZNuD23dgHFi5tk89AYXo30LjMK4pnPxsTRGwzrKXT4cGmYcXCrYcA/1cKncdOV
LEQe+TUyrxX97uJ//4IDQXnEP+LoAfJwIkJJWDmrA4qoLa7v8ux+j+NxB1Z/COdvadXMpy8ioZmS
yPonldLypM15l4N9mNnHWX5Vu1d8doNGPF+kd3UUx0LFdHBQn3T4N+hfObo1KvZFm6cM2yXDAaVp
SkB7zOh0sxyQYSR+f8mIuoTCsc9DcDiPpp0SFi3hzHevNTZyYHhLLIVxnTVvRTgx8m21KNrN9XCH
NZEO8sQYl0zK5gWvW7waZ93AgZc/MYPXOdqKOoSoZ+HGkqxubcl9R+rCRgtfSVR77hdB77To2cng
Ys27zQhY3xPlTwCeQXyiXef2waJ3i8g42eDUKLvOKCE7P07OJwyIhf5f/HqkSRiGMcFAlyaui278
hdTMK3ffKYKFg07kp4TsoIBPfUOc7L3qwGnbI8CKDKuQP4coRXMwrVsspGWQ9Y7cSeabKDYXYAUU
pVN7eTK01emEm37960Bb6U1GV2vq7pprev4vjkk333mvT76u68fA0gIxn6/HyeRatDJQl+6IkTxi
JA2kZzGCuyYo0SYfzTqF20dXS1kUGoaztwV5Qm1vJq6AkFIsEeFg0/3Yc/0haFJyBQvjru5LK6xD
ObAcCT3Tkfdz39aherBDo0Gj7EMliaAy5gOKSwIDyCP7rhQmhhcUyQmRq+xgzA6tbogRsFpFjxHb
PXXSmFyajnMwE6lkWVdimxX5OJKbawjRLb75etdCDKgMwjrfGvT/kHO/mQ7Sde7vJTZ67tmLjOH6
+2/5EftO6YPQpqlmtepHkVnwEJDi6FgnYfXCQXkYFqOL0OuaUQPmlk+Ex4zS2oy2MYlVDdFNYtM5
lqAd/a3oTLGvsacZCiHhJ97qLDDEUnmWp1jIK4+kXT+enaCFQb/R9knEva4sEvNSYpGaUXXpK8+/
svNjafzcZRRycgLYcqo3WM3eU3Pzr9gXpxReweszf1C1CaNl1a1OMa2hvQRY3JReEdJPHGoKr/Ii
8OHzs6ZlyNfqGJcqnF7c7FH9jYj3realVSoTDXyLtnTZA5cGRH+BvITod4436a50iTlrpIlsQtZU
RhLthXpu/8dOSj5WyjWxylv6V9qHHN30Q5fvr791SN23Dy+piXcSRc1mRkT8s7eS8F7ywfPNXoH5
HH6s0E4JftzSSowVruos/TjS4RLXLU6hUFu8HPT+Cn3t1M79icK7wdg7Dqep43YKGB4R0P7iG/jq
u2GrAS/HYIxZwZ+IA0GSC0PUBt3UejmTOfTiFB2oyYCR8AJ+WeTg07CxctG9jnQO/kvoKHgOzDMR
hDMXMOTzc5cGCaCZQ2hr1eheesNvXZOK5YjwXrOhRgaLGNjTJZAXU6S3Av50bl5huMDVTB1Puf+t
3kmMAXv73P1OiIfviyUUY7VdFjY2IkFnome3+4CbKAVydvXorupJX5RGmyprsyojU2koE2/ibi8v
UWs21RGYicgUmuPydCY84ZW6XT6aOAgSYD62CfInbTgYbGJQ1+os/oWYdToyCl0263HFs9M75qi+
uGL1mIk/FjBlgAjv2Ae/NuuYJn+kSjuaBsfhKVAfpPPtwb2HSA4zNOZb7LBW3fwLRD+VUn1rosVN
55YMR3DOGjzuisSv9jkgV/rcHjx7ZtX6NWnwAT3h0+PDRPqxRXkxH97ScIOep/9O9BeX3WQUmGHC
u7GXxOQ5XxoUo57ylm/7ZK/4kVObqGpz9jrdb/yLuvP6853uIeShwz5FPM9l4MscmwTmY9Vzu2kO
3f3LnBbuhlalqxkh+Bnwujg/Cg5mk0FJZLEgSJkkKrJQ1YzzUbVu6X+BLvs7GVk81TYCWvPFtV4m
RaaYC8HF4PoNIYiggtxVGzmLiomTMdlF8owl7tqdtu1l4FcsalhadWPy0o7Sg95kmdMpp0xKiduB
u++tu5IyXgMIv2Yp5uAMAU9k+dTelBPW4K2p3sI6wWh+fkhuNRGjcjAAf5W/Yxj8Mkygaoets+ma
AruEWPY1PngMdoCYPJ3o/SKsjxINXeklWg3bMIB7oEwepUN9xpdSOX2DS0SE/UmJDsua6rGrbTuP
tSYxAHJY2MBi97sG5Yo+As7C7wlhqzKqItvwryLTCggFsvf4ya0ARfFnvHUlf24HhHKa+896+Zid
ALzuEeJzve8cNhZMxYDqXCBE9TMGA+M3mNXO8bj9LQtfEEin7Mtbnxk7z8AzzD0AUr+xpIW6Bx+Q
z4PCqzYiNYGhKQhxUNrHX17kJ4QYxb9PKMb657pNj8Horf7TvG8BfX4swcqZRY37pApy2WJaQ/0O
D+yHwQ8D2rv+55v89ogILODoCMQ/Y0BzI5nXzeCO7+cdNz8Gw2DndUfc4UPTjn0/+Kvoi9TFboh/
Svat2Mj8/eiYSm9C5bVf0CgE03ruaRBkWg3JufLwdKkAq+Ma9T042B58nly0DFSk964ob94A2+s8
tH2dJmIcOeagkwn6J+M7MMYXp794Y/aQtMZtM7UWfHYXgsuLIygQ26gVTlIKdGERYmU/w/dOavj4
ehkY366hK7iXnnm9u+3YhYhoY2C5vyRPSchTr1CAWJQJJCPjCfM1mD2GyP/y544HFol0u4rJS/J2
6hDMC1YTWwAsojmZZGdjcFS4Qdk1DypLXtLJiiGb0M/3XIRGyn/Fz4iC8OZO3k0C1ZPgSFhMmxKU
N16D/jqVYxGXTTjWA2AvaoKUxWfzeJamlR/RlXpPpmUupLNsySDUJQ7EtbajPXx7psg9GUGLOxlA
egXkwPqGOmpV0uxHpfmpvn+Pv16T3aIC330HRX8TEo846QKrNmfBO+EM9DiS8hXpdSCqt3asYhg+
J+pqkFQNcJREdlfpqXAi/VDYc9mvckEhUscMqPs9CwpaDzCF9zhKdLvCnCmwpqNwaoCqtgdu4qxH
OHqWupZU6T25errSPFpTvbbC1tV4f02bmGxn47Q2Pvg/tFsDXwPr2Sy9CPkIQm5agKbZFHLN+rlI
5W48r5f8G3SclX1cfw431jqiyS+TWeosK/YbXonxQwF4h38BeZwQ2wHbUkLHftRydJ5QJQ79SJNg
r9i+8iy4tuC8069Cgp3RQTrkdXmOKEn0co3uQOwRhf1WYQPuzBeRCbRlVTaekjK65exeBLv8Owqn
b9FB2Cs5pvHRzm529zJnr7Iey/lKp36PYtuYGpx87jVnPnAcfziytVtpNjCCnmpHwPkipT2zfhu8
2qsJOJDZdX3zSZtV627qfNzLNE2zjAbTLTcSOQ2uqVOmj2rjWoUnsbaiGG737EYx7UxzIfJrn9gK
fmft9vZ3bDNHKztW4Aqod4Juy1DH3tu8N7Q/q0V1rzZU9Xs2lQ4TidUXUbGdErrTha5RdYodRlUl
NaPWvHDnO6FYt34FZGySxIZhP1QJqY5aJ+HHAeWd09yRR2WBGZFcsz6LGuwYz0/Qqsgt7HSzDDpO
9F511XTVhnHoYuqsBbIMu+w2XXeyxkloQ6vzvtMyG4egRQIo9UCyN17m0esGHe6ShUvCc9r5s70+
b/oxUgi5OZgNes7rdG323CVkgyvA02zCwx0RD7vgsBoQ7I91exOGtCDUe05otI+r74+bWqkjyVVO
oH4HRCIrgBBHI1iH31ZaAuTsPo8hytMtst/RvAIYEuhFxSVU7fTGhfZUuigOF8xPzAAQhbichrG8
kC/kJCKGn8pJidHl+fWw2X6OxTyauttL8OZGkuvcG9ZAiJdwqAtGbkbAk6B8qvQxlIG1jAawF1JD
Jq6hA1VDYlUYLPikozfjR7qkqTrXgXgCa4WlzEjmzUuonw2ZAkboLp3tevAtu1cYsutso4SCyqsM
a6l2hxBjX/9da/SqgI/nljjf/516PEduSBzOnWqSu6o4g3T2dCEmiIzsJ3oUpBVYoyK/jlHc0q10
+UjE9kmab4pOyAIIITNy8bZdcCAyUq5C6vXMhzBpYg90eQSGdf2pEwKePem2gTEn0CiN4UADejdu
tHl9yipOVPJVlfc3vZn8D0MzEErhsqYiLJcl3IOjhlt0xe5idvcvEmxoPhhR0WJyU3ZnrbCwlTkG
01X5AOSS59LwY/f52DdT6hdORH93yVVabr0rsjtrdkShYh9wW6dDF/qoiholFdg24AZT3b/WJIpH
8gkvh7TuVW4Qf1+BCQKfooOy2bWEvosdy8yZFijLw9GOpZhJTNpxr0yCsfNLvnhuuoHGIeYmymAQ
IAJBys8cjxzNh4eFwg/FkIzHzclrNk1bCHY45DfJEw5PlTbPycyZLw+r01Tlk8sBhPFbZHRDlRaZ
oE6BZhyBw7HSoLfnvQwD312urDo/Yj7POHFHVt4WmH24+C1h91Ol8W8JNx1qOQPUdoXCcmD+LQSx
g8J8xwqlq2qA69/6t/F/WjnpMHCCd31SDPhdRQLGZxvoulU+Q31drJpvQFxd92+A+aqGlGaJp8+w
aRC2nhLLrO9ecfZVRxxRNcXuD2O13XMfNdJ17Vzk2rbADRgw8DQXn+6w1TjOqO+rdaXW0iczF79p
h25cz26uBJiAhWR+7i5riC9W2WJj8y+Sc+S6BlHFUm2MVUHpi36xmueaKjDeunlPUQPIjrsjszAs
aMHd29NQYB93MwTrhu6K0zXA8R5pMuJpgdGJCr3uN1avr7uFXb/b687Z9fsdjMqM5Lc02e6+Kfnd
HJ24UZmpl20KoGxWdasWjnhP0zYwD+P7WnHE07OmSxPEog+USPOv9GkZf1vFJ3lkklvWSi2IIEr8
nhFP3aX+X13H0e1H+zfyAD4EWbsXVePpNqnyxyII1C94/+6cZ3Ar5S8qPmjUtqYHkM5gt01NzLmx
uiGCPIgB/6evKhfy1aIIF8pm+wCxvv+EVvPB1/SK3jo8QSD1visLvcb/FD3f+H1fN4V9iUMDnCEf
Q8OPVtWt+bf1qZFNJppu8ZmF6RInKBsAJlgMlEpk8V4nTpx6wZA5QAWaZ9ezp7ZnD+kk4/JsnrnR
ocQLVGyZ5O8b0ziOcTr/a5JvuDr59puH5iDcGfx5s5ZwUmi6zbmbvHN7nQdD3oGc9JDqre9gLT/0
DCcE/igtkJknsPa5p8YQjF0BkIhqjlEbcP77dMyxOXhvi6cFvfwot/jHGVvwJcrSogNthC/zdtAb
ZHcGsp+LorF5gcVoNRck5lbHOZ2BvqoECoksw0/k1p7xPh7CV7ObowUm/Xq0+dV+atXvQbnfVper
cZzz/vY8cH+DIO6e5+mgrApgzQjPPQKoiU3R7BjLFdkP9AIJbhhgujyEGMEQiQDFRtSr+la43PGP
3a95yu9YM2rXybo/NNkigjhb0CgShAWnFBvUsxLDQmOGyeRyF4dhcE0Bwvb01fJxfjDXX4h6iPKC
wQxJ/VcFN8JBSX69IaZAflEEU4131Ep7qa/GWfXtwcCuN3JH0lDoelRyGKeZkoCeo8yl84RZ0KwQ
VdqtxqgpNsO0znXfi4u9HDdwV3/5OvKdbibaC9KMlYspZlGIExMWs3qL7PO++QJxHAg8twY6g+rP
DFBqgWexS+Bp0Bfsaxcyhz5zU4gp5uyE4vkTSqNP9tjNl04mEGd+cLK8btLmRWmeX6rgM+J1kmQx
wOo2smcF91KfAGLWw9RThc5w/oEuCWatUdfwAaEKI8n2Bzoh3tgsXIYulYDMY3jgMNcaP04pIP7S
5mh6NllvW2Y079oX5huFJgXlScuCL+g4Byjs4cpP63dSZr6F6f2K8ZCCWZgbEm4EYWVXMbL7N4Qg
FYjLSjCIGzTC1Z29aruT/mnfvEoonSMI2P6/DmjCWYdzH7Sl8W++EHCgIxbk7ySMBkF8yDo4npHT
ybjTjPBdayebYRmpXU+JcOaaTt1+lbXX04ymF8oPPGX6/3w/U2o5w5+znYtl74X7COgtXnyV9zn3
J8WEpx224bo9ISxYsUrF1oo8RmpklnSa5XgNlwGjMFZVyZnIkitVLHp6eo4e70lZhnQ5GoDobwa7
LBYoHcyobqLxjZcAj+GD0NPh58rtAmjYWvs1RjRqS2S+Ik1JwIn4eu0Ht8oRRfU4QDbaNnMBC1uf
Tfa86eAorXTTzJUPNh+IO2F/w/GHmVqpoJs+PFaNOIDHrB3PHcT42V3Tag77pitDqSBlrg5tTy+7
bus/2bNCtmbQ/mPR6VdYEQjHH+UDMyM1Zfy6YeLj5eLbkOFQrHQauL6D6uimuiefQz9NOEZBuo9z
tSmSoK7g3G36n/ztbhlHK6VnMVvdO3wFU0VlnoJ+1/frLCCiudjWy0Ebu6xqsvq2IMlt/uKH5Uim
BGS0iiluwMQxTajnInhCs0NZQuGak3pPiULYoFIah3x9uKsMfmISwG8BVLWPsiyVn5CijssJN0vs
kpz/wxNP8yjH+WUSB2PNqf88qGZh2LmefqMF2K43j9fZ/DpSGQ0eXBGlnFOGccWXXQuG56QwOHYa
j8NX9prVBwK2MW0Qy3LGEXOhcPAzXFLqnF70uFAeI3ELKhAdm5g3xfvwX6pQB3ecWP6zWd/8SYVq
f+fFLxc+XX2zzaBWF2vzmsaL7NbxQANHukzv4ltkDNmO4N3fM0oRuBCRfIFSgJ8E8QOB69ZRaaIS
wtm4RjsNCrqJZhWc8Ljoda4d0FvCihabbvmGYYVI7PCZ/DqtlaCwqidFze6V+MktnEFaoz65THtD
2SRYEV+E4l+VRHSO8FxlWLi2K1oBmiQ4XRRgZKdvJN8RvYrm8lHEvaeNQGp+lrXZJPD0qcwc2GGc
sErSabDrqpYa0moMveOX1LWPzOWO3FlM/eXtUj6UWhfb954XxPIqTgi2I0CPhsH4QnSOk3PY3J9u
OTTjrkUJjkJUh/x8OsB/RiXN511h5/3nqsVncURNZDXjXtp/52zTF6pBJVsglUrKxuNPlyvh2/TI
j593uBYUapa/dGc/ijBczX11QqOhvp8GFPOwyv4Du6ifCz48kVY9bP3Rfdg25XAtHCPF/Dp7k/Al
5qHeW0B3c48jde2kTnqvkSOBtaxsWMBlOvsAUdEOq23eAgUHe7n4ERkQlBljLeryUHQ3horHSt6e
ZtPMGHb7wrJjIjZ36csvxYP1vyRycInvH4Fdlty1SqDaFPQpwmwGkg0oGlpCYfEo4FV76GDy2Epn
FmAaSM3OvGMUPF1BjXoLBU83uLBlbMDrdlHtKsMyuYY6mvBw051Z4LrfDH3FIo4f4B0AvwJJZ5MC
n+Dk+N5cNAbs5vb3I7hf1NtvacDh/Un3mOOeRGsveVX+cgtm5R527YEYCkCs7w96AgI5X0hCUH/b
P44eDZucBKRnnmWnW8LOh7FViExnHG23yLkXNqPMatFQ7IBI45sAwQwgmXPtAh2zcMTXvHPwIIQ8
TYDwv247G2wu9TqcflJUAA2Ngk7xfC3T6Zqx6cy2V4ABb8KFq+xaR7o/VwSRbFlegYQ+dl3OWsmZ
edC6QYIvM1wP+U9VbdUj1fLPeo5i/RwUqobpNACkLnhyyt5iOEtvqpabNssrHX/a4CzSlfiMMjDW
nFxmIzN8xSqq+Sfdp0KtxukaqQMRyW/qbvLCgr/khdKSESUSuUwkx7bpPiPDMrPwGZp4h8opn4mi
DGAL4Qv3Dx2/qsf8qWwnNzBlsfhD2xRY5798aL7WKdKPfn/6CPwaFn02MTWvmVK6U6u91mBS+1mf
9wflPW3CnYDUbvjqlWS4rP8khs1lI+Vrhd1aafeOpYjM7YLvy61wEIBf8bmEndLmaRQAjc9NdBql
hio3byL2bGjycUe+vumib/HuHwzV5zNU6X3IHcOFWb7r6pRFPQgxO+7UVP2SarNg9IYfDWNizURO
QaJ0BB6B3nclkJrMH/fZa/hT8gqKIojN0b6F20H2Ve4VLiSrgsk4nA2xYQriiEQ0ExD5UlE4ozee
bEIyjNrSidN4lQye8HIa1mzvgiUP1prmCIJG4oMYvkv6dP9do8O9bCvFhZowLrLEU9wXMMg/Iiqe
lR60mrXc85aSMFaXlexXVsq3jqt/7R6O5sGCiTAVkB/LIMwPjYJh8E2IFv23nuJDBWTDq7Zo4+fR
37sGB/CA6bIB5E3Hfr9SWK93oyouirkwJFa31lOfGuC7f7jNZ1UrnnaPP3rRW8/oD2jvcvto44Rb
UEHqYRmeXjrKrRN66katjNm5r8M+qLg/TM8x3WWrhv7C7ohuaSQBQjqbsLgt5T2WJne24SvQZy/f
xjB38IKyk3sCreesFN3eTIaLoUYoua8Z6kmCdpkaTxo0TuvYmWkU6tPmxZu1T4/8KtPIg82O41B7
2u9zuopNS1Bl3+AdYv5qaKpGGv7qhjD5T75pzji+z1h+Z9o1QyTBFNgfi4E6v9hf3Sze0+fVuIc7
UfIA9nTckZF35iYR/qf5eTLKsJedyqpO0tYvRRAZyJ+iqX775QpX+6XLJ8nlucKCZFGDxVSeUDFA
9tcM07XYK6iQ3Bh/3O937VBGWNzkJs7xqDw+WujyJgE4YNv02Xh8rmlYEc355I9eHL9bfAPuJIhD
LQjk2SzjRr7TA2SfI96h5jucget7GKkyu3eOxLWsR53MEdvqs9oBD5hOXlO2MezLbpBVv1ZWAxum
aVtzwXXbFmZMtgSREAB2miqjUAEcxjZyH49Kdy5I3q/s2Kxz6xXgaCAx+QCTHfAnP+UqP6gKId/+
ESq6DEGFmcwgi/f20zvb7WCGMfYaqxOsE5OIUBgBeyKB6yrq9obSWKPb9QJcQlQ6XrtCnV2UQ1kS
tbOCfovvpzXhGjpXqdTkUYrf5SfdCgvu2EY2KUDvHyRXGMU9zeDlqF0GmAjmF/fhYBF0hcFDmu6B
ijt4WNqXRq6xRRj8GsjwKqTH3+CiaheBFhquB4/nfLGk8A8ByScvlvHNATXWoQ1kHFDWnuitSOEt
RAO/GvXuf+k7Qxu5I4cnj4yeJ3FANiUqhUkoCKWn5t+Kc7Fo6j1usABa5XJmyjQ0GARkGhg/rKPa
rhH9YXSZtgKLrogF4ClMUyfqcx9SkM1ekcUcZ3gnwsNdAeiSxSppHdUMcpoA/DNtnm4OK3EpvJqb
rh6aPfsjZQBEkAQ61Q3oQ5DYWK/YwsyuyuK1sT9j/R9FTLpeJKNZJaEjnzuzTlSgmKaXZIh41/Zr
q75XkAcwMNwqCe0EOougZdX4CWMGpdXwLhPyGA34XzvNwVcK0aYOpXypQfqYlzOkHChS48ie3anW
7uCTTDdNJsibqfCcQb1gSLNYph42yx4+JjGpesnltBHUOc/wShJpOWckNxFff68ca+5LqEiTHB1/
P1iorSPQQvcptB2OVniLYkdwZz8nIYqZ3OXCpnWLIXCDsYspELId+zxNJEizIpDLcrTP6GbGVME4
8V26BprxZ9PtdshSVhstQqmxm1BOmhEK784EqKTImOlaXnpeIyFl6YYfT/yB5ZrcqMKbO+mmsdWy
cfxpAEWpapG4d/IqXuV2GK10gyydZpVtcONTvgHprtazInRkRq6IPzDnPcnpMHsuAwF5uAf5w9ls
/vhGOLinAhoA56whbnD0c+Ww/E0lcALv+ZgTewAGMxn+K73N+OggTOWr723W8NwQIjomh3RiokV+
1PFKjsSQCWzkic+djmDdWSITZd7rOHx5OIPSEP7TRObfc0yfSMStJdpzTXUx+4NOp6VSn8N0Ot6U
6QfrgOYy0flDfH+sEvYQmyp2FAhaeBtQ7RGiTMbj07ZMaq5oeB5RgLmzsNKZvywJQ95AFTHAPUar
uVf5538hiH3rKRFnhOh7nylZUmABvbZg4F+Y/NKE1qlmoiJBaLJBkjvXVMggw+tDjGGYeyS8DqiF
15/6DSV2eK9ep93nRVXY9FwAiOHsqBQOVm7UZNKB0fsJPqeuP2RO4ZbVoGcuA9sq3DkVRLKsZJrv
NlCzOx49a36z8BJ7CjAuAApDAcJtf7mQ7psZOOVGZ/Jd7hozKRYxiGG8MP8O5UNVlZ92QlDeazSN
TggwnxisV5cM+vIqtjOINPv2TloNOig1QN3t8L0FNtPih4wicwehav+xPG4qiOTMHUVXVuX/oamj
TYOSSyMmgUHt3nffPs1w9N6Ntauvy7NJDpnW8mExUsblL6qz1AMhBv9kQxr5Y2vlamL5BehbjyJd
iQLwRih1PbG6oBjMs+Xkbr/Tu4V2Rz2GhqZwplH96nUkiSe/gaaFyuIw6pOk1DORcpCIo0MOQi3W
HWIbpBoxJD6Ts1rIElNGNmqiofXYQQVldoUZmCJh0OEr8ktpMmlH1kV8ayRFr4E+gfK7yudeRUPY
qDpbn37/SOUHxz33exOPgltZ4YfjdqGthur+JJfhKlsv0LTuE3FORx2tVLbRQ2Wwl/pNWlQRG4V9
h3qdn04loAIuTiWJvjJ02BOOzle3SCFYzXHtLmRHLTMeg4sfhYzHTgR69y32xQaTtnb9d+R6Js7n
Aty4S712ye+UcQAff51UNvKRMsNUqRMU5Xn3HWITIVmnaLpX854dTj9+S2kWnBBMkGlzbwul509g
7ZNUKvDe2vh7NpV6KQq0jPHrkhZ1ltil+0t7SNWROMR95gubDSAst7E0seNvrgundt/TFPUoUW88
pOK1dpn4e5D1hNlg/esYMK2CVPl+crFQTiKO2dnMdMkIQlN/7siL6wCuA/7ZyCujv4lRYcHeaikg
nj4SpnWLiQAs1wTv/XAv2ThRwHkwDn4jEl6IkoP2ecfztPWYeAYGe4tIat4xSrCqdIpiwcY6b/8J
/gZZmeXsr5jA/s7AkhyhDB1A32WKKOWtpEhbbT+i7bLF4FWRnWUS+CboZTBpDKNnZQ3WcsGz19Ot
W2eSd/106zQdESIINhTW1WlbzLVG26zg6XSpq+WecsJF6B3r4W8NFotpMBs9/OqFpdNpV7b4ALF0
WF1gi2k9Ak49n79OoJMoKXqqDUvLoD7dZzCeIpx71qJsSnOgmaKWXYEVeTSSqJuC85KMbQMvdkxh
AYG7p2Jsi+Y9jwt0AyvJraSePRAuhxZIT0cysv2/Ge7pYXhFw1XfnP1ZqAMSKCUVem4Hll5pD4FE
nsa/fWXlEvetorWSxeimz++xZqQ+5JI1U+kbFrHkQURTCvtyCi0nIVd1BNPFfAt+3N3uBERzmJS5
7Ggj2PbncpX1EVh7nvnL+2UTbqrEnJIRvxOiIwGEcmvpGyY7O4i5d1lv+474duKubM71W4WIVxEH
SqUlX6kLzXvJrsxGFNP9ZnEwIA1YBi+HOhZXP+a+Amf2IH0j1yNModJosLctGHyLsps+uCZ/wCo7
NAJuABCOJftd641Hft2aZuzZTSZZaGF9Kz+juRS8LAQwsbzmvGoTj5u0Uu5c0E9pEtrIA/o22Hme
5xLEn5dOSCjnS00aG4XWdm+dRMb3xUvB/aTpvh49WkPNa/a36TbnSZQ9zPTSW8JIzQRugQwknZvL
qC8OKc6KtH1VT7FlOY9m+XlCy8Oer6fnsow6lIfRq3SHkqbps2nYZO1NoHrkh2R9/rMNP4+88+bs
QVavXU95bsF6PpnVdOL9CjXas92nR+UYX4dRDLSH9RRiyqnHC9l6TXaAe+DG8hR5udcQ4L+dcIWw
DyPwv4APH7LJ0IY+PAf01I7L/lItm122gFzSRAouzeUSeOZA1C6mQfnevDfryqMhYoKs1MxaXe+M
0vuzCKceP4xy/fh+dd1Cs5lBWRCKkycJDBXH4eQDvbTY/eqI/w6AIAz+Wiqdxw3TxmaQfoLXxTH1
LHf4z0GKYg4hDi0ydWnl9XzRJ5TIxtjk55kFtQkkCxBXNBROE8E5E2xhAiovkmNuzTwCXEEa08Ul
WMVf+iau/cKeScziPwS2nKN5saZLmiSWotkXgrcAgGi/U8qk92rHoldl7UMo0gSHDPJoqw0YRc3o
lPImhtEdAf8lE9P2iAOf2J05LHilpetHjieZIQP0ra7pxZntOHOxU7KZpp3rbB9WwoQFUPdgBZZF
BVV29iaEzKDxKWBWo4X03WlfJE75avaytzZTMzrY/E5I72a0OE0iPBhkadvz/9spUlcEabz4aYUq
s4Br1/AUpD1z+xSe8fcIcuO6xehJbg10exFPexuOwod4ckh3pQORp2wpSP1t+HBhscwUkz5mNcQW
oG2WKaR8DWzEoRmqD3KmqmVz4PGb0we5rb29yj99c/EX+JiUZbONi/eI7XuAUVs2+QB4KRhQ2n7c
4cGgMrgWFwajrNEXD/3NAFDctu1v6/oxwdGPoOICV/ODnDJgrttuWKWaGqGwGFJBArG+ZpGXP4ZG
vTiHBjlVUde0ghISVj1qKcwnM9U5K/Gch1qG9ly+BjpXuV2YRXEKGKa3IXPN1pxl4M2yQtJUFPsO
HknoK3uGS8sFNKD6r/VA9C3FSNLCpMCJwtnkXOZXLotOUy0xqSmCUG6M+YK8OA0BJz1+xmxcMDoJ
ACc0zHM5vNIswSEg+CUTeJWiYAPj0Q+T/qUnxjo6jU2R+5XqSU5PQ01dNnwTyKFWZhoX8K5dSzeH
2M+8jUmALb0qPSFSlrCggwaJv4BbE8MUQXivQ2ZPUHkV4DyeboQDmS4eQGRhA19zrzRWLEYbuWrv
bGEmgUVW5c9quLPXhL2pgBhL61aazwscu+eIlfkmcxPDsIJeJWlTZrIwd/fn2XIL0uoQgaAYtBK1
uzlrufB0vdApkPExiRZauL0j15YmN5DjrvHanmsnfB22rs5d1KL+JuJ8wgM4rMwGidwfREQfojVa
hQM6Bu70yT+b5wQnOWLGexoH+MuRLFhfn/2HdiIRym//OzEGqRsWLTlCREYpC9YxiDU8I7GS4/6f
LVs+jNLJSKvxwcsMcjoBezc0peVDiTBXhzfiIScGn0PTc0kykdW78iFSekHKalNk/e/ZsIn2m/EG
PKJBiRVtxPVb2bQ7uR+Fjwj/hEj2d1x7alIVC8l3EcySsWOvKQsEkulKtHyHnClv8nJHKQWe+KcL
VBOIOaNXC0pHSp1RxERNbNlt5jWH3CblvMXi0q+teVIXEm4ukNyHzevhWUlF/Ypiv67Dn9f56xR8
melcQyboqmLTCPge4USIR4+G4YfOqdMY/wOYOWNEiAfwGcfW0zch6xhu2TFHF5X71G6NVlHKad7+
qEgGnbMaunsRDqzicrPp2uwswYxwjYKoGzHvuEyOZDwWwstSIjX6/TVQqkmzEgbCveCaBVPbRLso
OrCeQqJ5lN0eiPnsrG30/OyFjqyNKiE/4+No/ngvnBFmIC7LFmtOSTkCvPJZ3y6LHQodjwwKg0FY
AmA0/J6r0P6bUJmmaSNCjqQJVRN5IAcM5gTOatw5i34dLJVf+PCp6E01rzJYqiFOXspLSFoZwLSe
kPcubA0H03gY6lwGWYExUQqXi0heYvb3ZHc8tfLY2MAxtrz3y+8DVXlDz9m5VPZZa01mAQCCSlSk
a+5kWRTv3/4nLOY+H4kaq/X56/HtkV3ssI+bm8bI6HQtUyXl9RIDM/4IAWVMDQwjJA1qWoFIj+nz
t6+4uuCpotIFmzMmlx3ZLY3JMcDb/UPExWGV2Qjrv+dGfzQCKh5HMaw0fsmzDtBAdID6O+NNhP/h
+smIJe4DG/hmP8IbpGinT/tI2gvA4dhkaXyit3a66ZQzLlg9XC5Wd3yUPgrwVm+pC6e7T6lyJoVO
duAkBr9A/5ma1JZVPGmprdOEoJKgoSHR3euYFaPAiKQvvgx43NZeAfi9tBgIWLBjwTzSbqMegoMA
2A6ZRcbEsOyORJ4eshd/XokkuLVKfy0By+x2DaGvUs+Fo6VWaYzGW7Ud/+xjxMofB7OnVf71TDtE
Se/4E0UNw5w+5Ipi/EE6YAHsHhmqClmauTaH93YgmUtCReRBXsqkGcBqsirGT3QKR+rcT6uiSu0J
xWL0FNJoaGmWWWj50Uw4Z3OS5s3ZdvPucPC2Q2ZVmnHYDhtAaJQHuVIvl0PP1uqZ1rl5MvCbJwQB
kgev2pn8PN3o75aEifrr1fyC2KGwf2YOsntPM3FjmO8cxVOFz59PKtOQgGfKeKOU4kN+0UOZ1yec
gagM+/sbeiw+EbivQ7N609NGv7p7W2Pi+VfbqY2Eb69N+Zuu2G7BHSYBtsTpGEKzSaL2nCe2pgyQ
BYMSpNoKZhnHN86qKZo9vwr8Qh34VrnGBAf1ygAuTA2MzPGzPRLzgt2XPoe3vluXiJMooW8hz4ui
Wbb9KaykgiQby2MfVSX7FhUFvdxJlbQZZ6MA2UB5yDOGxEyk821VhXJKw4D6hOQaKJC1PJXyaHXm
qgc0lPfraowJJhwq73VdrgMWzYuaraU9bk4oORcYrlRwXTn0vZbp7wQc1iGGr+sASDEdheiuovx1
BAYiYIKZW9zbyxaPnitOB+k/kTl5VegMYw8v0Iknj2ylvk8Lfn/YfmmF6ndm9Ryn4nIPNGALYLOS
Y5PrUkudY79vmEV7u1zwZoPbLh2zOOQ7ir1aSUNbVA9CRgpilKTaQdtd82QAA98M8EoyopGxd38j
1qFqjUKl1dq+/HwEAaVX5e8WnIlGN+qU63q2jFfSUk1NkEm0LEHSRluSI1dVeFTO6nLgkxCdaX63
hHo/XYvSG5sWgLvR0nVMSTmNee4v+DMK45OYb1dAYb7bsLJUADHNlDNeWT4pTEwVBCJrtk53D5C5
PGgtPUZy/zZ8o0xEYGuNWgRgdDP0Q3jfmkeWPFDQljSgtT2XN2UUVGXAe+wHdeU1z8aLCxFqlQe6
n0QXIUtrf2o1DfHg32p4F87DwFVdRTbjZv7rNkBdnRWHJxN48VagCYqwXfjhk2cjDcDvUmJOaxe5
tNvaRLnj+P0g9avgI8ZCOz1nylctwMijBfwiuTEXS9takdd+On58Q4LvNpg67zHz9Fvvjk3tlv9l
Objic+JggGIle8PhaaTb7CYL2zUyR11+ArjZv68mU17iqXdoQgO0LzOvEDcajwA4bchGxa/TlQQ1
pa1ZSYg2kclg9myjIZiXrjdJewOthVWdbD5Lci2Oa92XRwwIFXAUv0KXWwujShTSvWz1Lahm8Zzh
uemCuXUUyNQoiuHdx82kqjkLmPiB6nuhNxf34rRGgM3APSxVtVSHs/EvW+Gnxbqd47MnLuxQViQx
feubiuJtR4K3bp3guuASvFctBzPkO5K8eOFvJMkAwCSloXwoHk1qLP6M8PutOyvV/H0v1YnBEkKb
d5N7DL7u6colW5CoOSjUzqJno/7vEwIhGaNvbjHX5gS/cvwKUTJ0ljyYDT3MPxucabef5qOFT7DI
VpvnpnZv2Cp3Rm5zBQepEbvOp+vMtzl+l0Z+ZTkvBVfw7m/ME7pfyYANPyDWP/+RQzwf2JZFVOTr
mlT6SY++zT78VxE3VVH6aCOu5pd4REWN6MWHpVNduwHGrFUOawcnsJlb3J99kLec5jrm3BeCF/in
wuOyqsSTNfOk7J4VGEsX65DNa1olYpiVBv3RGt55bfySbe0hjRH2Ub6Bp64KScmuLpnVc9Peup87
PFxGpistkxPdKp9DLTk9hZorQ/zP6w5EQShEl1E9kCNg5D8gBGkWdLlACQBJKCUqaMpfEelRb+zG
CwYIqKSzg8xmwbNjmd1qM4dqRptkaOf2UbkCA2dO4Co5y0ww84gQZ9lUnGiWqAGqMfGOsLISA3g7
dDrPOV5mcdgHjfbbxSM4NLhoq/flV5Gq+6fPyJ49d+U9/V5jUIJrDXGJ/KfiOcvI0/gOoCcqPvda
Okqq2J0HN5RX9otSZRYiArVkeev5zLQxQTrfOBZLq+IEIIsQx9wBp6YEQTdQO1wsNXzxtuDfcDSW
s8mpdn2VivvMW11m8/AA9Rts77jG1AnurZ1TgKSty3OPmFHoV9YPtPQ7lJYa8yT/9FNBIPENC8WJ
0izWEElifEkMVC2ZRmhfel0hKnqvR4ipgx35MF9XmddiBMn7U9UPC7pjI8KJT1YKZMjDFtKPqoaW
jSpeA9C198I0h1UNtRQfLxB8WJA7pUfQgNTgZ3kd4HWuNitG32JXg4xgVcHkUHC+nMPsNHC+PfrN
7GAMqJWVhSZiiz3Kh0P3anwh9W4IWznP4nx0WmfmnbFfzhkxUZPPDPUCKwHl/y66UMCbRiKpaAP0
4cFgrGsy0E2S3jJ09miTVb6hWwDx33G4qCCQsr/S9J+SdxgBGL2y1oN6DRlA9RldpmCGIRr9+8V9
0YNSbncvPmLnpQUZtcvoNfjdFth8HSgDsiur53+hUiaFjd8OypPzAEeRb7xIYHCbP0z7wFw+76ae
PHWamTo2q5tUCdVmFJRz8/pNzanN++uX37WbKTkCQCovKGxv3nWqD8HdrLZvZj09UXB0kPrwNx4H
36ybwdqM1rFOvOF56OdRSjy+s+1IPcwSCwEU1WaWebRQt0hVw6TqxP8ZkL720CYX6OjKdGNlnaiD
Z2GTXau4JMYbxdjOxeSCOoawcGDeW/dVyq3Ri5l/8VTENI7THuXY5Hu7900poR5WVqOrm57xUulE
qKyOu9H3+jcBVFsxjQ8Cc75OM7I5cZPr7a+fAos6uJ0NoX0uBQy70VHJJBevEfBHVAocAKtFEtWB
HlxBF6gSZBUF3y22s4R3TNzJaCqyebf+cOP5RZBJL25gofS1pWxfBMNlw3c7IOmAJWI6syxASevJ
5WIyu5fYIGjr3pej0K5yi1IV3kqolbG0dNuzxEaw3/ZOBP3+hG/ZpmkTiQ/AaYYJJNo+mf/4/iwe
XlxiQ0VkabkIfNHIgAt94FfOLcwlL06qjH5J4EwDyIDRS3UHFyK120n9UJlFLc51g6yxQUrQc3md
9R5HrSTKeJjlLSqNw+yLQTwJ0ZTzkCMLmh76SBelEDH9BKXZYWy7cp53Y0yVKN4dDh8QNctOnxss
mte9LKudQhKi+LCEpokckWayC5T8FERqije80jpUCMCKYM8odpPwSb02mDBZimi2qK40EaJjkDWs
tujtti6bSDpW6tkudOVoc7Qf2bZTe/Fn0xYBv9ohqYmsW61FIx91HyjxsRTPoTkuWnU595Y+HaCU
PLehYiKbMm+8xFPPKTW/dI/dQHBWfu8GwI63Hs+TXypbZ2MAOaIuis2G/+1z6XFiUZBvcW7Z0Ll+
ZK922rrDuQIGqKUxNhF+B4ApqqvDEvK/Is6XsZ2nv3w8BE7KjSyc8rcEbf+lV97DXA59Gp8eqNUq
mu5vbYDPCsDOU6k3eJUF/OqiepWx7E7Zn5tKR5y1b4p0Qq/JXEdami7ZitZNt1+QlVFpLeBiDpfy
RSyw4fhgTaD8/7rSXzx87WD7IOsUFdEO1OlZmUP/FcryPHcupKW5M0/2k6u+TGJtbnD2bFrKDGvL
7GWjzLAmiRhJ08rlWffE2w+6reg1G1ypxH2incae986xstrYWzvjwsEw/vfaX3O0CEUcenrPO1KV
7yD+/Zm0q0tdajFlf0A1Q/d3xl7F+ZCi2KPZhLemR0bJCjrmlxMqW3PwM2597g/dW+vE1SZ9ueD6
UdzATrNp6ZXB2CDsNA5ni1dsdt7nLK4zI52yLFTncX3bKbGclYjG4CoVlvO/AkbcD78sRDJp1cgK
/CUA901YJUr0TsksJSqxTITr4rXsTaLpaGIqTJ03bmt+5r8XLXFxVi+aEj/4/3PeuvCkiljlCuAj
Y/O3Bl9MlSkWF3HY+fTpDIKvbbRNIr/KLAmY14YZZrbKXgIRDIGFWmqze+1ssh+RmRWT1OksgQWm
gh+kJ8mk6JDPfaXHGXCaJ9IOlUZEprR4Z7FRCl238645bAoMz0mHU2oIqyuLajjsSRFSfO1qNhfP
PqZxoRHCaAr3fMF8XAFt0vlBMaDYnC96kEKkwk9eXGgoRvweoh+RND7HNz+wmA7d1FSnLaiVQCnQ
IlGBJhi7gM+Mt+D33AMjHvBQ0SXO+6yUn1VYxrv4Cogj7AKX/EEkk+2MO86t2eL5MvrmhzATANMb
wHRzLOj27sApQAUhgsrPGkvkCPf8ix9dxsr1gTRjy/+EVQAaoAcwvzgYcy6+ALSJhoVE6b26JCgH
4S3jqDgRKvCg464jLc8WplW32XjZ2s0Q49mBNU1o/uJ/+WkVyKnVfkapnpuAuZA5Egcz5PeI2nKa
HoDT+jWdMPENU0qQicyntvayMor8RpT5glbqpLIcI5DSd8uLaMagpXFc/T67yySjNpAuB+0peZAq
GIBXNtr7HdyaXmjsrS0qxuKi3h5X/a7o57uai45QfRwApNFiwHAnm1Qju16Q0sFE9LlICtepS3/j
pxjCU+LVb+lelUbCTXuG+ytuvmjPUEb6o11Sx0PblsSh3L8Z5L7pjaLp6lOCyYjmrpH8epIwRj5M
6RtgQV3TsNrIpt2DlMnLDrElH+SzNmPuQ8UXyB5ZLp/W6UlyNrzH0Zp4MDMtkcUsnfiBHcxLj0CF
1p5Ts92MthJ7en0poS5v9tsJuyra5TtWlM/DccbNqsyAarMWuguWnh+aJ3NpzR5hYQ5MTfKyZW84
1ZZ/DYj9VpWWnpadTrsKKzXvDguJupGzQ3tqqc24aoaMjmDW7xfS0HDfomygMXmqEbKuoewwm0qU
Ubr7nArKj0aIZXvmmW8JHFgdd6pbmO4DU9gY7z6iuxcoKiIxyvpzI8Fhs8aeTzMZK0SXHIQT89B9
hvhZ71G97YJYecO2iyAPKf9tv+VTzpJQtvz/ZSEay6QAAH6FB0mwgmRE5wMFwn9BUTy88TSwUNBO
nnLZvZQ5820OWfAc656eEpamh4M1L39tc8MxLFAwwmDgSYtGliz5cyww8yAwF3MvXbbBgyW0u6nk
Ql4RW5AjBYfbglmShZ9jVafXQD02BiXg8Dyb+hOZnSSGtug7IaYPq8mzvhxI+54e+oBJDCimjZEk
lS9VGhGcuYSB3Dha0sDydBHz7DsFiMHngP1nL1oo1lJqwbedQQz96FDm9YLVHIz0+grOYdO32FeD
TFJRsbiljc3AMfvR1KCd2AWGBNOWCX0oCH7v7voV3NdA9dVOkSlXUC9lNGlhckpzJw4IMvhk7vTK
OfxaVWbiB/CQob3UGLC+WHaxKRl33+jTqMSDMp6gmTagmaL9mKystx8TqXVUgE5yBOX0VQJFbXkd
DelHb2ATdeu8WK/RKr+igcKYQoIOKNotjGGsiAK9ops5e/c2c14ZgL16A5Fzlo0NbMgOsO/dHvSt
4H7JXKHrWm2QDfhokczyIjrP7H1nJ0ad3wS1WmOINwP8BTS9SlU9O3W400ITTFU7dpUO9GQG6SKm
o5tlL9EaLt1tHHnqAnSWQXhlyjfafiQl3SSmfYBzA805uCSQZDh3SmL+wwiiykzP0nv0viSotVUZ
p37mIzij+p169LmRS/yQzLnbeutyXrNHP5wDq9DT8WjpITzNnCsS03s2HkimaT7ur6SN4hZcD+8r
EFFIsEWi8doIBNQhFCFRKlbVn++x/BGsmdKfIxY7QkIyGWLwFgNwMgQtjCyLDo9pVCqlmzT6kZgd
/mp607K5Fdufp1/4lbwazifQD8QYGkgEu4sXkgQKHfhZxwL9GwJsckGH7y7bT1rUnLYU/Be/aYgh
TYvUWk/AuJo662Lzp6ZpuCbgM3w4s/gGIjqIkx4v09E8BaFU9UkWhb60yf78y5NCmy4Fg3NpD9Th
lTsQdq3DrWdCBCw8IUgEWjFveQ3ecbYof4/uQoYR1AwZPPmujbI3xuye9+yOvNMqOwL78wHjR+SE
YoqOYCQEk6II5wm7mVIkB6wmUTDXWxKtN9LYxn6aRCiVfMQw+abZZ3Eb39JNaADNaWsrG1z6B+Uh
TWEO0kSnM8aEbADDjaHzX4riWG4eEoeX0TPKlZyU0BqBLZf0eP5IrUywGz8z06eECpu+o7AnDD6T
HHg/a57mODlG1yjcWhUULMNrYobZaYHf+g+2ntnMih2vixup50kJ3zvq3qmYmA93TAqoAdiWTGXD
DHKhBwTix2liHoxDwZq7DzIFY1Y/XMQg9tma+l2borHSRxFJFyE0nW1eGub4Al3tXJfytvpD2iB2
rlXhN8ht7vv0qQyRjhkOZ3TN1srDgRAF7EGXlpw11SH+/wxUwNSdgJg5ko+zQlna173AxzicNsT/
EGjNPFVF5is4GC1abRx4wQYO3ZivBTNHOtthBiibYtvLRDaBs/viQT7Z2K8K0/6fpX0S6FWWxKZd
MJOx1mdgkY2g9vGCGBqIjQMco2RlsSXTI8svnkvWMPPSdZNlsZNxF9BJv1HVp8oMLNjshKTJ3FZx
/L9gka1IwRA7La4uzdxpOcKXK/zXytHqmJ6uprYSJFb0bJc69PItRhRqQWU2y7GgwYT105LXQnsC
WwfPbq8w2ZsJTspZ7NnVw4fWu454HINNzVQBofQBhRHY2H3aSgy3If85ujO7mKLfUwgo+92DrxNW
nTBz2ukbxYqSmqkaTnicrG5Q81IbkAbcd8oRn+GAa283jcnjC5p0BvFcvmXvvyJyBBwAmCyJ0qa1
xfq6qXIXDTbMOa247BI7uYzNzsvY2K0G8aeE86x5GgNJUJ8G6smGDTY6/1LnF31nNJ/o48bjxnNK
DuS/MiSXlPC+z36M0YlrdJ160CNby2iU+0jdroowyGp3GOqd4KlmQh4iOgEnIfZ3go4Y/gg8baEK
sj8L8XWc9cMJxknyoqxOS9nJfQpn+KpJ3GSrj+iv+OnpP0agW1SRV7wqEdrtbxUMrVxhNHL44Mw9
zr8d6znFqiYs1AaT2yfennOJA3P0IGaIF3Qrv6BUsLUXAGs0uNQIFEheqQsnFmgPgw9e91x0Na98
GWReSnxPB3UOrmwUqa4GB4Oj2EvSVcKxddaZqsbElWY4v5jXeunmAtr9TfTlYql8QCNePECbJ4Ry
0Mao/hROkpYNK2I1fRNQVTl1uVJ9bNpedLkH61kpzvuDxkmySe8vL4IwyxacshXVG26npz7gVeg7
nrthvpXbcnF46Lr8/vIWXXi76Ukwht+P6bugN97qmBh/dhFXlTd5JCdh587+OCmYRhY70LNmVVYY
0s6g8qkn+BYqUJjAN35HefWxnjXmIHsaJS07x4ZaUPN133wVQY/d0lEn05grao/Sb/fA9586dmmJ
hkY+8809XdcdnMqKIJt6SGZndaQEYWHi/QC+dY9Vtljds631eIn5khtXiUvtKzURLZyaWAW0K9/O
Gb94ecvmzc6UXpEuhX0Adu5tg/3hGyr63Q5iY0R/I59YQuKr8N+aMouOMgBG+U1f5gKVzmZHeksv
m+uOliLBzBddVYLMFVm2v/JquJ4/ggz1NAmYoLZQLkZHst0dQf4C25zJAhrunPXhbjpJ1oIBmQ2U
yiFi49J3MDZ1lKR5XrI9maTHk7WhqZIxTHvpDfI2YLIjp5CL3ipEAq+/AGvJjcYWDZVejFS653Bs
FoWvWAZlPJHeN3A13isdYE/J+B/ICLDGcNGpx+7L4eym/gVRa+uGwpBo5F5rphCOQidbPsQOLRiH
V3nXuOlGR4gukhdkTXxSyFJnjdxdinNYru6OPhaEeEk7J4mt+y3bLb7e6c3SgQIEahfp6hweLHRd
eXw/j8asjGfzjZ/IBUODqdm3gXwxu97V3aIoDdYV9ENC/dkeQzOzOXjgIWQk3YyDOOftImF4qSGc
QmIk06qKwQ5w8tE6H1sY8So325qzu1B7YADf5TeDs2jbf3rjW4+WGhHIMjn8OnPiiX51ci8Cysih
I2CuGkSEg2wGMg02TCHTFPlkXF6GPgZQmA00qggzfS7baJhs9hz7ly/ljly0s9WgNewSkd6agkxZ
PwTbBud5hyEloLnkuAtYlr3K8eOD9OzhhFhAKXxKaVedYAOiE3h2HW325XtGTkpTvcFhCwicP1Yf
NcktP16lOZcKAuXeGMuaKXQ2/3LK4+brFTBNwQlek5pGYHNwlfVDrzmKinrRsnbuBE7KC7Klhtxs
xw4L0Z0ZoCd+jWNMJQUZZ5GhGiyRN7KTUbsv0zcHvlGxn93cju5rDcz7RrNzFs9IiOdyIGmgolZI
0IaTo33L8QlOF483uJI+Nr5LmzGhk6Yt/foulkEgyiNx6vkQ9rCqRPTmLd+3+of/uWC8PZkRVt+3
kshpKQuOxOoEUWN1dwoyFIcnD+HJrFz86jlc00PC8v11ipPc7ocbv5JFFpBxRyl4j0QZNvqinqj8
GHrpBvL733LQ65QgZei8vcSgEkIRaPRNFoClQ+1X1At88xdEEUxuMOf+BxkAi1y9SKANzQD9ckth
7Fi/zlJQ2fNE4Hou0ECYrYjytiXk7RNUcd6sWj6pGHmXoaEaQt/Qr0HafHki6jBpCaw44ridzZAb
2eGZwSHPzd4B6pCn2Eg2MxosTpH/NbZekVOtdeHdjlD98Hi3ArUf1hZ/ZqqrzJyAOOTglgOIhnlj
Dvikg/lz87etLP6xjQ+B8Bpp7bQno4cgsqfmPsFIioj+4ZCQYDkkH5OmXktElGDhOHKrUY4knlWU
DVD5P1ANYq4iW7BgdwDJNdmGclSZHBdpn7jKsNBGa0P2eSxaIUo6cCCTFVELDOcZ8ucMJPlaWe/H
CePofn6AjSI+t2vVben34UV1JZM8/RcNJsXIrSo9OPvJuowCcqbkSSQ8XDP5L1kPpS/3zOWFgdHD
RY3cVIVU28+ott0TYhYS+EvAHvYUWYlmr5as+VqCVvZ0aCOGVLsd80yxvzmBwdmtoTCA600Xw6sE
yi168wA+qFEZpIhGdqVa0zyM+faw/m6sjFil65DybNNv9fenvmVCF4r88hMIBMDN/ykdLnV52VoC
OHNuyoJ3PBXD24u0IUOkzTl1R+eGNBXbIU7+H+t8GHjN6YyOEQscSYaOtc795oF0wARmm74qFLXJ
6cfQDgSg0OKz+a1bfjR8TECkgG0+9AIx0khvRC2UpLuOFi4jSyBoUG3z3ZS5b93vWm1wrE8jVm+7
t//+CqV3bxMTSLO8Da092bW37le1YeUcYqz7LN+TOfccJEkUvaOJu+cSPZM7TFC9di0OerDYbi6K
5RN7sK0UWmXsV0Dw11BqnrZKldbt7UmZkGy7ptF/SOfx31ZzRmuUSifaFtrUe52ohglYv9CJ9YY6
tu2PvH038CNO+NZHB9hbBlShNpX9UMuIZiDdck2WkrLx3ITqrBnC7EW8G7oVymrSPxfJ6PDxW5XR
blqrBBaMNjx4DyUtiG1HnspdFV2e/xb3JiSmTCdoT07JgeLPgfwAQurLJ1SpEzsC6S0vpuJr4C8K
GyiZ+JEjZzyE5SlqrfPswKoBihN2k68yKOxmhFi7hBv9izk57ZE+aDMN3Cl3vBy1x9aXJOl0SUqV
ExYyOlkmsUzGo1OSVDWxmN5E/JIpxYB/thK3OQc9rWSA5J+C2IzO3NIhn1cf7iuYwFpMsviorffi
hKEFVlv1S8JUgTwWSyM2Taqezqn6V4eDPOHt/e/axN10Z+gAHK8ajkE4uMscHIKC1B1k3u5Gfvb/
RyLv+TKlM8nuJl8j6zeMxyxZvnhgUkJx3sm0ZM1EHRdXuv/z+B2WvEtj94na2i5KvW7QHz3GS2rX
IjjvKyysNV5ML+UEDJYLSfSRItfJpf2f5EQ/3kBbG1hkoEzcL/hVVfwsMIiyqMHRegnH6prvHES2
bOx4b4gPcCPg66lpwaGp/cb+lz4B6LZ0covEOZcX8OFZ5Lx3cBjuL4hdsHtITHTQ356paLtE/kRQ
Pu+UkJ3/VuJqZPoCqaCxNE96xcPYxgT20EkrUkoaB2e4SlIUQRUS9SIkUWqjZiAi2xixyzBsbhVZ
H0j74uuaDtBSdswfYGoJ21ORHwAAmrJyRsxUwvZvnt3gA22GMmU7XO2NQkFaumVn+89OFCP0xL6z
H5W3zcsKxAuR2Ck/P8ptCVOF1qpXub4Fl4rNh9j8VzEhiQt8vEDlsRmi3YduabIb+K2GwYPPKJoj
vTXErBmM8+U47NEYA/kOnwupoeuZEPiThoW5/rk/mn88+JzdjpPsX2MfL9BpT6+a3k47EdHAd8lB
D3jJ32m5E/dF8I4mVR7T3FWkxum6SKk92JqCyaLt1fQthlrk3NG1vGNeQ8HXuz6q+SM9oQ/28PgN
4Nh3fwTG9JqTjMhZKzK4KwUX13mzm90rC4kDXIIs7tPd+0TyDwCB0uLBke/6QYopaNm/V58M6YOJ
CIuE/Asz9gCPuACkr3jmapePd0Fuq63kVIcD94/StetbUCAfF94HXQvRXEQxrWIJLvOhsFBo4mNJ
wpJTyMpQHBIHzFv05/+1bHfR92GRG4YHnKOFaDyfSd4E7IQHzdj0pFV1Crh05pTdaJLBMTSKmQnS
j9JNyQMZ+cfjGDWVwFUXH2BiVRVOcvGaBvoZzR10jJpzAS0FtCrk6AXoYxkE0EdbSztDqF9wK2Yr
c8GH1Z5vjGvkHvAP3+QBiVb3pcK0EMlN4zCOX/dc3kZKCZSyks1Mr0yyFnpnjGdeaGHf2NpeLKKz
CxI2iCO0MmGDqsFcgkq+rdJPJtRI5BhTO0R20LpLwS/OUajUwHtbz14RpqWdh+B1ayuyYqU8BuYv
HjmpBDF4JVJkABhokLSPH8YSDvCdy5vX1fBwF5h/LqvgTiqGaEtJjn3H1dqzX3ote96XkwkPynF5
zaNKE80lgWFKa1+DifSp5OSDiS3utZWwX4aoNkQS7ex+CY81Iy3dYl7MbP/EPqy8i1giPHpXQEjx
SqfqzwX+NXR5XruSsyUCP5Px7smybdb4QjiRhUi6k3vvDkuUalURq6ix6vfoQoHxnM/oDK64O+0p
IJ7uksomEt/CRLFo80jvuLRBOcGpRnJIAi9fsNJRibDyRYq5HFqmJ+8XYdfuNbEK3e/c+kn+rzqu
o82NT+KYNiwa8KiA/zkd+L3q+54LV3Od8ezYZHCezR/y3oa0/TgNlxwuMD86zhzWuN3aci407Swf
hSGNF+j8BWV6RvzE2hddBXu1i7vVknrNVwES3lHzAkRzrkfCU/IMGS67V2pVTWmgsgBpLEFBVI3d
Y4gvTVr1zmdTKQLfDYEeGkyEjTFmMUrY1CFrpM4qtVvP+ASI6FWoFccbMfxayVb3BPW7+Q3h9pgI
68lY8MK80TM/DYoskkts8WptfvcVA/NDPyWJ84oRThwYFl7KfTgckCSs4kd6mN0N7LSmjygtLTZt
3gaQOSlBMPfBXVEPvnADIa9plHxU43KBcX6TzTwrpP56aHeZQR49XDxj5tcgXcmSa2JSizI5KnJu
cG+dpjghH7TaV0MV/o0mKkzw9ChRB29qsqrBCSh67k3vufMj8NwO5GWA9pWFYjuyaVbFO+q14VF7
tYGD4PT65YPP756Sjsgo2okhnPXaeMEJzH67gj1ZhVhLD6y0K5xskfmoKim/w/TQpHBzzKe4X2Y1
Z+sNsdIa8fB/AvvrDiuzKaf/b2vlGiHo16JBnjkN8SKMXZTu47rtay+SdLyGiahQOFXutWcvwHW1
AFkE9u19I5Lwta2jUlMVBj24SD9twiZpAY5AchVtlcAvTc0F9GYZsk0jEBBhPww2lkElK/dZtUq8
QIHWT4ypXf/h816ZhAN1mzXloGZS2h2z5n9sxdlXhnJqqxMY+Cfw16ARIdwY6paFKGVeCKbKuSme
eAHKSDYNkJWUjKbeuBIB9xInrZMYVE4SCZkjYw2QgBt9JEaTMF8g95oU8XvnbE7ZbbtbztAQ88z8
LVLYmnDEPU6pS8lpooNtsXqXByxYAKsmV4tKlSYb6yyQpuqjfpvwXxtVnzRKaj0Sdp8wz3elzV9F
s30ICO/DVXB/B/cpjxrey/qUeKwDFGZC084N4ovG3DdQHlh+h8eFTPz5L2VvqPKzUTtZyau5p8RZ
lPlyt18cjdd83XRQMZ8j6w8VdAHqkO1uy7+VQRYc2OT4FBTrUb2oLIb4oQCyR+m/wySfbSn7jYeU
my4chKVnOFulhRTW3/wHIu7qIhA3MiNSWohQ7KWuPs2vF+9qJv3hZh6aAMPhDSIR8DiRlLpvBhdk
qciN1Sb8OftIHXf9WQc+elGQdj3DZA+EBfm68191Gr/l+CcxWWcx+F2ecnRuqheiF2VaYXbMgk0L
8dGczQNAJt0StnHsDkCaayJ/8z+bQFO22SIq/spVc8wJvYSvQ2AovXta0ildn7tyQK0jTP3l+1V9
fZLvG36XkBlrYNCG7wE5nXt9dr6XqIovWiGk5LZT0YjlkAbiY8OgeLD12bNtfn64QQa+pp3NVNFW
RDc3lVNfyiAkdWFfot8UMfJd+7TfxFuIvVP5qA32eyHTv9WcQ4UEEmgJdaBiLVOUB5oUw73S5jSA
1imNSTfpmx3dSDONbJojCQwog89JZ9vOhhlLz+EU5qaqDk0GdjE2m2j00tZdwULJ7zf8brCeVj5d
kqt6YBAk6efcV+YuZAOsVUQXBDkPcccSHZFZLM/C0vGEG2Y7/aHppy8V6/OGwPZNZz6j6iDtT3kf
FAfKSoQZAXZ5Xg32QzL1M4uOdjkFsDDNdZzOgyYA6usWM+TtLSCYBQUgLaKRFF2hHBVyS/VqIj69
vxlZQOuXgpQxJ8nOcpCa50YP2hhZuDubfE7wbBz6XZ1SyLEo7nF/56Oy3w9KAt9mHMFAYRpEjkWL
qtVCR7Im1id7VFm/Vk5G2QPEBLdh66ZWgWejbG07wydmk1jJb9P7A+rrQ3LkYe9jCwROEkTmvWxN
cSmXtrQgIjq6jcNvw7F24VFR5hZaZ8HjgruE2dXjGtusCbO7KMtorTXbqB6aBbCBM8w5wSRIFGw8
BPp+iKPR39lxQu9aJrmJqLHFsZqs81oae4b3tVDDhXAW096wbifA6yJLvN8qv/cTZXv33IVlLHvS
JhmZoT+CTZ5lOc1oaW0zt0KSST2EwvrTWqSsbURDpFuygEHXIkbrBU7ixzML2fvev7jJuy6M4fk9
0CuDm9vgy88Y4a6utfSK2TDNBTMKXn0RUajLEzFaTb8LJ4CxfAhea3TYmYRhaJVXLEZ+rkyoZC/g
lcNfhZ25ARWDI5FHxlvRKtWMmzhKKzaqZI1y19PHJFJPgRVPRUkHTH4JT2G9FRZCxBLhIbSsZtvm
M6VZKUqQ/enchGqmwNDRckNALGATvutCiQ4YRyx/zDtKZbZRQ5ziLIjSNKS8EQSxaMFVJd1lOnYU
Pu1FC/cpjJYajvzSxYesUaaigHEuvwBRsKbiOpQzJMqaMOWhWEhVbA0J+Hvy/zOGbw97dpoLnBFE
g0kH2qa0CrHBK5TZ4MCofvEKNFNzS0h8b6fvvjowPj2Yx+iB3kgaE+okclpSH4X/iQqI4sbgTXlB
FkusopME2MYFJG43azInt3a3NR5Y3eK8P3x4fv5bj676VBQ2O8LQOUXI1p2ZEkSEdcO5s6r8QZOx
4bfgBK9sBLM47XAiwJs2wpXQIijI40kLduj7JwGmn9NKqGWH2lQIvL0JMxx48NygiQufziJHbrkh
IgXtLbhVqftCg1fIgvZbNbDJUDDTKveu57oAeoIfua2b8aSofRhk0p4aQJBotOVIOwDfRCp0z7nb
3N3/H7QI9PgN8qdEtJkUPTQjPzCEUJRf9y5B3KDlpBvAn914cHwpxsyu2wAhdDpp0UlTaTM8tq3N
nT9YVxwzKwnAfuBAoLk2PcnCYtqJhCDLcZmBDVtCLCiRYhamD5WaLDcIjz7fza4d9CotMyFkpSy/
gVn0IskXbOpImvozTsRCX5k6lSTB9t6ryk0WqCehOdFQdxEO2w8qp4F3dytDZEVyUKyE58+MlXvz
kWsRHnWfq/i2sbxGDREaw/v+F3GLd31xtC/K2gxgAwhFWecx93g766hXHg+z9N8nct6xjDZAGCfZ
ZgGOBZ3lPSQEDCi2EZohd4YmGaPzaImm8RN9gxpv6OIGJtzyegzRmR+Gq7lY8YgJ658hXdAWyPJ+
cgcgCtO4uaZqLWJro8Ig0GjRQmNnbeaoNDALK5iJE0PUD08modgbYKUELW3+1Z5s6TP/LR9g4X+5
BPFEv71aW2utgJX6u+PKi20AFYWpR5XaPa8LJbCeQnBIzn28FesHpJLvxQP0LykrqwKUFuCJLOvB
XYmS8p3Vuv+voqaPy2STCsaH9owbzHq2GtD2j8nPs8RRi2aJyf4On2rd5InH61+hoatOrdtt45Nq
b3/HEcE4rglBZF4cewavWuncbKMbK9mMAklH432JnIY4sk+Kjqfec1H23e3Q5HtcGiJBWOKuOnmQ
yJDw4CvvJFy/AGyGXMnqA6ZJCNP7UMBPcwHrGWhx04XcKEWYGZNR0JYyjuzodkn/QvNFy0/MudPp
18wNLOtcX3JaWjsHoH+xGzPTaRb7mXWMzkn50cR8BDsGK5mjx3XF7pTMiixLWX/zzIozOD3tvJ/M
H6PfQqnEPusTrhDtt8BfUEGP61z+vRKo5s5BHdaSkNr8xQrItMdyMQrI8mjcvcbEtfpM12uF0MWQ
pfE6+BZ2h5m6C/yaj5xz00E4Hk5yODp+/u9TsGwflVTYWeVcUo0u84nZkTZ+PTe1XeUkPR4rH8li
W5nO6YpFHpLD4p7ktPFNxNS5E2CHPQWJS8eMFKaPWn3T9zGXbt2A9eAQ6cSi6bAP5CCKulfB+jZr
uiF6+dEpJuHZKczDYfwNTrJQqrTA1ozekNVrpmRV6ZIAMJXH/m3bfbKv6wuwEX8I5t/zEjjtO85A
Wx34w3lN6muKmFs74jthiffn6UoFQPP8OzTFvnMu2JkZ/kw5qRrjoBiZ1K04Q7y+Y4tCU7FSAjP9
NLiNxvNaYxKSIovLnYNnu2PujnbH8Rs8BpcBKMnbXNYvuzY0Z7Aa4gsL7OtM4t5bw+vWIQvfKlfS
BbkdibRppkuYtEPJnPCBitOlLCTQWI3NEo02beyjErUlUURtru4wyTUDXbp2jd0t0kboiEDis0Pk
+3IIcRKUTjv8l9UL5Sfrf+vDjf9pfU5QITL+rzEYWdBH5wpv4arUWB56cSwaz7kMYlNBQZSp8+MW
IgQeOuDY41kvjTJGf3nZ2oEu3rPbuM4KKPM5uP8S+mhA884O2Jq7Hsr4umJMt0/tVYPc36pB9wY0
5gRR8bDptlQVZcLwH4KmGVHEu6wHdEyq7wBJdKBHj/dLuVYghqQ8Cv9yLDn4QKlRC+D3GP7RtKp8
YCqgBeXRSKAtSZPWVY6wOGPG2tKB+6oRNeZuOaLyFHb8Wg+XmlQXjDx727kzOneLdPLCWDp21w9z
GMuUv6+r5PX6Fmrz0j5Y+u9S2RLYHeJVp8v6/Uh7pMwRio5NWapRB9uxt8+1sjiJ5NUlouaegcWX
CzG1lM1lCJfdVkisUhyuKDrUv8ZitCMKWBY7mhH4b49BhsdVfS3OJB3myFcMHQLXC2Gqko1M5knG
6CCsgFvE9RuRbumuTcjQx2Gkbe5tCVINXvM4+BvhKlW4TS5N/2tUdu9S4O9z+T9b3Azg5TWqa13r
2rTrh/zKWL2oSTFbGW7BvaXzGQgjVm2efQpRSxklgVq5jqg0jLlA0F20vPgGBmsXAwY7k8ZrSfB4
7BCbG5EgMFKIzwFKPKzfitb8oS4hNYh2QH/fYPrOyI48QfhOZtPCPiO7+joXH4blGVYg1tBj2y0J
kFCZ07YdO8bruZREFEJm5ncD+ZuSksvqJaaf9CADM334M78CAZBaOdYuB0E77OKEEMokiFyZ/tJl
yfPmHcEGC8FU8e6Gzn284zo8YW0QU5vh7BOO3KC5As6+t9ULbSYGz/of1lCDvUfK9QOgbBAjnMjK
TSvWLtHl6/a2RUYW5pE4QR5Ax/s84rXFDrs3LUJw9ebd/+B63EhKCSoO8pGo21UA0k3vDE1Ms1/H
opSf4p/s9j2VxKp9DLjep0AommVB+p1SobWiUSSjinv3Ced5Q3MaoiqonkwAshRkIi8Wxzc+zaSz
Yr04DlF36/Swuu+cHPo9tZu4XUjjLvvfYDgb2uwgojjq+FlVlzRSmUDuL1Ph8F2kZaszlImGqc5P
FTyZ2eyhRXKJ3qXhJRw6UfYakMYgBkER/lNcXke+epE4MD04xzMTvvvsHw3Ovk/VIx1iSpanbT5t
aDEFL8aM0KliviG5Y/L3tjj69D55yjyhuyGNZ4/zNm3K3fiEhSvIosNogI7lnHZkCDblZXMKUHrE
lp68em2sR+4jRhpryPQcjkU8KOXs/52yqfXrZmSc4cLhliGRW8KYpzYxzqf2hZ1nStMFgI0q8+n/
wZ39hZ/qkp/ySZS2TlmRhjl95iPFshRkDwBV3FLycBCgy2N+qCUGZ8S4saIH8SCNoFmAD19vSwEl
Ub2HYz9s1ldVOd3/VNpEajnIioIKCpikn9PbpLVCopITzoecFWeeOwVj3CK9TrtTsYGjEHraMQW1
eUsDukX3Q+n5c5MqErvSqSE6nNGRVtx9VgndF9s1Q3fbXkGm+TN/kj9dpou5TDastxQJRPDnM+PI
DzbpIlGOhT3FclHNu7Z/9SiLhHqte3N1AK3K1LlypXenz49Zfy8yjcRcdR1pzwbbjhkSGeZTr/wH
cnl/bdFLLB09t6vEJobnd35POdu8QBEtHGJc3FOJTf1JM2ZO8xHSgeS7mX3NvYwz1CxqGZ3Y6cA6
N9qyA8ykftsZMcj+96tBatzz70q8wyiwH9WGmolBvgM6IOb018WGg1Qa3xGATiurjASRHFy/VmwT
iQEHavRqfIcRNWXQ1CPqSjmfz5Dr3RzHDWvjF5EFTTsUdF569kJFu9zdPQtbCVhQKoZHOs6pqb0u
cFtd8V/m6mfzICTbKGV/PNM+hR5mWs726J5JhK+/GdzZhRROrptP5Nc0oaFxPfLxQmKXL+V1j91c
IDBfUsodK1sCkbvcuiK6aRplycLiItAdmYPAHTIxYQwz1CDFpeseBfh/Zobel3M6rNmdN80/aq8C
uSdY2cq3yjhwRbH04FWa+HLqnHt7PJAnny63usRh5ODfzMKHNMfF5B/de2J1uvTfz1cb3FYloN+n
veYwjH6QhtCBATpktKHV8Gc6JjcNJIgQDU6Z9gikuFg9fXuGOF6IDT14VlxqMMhh0YTZRly5Yctt
9gwZwhQdoYLMHq01/hN63neCIS0uqmV1UrUDGFSetJsrp3TgY8pHtMgAx2XfD9Mzf/V8ZSbQHgO9
hVAhedf0C/RGn45CDWqwcZIDkT8JRhAh+y9Y7WntFW9Nsz140KC/QX/wuXqT96WN8D36Dkqgpd3n
g9iXcGWCf4RfYyh11K0CgQXY/Mi2QBijGzqGr8L6/Zlv5c5wkESU51OSvDGzV0eYETjhRmWE855Q
veZcdRXXTYpuVbHHaxNcIXU1nQcKqjiKO0KJB2I4LyDIteKbjkTVwh5QL7O7zwcjX6hgn3hqdt7o
pqF8Cc3Ldeq+ZDvz0YeaKsIcTHlcJCyA/RMBcsyDemCs+HNVfsa9ew+DOw8wNL6PPiTp4yJDY/7M
JaLBh/lg21dhGirnsr6JJmUpQppS9ZfTITuy/hzKcbgPol2QgbbafesiwO0K2kOwojGxXPvfWKFr
0xOs8/7SkvE2pR+xIo2e7FlbiLfWOcvV8KLEJ5olEc8LiM6sxEO58aYnEzxjo871mmLAgYgkGGNV
vXMGIB3SmOVs4/yOiT/ajozCQZpX7JMw5N2cs3c9PRladMpqN046qxC58XYZOzKGIgo+pBTQVtEH
zPRGvhAoHr92OtwoJlCOiIZ59/jhgZ53yHv3j8ylLcGi7rv9KVvpKSN6GGSNpbfOeBNwrhESU2Ay
a3H4axzaXIUBOxCeoVN4SeYhv+yni2k3umrow9iAYTOgtHp7v5VrFQ880kFTZTvGJm4IkJrNa0Wp
QWqRaM7rSPJi2xWaoqmqRqvJZhkZNVeKddPvKGnFI53MAua8rx7vBa/T+k0p/NBrNSEt2GzPF3GO
N3qYdKYl3yN6DD73aL0Yenw5gueumeYNrQBXECYmA0b5FEHlim/1qYdd7XXsPjKHS2BGmruvYvZ2
eSTQP0KPb4ok1u3mDD0LTH9V+Z3dBCuF6xlia1tM3iGjCnGWvIn/zzmyLtcnvkuOqQi9FuClGzYW
Y6ztVD5nyFgg1xv68ad1WdLZw4XxAtPvTaTguiO0bW1M0g6imQpcBWeQ/Wo0ocpb5otTJ6q05+HR
cmwpsNR8ZQMesfFiJpDlz7OAROy6af+uRfAf98cAHA8MIfxUXcfV5BReGg5pHI+HeHNhQcVBbjSr
tq4ZQ3cUjgq1xMSILPxHEE8KvIkC20C5sKAfwpJ/jySazAAQcpuy6/XdBynOvlFWMCKXwkpBzbYU
dhKoN+B8TzDuwKdWTOE2uld1rlCTSDXXXML2AB/S1f72z6050Kcp3UcnWejJ48lJ8PTmRoJicTAN
tUHVysV0iwxlXG0ddeYoMZzqq9xfLUGi2L7MHHz5Kriu6WPZsuJfoSi8Q/mcu8iu3AhlNHvutE3w
6jDmlxyew47zRjkvzfVupOY26G2drnGtxJqNuE40u0E1EFav9ZG6uLmnE6a5CzVx4jZNS1zQI56N
LaqohTT1+PFoyxugLPFvUPX14jIJSqAIR9pzXXUgHOZ3Vc2hkGvfJ9peoMc/gt+y+C69JgLKDgUM
WiwmTZd39plLZ3ZXnpapWVUZ3MG5rGqbCZm7AkElDGXCN3uigiIYbR9dVXL0woiyLX+LN1rw0qsI
dQHWfwtqSRgaCbRyu+wptJnT+4N8kQZFwpCzYvwiH3c/+5fkPhJEiy+Rod/oTzgXaa4ORtdHhRsn
7G6LeB6vV5sCBnjvBHlSiy6k7AQyqbOuhwzndy1LYySE3BsxNKGjXFw1w2AnMqb/NRGLiK2lWIZB
9I0dLqSO3F1HGupF9p0U5pMKgPxMApjegJ48KZ2NTa7Yv06d7TTby5BCtG3tEAy75E+wiHObm4Zq
9zn6ZEkUBhWgTXLvxaZEiVMr388ydVEmd2VY16RcioPPebIwlSGQLGtSzZFGvao054uJVGxiRygJ
AVVNLoa1vzU3F+HHvYroIo1FoCJKpvJgdpQaHIw+OxsdEAR82wV+y4+Dr9KRV5FJ9bfI0FCTcFgN
LchKux6xX5ccX4XKk47OGkAn6HOOaHKy+maBj1IJnqeX4YQXuYqqk2QIUylhwGkaej52UxZy98ot
F4USlgwmjLKbn7wcLF37EsseiZLyiCrrmsmJ64AdjTRuGFIr1BnJqmHzE6BlG5iKWQgltpGMB7Yc
EzoYNYC8CC8YJT6Qiq4WRPM9fcUSFIR2B/e+3Wu7bj1mK46+CRPqPQHzSHoV0RNNVb8WM9LRcwOx
YMdseHxw1YYS14JY4oWeHtVSkBcpLwakFOtQsOtbw+B34C8Hv1U5k2Uc573bigBeoZZbyfTsj9TV
ikTfQM6r5l0yucPkO0I5dXcV798zTeTGXjbwje6vihz0yYnMgA7Icf8gCmYbggGjlHTpcdq5UfSt
F15YPsWnHSIjc/rxxDjtInRkOWZfnnVbAzdF+7JzLG9hEyfSjsSxjr9bJJAdEC3iwPLO9/gwjd05
ZnG7MoOW1xnLGIe0YnpAwjjSxC/NczFguYQHNk3EQnftfDANOXYEOlgJ3denscQkVbtcG8PIbvBY
I0Y1X/RF4N9aynWuxtfRIdlZQNPThNW55jZNNpltP/Z6ITcwW7i/gtumGdnM2ui9sRkPdiPDoGRp
5FjW9s96xCfVQhGELtMz8OKPJKAJ4iWy5OSGtdw+35Q2Q3JZL1+whubz+2Tx00wWa36yutggo5r6
JskR0i0q8K3IEQvAQhGiUVgQREh/u0LzwYup+6qc05g3UOXk6p/K8tqZQ3owaaDthb2EMWGmxJvA
U7NjrA27i1ae+R+jgPUP/NFfcSrvVjwxndyruJdVTL2DvjSIlI8MOy/BO2pyWBUq+rchwwz3nLoq
rsIoMhENxr3Wd7UU3cBG2Dsuqx/zP2YgZ08/IPqxMlIMHEJwnsC2BFwf3R/VJJOOfFlxGPI1Wr/+
G39zKleYtxjWbuqCPXfiW2BU+iASlrWSfmljCP1j9mjgYc4ARssFvBXw7OpOcwLEuvuc5Q6QN5O+
ZRO/rK9tInrLZgHyhfR+KCPhUUKOjRHXOrSVEgKcL9PNVBThPo1JIATfA96eT9KShNgXGctrAr6e
N2dir6tjtyOgrtkPSIhDHq1hGuJUecuIIFgX1Kktz6cztgXvv2n1kuiShI2KvWY1mqihSIBElxRU
Yowa0XwXpZ1weLfa6LckCWqtC05Mt2TTXwzlYRIkqY1fIzQI5TPEU/kaPSEc8zCIxJ0aRKC4HXCv
53zrrrXtvrFqGEFYSoyWb+2RNxmqM2f2NR8fYfwhB5OL+vuugV4ZGLFizjWDiCa/JmHjIJhjp/94
/ExcDL9wE+A2LVDPxNnEtekTHwR+CnGB9iFjMFY5AOuGwrMW+qndvauAH/9aKZz+CSIKpTT+83ki
S73FcMEHQNHcuXQ7c5HVQu0BXN8x4k4cAUTv3e7mliS7nJwq0xaIvHJHgZG0tJkmeX/USsy4iInL
NAlWG0SHx9lBbImpz8AI0NTt+mXIzhbY5sSkQf/BfB1rT+6FbmNaK5LuBKdqZPnCymRrhe8Pkj+J
I2r89e4nu19juRK7nw29VPG7CGrELF41RUQ+NQtKR6cPM9Sxd+HJ12xliJIjAdMvFlh0tqGnmjkj
l6dj9HN5bY//DF789yw4OsDWid4rdnfzTY9rDRuYZzHlqv/SatW/ph4JwViiqu1g//71pyA6IhpL
oJ5iN1cYELRMwRwpgH/A6FTRRGFG09BwiuQeT7PbA90cnZCcwJu1SD4u/tn53e1Sehw7pQqG2eAJ
gcsK/JFO9S+yllAo50XKDQ9RvbI9+19jssPIVYatqpJqUOHzay3dxjn5TpQUD050PPVl1ARIilAd
6VT0g14QjEN8XFj6ISlYVP0IfM+2/rj9jwGjcNS/PmIBSqtKC5dpibAtHnK5Vh8l/MJhQ778Rxnv
eE3AOApATIiP50c5u8NA+7XbzuL2mAqwgv5yK1CXlXWN2Eph+5O4fcnnMw3wYszNPUVELmoVfvst
1CAnH3huPOqUm9eLgWfTF8u+Ix1qS/uzrMkihwTVd9P3NigGv7yatIkTUpcpg8sYmSlIv9gwK65B
nywoCDszQwRdXVJGcYjIBwaWSUw7RtRzuXCkQEk1wa99yhNB2sVpiHIjAcpW0QpLiM6q0/QxjUHe
HX9bS/Oyh08Yvdjq1N+qvipP7BxWJQMd5tONz1JdieUuhc0gPmA3VjPJwN6bImmqBmRpLHD796+S
fQeTwXBlprdky516RKP51HVdHZsYITPGt+bn0O1QoWKD0eGrg6qRLxddci4H6vTW8YCTu2kqeod7
AzPDyNI1sCykS9VV/97NG9fnvsbXiF70hdxhWLzr5PjvqXrU379reDsXOcbUTyrZissu96F3s6ch
mdo4D2tiPMyL2Wshq92lJ/3SQC6nSEE2jx/c/5RsfXRCyNKcFkajnwIReefOOAzuyiuLklrnKlB5
QQ+hMwJomr9BjiEZAMnPVKcwliNXwYz/sDRGP3sO1kJWanJ2JldVM3WNG468lmVqS73dKR6jVJaf
7gMGq7kPwP0WLhwRZUJFcKPsV081g+tWZFtynFZx2EfcMLr6n+A1V2av+2CCcvfPFO7YyvlU21Pq
LyxJ6x7hQxOmh9d74PEgR1q2SWpE6mSGr59Gbkdi0SUVTZofPUH8bS8d/yywoXiwDxlTDFeGBu58
Hhgwa9r5TazXBJrzkHFETTKTUrkkYUvbYtspho32p0BwMqKFzxtWHjn2zdvIGf8jcWyMdWrZM9Yk
+Gt9xE8B4ABbDYDA2MwvRjUsBEpQ3wh7PNFvF69ZBGXX6vPVmKe3HhMkaXYcaJ1wAGCstslw2/ud
bH4uys7ofuLBKmtqhL1Gmc8cmkXEZFuIRlAr2RcvQ3MWzvpGbOEFQDx09xLpjhWCFZ/iAy4P0B3E
KfIAs89sRGADdXHpurtVrAZOabTOeCdbLHIQ2I8pbxsW0MjxfrOpxKljflBnkekUZBlbAUf0Qx0d
AGVso4yD1sP2nJEDuAWJuoHc6FRStJzzisgY0LlX2hn6ZNNXkTZRWj3Z9zdBR9FDRkVxRr6V1vso
QbWStSwU1nSZFAnW7s/ZnKJE+sGnPWCC2PuEUQirNqTJvv4sADfYp4SvkYh3ZA3CgH5B2bIfPOol
SW+muT4I+pp0OW5RNOgEz8xgTWc3cX3U643VHPUlHUYUjDik13OQm8LQlpuVb0IC0qiBKsfyyFxe
FDad+eHCy4dTSqk+MveD8ZtcrTkzuWJt1LiTShZ9qd0QkP6OUYg7vm9DvZmn/eiQckOHHIriiasR
nYNqNf/B+Z1LH6Ml0dxtbJc5e2IJ53Nnk9sk6H611Ss0KYA14WODPGizeYgKQ8KmlrhQ6n4x8yIT
Zs6Sn7hqcHZ5U2adBDVl8vSOkPFH9hujdyOUSC+FCDhJMEppp6LIG3oOBXNH27mv9jS4shOVEXa0
roRpJt7GsLNUb0RL4RF/lKENyU4f2kuASPC5Xbm6ys9glX1DmPon4BCC+n6wFhqwBNFY3jEwzPCn
sbEfpW0L3iHC/mg72qqOom+XbR07E5qsIEucAH1WBzNgDo4kk8nRAFPdIOXibKUseW+gMm7gEpxE
bZOd+4LRIcDAfOx8svknk3Q74Gba4rW245FJWq9bph53JBasNeu8SXc9sTdSLlx4gjD0w0NqOGlb
Aui/HxGRetTnqHKMY0UbU3KGm+wHrMazUpdz9FRd1pKQd2+Pi6SBr+qFSwiuyp1qJ5m8Y+XVp1T9
q3lfUS3IF1LjBDDgAKDV15K/ypH4GqUAdHpx5/YXGMnijWkvMuj3uzKhRAG1PZG2VSseoVmWwaku
sVtG/Iy+Qs8Y3Q1BpU1+nNnke+kcNVM5s757rYeJ1MieeiKmtoDPNEq9W6pg2z+WO5JdSFXMODDW
VroVobY5M24U6Fw6uz5ldte/dnydWUMM7crfdoYO/x2WE3A2PfZvhiONVklm+eHkosBgwFhIQ+0U
mFx//V1vXKqSk41U0y6h/63xNP7CyT6YqIF0cGJf8NKakVYM5xIAwa34BEbs87z+Nq5eIm1MRFCq
wo77rDnieppOx9YfVtkIANtf2/sAZ9YNfoH2V2NqA0WUG/L+UNxAyOXUxboVhNrR1BVH80o9Mmvc
UFpeONOjJllbjOJds/v7zK+mC5dG0hKrXFPGdo9tZXZvqbVSWUtoCf3TVxNhcTXvd1GTQONXOnk8
zSPnGs66WSmKFkNRPdFUeo++VnDAqjRr2NPFDyh2RY9r6TzjXlKJkRCH49L98Twz1RzhkHwrWwUu
7hxJ7m8JSy4iZLqD8WHvdDZ37+H7rPHNbGhOzDUOl1NQ7R5lcuQbPnRFwQDGWD1nPo+XC79IJCI2
IeMpv5DZ3VvhPVQ5GCX7NE19F0RDFk7/794gKSaxGC1PTOaa2/nQ2x8oDfLnrkRof3KGFmUUBiy/
RRvS1Ove8lknhcPbc/vKqpsyVGOqSyBRwecjknpKQyGs7U9tnz6L39nXYTalxM7KBsNWIX/7XVWa
XBHMJb1puqZM+3aSlZEuNe+NtWg0SWZVINCD/E5pdKCxapmjRSAudWdqYDms4ZaKloZC6p9Gevkp
GexEeKX2FVSn88dHqTlg/GTTExg+eDHl6rJx8gOJSN30SEPPrXypZKMpAzXtvjDjGW/ZBzDrKCbf
A8N1r4uBAggUE4+Ua9xSZQrdmbtdLI5vK/zdtDRL4LylwHkQRz2gF3eEsjC1yPCW9uKndRZB2LFe
HM1gOj0BiZ1t5ec7a5h1XbPEwak3zre0lKC/fGh9ZjdiEcLKZnByBqMwxiC9fqCRWPMDsb7wYMQ1
/Q75MzfJmFH64DIOnzxSi1Oxkup7pJxNeET4yeTU3Bkqyc+SVDkA6MIKaks8tZhfoHgJ+1PSYH7F
WHz6FrXzoUnpOhGpBZoLL8v7xWbLmA7Kkr8/Wni1/vcg+FJZrRN6pXkUI60H27x+SuQlySQWizbi
uj4mQIZwSCgmcY9gRN05LV9lfn7WngiRZ6f2SueRp9i7EgMZRKfb02w+yMhdAHqiAlYUHrII2TN1
qdaMoEKuV8gxa7SMIquJhJo5Axygov0BPULvx9Jsuf3Ml2BuiLfREE+z+bCoiuDpnNj3uNqWhDAP
VgvXdECiaYFOjc7/tVxTP5feKEUCIfp9KZ652kx4z+aTfAmv+P+BfE9xQgU+lHaKWqa7yUFoOqbq
Cbdbfd2OdWsiD6Jp5IY/9kDo00QWvt5Mxd97vfsYfe8bSBrRUlMS/aYrVQPNZREtX3yuv79kcrTp
Q2Of28dbaPo6Gac464A5vZSSdHzc3HBu/Gf8F1AcJnlrvwoqweGMehStvRvRlHls3FGHSecKfSpL
+dNNn2wvpqLzr98mmtXth7sefr2Ia3r3AnHDU9wvAD4zVxAmIHaBcIyaNc3VcJvTZiHu2+z99siu
TojE5K00sk3AwSaYufVjHICZN2wwD/sY031IGFgkGAbueAFVGyIRyxVYKhm6ChPfpzQxwzXT4zjf
D0KLNBvtsmjvQrntGkLsCDnMVESYwU6etUXFGU4YDy0tyzXzKRJYn9Vok1ErVKnaa2V0A4n9+SR/
u9Esc8Dx9RKx7RdKYBlSGlcBna77ERiUV24Mb7ZEmocm53Om+hdvfAfStN9gQIok8HqsNIlvMLhW
5CaEt5J+qSn2noWHCEIPfaf1qVvRIU7N+tJzh9Btzj+HZOEgaehTftFHi6UacqJZdl5YaDlkJRpB
k8RX1uiCgIwpHIsALSCycQzQSVaXEA2jQDpbj2PXMQbgWpY/j7XtzTbTz4EmJbrT9Znd4lSSdMeo
vKnJyEtMNcqKrBMj/Un80wo58cIoa+GJ0TOj08GlWjRV3JFcGiEVlpGZeY6mKXskUnrjHRnMm25j
vFgil/Cq+zq5w94cOYR1k1HMdYgIVvBZMrt5hyUs7p6e9Jmn+vWFMXE1s17sx/4of7qaQkzJ93Zx
k/Kb6sRANMzFiQ1TtRY9yAPMOEmJvbshn9u3B0G9zPnE2NpPOsGJn3xevmXn+LdXilVv/JoB7ptY
nuOKU12OUMc5HqqLueH+SX/dsTK0oPg3VedFGkYW25nIy6i0yM9cRY/teyXKkwM9LOCZcq9KwDJc
3hTHr+4EV+BmJbGn5Vv2Peimmx0eA0cWKuDQFzK8t+USgetEn8GoEvIKZFgZLdgu2TcoEMZU+gGU
aPst0H4/kVYwrjuF3xyfucltnFNiwwwfUBuotxy6N0kgT52zXuxbGmREFm+5nz1blil8AlSS+WNh
3jrQFLNPlhIVWiNWlkywytFTObBgbj1cJna09uEjZMpYGu4KY6mbRwn+O1Qs/vHNp+EOKALzLsRi
sHHHmwj4eCEF3H3WL8T5jIy0FCEiF/EiiIR0i0L4etOoBwbFgrqvRZ/rorCoTxiYbrFVwPElW9G6
jZ4UyV3/N8mORHGj4MMczQg/MgRPHd6LhWLtfsHg7M485JS0yDtVhmCRgBucZWKU2XMMkH4CfJrR
45etjA6Juezvt6juLWnAs5TnG6/NdAahYqBbGWbXZrnkZA3qLNUTihkbhwzy48cqrdHlvGl/Nv8t
46j+iVdL6ynQItbBFFAEczDkE2nU4m+pK6zue45pg0in/+yhgaDEWjz3uQjin84XnvPdmTedL8CE
BhpfLnxhG+JJeoLoVPh77Km14bonyYohwmfrbpBJxSEOQxPr50gLiLp4SsA4ne+BpwHMjWy7xHuY
s3PJyni9bYcBPBNAhR/niBMBalQ+FLcBK49eNt7CVOe6jn+y7Qust5KjTky6SBt2YipLvgsIPI3t
HNo9RjXgDy4HN9lim9bto6GoKXUdMyQPEC27avwRZt2qpkoxjucebz503xeJTXJCLm936qVsX4P9
SBhyti47Cp6QR6ZcHaUApUksE8GBm2d/otyktn6zlnUH+0qPQ/LejFIVewZdr04wdS+Jizt2cwX4
Bz6O2lE9BXQr0E2akdexzgTjwojC7BDNbFs3hHiluQuWwMlvvrLd+ANecN4p4lVNFtUa+jWrL95s
puABrclPKpRd1TVKR/7jWO9ukD+euPqWXV7TBhVZlHdhuIFNpQWbPeiJrrf+K1oNjeFIk0uekOxt
sVv5o/JndWHq/g/XQAIGMWNwjktcyt49z2qptQ8wiveFOHdMwwQ3XqVPRj6Rp9n55VY1djHazOhh
b0l4PSeNdPRNCPbHMGNrtU6RqJP94L99qDWhzFrWswIqW/ee0LiUUnehBuzw9J8McIUGkSJLmdvz
W9Qqg2DSCEwqYpfd0TCriH3ROn9l3b4D+1jWH+xIN8WD0R7Xgcuz2fWhZa9VYVcYQzF/1w8jO/IX
12UvlKr//B5hoDNRe2Ip3wJGAy6lagx9LK3qDKjlneCCJUAkFXZ1fCsYl0Ce01orOPHDLxS9WJlX
p2qhyhwpWkf1Zilf+Lk4OOWCjk1a1Y0j4RaeGdg3OrrMTupNDrJWhMYBGCMR30YIdCZIZILJK17y
3jbO5+48U6Jkpc5vxf8UDbHc20kd16BD4i0SPjuLR19En9sl6ygUy2vH3dn/663BMPnI++gOMELl
GhG2WvJJhNYn0KgVi1zBND07bAbZ9sAVHXQFB76xyqArkHQGdqoSwjDVxKkvPnwL9QDvp/xjX6/u
LAfBOG2n/Ugw05sRCub1UuJcWpJy6ks+jtccRiOwY+I18zt40IV9iV3+F72hG/MQwyQBERHqaZTD
CWjqP+5lgh/LDVQ3qpmThSAUchespgnYqeoxmmUl26PP6GFfuAN+lth8YVr4VST6PjdifB5Y3paO
u8WduCwztIntkr+Ms7Hqwng5tHJ317DeU/5VMMK/2yk5i+qgp0G7f7Ac8QYDlOqVBOvSFXfxDbmq
XrdftWsUydJM7BJvMvcMUqhP/pvbG6kOflyOwCfmK2cj/UqE//K8RqAug4VwhLnqvbok2QRX+Vb3
hlPM1fVpkttOwZqGRx67kJXyKeTRzrRN5m1coj5604jlKYBdhshrFwnHn00TGW0UbuxpjB35ShIp
baNJhhV3IkXB/VL/qelkjlbh6Xny6ltTUZGM7dhBkD+dhFarEwY4Yb5J0DKMh4txKLFBQgpKM1rt
AH4KVS0SKTGMm9eTqDgdNIPgtaUUvg/yVTUccEXgSuyU5o1Qb+l1f+LXHzJHAJAJDqRxW/Ak1tDW
Bh6JhbfMtvBEwQ5FbLQgE74M6deNcSl6Y5pf2YflrgQTI54UpVTen1Is7hiLrOcjTKUmhOJrXVhd
wfkInmJ9LGR31z4AoSzJ0K/ybciSGnDFq9yhzFO/JGNzcDuX5J+ea2t5j1Z3Lce6/BF1V8JqB6R8
mlBk1JKg7yu5kE44m5hOvTFxuo/c+tsYB42yBDU1SFVo0EZQjlyr0gP5GA8QxckssE7dYIWTOyit
Zn/Xg8/G4XlVpsxod7+BOwOjn7esta7I4Ab3FlTLI/KvCMFxQmwtWv9jyt8koj1Owo/BlVDeUfr+
aCfdVhhfQhCreUytqfF9hFNN1Jk5/Bty/q3VulbXnFI96nsDvxUDt63dM+6pt7ExW4XThC3/pX8W
eXG4l7vKaFdz6cHDLxt8yevk7mDynvlvqPyKL0zSV4PGhYislVSmUlcEGs0igV5IlR9L9wyA4L3+
A/AECLMhigpxJbepyRMuRApCevfXlNOFfmj1OfExbcZWEQtLrihyKsZD36kz4l6VgJOk16X1t9dJ
dWnt9qbnxXukNqhaA6o05/bipDEzaSXvOpueX5DuEh3pntJfeI1VH6NThi1kNlk4ggxhGkusFxNE
BBaRBpnO487jotn9tRo5XIZsjBhw8TOxQmNgq52s5A2Z4oxMmzAgMZfweAM/WiAFXyLrTJRTyLDX
vQf4Db5sYJheBGqU04XM+fv2tT6xIntod6eDnMcI+BloJGjLqFpTyf499IuZXcE+izN6AAGdrhEd
nbkTfq31wSEc++E5IydUtNtXxnSWhQVp4vQTXCQRlC6hryVAGH3FRRV8fShR2WSomU2PkVDks0VH
lTE+dlxhzLmf3Kb9V0g5prJDLDCXLnbJBfTW50nwQdIjycJkYhAUHeYH7cArU7gMtqrPYZg3T2q1
8KYhgywELrv4ewwkS1dudH27Iief/PDjiiq6YxUs6axdxoRQT3YMTSPGn+2PC4wq1IdB6PLPgHNY
AYQHCPVUNysKC+6zGmLlqHskeQgwuSqSHXLwSJMRUDM8xdcxplt3mOZFIOFjA87v1TYPVzCSiM41
TAZ062gVVVEYHV4jE2BnibgPHK8TxKrpkSyLTT/g+oVLVVLxVCfqcY0oIMQblhOdlwNg1wDkTL9v
LSjrKClOOLa3g3XB1NIBS4HY4Z5sIeg27iGjSS02O3eea8mf8T1EjlPF532zSXS2FNnWjfk07L5u
FD2LpZXGqsx2hXUej9TtTWtlT0vzCqTP9O9mLie/zqLPIYMblp6v5J2YPxqnWn0Kc6EkyJKDtcwN
PHghveXSHfej+V9YfI+EupZEMGmlRRKdY/Lw3EqTKrfoGf2QKxxWo22L4Wz2G/TbesKQkTSmXMEy
O9h4Mwfce9f57evxbu6FRimIFuZhDr5IBh2m0/z2ZbWV9ix+5CHUkOwfbLYsPCIFvsrqasgQeEpc
gsnZ72oYjev3g3B71osOI0XcDhwZSfo0LsULvr+zZuF9llFhj0nlJj1Hfx3aCNx+z7NvZHCKC7hw
9QR4lhjB8xRO5y0yOzd2KhIVuozI5pmFVIkBDi64EFGuyoKdQsPcx5aH3PomWw4qjFT+P7AsJh3l
She272zhI46gH5kYkYwsEHrUvDW+arrpcCwdg/l9H71TvYPcebGX9z/4UnbUgwl3FsBTs/D4r7zN
gUS1Hf8dRNsglccWM8EQHlkR9uQZaW+b9TZHDx5/r/GAFBfjG+eoyz90XmzR72FlB0zh+scM3TKd
azQGdSr4ViGiJ4CieoaODXmNGmbzAy86MmMyNQHFRyC+ulOHwNH7qHgFECrD0HIyybQU3kVr5p+j
ToCdwlFl9ntAJqv0LtPr+uO4EEYUVM9+Zqbx6hG0wAB5OhrCGoPW02u1uF9p8x6W9H3uGi28W8Yu
4y7qpDShAMX3E3/JzfJMxFs4KYx7G7UpN6GU2nyTT3fO5gZTHRcnjgDdDjNzvJhS8sbUSyMM6dcb
Wr+EC0LwMKsfMsp/1SI6TsztoLqWbfBei2IfOoDw4Xhmzc61pahT9nLoo5fvNk4ZWwnB4CqJyi7q
0NUbpvxmE6v0mKWW3jto2wnMe0y3iV4sSHtBxt1/EsC/A7Yj6/8gWpUVtmgb+51xh/YiCE1d39jp
lDWhUaZNd1e6ZyuR2tBsEv21bMIouRTXvdQ/1doClUrobaWew2UUi2SerIfcO9OHr913fjANE+DV
opZzyTAr8wKAZRjSxoJpjxSQYEUyFyHi+GDynlqC+qID6BpZ7XRyIWDZ1pGs+uZKnsHnqfV7IlGk
g9Z65qqo8uNT8gKdeLciVR1dzdpg1zlF2lbgq0KxToklOP+13Tfdy7WgUlJ8r/xKL2By/pSkn0Fp
TQ13LytPFpQ5F0a9XjyJDRy7LYvTXFshEzE5H5m58LVATIN6an6Xaz8GFzFkL15hzixb386tL02I
ZL0aDHdUkM92WRwV43SCJvGOvfg4Ht5zDtp45+XSKTTSjjHqZNzJS5VVj52iPt8UtHU8iUlACFrW
5xwULE0b+zFiEIuY52MjLw1EYRTeNv/tRObElHgQU/pWQN5QXPG8y4Mg5jpvc1wx322DD+iTaDJt
ozRsOGzgtvraLH35i2LLQ1Hq4ASneObVbc9GDOT7U3MpaZPpUQBSp2YQecQ4I96+hKcIpLf14JXo
ImIwaUL7NBawxK3M1yjJUk/NcEY2DR4TPSWMh75Q5u349VLEn7XLuPsImT9xlpi+bIJbG/Pf6Ajj
fwNrCnV/qUiJyoeCGdzhmp3WkEP2J4b5xkXJKTNTiUj77vdVgG0EqcMZjmR1Y+rAmg8Bwm0ov7jF
bsKdwOWMIIEbBjSnrqi7xp9mRdxGWTDY4gCZQa7aszSy8YsAUmD1X8BwLmOAPjIwOBaX2+CuSWJY
gB8ZgnOpy1Wl0lsVJtlYnrgfQKk75m+jzOi1Pi3J+XqE2x5P3dcu1PMP+aUY61F1WpIFCpmsCwvs
8U5IZ7ioFxhWmwlsGOZ9oq5sdlhwLcX1YBiFa9kXp1oW8Sq+VPjaaQTHoSyy1IeR2cVeNtu7H/1V
Xbpj8pGGqTARbdm9+dx/fuX38FEEfBF9TTuDmo+tEQfn67J4qSYzLm7IywAy7Wme/RnWCwvGYdt7
wjy21CajMOnzW8aAIIHNuqqRVNX2pjntHUuvkRf0lX25EcXfx77+uX2F/0qfKrVECko3Oc/Cc+2k
SB3knhU0a3eW2FB+2Fo97zb8q3BdpVY/ak+URi0iedXqkJ6SoRbdGwXlkqoe8g5DBXfr9N6+UAHH
FZvpFcq+kNEu4wRkDP1EuVQhYOYlVoiilodpvFZR0FrDBvOo/iy93XmyqLAGdz7sX3ruh51vEify
Ry0woJ7aucKYVoKIuVu5sLJG/2ik90O5TXfETB/MdvyoRNtKRJL7Y3P9tLcgV01T4a0X51HoKKVJ
DR5nYh1QhQI7u6u2hNSZhhfUW9ksPxf8rVMkx8g2fxH67WSXW+u7sy+cAYxFX2gZnvQ3OzHJ27bR
Qd3HZfI5Ck3+0zVIofFecZJIbGpZ8LG+Bc4Zy/VS/kQZ6HXFwyHw+AupUjjTsqdsJpe8lf5Sk1WD
mNkbu+NlpuDat84p9c+ythix0qkVObLd3tk5xLaVC2Ez9R7VSQCkH55BcjyOERVd/fV4YmJrH7Jt
ZWhxES7RMXquKlFq9TYfHfT4vQZorLdk1gEjaKEf/1zdWcKc/l6Gm3TAQDTe2PAOGyoW2CBUrTt3
7SzGHu1GGeIp/xGyNUmpE+HycXWOmyffWKySCaIH+eOK9IWxmIhm3dVZdRwcUtTqHtOvOaUJJsvj
cTfNkTy3/wEoh3/0ZurnRgHESEYBqC4jw9iBnBb4i3MnZngPrcxTXGdTAYCFVTQp4h4tQ0KK4GLi
RbiVCsj9y5TU9GOIR597H7xk/cGrROjuua6y3qgOsf7hy74HiB7PP/7tkBsT3wmvolCTs639O9/p
NMNUb7/oZVhugbtV/OzAN7V45oVlHp4oi90StgUqmaUXTMXyw7GhKQaI5iRd2+FHVHYlnAnFufft
k96qRp4c66CBQnzBy2fe/KGD63epslIf4iJg5Cfv/nRA4S+A1DUmxtkmTO9LVFPpzVO2AB+hkfnf
lYWa1BbmCsn51jOTRwP3qIFmF3aM/vII1SSDbkrCLTjEVCID50Tdd7xSQstdV4WD9XFpg0qA3l8N
c6+LNlmj1nv3KVzpkOMViYLmrkoN0lAqNM+/UFfoYT+85B8gVA55XxsPVwK+go9192LLuFQW9nLl
kzFiyU3emMIVLr7uI9zIHj2WZDslA5H00Al32FLtrxt0G0IUoernxFmxFZXc52QiW1ddBs/QcFgw
WNdVu96FyDc6IwHh6ycT18nFdq9ru1kP0qTVGmNX0cyy0nZHwLTs3+09+UzM1L8TavzDC3dJI+KV
IO0saMuLrhgMXP2qM9y7i4qp9VbV/vExzKTlevyHhlRo3EeeOGBpHgRKdPlBBf3p8GRvtyVsOjhh
/g0AskDdt1jb7ZT9apelxWK5xw5g5zmsr8WVrjvc1/A2Oss5bCvZ8Ur5yq373rnpI/leFDF4Eey1
2+s04FPzWxUe8VYhajlBV+rXxZq143wpb4Y6WcvmAMfeu3a+Nd62aeyPePeo4I5AWoCY9FpzVk4P
ZAwxX1jC53/23Mxs24qgwsy6d3HpC7lkQqOFmFtOkV4sx0ylt5B6kizqan011fkf2v1jCliEVHjs
giGE84wfuuMw2IAb3fKwsPvd3iLhJmJrWpWyTmOWBRJUMU09ekQ3+ThNP8DdMbhDF5O/ZqSeupy3
/e2sqydB1DFujAZAhMsu+4KpXwIieVo1sDUgoIWGU1M/xbUCOp6+HmkCC4zEqlbKADp8v7c8azFj
aAs6v3hjy+vFUYu4apBILetBi3rqmL8zRUpanYgDFDZw8YBlRQ8dHfihUEUg2PkMh5hC36+aolr2
1rKvuikP27gvEjVBP72HvDhI3svf2hm2/f2pU9bdWpX5V4vNDSkyojPyPUaU5sGoQF8Rwg8CWsWn
r6vHPXEwv6oTbucMFCmtqwPlrsu/81ZwW6j42GHq2sYXRUoTzGr7bAfNoDrzzB5Q6uCN+mcL6USq
Zs72svIGdBk4ZNDToaufzOI1f+09NaEpqKW84G2TvZL00riDBANzXFp9/W3a1xSyy8aeL94O7LlW
3N+6p+9JhEC34oajDlkX32Lo1dGZ5ckcaYDjjlnMiWJT/hn51+BGMzMj1xBzejO+toF/rhlSIbmj
O1xWwBeiOEAcbxeS1EW9MV3VJNO73hYAp5UB7OZtGKLRNDE9hHg5o1yWlE1popr08qi1fvLsx93M
lZ+0I/im9OLKMBMYNbB//cLvYe4dcrZ0/6JmVeHBYfVGdGpA9fO+YE7+iqVnadfJdQyIe3gR+Yuo
skFl8MYXlpSJVbzrxYJqUSYPI3W9ecad8OmeHJag9xm3UCjtpw4hM9C4KmQWlxwHPazuUOPzuigp
R6FdELpAPJc/WLH4gKc6l2r/DsF9LjOuz35rLJ9KL+Rv9HFAF+wRWAha9lo48zRVYwjmrySpg22K
cmVcuhHNCZnS7q2dcT2wrPMAIznnK9/fgLYDFIb46baOFtUTaa7tuESffghrHMw/mDTTaHA9miCM
Kn9URBRJRzhKssccZDqMDbuh58vtyPKHOLY0NHrPOGVHGNzLOLGpY4ziTucK6/omwMUVMsmT8V3c
wGaQjWu85PjdjAR7PCLdFDyP/MYK8nNzncjMdM1WOdAH6zZ6nX/77fzO2s/hM6dCqj5/NDqwipoZ
FxZWDQNyFcl8mm00Zbr4AH4jy2wSwyeTS+F+BcbyWfw6YtpqojE1d4nt4Qu8ciP5zEIPveFrCqH2
ngdruPhePxOe+6dBh0BjcxH5ZP9tIIbMVT7anjj+QyY8Xo6P6SV/v3Y3NO4BHXZ+XdPup59b5wlg
WkPBKcGm7X1ueNy+xX71JcruJIAynpEqgEqOwn/zvrQaGJhqB+6JcxYNDBgAULn41qxGugSbnUs7
EyHcNgDk07SUREb91x/U9v1EbpW/gAlwDFkpo3jilfCup/lKGYj2YhvkRFeM6al/nD0q0aluDuxb
pCjq9kL5lcZ1H72eeVL+wZrBhCMFRyvJdGP0miQqoruVA9e+BFvI0jkyL590Nm3GLOWnsaOAlxJ7
MYWLNU+QJtHQ/KwrwyPH5mA9nv2kuJdZhBaRj54lvMEhp/KztXHDr914Uq/dvaGT+9zkG32ndEFj
ti2fjf8ihGx/MWGYEFPon70WkNnl0CGXZ14GO9vYn+WHaa5QqFf4NeQ4SmCo83Ab7v3DqFVMB6qe
S4qX7dKgK4ygNAO1bFOAMo9fLdEyihkiyyaLWNiPi92KlVcSERoUUO061J03QPm4MElSDIArghYC
+3iK1trwms5TAC6hhXLWVeplBrY1EK/LoUynKSZ+VyLQRHUbFLadUebchh2u5gdbYHEfmO2+EkmN
6MwN0cWs7sdn+1qZMMNpeL3LqFHerqFS6OVS2IUxLxf5QP0gs7ZX0moX5C8pFY+/kF06kFvinI1O
z8EJkKXFh5XiQotXM7UCsLyK4mq/+75ChFBRl0rDJ+/Err7njSrdwH32LPNrTmbStKleUepxCVV6
pdjyVh+ZLeuicX8OJAG9fTYuSwU+xjZVQAZv11piRbOLtbZwZD5hTfsmtkJ3fhGszDCEaSylBEuO
2fRAtUlpxkPiF8YdOcm2mq+UgXEBVHDGzorAWSt7mt6qfbnP026M4ZjkompYLLf1WVekPhnmeB9x
i/QLpdUEBdaTRK4rSNTHjS4aDygOknWGtXAdfWaW1UoWfMgDFgvkhwAMp355XC5d6ddPcEioyKzE
HDj8sMjBABEyc4weoTXzUjzNtUvIO0u5Wfl/XX8cT40VxNzxW5eeIjj7+1wmakRP8ZpZobTJBPqt
ZqIwq4rE9vyoE7wSdfvyYKF2rjzMZaweJiV+N/+gOS8yzGIjDKxw7sAqSy2S97Px6CqqtV+NnAej
8gak01uc+dT0Mjk62RU7UrPmzv+apFcawVo/xTRvUSVphONFbLUKzHcaiVNK8GQaPhCO2uFebDB9
GCvKVil7cbB/9hTnoANWOV+1iVRv2QpMTnAGtvCBjvcXiZDHSiBiRMIrdsSCYXFNn+QDA9aaSQRA
uqBo/sd/k6/QzeV89q6ynfd8sX12+eVl52E21Ek9SRts3sgr3mDWfakRljcMtAxII/3rKUZocp/G
t9u4v28M/0i7PKm0clI2PRQvWnt4+NhrhvwdqSM2A3s8lSC2AC63GmToiOIR82kclMTFqDqFt+O+
Cz4UjM7TuJjsqxuzvmNwNOf576DRkqM8XsBYMoSz0EbD2OSfeVQ3BhzCjf/JnlkgyUJtPJjqJnze
2vGc3JYNbrwIZ0/GacFA0R+zs8PdMVXDsEB+MSpIRFbY/aRBMjKB45FMR16mcmZQsOROsQE99RSS
hYDM+UjnrRYj+ukfwnh2LG817wciQ+qlyBBfTc5OQfGFH581EPEbovs/bj957rpyZOgn87+EnZnJ
90fw4n7fmEa8ueaJDNg/aaJBhwT6wzVXT/om2I9GBkOkRO8U4a6Zhh7ntU1hoTzLt//bRf4WsQyO
3fj0J+IiOBfZA7496aIJs/MQhsW/dGk9MB62Z+c3PqoI2zAQ5a+s7GlU1EquNAm7+9qfYmC96DoK
vPrQND//ZMw43Hsb49nIoPwshU2rKCciFmFEMK9gZzXSBFbsk/ZC6+p1mfVM+XpSs84erFurq2yU
LUX7h5djYj1Tkpzg6rReLQViR+FhYRcCRB4cs4l+yTRcwGIR5x6tYVRvd4Q0HCxzSWRByKGg9WZU
7az6ArWgOcCDNT6UJF7RSSU4DurJ/SU2zi92twgztX/kROO3/hhYiNY9gX7rz0CKI/gDbdNbz2yG
oPtYTTTx9yI5O2NVvFo0FnXOkIkANe4/67sj67TRYUR/Sy+GMF2AKSTQ3wqjqwxhVUQgK/uELato
U8YXCChSVLqBCcc3t/y6DLyCb3yuuNswaccy2GoYqVXH/O0yR5pDqC+vRrda9FY1oBqEdvfmOKrG
1oPXne5q9p9TdRaQqzu8oYHBKxRfFmEjRmWS1TUyNGlkH4twdLJmq07CWN/UhsqsmIq/x04pjWXb
SYeThe8w/2vHC28d8wS0NCxdczGTFunF9lv4QORmoC8Mo2lh9955WB2xcYSohkKyO+jYVi4nw0TX
sbKAvGXcoMjRuf9rX3QmeqTFc4csYa+yA1CA4G34vOmXgH8/K1I/hihfIUoZF/0LkOnOblE3n0AY
UwT/Q+ppUGvTw3SLJh9W47IhR/nw9nPQy1X56YBCyTMO+++s5BiOaYBHIg17YF/t28sPvI/PMMaH
y4oDfuXb0HfKtgfcKQvuVW/cllTuuOKQqHWGmFJXe5wAcMCn1fZu9pZXmN2PkfgV3cQtvDpaOmcE
nvhn0PdzNHygWx4/bpXseGgvXyPQ0tcve5lXD4tIzLskJGvqbLyJGN5+IA2eedXD2YdMlEA/UFwY
E7C9Q0S3td7l93x8qlr/Wn3kIEGAz01jrtOLrs4Kjg+GXFieskrXkloVeY2+Lo/5PsFuM4U0UfYB
rz73SGpk8fdG1m5yiy7cJSL7St/TewfY2MPWv7N+Pw+COFm7r3XlA66ricO+3bfhawD3UFEsuBam
bmBQ0EiwrVO9Vl+feZVaWsdL8qUGNTtCS5nnVoXK5v2P/LFhgIggOzAJ1okKRbL3COi9gQTXD7Ql
BKIg4BTiP0vEnpmTwZcOeWp8RhTL4vkw5x6Ls7u885Jnjz8CtRiozlEEn3nowT/NEqxYC1fMGkN0
wPp5kqypkBe4y809X+m9R/9kePnchvCw0/EYqkXDyoD9XmU4tvMK5pvPXFwSFEeC+KDd9XeUa3xY
FNbF5zsf2DZp3XoW6GEAwP/yupF8Ok4TR+gCU2tYiV7wvWkbvBY6QVh/PH6wDu/XBMYcdOCQ9KQY
3+e0ORG2KS1w009s0LlEoQ6SNvmswdX2rfaMO36ZCNU70bBKZ9Q60beEKcYWCO5McsmE0WNfhj0z
T7LTXIa57TcTB6yGzbt8cPPKGpoy8jV2f039qzwZaT9P40ixR1spgpHjy6W9p7aWQaDG68JjDbXs
Og3BBfimUrYDhOS/hGp0uQoK6MWRltZsT3t4N86e3wYNONWLskuNj8urdVVJcc4qFbygjK+J35vr
0zUbvt3p2K2PQ70lOUz/Zb+b6QEym0m+qdwEHMpDao02SKqDWohZX1nao1b7xM4L0pC68sF/YUPK
54NtzlulY1BtRW50dKSiDQ1OfOdGczkz2TecHVhgmZnhFSSOuxS3eFMKVT5q4XXLNFCeJqiKpPVk
N6BZIHyuLktpwI6Ao4RYr4zE5AWm1xfM8BJd06gB7fDbV+4yN92U3xtjRWEeJMWnwlk/BEOgmndH
luVmFBDp2VWwyOFM+qBb5EqdhkqhNbdiqi81ZA64CaAtSFU40nev7uWiHE2JrQC1brPZwpwLasgO
xShnAuGv/i4hhcc5UPRcpkaVOls4sgrGj5CTSCeSB+IR2wkETxt6Vd8ecTy19itngIzmeqS+E5aj
AiyK6hZsje2eSr2/KhRlkWPt10delwBQ0NvjQzxoqzoazixkFR9UO9CbFNAttF/0IXRbw/TvzAsV
ygBFwFVrzWDjL2qDulr0+iSpwYmp459n7xrmg8o1F6tnVUGxQxnkG1H2pFW9S0yM4vnWb90Go5Mo
TWKyltE27mAuNCKrk4NfbuM0YFJ/5YrYphMoHc9UJabqQ4e/Tkz3KDP9JJBBav+oizi38YEbYUs6
nHfS2ofs9oNuJf73cnJ26DU/DHLNApxjQPaGdiOpVi5B9D5h9tPBpJcfPdCv+RWdyJ4HGfnWPn6t
PHb1Ge1ye+7MFZ4SH33VDYSOcCzA/8nNWAChy6IaDdyju3a9cQcp8gOQkVl4ho0cDQl6azMp8pAY
im+5ba7RafMf2mxkaiqE2KMcoPJ2yntD8xHlLibXkvuYOOaero7HWkvFuW/Lq8O5v9LTF42Lefly
9x9ujjBcY44utIOXjZJuv2NUG4gHqbJ/1n0R/KN3SUJBhE2Xs3PPP8ccnqypCzaWky4WI0Le242T
fFtWM3v7IOyvkeam3n+DPc0xCCnpJCSx3wEhM3g3KX3zT5S/m5gobJprb2AdcRsUzlGuXoihMf3a
N5fK+VcqnD1qULCymBgE/T1e/h3BLnNc+OZhm6M4Vm5zrpF1Ls0vzbJXOt3Qs9J1xdnkxfFLWbDi
8OSpT2ok1b1h+FAJ6tJ/K1+qJcbBg6Fh8kjVH10FryLSyXviClGUkH68AJYNaUQdn/vgeiqlbt2X
UJZspyWreRAaU0LiZFvMfcQM2wBGF4vWulRevd+DNWgefd5toHXgKx2yBL4K9ObR8V7x+vedme85
FgDvkxgwts5IavIuYK6J0Qy1+RDNi5uKVs7ZrjAF/tKXJ2QMm7Stg9nrM+k+ZrVZK63I0kadTFs2
xiiVzqJ9jTXWatVjV6huF2OLQbWh1PF8hjZ+tAsYIvFFcGv80AlBpvQSvnj+z5+I12ulWKmEO07Z
XFpazND0AzLuobkS7WA0/ha8k1JfCilZj4pKDJFd+N10yduhcyavBjCzQgrMcgkUMVa6KSIoMeU0
uWQP/UavItB3Tvor10UmMNEmL0ACPmh65iUbi+jnjQFoyH2rV2IoiDnqBtp6zZpS7o07PGi/H0Cz
eWu9CUbzGU57YdyMcYI6v9Z+5RfMgWLd1ho80BQAiN+WhqsqFF6NG/A7gyl6CGbF+cTjGhXxca+j
VdLA+VSSGpqRTA9u2gg5lKOnnYLTLmFWwU2UpgA6S/CyrE5pyxLxudhzqs5YoZ+pF6xmpZ0bbL2H
TPBprfyQkjqcQuiygIB7nrfPb/dwqLH1J4oHV2E9X5AxB5Y+YhhPMWFIfoXrH/DtHcJX6QRYMekm
F9xceXmWz+v1RdSvgvf7NnwKphEDK0NCulaIjiL9cV8Vu4b8fxQRapAVrBD3tDkqIDgBQ8C2I2GR
rqcJVvDlq8aXL/00OfgdNGSFNl+aH9J64utZYFtlXVPtz1ojwGjetVrZzvCfu9WjcTnOKFHfD9ax
WOH4pKgTeHzvKwW3VlTwomBrnlHK1I6/H5iUqHp8XCWxzBH0sGbuIE07OaLfzfSdw9S6Rxqjqhk3
+S0zWlFjAEOZwUlyIYnxW2oSxpBnKLPgv0xNlG+/0puOw3MtxIEy9fMaBm9t9WNYa8zzKZDUA3x1
l3bDW3lPVRZfR6sUR3pAVxpLy/OejJmTLuC4Zab6oF01/x0He7PhcDXrvsJVkzhNFLYoJ0dJONuI
crJ4bWQ2bBlzz52SD9hEdyFV/C07fVnCCO/LcmsKSLAlK5xpWY6YLl6dFnyJ8sVl1QOagzJJ+Tbc
nTejfW6QLMwMzi/A0HFzY3DPKMFVd5ovsDA/HM9lUFYJNQQKfRPKYWKUl33vSuxZ6ooQDo7v0GTf
N6c5X+O14s5tf2QVfrQY8D0GhpFlfqGbHJSy2uV5FCcn7PUaJzE1rRLGYeUXUdEbx+Wobyg2UfOL
IbIOSd2Z3eOVcmRVng34pErlmxKXsAd6qkhkJRZqANi9yyjeqmXdHptEG1rZjodnRhAymGFP4ggC
EBplgBNwQxQgfrOtKAi774CRGyu+L3whh4feKV57S/8rz7h3rANSEBn3Ev/qVea5/vq2NNumCdtl
7U+JasWZU8+t3MOABlUZTJbU8ex5YoxwqlhP7MSSWO+l6wyBHMsic/ROS2dMGFCIb/vSSTJZQQN+
uGwWQXZ6AUpfEyopK7C/keBoABMp2ZJGvRgTm7I31XFf4a4Zjw3TiuKT52/lfIKa94oEvrTrwlOo
lRXGKiOe0tyBy7t0peQEBMr2ZavpvL6YCxv5aR7rK+OyKxie9/jHjzoPdxDbHKrB1kbI/JEMHZ8B
tqSWxZx8k1F5Lb9yszafvq47o7WHas5E+bY/yBSBlc93N0KJ5yCQV0C08AB5/0GX0pbWiIJGcw0K
zRKAnYKuxf8h0aGyveg9m1CGIlVDUYP5m3zXMqXDhIGX2X0W+gIfnVhDLNMqRZ1GewSNrT32Jr4+
s3D3cW0iRWM8DJ+LAteKd/J4CXVmRZ9PZDk64FNQ/tFb7VieN7Iwmw23LKOKXZd9rD/Dn2EdqslF
1XDtAio9y3zp5FUoepTrpUpHdmaauhBdmV90oBS/8kl6vBwI7RMWuhndvozKt+QcVbQ7O3iK+r76
Gs5q1kkKgx12DltBKp4k774NCuuVCFEf8Qw02ieSnAKjLXr7ttgZurELk6jyxPIf548/GPtJMtez
VDQa31mG+ZC/q+7eODIIfRk7ntokpKdk/AWKGs8tc5kYoMDy2fqvjqddRl+iN8eEILejv3zXesif
xXWzlajjhUNt59n2vH8PVP/Q+tfq7CE/5FF3oCpF1HKZviDC+Ze7QwP8NxX/xCCQbH8zffBCSJjj
btc+oH7sHtGfR95KTPb918jeLxGFln75P3EUaoQwCCMCq6HBCo68g45FYrwObfYHx3T4chCiguO8
N0atr5Xg5g/5H98fyZRW4G42C1sx/vSGcdoq6Rbuxz60xsXgqXa8SX+llOOt7Sq5VAealreQHUDU
wxbLLJBA4tl9avEyS1Pc5nQ10rDUVUPOiM/y1uIUlzniDTfp4gKENtLV6+McbUfPmYWxkfMD0XKs
ExxZgCXqJSMx8IP+uHTR5SDjJED5HtEEGQP5i9eOBcCAU+A7sHFYhEcqKlwuAFqXu5VH0AJp1O80
lvPZqUNSITl0xNW+Civlp7yhHUQsKZFwIt1xEY3uIaolmV/VtvU+EXbVuYVhx3XKfeUkwEi9AcRT
GHwOw4qwM37room9k7LWqCse2OQeT+OHhXPEMDqsmTyTM80X0wtK9fRtTyb3VdF9F5JBKIU2YOW5
n2Ft2XR2megCHSK71HQAOVkGG44tVnLBt9ke9ZH0kph37Nh82fFUShxllIxQSdAZbH99EB8idyir
uQJGFsj0KmVjyvzhSir1rxQfsVBHFv5TgK8K5yrNW2V0xReafxRJ45JS9mulDxOHoKt/5YAWvnIz
92ezGKzEgJhF712aRTL2DtyCGFJfTOwLt21ZveE2DyM3FoIWUCNIjsBqtsZiHyUF9dcIQY92Y+kv
WldQZEtQGfeb3boulDR/JCaMBMjp0fS39pO1FFMOaOUXmyGoTYnExCufFr8p7non2K3PwnQZ6IFB
MkxKhj/lyv+4YEVkfoo126nA9r+A1eHTI1lbpLIJacbq+L/SJKEalf7AQlnxWlGIuIulnbf6Nbn/
TAJTjX+si4iM945MY5ri/kQJGDHq9kqxLaMiDhu8emghbaTIRjShN4GJCv0fBBp3OwqB7izVndPf
bkZuKHog8TObmI4uhysVU5utyZT62YnYpdCVrmTf9hg5jJKAWjzotXFWYlEK7iLlmthM58vVJMhl
sUUM8Z4qxG0m5kzm28SdtwGTkp8oWtM1n3raCBj5XUqtV1JVOBJkYwVKZ7d3CbTvV2iUtK6PW0RA
wbqE/MDhwiNDx3RAorild2sdtMbGxan+ctkxtRYwPBgXc8wLE/YfILv3bAODBMWOm381OFYvmfxJ
Um3EhD/xbBJrz/nDo4DEWj24zE0Tl7mhN2D7QjhFlEH3th+npoASrA/dJo8RiJbQz2Nl5Da6k9s4
3FV/46woQ0dkpsO5FhyDftFrzU+KxBeoMUb7+4PCPQrS9984soZZV9HKv3vYdJAz0RLY42jzPI/w
2jgrLnFEGf5Kpu8/0pzbpo5T/33QGjrhx0+cDspHRKP4bpBtLe4pH+79Df0nNAHMfocTJyWoAsO8
H+R6MFVzKsqFjUCyMClx/KzsU21FVn3SPtA/iQLgOgxyFAO1Em6mUGm+bDSUUgQzyLJgd09e/MUn
YxeH81wtC2Uk/CCPKVwJCGIPEsKlXbtaMpR6GhvQRQCwa5DpoAyDAX/wZukPyb6rPO6fCtVVZXGO
R+9xO3VNfd16Hh9Dr6yQsUrXuINeGlnSOZMpvEa6gpv4v0cVFtm5a6RjkeBo9DcJgWIlH9CqojqS
fMtpKSB4/DEOig9AzDfCpO3Itlsq5v57aLG4ozJYjrH1jQucQEih96nae9HHCJypsk5CrifOlms1
aaqL9AqW3Ns2zUO7SPbzeNI0ZkUSnuEWYHcfMn1j92P9EWhAfOK+6hJHLUX2A2W1iUuyE1xdB/m2
xCUwof9eACppf+ix+LT7an0EXKRpAXPVzTEqxSfJfrhgDq5fhl6VJbDdRBKOc5agFXcGW7tinVEh
MFKZPPg6BOTSWUx2wga8X539IsdSIZtVonssEEAWDOojN57h2FdEcyl8hvlwOEUsEaePMHdQsqXc
r3yehz20FE8l/FUftSOZevZaSX8IN/4Tz5FQnFUpFSAr6P2SYgn8uUiFG93eK9n9++SILjVvP6iK
tiuyYDs+iwigR+FqB60Mx3rWxzbx4O+FeFfHcojtk4mp8mBBf0n0NDwBuusTHlTeTpPzveAoYPa+
DpnJOm5lL9OJOoP5gOwCt1FYlMaoZ6QP2857Ef7++a4HwE5CpqOYPcCXKbGIOEP2LWCiJgMzui9/
nRMr3H4jygYmdB2YE8xKqxMgTzfy3C9muMm3KGbQCNwmlpAShOKdWyKRWN5d17QYIkkvPmQBLmfM
aZ+e3qyEo5cRUFOgIGR3YPcKtsojeV4I7FpkYa5V1shQMcflJZLQIID1zsVGTG63rRHhNEYuVJBf
CN9IsEroI21mjtfL5GhP3qtXs6pL2hNbt0UUdx9d55QHwxZ0PhW79e4tigcJJ1t0R0ETFILdVdka
VMuC6RLAT/BajrvMZd61vGpQa1mj+IUKnSfVXexOMExXDLYoSN1WyusQmsE+TwAtEpTX6NoE1bd6
jTca7Rx4ktkSqqGOJaHaK6air3vCKkR2y9oujvysYUvAIGCtBDXXwNBIEC10jpJ44X4RGPJQsBiE
qDIHS/gk1XnvVFWUrPuDB2dhneax54XxR6MrIV3nwxzVKVIs2qF1T3IQR7l4Dk80FArqmzq7NE+u
yqq5MHowdya633vf6ldXydR63gGtGLyTqmI+q10eyZUdQ4HhqNWVjAwE1f6YHlOU8idSPJJW3KJB
omRlVIRHU1igQ4mZwkFPL2IjRAECsc82m2NQqlMFhDAepwHno3n4MPkPgRath3A3FHV9ivjGjQsE
y7VMSvysqOikVKPZP2ikdGbgwynyG3ryNHMzJGOYVgCbJUfRPfiSMN7+pwGacxHb8uJTlK5NeyiI
P9NGBc2psbEHaJ1JRElIFzlyOGikAOJhedpqzFif5QJZMaTthibYvIhEHo9WaCC4oOd34QDLCgUN
wm05O0fzjwBneKcwlTuKUwM30NRTAKGimlwnpy1XFs57w4seG9ddncb26I9m9KROv6/HwV0V0HDs
HBrBunL8bg0ZyAbP7RHCw/rYJjAPqzKTos6rJasRHynxWJvAOl/fE2jznuQz1UTBNSLVdbCU2vjx
zMrRXyk1VEu6sjPBRGCDZrPB5Uwg5FIlE3FBAwpjOFsxGRPgEr+5/w5Z6Cu+dlk1DZyikw5dv7VT
YSqIGmTAY2BoX5/5ncJSVe/WR/ah0bvXehtw5WGKitW0ZvkuZRssdKYTENEfPSb3x1gBVaYX7E2O
TdR80qGRk0jJ5Y2vl7p+cu19hYgeTHWI0j7iYOn8Rq1z50FTr14x3ktL8+FYkx8b43cFXn31o7O5
q9pyZb67A8Z4muCNAh48KQnyON1z4HBft7wNhX8LizBaDoygjs6KNfYv60+Q9iQcz+/tnxYkSqCB
6PfrwHpeUYxto4LONk98s0jgtarliHprIMTXToXt35hSDOD2XlBo9vMXqnkjL/UAPp/0bqUwk4Be
9iw6R1S2baIeYv6JiDEGq3Ip/LBSLJt84kUnZ0lPlIwFzSNVi2uXkkUsXuiAydrmrnBYNaK/Ja+A
bHIDggtNFkVrcjMtCrBvYrVTlZizCnz11llATiflva6sCho08Iv6tfiTAVQTL0GWvMqMgMaAK8j3
Y1DInCJjesLcmNpi0HBKf7Ua98YbSPs8b7L5YWHXTHgA6s/HfcNRJmPMBmn4lzb4RmnzYkLTk4+h
gL3iHXdS9rsM1SvAlxWJUyAjeTnDzg73nXg6w6huZxnJdE3Equbl2dK15+Bvyhnbszgrm68AlzpB
XPPW1nBFWI8SMjk6Ny2fOwTIN5u/DX9opJKG4ZT95u+zZqb/tduBw4Ju5C9SZa2D/NJ3hSV4GZ4p
pI0abQW50Y4xSuU5buivUsGnDbLmqIoi7wHhlF9O4qzCs0qqM8mM+AGIBKOh11pvHwt6KrdHfjRY
MIa/T3OG3GuDZyVdtOIqGC9yhjXR1E3Hyvt/YaO8+XSa6pYp07JOgC89OEoFzU/ahuVd1xMk3lUx
k88wlHtlxRbV15gK6cWRFRy+2G2oCjzu1RVffTEaR0FhnOJtM4/bOqvLtQRH2MGQjJ0InEljKDHk
j8wUNNXwbLjcHnkXRokefv59ME5nFQYEOXm77HXVC3VayeB7x+pjPn7ao2q7kJmHvxG9LxKBMA2A
lFNC87LXJdBDA4LycX+XdqC5D5T2Vr/iZrS/IVQyWeGRyRisKDFUgBXbNth0TtWcXqSyN8tB7+Ah
zZ867T6I3bDnRU3NPHqg4Y55VgPr5gfizIeEQf4faG27q3GNnbbJsgLAMX1NRJAOWGaiahUe6NOr
Qf+CZ/xgwEX5d494XYcgwRhYWEAsiaG/HKIaM3zO6p6Y+A6LUEQ9x++AcHTWkBQo2LoqXi3tpD1W
S4q66LdzD/RrySfbAJUOdUM9jrU7OcoCvn5YGHx80soh+F9GWf0fo+PZ1lIyK9u1YzBWYtk5Np/C
TzbYV1AFUWkJQFVPpR6g/KCeiXP3zS0ae7IPpm+D7I09ZRh44SEWCBdydmzVt5LGA5NJhBTaSAg0
uDE63cTUTxXHqaNG+0TkhAO0MQHs3cpNUCbDGhCqfVQBw/J1Qyfo6Ti7Uu5If/MrgQB1eGGpYRr8
Ol9VEZ/6wj4ikyv8B72R8zNBHboS7PVU8C7KV3yplokVBrEMuN+jHua6dpjPAjb8g+ugRG/TIlYn
sWQT91abp6IHczJnhMZwOyl007ZLXcfHuhMNP4y4y2nqS/oYheTyfXtpN1p5NjVtjHQbqdHF+0DR
4pChP/i8wn3vSiaFh6//G/TVbpIZL7lcETLuwAQ5fH5ZK9krqAUxr1zRuCPqk2u1hKiWacknrBbw
aSEKU+qGmkDHmeVQcFg+biuM4lMNrjuV+vYP22T7j+plR+Jw5PGohxoTqcyYsxVl+TadbvSOT5yU
CkbBLeKARFQejQYEcrxm/saZBj91DoZ7B2C1It6PgIqpl+TLH5EpFylk/02Y+xZLsEOdDSd0eo4d
EQTD23CbHzww8l6lD7QBhqDMwxzAMj6CHYgOP+E5p6RLfQiyolgT2Tq1FB/U1iNWA47jADLU+mtW
ExUaQXbP2gqEgjOLdVNa02ARnX9++gtnUlsHtUgmK9U1f7t9uCkphMlxs19GziPkQVmKroShKY8w
IzOZzk7+af8GLk0XFYM05A29Oi7FWKGJi5vO/+DWuBtMs3FJW60fyi/NsQxWEpWK8/BKPxBoXta6
/NMkvvSIcf9INVxXHPe2u+4fbCr3XgFKGUqDJl5wBpJFuMYr17BtbGA70tV0U285Cp+8IgCz9Zab
rqgZQru3KAYrJ+paPmoed1qGxp836qb7MlWFm4GLOjevUFyFH1BCRfnWy2CcbFQ7H/R/i3lMB5MG
TLNMKwb8qdbwU6aqcAdcNagz0vIZsY5bo2IhGWXF5ie4+zbcbh7B1/svRDSnIfU1Nb3f/p0j+/42
Bfqu4AFmk1X2fTXz/RvRqBCh4UCEXVYP824DS0NVj+HGbHTTH65r6IgFoZbo/5/W3uhi1ed97ZHF
+ZUTOdGoVxzzkYNFJXaP0tXjF24uSJl1rKLwIwf+uktzb0KJzSrzKm2ShGvBwE/Mpc+IMEwn66KA
KWAHlK9EMWg8rhr1qxgSI0poHym73x08inzaZmz+Mt98vntkcI1gHVwWxk6AusBOew9ILJ+objax
xjNsLs2zIncYSbCSJdvrYCrW0t8ptAv/i4qnqvknvjcQxlgxVRe9sKIT8XFopR3gfnvvQa+sXm3W
yixBaSQes81jYVyIKFqCGVlImg0r8EN/qPXbveYW7c54CWQmnzZE5kF6qxAgBfFutrn4i3CkKX0R
OLS83efNAZSzfoMl/5pJdaBxMcnRGvAaWmSnflxsUT3PoW07SCZ2dEUb1amsh37nfibwPSfefDQE
el/msEbvuQK9eva1NpcF7+D3sIhnow2lu/76H7Pmf5eqx1dy/1V6Wm5VW6LWNHZqEvoVQHPFlNFd
GX+/Ql+1WH9Bv49N/41TCj0/DAno3I80cNne9YzolUL9Kb+bgS2tXBeKsa7ldyNbjqReHxp3so+r
mP9nBkBiq51aBa3jahx6G7YHvjuKS6n/qt4XFVpdxqCnceX/qjW4nD+5uhSUmrRHAfaDilQymZXh
adl/wOBlZT0j6UNOyrh5JXFiY82MVDdJXJMI309HRVvSE66PGmBIaWoYpGohdPjisx8YHnFY6YMk
1FCOF7tZW73g1UUM74hFP9RXVcvfuzxQSjh+IMeTwP+i847znsMpIYwxFrKHSj5NbLuNBRIjCxI3
sP8XqpBe33peNsEa8X5W+lic5ftTqLH8YM70PL5Q4Ffoonn0fotK+QZ974VHMOgwo4khzmxgdloi
CTSccRu9fqcxY1099ym7wpyK/Lv9P7H9KO53Uh/UU2H4YVaGuUWZJduvBhrODnk2UHwYrhuAYwgA
6DLsP1ChXzrkAUGB7F/SbJbVp7l30/asS6DW4qOTtz3bm7jz1cN54Ff1tcm1YsWgeyyf6tOT9IIz
iGhzj4WBzNA5LAwXlXmonuYJNzO+EBjdF0v/+lMTWrPGzA0J6BnncUG3QWUhMv7kzPYbs1hbqpPb
oinraQbm535Zg1yj4CqyDYXfYnlNbkOJam/YV3txy+spytsi9zmFxg7w3rFQ933ryCzDOwMzmvqe
7/T1I6MjQLTLfmdkjtUP40IWSGRqupO9zl3cBrW151+nGvjZAfINDIH93KoT9LDFDH+5bTAEmvbk
Y2dK1w6sZehu9ukF1F2UEQXD6VZiYYPZ3yE3I/1BX5wilB7ipjiFgUJVecH+e91tLcOVNAdiy8rB
Syxk+sx82VOZh20C0QagC6kuWoky80LCtWoBgragVd+l3SpgsuTgnjUCvm86tS+6b+6gbqOcJ0/6
mvJvLTs17q1YrHScyVV7mLPwxfviZCKZltKfL4h+xO0ym5mGz/UZqXq5IZT9DkA9EbsGu6MOjDEf
wHlJFtag9Tc83VBHqBdSsreLs7GU5SqsAtIMXS5bmhy/P1HzZGKEhVbRQK8lFKFduKVyvp5h1ksn
bptZErEQ3SUVOhSxF8zQlglvgLJDDKZTmE89nROtofsOzF0MQbZTugAZ7hVwxupDenHStLZnQbe8
kMTlLibZysWjewuWa7yiKgUONXd1FyOU7ymGBhxzyD13l80+KaMtApYDEYr14Zk9Rn6X/4fx5TAF
cSa+pgPa1n2tlKMH7iad9e+XsnkYul9GhJM6eOO/awoRTEOzQ+NLr8ZdWxA26Se37fCiLmMiP1as
og0U3GeaVqwcP6aFKWWdIHU373CZxzzGqqUrug6l50XnNE8NQQmNxvyMrXR9ATc1hIkP32crm/zi
GCwC4G3thMChPhKHZ34zGUL6eu5e3ZJqzgNsIJXa+M/nuMkTeqr1HuECHt68j8Ck3ZYYcBKTTXZP
qugM926uPYZnBvZIRW23GOW4YHapDiaLKGBLhYb1ixzYDtLPYq31NKkZbmHxEniv2i/Ssp3TzP6C
CABKVs8+pUUQznDPi3Sw2yJqk5eENKnF5HUIS3HzwRbBnW3mjeQVk6I/mATu86EoOaNe+mkESsPF
1sTEA3EaJo+MAIlxXVXg3756Xx6P6NOKCC5RMtXDF5nsC9VIOxWYEogLPfsv3DUmmvs1+zY5U9rv
XgPw7H/2FgYEJSf5xnwiUtucyr5UWRHgrAK63dmyhEa23wor/GI6G4Ms6INAbWLaGqJbJ2dA2aE/
Syn64wPdzOPh4efvOxg4L1Hh6uXisJN44aTK4bHD0iM4mnh0nL4bLil8WgxPrvtwBu4twCVMmNxD
NDz7mUeLwTiBi1any+HvQQ3VgCYUUYVVYOLeBaaSsCbNgSxlIuv3ilrSChPtTk+CPYdvEld8BVkb
FbfcC4At7qIWuxViuTaOJq7d83bOdWzZE9R2i3Vch4Pk3DPBKOg6ch4T78pV01Um3UeMhTx1GKJd
EOLNbAcwnBbi3LDs3YlnQgmuOWEZhdm01y6HxusW60DWYmgJl9mA0QsYkJ5fTvgiR2fsJ5gT7ccq
EDngWBPiq+mDoP1BO5rV4enqmw/r4I2JVo1taUAPlmLGoVOm7PTJSuEhz7E6zJAMFvsGHhtPH3zX
GmaOBh0L4UOMVybxfgvTi9H5fv6QY4FcZqEBoZ75f4g69tS+9x3SralKD7LOazsy6yX/+/LbFfQx
+Y+r7JSmDWZ7fJNptpY43FhKjkqHX2gKi19hwzq17AcbeCt7QDkl5XBMCBTtNpmFb14HJdyvdV6h
Sbq/o3iUiWqQTbxVtds8+BflUsqP6Vc4ikAacz5SJaNewaNNfymi1WLtwhnTCNWeL88mJ4YuUVSc
pj0Kb/y0oq8QPljnUtOxBcs596oRYy2U4g9406TrsHVDlXeiNQPtWS3pT3E9yPADjCSTqPzm9VQH
E41PW70akSstjphxfc2qeHHmXS6+A1d6xDeZSOHYHoMu5g+avstBM0ToB8xIL9lfsjrm3cdff2uq
qkhgqHfYPmq2iMEscBZH2DEVhk/rqT42d+NNbfKDkCCi3TwMviNMJbG/sVMYelPHdZMmAKVKsS+L
RDn2Qe/hdt+JfKi+4gCJYHgEBoN8hIejz+Mccs9x/lKtEHjzEsJiol2HDgcqz8tWgBZfJVhhTcP9
brWEv2vIKRLItf/L7qydpX2AbaS/2WmOZ2ZYmiWW7EHqe/lVqGOfVQ7SZILeJ65WDGHQpd9xaPud
l9+SYdo99EEhX+4gvgrJVgsNDDtyttAJvK2GkMHFGItgtm51LB/GyyoYlx2iAfhQFJ3ODhGgV8tf
ZAMOSUPB5+9njalUv2esE07Q0c8EL256F7GfiU8fckuujln5oRjqtgnYDDSQtjuRLcgz8Bx+ptLl
DwSLs/ybigPWCAjKel2rJFwPVvF0GATFVs5tirQ5lXQAJCrUKNwTsQh5Yj5uacjsX0uCJiZzQrve
QEJYMEGvdhYyijvfHHk1tqtnfntxQrx780a+bGZtBK2tVTlzxxEx4ucRGpSwJeByNvx6XiuxqhuO
dFf1huaWCIzpiqrrvn0mLN899NejeeVfPXq/nKDHFjgOImfOM3iOARV7mx3pVhjNzcCLuYgkLDe3
vgfd6jhSFCgQ5ywoq2Dd5t90orLJ6XvdMaDeNFuIcBjXm/JSwqWDyBC99CFlsTv5dx8u2lNZf3JE
TGYKPJlc8rmWubQK8g8ed3UrDWhj9ON9izErb8TWe/b0zzNSY7PvTngjxIAQaVRkI6WmFzl6+asG
hocAuDU2471lv04BOralsQbWML9Sz5woSvNgTXlwCfGqOIczAx7w+RK08D6xbdV9E0CO2QR6Tg3V
x4e2g3zaPGNlTt6VqkkG+/cADdbXJoghv2jQfU8O8rWnp0Ri2P/CCVrHi0EMb2FlIUsXYFIFRCgX
RV2c6oRMHhNxkCKLK/Xy7Oo7GeAF5SiidSHj14JKLNM4VWTmu4b96yK3LQKkc5fX4UDQU48MJ5Qm
Qo4EGTAUOZJTZWw9H/cm4aXnBYWrBjQ5P0O/2rjc+8l4M1HGMMS7anTzfjFFcpqGk+PRvg3ePNrB
ePs71OoseIFsdShey+jmG+j/v+dkht9s+r0nqhfI481B83pYfptFHvLnmDpK6osOD/8BeqN43dX9
aF1VLbHn3hgCOYy/y3qEcVo5U/3OiZ0OEwFxVhOttFLR96FM7e7kEMM1+j1fXxhfC6KY3e/FHeWf
5SRF8XCciVpjc1SLGxENJqqnDtwZa4gz53fvp9mcNDxj94FVgqZ8QzzyRGvsDfZ/idq+3ZuJxDIb
/qylb2W97Nt+2b/1+UlHyTdtC8pIiusRHXeRxGlslu3J9Ba7pLLX3jDwDZq28qaJ3Jc6MprfWiEa
xIuDQyrkJ1mxCfHny3r1RSncSiIJrZ4t9cOTFnTGQNi1koKLOrcwvU+8KReYgmS4iEWkIDPDHcn9
Sch8tlKZaDQcWI3fsMq9Wo9iHyodJBV5tRIPumfuya5kh9B4jxWEBIYMYDUc2XsR4VOsvt5DE2eB
Kp1IYG3+bJ7eeE4gl4qfupTCaTtJl8f94qetEW4jq/2oUfQnCDVmZAxG5USrP5JNYeENL8l9MexJ
Kl5sFoyAYvT6FOfsuZ6DvUg8ujJkYsBVMaNUtqaT3Ic5+QtAWqAiuhcvVI+pLDAwDfBm/KksvILU
WReBhHRjemram0e3HrLpohn3mdBsQ6spNIntRoZlQGSNlZpshtfMB/vGaAA7MJO4x4vIUQJePExa
xCnxSxRVF5xYSwWh1AOVUqKCzNbwGTG1+u/y519Bc6lcNi8snA1vIbT/88cNjoYolWSbz4gLLfJX
9LKJeteHyjao6NcS63f7OF0GUWppTNXvkYgY3uBSTH+qOSOLxpG4x/0sMEJNbuhFobvxenNP54eu
P7FGq5xI0/WIOg0F87AUDPhg8UPity77SMnTERR3M9/mZn/UUrL0E8TmECJNPWJdXpWtRqKPOySO
/0w08p8rkHKA4u2eO+s4PNyfqI8RZV5dKKB79x/xXdtK633Wpy6yL9ESB7HUGthSc9dBaxI/nKe+
1eY5gvpJeEpSYjprZM6wy2nNcaHf4L0r4srB642hUtt1Q/GbDdtpfiIDE6gLtRvGhTZo7jWlgpAa
nwXfjTXz0FY06YmeCYQeFSVhe1Kbw/vtHWNOodZiW7nAv+qAU+QunhAq9j7uXAIx2vxhVZxgOgSh
0Mb5J1QW0rS4a4NbOwnuyiI9DtMDCwslvt3Izm7zxkswlAvam7CdigT5SP1vEsncPEnYiwXQoJcY
2BDt6lmyu1yr5NoYvzujWbep90gXj/RMea19HkzhAnxEz4xo79Y/VueXhnno0/xs5Byc9dWf/iWq
zLHRVpEkTssJUfTBJwbRx7do9xhARNR9c2tUokFDa1ZCLdieJnkbUj1Ozwpn3EAEGkI9c+zJjJFm
f3TYienhCBskBSNDR5WaSg1k8//sTQ3lyHdJ1zPoSigGJiSkLKQqF1+3+TkSNin9AoKzYn5Ta94n
9w3FYy6cl4/aV+LLokjw5JUlEcmaQd3RL74A+VAq3SMXTDFmopehTO8lDVX4uoh8PByadO9B3EFh
6o98YJ2lkt4imGufDUPIcO4oJFQdCgAStyXyc0TbORkCUTGvEMEPJRMzdi6UdbgahTd+5/NS+3kn
sUtI70rKxq4EUyeN3gxXqq4+ipI7kKRMUKnoPSv8RHvRnwlH0u4Ws5o7dYXAyFTm/M/fY/5BznDi
wsAFFWCjt4Vd9nTjqf1ioyG9I4Gl6seCkGjODPH13hrXDpiwI6I2U4L/QvPcGwEtIJzQ4AR+fPsH
2wNDtQ/B72RF+JnuH5FTnxHIz3chhg6+xC+phbXJ9k7ibr/kGhD3qAkq/1erEW/HZm2WVSxs+pch
pxJXto7yu+0QweyvXBev4hB19/G5OsZ0x9Yhpnh+YQoRg5jjIv5zQr8ucSJfazc8w9o14QU01Hnz
rWtPKtBCunF+6X4hKoAOjm6U22IprYnYB9ufwAMV7zlYDObU/EiG5i9ud9Bn6Nk3o/tXw1NiJd+4
EXnA9Wpv8HTXnbQVbnVduFpDcYz5x5BduWz7wsIKv3ZifgXeNRd5kOj5+wXZh5t/d2PwLYpeH7Oq
18os3MesaS9ZBWLpJ0EYcW+9i4zO4eSjFCDA/c+dec2A68pw7jCsIIFwyLB6K3EeRvJQcpQ46KrJ
1FgO9wvlEF3Xgrw8R27NYOYAnj6BxTxdQx97PjhJ0vy0HEHpYsm/osMV8AnDI54PkMctCkkUljqm
iSuRM5EuVBarQOV2M6OM4zzwrWOG6ZmqcvX0HcVojMr+rP28Z1bQbPei0rwHoYsvxznSJbAF7XRI
9E7Ea8Z604EvKAbUyoZjbpgty/tNXSA+fM7IfAXo4VSH3coBYHq5qglAZLIRxWtR/MwF1OPYelsb
35yh0VBAMHWgNlVY7GJq36GlkyVzhMQFKYUNSyxqQWxnZKIMaxKviZWY5FDJrPD6qI5Wm0Bbzd8N
ljrjtUQ5GCIN/ftOxMG6h/QrAqN/f8mCqgoBtX/BPr448kA/fNxEZ8vyCutDrLeCsIw386GwoABj
u4NPC9yq9h8KUaRsOTxRwmI/VKBPIv9jMd2HolUtBdLO3dnPvNPsxVkP+5nRhkQrKajo/k8FACQH
mquwH61SkFm/yRaWKkoSEP3on9cWCj6SoXj7kXPIBZQzm9pkdF4LdytTb0d5pP/KH/iPoPYBCV2o
zuQLmx8EewCUGDb0oyX1iDWRIhAhoy7W4uFY2WxMJyzhs6tPbeLtNvNH3nXKi73QzCyhY/SXiB2x
hyjyttSxjmh0B1OCrXsKd37QxlNfocq1YMjW8eyO6Uyr9jCRC63e7sUpjOlDZJfPpWggq+u14V9y
Ksm65QpHWRS89AGYdnsD3YGXhlIir2wh+kt0SpNAQoPcNWg/MLzJovUPYiuhjTaTtqB4qhBLSDZr
sVWe0RzycdqcYQf8Zb7K8pw+GyiLtrZEqr3/CEpn0h1JyssoWMxSknjsTkILvu2l6NWJZj2Kv+q4
plLcnVRroSkSVSBGD2GX2F2yfJVrWZhZT4ZwM5fVurqEa70cMdFvgfL5Pn3CtiAzMzABycLOAqEv
+t1rQ6OJjFRhhPHZzwb3R3G2NDJzsEnr2+JJBlZrBtXSa6G/8CKNZiXX9En4OJ24BR/PxK3vYs/U
/sJ1V5/NYuj9Ba41/+TWfKPjKgl2FBhO2AzgTiBe/7My1hPh27x1X1LyILGQ7yPPdcIJR7POaYtl
1g2im9jb4zAhg3DDHglFq5M8qtKrV2MhRL3bDVkRxSD2ENjtDjIoen1n7syxh0Snsnf/KlrhlHsK
7WKyV/mwV5APiIpwRIPaG8IW96z9p+zyRY9UQJNwhpQm14dkexZH5B2mY4wBippgyGub3Om42Mk9
IVgtPSKtbYlxNvLCADv5mJNVhf677nDB8/9wiCNEaakW60ofAOg4Az4zAT0AGBcrSu7qelw601Hv
nBxQw4THBkGUPXBHQiFX+BKVS0hTBdhS7orDM2zoIPm84GJCtyGr1t0/sLnFQkIlfCGAUzJkVRcb
9RGllFVZRUyga27Sqe73/Ga4uevqKBbjL3rxRKL+ILQtMRy4PPsu6z2MQwih9ydBkvdAL0H7b3xc
z136vIDYNp6ESSeJ9uVda6h5IXckDmjAwd+CKYRIqHdbgLlQM5XfeMSKZEI6REzwKAbXUBIAEvUy
DGw9IT3zTtM3DmFnwkvdGfYHcf8eObBEODgTOERn4blxGCrlru1V/0xI/rOFmUqeSDIFIienLqx3
RNyeirFkcp6bN7MIlOSvO7vyfHg7i3xCl/Z9kIZEd+RBWh931ATXmJ0Iymb1MMim3VRkL9EZPc8c
5N4vsNcr+Ksp+YhVGVE8FQrA38ybpDOSJ8IN+jaCV0k1pjyxSOAjoSTwZzdY1w604wqWa3Htny60
6b7Wu1kvaLX7EfFmJ8vzbU73ZrZoU3vO12jRCr5msMASktupQONUN1wimMaUMsF5WMPJRnW7CiNT
rZGlUBsE5Hb/gtxvPr0qwYLNil01munpwb2wl/3WLzuexxC5f/YRGodZuHdZWdrRY6QQeTva1QGS
fWhmkuNW2dYLpVKDvLMxH05qFyQDpkMXs75lGmwZwK8japu91THBKrDBg1/y5jPdybHK4fng1pfR
whlaU43x9svgKI+BktzljWKPanZxx/uTL0/4k/InKhFITF7HhnbbjY87aDBPYbzUznp5VyBqdKxf
1fKw6jIz7Fiv+Gp3vS7L0SkD8lFoGt/VTMCg+wjYgM4VAZsgB6UIU79M1uZPaVs5gArbRPP6L9Qo
/ifYb5sI+CUg2wcNlYpAEZeXgSJiuSP+lWjVVB47oBSPBPhY//TyxgWWIk6pgSq507L03sIsQ63u
myKwmR9PTR++aqE+1SquqnVf7vTfWXaK/CeLvc7rMpQUSt9vojKZ4fKjwxKqf5pOHSYyi/EsH6gW
7sdJjVlSOIiHeH8TL+V4wD2v0/BByX7eWM0aLK2ndqChvUI0sBL6aYLGb+UliuL1OP/f0o04t7hI
XWOShMFlr7//851xodRuqxAl70ex3sjNK3/cO+NG0QpMCsW0BItSruwyAnrHWCCgsDJRmbNyd8LA
XVVvwxa/EatVNxA1pnnX4rXBUrvEmYnPDkUVRsnfN2XO9acFU5f3GV3cw8mkj4jt1p8Yg2PqRpD0
eaKbKajs44NeHmOn2DtaxMqGyZGDjAS7vR9URjLtgFLNgpNd3wx9EuM5HIFCi4r2E09Y+wDZSPZ5
Eix3oHFytifkhHzfWDq55nEADCT2ZsjwL7YoX/pBf1blTVwz1VF9zkmwdcNq10imBc95+XGvgHg/
5o+5mLvudbggng45VKeUz7SKdlcz0dhKWdE0rtdif4mw7Ne872by87Gn9gDZgZrfxHVIpNIY9uFX
c1jpXF80GAG0UHFeDaTuItbG24zPsyly0j3bfdOSP1VmksDHWTRtnuOlu9ezBlZO4eI1RO7GpmnN
BOw9+TiGCL3x78BA0ei97GNWhIVdh2kHPOZGaMknGtfXNNMe/5gAiIhMzPqmrU+zclzdwnS26LZP
pmVuCa1l7hhMkxP+dDULRXJXtvmhWVGloYcy0uN37OrtQuE8hCkGcITcGIj74BLV4NcFV1eqeq+l
4t/7iCJonuGjQBX5UBvq5v1AGwN9MLD/Pzr5YASkH4ocvYlUl/6+o6/NvqapYeth2v6aWO+M3Sh1
MHohyLaiVKq2C3b2iXGBgE5P1e7Boiud/G0fw52xOOaxunIb6GTjEZj8MqnwxtxD1p3yYl2Y4TH5
NRWpmgmSXhGJbXvF+FLuOxu+zC1u/piN+99YD18QBXnPAp57tWP+LE5jUXilbStXix/LAi5r4p7s
DLTE6QkrXERHWpjxMEI/b+2XkGaB2b3ou79yKG0yLyKkjZDLEOyacF7wuMW5Tj/kh5B3JcOJ6Gr3
7lULtqZCi7urBs+FR+GrrIno92aQCDWSCfD4AOkV9fKT345b2oHM3+3onZ09HplCZxGuhs/gaMe4
7ikq3v7aM9+w2vK0VjYiYe/XJIJa/GTZXqORAU26k/wUf1SD0XAnbfvSUzeseWoXEsbzzGRL1Op2
mvGUb7xDsRbWYjSaw22GRreZ3cflvR+F4oL4C190nEjV+wg10g02OhGJ5sVC9H4rAoEziU2PptRj
f729wiVWcVdJqXbz5HozDQuCyunOmYPO/Q7jAXz29Zr6sXlgtDgDe62TAJ4E5LzzRrT8v4mbNwd9
GYSW/RN9iSGi6ttdlGelpnd+HsobXZv/BTmIAVLDSrHctiLau245vpAO2GJTmy9dRZtt7jY3jkMv
e1baMN/ewBrplNqF3oW5xdq5tVnBuZ6SEuiAs08u15TSFRrkPXkg8SIKT1xYBe1dKyiQE8OdG3KS
hQeeAB72Wr9vY1diHsYWEjtLH3Bt6GtlM3uDhIMntYtnnBkM6Qi2W3yDx4XOc7KtJpftsAi4ObB+
xjyiFOg2Qmkf6hqjbS5GfUjK7Xp1nfbhl90KlrUT2GqLWipqbhYbEGQTKWpQIj01y0RUiRxBwvC8
MZDs3hwajZjlLZsCl3zuuK6C6prezXPDFUWrKT6zwJO2MkSQMhD2DA3Yb8p+b7/1Co1qmuhmYQot
Zy1wSqrJ1j906UW14uki9VXJLTEKaupy7vV8jr3aGFArg8aR3sBE0PD/grNX1lSKfQD/4a72QhXS
QvlvIzZaANvDi5WNWcebxG2WtcAEeKsjfdXHUOlWobIYpqLqnde2A5SPERp6j5TkqAMKb9cQYoos
z6aJz1V9LbIAlEyZ/j0F/veAKnSc8TdzJr8NqzQtN9B6XFlVWa1/ycPD1ocYH3JI5g25dX/Y1eMB
04iXDuIdURKo9nW3s3SHy6its8Ova7hJBp4K0dC5wVC4685Aggl5kl8HdKIS1CspM7CxNeU8PnDb
7g/QFJEQ6w2PkJxHJx9c1s9QAuUqPjM/QDVbLOM3Ge0bkqZy3+PF3dbwD6CKJV+CcZ5v7OOJ0XGs
WO3CAvPRoMVDdnUxpjZOhWSkhEdmiaA1mZhdAx92PblxqlbkzWZu5ivwoSPmMUiPv6Pg8NPXBvRo
0elPXqM0yaAYwo7yOLWIHYVHcBF7qvnXGCXGKqE6zB1NcksTX1JXWIhXjFxd/yLIHoZMOk1xmlOK
MLtNNvtwnYoXUU+xJWm/npexf8l2wJm29mA0SeRNKQRoUtrRw2nxXvBIoPk2pUckt96H8Vr3PXLE
oxEIArZiRpgbxV4Wr/2s02lvv7ktUeckkTHu0ZFv4lspjAo33ELPk8kDRUtBThoHAM7ZhSJj688A
9aS+CJmyAM0zQQT2k5Rn+KG+K4Qj79vghfTGu4hEOwIEsuYQZu4mkQFyN3OFCqXEt/BDrXYKIpWQ
jvisFgFTRXxlq8gbgFjddD5GIatruhIOBK3CYST1yeaxiM77y2hOx7As5k4uW0XJH7pB4I7YqNPP
GvhUj8nowfV8zXen38A0CFlFDCQp7iaeHlDBs1s3ixD8QJXrtpSesVUNB3pa/rKmfXsnuht3zOcn
FTeMu7q7nkXllU/fJUbYmeIEbSo+o32mlam3yeWK6mPQy54SnbDKiY9BUc8QI2QIk8hOBxNu3rO7
QjvlaKuxamq8SjxBqrlhgchahkfYxDBJalx8yQxEgh9BWdv+FnG6ZYLp/t0DXvuHSvVnp+xnsm7v
Hh04SDP+jgYLovdKoxYV8bp5V0CMj68n+MTevlH8D+laSYLZ1Su8Q7BAcZXv+E6ndtrf9W0/HoFI
UGKacjShYVSTC1oFJbLu5M7CreBwKZolpTlun9iVnFa0ajbTD3oHG3i6YhC599BPERt1PAk5k2Ai
KPfAA6eQg9kvDX+bbRWQrefB7/TgF8N0/seGFiVyofhUBCwMQoRJOE8g5b+pYAMtpo/zzHdZ50fc
dGGBbKp3yUVBnWFgmGQHWyfQ1WlA2hUuZ4m7wZntatrfbyrQ8mCGL7dIsQ5AOE6DH9CihHHLhlwa
vCxjNaGvKANxn6Htif3onzeamJSxUfwZKKGfAW8tb5r8/F2Do9DFdKQPX0aElCQE45IJ4nAkBRO3
y7ADp1lS3XQYTG7nmMnn3ynw8qU3zAyNRTYtR1V2HfRuZk/X+QtyCCbWBTgLV3gdWR7nb3ZAZCPm
LeT7ExyGYVtES+kauywJp+JbUR9jFty7sFX40neeQRLrURoDVSCn8xyiuEIagXIyPMBCnVeENZhv
MYaoFS54zXbPaLepkLaLUZDpm4QN2bVVAbJgE8Q2CNWL7ZPg2Jd1WVSPC5C5idxgQxK9pF1c6sJg
on6SvkHQQpEgLU8+FYq/fnU80AiUmO2/dwMGhialOoiyNsdYdVxpn+BY4ihqJ+jvUCcEBmV+gLo/
wK5YLD1GePlM/5X7Hv2M1DOstTxyibONm3sYDIXXhDs1AJo7rxFt9fPqhVhjEUXrZwE+KaP2tL7f
gLTTXTXYngZAi5MISMDAEFGIOjUDWZKhEHzGNziXYZ09cWK6gB2kFQJjQuHChRmBQNkwN4nrUuQO
kTubqMiSICTLhbjmlALkCV4kjOIsZstkdm7wbUJZ/rc3yhMol2SeFmMmm99ho1pF5Z8gJEmGn5nV
21sVMNXvBKi2t+wYphsN00Zhsu5yow9VTDoescryw4AlPpnbULTyVcRAvQ1adFBy1B2NqS9rfbCK
iTQNIfy95548KAhikERsDmktQ3dJhKOIzhjNEt25s4YGQFtuXzySFtKITh/Rq7OQ+Yh5+SMCAkG/
8e56xhIFyZRa+9oUZBk7SmSqsJpX2X3mdcASqiVBBLRwf2VBLHsGy+vgMuqqSVsaLenOiMSmeNKi
3UIQGN9D7QOjvhw0xpx6/xvKIBl3nocZ+iapgtGqwQR2d7Bu2BbhaJ241awlcC48TRMbZCpr8nP9
WIjAX32CF/CSYVFQjzDK71gt5aws8wn+mdoe0A3IxQVMGa/ZyXnZ5ahfPqj1KMbo7rZnGLWWbzkR
zEE6MD7K1XgIBy6ACw2mtXAN30+TdDeV2/3VNGkwvH8NlIHPSljAURvUKjpkrl6dXTxtpHhp+mBn
Gbzakorw5XKnYz0kXIPjq80ULnjNfALbP1n7FfjB8voUR7iqKN0CEC/7okWYP4HFSLgOBgs7CuZB
Ol2ZB34vR05aW7N7EiiHau6dLeDcMHOhJitSU2hd010ywXPQFr5Mm3sjs9CeYnMpO5Y9oXlJQA+y
GzUhY0tzSWd8WTVh6pU8MWacPOkp6r7dJwJLNkMwVNgJ46hyUyHcmz+1CuhXirBwMshs+4KSfDX4
z3vh4NM3jY0dKzvt+zl7jGroL67MXaslTeXW9En3hIYnZGF/bQdyqLeAgQhTiJI4dvCeRggryuQF
YHyOEc4b5TS+44VUZ2hFKlbI9WUQkJbxcKpnMJlYqAzEpBjEqOwdPyswwViEEy0lRNxa5wmIOYkc
BVT/AnDBfdX6R/g6J8mHeMoRUYFtrX6hEo9ym+blTV4yH+ZJbo+y4nfSCBFj7mi7dxpqlOTW0L5u
PuQqTaMvXm8Sy8fFm+IiOi0g1n7PMIJ+ba47Yk8yDOC6xDgRh68W+eXAGLGvDgg7JOLzT4V6+vMm
9qAVNIstbOMEvtCGJ4jaRzCbrS5kWDNfIo6Pe1TCNzgTO/pfPBCZuPP7VdOQZl6YlXGy4vgifUn9
2uoUI5CYNCM2V8VyQ/807eEQ35QtF4qfg8nxZVETKFHIUXkZflfg/6bICwyyjRUnu/487rAGb1TD
IiltRt+EIkn4eAh3kNm0um/IT8ssnRnbExtrcnj0S7diR114MaDh4eeUZTlB2GJvsXdMxrG6+33K
ZPE4xzjtd33FkscyhT0NBMkyt94Cybrq17QoAMBctshrpcCTZTaG36eFPRXc+4hklLRSrDTzTQIF
iWacNZU0pKu3KDro55raTM05uvBDCNjNffGB3xe8W/8Luh88kg/saf4hHoni8j29W/mlPME+gfsq
0FCSfBNCuEjiYQ+aY1P63arQD3zFkGmagd2scKc2yxbzXb2mv4NTbWF/Z9k6ysMWmF+BjDret3Ga
ZW0dvtiwpdjfOSJuKYUgseoJHw2T+w5gBhlpMKUBFkweUKEeDyA53Y8b6yiHzHjnVVLFZbsE0l1h
UzT4Y2ugTSjiXE9LxVXaoNRSgRkGetZ40i4I4f6oYBtm2fjFhLr2RCyRoG1FPwLmjJlSFetpNqLc
pf6ursA5xiVb2GA4U/2xg2LeDwNn5CZXjwGiGdUif7oQ9wtwsjmvstU23qtjvmzfHa08aeQiNzKz
rJblD2CSjq/gXlsU3TGrhl1gOD8aQ6f5rWCAiHKSjQEVYp5SFrEnxun8oC5q1BmvaDc/c7it9F3e
fka+U3e1PNxH4DPWnZhDeUxfsS4gUDg/5o3TJ1aJd0oVCdQ/3Jppyn2Q/lgqXKLpUqVTEBALkOxR
WiJAjxKiFnoCxQhsfR2WLVPWIq42ghPr5NV5Wstga3DGxSu2M5bQg6VlWP9VkmBenCaus42Y0R0m
yYNVKrRkYDXWKxY4zenwp7xQf5NPR+/bXlfOC+9x6U7hKEB6eicVc+b5aqdSeEB9APa/rxRof82T
BILYqiS8iSwMbM+2c6IxQHvrtld0CZsvUlp4Fr06SoxTYQdBEIBBeHobpzisgBjsLWCCkM56O/W9
HHX1eA9tcppNncF+hX7TA7xQsI7uOTtA+LSFl2lJ62oVJnK3xii1BO47QKL9H0HKrgc2Rp/60mwX
XbtUrwavQfuikSqtah96yYPTONnGJdaxOGoOajo+ujn1Ui6JRTEAr86HlEZFdkDy5EyqVE6EGK9/
tXEPNSDA12VU1YlcJJaNxPsvN2XlTmXIKA2a8NZC7Cnf7OKz5OPJ8w4MmyNiZr7afTbTnZO1XaM6
kNjZm8ibOCx5hWV5T/IxBATU+hS/Tv4hDwVzlcqok8RST3Ngw+zKf3DULhHe+/Usiyu5f2DwgbQS
Bg+Oeo2JBqc8nPtzDQBN/+BVBdTfTk1dN1PfPdMMRbpzfUCBrQ4rgq4u2g2RwafjxHhVEBKd9uE7
4vCC8Q9el1X3ztrv4RQmh5o4D2ay2qI+aRhCWQzRNkkLtFNNZbkLKeOYiaN5GqMpGJLs85tRfRnc
hdFbho+nTGZBVlzcH4NK+Kf0Qjj0c2KV8et5gg9PJapIIxIFl6YQvwzSO40kgfrAnR1udB8qbpmN
7lBUBkdiew8zefFw9A9KjGt1Lj2DE50coD79wsJj3AVCufM9C8wVDMgwfNHiyYPyc2KQZnotaNeb
8pNz20vZyZZWWIVenQqil8DORZCrZ6iIu4EZ6j4F0E5avDdpKPtjzzNjjkXBRpdnekYOTbXJevr1
PY2os9ZdeuTV2DIJvaC6GIClEPMePp9J38rC/xyhQ1z+Ien3er9g2mZ0W0PKfrUrZNGji+MeToXW
gsc7CDPoToaigE4JD+/j7LYdtkEzV4TzMRrgypfNoJme5YI2pi0DM/+I3QxMBS65hI/O4PrnRG2L
4Rb/EQsElwXk55shUVAGlVhzDGsQx6fA0Elf24IwZ8BlfhiYWHgQts+zgjzxffSncln7o8mdMY9L
4LbncMDwYjOx5nT5cqNg2BX0RkLh9tIbhBZqNrQmzfqIoW1VvNvThZn9VZ4ESNnC9/vScjQ+MOcq
+fIorXreUo7u0xdo/80U4cJTP7RTno09NCCFDV+Ry7LQaLPEtwmmC6pD6UAXy+h8/SyvEp3FhbAp
LTx4OmdSwxnlYtDyVNvK+V8di1n5A2M4SOHsyDe9nzfRn8jIVONjRbCZ4f9bpdfRTFA6GgWTHMRR
NcBWRIaSm7zqkDMy02ZkQc0LNO9qwGciFg5XfY3aUmxwRk97DnWGdkeaTOTN/YoHyxjlnZmCDM+L
R+hn9FsZiXjeFfdhYvR9+GUIDv9OgSIqB6f16SauvaebnXkFHGvHkvnInIMCAlrXUwJtoYAV5iA5
6I+uIRWVfNGaK6lzGd0yPWU+kP8NoAYgHznAxA8swCyNwLRyO/qH2O9kkQl8IN/ZGrz0P5qY41EC
trMbxawBA3Ci0QNGPY8bg+tAFL967MzmZBN+6OgOLblhtz+fP21gdMUnOiuwzEuzI3D2rBxCJFPZ
uANUtDJY9cBFWFOycVUIYa7QlGwLqHdJMa1eoCIu2KAF0kcC7JplSd7ArxuwBeVxr0UdU2sB3xIM
IoF1W5fLVtNA9S4tQ3Yl4REv9Vf+H8ajzfRW+eQTLDLp9HyxnPN68+Ejp907R0NvpA7u0woYkraT
GfqCotFcLHwFg/+Ss0oea3pKPja3241hbgFJQ/CcPHQ4jWThnpMC/WAKy3sDulxQYNXKziIhnCDm
TB7mQLEnoKh7qcTIhXvAIjeYkvrSVA2PhjdswsjthEJN6sX1sIsEJmMg5B9Nnv/HAwDfNm/+vT9x
R27qerHlgo81ljdeXBYn1uCIum2fFkdoqx3kREJI2bAHMSgGY+DOAgo3cmGZ0QtPeuu6XaU4JPx2
3rP1hRmFsnHlhEsPB0vp1saT+CiiPrnH1uFFhzgr1zCYgDMFbsA1sYnhtk3mthS5YXymUqNAxg0m
yw7LuV9FaVMH9WziNOXzwPUaxxLZ3UbWEouPAqX4TGNha7yGx4JD3ojqOU+pUXV84hYuO2Uqco6X
wQv0f/xcDAJ4p/3qN0d0u9BLIFZXh2861tgmTNVhh93WJpRAeYruHFDZAJ7dTn+zzrHsONIlg1Ig
P5KFRh1BujfOt6pSTQyiAK+Di4k6jskEOrrDfUFIV1qy82RtYbydWAE21h/m6qP0Wb1x/dsz6W4Z
nvXuJvoY8kCGxafIjvxiO0FJ9V9z9WwJbZY3Zrff3iyM396dN6TaoVnia8U1/nWvbXWeCou8yArj
tqSygNiOTWhJdWIIz9dBWJVgXllDsHtEdMz67kZau5zH18Jws7e1QPpsaBFdYvy2uyCeRudzddqu
wDQB8gIBWmpcj9cICoTEIUoyF34Y2r1DBLi5IMed+hhWSFpz6RKYy7yoa9cKujtkqJ4HbalweDmQ
fY/bgMkbXUIjq4xr51XUNUo0qhewKNazD695guLF54Z7qCePDPiAvP21DVQWL2e/d5F/36+uHXHj
INceB1K16NUf2kyqfcFFbv3tRX3pLN2M8nR1sNnPppV+tvm4M7NuKdHgJp56oZD9ExIZHAbSqrrO
IFIXY1U+BpjPAdIUUcyWRF4QP0v3c/FyBzKukFLzSEx2SUzQUkm64iTZu4HSQWiidPX32UslpaJ+
9pp/d1jcWT2RYHmBmk58uC0dpwxZUMhjlgICUWJ2BIkBeQA8wBYELnF7D9AX0dqaRVN8iUZ4dtAq
LQWWgPqxoKGrnYPzn2PD44TVeZs4a8AqwzPEwLB4DhRLZhxa5lBL20SThXQdVhVl+lv9QzBs5RPV
q1vkJN33bUuK9buNhadnAQIFvIrfjx52twW09CLRad3yG+NLKiQ7aNB64qJdmYBTzpH+m/yiWzM/
x9DNdDWdBuCpQyDylXzAXW/5nfaciHdt2cvIDzJUti3ZDEGbBv6ujI7TO+EnecQYNa3a3yJQ+fmc
G5/YWgIQ6V2kTE9kmr1122NU4Rm1yrOczIUUBCx73ZWZI12b/mOHT4IO/Tr/CQEbvdFHj0e9vloD
qZBV89BVgAXaFU4slMHD3hfkdMtLE8BMJS4O2mqa2slTgzaNig1rt5WRJKcbNkE76JHNFlVtDAXd
ja2ykADulFEzM3J85jj3d0xFWPYdI7PNsEI1mZqiNkc+sXXPbl0eY+xDJQJ65hWw8XJ+FZZZRBYu
KVOaZYu9aoZZ9iEQ52+hfGQ9cp7cufk8N9ngbiQdFU0DFDU0ivpHJyBHRP94UkGMK3y+brn/v8i/
5NQCji+ITMsY5A6ediL7ECmzaRFw7h52jTK8NgAjsQ8VIx3WQ7vZfZTnBbLT1KgQ3ND2f7t1SXq1
F0H/t4vZq/fZWEMcSWHrrOoUDD4plxZXwG2cmRNOL47Fecejoh1fyIqUntJxC0t5Yf6gf3MkY+gV
zib0+E+7RP8GwbRbFr3B1/FDq3bi/Wv9SFBmibn/qNUg61rVSkVZ5uRbeWJwt2scgDP01tocAjSn
4vS60bRPZwNjSMQdVlj4QimaaTKKIqN316PGWGZcmVId7szuYUniy6iCtiRKMI5r6hHQ8feVk5O4
BoyEFK6ZZUhH5yRBrHaQRdk7T8K1qhbTGQuo3DkShQ1Mb423QZODtnN/sey0isi0DLOdciMs2t8t
jxbO9ysRe8Bu0AT69HtC1UtYW/zpsrBpVal1nSfMuFHcFFDPrgJ+xBzoiX3RfW6x4g9uMdwDqJio
TOLSruoGXBRrAOBBKuM1OWpMhhPKdWyQmZ6BLDFBETd/Bn6SuWn0to/Z9qZzqcH56BRuuZJKG8Ci
k5P4dSN2bzCDBhdxurfTcDhL+eXqwh9366vFwi5DWq1MFycQ/hNFcjFa0/QeSL7CEmaHQXraF82y
AkOKqKpr9/nqUUWD8+logrxQg2/F/apQ8wbDPTiNJSNXGnlasyLzX6ufbpGSLY52y65UxJ2e4Ndf
NVQJlny0ETkYp6Nwrplu1QgQlZCbj5nBnad0u0v3H6ZQ2Lg1/o29wL7ZaFH9/SRX9ASHo02zZmWm
okyNkI7llGAmfsz1vYGFEE4QIytDv+Dw4WkAuhyvjw5yQGWwWsC3HhmAx7BIc3zY5HFD+QUOmW0g
xrd/jTMUj+0+dzDGP+A88pJB+AEBU+ATq3uVtDypyBTl4WJ9ohjCEGQQI46zaibfoxHilpTjSwP9
EjE2ZOFxfMclLq3SSzmBShWhC0MchlqRRg4m9lpxkBIfE0uCC/8NBmyj+k8GK+mgzKQSO3GjnQU1
WKJF4UJkn1ZjhXZx7y2GflHq4lOy7nCFUy5oVU7mtlXFHTGS+zj5ojaw5caIbi4DCDJFMVFV0OZf
go9BQ+eqSDAq9ZWn8X2yj2AT0Xk6Log8SNIFCaxvNxP5mPbbxQdmLrO4agA1iu91gib84M0ErWSH
gEtAXpoYv1nP5JdfEnyX5STt+Vbes+uEVPnhHZ2WWbyAROsM4zUBXWWPi9R8THBH4ZMOGn7mkj7B
40at/Rw1jFhFdEc0eggQpvGmyNWwGevqQbH477B4wVXkfzHb3GWBL9XfeLrjtRsz+dQRz9F7Is1m
zripQbe3RG9scQOdV3f2vMF9jA62LPH0iHUXK7Q8428je3i9f8a3e4dcA58KewOsuc6W4deCrC3C
AsxXlR/1pEfZOdKe+W2XXKr/WasqdSfM4D5w611rHb4a/QozlFJB70F74KzUzkWknx666zt69p40
mfVXSwDnEaZa5eUUsyszGl/ArLmZJx3CY3BS4dbhv/iOeYyawOzOgTmnIJBtmEr5/0mPIGhYFxOp
3AlzyY7o8iVrcdMUVW3beAUrzi1XADL5moKTyW7CWXg6hyS1x6m4MoNs2agTda5QORgBCvIRJ72J
0kcYy+MgebXYdBJUNr6fH8VJYvOlcy/j5tVLQkG1J/uLySNrGY6n/mOZV8pnFBOIfNlo2jYcD78d
FkjqpqsJUwZff5ZiOHGFcVMwXWYb3vZBkFJLV6xemWcGhXhQnG1/J+SPnPZmSlluC+grZRE5XlqQ
W4GDuw2md1e1osAyeHAvIt87f5JyxG5O7Kv9SRrWwlE4qxwUQqdkBLgQTaX4jejheGa2mVDUUPys
om3iu2r0nuVVymH8zMjTUtm0QQVp/d5F7xMkQMMJS+WH+EHaRRo0f5zQfwwXRFLFCuwRhxfrxMJD
8tlnbNVq7pMkkhZsJUvFfeQV/SWagT2Bvu1ni3Kykwke+sty7EyijgoKoPnqQ0nvm3wZ16tHQq57
fd5kH6yxAr0TPPdwfYHE26uu23Spdnl+4K0QQNU97SrN1nFQHM7YpRsBKdMOd7uVqEC1jz1oCOBS
hEh6PvqYCguOVzP+3VK1V+iDFHLJHUTqBioMiFHnchEMi4Vxdtcqbui/pq72gPZjUcm8DNV5kWaq
7RL6m6C0a3IMSv2AjjOY2cY58JMANS1MibNkTShb3711Ww8N2mFzEUvezqXHizXtHOvT9Vswse1d
HKxLsEPe+YJA3oVPVfr0AL5zCAVsdjTLoAVR8eGFnK52QysSggOFdq35kksYlZ+epTdV229Fvi0E
7IB31ik9qpOlcuiGMGh+xsIznQR3AQZC+Izg+45quGdk+v1jRTsSZ8hD42wBpPzsa27F7VP6gcw5
BdVJF+1C1j24OQJHeH7yQBBRIsa4+f76mVoLtlxRNvYJ1hUT1rz6WrMc7OXJMSKQZhHueycJoPeg
xSm9DMLXH8XoSnE4aYtmDNT3y6feR34CguJnCuxyC04Fe36bk+DZfoRbn0uigb7QOGc3zKNOmPF6
KrkwGhoeMXrzV/2XeStLGNL7g+OdmyvJOlmumiMWVsYTv8FycLkhDdUj2mQSfoqQXt2qYveK224W
Lcpf71xS1i+X1AwycnE3dg0aGwQRpN4fwDZe8x6DuRiy8uvMAXnFcY1a9NNECbEHHxIo7qAr/2Vb
MFNRvKzwPgn2hlMJcLwPloW52n+8JuctsoIrBTFDH0i3qNppxa0HHOHgiS5cSewK7EaUFdzMYDwx
ascQwvo6wG/RreaNuAyY8X153rxSeK0Avrj2m+CmcexEV0HHJBzN6x2V06myvOSTlON7JfZfKUUK
gTJGYL90DmDJzV63eJNVxadFXmJk6bjiX5hWtgVhA0paXhBeeyX7YZALnofNGpQdSgVxRdvNq1FT
ffveyWMP5mWIG5lh57TkB5qAdZvFu9QeNwkaBCkx7Kzzxs35t4P774Pax/h6esX8KXnyF2o0vGm+
lvIswngSpRtx6W1NV76HAy2jwLAAtZ1hU9lOAHayBgEKU5p1AzEJwTzTUAsu1vNh3JqhbOQ4DWT/
6FSlneCducII3r8xlVU57x+7N4cRWDRVzoHG2COvNC3yBKkq0Ph5lwjgDcgY16SAEMiXTbr4pj+w
g6mQ5jEwFNXjR/JmZmNRCz+XTuH2kR/WDWuoiUgA5t5Axmo3LMWcNDZz/Tz2Qv25Bk5G6JuLI3RN
brH/bo17JtxiIM+1mdLKgJh2xhy25dRyZl3PjOfTpclYOC4xJmYpOYrVGxv3H3iAxoEf5Y8ToKv9
4+SMqDzppf+Q0sVfdKH9kWYQqtYM25PnsqqrupOnrtC3DLGRTYwgmfANA1qWEiuOjULKoEO2Y9rc
OE15AU0L2FBXPR81zPrCO55b1AKAbaO7QSpttTAlHXIhD1qMeYWot5mq3X9nwPEuG1tBS4N1mn+V
LY+VsAT1pj0hXHA65VLSSRMOiUVj0SQY7S7xNyBngejt8DSZpVmBM71fOppnVIg7aMKXRbUc0o1E
zEJTtLjrbqRFihcn0ubVOnwJAay4zZnkPGkDa8QdHEgcXreIpDf8ZxyWB061JbQ9Koty8Gc1sgIe
VSyszQPv/AOlf1KoROPOvIOPthfTIvKCfThy2hKbN4Glz35csXuEAbU12bQ/fERSBdKJ3ueZtsmG
AmcpdBkWwxwJ3mjseZ+C1duLivyZG6UYRG3mqep7PUDNU0i38hg2r4rPujli1zPujKcJ4SALO9g/
Ax/PhL45VKucNkwhrdNxoQJZKlav/7fXAdO4RLuEspSpISzCNZdeftGA4eWY0zr6k9GpWv1xGRZ0
PGJfrt3GKxANwsFsUrqOvomJpNsLxe83bVN2keqkj8VorlhYBsBpmmkIFuiDqQRC38TcxlvG8rJi
ozvHYa0f1smWG0xGGkh7PbW7Sz/XTiZpihFzKAdGrK52VIbrM8AeAAuGIDbbC94c9VaxhMNrjg0c
gG+7cG6phgo49Os1xbzk2feddwEcUB86S/wrlgoFvAB6jo87HtkbHM96rxtw9PO7sxTFiGtLIOiS
P6rBwbGpzORochLXm7hY7T/MsMtDek4Rile/ibPaJaxfNnKjDlRo7t2sxEifKjxSIAcyBDV/8Ve3
T1lzDoGLhDdXBPM4YaqnjHzpprRCoUWxG+MmZjvXVeeMr/0OVj+LGVK/Y+K6p43GCFJSnN2vPB5t
jf4c3tkCsGbNj8n0IG7YXE9AKJbMgNi9Z1lzlEgDbT55xETQur8pReHhtcXK02sNzC/DD8x9WOxv
dgkFh/NqHiGX8ZjtOB0XKl2KG6/eMzLI7Hz3KC0jtnmU3JtgFweDcYOedZ3heFqvGmNkbEJRPOC0
RecbcO/XBEH2zQwG1yebzFlm51ynRt+YM9VCTcxnOD3P3WZT+E2kV9z850LGvSA2FBrDPh244Cym
J1n6JqhM4K10IEMaq/4eZKX8/qSPy+qXIpJcaTiZfukSBcF87BerRlaELA8Qr13GD1UBRYQPzTzN
KxHu0v2xOJCqyx21//c2rOEBt2Av78foS6vhmhh95Vd0URRmHs+OCfwKB2DmTkeaZu3FeBi0M7zD
+elLE/t0KucQ1A7VnK92HHb7K2b4pZQTcyvw8BUPlLMfFEG9R1OADVxcRWKr15fFvd3ngyqKmNMF
ucq/3RvFH9bvtxp1v+sat881zpEdi5jHkNomrawWWCmn4kTVmYuZiU/FtNjIuQP9QfeG8S7kvVof
easVHIq/Kw7Anl3+edxZqhNSdjc6dJAr9ZA0+5cGEX/3V8F8xlKxkz4rb73bSHASdlVkBNwO8wwo
FBWwwfijwYGzV5oezaJBCgLc2FKXyM/tLt4OWdbSPbyuhXFPDgAxGq25A/NODOrze1p3EWErftaZ
ICpQIsfBlMibTZh9bS751hD/onYLfFJ0V9it9znJo3jUIgiUN7sdqiQfm5uK5NG2BEg48t1Dig68
gSlBE7pHEfWcIt7m6ACN04O2PINyBpoIN+5wkJBDCPXbXVX7VcfEIyTOUP0S+Y8j7Y27mvJWtKNT
/sdluC0b/VwYRaU61tTDij7j2EtGIuUQko1gWJYIgPUE2RS+MD+UcpTnPKPt8vMpw1MnEqC1z8AH
ttAnHiKdOOLcUejxm5zm9nSrjI6NB1p47Uqop3yny0B70LviSKYq1EBljLzq8Puax7Z2C4NeywCw
yIFir+s0QaXt9jyy3c72NbfDsmZ7fQlTxycog0XhlwD9HEGBg+DGtUBhH6J8r0RkrLRS8gdbW4hF
fGNlzruESAfiFctmOn/Y17WkZLl/AIPgaLpOVBaRROqElTEfmcSXDL+g5zDl5jr27JfQ3P7JdlUY
9rJdtBj7uZnqLgc4pZkAvJWLLPpPsVq0xs6tBvyY+2PGCgC4rzTQh6DW1kGxvxMNlHb/wygVn18J
A0sjxZKh25R2+gvCrWk4zrlZmlMKMBgfKf3AwaV2Hfzqmlj76arpCsIqvguDGNbXT3QDMlzJFT+A
a61SHtKSgGhcN6QVsQnrpW+VYQqQgYHfQYzO4bBh0A3teJaXLbqSTgLesOBIUQjGRZlx0mSc6JAG
YBV55TNAC1pDSdcj+KmaO6l9+/Cfzu8CIhA362oM37eBRvErPUVJzykGFlE9eOvvExwV7Gg+d5+H
FqoRrPoWPDtlkdQCd5ZzeMYhAFjeuL8s711gsCKqqUC7+/HgcemdBL8k6GIaGy+sF0pHSSDPQwaw
O2rOLA+i2IjIP8ZPMZssKhsQ2SerC5J91GwxbCVXSNGxNPF4gE+ZbBbklVSO1Z5f4cnr8lpztRib
GBLIhoSYtm7lBpHHzfjjCmnxovfaDrNxrHGp3Nfe9fKtz6Fzr9teM7wHJQmhFYivVgaisD8mN7CN
r19N3UD/rHJzPlZGD+MnwBzDdl8vgZPfFqP2M5a7AC/BSUmJtufMyZgH6Y6GgqdEmosfIfW+7zzp
ynnoCGN2lrOZAEjU/loWQpcdI+VaUpViZNDAfh3dPTIvhONyq/g+dNNg9D0tuElos2DmQesFR9z4
Gyq+si2io3YGIVAMExJvXR9vVsA3nuNMiFffh14PO823khs7z8T4r4cXhvqsls/goE/S1LPrCLy9
JZXU4vKtyl0CN3msgeErhc9N3MThXmXZyh6AkGM5bfgoQntWC08zTz6cfVzYl1rbx9/WS3t0651y
8m4iihdBE7yyhJcIZK7Uhpb1HQ34/mLKWCyLCTqHfWtxPyUbWNmyPgsbJCPDOO+bxWeBkwUVeuRN
xL1CZ8pDatGGlyoJ6+NoQsFNnjc6G6tFQyLwm2AW4IK4b6x4f+eKMPufyal1gF9DcbMQr/I5nzHz
u1QYBILfObYsD+Q4ZZa0YBbT3aDF7M38S4EXBpqvcil8jMLRzcc8QW1N26+VO+JakkGIM6xrsoNC
9AU6sRNJeh3tp+1weXCfFa4d4Za/ktU6Cu1W+AFb/4pefKjagXBiLFFNNVPaVwOIXWr4cp+qPQrA
bA3NnThOwkQtxRfxmAJ2UnK4SatUXRj0iK7mTP4rqwtDpd7uaLmQNjQqa30TZ9rH27pZfLDLR/Wz
cAlRsiut5uM0VlRfX2DNVMOq0z5xyACTe7In4FXyVODgbkDQwWZ975pepHgtQxkekdvOpo6OOvHJ
6a1q7hFIjXUDTLcL2tHSVOPJbCynf5m1/pcctlp8rzrrgF+yZjBYW3qKiBdV5BRdxnV6ofpVsJYv
LtV6GE01gDcvpy1lvu9AWkbRhqtLtxVYbtiyIVBUFxJGS2dI+Oua2TrRec3VY9kwVeqA69OQIC4n
G3ZVeXdRq3Brhi/IITPK+LQTPBLaEyCToQXbSt9ViwwLbn/jTqBm2L9TlwtUqP/vGxmEFT81qLec
gLWSXyxdCyRtPKjaHon8WN7ZyZdicyOcWksVfXEWrlxSrQMq3pc2wbqyq9dlQ3uoOPGYUiRyd6sc
GJuPQTeXz2Tn1Hj7toZhVF+d4h8ZRcjUHIcSRHRKyzjaztHhedLaY73rZBw41z5TvkqhvN7iGtfE
kC+y1lXQgtpVP9VAtjFBrBHG5LEkCGLxehCximP1Y27inCNuzxt/KaZ5IVSuCiRyHyhIWy1eO1Av
5j8EF5ynGwJuJsK5RS1yvqg4QScNfMenOCrgWXtEsSrWK2BqquGxY2YonISfxQ1z4U7pCMqt31aa
WXs/OocenHu12G9QuoRoTgzavCFb+hm7rNwtUR6aC48KOTkL0A/RHg2CYU9U8r3KKr1IQXaX9Bwj
WgrLji5URgqTdSFPISGVa8Ed0JLM043g2PQkgtA2oxf0cqPRL2p/WweOV3Olix04HLkkxhSI45Q7
ySosIbopWkEt4yknvGi+czX3Or+5PKalV2r7rE8WQmmm3fig7WUc3V4vcy/f2yrUpIH0H4EwSE9U
0ylvcUdq6H59y+stulOEIkhOYmCfqRvcw0kg432/EUhBv8D4968+b9FpRR3WygNzqGq7tt4AYarP
lWg2Kmno4zBVzwOpGkYOWz2qBgRYyHyHCc0tO4JAXKxSKiGUVNZO+yvDs6GHr2h9frCzHzGSv6RB
FK3XZWDNPgZJ05AEaoM/uYANXKRl5HEwraO4upwERvwETKGA4zYfAkzwufWJ5JtG0SjxUkSqNmhf
LiDAc5VhGqvTa3s69zmYFvxAeJ2LQpptSkrHOfYdWAKaqNlRA+bH6xHH8dA/Xx5SUKDPn1WJtDh3
ow157n5Hl231iT919RjG3QIce1i4JJf+557i1wIIw0rall7ZpcaWcrxvzL+Ck3FSqdXSjC7MmJxx
afwslPE9H108iwN9hgeAJqkwzaAcGK1v0xTW8LiKEJgQfgDJLLA7of5PkAn9bnfcS8Q8ac9mP3TV
MD3+ix63UVOJjHQKd6LSAyonPDQF3NTGS5DsueDbDE3V/zuEWSPcyyaaLsH9QkpllyRnQwL4t+CO
3pJJBujNtdwDJ8a2+bssgGcMBXocT2Vm/G4/lHbJjsIoHOaT3C11P/dXuxIHss5JeYbgzAXAoWOp
JCvlxW3xiMf45SyuNHsBQmlcQWO6AtYGGHSjpnyleq4wIK5QO4iC1GgAlSfgA0jmqSb6gmZdqlap
1OPo4WIInoRw/Eho+ewYtLqIoNlsBWzEFN8d/xWdh+MbqtDU0kQDXywU9KyQHzyycxzXbm30PoDB
s9ry9WolEhWDOgJ6w27atuny+9Sz//RU2BHdOyLx0+c/zKWMOCSMx/HFCx6kugseh7+ilpdEt6+t
ivNiTM8OUe1OAnajx1XJuZXPQh86z1dZmUCm1oMmhxrg1T2yy6GRPhbuEJaa4UuC5jXVvc3UB0Yp
lqFRBEOUW791IebXzKqDfNN49+LUayXHOyjJAIcFfSqF9pd/iooEyGufTNIHmB4oQQPiF45nLeWm
OKx7/tXI+48HkVrKQmqhxjH7eC6JI9BWGe4z+k6/wlOPl2KdYfta5o4BwQ/Ipfsw5pd6BMg1FbsQ
wB+6yUyVayzM0wwnRW4RSLiC9bTm+L2N1Txnf0qoDBP26lgNgoi+jRw0fZYEUNL70iZ4SsVhYhXC
zWgFKzhujdzRmeE69b+nnZwV03GfEY3dOOUSoOedmYK7mGi244zcqH/EArn+jcK2CkGud3qAn+yt
bsxv8yEk1BEcoROCeJCP4z3Ts66oUhDeNZujoPIslF+mbyxglEFRY7I4x7+H2DmdTDblsUUC1ypp
zRgMRRFbZF2Dn2+29QcWsNCNJTJi6ryFJy7nbGnYp9RSLtL5RRL+xD/1YYPTX6gY7Autm0rDrVYP
+Yr98nGwjLuF32U+eMBpoxz+569hCnAusTwA4yNFXViQ0MTKUdFEa7Bot0AaTMckpXU9UfaCKQIK
6iLFfIyy564cOCtFhh+zmc9f2Wyk4cBm3R/RGYryOIMYUaYIWlnZCYmBBHYayKd9AvFhVyNcX505
0zTxEj6MZ5nTIeRerlvHqjVWv7rUpVF8Z1k+6/F9UQBnve+t15h+KC4cS4uhxQFvFN57I5vD+muS
urHZzUtPf24TVMU3CVJpJfLgyMlUBT1sfDfh4es9v7TB+4kmSd6XKZwq+ljgqOf4DoyUbuPGzXAA
8l3p5E1jdPaQlaHXlcP4BxlYpHP+j3wpc3e4DsLapNbP9YOObFMSsjwdXB/LThh2n0y6sbZXxGuZ
0OVjlKJEE4/iFUbbTm+JT/xovLx+K4GcyUrdxOiFjdrdkgaOVAAlf72/h5siwqCC80s+jFmuFpaA
AQqzaerFLKEMNcgCn80K9Od8yDSSDmxq7VVi2TQYGAE2UUZXwTejalzvJbYEhnycTqHDv1qPAIxj
W2BpaNkHEHnF1fawdnUKByfDncHOd7CHnBgoAOyUUynhSEuTHfvlRzD1elox92hY9B5WFFa7Qw4l
3WaHNzONdbs+Wuc8wQXH8lSviIhsQWOdnIIXXNqGP9H/P/KH64y0aO4lAOn77qcwQtLBQiQ/0ASd
9uBIXpeSLs4Sqj/K6bgtJIqkq0nIkLv/5SUnnDCmRp7NFKCML/vx2X50TuK3bb4+Ao5ynw4oAuNA
hIZxlE7Q3SilLagq4qcl03BX4T8dXatG82IP7lET4kZCmfExH7EZGnQGO5vvx52mK6/SztE1SBFP
sxOGVbhwCtReF5ZXCVS5EpZZQ+pNvTjcqD8win3fZyKLWOTdx2qZit5TydYxVhIZLGKeij/v5oPx
CCn9gZPoho3ANBSSWaByTgjdl9j48cMtDlgufNJqtPU+YWCnm5nIZfoB9HFWCa0H9lVSOUpezN6Z
M7VRMDSdFvGam65B14nzXKUH/zrmAt6xgZxdpbUkFpeN0VgkRia5vF+VBHKEwfIbPtOh/mwonFm8
R2VLM/1A0GnkWCOVY9+3RMDt32B3bU0X6ThWondTz6i/7JMcSewTmqFlGEbmPYRRgdmQcYZPHXeh
b/LNCxibC+TFY37v88qddsQe4p9T/ODx5X5ZIORaoFINJqlsslhuLdcfam8fjFazWHFmjS1zH9tk
bRKdE8z1UOmyD5987iCy+n9tyJnDfcHkY/KABoOK2wPow/zPbuBivRMcpKbxnJ7JLN8/mXmCXlOb
qCxFEWlOsvcSzlxWrkJVHGFyRRW9x4jGb6BEVcbO+W9VGbwY/SBuRY91hfqyh7NuiJPlvmNDmz96
kL8iQ0/t6RMjxrlx0Gqq2qbgXqjP7JYHZ0Q2M76AR7enQnIv+10qnElleKKxjkSyLVJV0MG9Mckc
uf5FeePUhPNHv/LZBXU4w5n5HtrJQUIPHx2wi8TDXKmhJqLvD2THVPSRUrAvz1cq26Umo+iTIngW
AGj5rPYyeZoQTv5RcfUHTj94IWwgiJ8DRHcwhmRHBIH575K1v/ZSRqR09oG6tS/lwkzRyFWbki5D
kvQHFDSFZY7NrlT8zpIEvxqPf7bf/wv+wdEB8SaRmwxmQTTcL1iJpjlmPfsKdwREUscc5w8AQKyg
b5fbaJrEdDwO1TXrd2LgIoIHSevt1VZsdtTm50epjGNfVLV+EeqnVXIuPB0/D529DL4e8KBOzMbj
iy5IqySTGc79TmEemGifzdUhyzdgW0s+797fIu83UlHja1FWB8+igGkJ0kgQFPfy65GT+8DWOpeG
U5f39+r+Pi5X+0Ay544mmPHZ4O6nkjJ+6YZc+WIFd33BuleW6VJ7xJpyeYlvFn+4AcjKYBDzda8S
gyVCaTWOm/OFjKchY2/3grD22HHnVMJz/t3flbFysbsiepM5vVupAlLMWTDr4nNuowikkTH/JiuH
PiTekrIKBJSs4kw6Jxgcv20E0u47QwrHQT6qPpmnWE1xzFhGSyBhmEbyhLu4ARWhOHZFOy+Twj35
Gx328L2RhbvQ/g9K/FgA/01WAY2VVyrqcO7HyHPAwEKxkTOU54YGvmV5rnVY8pRjg5ZlZE5c6/AL
L029NlE1Pm8JAfb/YrG1wqhClzt6FY2g74r1H8cx6bgO0jdGSCwNPeWmcXpHj5y28e86pF0RW/MH
7TzYZG5wRJ4cm8Db+/eRWV745EhtiXTjI871978nwSbIfKJ70yuMOW0VMI519S5AodlsH8CCIIod
nXdWCTxms8TT2O1ghsxlZSSg9YKHUVOQR0w8eG0vhpfGMHjww53pXarj+JjlyudIUsMlYBToZwQZ
Lu2m6+8nwDl6/8YLCOdWhhn2mQirSvZ13g3h7ViICWJLtOvAvBiTHWi5MUSXJxhnFJyaSrZVpL/p
eS6MT1WoigDy1Y2+nnsBP5yO5XsLP1mXVv/H4v/UuK2BWyYwcksQa0Hd+Je2jyRbrSXKrla5zJEM
Mi6Fe77WHqv63rZMD2iUMZ0w9fxjLYPQB6O3rv0loqmS00o3octjN7V8lrs04RTM9b+EFKMi2E2/
yGBqGmNTWmwb4fnBh9xsSzWUlENsCSviCBBAW1hokBffYfPqz+Iik1Rilru37kkVXoUEKsNL+y1A
RndqDlJsCn7qC7labn9/0iDLWFc0r+yyhA0gvz/1fzKxp7Mm14eRaDLsI23ac6sBBOqNIc+QqzMW
YsZ20Zxb4XdDjXoMBpY32E9wtPWHiIJVYgNLft73NcTIdYU4NuyV8QJE0otZQU6t6pr9TAw8Wds8
hIKpM7Xlqip+BHxYwpAfby1409TdGCJP14M7NFxq/kys188yXhDzEVZbvkU6BZBxIs2SYVPUT6Xz
+Rszza4+y7hdzduIUJsWrP2uuq0juxbbjfzA5+VMQsUaJBkCHMBBlSI8bWQAibPNOFwoO3qFf27f
gBmX8YbPlw45FJ0iBjbG2WzVJB/SzPlqunozwOZj7lmN1P3pg28xmqA+dW2YZIHe0fAwOS80OH7S
IPjbrTdadlCwUysq5xB/BMs8qERIIthwn4aSIIyAbb7IY1I1cnNj0mTGqb4PaNW6vWsjYDAcAaN6
PjOQH3YgWddGTtVQv84q2TmmAfB/CQCxY39t/K/fAdu51epJ8VO7dFbyCUod90ggDyXjg71R3KUL
CRNu96FWck5A8sCViXMut7fqL2o4E80HD2+yWOewim1kHxsgQoHzo+5yeCzyv40WeODxuRN0pdpc
KINhjSg4jr+ImUDDw1D+ZbxjHT6IS0ZlOZaXwH56TpBWsyGfyM02dYtJ2/Tc9wkygvYY7XAi/bCb
UzKEyt+RXrfy054Hw14fk3GQw4lsJlZ92houvc2U67aHBD6BDqBOkv85QIF9goZER+ANT7IBADsR
N0JwBe78KjxAWLrMAl+WQcc/T2H5rQMlvcL3xEb1w1vyFmzot9GeGTCwpFN/bkXpoHASnlNIjDQG
sYn02A1NazH++AbEWHYHMzf6GJ3+uhZx42KeWSpR8cvcbtZjoei1oIuMX+Nq6MLC+3TwN8uLjUx6
auIqujHh08a4rEVRuZ5fBOmZnnonuzEIai1Mqwld21Q86KVaTIm0Yih+XVeUgTeM0f+SNNwZeAT1
raq4iFFDO8tCeiKl6/zVdeVSyECrryTAuRUR+iDWCAVjBNUlHCC7N9bWf5aU73b4B9PPTtCk5AlE
2t81Xc/O9u15Sggl3niHjPjwx8ykHH7DbnPrJrZ9m1pIf6C6jDKA2CpRB/r17SXGszqs5B7fwGA2
8YUVfL/tWwguzT3wCxZQki2FVo8DFTFsn407cji3Ej9EXsUjWRLYV5AdjUKRq0tWeoP5r6VkWEe5
ZQLgVy3SC0yRHSPwpoir9IHq7d2jvVXQTcE5kDmMAz3tdRAWWcIE8H+gsn9xy3wZv0kztmunxGzL
aUlyGk0Nvmq/QD7kg1tv/syxFvD9dpCgEgqZsQEhoS/ZdXrwtAYZ0g1QefoAoI+oDmT/wmG8bI72
Sd2I2SUyAkZ2yZbxoZEucXBV/pj0CjSFdMrGyGhCGDP4X3zbcXUyhP/hD0qgxrIjqdODSkkZJ/R1
a7AqRghrStBbiqBkynLD74g5CFnZFYATUD5bp3dZUXaUEXKUNH7QwgO0ZuP3e4y/EUJ5Lu4kph9J
8B/uBDM5q69Mb19zjddXNOSzTA394fx4tEx7aL80YGq8Sqr5DikIlh2MYkg0pyTgNQKVkkZVlRzh
VkNOyo0mTxzGAiSbQkVoBEe0K2nBf+qbdAxAqwdat4vXq590E5msV98rAe08pnuilMCCaKQ00W+m
I5KvBFRAX0K3UvpzDhXuXwiAveHdpEVCbVF24lHqTg7OkyOQwI51wshlv6RYW+QSYdSdP9ouBVgM
VwxLvFlqcZGJowaaeczp5UnTH8YOEA6n0jWTmppq5p/T0pQn5fsOhlpOwWMnmBfoqpoPjV6xaGOA
1w/OLTnCufg3ntQ3OM68pRYnK0k//MAnZq7fVRUiyBs1KcXI3lUp68n3CCBOPMjiadKiCaTxsYN+
aXe6+muuCk1u5f1NE0ppdGx+IaYen4COyLsb66DgGhEsj9aBKaoO+u1bafCcvK8T1AKR9JXhYBn+
MQ2INfe84TYlOeeKZFVPxYIXPZOWCVYUa5nIgt3ZlHe5wKSQdk6NSGgFXTPTDuZkdTnxc440B6cK
vuCQ/pxZOpFcgim7DlyeppwkOVFHqb6b440hr4G0VFOuWp2wswFnLHuJHfvg92RgKTr7o5e0+Ixe
vdBqu7PS2lv2N+OzU5Xy2NDbXxnxRO+mU4EpbEHsSX4LcN8Kzad7vUJ7HD5Ke9FVey14RyDqt6N4
z8fICz2ezZrQnGC3AzU3DPqK7Nv5E/lS46ZfRp4e0Ss9luCFYaBfhYkHiKdxIs4/07xlvRZyQq+h
XMUC4v7XRupuSAgERk1HW30xmHG6uUqB4U8DAevNeFwrtfgJW1aZJrZxUHE4S+KgH83wAwdRYYZw
TvqVZ4OYt9UYKHBm7rXncp860rxKJ27H/qhlW6rO2cI7h+M6UQuF7qtKzQtg+hG0rgrl02+sBsjD
5aCTvXfTGzhDlVILqrx80ZmAbZ3iNbllqf+Vt0AH9XEHj7i88FxmVTTq3/hFO3+8NF0NF/lKLmIy
yoEbjeNcLvNmGz6Rfgy2usD48lWdXUHgvBE8HYgJEvYLuy7aHXKkWMa28SnSVcL9LShMRnfyl7Fv
h2FQHM6vbBJmt28ei8PVVceItJXy4Y3o3JYwphajquo7zj0RsDNt/go0PlN6KWIpUm3eE9cqQYce
71ag0yqrSXsHcUeelVhQVkOSEa12b9SdGlVNA839Gcui3CGSYMvVgOs1Eh1bZatxty7fSS9j0Bom
KZyPKXpEqgQab+J13/BFluKKRDrFBsx5qZ7nGen7vOG6XgCdhCxCyTSLnytGfP6gdcbp9FFsUqpf
JDtXEs6PdGGC+b5plX6C74zICx1eXtim8ViCmX+HW0poudvj5Reo1Ugl+yBw1U55rVQSm5aAdvYB
yKXyzcCArXIsIYVvZmhWbBfjSrX+An2qQzvFGCYJbfovqbbL0MCDNXeJEuKsRt7WH1FAY4B6ZLF8
Mj1y6hVpuMHojnoijckcTeKRGYI9uSefFLXxuBu3uhVxTgbpXKzjz61XA83qCIQ8sdDk/X4O4NF8
uanVprRghYJwwGbCSyNXV75MRSGKgqnHV4pw0P+Kkmaf6DzhC9SAK7OVPjo2STaJyyzt1t8gmvTx
Q4o50e3hAw88Qg8hYw87/W/DwO5in7P8MS1lB7HfAo5dLHqjDdmXtk6rE02rja+15PdpZW2ZNKrX
J8W5sFnUOONvOpF2eZWown4128x4Jwm3t1ON9afT6ZF0RzEmsrcnTYlh9UP6KfYJAcg4OHedTZaV
eBDtKAupMBwBwaSR1wAyeHMQVJu+ZHVAmRaLp6ft9/r+McLLBMyjWVOkFkPukJ4UurDJrf0uZ0E3
z17hyuRQ38Ch55zkaL3VaGZIrHOsvMvtWOirLed0I4bt9qAOp5IInitg1Fm/0/UIvM1AN9QS4ah/
VwMEHpXm4OjwcPeWYpmA8euQ8a9E0JeDGR7p1EygnLCnX9Yf0hnn3UXM4UFJHknp4Y5S258lqc+O
7XiagFqaVEBkomrtKSYUCIY1/07it6QUxw0/4C1coZygqHX8sCXE9bYXcnjsxwB+Ym3cpkMH+xIT
512SMEc02vW7xCTrdn7Zyajp6a9TmLdNQ1hbaOGc84xHQDByGa3961HFZXv7zo62/tSOLy632EeD
JB9lRnji4paB9rhydsaNu7BJ0OiIQw/Txith3Andr0VUKBOEVa4aESXcJADzWw8ffv5xXapMNp46
o0jaJynzMiIXny+OVouRkrJ+Z5IoCgg3OK/+75JzPjHb1v8n5mqKNC8/+ddxbnS//ONwoxLy4dgM
5ZomxTHpGBLtbzhfK7jX8uEGmteafqRJqdtsXX+sE7e4Bz873OY74sMNzGVc0jtlvUXMzSWgBoeA
Zz4Czz6jjcCJF/4Xs6UcspN3jszvUmI/oFP4QYBaVUZQMOOAgNqTgkeNTPoZEA6WmT7iidVV8GeR
mNkt+5qnoL1Uqos61ISRKToawexwrzTBJAaE6os+5O4lalwAiT6qxDmhWh54Hw8YDHPaotBaS4qi
GSjbndDznxDB7X3vD20cIi9FP9PlQvRJ8tKvI4KZM++3dlyiZc3yxQMVzD/7TWGJxTG3pdt2Bq8A
wa0XZma1Xdbz56n8YeKNY4peuU9ZQ1qG9CstCRFwaoA149QqapK6iVjcpOwafQniqeCwK2HX+76g
4+19CHZVSzG6/MgnmjrqwBLUvYwQu8OoBB96CPjYSCw5N1oNwrWmtdJhQSASOVMBDYnmJAXTQz2M
DxKAc8kw73F5pHybpn1uSeGPMMFrkMN4v5Ikm5qeEs13Aa84GMhvYapi38OuMT0Bn60HubLw96Zk
clOnnfAE7BkKykxUKhvSg+61LxKnR9BiLFCuD6Rsi6eB/tzB00/1Br1Pdrse6B0C3d+WPufygTjU
UvGkUzU4nG2mhPs0aVmU23cDTf4atjry2ivKzuP96Fd7s5Iw2PPB3ZnGUIU6XI8tuRV+ACx0RaAn
grIfbxDf9SK45bJ1bfI2RhnO5fpTo416MEst5HPN7dap1+nqT3Ot0P4zR6XMveopRciruCRVKvFd
0VnZeCazNZ0AEJGubMtFIvqGdtZ/OLkV6fXA2O2eaJIsktOXmWUZO0yXM0IU2Dc9oO2uCirI1ujI
WPjNCRE2nB1dq/9TAHzOKPR2M9uYKMBQ/O1wg2e+HGGxXDPtVxMqDKm7kBHgV26hxyddyQro5zMK
wg/6//k7n43TCWW3lbGNtFR7QmLkBUrE7aaIybyF3zoVt2pEi6miUk5I/JUgSCVCJnsThGypmaax
NDxsuU39+iQGKGOXeobN8XDBwf6n7oMKUM7B7fdJpxGI/ULNcPFmdVlsC3sO0XAUs6Jkg+MNjvr9
V7iV0elK9c/VpqqScv+g9IbP8qqPDneYTaSKM4UiLtyfnw1l2CHtALRzX62g6TPXD9bvK7sR+bve
rBngQE2Ypbf8WoljyYvGd2XqYewtLVePgL1akAvO+rYUY7l8BPF//kZHRG8OIeru0cLyU6hpcwWq
Jl8NedNO6UEkYurQhdib7TL1lyyK7LCb46erlBO4l7tOaZdwqQcl0dTU9ZE8ZCgOfzaOj7wnx24o
vrH3jpwCFc4ZtlPsOUeZ7mF8LbcMWfrGu3FJGAJP5D2NS7i18+JqZj6wjBhFXUXaKl3uLA5LIyUb
Am7WaC8YzzZjQhkJiTabf132+qNz6uA9Z5hnRpjHSnkc1SK5yLnIqOtyo2P56bW0ThTv+nU7o/Pu
54Q+SWwcNJh7qyOh8norBpdyLL5L3f4mzKwJeoijiRNMjtXQ2/vuhig8IP0QFA1SnAejWO2RFMSM
aZVR4hYzDmreIcaWoAPJrocWtUOwAfZsmKRLx1vTfceTGaG7WtPckctvS9mEXAmNa0/dn20Vyx6N
ZqWoahwKYWeEmHki0UulQ1+hDDyGBgdYR+61P+umUNWvSCPNUGT1Xz8iurVyN8tyBOx5uV0jtXiU
x5xrfU68dYUcuR0UtJsMBBkd/I0XrijVoqyTq3IgJx/4tvBOmm0s3kYDyw73qxiziDpDy3u2lGW8
I+ZjyE76EqA8g4k8j0JLCRhAbX8jS479O8OZAWF1AuAaqbO9b6CCRo5kupwxACc/P9VfRsIl6gOi
HnSLyOioOR+JxFI9lEXrjHoc2kJjO6qzh/m1yZmIN/+s5TovNOr/3FT/l3zbISkXL/H5qPM3BsZh
RpR/31iIRgKhPcrE00bXUf3p5b+y0okPNcDZdNH1XaqYjZFKYmRHTM6KPHL+ucfVZZ7v9Ytc0tB4
pDGnsrn0+ISDX/QfWuKWEik2yhVdqsaRVuM1d7efoiyDlMK0qo2KLpP5Jd+w91lg93RNEMznB0ne
0R7AHHjBIEwxc4jELUabQbmt7i6u8DD+JMEqG2rQL62Hn2+zTk/xEf9CS8ZzqwoAFW5IeoMsnAw+
WL1kZsc9SRc1RoRXulKJ3yiVU3hB+URe+EdO11xzv49RB+y01b1FpPjYyp/7ceUO2UGNZmXhvaVU
usXOfJYys42jkd5eyce67zi4qT2hFK0XGO8pdcnQfUgCBVTVed0Tvp7hOi8Rk5HrbQ1sKcnxSgMP
63dFosLt1G9huI02EBEYecMyJ/XlmTR/tAc9Yav3jc4VxuVlZXnlv7v3LjkQ9LOUWX0ouf9gL9/G
NWVuMY01VucRnfm8v8/iExs0Y+t/YtRbZPGjg8qmMliil2KgWV8R3vkVgsXlhdrpyMumAed/09+K
dZFPjDuHOFa0HgqPAXFNMuhUZVkkPlcC2Sg+42KcBZ1TKKfORlJXQ0pmz7M6LzBNGy1BAP9ddthN
aa696SvUAhy4OWZkjD7OglxkwhLGuhuL9bFwi8mVCJWqUi9N7kWndVnqX17zXLtq4J+0fAxtHoLK
U6m3d6kVG2He9CvNgYFnpPZ2TF9Au/5fUtfZeNeuoGMTSzI4h9S6Tco84uCRFCjo0jOGk9OVQZZm
61TtW4yFZLO5HY4wGCYjo5iAZqJnGMNx83U+ZVndgPMdI9q21UyK0VN3u7ttFD7lGBWrrxr9xwg6
0JSeem2RtNWEvsbzqEWe6v5wOmg2XXvwQyxkk80P1fPMRnDEk3KfIfighKdGtXGsYbqqlIh5sW0l
CaaaTX7ksmi1ShNBvppqBaMegDb40kgs7SBMKe6QoK85WDUXmZWzboTYnctwJNpQjF/M+ncaVODz
ScwTdpgoIqjHPaGtAs9y/liSDYVoCWr8ca16N/XaYksW9yDNS7iA7gQAhEFeJZLQEjYWvofiVV4o
m6y2W4MLWTQ8K3vzF3DskyFj9y+HvqT0anqGBHA4N/fKkTzKGRssHtwVn8VvVmPOl0bDlC9XRufh
0zbB+5Zc+7rJbXeqofLb/oO76E575javNLmDpYBOFWmnQKk1DroyIi62UXfi0tbhmmGmuV6kbgiu
Nj5RVjivmIyg+Kgz67tl6R7EMC9Qyn+cApXOGFLpbpqEPoPjeSt912S9yCEhZSeHgPxDvG1Xkdz3
aRdBKA8fymJc6KJFrx6kcdqIoq0/tUTCy8YIJcmtaV+7FvseXDHR6/80NAGs7cU/t3NTwyCu33PA
jXHeeuPi66mbBzgWbESnIrQtdO4Gz8xdUGK9t5qh+wJprrfXo87aVAYWkOQ8QtZ12S8yTI8tJi4H
ZWWrY5f/+q4upSADO/t6u0AlJBy84ayZQ6SKtSc9sPCSnLFPCb7LUTU7UhYsv/PW4Kay9k3JoO0a
H4hl59fzyf4cn0cRZfFcP6Iqdbo7bCjscP2WXzvHg6rRRd52v717O4qHG8IW0NX98OKp9Ls8adES
XyNpTNWMplkJrK/vkmjr9uUngUGsXexOVRivzn5wnl/UAvEZzEluBVqxVWAIUz7bDEgGo+cHjOGt
V2CcAHwpY1tMtiFP1YaucYBQAPQ6r0+Chq9aCOMYav0lkLOL7fp3rBCe8PdMsy5Lb8iU4k3whgz2
X+MlrAKfbhL2tIufexJ46qe8b+oixSClUmx8Vh2iVnTAuMJsp9ojhMYpkz11d9oZ4ck0yrWHura5
DlrL89tVSYGJqgo+M59YcgoIalv7nLiFUQ+7Ikf00GStrZP6toeok0vXg0mTomyLZ9D48KGYxkZq
I9KzHMxJ0fbaV8/4PIe/pYzYMUUQ482ZUl2rUhI1mWFdCsNpWYz33kX9Qu06XVDPSukgY3qrl/Ha
biuBBkqPBHYStKnYHhXKJwgsc9qTbvD2h9hNXZEZK4d8q4Evxljg6TpjTmx1u/qBT5f10eD5+AYm
iGwZtq0COlctHArMJDo94QXQmF6mt50dA+8VcEc85GHQgnQIsrSSisQUXJNLV7slBU/Y5q3VjJBy
mihbu+QFE6ntnjjqCUT7ivcQWQX9HQVBjxhKEt25FfocB9m6osWkSklDKNeWdwEY8Ki9ev6tNDmL
+XxVUHByrhEHFDQX2uVJC5mj8EPmvHuH2E5qkSWgUlcJlNYgLiprmcQxFnfGsu5aNtw9QiL3GYBw
HMeuseRW3ptHOx7lX1CSd2mP9dX8CyrXUGRHKd9rKXphB8Cln5CpLcPWN3ytgk9zapN/TWF7uQOs
/W57IVwQQtmKz82ViWujLGK2jkHNmgmgpyQeFElyHFVLojbEiU1iCGkg/+m1YrIY4Mr5UohQayeb
HLddl01fJprIDumjrdn++NnzARYFOUFZ9DrgliQVm7kaCl+H7onKDPX6u4cchwVIJ+bHnEW+6eGN
TH2S7/aQ5wNzJdjCnIHRbOZ5fdw95IY5rn6Sp/d80eThAyJA13eYQeGttqPKx//eAQoRG6jWWXG9
BviV7hnvyNkpI4OMMY7XUd/5K7DCLKXbWpWIAgL8zTzVy56zZYYCrwLsGbjLak8toin12+xt6D/6
ODzJEoscWQEvSdXCQmKdN6UjPtNDBG2TkRPJiI59ah62V/rej5JG/vZezV1tBr5WMq3BGe7O8/AO
h++za5J7ZDsi22Lk04wKJ6TKvp5036j0zARvoWiyZzDDsBf+iz2KRA+82iZfFfb01NpSc73MkrNp
g+aXwduOv1jj9OhJgCcxzu1rtQE7ExFhq6GjBugSgSC+3n4qmwhmPtBoucR+tbYu93WEkFFKiyLL
efGzgoe2yToPhE6TIn50o8vrLp0xpYzdqtlwtEea7c1+L/6Akjwv0I2A9PpOLc9rLCOGGP4sjOkG
CxheljwyeSsjsKKlcyrtY8DWDXE98XIAo/oiDIbfeSqW6h0L22RY1/FGg0CtGCgBID/wXOjwAj7N
ud2DPzHTBsvHNrf0EK7r+8qN6sMhwoecBvocoW4o4nefaAjYdshRyYRn99rPJLs3z4XTFhtvVAQP
ntfH5e1zJmvZoy1/0Uh1w00dWZhmmWWupLJk4C10FjlSVYT9JFk7FFHRftJ45Ggg9I0UnhItRZFZ
TiReKgxkhxOrsWvd1J/FFUeMpiGh4ICtUnk8GwWRRCtWCbxvDyBnz/u9Mu04OTp7zePKOl3F4n6O
7FHEAk8+eThcp4G4D68AsZ+8FJHCcpbYG/Xp6/30NS5ectTRCiSZHEZ2IMIuMNjQ6Mm2O/yGPQYO
cXlUh0g/YSzcOjSHrNtFu/8GwDu99N085U8uBjMoKhUAy2jB+9SfsTB3lcJzIMS/OuJxzT0qAjjY
wge67ipYKnAXLWBT5T7Ckdz6rYl6I5n5S3WfZdBtHVwwgjmu8UuvXIWk/1kvMC9Sr5BlV8US0d5+
kE8+xV1xFc0Kae8anOOgFK18DoZ7MR76/0suTfzlDSY59zfT4QgTN/5RqOg7rz2KOU96lh7vbINg
DZism+zWTHcIv1jNfPe2JJzU907COSRHQaX6WP83VBkCKm/JNDmmquiqthDxtFOddHtRklQMDCHx
lVusaZcH61NCupc9MapjV4Sdj4m0TCyhrZoy3/i5XvJ1/wFs3PUKFzkpI1E4MyHleDBCDA+95ojA
CelQrtG8mCxkWn2osaYryQ+5G65655O7q9swd7JmZZV8jT2BUXXz8QaLphUGVckre1AFotcqQpB2
AotpFCZU0zK8UygoAWoahMTmiJE2YZN3rVeAOwBgwytE3xOlKPN20BXzO1tLqUzwVcp5hazN6psJ
hIKbm1doV38diPJ3cNQJO7QRHQsinsLgsHni3s/b6dYHzUphechGvA0JrdWz1o/flA5Scbg068bO
N8XyzzeSbRvIti+rQ97OyiS9F2SNHJCHc+dPLJ7DcMw8kqYf4/0pOW8NbvYni/4ZRpKZUQHYdR+v
cW5tzrcAGpABQa9p0TUike0+nbp310zobDxqCIugre0u3cSYoqoSA9aA/6MSZWvRXaeK0xm5hRIt
rM4Vw+xkTK5D09pzVMb12zcfzsBuzHfvHEo54tMeEXebQ2tLBGPfPzEPmzmrjqFpPyWYHs9W1gH1
AJrzMQ+QtA76Y5/U9QcwQ/47O7NSZ0wXYObZ1j6oj02nuMo3UwjoLJtL+50qH5J2HczrkP4w3/SW
slqjWzKKfHDtrY1HaU0HWEvu8ODi6YH55QhunRqJV4ixHjDWPXacZsMwoD/qQpiJ8JY6GAynohyj
pL38IYzdg6u7oLIznpi77dA/R7YuuLoUsUhsi3LTVUrqZAADfOHnDqBY0GqsSJwfaK4ayXZKNt1t
pRYNFS5ynSliYtPgofxa5Lm7216V32oYB79gK2mq1Bb5kEq50wZdjQwPrhufFke76PnMj4JA3ww5
9/hiiypdXB7rPMwXT73drv+LuS17vvS2L2Qew1ONjJ7k5w5EKRL5X9swyOVAIk1RmCUvU88zqgPK
JhY8j9MifKRiX6BHkvAKJ91HJ6soZg8ufxcr9VD8yE08IoeW/Wr81J/5pHAAsMhi9NGoKwKyADOL
2F/VrKIbx2lYarXFKSolc6NUKtEoZinf+8rzWmvHxN0e07oKrjgppdUUis68lCDFBdLK6GTi1PVh
iAr0Dj6psSXPK3kT0nch5CEhSB3R3mpIZ6O9L7+zLyulOM8xIdPYo5HLcbfUmlT7jDxktZYAie8/
iWW9ofvNAKegvULsb8j6j8SUY2rdN4aKV2zsokQegQJHrQDTHHcOetgYFKk2piEbNuyLTu5Z3F2M
DuG/5a9aB/zoUuNy8Xq9q+qnNuE/2w0tR8WDO+Pwt6FrfwnmB1QKbHog0n9CGmtU0xPewBQ0EgcH
eiFgcJ8SsnF8s2N0ZjKg1BVMgX+cm9UOdVUx5M3SVlT6UJjCn/ydcBpLLNooeIUM7fqcGD6vfz/J
dplOdLk4Qadqln55ajofSWcczB4Voq/nRKHa6E0UpJrfMhMJWYv0X5tHdsIILt9Y6V7j9qmJcKWL
avNW0cl5EmicUFa0+L0nnMWwY+WBZSkwrDGf4a/uFx5goXF42C+pj4GHYRIzDM43evlHHHM8+CBN
RLjT4B/8NR4lylJwKFiCKYJTZ272Mjqob6s60r5kyNJ1C9NsJfS/lApxb2D7U3dJxN7yjc8STmX7
KyKCILsjfXjnMOYbncQ1JsHnBsmKJ6I9J8a4vVWIdxI/OljIsAoEAVUzyZc0eMm9mETCwsMXZYeT
4VJEg0cJf6T7Vw/SpUawC26ASyPUE7hmh47MEc2puu3XfEkU5RFC4IURlpMigerO0U9ldDDPG4PI
nmJHHIMT1++A8nrh9A1jtik0T4cCgOSv5bGDwTOxh2U1Wy8K5SsgipVWnsBamGk7Ixmzvdi9D0bo
1/KfEozujST9B+wZHfjrpcxKo7ao2xcMkeETWj34707uPy005JriB3t8QQkp40t+b4tt+5lKgiYR
A/utyodsMBUSxw+h2W9zqqlqHSxS7aQVB5PkJ1UJKhIJR37vhu2ynFi4lsoP8LbD28DGvetqnIKl
dFiZRZPpgHmskDeCruZWiFc2dfhXvnSTiT4351L7xYNKwYrjsvri9JhyWSEamtrU9POXaZbccbbD
WBrai7R61/M3hW3vEUPKsEu7NHBxq8yMgmg070y3yNb0pV0UQSfHb+FJsdPksEenLf5l6B2UQoyS
IWK56odO7WNd6HNS1neh00t5bjdvg7Mf5pmVimTSWV9dLdONJ3sGXxXR9h57wGqupzim2z+VL3Ye
t+cYNAuv+2T/u5T353hCRshok/yoX/Zug8wIzukoVw/VpKXlfEBU0rkiyzo7yFAk/2M2Ckc9Meji
lbzrYa2hjHtllirivuDjce4xvkeVI+ret/pTdnDWdX+/84mMbGxTFwfqUxN5zF57EQpfpn+e65T6
IH0VAY2s4kyX75cny/c5/mbSBwsEtg/PU3qwDbhxc0dtboJS5G5SG9Sz67S7GXpb5iGSA7LeT96U
8oqCSmndmhBeSIUv+Y0UTRY9cgE9sN8O6VCUGTnNRh3HaIAY7deNkbNDqhMOJimi+0F0FWiAhrYq
qnF9khvG5TgSg8W6bLrzexu7BNqJjzc7YvWwb6IjZ3RVfmnxiuwS645UPiOHthTuzFCf5iE2gRjp
ZIghzz4xO9nNcKRrmkPye52whacV4rcC+cUOnhL6JH6SBRmElwBk71c8uVpEbagOiHaE4Zl9nH9z
UmUiEfcWj0w1NZWX5vnMOzUdCKO/zv/WOM+mgIWOX53sPFej4PujpQ5AJiPpKuzaFh87pMG+4oG+
EUe8fHqTa++JBCMEJGI4l55i1DjWHby69WfwLkMMyZcEPu3O9cgE2LGtGQlK/k4LCHENf35+sXcv
kjWcAzFK9nJRXqjlGV9QEPdp9pTS5z2uxkSuY3itaahXvVGGVxpZe0LBCs+Xt7fr1xGo0apgqfqW
LFYBkwmoqzWP6mmaIyaI1lqDdGapDvkc7XIDBUpMWb6/ashgFGq/i9RqVYJoV52SWo/dx76aLGQE
MyniTgGNilcZs8U00MHTAz5EmkoB9dXhG6daEucAanHFLDJG+U2GZwS9Gn3sFhzIDEnC7BGjx8CV
+P8bQxFSvV6rsqJI9gG4WD8nYCh8zi5J4JhsJjmF9oZJkIlPWucVzp1J4XbLa2RvomsGATjFicAc
+4EcsxAH6GK/xcZFWAvj8fuoHryaw+4/BmmeeSKaMfN3maHZ4L48P3D8pM876j3AEAH27Q0aPyfx
PaER8HjAlaZiydFfJpkwIuc1hVN/HvP3e3vI1a2FXi5fCB1ohzzhuTG9oeXhDZJlRrTE2ZchefhR
v7OO0UtP5p1BhBiBX5VzUQuLQQbGxaKjGKuEAXTYKXqjKzbsnotCzFz23hABa8Vf03Q2lpl3nnWo
QRFTCg52Hp+dxDNgy0uFxSCx5pGd+wgiW/Qeom1l23a66qPQzdaJiWKBGcJDdtViHRuFTgVrtO6r
ceIgnXwUtc9Zpk8quOnSjPOJ9/3D8Cmjn8wF/7WA6UM8H9Q9InL4kjFxLA/4eJPSs9KUxuK6JlXU
gBXX2N4H3fndQIlgflvJva9qGFEj0ZSB5t/VoaFkIcIqhfx09Y/xyjzJSwcR5gPXj5MZRRjuYTwg
sgUUhXIOpJ5xm0b43DiR6F/xQfzD519k09xRrTj94w7La1n9Nc+Sr/2kFuFC5wT/0ZjEvbU+wSlf
9L2j10dSd0bOj00B1B6CqFzxiGDfuiBqTGiajjUwcAjqBjGy4VRjdB26MmdMII7OE8286qcBpclw
hRxkFbmC1DQlS2QL9MqBucKMH31LikiCEDaiyIiFB42O7Ip4PfTYkzNvfdc/60cMSxhULrZntaYg
VEN+xq/o0pl257axqrZAxaClCnbkjwjYPhq16iIdMpjlidTlFd8E5fJsksb+tOK+DZ8+hyptSwLz
AW+hwe86t0YK7q/q1qw4AiRmzWX1mpnFZ6yAKO82yMKmIgYvJUQ7F5g3hZWmU1JA7vl9p7T93TYl
kJT9zLqkmigqX3zmKd5PyvRU1DSUN+C+W0AJN2lOrJypjwrIeD4RqzL/vjOoHfbkJjCUxpwP2t94
5mMLHcLmsGj/MBociFI5g5YKc4sCRn4zmZhw0mKNKckGk3F/SVRR5hQwfyNri8fKCPgEd+hZk94o
4gYqVtpSeFS73vj2RAle98iAlvjJkdGOLhuRfqTSEzcFSLca/C2q9lr/DmfNSLKN58jLqDoWROGD
ACBbLFINmeWx6bEGqY1x7aYfWQQzY5d+RJmumlSGJY3JHJaDyzWTiSR9riLkfxMTbuZphz4fkjOA
Once5YuN7+6hexOeQa4dKfhNIdzT1Du0SnbigmXGB5gp2HC6n/N6N2RRf5UzZkB/ECnUmi58nHx2
3Kg92S3SgOxJoPQ67MinpLQgNBqGNj3L+eZK6vohWlyQNY1dUpG3fM7p/CN25p47Yb7vQpBkGI8b
nYD4sLKcywMi+1SdQ7lRkgOagSLwfGLMRkXk1gsKMPtDBgWYbZnWcT4VEMU8wPglQNrM1bOlTiS8
5ymNJbq2wTZuI5xt1jVyMTMb+yxdy+rIp2ZS9c+a2auqPHibdQeVsnky3fFHydP/9cIB1LYGC5CA
YWCYlpfO5gtxD7+HgD0m/my8jGdcfi2bR8qpQ93YiTEz4DVwvbF0L3P+rmpQ8AVrBucmMwiVnAQ5
BtcPt1TY9xInkBGX92Es7MuoUND0Lmj9YPWlNR7uNvvXwX0pX34VMkGh8mT4mxTS5NvwhlGoBHHV
fzCKKquMnil0tgRIqzGwoZvUmjsVeuMrK2kquSMDD2E8Kf40t5Ri9uTbUx3C2wn2fbRIOqhOFLfD
+TgarddOUAoLA9UIsWBq8+GcjfFGsAy0XjZFNWH6deq7CtfITO4WomsxlNWXVlH4fwayGi6IalBc
hDhr5KYiCScBHKtcTFzzYN3C1uoPzc7QYQFaEN/LaMthohbZi+xUIv9qnDwS/vdapL06vKh+J5Oy
lkBtOEkIneT7d574Ey/eur8uk1pO1qju3LVf2HUaOoDzk7YoP8crE/aVziSRQLp70jTZjE44FkeS
P4ftE7uUxNPcjco/ZaTTl59ToKEoQKtPSBNbkPEpE+/0WEh3K8pHP/PpZeuJ3VyqFj1QZd7yFj/h
73wLV1AsESmla8zEfNQZ2g6JbStr+5MNrZ+WUV2c4fvvvsVVv1//0aO3LYDt8rwfQ5ImIufJe968
/fitryZvGKgHOOvBgD5xFPslM/QYXGte4199+AKS10j4E1pnBnPcK9WtOx5cGzX90NMONma1CtSO
5hsEC2wTOMy8idA0QqhdHZZVi4hGJV9M6iSgOmKyKvjIoUFXdVe08M2Z2bbZc/CFIuBPJPthtFg0
WVObB+74g0a0m99UI3OgRY1GNF+y3Tja1cJV5B9U6emFxOyG3uSX6s1S+hAc0CAoPeU+N8c/o1Zf
mUPf1TR1NjzppdvNQpLXzBTSp4274KEPq1tnIannAK/h9Njzw1x7isfEgVGJ2IPMs2mNkmRBbj6c
CR6l7N7Q3Dk6tPz14lOkp1Cgkui+p2+5mfEq65bpa4t7cTaCJRgHm06Ed8hov/MHu4d6Pt9SYKUb
cG+W40W6pUkfniXxW2JqbDhIwiqpfvfOU1GL5Y62zHmoWD22VtbeNoJHcV7FV9m3OBRWKWntFh96
sbAD52UiNUi7v6zpSI564OnEdjsagvCCwnBWovYWavcxJVvaXXpJfZLOYJ5tbkxuuyFE+XSUpS1D
vpkm2CwCPCUy4TAlnkH9lg8wLAaswNJ+n3UxOi1uQINMONFjRscYQHv7hf6saVS7oH4efBQ+JCFP
r+qoMAKcsWCbIkBlMIazj5/vJZnz6YGFyFuV7gfBdKsQkpVdYx+DpMxpRYyQSUdVRQZHUImmSF05
pq5KpIIMfekwV7lBXpxGBpJUofFINMPZoE18TnJBvAHXYMfubyIioOEHAk3F16JbbzuNPLBedCp+
K+Phyzdoy9AuWpZljlRvBJdR1Eg/pu6GmC6L3CoNvINHefdutSWntIjXseWvzk/gdNMDD7Bqw4OR
oRUSDrxdEiFOrR4ci//Xj+mWrHRgnRdqSGPkV2fv5Lia/imSm3Cop/F5Qq+czmCLZ4H5NStoYiFa
NvIQB+Yc+/ugqcdYZWFLU7s9XmCigj20yAK/xC8v46I6A2/vC+5eGmpAPXDWUyrRXNOqOJXDYdxF
mn9FmpQTTDL6yNf8xAb323WwO+bFS9yGOHfZ7dbQr89Gn8b8JX5Nb76LGRNXf5+RjzGhaady33BF
KISUjvfHXc1grWN08XDUDMZtwb7ZIbPYEz5IvXIH2Q6dJKaCTcI8QMXs0NyyE379fFhxxje7+b4f
+WRGDw+ys1pjAOhj13aul4Z3UoGhdhETnQOlm0nFwjsEa+hVgR96xAeyr49GLuHm2sji1HZX6/6s
skEd3JIviVptK0tssUDgl3IZ89r+0nRqxwqlnfon7wZDv3w3bPdMtQ+1vIi1kkEr4RpGbeeC6/kp
H8e6wPn958Eoe9QlxE9PK6SaDj8wXK8TGraZxz98IgmNrT1FzGHcU3xNye6MWgZfdqmJKTdatcsm
os+AkZR4gdDDby2NqMWBRcnFAyGHgwdDh9ExzLuXX4dP0Rx6bsCLqI18vyvqRA6pxZDrQkeJ0zkT
X3Spu1RNmC9S00xrnzx91zkT+jXXJANjvvkdhp9NhyQ79XCvveogLR53fIHFvAxnOYGZTDMlS7Ep
r8QgmNNS+7uiBdWl2I1HbbQmEiClK+B3v0lFbDEZVLF57eCHnW5YWzYJHX1YtKUTtg64y1xyXv/f
mWuHsA/wY8yDXC9rQEQjFx+aBvlK/DOn5gGZDbOR7oK7pUC5EYSGXPfE6HxAAe7Tdzuza/9sxtuQ
A2ZSpboFM2Q9V6+OxptBHHfcpn+ho5uapMpD3rpcdPwaf6VAQCYFG6Um9vXIhIv8N8b17kX98zri
fSEldlwPSjWeX08KvmoHriUd2TFqXSeiowfZf522TlrARgHlEuEe5msBh0EpqY09LsPkji5XdXeI
11HnrCiTZcslMyXsFI/JPQdcCMzktgnHcuhgY2V1qZqOEXSJ36gl8OwcwWu+PijaT8GY2EpyzbY1
AT8cAd3NKMgn8nWlyX3Runike3Kn8KZ4N0d7vkPQpgjln+z+GDr0fu//PfBenWdm+rOpkYUT/7Fv
zuoWE7Y9TnOM+vcgoufyuVt2mBNTc1VgbgQNeYmjCtQo/+AfeSt62NoUwrHy/dNEi03QG1viWZIq
eisZV2T8BNniIKKiX+tBhkEw6aPw4lnXJlL84uxQEo5Or5X5+OSysH/LltD17QfxOnmkl0/lrHwc
NpB0jtZpXVhEZbcq+QsnRleGqX3Te+vg6b6XmpwUkpb6Rz0197f9XnVUREGi98tnlIoWizEFPoKr
795bDVOQOKVoFK2w9qqRA1jW85UOfkZA3cJmMZxKTAJ6zNULpNHNxY49Tdm53ah7xeutdJK9cIEa
E6w4/6wQc9YMjM3YR1HQIjHbKmnmtaF2o6H2hFpPgK+cDoNo+9rAQlnAwx7o5ShEmYgcmyPQ5/E/
PXG3BHqWtt2Nz3bgTTKi5Gn3qySwfSVYRHUMUd5FHsVEy4hc1T/LOSpC+EXNaSJzOuGZHvKqV6UX
c7PvKQgKv9nqRDpd0bboENUrCc/xVKLhFhZPoh2NEp0VB8cyQbVSdzH6F+ZTNC21HJZmBS5HRIff
VWSVeZrt2V1dhL4anvksNWBtdnaEpZ+CI40Z8dkVIQUw8Eke5Qx74yeI4/TLpnzcezCnwfruVjMZ
cjqMjzKCsCNiXUdaZlWCMduWJosAylujrzJnC2P1DINjVQ4JD+SyRAzjW/orzoflnYCfGMZVLaOg
xQi+szhPzegdAx21JbN3d9Jc1ADtM5SbZawwdtrSfyTVLi8uqdN2NSIznCsSPW+Qbd4TtXlOKu9a
7JhuCrSuxMIjiLw3XBHoI2n3hz3A5YWfJMwAdYshH6rFM2P2YtiL+wfBvsEFHaj3Po/Byiwhu6WO
dvUQn5A8otlz/en0oMtaN8v43OKae6U9Etcmy87VAqQ863e5a6smO0Pv75aIy6Ug8lTP2AGUzXZP
ZccImrnIaUr4fuIVuikWJkahsWkDZkxmNeSuw/sODPlqJ5Y+cMoruMl0Qh+FWeMByNsDgIYboJq8
6soiNi0ZgNsSJkVaaQj1kRvoJlpdn3p2iuTY17DEDdIAuj7H+MqFrNzQcQtnfD37KlsHkkSit94x
OmEW1stAji2WqeOwHD/BBrcxwjp+O5fgSIGRMG/9mGDsJLOdf63pbr8cHd59/QbCMcMjGBMzL7d9
hvCMXOQjkDq4nKe/ZgP5DAC1tw7qRNUaihakw7ENxt8W/+YGncEOwGd4DouAovoActP8j5y9RoMh
LroOeENdM7p94pBjo0TkOAMDNCpKT4BUI02g+M1xYLniOBk0pBeKsaukG2YH+NU2WcTzRNikDaHz
buQKY6NdRDy9ntFmPwfMd1nmm/vMPQn0maqWIYRcgMDcnvOSfDPBxs3TZX/pp1JrpRXUWouub7o0
yF1I2Mh7/VMv3rkQPC5CZJaIjW7+TxnoKco7muJtK5SN/M3PRS2HJTAOCpapLnSOdvJk623tcJAN
WL54bGZCDe1eb6IymU9u6W82ENfRF9vVj2BWG6Aiytj7Q+HtZAz9HQK+i+LsKViU8smqw1xioZCP
7YooITVfu4/OmytVa6mr/INnEYD73AxXPwpEJjyY9VZuUWdkUZnyap8foIcGOxD+R+xgm7iSmTIi
r/ztye/tG5Grldp4/mM7XcmBfeIF3uGTOpxexuAkPgn8baNj54TwRKYmENMPdPTYFzr8MdEIHWAy
bGxUYeaozemhP8WbKlX/j2dDS0I9I2X0DOgRkowwT2Sf+Pxd2g8TjteQohZJMi57oth2FjZatUGW
X0JTrBQapvdMhST1F69lIa3SDDjHOR2QJzxeRqzDZy0rY4BHw3lV/qqAbQoWIxMdgIHQb1eC5Hta
UP3Ykht6gMPyMadjMZmndRQmoQwPAnhO6F1DErg5Zy18yTs/YclDz/qskdZWXmlS45xgUAeGfxPE
i5DfbdnNHBvZuYWS8tpKJhmjPDskEKgpUekl3wG7myX7jsx29oDTBFVsuq6TtpftgregObfP0c7I
i6bzvqHC8bBIdcwKKhqpLpi467+0zR6iDUhoDh5LLHSFJb6tb1cF4uDl+x6K+J9SUzLYkiaEXuYC
SM2AZOtiTeRcFUg3MQNZpQVRVwNvgne91bjDjNQetUpQSnSZV4l66R4TyoolfktcnN43/13iVC/i
VjLK+XjMksj8shGJeLLb83+eUTj54fazqi2qCNsHorMu4SYnGRdB6kO8nnS+Ms9er+2HvML0r7ma
TjchmJWSzBRAQMSeZ+OUvKSouhkwfXL1ZkdzA3QuJx9wvzBp2IVKe0GN9rLJrOhJCvKJIVfrSBDa
xKrVfvB6yuvzy4UJwji3vOomvg+aDBAQwjRaAvxj1OxoUmCtygklmvWrOZR3ut0KZGSaw4akdZid
R2diJwy4DpQtOs2yrDWiNeZ9ShW2GH4IJxmRkVTTi+xohT9GO+0Xbev1/q0OiLJew1U5fcAG4v3i
V8oOLu/jJmgsijehjzuWleGIgPGkjeqmKToZKq8Ch0OBK0Kw2YS/tB1swjILVnuSipfJiFtZj6xq
t1ac5uXuzcfuIxBWRR+7+drHBsjC+Bgoagtt3Br4pVM1WfXp1yAuweTf8GOE9FYsKomI4hcWd7p3
stznGR7fM+DUo1L2X1c4wFYZTgaLdhAztq2oLxhTgDM3uqmKiEjnlRy0Yzfqr0gX7jjpAxWxOoNo
PEi+3honqFZCxyOUd9h69tYiFSsLq4nbcySl2VwPROzTwJvoSgF5d0B+1z9UtcWc/zEJnLJp+Yc1
CZ5Ztv3HGfw/SkGvrAba0NaMxNG/vQXeeWavUa3ASAg9JCzfp/2l54861qGNU+OUfJifsDKIdXni
K7nFnCYTY3fWZ3s18y620cu1KOSjRL7ioJQpi69hvSyTsJm312mrUp+rDCCjbeIBxCWHYlvXFlfJ
NpBBaBdy/PZ5XE6jzPmqlxjaOJw3VQBuydN3+HFkEnQ6FFQei7GgUn6S1jylAMNl2U9v3Cmju58V
GFO7fXNhiAHU3xW2aZhaYG10qV6STIPiZLv5NoPqDMan+mEC9aDxz3iTFRFnVGjxZYyoTvlJlfMm
f0pCzKZzrDmTaq0XLKYIu8zHjsaPI11hMl/eD9Nm2SZto//uXkdU6SXgBtJMpVWiJYGSgdfPkp3G
JjWpuoEl9WT2TOQ5r41fVCgSzY93pS48Dmk26aYfwPSk4OiCRmnQieJPG7otw4cz3PbmPevYCXMa
SbSSBO6KwtJ3fjW3eteuBI44q5luJs12CGGX1Iunb2gUE5QpXyg91nPQEmtLP2JQ/g9HzoSL2b/q
6jGD8MX/7wWWnVynwn8iAcdJHvnq7ohdBporKTkKMFHhX/MDJ+qgLDnLsE8HiGDXB1TytlsG/8Sr
7spZ2CHOn004wLTHQgt9I/bQC5ixFiywyTGk9DE7w6pP87A0HWshbLxNCSPlIGTEMX51BS6AfNWL
NTOC1nmdhDwCPjjEOANbILXoWPXEAAyBYekd5R8JVnawvrGZmZoUXASupjFJIvFEmkzpm/sypwFz
biXFts1YcAizFK1d1w0RyCa/xN+7EiCm7bq3yN98RLIMOSmchA4qdeWcLgkhThE6m44GpBOV4e25
+K9APAplxsN7pyIKNy/JiGzqPcBiwpoybwHTpqc1edN6NEh+WT7VEpS44M58+1yXMWbNrYiKwZYG
H9HC1zbjXf0O3+gtEIQ9wh6uD8A6Yh0FDckE9imsxJE2v9qeBATV3nBLrlxrfO5yOIodlgfBYfBh
vvum5i7C1opQRGq3fVKwo0XjNxQcSIqZ0FN/Odc08vJGM3rNFZusx5ShdY6gEyuY9MT0XGHwa65f
Hby45MH5Rro6ZH314NSf30ossSZaF0/sLBpIhFgV3nXX1Kwh2zAXViE0BKRhcuVuBlAlVAZsMbVt
bJCSiJRbDts3sQEe/GXsfF4p6k1F6i83mKVdIK0zArdVb3C0ixL7LxK+YjnK6CGGfZtGBHoKU2Qn
BKpRJdhFSQXgi7ObVxyygWcdqhTyFMRgok/xoxtdI0ORqHMkkLiCNtBMcqUN3F23hH9CfMzv0Mac
j0c5y98KdecgM/Yoe2BLf/EfckUHRwIhHn14UEmmAJJ8gf4c8smKV8pIJaTeSKAAM2o6YWAj1jXg
qWzjR57k0NdVdWNe2/6y1/80wwmXlynlbhzAk75Zabvxfe3sC/sV9wT4sYXmlGkMubwAiHJDwBi8
Fq04nNIy3azSydl+swk51oML7QvwiHmZ0Q08HqKgfJ2KjUwVttU+qw4bTQ7B9uzYXoMmrtUPUiNn
IuJ74X3Dnxg2viVEFuUB1FYzR+2yVu086U2zeB7cn2v8NlkYwKQ0yHvmAqVzC4CuV6mQZg7KJZIA
FAa83/d8jfKaRkoqh7XBWiaHi7K+q1LYPSNGWCNfFWbppyvVmtYsevrCp20rtUvjKXgmlBxtNQOF
rvXRKNYT3nU/d4/F+V9CwnkqltuxyZXpsQLfqov3+ftPSBXPaHt0WB6dJPIQjllpbD1/mnCXnSBe
OKL11cbMinxrEev0JA/KbQ6Ee29WpKNFgSB7+I9Lj2YcGg6HLyst1gLmTVaAPFl5YWOVIKjRzEwE
/2wZMo9KlhvLQJQnKRchg2l6ti7o/bsD8MbzFPmrriQeXRxjQcYjtVlagv06Wbn5gr+38y021F+D
xBdwxOBCxyPPxjt78pfNVXH6XBrxnUBZrDmNcG1C7eEhwilSnw+O39ak4PoLNP8ANAJeyGiq1nxK
8i4HAHAqhqM0AKiPyB+8FFZGXAb0sbugFWkpz2VDdIilXUoGLYaRV/MYq63LYHvx+DiRhH7YIMRd
5NcGTBWedzSTIvNSgUgT5a4S1EGzOZeWv0vnv6tpB19YFmivYvet1zeYjLcnfM6n5a6mIPiECDql
2Cf1rkjjkvzHX0DuLHAshgy5T+40YGcmQVeSB5Pbw0ZKXIfwlTtGM4WlehApzpTJP+HUudpIENlT
a2pB7oM2OjcVxPBrTDNf/wTErnPUuWBTQtbytGk9De/ic7vwtixxc0bGxaylB6GfNbVKaDDakT/t
G7EgiZyjZgLAF0/FnkA77vLpiv/4Vx3ObCQAzuXV3uFSLp4kSw2TzrPm7vInyv8n4wMMBcsz3l88
gcMCIdzNmg576i41v1Wk8439LOQL9j2H2jT8H8OYOa+1W/WDWXCqrns2A9T4/e1CnacqqcEUVr3j
kxA7+1BZM6idbgpXpC/0aTY1oA4GI4Hf8cwToPXcIiLcmALRe4xG6unoXSk4AaRpHBKSdsZqWr7M
ktDn1EbCi3ST+fL+gBI8MZji+3Ylnxruim9/rMVbaLHQmCZ+ordq07M4taEaYib0w5HggOeKpTsu
VJwWWgrPQrIAt/RVQwcXNPdyN7v+ObZvCbZhuLyFdVyXyGbSiwIlsjKO7JrjlahdKvLU6kp1AbPE
fgsN/gtzLYLOT9HWTdvL7BFnfu2zNwPxhTp2pHkFShTi0PteXp8ANlKxjUqgzcNtfgyIUpEt42Qi
T8MZRGhKNwDKLqtlcWJkpKzqT2tYdGwAQQs99I2x16DIFmCnUaNO2l7vwKmRWsyg7GLIbsXU+Rzn
hAu+8FcLKyDjMYXCZYq/yUg1FRJMscsfLDQOjw8U9fC2ICd+reWyzfQVwnSwxsl4cE11tQaS/EXl
MfQT/rCuVlLF9LRU8NANVBDaelMF8gAclFqPhx2uL4NBy7Ck2kVnhQLh/GqNSU12OiB+MOacBlLV
HMuhAokZgFQWSp2TYFMpjQzxEdpfzk+DjBy8RZUmOCS8OqZobdD502ruPS/EjiIqG4+mqOflbkdq
EiwKBk/oVVUDQQbB5WUw30C2msISt3HuZDnOZEvNKqkgx8jqiUVaWtA4fz7TRY76GX9TCLUq5kt1
QeQFXdbofbecR4SyrpdYeOqvyyxk5KzKytUQ+zAcDRwOn2MWW+VRjALZBvsYsXFoVGZYGmtdWFWv
mwWvn/iawCNsZzBx8eNZQo+1y2GgYTov02P9uhZHfXi17jSCs3VoSHZL7xU2fBbCitu0Ll+whE8l
cJWJcmGNNAQnjvU9osIEwBmAmvRabkyCa+Fd3sbN8iMkhxNsI0zd5VfzgXBNm6EtEu9Ev99bziW1
4rXCYJlh85zVcKZtuXM6F0OVw6E1FJmMX93JFXhELu1weyS2vhNCucxQUN9dXstLkQ5lJAgNXxm2
V+YpDzFdYG+0R+uNLD//frmXI/WY3eWgHfr9kyd6WbExXODHlRMa7/AfrB+tOAgGBrZxsx0KRk7s
Tk8bdrF3EWfrliXHNG5DQPZ/mBoVsLfjzpylKjypUBxCMP/4xliYb4eqZ5Fqd3Hcqi7cxmNyxzMn
LgDg9RRvvkOK+H0mdIjz/SGVJOyYF2Ly4yxoC0Ots3yERB9cfoFqPWtOoOoG69GQYOXvbChjxqeb
GeB2E1+hKE8ln8D6v2lRYtLgZyxuVysKIFhob1kmfiFM10fQDkChXYgVy+r9hiQazlbbOgEWlKKW
9vjdawIHFos/UCe43XDhqTkxfhvhKgTuetNVhi9vAk1gLiaakhXHmbAEpsLNvObd+J+959z/cFN3
NVPFy1SH/Z7n0kG7rr6P4Utl5KKmMI6m9VbfspDmUetm++PkLzuBe6pKxXymEeQVW60vp+GGLqgy
7TADiivKmPQ6pOdnTMqVRlMXNexBrsE4IE7vRSu2wfL3qzNDX6ZPJlfqvk0bUIfusflkxlfra4ho
WFGYgSwB/LIgbpVPf5JKUlOKft/kNh4t5asE84ERjx4QRCZ/dMArfITPvmawFU1iQ4fM8pVYqlpl
csKqrXg+dZ4liwgje54HzETgJpjsoOJE6ZQX3ohPkd46GKMVJCUQMAxhl2w2OEObe14acM5WRcht
e5SkWj+ruwHWxzlFIzicsducapViHrzmnFE7UdJu0VkSZXimLCQCfFzAzJfw3OJ6y1td6u1oJ0HO
Q2d9FWPPW42sifCW+kaRNz83PhAtMGCwGyGH/AJd0iB/QPZN9KgQePlRGwIfF2Z7er3e/tU7FgHM
LdOjaM53DJYDo0LN/RO22TtXneltCSxtqDifUHvlHbF7G9kbE5IBvBjMN1xPJCxcgJdtzs/rwxIO
7P4Xj5tEeDAcgpUBIyGBuHOpGd5DzSTYmZcULGYunDYkd5H3Sbzq9vfOIypA9igEkR7qTJHpSkzT
CSKx2oDgqFUeWUNxiAVvVJ6IO2+ImsUmRvY4So5d0n8bgi4K48KXlmx2jc8F22Zklp3PTsOn6zFq
snD+ECNGjaqTxAcaJZCQfZG4F5PtvXJiYXV8O9NnXsulhC44KqBpFyLVDAjo8pAzA9Pzt5UCiGBz
22zNuAHWwa638wY4nxChXtJOa8myFZRgQPQAmX4joU12sooo8sYxC6GHSIHcwPqEo3fhD4ZzDcmO
XvkjkbroWEw9SUPQklmDzNS7NwXR2ecsbuQKqonGqbhYFiWhc7kjUwkDLhNGExlUcV2lJxfQjtz2
Y7emqYQIIjyYxIsM+1hrkKYe5j5zHc7DOqCs3TcUR0KrqmucWKsOwqNnos77Ac+RAJ2UfidV8N3S
SfztX9wFnqT5r8W3aE8XvqKTX5c7AAg53AkVMPPaCa4Udo4tyvc5ywhQBEnZdyrRmH3UzhaTzoL9
FI6kO+036lAEkgl9RbJxdcdotvlDac00887W0iSn6RpSGWkdy1/vy7xTF6E7YSxXTIYLvVJjWcNp
fBntoVH5eoA3JaktrVerbKsl5Umz/oXDbvCnALOPaIl8pkU+XZD4eOQLohbVFNZYuBSq0Hzm4W5N
tgdwYf+uBnp4vpbrT4rbF4q9hmQpfP4W0+rdYzq7JHjWcQBZaK8zAtIaFWibKEfWlXprx4JychLu
KLCgXKkx5EsxBUQ21QvL2LLuGN64bmMj4k4b1MvONQpMb1qtDZl7kGs96ZWMhWEl4VeuqRpoOXei
5RT12t9rYyuenNDxRFJnuqw++VHGj6pnc/IbbKw//dQGTxAR1jQ39jpiUPczPIzlhw7P2/IT3qK/
TYKzZpM1wvTdUZnNc9ZgZEY+0yrYA9U8FUi0I4QlEaIS+mmg5d7mg27l8/9Ql5QrHGGC1sfWJO6b
uMyhYBu9B/am/T+RiNnLwPrGbtw3M4CqQMUWnmvP6SRCwJnYhe1Kuf75OVAQl5HQNSlJQS6l3zwf
aKcb4WTPGwjYdrazIUSwPd5Imz/fkU5zPkLwtGW83B39WfOdrldTRCQCarVKjJLBcnJAXEUbgeSw
MYGpPWwK2bTK61ZhrSgxnZPm4ZQ5Y/YmZT1Qjv78qLB8taCGdq1BrcPbuMYfSWCR7v4m3cGUC2a9
Osmja1h+9nsjVkqm15O7hn/BbRuQx/YRUmdtq7j49NUQimCVfG8t9qov/VTApiTUz003ksj2qe4B
1+8VvS1qUu7D3AH++AzL7Oqwd4WTRE6sZHAhgJNRgs+cP53UaGG1R1X/kZd4zTaIkL6Zoi0Awjw0
3v7e70p+Qi749jw3NVDKVS2EGiddvm/XYhhlyjikTnv87hZWu4dK9Mtbdvb4FjEQ2bxksoQbc17Y
/KA9xSmFBR/R2N17Y3QHUu05R2OJGFp/RT0fKlxcqlpGrRo//UUZK8LdNst8Q3M4gTTYEDTyZon8
nI0/vJR93SsF47Mo5FtcDEmemcrjSB/+Z7JyHOP+RCLl7EOuhPGFr4WbzmJO2qX0w5CedhB1cObh
P/I+oLFyCJTJz5KgvfYA0LJtrE8rp8bS95MQ7wkCazkqRudfkLzB60TXAxFzMAyie7StoZ1hUx1g
vpqhh/TO6OXyOw4GPhqfobRx3ImvJ30Lrc2FF0sCpa+2Jemexn9B5d7RgIEFgzMk/tdfMsLRcSya
O3bcwUMMdkdCmFFDXlXwOBgUPDPGU4MDf54DcT73aHtZcvtMVpk9Bd6GQv2xXH0btT3yE50G0aPl
xJ88Ysl6jgnmPFv/w2ZBNiQf2Q2MD53gtogZ98Pflnb3UwPhRW2MDW/Sps7hpGzCcvAUwqNF25tw
qumOvQy0GmjkrH7Ep+cRXfZW46+fzfzrUWy5Bm1xvnnPFDAWtzRM3+qTF1cqJ//DJk0dQC29I5ux
e5Rn4BI2HWN51GQsTy05xvhlDkZv5ceFI8XSDqQigDpnF/XBX3VBcaP/XVgnQtaIU68f09avafWK
G6brtmO4JUnLE5HZdmtXiPufFxIRJn6UGhaguj9eVsX2BI7X8NbCwtTTo9Mij+E8/Ve/rYq7oO8y
OuO4t/1a4LcIF3wYRBmTLHNiCCqJs7ZUxJmzC8AXrDDNXlZWOAbVJ1DJL22+idgjNkopjAhSSEUs
cMMfDccdBJocax7mgH/Tz1w4FjllmArKXCB7NLQI5kYTB1egy82B5llN/5Q4EBE6ODvBBX7sD/1k
iduR7l6BGH+EwwSbMl9nM0LJx66Pzjf+kpKJZw7Ll4hnIBgydj4NtkQt4Hwaw+JLn8mqfjWJPXt/
WL5K0/6mWcsdlBJBHDEKVh05ka5aK6b2Vi4ZTdHC2FTjdpE8Kvuk+8Xm87RtuI3iiXzPlVHhlhkY
3g6s/pOUfYIbOQoETY9qRIJ0Wr+JJpccUmTMQqvB3rNNOgP2VVSf65UJ8CpLsPzpqcfJy26AKR9n
6perNsSIGP0rdTsaT9FAzfzCyRuz04fQMwtRcQgXrjIJ/RjzKnfas0o5hjGm9tnhQ8zPNt7+CKmW
mM8SLZnhd7BBojsrgTYTc1ZRQBIKE+IReohAspXfSBNzUxlCMxrjI4CLThdPLdTnMOXTNuKQl75i
Gj/qmkkgcWzJy0iIQKqU5ovCtZQP1e0NcBlnxS30xxF3qlyY6im1tqJw8oAWDFUQ1hqsQoh/GxGE
WbT5RSrrTZZwQtmM9wGlgo32Kdg03dICGWLpa25p5L5XDyBRn37OlB9n6Taww1tdpSaM//zv3QIh
SRC5fSjYwp/BKmJ25Lp4ZuGuCafy8HXoRDiFHSX2ujgUvmoeKqnq0HvszVgXGTjCte0DQS5e91FM
mvC1fsy5d7Ut8gKw8xg3bWx5tTAxUDM7P0KUCY83lPVolmRTNxWJpyBZ3P05BLqRDoYy0G6+QRM6
kOtmmL+sU/apEdytLATG9YD/spbxXC0gYhQVAVhDAQ0WEcrnn1VMrIoX1cg0Lq3udetAwbMYTTMO
j4yWGFPsLrSQrfFKrbt7TbCF5bkbA8WVpAqoZdSgVvXpEEGY7udw2yzsrzDI0AF4dapu+ioEiiey
FkmEJWbrduvCTReIqbofEZVmzHnu8IkXZXGTIsf7OutId5BsjdKQhsYdWKCbcOzO4r7ykxBrv7N1
4GLNo4GgDYs6cxmiJO+NEJVAbpu9tsNhwlo4gNaM3qiZ6myRUuyoW7A6p/EYujvz8ElT32gYwxJZ
BiJmxkNxPpEBB90Zn04putNY3fHXyZWWNsrn0dEAGXHXpCVERq5Dzy65o+WYWFZsLVZvNomIRwkn
jI7ZzmQhgZYS1pp6wVJp5hG7/XkGHmnWZGI4QSSGIMmHtWrrpuAyouw/1yUZ0v6hBOhd2bRizHSy
/PW8pBduEcaZCHX14RebZJable+v9ibEO+WYaabp2nNkbdpM3Spf0lCGqp1mgkv6DYnqWx63yotC
ejUCSDY0h8Vtzr6PLgwzO00RaJpxJcq0KLurJnQAyg3K0jaMHrEgn7UKvTvTCUqwj4083lvkXOcW
IgIaOt6Bo7mNLdVJg5mgCk6mj6QllcYClXN3FMQ/G+/6sHrxHweSHHXGWkESli9U95teExB5V/0p
fcIyl5fhScMc4xYknIxB3K4MN5/v85Ba/NhTjOnr8YdGgmsSnUwSGZicZzqvyhylo0IKgkjtUlF+
e3VRwnMI8xg2qXI3C/7HdsVRD0GS4J+Wy5QcEyzJAMAxAPi7YTLlWyWjinPfUsE0N6wMlrbs0+RI
uUaId8GF/OBeha5oDgX6+EI+nt3irDOPciInSJYvfI6V4QvAMtpfK/W88EMYMofowQ8+4r0PUfpL
9bCivu9c79S4vEax9NOr+j62C+RzkF9LUPksSv0ICa4u2KaNvv7HKzuSFzsJDlUswFzoKqlwqc+p
I502kXJKB6lxOsm1oWN+s186+o5XLiCkIKmwv/1AlPUL6XopEfoNOyQbn10HCNNLKM12fMc0237j
C1Xb8/a7vg/V4QODvN3asbUidRXgzBabxsni7Tenue0GMiyiAMRbgtyVoEAAr/CgVBydMV7kMo1U
WxNk5BmmZzykspwp7WZLd1s3wdo7VeDhm+b9Vxe4HNbJ7TG+aifElS8B3Zd+OQCrjqO5KMD8ZL9q
DIPofxK2IhrDCK0Xv9O1EItNyxUFCCZqqbOk3cFTnV92yZAVTN3Tg/aVequuhs9vyXkqimDmSEag
mJfUdwRjp2C0Vw292Rqceq0UHXo6TDqtmHBEBGuhtqXqOFpWDXGGwZ815zNQ9IVVQaQY0n72H7Dm
77gLgiIyaEGfbZE6ObPx8NC7DO7B0/DAPsI2w5q0NXXIWE2UYj1FhsPHWqLj58xsRs1Q905tf7/P
/2ezkImCxBGKcyWttoYUrg7rk1Fi4Z2Vj+6jQ+yR726RDhNa+a8UwZ0PhynUFkLBWQoqCv+AKj+6
b5Z2xi85sVkxMrvERrEwzh9bRQ84DnQGADXsqqRE7FBiUVcg+mZi9AfeD9XRVW8c3s/pMAHurGFc
x2/SJRU7+qwLQVAbCXLzxnN7ExqgMlCu5sHtfH9z2xbiayFCUHu3/jRhuaIlnaar1qyMlwrWw27K
u8AqOFrQsEs2aenJcoWRRCCvL8lW8iQ3wKc+5cY/We3t4zweexSW+Kty9HZqZCowJSxJd1rYMTzH
aVZ8JUobYEh/nifgEHXirudZUsmYJZdFHtj9hakSeD3Uf7g7tjKbdnKkKcIND5hGFVeM8z/dZhFa
JsZY6YFpeXxiDRtZ/AKGOFWpA6iPWt0ptUHNFQSXKZ0rZH748i6yfk1uoJ8FB6I+zmP3XRzALo8y
fP690hKVqESFs5yP7pugLBjsHI54pXE6wwHcGkMTHyRAVyxk3vtM5yi7qD2GBjo7WVTuK3n4NCid
HQTjM33oxctnmI/gizZFoNsRVw0Ep13eo3j4e1YnG1+FFSW/s9+sgQDgN/M5ZAop9wZL0EPElEu8
Mhhnr1NWSa2akRYwMAZ6Ba/vlqI/4wZ/SyWd9iWEUCU+/2wS2nI1iuvXBuAiwgz0dEscSwZuVO1Q
NRO0kZrZLoOJPh0gDj5i8DbP2oKKuIarB5lX/ubypHZPiJoFSjan9Xg/aOzlAmSIgdfsVLE+dsfn
EHyJImMEvhYzER8xUXtbnxU0jGV5vW7ToA3xmCwYiHAr8YwyHKtOUGKECJUgOFaOhvV+5yuwEVhB
kJi7DT3naMiSQvd4T1MibZYDq7WEMI2GFcqZ23qFFLlpD5Yea4K/2g9+XkzmJKssUB0B7s2qaSwh
sR7v8ruNGRxMOcbpKmUdaj2BE8HfIKl5h2y6nsZaRbUnW4LJgM1CRTHvVEJ7mLonU6Gr92rMJKNb
xm6LB6tAj5AGDgSw2y+CyZ9ibyDw2lYE9bqT5aUoX/2+B8/MuYU2Jhvpr76dsNW+km1sI8E0VFPl
AE0l+vv7JpPm/Crl27gChwKTYN2mjUgEa7H1revWTn4YqIBy29qBsfzOf0zw37YH7lcc1Hwl7EVg
cn6zWAtX6xURo8GPcxJ+Y71k3fV6Gbpm+Me2FQ8TkEmdUXQTC8sJ3J6LRMSLbfDCQZW2zuV98Tfm
JuZWkj3dW4b0rzymJ99V6EAAxFDp9xbpFmoJnjrbYmYrmbsCw4WXY9Jp8Z1F1DE1DpC1pz9wRS39
6fUzKhvGnywaMp9ZO/A2Soc8WHIdhs6lxuwlzcDxLWvZMZB9mKM/ib58feltiRK6gwIHelYocgks
AzntebHJkdWJjT9nhqvtJ9UyugolW/uVnmDwT6u/N96dDfPqx+/rOzTz1gsPaSK0FWuVEHM5e/H9
Q6P7LDmeyZ4h1oPfl4RLtm5+9uWex8FuJz4sUMW9tgS9yLL5dWSSYQNOH+ub2CUfv/kvKR2Za6NP
bopNhxOQhNUPGQKQpORdB4fLX5tKWm6pJhzzxMzE84CiIf0gpdThQNjm3N1c7U5jKuD8tVKnuPGB
Oyltfu9qZNEZdT0trFJMNlBy7uaBtB4j40hzJy2/451uhNaMwu/gOYEosCBJ+P21Y+H/8PZ7G3vc
grbncjVfgy84ikuWiwYRqJ+4bWNG5W+pTy5OOQTa+W+oiw7sPCdLI9OFhN904ixLhac7WG0UlReH
VtT9xBNWPOl7gXx8J2wqbCqUd7EcFojatdMry+3QHZadDmLfVXTomtHQ2s3gXiIpkZyYV8Fiy8aj
8r0SWOKYM1/hOHVfqoPRPJ/33ICx9veQWyfL5QHKGrhwjWYRyUUcubkBPF8oCOXJqiAcr4xoP7Yf
XxTHlxKj/MJFRWHcS8gH12wzikDRwTsjCjX5jDbSle6W7wjU9jOxRos1eGuEdzvPLJxoptULYWjR
csREZN/0eFcBrDPwIIH1ACf8/dQ3iK3cf6OlJf7dEVHzwvY8HvhmCQ01aYexI+SK7MvUmIq8QPO9
XbP2Tgzs9rx5U8uI4nVaNxQWOVlegNKmQKqDqzHzGRbwP8nopah9uuzrRmHT2JoJ1UpoQ8iZebzz
KP5+eAQcmQTD3y37NnNn+D+KdXcK5eKRE3NNno1y6hOmhZTJBwiVVdNtA+KlGghNKMwWoGpnVI8E
dYg3srCVEdoXE08o0Xb5IJtMkvqDXbd9CBSSMiUW2uNBJ1jab/BHfG0YGusYe+oiQwfMmvcijKx6
5FEgvOysfxVfoHF+75eMbBb6j5+i51WXpdXMB5HujcYOrtD91vyvxWnhA/tWdWV1rml80d5YX2SI
HQ7YGSwTWIEW02z2WctF035rtXSSIBWU9EqrctjXw4mu7a1U22fg9Au0AGjy7Mjd01lVUBTtqv7H
JwwxT0kOeclFZlJ+kVAtl3druoGG8q0ARLpJ+nB3xc6ZtII+oxZ3s0Ge1EgqVYPPU22CFswV8H51
S8PHklEcuoKSMBXflQr7CZtmyG3cejcDv25LRqcJk/7KGU8wQOC3AHIeSEHDnBpUivgqghPnoEbq
MovK5JHVRfvy07veJiy9KZ3XuqQtjPSuHfjYm/0rgCTJsqKZ5K+xWqhZtuHdW9m6v93zhC19qIhK
2ywNgt0i5iz3Wu35S1HVUTIat/vuE2lMugrm/yqsdTJVrpxgVAKbGLUq1aN3N3XOR9m8KgLIXAY6
GrUVlFRDVFGKn5zf53eEjhOeYXzcc9A6c1zW2DDiZTyYJ/lGoEBmz171d8Jqm2mOzqXrLbTXlwEE
RYEscF5xplOqMToWrgOdk5KXi24cx2Iw7nE0Gr5LOFX5L4ng7z576lG9u5bQp3WurapAUhhCDDSH
5Rf3fmVn06oxjA3IXILPD/8NK36CJcD6Jj+uoZm+a76wRUYaWTIIwkQpilvKhJ1QJF34Tiqo4SRP
50+ox33qb+m3pnD9J+XwQrQ2Wqma18G+50dam3txOmDmzKhjqO3AwbDldFg5mJjBvji+2pnC6nVQ
ZP3bLOAQQ8NAZMBKBsLZD4gskTpsJLyynMRpmQ5f6lLxHAcZ6L5loGRljETsbPqYb7N9ETTDHv0Q
gUlKQ3MWu0ra7Fu4FHJS6YVcPfeUiGdlcvpwykkMEMdQ8oEz2PyL95p90vzT0iw8cYKbvlBjlq1q
e3QyuDjxoH/lwRGzXeVHU7p4K4lf1PQuyeHAgdQp3HhCJ8uVwRx0Hl+VjJqM2SZ0kbwZ6yC1Ho4J
VZM0nC+wc7bPtcAj39x/0ougdtoo8PvUQ/Qa3eVBBofFmtv3xsiCwde345Ztt9H0GppIYFUv9Hvi
ns6Thl6wzIXaxf+PTLglw7Tn3WyFMIlGgTqSbOCchZAjPqwJ9iP4wEE6zMGsOy8fc798Lf6zSv2D
MRQr6Koe6hEduasi+C3t6le6lPragg7gPJq6zVgvp55OuvwforPGSnGWTVAGasUzLGcIkDtSTBGo
Ly5iPzN1U8r2Hs2bJkd/XkOwVwHeAlvjsMdJ5G4wChn+Bri9serstU+6pWv71UNvx9YmQ5q65Qpf
t12P4zsNfqsOtrG/JaU6gOdV2MmoQNPrNn51EpWhPQ9H9g5krwR2FumpyLwWyZhY94XIMtugXqNR
GrtTg3WUUy8PpZuujeplDZELUhn8p8KgUiQA+8ZMDgP2W7MDk1BpGqbdpzueAx1pPjqisrraKQ/W
AqXnYDbK6yYLw4R7jetnD7WhZzNnUYiSPVEPTJr+PovCitTpggvQA4g5nCFvbJPpM6s2YCLztRN3
D2CkHB8ISCuKs6NePL5Pf+s3VyDgQb5CjdkBZjpW4qXY62urhHVSIBJQu3qSkarpR0Dm0aQm3e1u
uXTyFEEDRYma3s3DePXoTDE6eBAZ/gpHZ4NHBKcYhTCN6fx143nIMmUobzYIATndKQ5v6XE/480O
7X+7lPcxbKej4b18cpMUJATj73VS0otpTkgnMuvuQP6mni0CBxgo7WdUOGqlEZdjGHmon1EkcTVW
NgAyVxON1LfiNkyBoqVwhS+bykAzQaRqA4qqWJjUAI3LNINAz5r5zo0eF+FDo9M58bGI0HgesZBF
rNWi/cuZeszBkme3jSEt2a9On0yH6PVj7f/DyafqCrVs6aNh5nDA5ALkhToic2+yZYUhID34DpDH
mlRuuzywGTsBustbu070we1lMWbonAfTOxMtcu8D5cU6ceAo3xUGTUYj94LYGv5s+594+oGMuSs2
IZrvgL2SBzo71mv9+fulOcXcbDE+T8BV/aXDuXlkinGsXYbEV1gAD1tzhonnoBhS1g83HkjHNaED
haG4uX+RIpWDeDOYjRyd+uwW0EM5oSvmxMLjvxXY93ZWCGsP3ANOifcpB5rQwM2rtraaBsJULDW7
LUZHFuj3Y2bdPfL31psHl33O4h9mL0ATTURTkZ9QpB/Xk2ZElyAyrWNC2LlT95D8LQBVR0tWZpv8
1FU+WM4D8PFES3qwOjrxX6rvbsLMgUytcW69QUY47XzZa+QnlENI2m+jzDOc+JfEg7cOK0EuO66C
OdaFTepPZ8QNggHZXWRn/rmRBy/2MN4ukxrCYZkKf/bIja+smLIfogGUPyLzVPxiigv7aofPc8I9
fNKrw+z5dmRiRMK0xV8XFHvFE5yvzcpw3Qw/SSAIDmehjNeG1FU3psQMq1GVICjm9XHlMZ7PWWqG
sy8rK260A/zkj+fm/HyM0Cti+X6Gxjs6SWyOv5eCodAuk3NzCOGPB7CC4vX2CEi1D7anxRtDoJoa
YUhH976WejH4d91rlZn7tR3uU3OgCOe6ok7aBTrKYY+Q2cBktkd8FTXdnYFwJcNvOgGlWub2sKuR
90ZJK14Cqb2wn5URpSjRd1F9b4fB1kn/KXT2NDasziC1t6ODExRY2dFlMXf5j8eESDNrjxU/QSFu
6Ggnq/WT7B6aFpfah3CMe2ET0eDNtOr6opfH1XmKSXOeeBDKCyCbYSpfPJOiGrK5AnmcSsiNM4Tm
1in4yEuHafyGPBR39qEAzo/1jU5TyGwVH4nQ/UVM9Qbpx1TGd/MW9bV5s59woqzq3rqW5bwLiG2j
efMkPl/iamZTyU+mRLg5m9A4VbtuKpPDnhS/3Za4DzUdkRNrmWm0ixhvZtjtaX2901U1IZZ/N7rN
fBLyy5TJN/HIRO8B1NUKxID2mjJeYYopD7yLZyMAKtIdpg3EGT0RhKE5Ou5wFHSa1QVv9gXDp/zj
Yiyt8IpHNtEEzMcmn9ADJyLD3gQMZ3LCpGEiikG4OZPp5pDGkjcmZt8Do/Ya+I9XJvp7rIljW+4K
wNKRbyl743VY388UOiBCWFJG8NmWsuUjTh45q+GThYZVFtmpivU2Okt+Nhxi7rCdNI4Dg2qBSBWr
4KI+90pzlQUc57QET6aRznLRfGlXnstsdQLWIhYNf1G5HEBHMniBMLSK5Kox7ffwX6F1+r3ep097
Gtg7rv6o/fVGE3KJ5dJlDNOrAg6MqDuCs/V3W/mKtY6pGgs0YwISI3/i08t984NnBlFX7DJYW9h6
c1llK8SoRVwjAcD1RV2/ATzde/XU+tRb2VnzZZnRWdXcflDLLalURb3QgdMnm9zsPEOpyfGl6y2L
pZH1ClIrTrDPZJvmo9BAD1QX6/eMqQu8zPif4dAJdkWB1LgAxVCNhODdF5aep0FCkPpntAgVvYIG
ZjOa5Rl9M667X2Ac3A8sHoot06m1PQBzdECGnWr2Q8c2wpj6pJHmgMO56BxwcTI9zDMcLyKrhn7a
5L8ojo5uzfbDfAAEG4pMGo2VgreVJb2u+odNWhukxFeTCk0QXMZeAJASm+tY99mkIGXuFyZfcrrN
W/WxIC04x+no+MoxVstMJE2eFJTcAaPj1GhURroOyl/tD8/aWu7RVCR9LDR78n99FBGzRTxs2+Au
VMsmUKjsGMFZcbDPDRA105a2H2bNlAra2PHGpVYkO1FBHmFKKr52eTJo+57PClClVNiC6CdzjnuH
Q4M6DzH47QM3DQBIshKJDFsMiNXSX4M7mIq2sM8blyMn9dClTRRf4yPGeYocDdOfS+1V6JS0oDTR
BRruoqNPKHHWiH3m6oZf67pBCfK4zyuNV1bpkQB1Y6IayACIMUKwUdWnQOX9SpZHSWH+m/lA5U/E
Y2b9EpzKr29IXjRejgw6IuzkiL+bIRQqrSXA59IuPjtjjvPTCVNVgNKEwMfcqxyNhKfFXZFNCUny
QaWD3lmZrtbD/Rkvdsx7khBS4/IjeFB5+kj1Ls65ga1ipccOd4VBz0UvdBxz6ETryqpWBBbs+bhO
cvryE1yjhz96u2wCh0O4QPuUN970jpSQncCA4ux41+SmL8WZdi7OoC8ywUv6W1g50Z5co7p7rVwn
P5jXS8JlZfFRqGnmjH5qjOCz+KTnt+UtmkPUJ7/4NzwFwfTFxAhLVC1uJ+OsahMEw4aFGIuC3D4W
9ZpaMiZHPfwv5yzu711ahinXWW+QHsiqV749Pr9K81Y6/JW6pWhXoZHIFiOY/Fn9PACK6ZJ/zXcW
U3GQ65coAH4GGJlFJnMXyeaCW8JB6mC8GxvkDbVg3360+eHJ4N5fpzyRSqeYNjd9NS30It5F++I5
+OukIBCeoW4u+xwqzu//5XxqFlt+bX8OHHMVNtj4rapjGz8r/Dlj8EdTRPO+pgdWeHO6dfjntfDb
RcMjZIAwX7veHz7nT6/MUZcObmPHqToNIgJu8mIfpjUAOM6JqVwcGxzljO5/vTPHr6HEfxDUleBo
dPLaLRT1uU1+RG4AhdYREBjs/T893NkzSTH+815ETtXgohLw1zsH4TfVIB9oE2X+3PsquN0Go8I4
diVJNmuUPDOk3v0acgGt2GFW5z95onaeXUxo1HZ2wzVlwqlcz6q9qdFo63xq7cyulL31Na7emdX6
I1koFHF/3CduIddZs4QrpMX1zbVQOABvMbGRrfTwY9PUtu7xwf2CkgGocYsgj+Pb55mCydHZ1J43
O0s1YOtLhDf1ehuXoCZg55+QKSknKe+Cc7k+2/I+RRWHXe4IQMHDv/ZKBtxKjDcE0fEHY7kXaFbH
Os6mq9G9ja6yHV+B4vQJDLe4ubBJg0ZDKquFgb9VxFC+b3o5mZSEMxC7V8m181//kr8owm26cSQX
Rvam1VFMC6+IviYvqWSc2l+aTZk2UjxTCix3ouS65riquooc+JvaoGKbwVC/JDZcM4we+eM+mbac
31/x4w+HqiZ8Qchwpg+5i7+jOlnGzxKYM9naMH3CJfHKvChwucmOLeaet+7bzk9rUylWQvBWZGui
RcLwg63+I62cV5Z2u+8V5Ho5mwE2GLHE9kAwd3PIFVL+uymAFE7HSf0mJJfixxdJu39KN8/frxRV
mA/MhEZhK8piQFRaZfhvg1UlvX3LpEMpHZ+887V+oNfJM2WD9rIxDUajo9rB1QkO0diRRKVYm2EV
8LgSVnOJqTmRaYwenlfMkhqWCiP04eywzQCvQ0kEO77pZKW76tUZe2I3Obdw9A+RkRRJrDrcFOBb
7ipmGSS9gWzL/Nd5dtfA/AN32tYnzDOyAtwvI0Ly1VOgIKsd3s06NWvsQDqk+ExaHK2wpGCJWiAi
GyneKkul8KuPEDOzXXRnyKWufj62a9+4IVq6MxujSPfa1KoydibhTONaqC+Qi/S2PqKIQxzw0zV1
6Y7/EKRPIhn1Jsx+v3Ou3wzOIKbFvMxbjHeEawB2Nd4HgfDUXigwlKUNSH6FCMP52v0ySEw9IJYs
leOYmFK5Dgfn/3145omO/6/sizKdpMc+y20V061+lOLUCaPxh8BhUn5Hm1A1BULQYTX79lnlk8MR
IhdwCb62Z55e4qeQns3dmh1Xver5yqv0kkXXgr+45Od/slrrErOn4rMfz6APhMRyCOZyMUSv+pg0
urO8kuPcmL4CCTb4O+kMSJVNY6IgVobD+05OKPtOoLl2JpFYtQkoHZTLfklIAWdI3zc6cguLdc9Y
aIQ3MnguB12TPN41C86Ko3PbfawnXPi4dwxJayWH9uN+Gdz8YwWNAcFPefU3Ob32w7BSomOoyT2P
UMBgrWhf+vpIE9NlndPCbEjn11uybru4WcjrnmfFiHOOXbqoA7EtpA29FbggdSUCoRTfouMCkotI
PGRkcWHb55WqSpHj9T7GQ6YYvm44RVIaeXvrnw3i1yHc9GODsIYqBWyJGdsUcwpbW6xOultH5aIQ
goreQ6i9NG+w7w/QfyMfIbPTdIA2N28twAdyAIAc+WrM/+3KM6XUwH0IXu4ySu51VPmvmxfuX0i2
3juhp+v8tYfUtCLUOlpwqgTJwTNStysGb1osdKgp9xMZToppyxRhdMOgG8TSlX2x80RJTb96EBwZ
nCdgEvqVfuMqc2XhZe7US0TgpcdsMRVSp3qmI1FadN84DyVz24I0rpT32cUxU8DdKtEbieMTm6FU
QG+Kwn69cYPTPPKU9B6ahZwcMHWskeKX2HM/dsKUsK6hzDpltvno4mwPs+6CGuGjsmGGm8VuEjR7
zxcWwjeU/2kx5kZBc3GwF/CZAaI6zHJRD/WOnOJ7c9yQi5Poo22wDrtLRx++/rrSaDwRIbNSDfxD
9pBi+VAWp+LE8yk8Hf6fVGSJwhTNFjK9GfR0XCcGmXRVwotZb8JapeQz53Udht4+HLcU+NVsxTQx
xvBecZMoMKn/fGkpaH1TYuVznicSWvRgPcbypLNW4kSFwH64ZEvUisYE7cR3LTMJeowz+nop0Fwu
CREEalgM8boDxCd8zZOAi+KFCPYsdzBHvNlgtSMqmuu4AG9Plea3CPmJ0ut8AZHOhItAScKf52V7
cYqlkLg70JEflrdSttOBpZkl+HSDe/kM8ua2u75ly0Vsz3+y6BvhREPWuCZ+6Qqvz71Bxj68DsaF
yKvP1mYTVi5RsXDuIZTMqLt1auMSAfW26DGF5DOzvimIsjvZTYVH/YU4DUzy04bfwdSoQIU6oKsq
9VvVdK3TId7rIpop6yN1Z2/YsQGvM/vQb0267ORxsH0vJTpn0RHaGGHdMrko17oAMmVhHRhP465V
YoBmDzhkPbv0wGsom2xBEmIWd46FUgKjISCWxJK2Jxd1xQ27taGes2/hJDUTn9gE4/YNIkF4OpDu
bNRn0QFDaedyuJ52AFqPVHi02cPflqeVOooJoA70y3cFRgzFr+jotzyBjREtLlX0gFIxQiXO0lMh
HY/Qw5YdDZhv8NBB/P/kXoa3IUCPalgnZAb0TPkX4Gj3y5yCSECNwDZJLxb9GRiX9V5wSqhPWb+i
ops69iIAcjeQGvJG0wlYRisCDYwShFD1EKj+hTGPwJcNBcMnbLhUjjM85iDECvFg8ysy5H+Vn3oR
88TeZjE6ePjvnRF/dKS65a2PuYYZRfu3Gm+jPfbNHwP6rj2hB1OMBZsc5XXM+bIDZuwKLx2WK3vv
6pq4sn2GtW7qlVJpTJM+7h/wTBv5vh3hoM+wTInyUCVhdg+hWruJFE3F9Oko7+8H2Zsbt3bcJ2ke
xNtWYjai5id/dz30VPQ9J/7/WqMKdw6iqJu4XRV7ccF+9NpZJaT4RT9OTTOlxCFax0wi3PgjUp0p
u7lWIUkXxvhWPgdhRLvhacZdw1B4AFhBLKzx5yWGpHS8+nwBT1hK1sl21eYAH13Kvs8dZAeQID7n
peqMhv0IV0kP6TEr6GvziERyyQEuDrjs1Y3kBjk3kJvFdU88dqqMEI/oMK0TuIutybjB7/Ry3qMQ
UdyDIGtc7tjXXihASM1BLIIF/PJDZRu521eCP1Fvckt/VOuNV4eBoo8K/R1rnewLnCdJcWQYiC8r
c0rcvEbkj3go4mN5pslzniaoO+gHEA0Pnec8GgGrirdlrlcud6nuyZORVUFKW4gVePJtcHfcTCNT
BYmvxX4fBHOunB7NOB6P3zLkqzGdTW4sZPS6O9vg75mSeDeTI05Ge+vOJ91KPTWOL1Z1YtNcstEz
m07QvntIGEI/omA22H5ux51kjqB2q5ZNvZ1EhQOZm00zHOx+HfKBGBFvxslyoPPDLZbGLk4CaaPq
+z2008RWuYpt1FGWUYVg83QOoUI11B7lbsK97rrqd4ZxFiKyXmzcFBXzY/CwvzZCWrfXkfRzrldt
EW4Qqfk395L5Z+Cfje56YKUtv8+JMm0DHyk8ID6YXdykM8NYWiXy1DMbDmAPoMQ53T7JZZcHBWZv
vVrF83p2JDXqIC4Jf5br7vv8sivQNwlz2i311msFjvm3dkU1KLqDqVDJdySL39NZprzT3nrR4mRL
64RjjrDHo3W1CTn4vtnwvbHZdyMgTHLRfoXN0ppen5pEtH9efFuNzFNmLSXxVyWXlkZmXQDx4pL5
6zzg6yHUl/jIgxTGgyfDou6ww4q2fPmc/0009w0qM1zPy5hisgcCzepdDgCWejd7B9zg0TrW4bgv
FCAZ3Blhf1xi9YnjVWNvxQq9vFAyofnjFd+6qKPMy3IPvpWxtBKxri0QuFLnvIW8fqgiChnI9SYc
3k6LBhbCRTUx4uT40f+zgDKkeFUg4ikedGCTTQIBjMC9x7pskVkCRyVpNW10XT1kSWIMvCJn+/sC
eAVOwd30lUGQjafVmhn2dskAVXABHTGcoBdVubXc7BFLHiRjpbssn9SQhs3zdHGQaLz5ZUANX1Zv
w34fxMO/Dl9VeY/IIxeibfmk4nsQo4lCqO2lhjrzEVPo5+wRSRUBB6/7jQgbIrnIgjNL6oHT73R4
HrLLlCHgvccfquoNOUIdONQarfC8KlVDR9iIxyC1ivmxSgXnBmLYvmx6aBQJa0DbK/ya0WXe6V3x
IjNgJl/VlZWJqNxcQHB1OWEtE6gkxKVixt86YMK/0usHDJ3+pqTPn9EeRRC470eCjVJv+QoR0VCT
TwjoeNnyqKFDTEN6vT5nD3hs4mJi7czvo3BV/YKqDY1JU+LpgvC0bdT/aQtIGeL/qUGjxyV8mK6N
2n4IYdv4vXyOpws3JkI0Q/C4qtf3szVngSUaHATEBIz/ZIcKpnXGNfEGYY5HuYhGYzk9/mBP8gtl
m7Aea2UfTkGuy/KtTIDhZirxZqgxDgUm4A4ES2FGxJGzu3wR3PW/5kfR94EYKPyrieApmQwDlgiz
i7SQdE9Rkc41E2HBopnatOpaKzgSs6oyyNi45PXVOvFM+S8mRYNFJy9zLbVapEu8prSHzJe0KlfJ
hoAwAz2IVClOUK2CLG/F115E//oI3G8613HygWL3f1W4cGSJDRA1pHoddR5RdeSzQAEsbwtcZKlo
8nzCwRfZ2eg/VBEqVZvx5Lqw387gJS0rc8v9CQDNcFBlrvIeEG+aFM/r2sjJJls4GC1egTX0frRa
k2iydyWZIvlzrBQNVhQqpEoip1U7PJ29WrvHPZZw/DsR7NWE7Fy/JMhAFIUTi40oXCZsU/Is0or6
sN1U0ahnLZLb/IcqzT99yrhcJ87V8iFlA9smElaI0UM7E4HRnrHP9sKcNwxaoR7gcvv+McYYkQgp
ckHEmjQJnJRcxs7OIuoqHUSFUV4/ryY0QoXMmxUUUkCACVzs0pzkJD188JHx2JBdo1I4DChbg6t1
W0X3jo4cbUKBkta8v/nmX1Bofv0TWvNG4XNSuXOPBCweua5YEV48DNwnqKoHDVfl5ZMB0zYAcBi2
VlKktZ4YOhFftl8c3E5TwO5Jj9eesIXOmmUecxKtd2KU9d7qaUxs0tGLSWjjlCIzE000m71SUHYU
x3yAPnjBsAjC3mC088IN1FNhG5NEIVsONFT+U+fu3+GNovNjhsINBqC/l0TQC3zQsYREJbNJYqnn
tNjXnlrko9gIKZ0DMn/0HaizcdEJ2DvD+9h8Z9L8zDmxYoOiJdbLq1le/kjUTyG751GQmFlWnKB8
3QjvHx/xy8jGwpgZ0PdWqnRAU/qDA9BJgElRPtZdvq8TaRSJUc8W9dLblUF0BYFZ5G06pgCXrlE/
CwiFmgEkN9n4lw8oavczqLl65ZDEfnDeRPxqNuaMB16IzMlTX5ThnO9NCKZ/AznSjSLta+sa65a0
K8ks5tQJ9Z4cZ1xmbRdF0LcEEMsMmDziovDlJE0Ww5GQZ2eHlu+DCToZ5AghgAqg7QJOckfo4Khf
vQ4wU9ncW9GkFKG9Eg1j9xQLuj6xh3wpKI+Wu6l0B6T29KyLoR4UP31L/xbq+P013GV1cO5KLJCc
fgXVGDD6+5d3wmovD7JAsPY4ZvvKj0E8avaI+McrVUmUjZb444WmdBKQVt+e+cq7iGM/SFIiP3dn
ek1vFm1hFFS7b+gjnY6AAcqxnI7ib70q5NNB0dhcuk9zLq6LXeFwon1CiC7rQpHHUt6uQJ6LXPhy
D9pBBTb/EA1/P8eRjnfxiSLAPj13pDljXOHym9oaqwiCIBjzXVxH2BArqNQegUfbrM1taHC3myMR
aV4tZs/ZiKRPKwO6p02TL8dU6RknuUXgR1V2pNT89VETmQGXeVnA1zNf54Xh3NRoYfaiCVk6oKwu
eXhQcn2eooSgju5mc5wLdGH96O4F5832FYrk7FBm2w9YG0dsLDckhkPYplAHxr9dx+q+j0NzBugm
u/zJLW3dNocYnMfffdaaN4eUrLmG9+cTc6TlAzFO0s1EFe4IR9gWtg/d8awRPCKLo4tePhycpfrT
v7Qx/clBw51uqu/uREaHV3rdXnv2lydvGtCjTf2PgVE8vogGBhqGO70RWTUTMtlsCtqZm6Fwlge0
fIESd+zLAvIlIH2hMCvsjrR/5N4cY4+o7rMNDTgH8MokvCtCDrwWEdLg4CB2YR8YcUUnw4ut0O9e
FbKhk3Vq1W96LG4NyazsKQLLnU2yh55lq99U9Jt/tm1GulZgPK2sGkacCM048AHtgBN7uf7GVHb6
EaK3cmeO0PcLa8uCeTVqjTgRIKpq/1wMRBnSD5kl2vDbGXSOcBsdL5h2zwG+hBSUC69Jiqehy+7h
D9mQKTn618cZU77U4nrodUD54kqfYVwJpe1dHpe9OodZHE52eoUh6K77fo2S6VEF1CbmBynQ8LLD
o/xVyNRK6ZN8uFNXQSyQ1BFlYgwtV0W4SofWdDCkvIYquO/ZNITTpRxhBluu5a0dMIskEy2xm+7P
DCuOSXPdZ5oiiDl06osdxkYWeyDfjqmb1YwjQH++y8a8ZR0Vu1U/IerH9Ur/RGmt4eIlhSfKuxTw
REuCgEB0Ggm/+BH6nelD4UjnFXWTuM/ia0ctkOTy1HPAjpFIrxKbKqGUUMGmjxdNeB48/+3k9BE/
G2CJLVnhOYD9JYnNxhPqVJMWOPaAKd6SDRFSR8fhEIhoFUx7/Q+l7UwqquRBbeELLiEXAUwjkK7l
l1beM0P3SS3+Onww6fsIWBAaN+DEht2PWqY1V2Skg46GYS9FMZGvMOKbRZ3HKdnENLQKgDmu0CUM
rKrP8ssSxjYKJz69W5NwdGC66fxGfce+MGZRbjvzpxnoBmku2TdNgIjSy4kSz11lOTDsH2+kwty+
ZIXlizt10W76sT9P1mrBrqFN9gI1aL/c88/ONEv1fbgj1gzUY77H8wCggB37kuFsM3daQn3c+ueU
KJhIwYuMHxzNrolYoGj1tVT7UHjYJJlZ77gaRTKYfsrrCfcGdYlZCXyseFr9BmyG8DNhrLLa9a0a
8RIvbmFGdgoNkj0YVhv7ciHTjbtko3Dk3o3wpFOHdye5r+BH6O23qOcQz6bD+rkZ/Pu0mSwPK3Uu
y2dx47c3HO8jTKjr4zWr6omFypicL9si04swa69OCVhqW93C6hdl31KLA5qTZ8aXmuJJ0SWquhFH
K8yvLELeLJFIrTAtooC1j4NB5H64bEnHDbxUUWW3m6HfW/9E2WDNX3UKq1Msy6iAKMbH3h2ldXDe
/x6pF2Q2VC1maWado8gvGzxodrTrLTvTbOuENEisPmmPctH9ssoVIDWsZgTiLJqbbZ9kpU8U7K7T
9BdJWJ4zUQyZr7zczohbxDJgjXVeSdXwW1dVW/ffU/vFf9JymD5tRr2QEUf87PGdweE6sJqluVdT
MGZH7kI9mn1STDEa94c4msCZL3SaFsirT/WgCedcC1fcIvOtyE6WaQC7B05Zw8DwDSZqBp2crVGz
DxaOomrbm9W1m+gzUkXforrno9/sVfkB69dloCn6TfAMgewb5i7Tu5T6A1niJYWex00kx44Xc7jV
jBvAutIAwWsGcXCKbb0osOEuPBfTbPQ9r8Vzig8xJEq0XJ/OlzJPCAQvlk9JSzr4uaRXUxIcAnkY
285DkQ9WxdVMclslxFU4OJ/ijtysb4h895p2US/AcTThorqSueXYPOfMRzj0Il5V1babRVMRDHe/
c+9ZfmOUWxbKV83EJKdQDoTTefMYI/q/i18vXCyWb/Vs0XK864KktstwSp9MIz+xCfawSyJ8oUiF
e+8ZZdvfVs0Ic3JVEH1M8HkY4PeJTIegOUr1kyB7hXgm90z6+v3FN9iOv28Q6phove+qlg7gVQm8
yx3xKznyk9Ysf7BT1LCs95xyXohz869AByuwAYksX3FtfKlsHvDVZaxZALfpsNBe7wSofGMulYvs
Vi4YebzMLFXlm/sC4PcT2vdH81fYeQeRT00UBVywx3pdsnlTKrjNeXKh/CMX0oODbcH1AU6F9lzq
J9soWeWAmmGxWtt9kY3vuCnEPIe5fElss6ysMOcmHd9FbU95paVEBx8f2Wlsuq28nBrOTjvhJWug
rnREVDcQvdo0O5QcnZwmmhi1B+VxYPO+llLb+tx5vPkn7SgpkIl5DrJD+jPuesofYjcm8hSMUKg/
UhwF5rQd3d5pFdAsQdJ6MwdCkMnVUh/ExEvMY2U6RJ06HBCHf+qvAt1zfquPmmPL7H+/lVYOETtH
xowr97k8NFkOQ2gp00rACajQwdRmbZoXXcPOo1Ysga9DCL1EOMUJ0UcINtKuxPcuOVx6KozCtP5Q
fgevvtRZKn0r6OhrQT+M+dHHOPSWZrEeCGhNJNiPHVdIv+wNoBDzBg9hJbxH2hgqYPPGLozlb8hW
VUs0+jR0mV37pqPl/3THnmFWPhNRlS1F3LSBGvox5apjhPhUSvd9fKAx8IA+aEZsevRww/oOOwBd
6KE30tMrDrRbuhyRntbiAwBGPsBNUHml9a9m48Qqp5z27sOgQFKtwQ8Gk1a0FVDEZ7u2mI60J7lZ
ZupzK3DCT87qMUMGGv2SLG61jENiFUAK/aCmPfINX1+TQa2nC5a3SZ19lDqdKuJCk7WF+SxBwDoH
ILiP5nBsDfoYKyCnlGt7pfqoHjLYif+gPMvyo3bYdYcMz72ME25WHqyhd4fq420y4Z+Fxk+sT4oo
YS37/RYUFx1q8Fqp5ue38yQAn7DLkAmzzRdcqYxmUOqal8KRLrWSNuqddLlNWnrOVxf81SjzYbcF
uX7E1K07IXxeCxZv97Jv0h7UWT6H7WspWaipOKQfmMtlxubwMqiXEopbCp0Xo/NtEWBngrsJFq+z
t6/iUZV3Rj7JN/CAsmrr9KSKBr8zaf3vb6xM9Y60mjPmtCmsXQnN8tpj0SPjy4n+d4/0ofPEDos6
hqD5uRuU8KV7IAVr6bRxO3nb+0fwurlGnBg8ObWOWIbl8oaMBvZ8GoEeXC1hUoWEBOzD5Nqojw3V
EiDucjq41sMnbC6id3zuswqh+HBcn2uhlAUKRg6XWQfmX92/PqoPm7+zIRjIrhVjfMGrMUiXthhH
V2qdutMzSVOk3k9Art1C7GdA9CBOkTXgVRVLYQUb/5GvrQTw9GUbBmxFfhwEwup/ma2zPfYxjeiI
/vD1GNPvLzATl0t0X1bX+OJeeES+jDO/fZSu5inqjVe7ELZ8VBKYmEJF0ZFFNhMF4Xl/NpMdaack
srZpY3dlciG9o8rHcSkOWS1+V2y+qG66nwY6V0WX4Hq0T4dK2Ml1pp9/b5WoRev2GEu0dZcQQO9U
SoO+r7qg0CBgNnhfv63nMseqwyOLuf/afYNL8yeZdfg1bfPoZ7bXbUfxzqtqlRIPh77c3TNinq2C
+aAtnnK49Vtua4eyNCyIKFCP4d4cNLlW5RAElOcbWY7et+ucQjd1EbAztufZz3oD0SKzjEVG10l4
/G6MsndB7chSD9JwU/wtbzJYXWl/lLdQT2WCfeRzhlWd/jmDP6bxeCZgljtiMujy9irHnVemE8Xc
pBnc5eL5g81QqVGBMzGpfoQgQnDBfjY9zQu/1LGLVYYqhxrelUq6smFVUeubHF6pNkW4ZVDTST7S
rTZpKAAxGGhvBnSWudYtoFBYAurCLlwgZ6jVR8Kv9c0LAszXTCC0XjO2Du1UbH8/I6ZODAooCeSk
VbMW7pJ0eTHyl4qHJUPFS2F3ijCJW+15Fr03Z/kE6TFRkgnEaQUSykIVtjUB9ZjdNWeKe4lkrL2X
dhdUPZ4FT/whwP4gMWG3uE+6tPSmBi0uvF31Bd+FopzufSOJ/tExsC3J+jT2+5f1xQrPR7IN7Smr
+Pd6VGY2RTSp7eUHsZH0R17Xm+3RFnoyKFU1iNq7LeHtn7zQsYQrSWVN6wdO9iAdbHIrZ1TigCzP
p7+t8offe8zVnrzVtDSsiJKUsnamlSb9O5OrFwAjJCM0e3xrdYn5OHvkLcHV8nGW191S3gZz0EEx
n/0dtcRFnjl0I20VqRoN6IzQ1OhWIQYV7/00prmSaqWAVAz8vHwydySmbE798tPlJWOGB+vvthgt
Y9kawtaJ+CCn/SdqWD8TekNOfErLyA4L8BkEhlP5aq0TeTNG5BUOIQNz0li6AQc+tlxjkiMFzBdo
z5G2/ZLn8R5Ll1LDB9lmW5VuFM2O9IpAnmd6nu44KASPeowd4AnauVLkg5dnmL90+29XecIQuVPH
8aicxRexAgYe04fVu8n7PnRuER8X5y3ek3+NzW60T0BbMWKJ42STqhbLDnvPFfvMsHzqJXrIpTJc
cMY3cLZ7fIL5QPkmakB801d9IFojHQ4rVI/UiD0FfzXRloQQ8Hbsm5e1EdcUAcPoGZieVB/BXrou
50JtYNNcF1iOehIu5FsEP2Hd1tzyjw5gO0Y7zTWq8rwC/aPD+/MsGwA6pbsPZXNzRvA055HaXlfr
jG+IpUrVlb8O7NOXf/p5y9qxOyWYn1odPXevv6W25hqGrAY3ZpyMBhD6e9yx3TVoqghznY5SxTMi
jSgkZYP4sBVyRBz+01suHGfBVqIP05EnNIVuWq4QOQg9vspEkNDranwxtbyq0Eo7vM14XiM9YrGK
KjyXKqJTV78krbo1xUTQ1PpXB+pBJqoL+PdsCEjo2K47SATgYStn02NrTItJBhvZYCWJFlhJMMnt
lIrfo8KbWfuqfZN3SIMHbA4d/LFliz0EZzGJ8rIfuOQjqSuA5t4msMJqrh/PsA5no+J3SzE90b9a
sjvnu69fjYFPF5aeIeNg7ZI1b6h4UZWyyR5F+T2ig19MrWgkKBiHy2qUtO0X54V/QHuAs2vFiacI
aIdBKfzZ5jX6Nmt03RL7GrJjn2WX2LC2OorudCpxcHjjeCmQjKaxBfPsSHIzSaXxMd86qSv3Hzz0
HSZrIBBvvAetkRVGAuFT7qmW3zWLdjwZWhNXHtVWlBaldT4JUMvZUGku06NTudgLTHBu4m2yB7IU
b67OD5fix4Hwn+KQSM2rEVSexNMtFumY0aHWSBHEDyY6Exi30+gqBGuccuKgFqEGs+HITRqpzNb8
Z4foWr9ZxFqNxhDQIhV7wW2X38nFm6l4nBlCtMhniUJc+g0/jvfXnd2R7lAfwejUzZY1B3npHaGw
Tv4CJAnnP3T2EGkMBf5O1e3xjgsxr1CAyRc5KmJ+bb4Ft7dYAKAcklCVMMVjsvLy22B8Eg7zVKkv
C6l6AjhL+vOZcDjMwLozUNUttiF7SoThGeOPJgmaRP0UEFt6C2biffwYUTz0YBbbM+lxPoixY7+t
gNWZxVGWY5l4w2qEYDSSHEdFSl97iQu7IuzDEyWj+Z1P2Npu5+XY1hF4zp5RvjPMPwRP0rfEkmzu
qCpj0fd6eTPfF2R+MELZBXajIxaF3pZ3Ep8lyjx0L37fksKMPCK1wAs4yhJwpCxscySXg+6trIux
BJgzm+mLeeOr2YDmMyk8hEqFwFLVWtIEk2PkU/73s87mprYo01lxwDmvLUwM4BymLgzmZO1Hb9Uq
kV3n+Ye4G8dfez150AZ0WIf7kW+fUxCxc7TUCo2OC/KNawxRs9y5EbHqnx1pQVgGGDHTCWR1EWVy
Onb4UfLuGCNHxX1y6xk0szhQf10jn1pnMoLvMqAkVkmbb9ccaVk5KjCfAHQgHEVVl/gUAn34vCQg
JQf3iZxvuGvvrKCaRXAbK+Ai/7y+NobL5+I0Tp8jlAPYLvD4z0BVMj7IgYUBP+pPzs5mtEBNMDKT
iExfYpOyCe3MGJSWdzq80moIKviYrVowGE0awhRH3Y1S74RAj0VaLfUdSstYdyYsP381xjCR0EiY
z56R7amWLghMlcAj/Wu2BbB578ZX+JWsM+/2sVxlrdh4ifdb8noJe38I8EZgjENUT2NiQjPLeWvk
XC3c766dmoGjHGmYyNESnmHVA0mmIY/M6vkt9HnCxwO6N+elIrtecjqPiP0L3ceYsQ74+63XzKj7
0Re2EVHGypwObJHRRlkn+waaCdkQYvzPmSm4X3T6roGBJzwNsb14GWXOswPOh4xJNyWmqbi3uKQG
qbQG7HJ+/woleRAfFJv1Us4qowM8AZK51janHcXBfaDQgfgINB0hTSuj4EEeRg/UzRXTAZtAECr5
CAyRkA0HrJFehnrdyFtTLH8mOZb03sOrGaToHkj4/a3pKImsSHEMpwV1qxrgTrIb2CcSM3gVKBK7
fyIP9pJU/1eQntejQFlWE7m55t6MbaxFvoUv1VHW/oHwhBerdEe+Ndd0OM0N6pV6bPENJMgSUrJh
niopsZoXq2VzEd6x/M9Lg7T6FPznxgn7pR3SX3qOV4mZjRBl80ifa4j/e9Ezgmen51XTKIm77qe+
ZKazjGgrwI++hICCVUUPBBWlX4Tx1aF/2pi5WM3rY0hLq7cNd7sqh8mPPrQqE3AfYkUG/9GIJEI/
kU/XK7CwAFmh4nkdcf2C00xPKXe2O7jAdWpQEpCnzU8FyW+4q0sQBsXtT6ERbVkvqEJ40NSYGfA9
ktccpHm2LRMvNhqbSpzte4NJNk/AaA4Eqpd1JqocM2Jk7FfxRemgsqbOaDzCKpluR9E4q3PDnijI
Mb17qBqOU0Fd++XLmXysxio2Tr/+N5VypsxVvvHPWu2nlxvV0DrlDbICqm4+HUTGfASliOjgAyYe
wfpMnua4CWv6mpJuX6fyuwC6LSjMNQW6DqndBGvHzg24IpekG34VRrWG94E9v+4Pyl1+/uahMGFn
aBIKqz40Kk2B/F63GfIJ4bPxiDPNaKr9I5CFC3FhK3C9EKylEq1k1RgAUJ14EJbXyS4o2TWDrY6z
XTfIQ8xbNsp2K2zsQknKMWl1utVQV3BXhmkISSmc6biwiKPj0OeeBJi332ni1E8s/CSpYjykI80J
JFWoR/mFjATQP0e2k+djpIrg+VVmow5MLuk3Gnr5kALbguyRDne7XvSzscqamvwDMHzSopPbwJmW
KQdLPp0jRU7kPJCvJi+R0Kg3m/H3XE6eozYON7ZFSTQrsuvD5Ab6UtKSH1cvuyivn9yxk/va/NYF
DvIiqQY6i6+ir5W8gc2HASEPhIW4gmDLacqFvO5RKI4m7naO605kCPLv8QJyfisNlL2hV3v+P6mQ
wFELm93savQUgm5k/8v9v6XhXsLG/wp/iGWhJbsHfw1EFLC3HA0uOx8h1o78NYszLCZCfR35G53w
yr6V8EsWGUeBRmEuduqamWu+kT4DX0htxMEnspVW62CxB6Mi6jo1qcApliENOR+ihnSGhSQfEGVh
BEtzPHAlj9y7Ub3rlV6OWuAhfMCPhi/cGwCMDRswx0N+meVsO5awYLegRXaD+T/Pk78xOHT1clel
EVfBT2NKcx4BbRXaEkv4CL1OTat3AFHASrbf7aARafqxf2S7oqkAJk6g1GMuRofSPr1KlGZfdLM4
1r6V1tQo9r0BeOdZ8CL1AR620V/FFAY1og3wcw9YUi/ExHMFI4UT+NAWcRYgW5D200SvKFIDD+px
D/Nfu3H+UFhsZab7IQklq6QEYI6Ggi4Jt/RGDjn3toAIbLbPeQOBALN9vk0EnlufENxWbrWZM66R
VP7C16nbGzVNmEKXEhQ0vcaa4NHcXhF+32KLFdktAZSbm5cQ6soOmvVIIWeKtwe+ONwuzF7Jti+4
MMHM7crhxmcjLa29or5k9sLhieDPhH0UylmNVSNBY6LSl1kyZe5D4SuTtgqIuRaa6YCjMfhvbNHx
aX5daj7QN09l3kYDKfekSuabY6CRMIhUahiN9p1DggWhz4wvmKwkrjJwsEoBbgfgyzRsgJ+rYDkY
cPFPki7EaVaNsDSO7hsJLBOc2C2rl1mBe2hrJjQ24UKgPPXAbWMLUCnM1aVp3oMH/lHkvnVIPjGb
exEHDl4ogLfph5095X0U2g7fZIRY/S+Hq0+eIAeSPAaJCdg4yjwGWnEcL+2XXg0Fqt5GgfMHqWkQ
BPDYUnRsgVT9ySvkYBIQGveMphfzpv614iGoq6hY3Mn+78CEFkMBrwtIdr4HElKZG4eRhG1prtyy
4y0UrjRPn1RQweQ1PW4ky2o4yqVJjuuQ7EL+wC7Y5VZO7/ao+H3oxEQYCxD9fvNcQTguY4kgkBs5
onMeejkXDpsYGYK+x8FbKGLOAfP4FD+pv0VOVFTE6rLaXMyecXPq+vGLGdnIkpf/48/V0fQBZwOY
1bCPRiwiUKcrERRR8mIb45TWgkFqdMjkdY9azxs+OoC+X7MXP7gsWzG3xumcGibNn4wRJooiT7OC
kkdQlicGT3d3mzMO8yBbahquj4hRvZCUpNEipwpGyfbZv5LrSAOcq35C8ep8FAtTpR9n78S5iMJF
WDsOcPM1xoWTrbwW2U92b/Yhn3dfE0MXuAw9UtzR3UC3KEGQfMmhHxN+xFm9+DifYM4AFm4wA3eA
eSzn0eBGY/bPijM8gwMJwkpTbuBWuYsUZ/r4kAGk8o/TupGbdPZHO567m99nYu2hUrUyxaJh3+h1
Bv20bhrEmjJ2lgJGqJxEK+K+fYcGyGNl7En8bsOc4nmrisdLKB1rioF0IqyeCIvoiOh1vVWozUF/
rCzNiEqcWjaenhIbWIQ7KNfxtnaioQsXehON9lrs3rooYrBYhEUQYeoUXazFhI+yqOvx8cG7Yj6N
EfOZMVqYJiWhIhQ1/bsTNQvrtkwkeCBLjufGBdUHoh9WAfDYh9Xgj0uyviB7UuY1OfNGFzG6LmLK
xpiQj8/H+MtkDX24diR+NjAGuMe4NGic+vZRmSpWKmUIsJnk1E4umOF1HaKI2+NKnZOPq0CXFfEU
ldWfytzoEBBTQc492ktwe5E7nFX4+ff0NNVehH0n5jW2wGGba8qrKMezxTc6YyHNiqvsAuMr4ORA
+EcjsszOGdPQLbLh30eWpaYfvKPrEVLNVwSEVbDsymLFjxMqLGyTshjh5lpgB03tNgvcQ9oIGJGf
WNolu1VZF5VoNSkvYICA3gONKRLFPZ11058pQiry+lfZr2UbcU/LwpaaW0Z+mwkRixWbdZwTVV6r
NzhA07IUk3VfGsR6719HvPWU3AYYknBdFaTmMfso2a7P5yRiAOKmj6xbJymkHFVeUQc9/YlMYkrf
4iPtEaI6g1XoMuNJvWPdDo9Q+pQqjZOp1XfgJnhplavYdoPAlMmabcGZgipAzEZ9xWIUmDmld9Uv
q68M+oPQmmh5zW5+Jr6nCgpzIy8s0A9DncHITWvM5s0aDUvSFnoA6Ed3R/CcTgJ7rZl5jDzqB//Z
WlfnnhEjdyBgXOtPtNCzW7snnRs6018kFPuovucpbtVr5fk0dcrE8LIjUh2h8D1LyzgTYN92MX7w
pvqexGQUR0TT3ZytJFEqhhuSUJ+EWV8X+b3IybbakSI4sgKaSC5ZZv+AMxO6hTq8AM29H202ZYx8
MNxJk3qKRVDkcWP2VrAljlVCMJALSkKGQRFvOJJCMGRgGVEHbV1TYCqCBg3fiFEWklW5fxjdxC1W
a9wb41WaByyLd4zEZVwzoV0Y3qlmiaAkavETDjIdnggXP4DbwtiXhf6Uln/HKsCxhfPlg0b+nGx0
xFQGz9Na2KBpGICboKmG+r7YIntMbLGxJox+RNCJNJIIfzS7+fCynDTG2nQP1B99miwZ6NFutwhL
oh5xe6zNRffbojBWKjC2ZB8TGbjXPkX7mNalewCDFktCT9OcTgrcsfqTzH5FJKJ2kpl34+MtkIdb
SUtVZMpdNd/hkleCuz4hBdVMobov9f5wRylaqI29UOZ4bh7KFFBbEwpqWTjgaMSzQ9qEsneYk+vK
tAg8GSgzbXKIacwvLhQFDKJJndEpv5+Fk2UxEFx1QJkW5xydVmpxZpy5FdxE7qgrhB8O5hCuKKyi
8NKWLqYQ3VT4YA92nHfACJjT0g7lfLQh7gANbbUIFsX6wStk8S0okNU7Hx6UXTn4S+8vWBKE/RxF
+opnIyEQYkbmWALlWUfykNDMx5BsCgqg+AP+dJIWXR6bYgi8czEZoyqjxXJJz3TpPrHmVsUOQDFK
Fehb1xuZQAniPeB0mE0KtEkAFPupyQHOh1WexDzzqRfvTOwKjGsdsybFTh/oBKbZlH2kbpRpiWl0
Q+9HZwa8WtWV/9E36c1JDSaLFUWEKSSKzAj+6DK7reSSgWDH36QASfXs07g6VgsbxpVsMZxNtVM2
JYFrGAym7miVzeMMrmdqkM3Mg5m2+ugXnbYvZwfONvmlBwVIk6QhFB2IzJ8amrLJ7P/hb60gWy93
EdqOabqm7P9qunNPMnkiYLDdjbpSFt9Q7l90fQVtPnTQbL3+i94QAQuGfYOI/isYFy+j3ELaQITb
UDE7DH50WwnFUMKBap44Q8pzhpkiPj2NvuiaoNHrRz1F8VNZ7fKL49lxKixtP5icb2Zxr0uAaErg
5yoHU1QSqAnhBkQWwO4rl+rglK36hX630ZeXy8e/utKr6hadwCvmRFVS91mJMHgiuV962c5iW60P
xStmjTyac3dvipsPLAvlOTjSVIxDlprkbESEKn+6fM1DApD+D3dg5cpEXcRRjBctwMo3kDIYAgLb
u2ss2Mqz4gOog+P/JmcGpWuYg1JSaicxw1/nCgP93fKT1cbWUEAYBnCokFpw9Z6fCpZyddYIPcwo
3MlQMtD3nL59tgRa+bB3B+NShkYVMePdqeURuhsKtIrLSPjbm5YUXMVmufc0GU1uVISCjtnpyILj
Up30w/yRYyy+sXaFXRrahd9H7vKiEQjvJMVnEn1nj9MiuMHfgJ1NTV5Fgj+kgjbDZlWCvG8QlAT0
mJlCo15GueOd2tkWg/jkoI2SI0d/qC01FqHHvk6gRjh7rSP+zPPdfegDpiQim55DcYED4ZltNCvw
DfLksI57IaUPbKWpzWLNxPLBKMuZfvCTeCrd3F/zI76Yb0sTKhNAGsrC4YcBf9mNizwTy1lL3Elp
eqOnABKg9b/3eR2oMD0Oc6XyXEJQH5MMFxdfSfX+tC9izy1eXRtnEG6zF6Ncwu+hKMRJ/gjrqGf1
vq3GqfIp4MxUKf/mBZ2i02zvw/qgjhqjU2Go3fwfolYf0O57sxpw7WyB78gf1LzCbjs5wGHxW0Mw
qnqKh98ezMAtoRfeMy3SN9OeytunxJ/ykzPySKGnWZnFHUprR8kMBQ+9zBZ0OD2T5b0LnetD3Mrt
EmAPb2xY2dbBIlgarQXg0FgJwyrXSuUt2n7rkZmkTD7E1+HkmO7re4y8ppJIELedLICE+TWe5UdE
21vyesGdiS+TCe+dFAKFapFhAbqzRRcsdCgAD51tvnYsO6RW5dww11DorYgKvlpLhMud7Pwi2EzI
5RbLfi60lM/zIZgX6GsWnshVxZiOrixQH3WJlEdpOdh4IWSR3NwepW7/1TbSW/va7K7AOlJw+jZX
yaO5zvcNMf2B0yIjzUVyFjStbD1FufrOfL+BaP6rfh9Fw7Z1/ujHQKi8Hdx5o9CTnT1gy9/f3lne
fNLWfK4B2IMqmW7Nddf6l/hH12N2FEgMbv46crMNi8qPtuVSFmsMpIM89lI0BN1tCoRE1nrr+VMx
9oVBnzOUPsVKFdHUiq7e7DNZBdv3wbJ2g/V73kDUgaUkuubOraUzH1YS+6ynr8eBHZBWD1afvtt5
n2eNAeUfY/BwTtKjwjXhe54AEA0UOo7ckCZPivHkDBXRFaKExq/oQmP64xvLoCjScLEDELE+edhU
FpY+O0DMXy50QCunz3KceD7QDhLliz/U9mskfAATBR6+PVPzGPCq2M3dDOUoAXktZ9tB3l4WmWwA
H/4PiGZ9TjxlL/0IZiv/XvJ9FgiLRRrWiUg3tOditMv3ai67BENZiUwgTzTVpm4fDvynP098sl9w
1Wf++OKjHliTvDjOXiH5metEZ/2kj/vjxv3GRBwpsuUxMyX3/uw8miUHpOYmLbsCJZDNHax3PvIR
G5zeZ0qJBcvHzEw/86fQwjNkSGE43s3LnN3dK+qYAwyIw66RxxeINVoNRedJ+WYofq0sCdPUr/jS
amJat71I3/xTnTsayQ4Q4mCCYguSxHnE8vyrQPdERemBuxqdDOhSI5+dOP1Qtp/v7cfhpWn6FEKQ
ZumvVDzLpvJ/gHJRRsNTYaWe/GajiVTIl2cHXNTZKqGXadU5yT06jaZzQEJQcO5WOhZJXY6fJaky
pGpMA93XR7nBznJD9CN0OruBVGvoU8cgCf77UJaUksvwKR1CSpACdQn+F3VMah8A3vo3/SGhOG4U
hIctAOTJGbl3wiSklDWTRzNIEZi+rs9AC5VYFj+TL7EyEvuhVFFPVVKSL0+2BeukY6bXyUCLnwKE
cYOzLa65tFJLA+cz6HQNRa/+E0EOKvAJGqfjVQo7l98M9VHZXOHNdfHy0NdnXpa3TC+yiVdF6lkK
3ceEkrLw4E3CJ8z6GOfQvyjxVdCxv6Xw2te7x7DBFGjzI+S97jEJlkvk4XRYzhma2vFhfLle0K1x
3jAbPYsqRS8GNTAXYNB1Fbiu55g+dE3WJv2/M738067LqdaiaP2uyXYROyeZPN5/Uc+nWOEHnu0T
0sihweK5z9cp1Kw3L7c++J6eA5uC/lGIOfOwFflyzONu5LErELzxpjFn4HU5U5Kf9y7Ivx40G0aw
oiehXsKaH/JS1QuJwkvg6Eim00KMFqQCb/pZ7lrmQ2JIOPjeiA0thMpNE1PIFW4xWhlggcwxbeqK
malM1x82Yc6d2oC9mJeh+xwxp6vE8U//7H7fobqipTDOaUzInMZq+V4WVcc1YlU2s1T6OFl/4xJu
PGGHFIvX8eXrX7U2NjV08Sui+GHBD296BwyuNmS86b99VyRKoj6aIqPSUs2T4dVVVTvZpCIisf7f
lZrVzU2tHAHmbpoU/yzpZXbzCTsRjNqHy0i7ZNhcFDrmyCIrhZ8EK7ldqehigrz78ejNwebfb1/6
cUT5lH/9rNawJ+GQjRfSFnvlt05rL3VbTqusNwArukEIaxzFNnm+adumTKzHkQFcEfqXA2cENzfE
J2q39zLaDrTdyNf7c07FjEr7WSnppUsKam6RG/9u+4auZ3p83Xm9DsLuvHKb0C1JOuAi0gjxxIpI
Hj7s1Z6vcrhM0zYm7jtKC8f8uXQGsfVtA4cDH4+urlGJ0Jo+XC8wleYGgfihr/wupswibF9KSnAE
ArLjsA7VhDUe9PdMzDpoayqcLHkoG04O3UcDNWjVNEPDtCYZXJ2mlIJCWdg3FykED+d+JzAGJh/o
Y1bEbyk4fjFkGxA+ADdYfKj9D8wbd/jeRfBBaSHhFBu3ddYSEpmru2DspbxojoQL2Nob6IZ90998
r2oLYI52uY4EZBwuaotp4lnGEao4ous+I8vWvc5As+91TeEanZadgbJ/69q2LEeWGxfzGlBvdcmC
/uZsOXkQ5g1UAOhWc0QGvwBw6OKoFxc2q8psZcfAKwMTPk55HTXDGo5pih2c8n9U8WWWLtvI4XfI
WNtAjHTJZiX8BgeFtMv49/wRBEAoEaSK5mr06j8AyF0bbl8XIVj8oXIMIIuymzqxDp4Nkv9vpdk3
puEDvTKkAIkip/ctWX/PNAoA2oaKJ3LWN5y8q7DT+fsMb4wZUyg+X+wIWhA91jucDzUUXq8FFh7h
B1oL82Sy2QVdoHQR7yxX+/lUVEwbn7gTzmxKAbS6ZqOQnaZI11nuJprKFAEDVS1/QOXCfwbTwTQ0
85hDEMo/j/kBhKjl5kB4sxlQOYbsRMSVUX0l7lKbrVpIeAVlODmH0zyIoQ29a9ZE53BuyZ2iMuFr
JM6f36M5mHN+mYCrAVofdUSy3zcRg2Jp9K6Ij2Q1jTUCsXJxnKdelauOHLIMWiLFWFGLhXoSPkVM
Qv0NMh0sUqLpbXb75s7JtP40UtIpmNzWVg7YS/tUCiEbFB7LQcWGbk08EqGfqzWQhTzLaH/r/kQ2
Ele/jt5YCu3+ZjhIROBaCppZLDN8dIUDzc7mTrHGbySTzEcSWjUYmXl93BN9XLqe053cr/sOW7kM
1DtfSms5RF1CFQVVgtfftVh8xCrcL4Xwxdjt8marCsshqlA5g3jK2VQfyHwU8A7Q+l/2P8MtQX2t
+Kl7401Cw6GsnimawBxWhKdqXBjpVilvhHfo/oD8shnpk/rhaSmgvi9FwAnSw64vlo6vBrscC37V
KuJX884zhB45e/rxG+1MjG1P41ZvA4dn8IxBNhvW+jNpRand/h0e1kGFPULmbT74SXmJKc6u6KVe
kyepjEM74pV1mqF+BavYMXFCH+DCbou4NCahxdVsylShHS/qJvWR8ukbGGmUkSJfzDpxhOZBi+OB
n6aCxzRzC6cxXAWvjs4bCm+2pINCG5S/e9UFO4AMcqViz5waBogG7BKVlZhI7CDg5NhjBwBQQaW8
zCzKZMV93UdstkJEeLGedWx7Yk0ChtNvUxvL5UIOnF2Wn4v9bkf3ApIi9dWoxA2pJOeLvyq2Y+aK
ErPrJw2ELJFTE6eoVp6Aez4C+MJEg3eR6Gg+5opd61YKw0ItDZRXpzH5n7UAK0q/I9ioRNCSw4V+
9oOZQF4GsCoFkNtUCrNH3S5zIqLYhssemaFqjsB11trdLkDR2qvsNLKLbp9MznejilCvIjQyVA63
Lb18BPq8m67DHAgPlKIBBrDEU2gppH+IWmY7ycd87htcbgHw54gvlECpthvHP5rdi2o8HrsdyRPs
HWpIGpLmyQ48Ad65Csj74DbZ0ZlMBB9SukLHP8jK+5/sFdGG3gc6G0xPSPlEq5gPCD04HZyNQ0oY
naRJP9jFzxOFVFVmcJ6EbWIUc/XpgYszWT8ijFy8t57B+GOXqP6BDV/rfLndQbJkHwGveTE7AXCy
JalaHKzuZ/3Zl/MqKq4LvTiU55sKYLqGFo9LXmwnLb8X9YeXYedT8X42+7nX9scjr4dpt3qhyMKY
e4ILRJpdUemxyXTEk5s5h2o30fKWSczitskxP3hUpj2NMv0TpkBWQr8E6HnoRmYNnlJ3VRgsTOye
sDnM5sTYBNwVYijJiJr4zKB1KgiWgyBkkd7CH7HIW+KFr+BI0DlTq4eIvay6L+dmOZBxw2QcQqam
0yijzDzj1hZ2+0cgCeuWgTWKwncH+khV3sbH1Y4HZVp8NvnA9tOHm5iLHcYdcR+qicmCm++LpiHV
i7fKb2ZQuoaaQ33Mu8N2ckcWyTklMmUXpGOatEkDG6jEyk6iusme0PDcki0HXe0X385+tZQXUCI3
FrGONIIdosMU8A6qKhtp2cdllqDpUAjusejhMEsMfvYGjhUGHZfx5o/1U2kgWtagB1+wveN3i9RZ
kP9oRO3nvc9y9uqn3EQpKOSt5fWKaeeaKb0Zf+CcGwsql8c/ZQ9mTHvDKtw4WxMS28kyOsDQp/9N
mDMc4CPmirAJXA8OnEQagKrpEGCiLknYsRlNVLMqkoCtMQtp4MuyQ7WmPCzJAWUfw1jy7aighuBC
i6YpLa/vwb9uX7dfn+7sv6ega3nY8GFwh/OawUYZtoyT4uh0ePyhvukYlWrl1b4OAIpIkuE4/dp6
TNxVlBmsOCU5F/TldPqMOcQ69kPAT7sOGUopAhBf1h1LRR0AgKJyILFKub85EpbEr14lcbNFPuep
BfWkRJZsIq2cfwGTHuzjiRfTJhPEFlbbDMCPDZeJLYEmt+tTsiQN63BiIAxoD/eSIVV0gheudVf5
UNfzRuTaONkTf08tQnsS9AO6Pccan2HZldJdhZxG3SlM/GinlnnDjKRLmGTdoIwFOiLiB4P0zypE
KRDnef5P6g7OOEa6pZX3B82XPm9aS5PgszX3dsUXxMF+2uO9uFDO809M+cKCy02HnDgP6sbZB2IY
ZoE5wGAOmIEA/lxMd3vtxiwVy4LlF5tW+b+DGboa/HzZvDmMoRZ5YnuOei/kfGVMnDUMlDfO5X4S
DCzDXrNs9w7GuuP10A4AJYSXQxjiM/UUcSwwYHEPS+sj43/QQXLaiqz5+FDLFO9RgQyeyp6wXXni
NvSfhu+kZW35isjL1AIS+Z1w/UzZu/ecrcvZHQYHid22DB/1dTGfoDu+kv8j16ZDtaDed87nfI7d
tXdSyFHXUmmgrB+8Rt23NfN8buvjEO/i/KHbzk2Aj7+aPkUU8RjBKYhrx87wQdEF3rTxghSKc8/g
+lv/XEy2tQ5ZlqxfG89/MVeDfL5u4HE1nviShmtMFPZNn8ZcRG+7D0tTqAtDWfPBje4HoGGQagLx
yoKQE4GAm7TB8vuRF7hoSQay1Qk3NRwqg3EdXx0ck+gTSTkFepvaAA4RgdalsR85eLQ9ZM00bVKf
TVOghC+HMt4zAzpQoMAS5Ji14O4wsUDm7oWazAdgmv0kHMa0sngRrziTNEqSdcllDEh91lOJbNKL
jQQwsOc8O8wAKGwNuxiSTDDPzrdp3fUHW+QyGMerlKZ/yhaoqGYHmdYzAnNJ1tz/C5F+2GD80RGN
jQPFLBCLuDGQGCSKeIEiYNnpoiVx2KlgU0l5m6t1SElTY7U4O4EKQOnFdSUe73chcA7Y6CbsilJG
TQ+EXdt8QQPpU36uRV/Rp5KCLAvWDzLaHHU+eVtH3GMiXNstVT/vloBbAIr8Y12KahbZQcqVuS0U
5XfsF7lfMw7q0bpyqe3gEtH2AJahsBCV9TupDOG0x7H2k2FaTIDFGhZcKvsXdgBlSIG5I0N+OrPY
YUIyxcCsUHmiisnjwj/uM2F/eGhweKdL4ie/qFxie4N+a/A+9583GPN/EmtM3vk0dLVnWkDzbmuh
dH6Nm97gx4UXI9tCKjWRE4olA/3FfnyOgaplsZLld+tO4hKK3JjfuhoQuXmZB5lopJ1BEawXmE9Q
irRVcXGRhr5Eeqn2BOZm5nTg2M4cmHbA7qZibt0xtpbqagaWwRQTnlYAviwQJQH7nGZR8tCCnSf9
CekGJiL7nh5Ckas5SNTuqXyE5sDL7/q5dh7iTKguvS2Hsej6dddbq1j+j8aHAaJG0ujMEIi5UCoI
PlYgeqOvjIsiP+FIMz/ZRbZuGLlNdVnF4d1Cr4f5sj/nYxa9WVc19cKOlhf04P66WFpBCdq7fanF
X2WnvBqd9ZvshTX7zL7P2rVny469sbymbHsdho/x2ba8heEG5rpDL2ah7MOocBbbq2RJMlanX6St
ytrTM8BoqAwWRYBYcozYNrD17j3xxZod7xbm7HuSYTK0fQ4Kr6knpNjhqwua0hF0KcUEs9K3PWKn
sqsmr5YRQPMLu5PrXLIjiCrspkfCXzvONCcbeWNfEUs5C1Q1zQnmbgBPh9tq1xqdkBZ6ncO8HlV1
o4UzIX79WPY5MbKVK2laVlhTDwloLOwdHxxsiT79tj6Y28LFaiYY92Sa+982BO5TrQMux3wxW/9h
O26ExaOH9ZCUPCAEAsJV4oU/eMcb4jOgdm567iJMZTF+wNYIP5cBHM/BhDpv1erffOfTImikqsyr
snfK0N+iwwMyGLm6mtCWE7b5c3NnQ23yfsfyXdktRhxq5nGki4n78y9//Ee/48gngs0cQxmjx/pX
AnrPIPsbF6Aqy00nff4MM2X/IcDDzTmX2B0rHXWHhgQqMc8Rh4aEDJ4GJ8ch+mXzHp9AGdZFQjNH
GNrSRaGlHF6fmmJM+xLj1+bCjgeh8x5VWaY9K8hPFEr/+5blKE9o8/8IET5kVdDBYauEcXN1qD4I
Ci9NJZkAKE5HHm8DeiKzK6ussWCy0eURekF5s073bKnXLjYM75ulekgf5qtaJrb7KKiqBU9nRz0o
Ncj18W2CpVDcpSFpT+Wq5XFwOizgBd9f8i1z2uPK8rt5+VTNopwwiUoB0y+XlcrKSfQWd9Pzc+xS
49qI3hKMJ+iW2iR9A8YfXEYS8O/K9OM/wvWk0XjNLwjIOZtHNlZaO615eXfHH1yv6OdW7UYeTDZe
dolHc6PxBu7CoOxvjq20nyCorv+qngwzDmm+VMaCoLuwRD8zuJVrsM2sl19uUdtuaLFmyAuKuhvs
Y4/PHLS8axA/RSSCZHgXctnTgpoHPkhNsYzZj+6GB9jzZz/3rZDXjlDiQh+7Xwiyx2WW1wbYr7N+
ee+qPbWh2DQgqdQ55yAODk+i8OEjAwyik5EVZTpwF89xOJ60wum2k78PUXaCR+Kv+2uQcZTEGREj
0+tQueNZQTlxJx+k/HCXVeex7ElvuzAOt4eyPItOcLc6AjE5U4pgGyFdAdg2hHjZ0unPdWOk+wta
mvtIlUj0mDZrpsbOXc7fBd9dZsVGm5KczcIWhHwrv4nGd3vsmhtnbWxxb8x+BNe0Q6UgG6tj8Jq+
t3fDQTkgZb9nfJl/Pp1S1ODalyhh64qIv4iRw5efSiILy0fhZdMRP3kE/YcsuCiGpaNC69sy5CJG
1UU2ZDMiGEXgR8MvhjzxcFbJn2L/Q7/DWeetg0397g9Bm8r9nlwwGXF+k9MGkNrYXHup+xB65SnY
JrpoAk07WJfKXnWwE+tOKdkd7WN7sEULKtEmZnelZLKDDbEc7g0YeSmsDlr9gHo72zfumVzlt9tA
f5CovUv7Fs+wgt06K35oI6OOVr/BdyTHDkr9wH7LLumrnfG6ei+IftciS621HawP5yjc9Ku8sbrI
uRYJmBavn+LeX0yQPz+PlbZZH7QqysXeQ6mOfRmFvVno3zFeS7VWrAoitBKAxjjGjXy4c4qNXmeS
Jy4RUuu1qXhxPB7WKba1ThlVhww0b8pQOQDBTZMjjrCDaTVg+KixatUCooC+Srr5MjAaSaCEicMB
rr5IJBc2ew2qRgIrbUgFWwVfAQB3cI7SvrweGvzxE65uVAF8yGzYxckuWvQSgAingUnVM6p0aARj
k4RDSuWLcmhDinydDdUIBOp4+jUNErf8CGR7EyjbZGkFkI/RHM8Q/bmO7LyZecI/N1OtDM0OiolP
mv6K55AJvlp0MxpI9vQCPyTotpr220KlJZzWKiTV1POtjMtHqjDJ7y6S2LYM8LGVoLy2DDRHJ7LZ
/iNz0NkU4El03n2m1lSrF+o1iCmxRsudHZIqrMHBXmqeYvxocQxLXI4tls/TpJMqg34wnZV2abq/
2g10STE/zJidxYpabw2gtQ1f0Dy84mRt5hCrPzuf3vrn4LIsa/ebjW3/n1TYwiwo9X7Zk3jd+JVA
vCHnIkwWi843thkwSXGvQDUfxGGFBIsNdOM7s7MuubDn0Jgyz5Q+Wh8FSWkZCDUjhP+vUImV+1+L
RF7BHYESCRTDVuijzi+xEuT/ff/oV8qq5eXQ+nBrF1mU/lfHaROGBVCWF/0WDQlfOeDfpGgdjrxf
4OOV5OakPikhyuiAH2T72BcJRr7/EBPotZXh2RdAVufGaaRD1e3DsjeJ9uEvjRvIyDU858A8pKC+
5W/oEUOmhQFBByXoDPpzeg/F/y/hGOoNm8xFLT1H9yDNZtPzbA54pPPaYY8SlvQ1LeynhA6H7yQs
KHoeR6GdqRsK92lN2hMWDTz+3RyvAyaQrZl0aEm0S1KxLZYl6TfUx6WiDQquNx71s1r0TOX8zlFc
8Vx1uT/2LyyaTnxJgfIwVoZ38TPBYIyKV1GuRzz3R+VaaQMUMWnWymcd+azrnZl9tEZRxOTBe7Kn
cxF2k+Re+vvzaHTyk3MSxoJk5vGNqNTQWXfg+pxeMLjtHFcnh2G/kFDJ8KARHUNfGOFUlVNzuW7M
AcAEAdSlmxz+dQxQu8QgimTrwcIur9BHp6Lx0mwqCNgKYf2bDsvW+CWlRfG3bG5s7C3tHXcQUpMy
AjYP8veWuh/LlfZCF0cBJ4X01Afa6DtzqRGyGeoz6C9koJJYUFkHH78W9GZU1GR+tKNOXhEGoyuC
8t9T/zGMsch4ZnQR0X3x28yaY4qSFHXw+XnqmRsJ26yK8vG6M2uMQ7IdV3ZCMpWaYitCdLi6C2Xk
0LTZaEsTkBXMWa2VAVDGaY2ghWWaYFMwUhaprvR8/BYU1DxV4/jzuth+WQWreD719Yt+j6F5JIJW
s+blJ4BzaAjMSKUs1Zacb9hWmG2ijA7M+pXrd8x8uDDVN34YHwAEIbkINHQRwgKWmmyOSQcGml43
zMaZrp4fbisV8TZePoakefKwRIn86GftA7Nqdrzpuf+Kur2tN7kGzfZuKoxrDy3HN6cmRFiitJth
lHzS2LqeQgXTId+bOkaQJN38e3M9EggnjnEZxWnFpU/dmSFqxR4ve37cSanSYbVuf6zlUNEmc0bX
alYf5PDA/jxbEHufhPJ1P3MK06L7KofPVnq2+DEiUuD1D7/LxjzWL0Sq4z8WTpVB5dveA305p6U4
p7ATTd9Ol2VZ+T+BvdJdDqipPIIRqMkMGEQ2WB5+8FizU4u8y5nZA/fQ9xyyRONrCJ11fGMWmCgJ
ane7IaJJP420iGlARXLzk2Ox8GmK+OLMYdY6wbfaGNefhDZFCBW5ISL4sa8gYvHKbgG/jFgx9qMq
U3kLKWNaTFVYBkyESjzTkh2F2cQGiqWquD68Gdgvuyw6Jl6XvHrYyBYlmdBZ2QAjlQNT5jXsjgpz
p530sCmXkVFBc02YPRnXUu7WQvIVw+uRiarJnTI22Qzlr+MCVyhJCjEVvxVDGX+YGIhGJKIiOkqn
490Gf5ErCg6I1rsYAs4vij+Wmad3BF8B9rmswxuH+tO5lroDw3HEkGTsrPTeA7FbNtNv74IabVLy
N7I+04AVnmjGRT90e7+9L1SY3Mii7VkDvhWkmQCLqyp/0/djVS0yJiXxx3NPSq+t95ciYpm7Qjoi
Akk1zlvbnnMFiWfWPnVMERyM06deObkvcbEQ2BnSu2O8trp2qdz3jSuqJVYUl41XP4Rh/PCwOBHg
06TpJvJa5dgj1uO+2Ihzs86H09OoQu9z18Xys/TA4JqAYUYaJODyi2wO9Qti8Z8aSThdgNgjAilK
lwHB59I9JRuwPAx214UvrGtPG1B2BSQ6M23I6hxq7rsC6AM0rgVb3SW0P0P+tAmKE2U+7UzprNQw
tjopAmD/ebMg+9CTUd2XB6WOHB8KK8rqTS/lZ1K54h0sidzN3Hr/8wErkyLr/tQXm8ahI7zpRSUl
6I57KuuWmHFF1BjnYfCgLlMBn9f3GCQ8HWz2sd6axh7NKROJSfIioAIEHuVbuIROmAOWVyQ2eqeg
24PL3dPF82qo9PCmppv/kL+6kz6X6Q+riT80oWZMLs337Wz//v2lmV1fDygvAZdJ4JiBI9E42XIc
TX4J3Yg38fPMZLMHEhOVrnGsyqhqCWTvb6hwjk30GbidlL99xcaOnciTWI131QE/YYtLf/1aVnUE
dspJPEXMJMdNtHYQrZ+GPExZesLcoxJPhO8cyomm/Ho3SMAXGbUsr/wys1Ok3Wde2nTzaT6MlnAi
CuG3edLuSMTD8cHnX/ai1bpQ5XvViNkpKRzbIiqu5IYCAO8q2+Zb6koErBtu5+k108JDEJssxgPU
gBgOPU3Gl9B3R+I199yedXV5VeF4lWp2wB4hHmlkDC6S092IbVZZ4KNAcjrgaYvViYFwpZeyueDh
sWVX/Qr1KlHv00GgsXQtIfc2tzimqr9snSvsB2RAV9a4/iZUSuKcAYbJpIbRoki3xePW2kskQwkW
punOdj7b0xnHr6rCtcYJyJa3xo4Jn+nYgLRH+XL5k3ezjc4zgWfo0MhaZx0TV6fL75Sb4FGfopl0
SRwCN0q8PaODVhdcJxHyrBlhhkaCdfvDqBvKI/S5ff20zoKMFUHQZPDuD1RTORBkA10jVA3c/KZA
2BZPrqFjoxLssQMuDDi3zL6D5OJMAuRYyCRcu1LZbpXNM2gXe4TPncwDYa4UyIQgHmQz+HSrPzf5
jfDUaKfIuB3hD0+IRYgBvZb044aFLnwHJAGiAGgBlHOEZILBNa3lYAxbOUakII4cqbTVX0gOaJaD
wgp4beZedaPtK49NrWz/Ox3JvkKbU0KLrj4UMD7lyHyk/D8lWo0WcLZxPCebG0t+loehKIEyrin4
Fl0vQ4y9sAumAjpZL97+xnL2ZOVcYxJQu0Q2a/A1sQu9vEjEjw8PZwX6qRxiL8gLGsoDHp7sXGQg
zoaMcRCcFlmLyhtFIbDZhO7vsrsqjRsl1Ew6kdb2+AG9Oc2GO66sfuGrlBXHf7AlkhsAS20+XF34
QwKA4yRxY4ObCjudGqsIxa4wcciwQ2g9RjefKa1BDYiOVdj0KNQ3lqEDsKHPex+Nhn7ULeVn9drF
4uITkW6bAdS+SLW5acxJIaEsu4dkFNLoKBrFmsUQoxtyaRnSN3x9ACx70EL6mSq9FvjRiMEp/x2j
5o54c9eJqCRyhdmJT7WId6RQAUYi1LT0jiJni1JVCoC4tRSmxXRWsfca1/cARlpwyNnlpdTqWxBB
nrma+4PESAceOef42VxV5QuU3qf1lFf786U/ucPDhaa+ecVz40lgDwOGCAxJ71aXCKSxsPrR+8ai
q6+1ZyAaAoywwcm4Opu+0iKuUC0zwX9HsxdrR1PkBqagSmDx0eYyVdRkhjBtUXuBoJKdeKVHjb/h
OSZPqkQAjn3vpx1IOFE2OkrIJubV6Z0wf7KudokBPUpLfJulpr4AeSrYYflVz+yNyzql+mHPIbVu
52K2N5GaRynCS5D38WA+6hPItc/Av0/D6huElnCy0MGRQVUvq3j/ICq9DrldiQ4hQ7anmUgQQP+K
qBOIa8tZj7vurhDZR75GauiTveQwTsG5STFjZ+xigidoWhYyMq5tSmjJSQludzDT7SGqIzzpIQWE
bq1guoLGCeeVtIvt7VHmyUSsD75ICHm0xZ9na5WgMKKZUB6dEV+0yKOhI+9gNnNMT+FgEvFUgEcw
31OlNyjoSbF9e0zFY2FKrOt1fVLCEOK4c+gqmSRn9PZ48z74O1fkjGMVkkTlAt4L2WMNQUhP8ksL
z8pMM6UxGMvZLRrxOwDDQURivuHQut5PFZnc+YQMYR8JBBhpwxNFMIBLF9cdpUudZwZxCQb69Mn2
r1C8qUzYcKnZmQ0rLntxnd9uYqXKZmG/GI6ffoGDAyzN+Hxj9nd/2955n9piVzC7/9n8S7uC8nsE
Brdp7jD35YNMJ1+vaHhB9ohV5Drsn4FKF65K3POLkFAZ4UAHl7j4lMpGKsUAFWJb+JLCROoydF9Z
5OYqIFOaVX73Pi74sbsVi69JbB/v7YXwp1KdsqVQpMt9XHTYaN5mf6VwBW1BW6jJkYXZ68ebIbPm
lQBY47U8RZVnx7I/ZHylcZ6o8nADrB34R9GBmPtlVWyeTs9x2jo9pAIwawAw8x8WdCixeHxp+oWj
QFDWVsZQEfZj+zbCHsMPHhVsMlJlax0IEP5JyyCuEtJ4XEg+qRxFNf4Y3szCKXIHQ+et25z35RYM
XW4FRpg+T3xPDHv7i46HwB2YUbz31sDJ1xXxNRhpnyifOGyq5npT/37LX6NLDIFyoktUy2u1SvkV
Ls1659T4ddfWHqjJg1Zo2jaV57zdg0fabTqVX+dr6+LIVkyv9+bHCGNNoqpnpmFbRrds2cRl6sQi
6ClyFL0UURldVfi34MgyJM640Py2GQvlnovbCad0O8vixZG2fXyoJxRLCqyJmE9Q84ASNRR+Dlln
qTja24jaahKefrFovQT2+xU5Q5Gj8XhIVxqG7LIpdKx123GbeG0a0BIgaq1I+Pk5hlAi2aEzBkAT
gDkrUM8C3SA9Pi6kwfRatwZkNxuAQU7VwSKeQwB2rqPXHoZPi10XgcuAmyZiCI1W2YrXqDnzOxkp
oXorbFA9OykP0hoCRMORfTrxQ46eiTLBV/FXUAxYc4OTlximds7anRKmnenQ4lTq0J4/iu0ahSTG
PdHvemFcBTwccikLr08Wask5TNch5urxnWqWpIshenKR4C3xpfBcra14tS5R2vI9qJijVE7k/7Ws
YIkRl+T/uCbypaevB76kSxTU6pStWkDKlVf4cQSHO30skK1L30xu+Yaxn8EEhZVAZWiYGGazl09z
6morRTfUtRKdiJKx9CM2IHFljKhyg6mBCxfyAVLN88a3OVy1FRmW7tVvsasqAmMSTz77P8bDw5zq
38/JoTdJDlLXo3z504swQ1OSiq9HMFq8ZxZAwwNdR7Lhe0j5hqeooa15xRFgSp3uYhJCug36mnSs
8kxC+Xrp0A46aWs+PWeV3eTNNmazmdTu1jAB3e0dNB4vgeJRItxJfvwtwAtpQj5SGnoQaGdI6na3
3pKYusvwkxdv1X98BiwWLAdJ6c1KtJ15IF/VbZvx1YacHxbvPmcfMRooWqybDTPnGn/AQrSy33FW
AOE30uN1rVwhJIPif1pWR3a19AeMh3lptzBZtRwkeT0BPiWyS2Rll27SjpIHDdqDhdPg0ihQfpsj
1FxfArGc/if6iY90qw96UgbLRwSpY1LiYZMJEbwgq1E8+DEPKvdCn5BvizekGf0afXINgzbE9BRZ
5fwviZZyY5FbSi9nnkK+V1px6nnl9iFX595Y5hKQyDoYqERVBsHLTdAOYz5tFghZF1UAIzsMfk/U
aE+dw6vM6LpFfsKYsuYqjyTR3hHi22n8QqmTAKg4cFpBspO68kZADKS+aLhZaDQVm5II6SMUamYM
cY1GuH+gyfwdOb7qDpRU35y35kiDLWr9pxbIsgvnU2k86Srg2jwSkUJ6PWTJBs2d5tfcY6j4lJhn
7ewOLmjaV7xgqcDeX6+7XmeHlkXkLbpWI5DoqrSfhGHxx9WNRunS5o1GXX8T/0pi8t3clsaYox/9
yq4iPxBLvCEC9o5FVOj5/LfFrpa8nlg3anHxKp4722gLiphRn8JrBHcaX3rRiPTwm/HwVpwOv/DV
gTeHMPQp16CwiK2Z1UnMeHnJmIg6PdcJX2cdzhvJoWODsDDohZmgM71r+fgEKK5dGSohPRFphWl1
QM2gpLCoJqlN1L0aPMZ9Amjqp7tU0HT35CMQGq0XuxICmmBJkVzVphxs93IghNddbXWqj1QQ+1G7
3G87gm+Efwi7bWHLuRuqgYZtLJtAJs23YeWvSDqflcfpA2EMJustjjq6xSfXEYIN/MK18dXgERiB
TguUL/CNUZVd2f+fdg15aBq5i+sMBpW/xZ2EQqT1FiUGKdSpog/LMW/Tzw7n6iedcDtDseLitxtb
kccyfHhf0o5V9Ox7b6J13IbBW3NHoav4pK9AjtshCqB49I7yVl/tISzFt4C1UvnLt9y18fGUFY1d
iyveHb6aQBQuBe3mVfjVCuFs4jLhkgzc5yCnX3p6lRch3zuQTWYgt+cSmJSTa2Rlo0bYWpYWbO/L
6hxzfuAMfIE2cwXVC3QIZ2g71zmUhkPGOv6G42IiuYRAaZ9QSmRsban3K9cKb6TrmDQCfERa+rpb
TEidMIWsqjGT7Q7f1sH9Z/2TCgTVMcxkZwedyeNOWkfNHskiUZAxAF7djxlZUJCn9tDWjdQyVq+w
o6PGR7oNRgfyZf+kQcfIInPbK8F3oUDk+9ntAL7VR9Du77slFGBaLEnd+0UgajLFXi4e3irsgM32
qkjQovbhQqopBvGdnaUsa3cBW+CsgFNRcwwj1eCqzhSCa1x9iX8iN3up+qjkhsL5QDhs/OFich6C
qSflkQOFifSUmI9k/zAa8+sVtKjAbhc1rFdkgZq83Kn2ZO7AyZ9bUKcfoyzDv5Ok8n3OjnJ4cI29
8g8WePU7N9DRarGOvXSg/MTs8wq43V119HI0sPzHSlfFDpenZ8DJMbX5LndjEeNiacQp0GvRg2iM
3PGx/BgKuRgcJqP87T351CQv+ivq+TNfoeBaICt/vVLI3ZZNVqoD6paFqZia4bYGUmxksmgvdtnJ
h2vdHW5AkfSSVyR+G1pp7mSbmmasxFvmR0il0/tAXe+0n6OnKQn2d9+An4+6n0na+/aF6xlXDC0+
sj3aiqFfrpT+P6KirNXHzDmC78CqKpe74JszLJ81ejgi17OgrB2GWZkyvDjFEwiMovRcZSI1VaB1
gFJuWG0S6Jhd1c18suZzEkI1FaYWbFs4MnAwimPFOhguBOKk8mYw32mRGpORiP8VATjHaUmlP+i7
MfveHqLVxVZ1OB5nHj9iSLdK6wtZf/gzYa4588Cm1dcTF3CFh/54o4EGIUB6kJxC0Qfxwk77Zoza
cvj1rHX/dgPOlPPDPPiRPap+FJtcBD1ZKWCPVi5HbFKS9xpklXgBi0SkZJhxhFVGZfaDtMxVVBvU
uuanp199VMPSiMIhdEIB4t+mREoifo3YJ9GfiT5kJNU5IEz7Irjyi1rvfnmLmAIRX96ICeDysTe8
eEoRrZLbWsKJwntwhN8k+ycy7Vxt4nEXCOoUyGYhbXsnRV/I+8D1uSxqXOQrhKklqr1roooAx456
WACMqI5masY2jhUF1h0MhDnSilYDglMVZHFV+orrlFMUjofvyy3cEWPmZI/JTFTTuRfn8/9E6yuu
gRO+Zlp/2K9IHfXiMHGBG3vZAJHf080vQ39RO3nVbWqgYzGeRcn1LOfr+tydi4q+T+4g5MCUjVap
PLLsn9EPrN4k3wrban3DBhjsoEBScftTHDQsmaJLfEVhs17Rn3pSyKAZMsGMxhp+5C643NoEBFvU
BZFvI7gzJXdbtNldJS1d5BjQHpH/4+01Ig7Oc4ixwMaxBQy6tt2NIUehPZI1IZhGEIB41kwHGq1J
AleUMOGFnY+XuHGWerfP0vyIL8L3WazTWGfW2BwEA1cA3ZIUV/s6lTcqeZOX+VC3Jyk9HfTerae5
TaQwP19dUo1FOBfSRi8teMR+VeyavpaOirSp3XHrN1XxJWz2uvm42NBg7K8DCx+SWORHUFok3ms2
3H/UOXwyI8C0+UifgZq+Iofso+waZg0BdM0ryv1DvoLoqU4QCswLZ0JafooDslbcHjZpUfgHRYnj
NM6O2STlOVyptRJCCWJaZOiricddXMNtAH3kW6oU5Yuek+0pJ9AT70m8bReZw2ExHGd4hRcGB3x2
stDyfqyZMpd3lBIBEGqE2/IHSAgJx/1wsFv63GPDTv9l/ftDF+gEUr/b0bFefPIapL9/xBmXEgGk
EUL5dusqeC4KJnjznH/yfKSJ3g63smAplJ9b79Z3T5k/9YowlCz/EvD1S+c/BvpXE6Wuw8H1CdiI
7BPkNU5fCZ0XH0bzeStq/2Bx+hx70xUxeZgL/qtkiErJpiw94y7MTQbnGN2x32ynUN3CjQd8eGvu
61BOvyJB7nAa1jWvm9x1BEIxl1z8aOjZID96MbxLM5mvD6VAUKythZM3rrk16K3RSVzn7DPuUR6r
K5+sJeWlECU6Y3vtQvRXKnZsvAo4U+/DE+7EoQ6wBwgQm0Hi2dm0At31tPlafGXjQ58JaXBnexhD
OlXYDzZtYvEQd0y8+L8myzwluTCdY08rHPgnl8fugBOLrTU1H6jKIAiCuNg1jbiQB7NoqHZ+aOH9
NI0pakyArZDGS2kRFJ2kEoWEJh+15a+omGgQFN4zSCsOxAXyLaktCXqOiunvbd7Sfll3c5Q/ePJX
8HeGUFeWrahMRV9OAYc2URG06tMBXuGcFCTRPA/U5reJpnAL/ZG28dVtcCM6IoVqOIO68oDSi/AD
WNb4GtfV+ZpVThEMCrwGZQz/fzd10eMZDcyqwW9yqdG5nApCX6tmvcmOp1w2dNF0lrldJNPNuloC
SbiHAsHjBR03IgWdL3zwVBQa/SyTuYUy7jAgn+o3z5a/ev7fdOJ7WHxt5Enn4m5yf5VpBj/W8KTV
oGrItSkbKJf2mUXZuTO+ziazPhoeDsy5/fP3CxoBexI6rIww4ns2FDBUPX8/mxFhguy9R7P2nQFN
OP+BnaMBr0PJcvBpLBZ8SVJO9xozjhGSE2FCoPvUyg2q9qW84upL3YDzC9qf9EgccNxS1RPygrhs
a9jCgqNZyw6cK4l9XURb+h+tWx9IfIGHdq4lSp5apgJqk8xFNpvz8ltDZMwXt6Tc6yyd2z95A0kj
d8/iMnn2I3fNfwDvQ8LUTkg1OPAQSAc0FWeZe8DZouRNek3sG+An0s1X4hSHS6SKuKqqEPwL7fla
QUCbjNJHpq1g44cmWaTGcQ0RRTucEAU9rib/ZxBGYvoOCm1++ZWM+7MbX4emus5qDVKQwyuUDWJs
enWEO1MStlHZ+kHTT0orISKkBbekv/hHxM0JiK1icT8xus/FygUNo8gZB1gDlMOmiTZobvaAlqMD
i0hiiDc3p6+4dPpNEWU+u1ewKquqEjxi8ydf1vii98DEv0GYkjThm+FBbpj3zEe6VKXWIKrnDw9K
syZFdFuem7alZjKvazjAsxmo8Cpqf6GWYFUXBBWYn813qIvCJz7vE/EldTl0MH54AkGDldzHhAlF
53UUJIRWnHKCcHNQ1/L7w+C2/fq2W5cIDviSqQiyk3abjaCQ6cw3ex98kdSjLtiTyitRxblT5Z4L
iyiD/RHXRlU6rhXP2K9bndI/fq9XOHQAf9hVZWnxYJveYQBF4lnD8DgDUny6UeOosRi0GPaAM0GM
o+27Qv/ro0s/luqSH+P33eYippsMBnLiKaoFPlA3UEKuP8evROnggv00TW95oCQplLnHzbuw53HL
Mm5FF3OxJix7l6AwhJr7XEUf9a750ueaWAaD9/7d7mVKCS4bbCyCsTP0NjvjvZw71kM/tb0yNzWQ
xu9ZAh2RfPhySRdg4+/+OzFGx1jSk2xaJqvFedRUglhzmc396+q8nTPqpCrx84tcJ3HJ9IWKznbK
1pBQRHSXiYk8irFNuNxoGvome/tCG4AIq5icPUpSSPr9r7a/qyWrp8Sil6qhVFIhrWPyI29ZrbId
+duQpoJgVeeVnrnjIR7vutMIL/GL7oKmCPS0ANvMI7PjVtxySc8rTwbyU+0a4WE/3aq9OHb+Wa9j
g/I326ZIvq/RYJ6PPqZgfL1KeB2WTI/lM3ynQN14qHWU34+Vn6NP9HzHC6BTFoYGvKMf3YpBZ9mB
1fyP35eHQaRJ3NHYvVORAsdJO76b8Ka68PNz2ymwrowb1A2qDbXLA8SWxFX649m/gVwk9KnfJYgj
6Cp+3fEtpc68HMIaCsPcdFJTDs/xJckrgeSg4OZYp0nRXQkWFzxjbGcspu60YRmdaiOU8pH+5O9U
W6aPeR3C78/GiwfC8xiWk/4mukjkwOmPKYi4oXO+k86Smelw3PnEO8WJxdcMqR6WwxqNI01CORw+
igb/ZNMF/e+GPmBaWl1KKjk3x5aKlqcFMDlroma0sGRA1NJD9TxPvj24OCsSU1N6fYHmL0xBJoa3
bV+oNJvCQKz7tcvgUwet5cjiH6CESfKvpIlrZ3BvT/19B3Uwq8iEtWKluB2+XulMw5+D92BKjpOy
04puvDd/+Z/XdPXzH7lsvnJE/w+dfPe9EgbMVZxTklgLWkJMJFAcdP1rjbrhXWt2Xbhok6J/rmAG
3Y+D28FyCfYwOQeSji6kHSYRVuDbmdFSX8b3DDAoihfcMw1pV5QYdRD07CVSUDNjND4VQ5UAyzzS
vmv1Leg6rW1+aioh2AqT6z+Mn5PKtmJMlps0BhiwbZeXBtpom4rl+K+lln/OYP2I9rjOJPF6vxl+
4l2yfh+sjMeypvMP12wOVNiytat5bTZXEgCivu/gnayUauwNZGE6p6bGXiZgS1MKItGPoIl/xf8o
y1iCmWdpharephIAYZxhMyy/9R8W86YI2FmyZQULSOvJKaTB032Yot8ftYjGNk+BoUsM/nMMFSN+
ueIvGxVRasjY0eaZm1OYAW1C3pNXqd/64d7JMXrV2ebsEp6P1PqKE0oI5wmuS2VkkTKXTl3VuoMz
nvuUQH8EaldC39lajukCNbn2iN1zI81qMT36qKmOqrNticX+XtUaXfEme+Xyu3cwBZ9aKzWdlZIm
+7soWmACTbn267gEVXgsLFatsbIOfpzWQAgfDq0eDxcf+B7G+ekHunfbpZwKlnIQhob2fBx7H0y0
CY/4cZUJoHpUZDtc8EAgJTUcND/cG/UKYY/a6gGXx4dJNdfFcuO5JZopmOmmuTfoBWZ1olOtVtv6
CmehaFXG/hjTxjRYvdcxQohsOJuwxaWKtvGDsu6KW5u6c54PY8h47wv7+tbyjmrFKFihPi+29rMw
4i4hQ4A31LrJtzqqqfAhdHmXSzIJ8GmLx+8ogNi3aQljZpELYdgLGYvneH4G2oI5dwr6Ud8O4Du9
jFJWAnXNy0f0OJWUQ20OBBGMTQkMD+2ZI46Yue/XGCk6Jv4OnIj+CXdF7Ka5SORlhL8JiYjOb6uU
yg/oWmhNKLggtqPGg2XHye58BQL+JJlB1E6ItwARSWTsolf52N9JGsIA8/hjK05+jLh0Cbxx3wiU
oeY57X6CRfp3rAWrxArEmLKP5aidgTvWpVs73mEXR120rqVXMXr1RhfRtYndWgT1aSqyjjI8hFBY
g5dj/W6JBSHic6WfGLqyxwTgR0vOtf6bqKpqGp3t3mQSY4zG4NLAfS70NT7QG1HVNxFpg8aUgl/x
EDNO033IjRLEsAc7Tbo9dN+9m9X7IMhEk2uj6CXu3l1/i9wcAz8w4By3JuBFeVPBPoC5mf+PAUae
SG6R5zNFIU+xm71HnMscGjQ52ATRyv5OSJ8BH/OqpzSSNjmQlywh02lpAfxTzZ0U+/jmgU6BI/tR
mMxVl494YdlesE5uDrbcGr/pUSYVt9kDDxzEuxCLzUORsfvtcMWQWgaGWpXXoKwdL5cK5D0olQZ6
UKlU0mWZPctBJIIXEXeM+2Oo8EJP25gmnSg9yVyGsTGIty7rLsXuEby2sVM5pQA+h4RmcXQQ1Gye
5Tvb/+WdG1Xm3sBqicaiBPh92ujyBbJ6sbEAckoJR/lqakR3rR2eWEwuIFlXTeiuKZ4HSe1t3xg9
VPKPwX07hSZHYBXe892rrSviTRjdvBkqVoHKatsTSpuPsvH5QPpBRcXG9prVGKh5toQKHctxaeUo
0p/hDPM1wHHxOrYFmTSXdUXXcl6VddBxm5TWLzlhxU7bQ8UETYjl583qijm6WehLGGWs4yAcLQca
a2RBpyvBfXl+ugwwVobqTAhiz+jCOnt7WFPFOODUXmcUX7HSRHNU0BfAbGWYU6e6B7mhuDf6b5LX
mRwlqTew9SFBR+8M1mUq0KrhzsEw57yvHij2MkBIE5UjrL/JHnsbJiYRNXFkNXByxr+EUsba21Mw
FVNfPkeG53v3jFgZLRId3BDkjbITWZi7zdwsySSfGR+BchDObFiZjXZQrlVZesI6IQC1EVcgCWB1
vH/5bFAiJrcVr3nU7PRJgTzlj0jh/JqU7QDu5/HVGjKStAijCGD4yCKRpMx70jHUNnPAXyG+Lc26
xtLZJr1zVhINmjub7EOzUYWVwmAxpStbDyAA+9SC6Ws6mCFvkfxnHA6R2RSWoMUGFhfrLXdCKhbC
3AFwCmCFd3nxpXl7DhKfCFgL+2zLP5QpWWOS3r3x14IzoKWa/EYAyOk0K1wMTXLCRGqo7m75XPyv
14Y80tYmno/mW9TIO3w3KgU+HpDUdVRMs24PXpjwdGywn+EY0B0BP0SBwd+0mlzEF9riKhRDy0oa
zYnTHCguoDRz0SsNfgPrxp308He/tK4AFRfmsRr5ucWBeVDaLZPXy7KgpnZ7wqmIlepaEjhH3lMS
sB9mPTrQ+5UaFptkcYswniAzB6FltfSrMv+DDoa1B2acrY3STafQCVmFOk/SYiOKliSck+Gt9O9t
kljgg2cD6L5enIGK6kHDT1p8TMeUcRNYoDDS7IK3IgUdDSqi4vNXwta6n0qnw1yhMG1zzUi8/MJW
I0n6PjGQCnsJsfXKu64iRPSa8sByO0ODUoTEfe4Si7TR65rwVKwBk3IV0NVdHWj4H5+lns+DLuWs
V6KQnRuMg4noXhHvQJ5UNwuD9VioaVxDzc3EBMyGUsWci1enIiwOfXCBINB0Wvbl9RBsP+qNHqkC
KuKH6MdsDidb56GbV14Ttod4wjsOquD0ooUUqlct3N7XrKlVXLW2rlXrlWFkjs5nJJZF8W6hgbwo
WdDToqiznn1SKQy2KPN0jgW2CZXbWjsaWcQnJh1WPSShbGPy8/ei4Sme5RsnFn2nn6+H6KOmFkaf
YhPGjT0nz3+A0yuXsRSXWAFrqPZp2xJ5IbxqAkHWEd/4+OwSVhSZ9A4aODwjERfL/j26bVQHDeJ4
sQm6Y7uXWH5FslZJOE4wkl0xPRHYlzuHqWJTdxzLL/rY+aG1X/UCQ1AuIkPrCp7XA5g3DeGiE85C
A1vStlTYWQSde+f9P0+8e5sD4NkpklquCjvoEBanjaIP3jz1YXNYUDLMhB7m+7ZR0sp9e0U2+TqV
EkiueQdyvOLNI6OW2uG2P98YcYL1dcyO8nFSXkEdTjibvi8XlQrQVTPo+2qVpPwmyyqbvTWyDYF7
A+GnHpRDVQqbOM/eb4dGfUeVwY3YwCVEYggZA6tzoQ3ZPjttZ4stT7uFPcftOUCE7sppdIBAopXz
mep6/Fpm+6IF8dyXiLzD1BF1lXl53juJUECIIItQqfiO6G4FQbs2mYLBiUEpa1CFCAhBPsk7MNg7
fddXCFGuNbL8kYGSpIB0wvi8ZkHhItxBWC/JhUkL7unqPm8t6iWJnWGrao/hENf1JPalnRkf2SLi
725WdmkwSb87kohyOx0q9vj+iSxNh+QUwfdCK9vODPq0Fw2fhZ2Ibz0/GQZfPRw0pUEk1hejhIQz
YL/U03uR/UU1CykEhf5neK2Php+w8OitvQ8JEbpBBbWUolg/ydjMM7YElrSVjEHFoOcJMfBB8XaD
ypavP5FSBnUVvGBoxG8EhX3PaO13nW0JhUoJVOPYx472pCEla+Mid+CQFln2cycV+IpQAOaq0iD3
+8xe+LnqqswWfcXlmDSGlmgN0irBWUCLXhIa+Iwd3JYkwLTc8R+r2DJhmqMD3LFjFUSVcTAIqFss
1KuSrobtDDTbSwdQ3mOQkIQha1Rhim5mXSv8OGmqRiIRhWQqTtNo/kgZ/4DnFtw7g90cEPPb42K/
miQTXQuOTjwK+ouaU/2WbVzvppiWmxSxLk9ynJ2mBoUYglqpkXjXWa2fWoEwF7CB9eqiA1nJtwYh
qWqJnqtXEx5kWktX5oReJwiiPHlNR/yUcKbJZpzrmBu90XB6LUqOr0Hbwn7S6uTYexLCEombkVNT
3pm2te+vDBfLRlVRSD+YoKB85O2mRVeTEVx2id9gKAwCuhZaNlzdQc4zDr148z5OWL2a/AJrKcBt
uYX7Q8RJRaRiED5xG2p6Td+XN4EnLB2QMEl4xYMnugWBPYp48vVYSyFuIOqPBwJRk3W6+syYl+Z3
ZTIyG+uUvr8nxYZe6oj2K0s/pfOJjkM3Q3Ws0sXMbaSuW8oyO3zlOeee5roKvdsbGhFFMhfo5TDU
jd976BAABOZmZsXOQaEmG9iXzA2FsXHFYriLT7h1d9EQohsvjdyRR7oRtCsIZfFKGCk6InlS0ZD2
/cu7I09sbwlFZz/eEpX6dyZHZl46Hf7dIVcV+cHsi2JnINJnbdY0SjIqMEMM/3PueJdZzilql3pU
oqErrwlElaWEfW6O9uMyMRyX0ssO1f2M/Q/mDCdl5Ifft0PfIcogTei7WlWfjMTVutot+sCgNg+/
SNs436+MKr1xzvBMUV1X/7bfVgplAQTBXNDuMnXOB8it3wEbnGrsWlXLB3m/fdcWBu5DEE8fUizI
Q5hSKqIjhWw2T5Kt+9MP7Tes8hg8SWyLsW1t5kbfQvNZ2WcEENpFcEVv7H4t71mxGdIv2GbJvUot
hitz8PM+wUFWo5740DTRGX+9lfXA2x/SchvklUGKyJHFa+Z4AcRAtxykDbupHEFqvkkN9NrE4qj5
TVFdVY5rX9p9Hothhb4m7n15ZceBugDYhVv3R0J47y9mCN6Ny76cMHXHAQxS9PQb27vx/9SlEykJ
1QCvPA/x47LrfUcc7ybLGDYGjmauaIBurs0PvOVVLa2xsEaViToSO1DmcKmtznliqd7axwtJCvTU
00RAmM8uwKyFr9ns5Riti7iJeJVaYgn/OcFGIh2ysGlVOcFmJkWyX+NgJGRCXH7yvv75Qi22HKgQ
BGROa/8zooL2XeAiHgSt1TBVv7ur11EQ1PNZt/RMHKyC9jage3ThotbbbYNtO4baVXEbFd44QZzD
Prbi0S6S0dBqY+ygxOootsdaJojhlWGGmnJseDkGz9Fxc5lxjt/ibYrgw59PM9v9KcTHuwzOJpQZ
YKshhqyXbc8b5w3u6ZQGmmOjlPotkaeESYANaihrURKJH0gWe0yIIUdv2Hw4+r7Ts8zJZoT7+AAr
6c/qApXwIk4swoKpwoUtXFQghRESrhcso9Ouyf0hTyn/Rob29M1xfHxsaxgiHKgCh1wVgkmqI2/1
s3p0wnVuPjj1+0tUyMyB/MrXeiUDWckFN0o1xZ7Fcvw7Q2KXd/CG54Z1fQB0dIDbBHv3MktZ+uXE
Yu2ngN6F3gWeV12DFJLGdM1oKkMOYE/epg6YrqKmEvxChIhHrfgBabDgvvtmwKoeqXnd9Sl8Hjh7
E7WpYFYyPmwrhrFxzH1RAuJk+ZL+4VwjsK4E/CePPuOYTbrEuWDhmY1+14xEbNLXM83JOqznstUc
k3Esaw5cS+/5yxBcO+JieZwdTXWIFXuR7hBVDoZm7u7f7YhulnHUGBoOVMvuICw8rCNS95VlQGuh
diqZSDG1tKG18iFF4pEi/UL7XuzPMymiUgRgctYTVc7nyzhY+9PmqFI1t9ijGRpFuO71pBihdgdd
yyKma4FzSoSyRb1x7ISYQQrGKnPnETywiRl5TsQ+Awxdz19aAzzQRV52f0+GQS/mwGNCAZogA2nf
BA5K74+aDmOCYqT3EkunHE5kPJr7l6M+zhvGFsTUdqpW3oNPM+ATz7mIROPq6p3/VbLfLilZocrQ
/H24kq94fE2Pe1osiB3eml7DGUfbszC91VjNuuBTxIEasxS/Oognht9DFJe6zER9JlLNIsY2uzEB
h5bOyswqSLD5Anc53GjPOfh2leSnrpBDTqQyAkeqX8JGyvgVOIbiJmM5NfLjwN4+AuZJvRf0CU3s
7O4JrceTWsEkz06VHDxbnVSawIKBxOIMR0eXGaIG9qKmLCZD3xQEp71mZXL1+8RSoBKUmCgfyQ8Q
VolXw2ikqrRm1f1p7z6qVoqCljZQ1ua0eG2pojl9AOF71UJYW88+/xMBWMdDz+3fXO19twphTLRJ
lWYfdZyBPS39Mmm43U+M10SL+CinbroaBhYsNBAeKG3gzy6cEfeyAS1SfCJbzbKBYKtSdY1zIImz
oq+IIlxLfXOHUTiiyDgwfCKuDo/OeVv/gIubadTxE010MLlMaaABWZANQkUV4bElQcS2KpgYEcC3
iuAMDzD0phqQNXeDOIuGn2jck1C0y+05Tx7IoIuvaK0aJplKW+qpyrlM2/nfPZ7qnzuYnkIZay3D
vOgky6/xk5HSjXdWxe5jBEB04RUBnwzBN3DjWVC0W0Iq74qIXivvPEK1AZ/FSEr9gQrd1iaL90DV
sbnMn7ldpEVG+GYNmQgzc7uwVCeWGnDdDbPfwgZVdes73UuXXxya/uwt0n88bDHRFzeKqKtou9dr
ISsnJINTKX2f5u4jn4nwgpGoenMQUCEul322RbNwzOUc2W4mSLPEOgbhl+MDSmqMLpIteQ1nKPPI
F9GrG3twr6f/JnQTR+lthHDPok23M93GZ4gtlf13Cbp5APH/zRCJi2KqmqvgTLS6+5NNIqFxVrgX
/o8ae8//sn26v2P2TYCsyMy47WrH3UmgAsT+aCIC5KKnrM+FUezHirn1wa95lezpv+/OAwY2rzaN
+yWgBAEekP5WzIs0GUKhwkqVJl2qidO2kOJQzOfgZSis4/K+JMmVAcD+XhRNRlAkm/bke8Jshgov
yNlRm5uhGoz6rT/0oUsz07yqu8N3DUGDFhWMDNHbS6KivoTFC7kwEaPMzvmKqYU2maju4p4Dtsqy
elNqpUdpofqeBy1QC06P72rdCmfUxES25JdhoxyqrCLPVlvpgIQqsyYykH+irLDJo64GvBJvAm1R
9CJjGQUW+VG0IQq0G87dpiAZuZvogXkHgp+720+ehhH8j3Q1GnH4mFzqizg73S7PrFlAxlyRCSTt
XvY97Q/lsu3921jiBpK5ILjydd4lRsj6Gu7r23tLXkxEyhy82ylFck+67UCcCR8fTTfGtEt2DTeZ
3ZFXqMjCPFci7rLts4ggkt49RDhvcanEI652/L9SX0dpHaFj2WO037b11vBHtYsvZVikl6veqi/Y
TUAHQ5oFKo5ERzVdyqLXY4CsQoFdGV9GjdA0xKUumihAla/OYmScwlzHul05wo9xMnbQUDqqUN0y
bx+pyTsifrwbHVoVr9OrtO97QLc8sljz7FBQt63vcSUrcL/BiycB6M7Po9u7fgbSCcZmBotfC+x6
Hc/HUBxDfnbq3uZJNNphRB1qhqQ4Xvj8lvgXNlcsfA0HgwJ7pJbB9nmA3DZjeAt2aVGozxybFN0P
Ns+0U8lAwBN83gRUekdVZxlcsz8E4lCpmRLAUt4gHPBmrX4uynTCyHHc8NJuLYXLzeO9N9NOzYkK
BRnO2bn4ON9diDlRg3erjLNzMFj+OZW8eNqBSB3mYZOySDcwMWNNVouxJncr76AaY2TIOvHcjxDS
AHVnhfWiDMOnLicH7ZqhyiAPqitR74g+2BB7RWY8bWjSxeOE6eVKZbiYq8w97of3PEyN6a0dj7S2
7ibCXeDMXVVaCnGCs+raPEsUT6mTrWgEHOvsw4rHwXi6ya37QH99Zhg7DaY8/wR0THkaX0EUSq50
kSV4P8J18a23v5HLukSzRbIDxoW1EbG61u1hrXuh7KGFpwBgNcUToQXstFp3hSX2ensIx/XY2eZM
abNQEeZ+8bm5PvwnaL8kLRUBUSJ9q2HxaXQLhSHNAdFIUq/KBi7Fr65E5ugYeLH2xMrJUKPReFFM
Jb/mOcRuj7yw8KNOKrKw4qNDuMkpQ/SnZmscGA47VxwTvbEDHd0SnOHFpAX63tqGjvYjk5+SQT3f
FngjFT6ZoUZyJgWuRIhUoYojXdwkMgbdOgi0aJVYS9GmFMxdBaOYzw1ON3/DGVjE6fC5D0WGINoj
29ZyX1ZYVVRF0IXweFmxsd0RQaIe7ZfhctnfUa0tyx6yz0Nd+rN5nNwgfINS1+4SBMsfvQPQNc+8
YMAMxxpnD2qV7OghhFQ+6XKXI/soE4EYXA5nZr5BvrxeizoxS2+ZTXVlj4fIqZCofI6QXExUA0HJ
iJ/C16sV5nedpIbVeaaBtFgr/QrLhhXVwIByqPNOXBA6if0GwKmHgoNOCwffQ4XXWIPgM8vlVbZs
galI7rb9j4tZDqbaSR0Z0wbyjOapMo2ebv2DFHitMjOOUgClvKbJbLXWf0/9axctXqXjTC3vtAt6
j93nfE/BQrsItZl6iPuLTRqrwlX/O5j0HHn+PMQ5UkZB+XL5Nih3ybmtBu/S1kt9PxZ3bkigO6CD
odWJGg8c3MQGaNf7glcC0X3izkqkVHWXpWw71i59hIeNM5c4QIQpojDalX74GZy64+E0+jV51yoC
3cV9OdiK/95vP5TtGQJxtT3yh+gdp/E3yeI6ved03IXNetirifjEkETRXx30phMKh5INRyRbHwXA
4Qszm/6OYED5nCGKPhwrGeSRo4egjRsJ8yqSORPZMuRcaqh2QZ+yRIlYYOzcFe7LHCEsQHCwYvkE
hhib2wavjlN0iIV+F9rxm5yk6hdcOMZmwd3dpboEBwmoc2KGi9A/10DZhBQQMCWIWJuGDjeRR3Lq
3N+mNXHeprHyWB/QITA6/l7qtFlSiRKPGhRWlg0ZdBr+400c/nUOzpEWIDVmJoYMe+M7nrjb6AxT
WrmHT5vpinLH2c9BuGgDW00CWSyi1ixDfmY70+sRqHssZaBvlRfQgr0JoVORtPSYPC3gWhQwdBZR
5T9O2cG1whadJfl/kUskcwC0kagEGo4rtnsfN31X2McyPjsyvpQW4G6tFlBwxjFsE193iY8USO8d
Go5Ru9jsvplUK4nWVYiWE7nL/QZABHSO4huXsTOqYNRjmIKzhSFcCe10mwRm2lpeHfWN0bH80spn
wxhooapU94uFApHMhRFh34kYW+9uFhnjvioA2MJ19q0mF3dqi6hoE4pTxkeKDTuzVsHpYBamujPH
0EIEKXlrECnwX1D+TJZ1SV44CinJbu49BE4z+djsgr76+wMLTWIWE1Rbx23oLUIAd3Pei9FvozNi
JBXGfkzcXFmnrMGMyHr59FuVFx1sgZOmuyyCGr6eBzp4oxLTbnh37QSVS55p5ziX880jnSYew3Vg
Pth1p3ZPfTz5Wpl9xBKJDKJhc+yeoXthwJu96sq70O3mkyvrGbrWb8tLTWSciAhgq3P8TtzJXV/i
HfhacrjIGPoTspdCQbrbeMyXSAOmqoX8qpAtu4BBOeFeQfEjvYmLzQcS/mWDox69bYkMn0/A8A8W
jt7cy8S+IZJCjv24rYSoJfUXi/IZa0Z3R77meImSkykT/VGCEbJQFG4qdH5Fj0nDt5clKvNxYA+8
O8HRYjvfJhg5FXg8kMHB7lQ3Ta2mrfWi4ovxmlq/bfUb0kEKlCZtN9c8aSqwdOofO5p1e340MT3m
GxdF26df7fLgmb7U++g3adOhR8+93ptit4l+SnqxnsxfyHcS+uuhtscOM+RUIFDF6EYRpoxNAaWp
b75/kTdQaDXCGkJt7G3tsQ7iT1awETNDQP6IEuxZjQgKr6XD5EQal5L3j/MxSx6WkoOOVYNoP3mj
E3lWeh8ikQhM8PgoHb/ypsKDWRkBdQ7ieQx4GwgS9ygL3QNbBOZ+v636MRrq+Srkr415PF2AAckS
z54jiXNPWNTWUf3YQrBzwVNUeXO8/H1khcKZrnkjR665TlL1Orh/HkDM4JLg1HEToBjeArGJj7Ph
CMuh4Ne3nDtnEg2LkDoiwIYNiLoPYkGyV/MxhbCGqTfOvLl0o/l9sIaMWw79BNw7xn9EEPgAEdJ8
5Vcw4RklKc67v2LoC7nGUPgNq3lrnqDY8GNn2Lz8SFD+uk1PvveB+RHNxmfWVGwrQUr6C2ntusm4
T8bB1QDbGhlIZf8hCUVY4Kio41KQiktn6QrpijfNBswkDPgxXr/FXk7V0iGD0P8M2u9/c5CjK8/D
mE2qGc1t7hToqFE5TXp4YKPAi0wik6y6ykkMZdPW4BxeYivJNRL6AZq/IMET1gX97TJAXPoSR4Fa
kGJe4/+zf412RDrucIoQ+GWbOXsQonIN7rp5Meq+JXQgpedLrM6HYhMmySeRByM3yDabJK74cNr2
QmHXBN1BWuyPDx62GFDso2hGvS5ffxyxGt6jymC9geuWSeQOpR1v7J3QQN0+DfPnDVe/nO1f6MAK
w+UvHRm/RDFM4IuFr0AkiU4mKl5bS+ckG2fyFBkeWdMGvfezUQaD8tfs92b9dEKvZA5Ryn1bIv61
SX8KNXWC4iUMn6sqF5adakCQll9D1la3j4jsubvsTU6C1MPQXnfM4tnN/DH++hPv9oo4UqXEBCZJ
ako1gA9MMRAUyvHHnmdl3uZtvCpdGi+SuVSSuDr4VTVbx0tV/FSavzdrUlMGY2GABnEbes56PGEM
7SxM6zQjn6dMpbTq7GnKrGsZssiEDRCt9vooF0RnJdNMnOtVA08XWr7d80e5zmRxjnSuAAGseQ/u
AhGf55e5P/dZgSkAwsZdtSuoGOFsdMFBEdHqwL2AxHb0dSvwN5qjCoYLgh3DhYMLsKJUvA0GuWPv
aa8Je7utNCgvwLIF2l9bVcDSojGVmeXyO07DZkPli0ccPsLwH6eUHx7DXHWSY7VZvQ8vlrEDXnLO
kkp5noWa2sGrQOQgphB8nPWdUTl8rtdwA/YqG/Wb+jODhdhsAU9R2+6qIbcrRoRXR0Zftv6iAMPM
BQLO/VATZ0ne6ZTVRyh7ZSpUmISst0lpZcxM2MtAeVw/8o0ko5lkLUYawyvvTVMafXp0bzbbSuz2
qbSIm8dQGQYRZhLOrH7KVX1u3ahyKUR5Abi0JZ3lNjaTeSolLHyFN3ItDSksGoDfEMnxoFCs89zY
SHUAQw27/7KO1E/Zixpi5p5ueZxZE9PKuggpul86FJ8t7ZGjRZtyybLxoYv49sIgC4NtVjCm9n+d
m72tEUDMUTTqH8Wf4/BbXXrLzqERBggS3PzVgBCfjNjIdgHU5nDpH1zXoI6iSDfgY9Y6Gc778J/w
STskkHIuvO4izqyJPZo4XQKSEkO+T0A3a/Kw2Faod2kbyEm8R0v2mSGRwOmBcA/xb2gdhh0Vk+6F
YDF53URg+LGCoKf1eLPFYdTYnKRS/TAmKulZfbc2MRXbNaMUD48MTEkIKoCyhRFVaPqyyI8A7hod
VXfvhkL0TrlXKK2dxmRnLIs7ARAJDEWj7L4otKJI965+Lsl2ysYkjGgIsjs9GYsNoHDkpncoOWoX
bTIV2btdHoh1w9o3TVKiGOaOLyxSEHNXr0A24kl4TQIBblAZQ2uaCGkfpGJg1VkOPZGKlkaq8Wyd
roJyPn/rHN06Tyc2vfPQN9q3vPtJhMPRHTnOioB27xKdH89ZGuMcUk4Dou6thYyLzdONMx6YDavY
99Ve7Nh712eKhyabsAOOETtTfr1cUFgynS2v2iKrKdFv1Du8dyxL5h+guMB1QJUrGJ2jep776SWb
TvNbt4jMogqenxRkGpuyBN1SJzZZHGYZItpmHM0922Q2OB0DgArY++Vzb2tSsxLzL428mF84I9DF
55HtyfWRVLfsZzfSyCmu9ipgYBdtIH1I4kBB2iQ+wn3yEaDcvJ1vAFXECvMvR4JdkztCjqxJFm0e
Fp7cvE/fjaGgp8sJt+kpOZySnGSnMlu1+Uin/JSw7f5oSSfJ2w6IAQ5jp31r+GL25Os7hT24BusU
hZaw4ns09a6wzLbzRfZIXyns5EmNrPtrBVCt3FX3iGJv+XvDBn6Z57lW2qlMAtwWL4XSPcYpAtwk
En+r3Mqa95HaiCluLe01Vw6foq3qw5sKlzvLgOij6mYCrXJs+Z6DBxOMEwUhMe9sMWaGOT8K3uUP
MVsgVDjGoAyYSQZXI7BuBwXJ7WUKWam8GDQWJyXxtrPMlQxs0uNicxBBmdbi5HaTy+J/GwZBjClZ
S5cg8wDwSPcqo2mi/lCpULSZAT5xFMT9KXRT14NaRNJ0Mr/flBklyYiJMPfroSZLWfSqqAQdsK5G
W94V2qLUY2Q7isztlvn++z9n1naQ1Y4O3SOy75nFpz/uq1ScxpReueq8mEqXD19tbbkr2UdQx/ll
MN+i5k+vqCJELh9Ao9fZ9/1117nPr+isDVOTnVqU04L8dk619dQ5yEU2/KUR2fbTU6BasT1nWHOl
/qlPk5EXk/lNIfV+hJDlluxZtnNhnH532CAwyEg17swGlKtJKF94a+4lsh7h89CnLzpX8BV18AEk
vS0aoKn9zBg2uWsyl1lXLCAWG9HdC0C12tatD06RJt+B8codjZD3PbA76zbrNm3qAe+pHlR5lYRG
j8NyAhYMsOEM0h315ogArc2Ggsin68Nl+Cw6iLEGH2mAfYaIr9W220BJwLvU8+QeI3cS3qPEzijt
pH5RIATlJx+3tR2sOBQFaHZWLUdSW+hXB/sVPBRnqaV6RYBQeGWQH+btxwBtPzke3rgIw3OU8Jxv
2Mx7tcDcWlv/yms7qYtniFfyFPisJDf+VZdbVrmZTqdgEiRKYcyBIK951Pd2RBpfYWkUnw/Xil2d
2bi74hGWS8mMpZvKZtBzQAQaN5lm7gemYBgs5zLxqqpEcn6iJCHR5WIvzjrd80Cwkg7NTUGWn0hN
j4h+QHOYcxjfcn6+nyP0xn3TUwk8NnsZSi8CG9ywOrzpFCroXwEbBgKKgJjoSISixcBpcIURD1H+
S3KYhDz3m61uSFC3C5zxWKR/U/EcOOnWc7MrDbYA0Jqn2MslRN5BsXSyrXLLhHRoh9zIrILwK9Mk
hcYvu1+u4NH5N6bpEWoiOxwyP197vaz08VkzRQXTYDaZ3g90zuVRlpoc1T9VATVBhcpOxbZRg63S
yXTfaNYQwlfi1hjBpmY4h7VjNneZJIBWkVoUBsnMaKH88el02jnBfCHHt1G/6Ltsw0yeyksQ5YLG
hnML9+D8gnsfF94pc+It3O2Ka1+limdHwUK8JBZmAA202suBfOIwldSVxd5KOWGc35p25E/jQiZF
KK39tBkizqG1H/ue6xsdcL/YYlvMbvhXPEGI3rtYmWys9f58DoZl2YVV41sSYRxl2UhXfFPfqzKt
pxM3NZJSfQLD/UKWUJOJFRUOjQDBqMyu7uO/ZPfLpX9+Z37ilRQvP8lYAU5q++sJYNz6e5Hvgtuz
KQBG0Xn+iDgi7ZzOrJfmKp9ZCzzcAMzeuhjOI/VXxYIxERkv2L8nIOEcrpL8nsSPXVGjnJa2Tr1g
dNkgLdlmknsb4VGv3WdV/ZRXw7DS1PWAiFhvXmrYn0Y9MvclWXyZ4DXJog4MJeNJK/kjncmmRsMd
ieajZHkL+XvMN3fCbBG2KbyAbkI66oYk2ojTs5cwNmD4+iXCjlu4TlU5RC+pJGavMc9QNIi3UPK0
aVqC5aqMlMXr51HCg3G1JcEk1DlREpP4eeGlylGv31tCelWSUpmeAp0vKR3SMZUV9w00rYFNdlDQ
0NGIWBZgtGdyxK4KsYD+BFckDDnH8dWewW6LfnuutzWjvFu4xLrtPLKeM3K81uXl/NNjeTHZQhBk
1SZAA/RH/XA++qD4V3K3sIjbo37WXVsikBbeQLAVLS9GN/8I9DVYDg02IQE8jcbM2hzvcDIMIdWf
fVvBZ/NvIDxpdXOGj3rI2wgTF0MVJ6VYlnqqvXqaXdZcGGYibmqS4RD3F1fPQXhrhRIueC06cbys
n8Pl8ntn/f8pVcUC5ZD1F3IaNpcjXpGS49yH2lfq4mw0odR6HV9KW1+FfHl1vo3rSX/DTq5tjO7E
ibq/l1h9j6lj2qaunumd9ZNkuMkkHshAvQ7CGNw+6WgOUoGUSLM2l74YZjXmx3MwI4cX1gMDJq4v
n+C2wjADvNseHsT1usx0heVT+Sppe7hPWy5iCH9Rxdh+ALj9gEvYqn0Yn+Lse28fAqWi+IL/ucrM
j1tJkAGgwnYw9/N/gRbioCLRGBJEgBa4SDtWpMlwYmukjCvUEt+aPynn2inUWDJJdDXctMOAEQGz
F/umnipL1FeZDD6LGroOAiCEOSjj1OEMAvc5YdI7g8jil5v33zJpYXWAU5meR0nEDxG/QytHm/cf
6t/NJx/kJZhn1QjHiStjC2QGDZ4xOovYyLn0nxSB7zp+EkTRGywib/WxidTvYGjGQZHDXD+xT1HP
3OX7xQWlM5LH2XVC3lQpZqQ/kabk/w4YUgiYKTSh5lHEDC7nzXonL3tOvxaCF7/UM6nm46r21Pvp
wn3chdi93cDz9DNFt3p/hX5WjFIhbAiDJULP/UgWXzHAh791lMTuISIA4Zt57ns8wm4liIilSn4M
Et/HgGODg2wNb/GFHMG3xeZx2B5K6de90bqlbNHayM6ORbNPGjnhY7AzPi7mM2TlxGtoxxpYpSDK
h2qOdb1mAYILPR+GgxV3r0AqaqsUbnUsQMfLN+hxbrkt57WvRbhRqnmgAGtu8knCR99tyg1SdRZr
SZ7aYWvjcVpY2fgCvMs7TH1j21tPWl/e1XZ0oIFuooOaqIVV9hZe4nJuyRxJ2iSpiMeXWNutX/G4
OH4Wz3TtxccwMCC6jcHX7mILy4Yh6uNQp2KjnOiKverUCpuSjpYEoF8NRBXuUYx6e1kZPjZ84E4V
S+15xklcL/vEzd1v+s1yBCQE3l079G466NJd1iCp/CjiNwp4l0sfeO8NJBbH0heLFC6EqC/3vE6b
sBrD10CxUYvmOVP+BufdRBX5g2wXKqpM3Es0n8wD0eKj/EixK6rZ0IczDqqc4Pa249eOKFktGXP7
zm+IRFc3rEMqX50sa9V6bCdTzzeRGrZeXb05vET05osQ9d+WiWbe8gPpXLdVWbXadmyUJpw3soL1
krF/Fv5p/+mAFILb8QPGmHtKBwN1U67wTzeQCZHWpsXpC3vKYkczjU5Oh+lBOeKrPRiXok18K5eE
1cgoJ4F7mKYhwSoN+PS9oNYdjwIlHoCyrWEts+9qCCsPKTBsICMCJ98JfGX9kXE//5dNf8+4k5gK
NWhAIoLcnm4jDkoj/e4dumi7+KJg6UW2Qysdw8OknjrGACkEowbk8lcuC+R+skCERHdwGz2O13cg
o/olzGqroEs6woz878FHXFj4sIT3TVBB8aYMoIgY/xLL+jJYKR6C9zttWaFAWWqr/f+R263b5u+g
6gl184MGgItsh5rcNIifJ6CtxKIEr3aNiV1qQ752ct8//AjBpUq8NFf/F3FyiuvYSf/ZixJPqpX6
xiXvI0qSHRy6syghEKgVmgk4OVSmtnylSDAcc1wg43sB5uFGuFYiaRSOAtdUGnYiuaksa5KIgWqt
H0R/6MZFml5SvN9qYBZmW6/LP5lJ29R5iM/nssywR5QGbk1mYDfZntVK+G92YcvLzvk5Rc6Xk6Af
C3hwBw90KeYScdDJT7NfoGt3IL6X64vt8Ypq7gk5yxZDxFooHAkH3+WhkQEDVBcGsJ/yqlEQW4/v
YwOeeuk83u9NUF8SK+E7NNqdj09QPpkMlXnxU7Uuw5Nd9In9HkoKo+jSUUZVpqQRIEnlPaZ/bGci
obd0vCZJxroDlYMghv4X0P7127ebV+dNq1O4dfEqAJfhyIcTtJjAotmLek9PQHuRvB4l3gc2rl79
HU/Pa+dd2HiOgBaQ9pospJVnJkS+u8sHClu6xH+68M4+DBE7hehO0szJx18gaZVeqxxWXhBWaT+B
nUw8fyo5NAOG8IXYX/CHQ4C0/FQL209EqxvtIr7b/WoNvpybgt/uZ69N+97plbUcqrLsHVrpos5C
GGHU371QUpRtASetmy6e7uUavhnHomoU7dnuEm8MRavkM/CFBksHCAqPI6nzhXduXniHYfR2LlrM
g47BR4ySBISK1ickFMD9gl5Bn97Jp+I3biqIgIhyqfDFjJ7lEHfCQay2vIzKxrtS4mMMQjdHs6ii
Pct/W0Zkd07HC1LFAxWV6vmmqCm4JXCo9ix1eQ5cVbilX7BCrx+ko7QLRg3AeddEIaUfhD7yK9x4
+WdUeghzQvzpaoNu5IaB+7ZYnPzDC8m7CkQ3hDMY4l7X+1Ci9iYaYxkRB0pihiwOXuzBjGoYzpO3
mDWHvkkTTZYjaWavB0VzVPFC86vbpJLxaPafQDaqQwSVmeR9lSyA835N43DjYfonJy9OTaIxWA+Y
DNojqqeNiLZHONUQcC0UEeJLIgRYeYhy2WtebwTZTFQ5UeAaoXNYjGirRFVfPxkIfWVxCGnaUild
jB68XNbim9mGx2/HoF0QUDdhAhSlWeLnlEEE0ev5gc96CKNN7VrAH/E+ziNEs17fhjYNQbPcSqoD
vc7dwyYGrhUk3NgzbArBEeXOmpSIeKPZywY+R+3jn7Y20hwz2Av/CqssQ+7nJLehWL10PfsGF9Im
7QToTrOG8whmsYLSxC2WPFRKuyr745kxAeIvT3O2yCFXAp0Nu8Zizi6TdoPnFeFV7J79z4pR/ZFZ
LRtXkPXMVhRFOCcr5ZqHpEaDP4vBzbXQ+GQa2HmVOulcrsp4wrXqPvGulAN7sxEjtAv8pPrsitEh
6A9zEJZkMpnUjVFbx3g1S9DhEOshGVdnHV3d7HbdAReFfYZrDloHn8MOhcQaUfwMCu9+EZIUOLzT
iJAj7NFyIwN/7Ab007VRJPoQ9lfK0iTsvGArAB/tuvk0aAFKTA9x96e23N9dLRI1EIH9xA0bttXc
KAFOdQC5lH+3PvWa38Cn50HQEhd7UQjLU6oRzp9HLTP6/jtYd+hw/9i6gy+n9FLfysOdzHf/nC7t
SFo/mXwqptGFhfuK2DqoQRsjmanKZ2laDKWJ6hfwIMdJDl7NqtRtLm5dq+3PYIWKZ12+OOD8wAN4
seSlY1FUD0sO1nEzNJtGI2ppCQ4nzCEdS17sTsN3cHheFuEVaa8ZxVvp27NZVk8wd7duwp7VYtee
11NwG2mvHDxz1FlUHnkXosM2dDty+zsoB6SeRNabOvyU9uvQiwlasI6wr8yeWWAGn+Zp6dEbjLbc
SUEtWp1VdMv5jiWWAqRUfzDV2drJPJ7lYXUFLAULLwOOYlrn64CUoelQiSjMT0ly/SQVOl4ZEziM
ZOusbMc31ka32fLki5zHw5RFoTQVbEfQHgG2fo7LismUyH3YYNiCjgq6f2XL9pSfxRaHA4wHmFHw
bDybKM3YoTaveKZlK7dDFyZUjRhltF2GXRsST04IGv8ncI6OwQqAgxAVcyXplS7uZzQRMUc9hSKp
iHoAc8FietK8CgO0IYDTwIzzAweTqX2FS/i0+tbhbSpGDazNJ03qnghIFP4VbZLrOOumrWKkyAdN
r9sqKbbdPdPZmn2g/TxnYVm7sI0apeZ1ZN2S2KR4NshrcCLMbASmmqNlJUf7MGNWeJlS8Q/2a37l
+0NFzbnqvcFSPXCElA+gvGTWKB4BAOF1nUQKaEUgYwLfhZJpi361c7Q1D0KzUJ3/wxuDrxIk/Lmi
VVeVMLxnAgKB7egJmXLpyIuKPoGK13AzVrjDniL6vKluG/TOSf5bYnRJW6spByUa1MmVrq7iWL1q
dExCkLSs7wQdf9SjFnj+C9rRvrl6I9ynvsphK/g+ieXwFgVY/qoqd2UXA7nDs/2IrvxIc4fQ3eNu
58f+oERB+zIWF1OTBKNXUiz1grgpaGn7jYty9jP8x1UApDtCDx1uD2xWN2c9PBepTfrGm30U5mLC
4KFZnzrEqIlF/PbMKfFgYT3nsBeWcXJ/VUaG3MfkNChcjqYbluE90AEjCBVqdUGSf753UWmmdKPj
a54zUQH25KtwnZ+omlMrirQXDNw1gxCYOqga+I4x2lfMzNgCLp3PzHRaP9GkhAwZ3WDKzGW1XZEF
YfNoHsEM6yLSWEM1Gu0KBBvx0wnIGfKaXQj4vD4naLROuspMCk1sGES9AZoTjh/Z5Sq9Np/9fTJw
QED1cF9I5uewn2I2MWKaPbcKMb5pSqDQkGNix5csqSSXR/e1n3738mIItnjMQqfZX5SRGHib2UIh
tv+Ws/F7caNQ/6OI3SOIA+Y8LtfOESZIdHobU0yzS9Xzma/xhrz5lja/shQqb8/1ZHOHuRKrAAfC
wmji3VgUyqEjfcaeI56r78xU5GbqwJMYHfW7XCj54GZhkUKsA3MSNbmP2fEToy3u9g1W76YyYIqF
rE1s7znO2wrHV0PEvB0vr3yxA9lqLcySSg9NWiwRkUW31LNv3BtVD653U/u0vXnB38yf8sNmlXbB
mECVOE98W6m0HVKdkXBxGA9XZDIakc44JRetgoJh8bmPDj6ZYuHx+a6QLLd7RKPxuX2iit5UDvWm
QETOzlo6wE214TXA0iGVtl9kv53s0n2KGPV6z4X5CHyiNSpjzN1EHWHUaROaw6QwviMBjMPL51TX
iqfs6FflmoLIo98a/4UotVwKR/6RbG2t7Z9EWDXF35DAxSj1p7qy4sxIdIELweWSkuW35aVOIq4w
8l+d2GwtOS5J9M8UIW+97b9F3u1y57NYy1ruEPI9CrrMCRZWYWbkikeGG8Y7oEBSwwBMJI5CRTSY
uCpzZfUZsAljAxearO/AqCovOhSBW/JAnAws1NxFK97SWGmLC4DSIyWJfffb06x7IWvORZytXIdz
vhMBa/oNSPp7Qy5Q+mBEuuOtqcMbe/SjgtxbVvtLCznQVTitAhpbICN0MT9mThrMEveJCxnq/aKo
ykFC3QEdziZ9pRZG5Sa/Y5JpLzYp/n/dfB4+3WMP5crv2Rd/kCmMfrOZmSlYbDu6kwM19Ygxfuvg
zxp5YrY29HPHWjE1Scl4+QYl7JEIdhDvWEr3JVWSgBhnfnuiGc7nZWh5xzhiEwu/lmVJuIbZ1haF
KTmmxTWZCMXdGDeshcO+c6TgXrJKZygmxhxNwsJRFXRrI35e2gZk+yZUonqqTUvChD1DY67ttjnn
yRwsCowaL6is8JXZ/qwqVcsZdyMl+P+1jK9l1hIFbCSuhNwI/I3o+eBF+QUdvMKPGBSF92H7Emjp
Xgk1cvOUoVLMca/D0ifaEWm74/dZjJIpsJKO1vwtk75yf9sn3ORSuFUvcdM30lgXvYO0c9nmlfnj
ESzXJvW2ASpNkogPkfPYv9LbaUWOo9trOR3CsB271kI8JQEH9c7gLbSnUZh9Q60ZHz5ZBMa5uVOa
KpvwZxpeAopb7LxqUJr7sgfaAi3oFymNIVJLaV4aqsQOOTTPhjXh6pbq/AGK9r5HPFAqzAlKD00O
wNNe6P27EP1lEcAkj7eclQzmOmZdiqhMAYiKA5Zp/SnWWq8PtCmz5Fm71OJ5Ax2T21JLdohpkz1O
VXa+K6A+scf7CE9fZXouE+nBz4YIq5AiQDrEJxhG0XOdDJCHRJIZsDz1kH2RCQ4Nrcg5ckAZPPQS
jcCaybZgwbhf5iiqVP7DiFiS/yCUCkKB3qqM+kLGd0RCPKXiA9H389NYK5s1OQ2d6qmaqRYO5HZ3
wyHij2brZ6jYTqYy8xe1NBUll2/qs0ypsQRWWGIGjKxP/SOWAF2rlxmkC7Wj+rfUeJQsUCBlSKzy
x86ddwJjItqD3OrJ7riMovo/UXr1xesShnPnANSqdcSlzNXeIeB+dPQz8MhMFyo4axPX7yzxN6Cf
lnNWZD/hjG1BUM1OyKRa7OCyKiKL8syNO3C8HxfglHtRHZiUjClwa4K2peYTrTATzMaMd7yHvBAM
VP1hzx3fnh5X/jmHcm0//9Uj0qkxVxATzpgLIdg6feKE1fMhfv4ZTBQb/b05eyhvrM4agRpexQ5W
H321DHB/0ZAfPDpLtvOke7xZT9XEihxec0543ivaQQf2xgNCj1aLm6IJ/nAdl15kOxPUr0yMlPUj
LgYaNFAKBZ0Uv7NLr1pgZRfa1W68eM6X2iZOjq3Wturs+8wkNkWuG7btfiz+mB9lQ/q9NtyVjzTp
T5fKXRK8zxWdBH77rv5bA0l32QkbwqQsy+x/LazdUi6yjcz5s9ZvnB4u7kraLPQAK7lIGmSypaf+
XhUOdVqhbpa77oo63IubQX75X+431UykIgfy3a33J3A4qCP74vtSs328DSs9ljXZNWMy6GDgSrlf
iLWpE/dSmQfbztYLibSMS4r58Qr/DK+hHZryf/BoQGYBJeJvgwBTFl5ESshfgGp5t279A/C/88F2
Q9qyYGob4itBrz6BOQUVULvjjkvTuYx3IinkMAvS/tXLYzCurZ4f15M2JbLKv9iOfR7FZk8pu8es
wYyWxMQk2/tyWmfqfC6SSXjKjHLPPAilMcyxEod9gE/trYOPtihJ4Bn3X/gsQn4/OhD3JFJLT1T+
n+m+qyI9noseT+0swHmM+LdVO+KUvorRj/LIZWKHCKkfuolqyxf9xxJ32we4nmpgtgQ5klebLVj8
1zuJ4bEh3zGXhIsvzjUFAtXaPIUh5/Pgm4rX619QOhRJMgLyTCnQEbx4F52SbFmZ23hXhHtzFkRl
9cq6ISYC+qahZG2msMbrD2W8kwDWLcboOcc63smYxYYpWxtzp6EQy6EFLd4EPQzaVTiKhxve5zL0
nl7B3X2cMCLJD+1tnZ2l7YpyybKDiymXHHW3SbdAAo/H5ivFbdHSyF0ew3EVfBhrbrsFbP4ZZvMz
l20TcZ13Md2j7SsyuZ/u9m9jNiE/1tyrihjq6dZIsgUEpzn5s7NXxOVNvCGUY7j6nybDRlgVzfMx
/kyirdaCd0sVToWVYDK7WMxUbb8ySRoe8y6HvB2he0YlT/hm7f7a0+GuqCkrUb51OTzWrNweS8U2
DCQagieegwTuwYG28Q/Z0hGFj626FHfATsB+aj4I1eYf0OioK2ovoSB/oLH72nPcZyuGPNecDjbW
jEJkUCepwDbqprHJBGf5MIMWjTgpW5eAvoaeQ6Ef6vS4hdJPBxGQL2icXaT6Z7aR7vdu+BL72CfL
U9b0CrwkvYwC1EkSDBCz1+YOborhfiGoEgtvswffIZnprhW/bgChI7JnGQdfR8XJEbwPocGmR1QS
CvKqtBxS3qUD7p7lreoCcJkdP21LfW6MkW4+zEvY0g1xoJG02/fKWHQEfl2H4bfLF1gPKvsduSRF
OpZofjSuvY2O1RKzA5lBGSpuTzMeoqzlNSzQ6wY71fD4NoH6sX0uLYVGT8dE+2PuRGD0I3SdlOKp
NTemAT1NGfh04Nt7/MJdRI74oORXf7SW9tivXQjMk05/7GNgLu6+pNi/5QO1PiSAtYT1zhMnDfK0
73T9DTgRb/kfEJ34rmVU0qf9fGjrydKpSi+jr25t76Zz3zmgXq81X8if4O5AyxU7Tq44PVoJDZmV
VxNavdvZ2Fe9JuJz7xhp4LU+nr7IhhtLcI2NEbsovbMjmSZV1N6BIf+Y1qJ3Ijd4L7HNDwZxS4dr
vPU/ziWoWXufNoqEll11pM+Lv0LV9B0mWAcLWMu96IfCn93dlBQWhC7QEBbgADCa6QLhU5zqfNKn
dvTTn9xJnm72LO4bNA0lwyyYJlDTfBlIPoCqujtJagfpRWJqYtYVimzHMw1rlr5cu/qJgmCGdZ9G
1OoTNHhVrjNhtZ/OFIKBws/NtqYyPm0FKkCQJfO2Ak2hlT/pZwys+tGq7O3Tm370ace5rB7KeET4
G1OxUntx3RT0UWPe/50YpChnT7DjNYJ5n7lFB3mje+cVYGeQ9c0QuVxMOKEm1D5Kj9o/3Kji8mTD
QauvJ/7CXuMkpDqKHQO0sgSnxP9luqPo/iKHTsHh4DgdwP58IasWWyoFWay71xYCuDWavH6F7YSo
SlNOgg9ocZL3jGg/wE2EH0kPIhx6wDTaO5hzrqmLg1Fw7zENi06IYTCLGrkndcdpTotX4+H5lnUT
HNsaMBGLyfF9VZMZt3G5xqhkS5QlbJYrQ39OLKgXQ8eHRHaZZjdtXWNRPVUQZZ6P88q5fTsGHfaF
gT7CV+QF7rSXNYxTr3O/lpFo9THsoz+sH21NqMAynhk/TuYdjl1D/J4O+xk1og1C/QwuGNqqoK7p
8U3arACDVLOnTjTqWycQoclXKVLuVZIsadD7ecvZHj/PipzJocs+NFEX/oMlQbFFBy1uWdC5B+ux
MPtenxHhMRwM4oPnbut5fJvfClDvV5oEXLA6NQIwU6uVMXD0fWng4zG1GYUa36CPyZHKSIPLejg5
rHJZiyt8/xEMbD1UvWYfPjxvfODNV/hylej+XYe5I4W/mMpJk3s0HR3xtUSR1MmoWwzBR6+zyRQK
ntZrXYGe1k+k7Q9WKZ83pE2JWYESPqyIgosJQoq/ne3WkKFErQHS10jPkDkWCFhEc3HIuWOmyXrP
4K70fNYo8s0Tf/LN9N0RK6gXJ9acGsQRQrdg2qO5npQiwhlDwHFwJQNUVgRe7cj/fmB8/lz9D4aq
Xo5N/F7NpKTy5TbdVNzikykSBTtvzvx9UrCbaPgFma/dxp+xr0sPAkHapnsP/qi5H0LeB/Shr+hX
JzdnfstWm+58ry9dReBim0v3zrtzUO9PCti6/Jl9mCYDKaPy5UyyRUyWdIqhNK/vzcqMy2LPnUoH
KvqK4XzPah6wTc+06XJwviMJfw3O+nkpE6yw/DgTpUOuo9rfmXEiELhNOudn/OEJQSE4jiL4Iqn/
SyhreFiYiV7sHj138zpY+5evUsQANHmUs5V5y5tXgB7eYl0jRKKg805T4clpL1XvwodvEK01A/C/
/hQi2Kc/8+AeS2aNeVxmvYH3I+8B7ZQMOrM1zn50oSp9cgbbFcGKKindKZ+DPe3GPB5iHvmGV0UB
jVdO+Xs27jg96uvCY2fzZ4uI8f/t7Btj2xIFAT7gT2DojPz+v7byEbQFLqXCSUeAX3zP20raSf1+
JexyAo9+kpVLvpRyUI7Su4GSrQ+I/+sIdblTnQGY7atTVY/CMvZto4aIgtB7SE2vB2heguqbNHO8
UzEPd+vLrO5IRc55tGGgYSY54C7PNcBSxytlO+aZf3NgcLBwkYcqMKMqReIhdsic2Vwb5VWzd9oX
rIjw2Va/F/lzanv8p55B8VNwWdDRo+zFj4EuzqpwLjhYFLw2ISOCIL1spMksZIyIe2sBDqZbuat+
kKY0uIlA9YxHRzjhMIwOdyYWLvKuJ7TTADm44SO0m6aQ7+dKgYrxVuoj+ZyL93H01eMq+SXlJGrt
k7+WyY4wnmJo97gDJD1LtAEoG8fCROsIJfB9HlzUxyGRtIJ8CQXRv+poxTwHaEoOocwzsujDLkLq
uVRmz8Mo4qMBXoku0SK4DoL8rj9ecxr0fEwni53Gdl73ArN86iHY4j4f9LyFbuuoCVFlJ3mHc3K7
CbkXiBkpTQYcQGMJb5nL3vBwEUpcTN/BXo5GcbiJf1zMJkN7Ag1fwevg3PftQZ2bBK+YywxgQ6dd
kIWtsyQ+9GtjNvSch3yYYopcfaD6+uR6gP4mXTAPA7+JBNi7+bb+YWE3EnO+YpWApkHv8n+21nc6
bhV/GC2wZBDYXW8ZLYmfyVdhp/xqV8oT4/exBumv1pczV/KcWLQqpWlsqt3epjaLj5njGqEyhre0
jc0gCCs3fQgDxqhSOvJ9Xc6LxwNNSGnVMOUfkRbt5YSIVkWpccigEvIHD911DHslFq2AkGdcm/mM
h8KBZihuOlT6+a+Tav/Zfm241oWd9v4SusiE3FaxIguA9hVAPQUoH2Ck6dC4dymt+pQRosAJgI47
C5zDTE1JV+t64vN7Zd227SYbBXnBPcBGqsUIOQ3tLLpvMbqRp9UA3S50U+riTeH3eiDBA23kP/Je
+9WZfD9QRdQNLCsgO1jMVj7uAOF8eI97ehUz3TemSK2Z7DeZOuMe1rqhH8k4gbSnjIFtl3POAY6g
TVsok+z2H6aTjV/1hhgIQwei+h/kpedcO8HtwJE3dgeCAApawDIqSenaKuYwexOIfiYncKJ/ibr5
GuhoqL0SObypHpjSYnfzVr6I5WKesdSh5qJ78wM+wPoESqXRuy9CPD7rQvFo8S2lOmvSkkop88M6
e5VPwG2iF+yRMQfPOw3aAI76eovZXfMpyEI4eFM15ijXJ1DW1tUTBHZ7xdIe6jqhQxy6hc34/TBQ
qno/LE9yVCQGYB3fgf1bVtkBybgfBXa6jWDKZ/yo3h8mLS5caAqoGg3XSJWVGTNE1RuxJZQbcRLn
bvwutDJO524+U77zlrWQkJuu6O/kDjOaQN4uqvqiCmbLMYFWc+9YeD8DIfgQU4lfqlEV8WQVUCd+
mtJ6+tVgbtloZQ6L+ljmHDV0KXdDZkB4VpSImSs1EtlKmjLU+bNr9gueIyI937Y3PNxP5mt0E4gw
sPkmIN4+6MmzGeMS7dadhB1x4U5M1/ln1I0oD+IydNd0bbvXpN78Qmtcs1UldvXONnyn2uPqzq3z
f9E1x6vrNhKtVDQo8rzs/Oqr7w6TK0pNmXJQ57k6vUiwqD5KT4bj95yKCRuKWg/ssHdPZlIWvqeQ
x24z7dYcLvDsfbH+n3TzQyaY47rljazmHFLxa7MWYroAFBZFQHhV8WUSrO2/8EDpNbvAI2+auQkx
BUWm9GdRCveI6CUxF8fcFcZPXT9LnxjuQ9hzHNDphrmxss/lNJe20mwu+MUFnqK9uxMQKi/RNKjI
m0JEPMMUk0we5pga9pEkfDvncjoAVVMOReYfmA8L7y4NyifO2PKfH6MspZHZHt5NzLZ53OtLxFPU
XpnARnSG8IYdmcpr29EcGAZFC7JgCGH0WXYRA4Njzk0FhcxpzpRzd4X3y5P89m1FsE8ZTvhXjpNp
X7egkF6ZaLYu8cXNzGg7bn5dxNDUaTrNEghetk+6ehIFn0m8DYKXRFTeBSUzbzhfD9b6gmuyLoE5
XuqffyW3qOo2fTnwGQ0pz1kPQJhnZ7jCLYOYz831BQ0mQYMAE7jCPG8hZD5uWnAbn1mjm6qAah1p
bRjevjeFhs1rw3yBVQ/7ZjICLGH8kzUUtaBAJYYZm6eDPcpIbSpZtmyjcyO3yRvZos0ExXaMEG5i
pEpvcCQr2kV9eVkXN9g5jAxXgclV0fFkcVtA0f74rzwavwYQL56mWPnif9P04ARtt4nGy5HniwKE
bRdN7HFoBTXtVzpiVi4COfihVX/1Tu84k4yUjJwuHmN48qgXK28H3mpVu4QrSi69RnyPlQTPKfq3
xYcgqtNl3znA1ENvXP6CmXecjePmgtS4ufOVFcSD4GwHHLz59fAma1tl5DdscK6PWQLcrDe/feku
Y3GT+svZe79u52c748FQwC/OYd1N/KiX6KUXIdpxc2Y94NukWCP2wJJnRs5IrqdHh/lrnJj+E9NZ
8TfRgcAKfozBONkLt0BWwQSKYawi4qVk0yUxleGj5lwxpE/Q1Tr10ZJSJxn63vl1PundchWJfR1H
AL1IHLoDicArUT9vyxuSNDV/WH//kV7PKv2v9hgTYovgvfpS4exsoQB4pR9gQ1Tyve46NR0AKMtA
7KnfYbqzzaOZ0raH7oBvRujcD7m7D1tj+ljBZuC6lz9uh2VIDHdrZ5OJOhUvKJWTDWoHZrTMmSAw
IKmy/Haq7zQKj7ia1dqpxLeafuATriqH9kLcuyv6bqb3oD7izzJwpR+G/Fls0XWjDLM6bjSFQFAN
N+mPvEbaBktYau0vm00UmpZrkbEquJb+V33Bl9D+GH8qbSp9h2SyTMxKR4cbJgOJ4L5sRFFxjm6Q
mnIB54OSSGzce7eJnlqtsVsAalFEdXijsV3i0tUUhOyPHrO7Q7sssJBm0e+jHW3L85OAt88wPJOd
uT1pGSLt5Y1dRsSZSiaKtQDmKDZUN8xPBQcKHfN2cf4fZQEnc2GPSKdVuKslb4cMe1d0jYtNrMfl
10a74gO+UB2JPtvI7/fqKpFUWKx75feDSR0fTV9TzSt4/du4lUhB4Ha3Bpmj02rIMK3WlLibqc9I
5ta0LdxGNCn8IQZXM0OcGADt05QtTZanHJuRNrbuMMIfYYnkw61p5+yMwh5ulrequQnXQmNlHffz
YtvfrBKX4pDXezflH3lfU07N6O0f4hZFDJMls2g+VYhBMuPsVm71GU/MglB6hM7muZ6jZH03Ii/s
2Dl7ds4HliPzIYA5OIG+KWk/WOvluG1TGdK1cJZiaadf27WFGCX3qIiahpDaCyBY1lfDyZ/Nqvi/
bvYWs3FRDTD+smTyiPsugfVZmWTy4IR3Qj28HzQZSNxfpahXoRKo8CUyA814N3AYy3j4vT4vFinn
jN9AUchLE23KNBpP7yuwDWdEy6OjFXzLr/VA5L5mTHynnWiYX6NblyMO0bGh6dMziZpugIVKXPIA
8UPOL762ZS+umhOuLtoYfSyVjsV6ryjgmZVqJrb4BIf0pfTZNxYOZ6dVBSc+xWddeWHexMGerdZV
ct+L0bzw+hJTHVb0rWpyDeOzkTpxbylyAItA27B2zU0acbZW9NVEpdas/VqS42g4KauQNKqJ6cew
kTuf0w30Q8WFXNZYI0gsc8sTV2be1/hDm4QNwNou+osHNyGkcG+vEPwMJ2HyOuE7lo1iZpld4Xbr
QO+j90c9m8EKBzWfpH2dKqgxmAtjN1RtfCtE0pCOIuBLdQMpxbEfnqwp3E7MPNvfkLYj51LNMcMS
GN2x4MPX6phczMe7F0M9Z5aKTBPiTMLNm6jIDVg65oJ8X1n0KM8JupUoSXYvj/78sAMv2EuT59bx
4DIj9RGNnKqDVzHsLMvvXUC12zh35LeOGa8aBAH5d3T/4F2aRqc27gopiwhuErCe70iCq9Br32Gu
/lQAZ2iFtomdpBD+X+I/vXmC2kQsyW4wBZmS2/FlMrTB7HzZKR3Mc5SOL7GiiaREjxnIrAh+496N
4Vh6bgxb72jIncXPbMson4YdbhVWBY3QhtjjKIEUuuFGBjdMkTs3zZendCIN/U1VxkW3MydcrU6W
3Wx3QR/PtjPjE5OUS2VEHQWEoaiTwXyWvDEA0E2r2p9knO+33WW2197B+Zgvd8FOZyzu9zoI3jlQ
dT7Hx93y+WtKSgRRvFUOy7cZJV5/4L+tUfU5+a0OyJ4/wq0AsGH1irfAcsog/u4u0uHKhj6RiyGK
0KsgYPr1HFs5muBjpwrdaj4gnXMsTs1X20DS4y/OeMsb0OIibMIko9vLfk8krJo04/b1PbGKoeE/
qymnD5NMl4zM4h4gVgrfUJftXegOn2GXsv1jTUnLem4wwU+8p/T/nBMymf9af8Oo0CV5+9b7UvJJ
JUTFqSLJxZRKxk6qXHWJOJUQFJE9tV+M5g/uqJcDQIPJ0baiHcF1Bo+CBEp72cozRpWiFKfQGSPk
S11XnRiLaoOO0/9RrkRW88SQIpV9dErpe70Wi6RJNn/h6wA+Rim3BCp3hDyq2jZX+toqW9c412iQ
e+CKIjSYbfiZmm1TnwGwVOly1NX1Czc91/V9o7cBE9Q+JJwzk0mtndLiVVy39mEWQylkz2ppKARa
9klWnAgW7Imf+myL4ZNomAfJsbum2FZ4efaTUIOTHOcwVYZ5BSS6yA9MB85aY8wN+x8WuD4G/lsF
p6WTLhUWeIidJCKe+aegeN0Vyr+Zj+3dSe6dW0A5TprCkmZtFqL5rN+7ldkMxKqkdJFMQNbTauiI
IOu/zuFWRfk/GrqaLAogozbNzOGiwTTyl8KDYZck+nV7WztlfhHZAKEjqZlz3vesxIffcMTw0sXi
IBGaMCH3l2UuUfsXIJ1AckFuchWcNFWEzIwWGrGPVZz0iP2Bl2HcPA+hG6oxJPj4liqPWF9hz9GO
XOzT2gcPDunGTIgH69Xguz7gzi2ZdRkzD9vULMmP3++bfqO/aWv/oecTETn5aDf41ZhI4fK/c3wa
fweSy87cdbH/1RAtAQxvmMYNnCLOsKI+6SU5EOH22M04zFroVsXW0kMuPdo8xbDZt5ly1pYaUGH6
B1gIjbBdFXkByZpV2raiZI8JfmLHd7utcoPxRO+qRUTbG3oR0Fwx6gyImbCCLVU3FUPp652WCw1U
aCrjsaw+TyuTWhD9TIsP4A0b50Ub9AIZFMw+zmX31TwVk0B/hHMnxgUDb9DaMMId3vajR+ANjJv5
oiQ4KZBkGEBN6bzApIYNCq6SYD39OSDM1kJ+lNwx7JVOvBEa+GUsACSUo3vprPc3gUDq3ELdH73C
UslykGIH20oZqqqtQr1zkH14yiWE8UbTlHlv7Eja//2zdkDeF/3GwL+H9jd3ZuBbIiDUTp8Rcqoc
CCqqtcMOKRMUZAzxOb4ycBD7+Vs7AEaRBE2eYwnYy2eBCqZRO3uEWieInNozhe6GbD//Yz83/Fjf
DTpk5g0lv9gAu4oaebuThbYwzmj7JtIujMBoJwnkcv4BeEgkkr7z6DHJKm4n2LbYyJB2RyG+nw9f
w2VLOoPaRqcabqY9jxy+mezyde+QWuSNAnLSPzsrXIsUgBqs19wIGmAJILLVhbni1rePgxf9VSka
w3QriBOIovStyJWAvQLP/WPbG37Y3w+C3FSUmFZpHKqEEcqt40TxRoo2DDB84rrLjX6/hnl8kOXH
wAqWFBP9r149dZVcGg7qoRRzF2J6ZJZsyaXzHhKrJEyagsQ9XieEGj6CqfVisuQkRwQ2UtXFxv5n
zx6gluZ9NyitWh9dKF4EF1GAlWlGH7R9kVfdBkeuS0gYCImQE0JC1snCd7EDV+H+4aNdEzcnz4vJ
zN0eegPL6ghrugGd9K9jgEwjbXPeavf8MJQDS5D6FE7XZjhJOmWZ05C45z+c5egPHT7nRjc7tWtz
5ANFSpviQjuOfHTR/ijp9R1ygi2QuwRwLDqizDL7X4cE1P0FivSJN0Pzk00RlfycMwz9fs20wFPE
avuG3Tt6k40tABG2WXTdu00xzvI8bTNbLsln24mUg/fCQa8fCKRlOk1FZQp5RmwWgwlbQ+rtd7lI
DP3b75dQ0DmvmqRDipfJXIayn+13oXP5rdAfBQEn5Xtu13oifj59xOa8N4a7crrIE4l3cxA5P90N
izM5U8inwxJb7A+8MEbOiZXLAthDZf+w4tjDx/ww5VAdrMeOoPMW+ULlaD07+6GvgXeaYhN2ruBu
DG1EtxcrYQ+hf4HXtaiIgoU7HIGrRG5v8av/5BiNScDn+0Fv9aD+fRmCYQR2V5Hs1ZXnCoFAK1Hv
46swvv8Asursc7k4oFXLYCFc8wXNzldWPOhGSeXlvDhcMsD3lOFFJ4fdCW9tftSf1QK5k8msc0Yj
/9t6a/85qJmJvWfhwUbtLIKJ26Soyr3ZL7dQukUEmby5wMiJSx5AgOgTG/v9wNGvvsAGzg8mj+oi
try5QT5XZbr25owDJisBGpCcxkwMs60vEJ90L5onpWLg+sy/aZkP3p0yHBT3pJcgHHdh/eiYgcfQ
kHDCrYgr/HylPdrR4LZIM2ureyJ2xiOUED1p+jQwz02jzj29dQfA2GXo4UB3XqqDkwclHvFaJY2A
GsgAzbLN4hXjnwRFKZPLjcDrTT3KHhnUSmZD+BXXm+jargaqOsuLOv4dCNsLolRmLOhylWvWJxvE
59ChR84ydG8AGAqxfLDgCZVP8hy/iFvh10heqecCuldC1vXVLxBnPrgoxHBPv0czA7R8z3GX0vB0
iRDffAlD/b5qtkq2vVuBukif/AmMgk/u49VqmufBaEAXXuuemQPMaNtCiJ33l1AJC51KXiGqaZo0
9F3Ui7TzHBmUpZZBpYe14j+Kv32rKI2CfqE060DufqmPV+CUhTGjmD7oudUA8DpvFvc8pu5YWOdJ
/LP9Yhwcc53pyKnMdXU0e9ckcGUvlJG/8XspyDSDf5Uc/prcwrx1X/BcR7JD1ieiVEA0/h+I8v8F
d+zVuWJePD+YO961YlQciRqKaoxKwkyw4L35AI0vjRUR89GiQ04CFHygz6wmVmosU3CM+eK6KTsQ
vt6Igp9xEwXCqpWG0QZRiabhlOSkV1DoIgQXApXla2k9DAHI1XcWMZTPeWhFPpxiI1miSzS42/6M
VRTXNIt4k5GRNqa+6waf8OAxALib09fmxPs4TTCi3gYfziG/XF3lQpytGrkO7jF9QbFYaUcBsxcN
oJIMzoxpiKOPs7TyBw9URlBiIQF4aA0P2zxXdU//sKol2IZxJRj5QHG6l81mHgkcecKLcYJ5T2nZ
sQS3bd1gY0FbW02AnBMaT1dbGTJxRoom7N82QHO1Hnh0hzfej1MG9zwVxIP2QGY8Z/Bpiy0TuYru
JQYfqCstMx8DoFhxy1MwF2CpqJavgBuFAUK/RZIic20zqRTnAERihGPJAUxFuesILrI66QfCerDM
f/yPtPAhcSVqdli88F0tML3Ls2I5P3wjGYdV8HiKR2w/0+XmGmqL0qMxf1XQ0McP6i5M7GHx8K+o
DfjBzkQmFOViKyYaqGn/2Z4wqSxpBnfO9mnqnrrxSryL7amljxNPtJZdco+4JLmwvY43V8cfEJvb
PCOr/5SYu2NtUrDdADMPq7cItLfTlRsoz1sY0cHG8YdOMSR5bj2TaOWcccUsXi3HIfeVvsdyDC1s
saovWCece6ebK6OEdBfx9qfzZT6ENaqE9EAJpS6vSfEkw9IOVdk5c1qT4hnhZ+Hlkf715zWvgMJA
3+wYCQcnDg9RSzYX6/zy5wwHBwVI71nqgAgRECKIpdtqWv2pDNGiv6Laq+GphYW5gmvEeRsyBbb9
uevYkEr/2fEQlSNfZve/8mXud1bDtysTs1dnbbBMZan4W4GD5StlmwcwJoKbkXFPEqLaiCWkascW
zaX/ZjjHahn8AbDHhrjwdUA4Y1kXtb8AB9/weV+8akNWclPhqzf9+Qti3WpHyJWQdMtp+kQKuTVJ
AgddIbJm1geoxMRbvjIAlNHajkC//CK2lmQ3cTYeNb4pc0DykIauXHuF/6FzvxmZORlDiQP/pZR5
AhKQI1DI2ERas4jrZwFbucCILGTcO7zPOPUswSYxP+26G9XnbdDXHLFwMiUh1sxEkin3CEo5d6lu
0RXWbqjG/pCo4YVOcp+J1bD6Pud91j01H1u9C7ZZmWMRIthLbimEOTnmipRBS/vkUaSg0GpIFzPK
RSW1qjyXl2Cjq9i9bjNk2f90f1tZe6QC2q9bCeni1H4g8gPj/YmNoFEb6CXk0iqK3sRAwZ96XLnk
9k5D0Glb6GxA0rw73Z78jitx4RdhYg5Qr58VDfOvO7Pw/nGWYHDrcX7sJk96N0AHoNXX4hxctf9D
tgnsZiovYc71W1XkovvwICyEr5iEpfSRH2WuUMhSM9nSYKiDfiGny7Q5wdCMVxjDwWw5egUgum8E
L+y7QdD2s8eg64vVYDIYbRRBNkC0wh7jZnl0P3I+3hCgtIAMfvIF9Zhy/FChdaJgl23zaiLYzC95
e4W8TI/6WaK1TvwYs+Nr+UjwzFJfU4zTWW9PUpAczzJGqb+/XLsKCWwYg0l/Jlv6SQr014jT4eNR
p5K9aiw5sOwSoSlijnryBPSYNovIhI7toIZaUCaZDf24UZnJjhAk9cRFMls7kZwCgA7rRQDek+cd
dh6HSNr1IiuZFYk+3XfWoe1a1lM2QvhK2OMwyxOQm91vxwcRlgvouh84UWVKVo55fA7rd6M/rH3u
iJeJwlcSf26N3jSPWswplXF3vLRHGGLD15sO8is+k96RFtw1D9CrFg7RHF9D7JUY1tmtSsG+IDvx
2YIiK/9hdsVoRx7li+Xmnljtqs5LBG/3UsSkYPRE92omN74KBcF46GEzg200PlkdegiXio2PrJqZ
ntBYlsKsSOhF3KD/qsAHw/9rSYGtDHtHwVNUZ9AiPOQ5Rnz1IK7h9mM2qXxtiIoeD50Lukzq/sZn
qDMd/tgv46EaMu9dULwees5za7mUf3Fy9GXJ6HMnKV0S/luUDHIymPjUo+XyzQ1wG5+tpezavwBR
Cv0pIBAjbcHqI/FGP3HNh647TCC/JbfivoO68A6GTQH1MEOswm7cy+7nU7BIwDZUd6ZEGxH+T2wQ
hn5RronDbHTtB5qbUKumRynXPigEEFGtjqzcRXBTeJKU4z0r28gXdyoMg/QcGjxUHakBbPJDPDWT
rbd5tcJaF+UrcktYFC2lqJoWXIW1oREtG7ZmzBur6S7rKAPRzxjgjxbE1yu1axhvkvfSBxBpe6Yc
VjZb587IOEo/oRdwCqg0c/BU5u9vnjiuasdO9i4G/nxj/R/0yfKcYMy7duXznTBHbiLC5a7qr4gQ
LfIk49reI88fFmD7TEcM2cmwlxRF7B0CElY5fZynJaKzdM+uSxDI3wzy1or8tgAm2UivuctSNRLg
c/1cAvM/vjj1hmw31sAcna1JSHk4jao85WnnVnPJXrcyTxwuZbHaAKqgD1GCF+F+v5OAzTaYZK0u
ykolWE5T+n0du/2KV+TD2Cgs/hpPfmPUMMNR/2NZPl1xMLX6m3NT0gpVtEZ6Uk0spUEwdjYFJWuZ
tycn5KrELexUwGgt1MsoM50k4issBMm/NjuDp+chr5TnU9d1mJt6osJlD7aAqgUtF7fio9D07sIk
e3mAG2O/nuNfqHQINAh/jzS8arHyfVYm05DOhY80JsAF/2h6Qob/kj9xyzqiHPayAL1WjxnBeEU2
8omchqNivnAGg/aezDqPN0ZOEQqj2IsRXHIYlFz8JbR6x+GipLZAyARsjRXkkvZXpzlE4yHLpHdS
HQ3MAoLZWgwgvy9Bnynz+hi+Ro0Nvl5tgzHuhvwf+TohdfyILvpvNlPek6W+6zagVMr2TdDutQfh
26bOqlvtQwOsWToT8U9J2FW37A6D4665tnW7lnpNC0bNqekbswTyXJcqWyktog713Fba2WARJI0o
rpSGRmBqT3CAJSWU5Ma/RynMwln2c5sCnx7/OISyl9SGD75O4+LC7xENz1b8nQg7oX7k6RdjQph7
PVlq5dr90CMP/RMPYbSFZpmTsIPzmPASQX5I+waJalgQKTUNE1AxrKfat2QHA8CGT9B8vINR8iOx
XVbZuwlOKHTKGQkfqID6rT0fC4JCnQQ7ODfaCI8FwBCPxRzwjqtk1oUt+eRsS4GqJLKAJpLIMC/L
a9i9NigwlvZ8IQ3NXR2CffpOxQ5wRM3M6//8HQyEIWnXeBj4OVNfQnsvyPCqYK53BGL02oHYeSFt
AmPUxrBTQtLAfe70JFJ8NvMAtkH+10YyI1Krmye9ATWoQGud6dcKURakmdLhoQt9Te/D5y6IGRne
+QBCK5tuXGJsPWKaOvr22APw+UwoYEqxrz5O0LaSdbXrXYOqQOMiu98vwIDD/mampOVtLW+lOQAW
ZBxgnjaAU7TbGtG7EzV6Ta9zqmWahko65Yk/FfJwunTjmqc9hehYBkhtP4ixrH5ozFkN5nRePDNT
6BrLDQAKG2NZz+XaezwnWOfLloI1ZJY1Vgod7FvQkhRdGlbyF11YiQhsznMecAdLYLerHDPzJu+l
t5ZCZMeyQh9Lnd2ES9nwb4REWgZivuiN1HAfk9yZfdazA/RmhlQgMpk1pHDYIRjmGU/Kz4GhO9x1
liAe33Ll+kimTVZgRDgFeqMKWQnjsaOsxux6Ir+tBS0eEIO3VjC6R+hGnmvHYNkmWk+tYAYZZ1vS
vDs4ETxR+WsSe6Yev7PFKxt4B5m126Dhsa/5aeUVgX3gFt8BcN7c83mKVXovB1L93w1jBDijmrhI
gPbPbBDy8xYxxvpc2ecGal/wfRy3DVlJudpntko0KZbhWS5Zf8c5NTjlBNZf1e5C4X1SR840TGIw
ByNnMC7gbYfSVWLnynIRUHLQOVeBz2A14tGXbkg/dP5jlC+VkWWlSOEw7I+Ar0rlw7rNGNXYMNBU
+NTatVVhxYaLmnu6WBKQwxIMhZ/ZLfllNW/R/dBJsDD2MkOqzj1EpIo2aTM1mi+FDy4G+GsjiCXy
6fXrcuv2sUnf1yYuQT7aXJ2k5s4nFniweFEQL+8DI3ISd/svY12YacsVm1uwqX2WnKrcuBle5Ka6
k1jflGLxjEy3d95nZMRKluJSU49rENoS0wCpxyaV+GMeUlZZifJytWmX8TaUW2QcmjSsnfv31Yyl
rjPG/3yPd9FsP3EGCjFwOFz77FsutQ0xMWOxI5vXnyLaOPXk04eYd/A5F1BWuNzdPRw7C0Stswxe
ykpxp2EiruP+1ho7GLnRRtdg14Sstg3rxxlA/YiM4+eqtxnKpETHD53oF6BOSKL8qBTS9Il3FyCl
LsybYzVJD4tYytthP1408cvb//j83wSV6vLL3SUSbj4Q7E9/eC5cBTGhEtZQ5mSbSUzRn6Zi2gba
KBl84pL+AbXUQ5GcWZhjN79cVj0GXfTS4QOH0yIh2L0YZeCIJXArylioUJr5FlDpPszPgw9eLMVA
/5hwhdlwqnz8gTAKJ6+JC9fL1mg/+qgD797zzRglgspqGcuXnGzMLxuiUvZF8u/q5heoFiKR8cly
rjubS+b9IuQOuuAbepCZ+153fXM5x9ytEOtf6VTW6GShqqKHzGVKmxF8M0+WEKUCRVSmpIH7GzwS
VRvdbcmmPKTobFgkaynQVw/b2wHMT9zN/hh9emXRkrk/rThfOUGIj548/THZWeCUE6LtlyxwTcyK
SslLAwzXz3Sv+d4ihCsci0GLo38SedLH7sw6szJl4boIsXFCA1lKvmc0gUFBadh74jqIVQZTxUqK
ptbQL9pfSZLauiNqRKERa7LKkdxOL3ridp2SungKAkXIYKTwHAqKXjv0PhIfHpx3d8wwOu/eJJO/
/DSIMv5cR8sjkBKWjJnMLVH6bLJ+kQRx0A3Rim7DNxB8p3+VWGW886V4sDVfh+/lhlATQnoDUzmi
z1++bV/4aCkn5rzITEWKrBdzgVJimXl8fNjvfcfyViP7fKpNP6MSaoeDUrjNh90dwymNvfqDH6ui
83i6UP0nXd7QckTQWOg5qNiAYCCIKKQBh3wGhW/aAollPjIcFYIpYLsRPpwoWnJFjw2OcCDgLXAk
h6JjjAzE3B2E3adHouGrF9rkwBUdiwCtcZ88xyNJWPyRwcwuwkxFrfUcyd641JfSp0YD1jNWxjwm
ZRWAyGwyIhh/OrGJ3e81eaPFTrFjKBqd18lIqCpl+ZtJs6EQvOgugzF6M5Q6+x3FMLIxiYJthwiW
3X/lGZy8xXA2OdfgfMWHBqzhL1u5YuqU9GcudZp3KwUvBdZ1yuAdNCdFn+nAyy5gLHlD1yfwEEhT
0LK+1ARAnHFGCg/IxpBbUe+EsjfovGuy8mItNbTGuj+WwfOXVZxnPyufFGi0xN0PfSHbPyMt+fv9
FjR+t9LQ9mFohj5RJEePQU7vbPI4rdMPGToINAgJ5HqXrG4TfCI2XB8e4B5ErHIz1aIpJ0qWYiAT
2Gl2gYrIYO256NTdpa158IHMCVt32QPaa4tnmXmuWR4za3EMpUfkdGECTR5UgiAMBlb/j1pJUO/j
x29QrDuey0R25pQVpzW8+Ca7TxMgkXhGuC0fIcXZdfST+j168P3EqlPgP9RPTBh08w5LYMHStsh3
VyNd/9zquoVPFTWyz+Th7usG98aW6eO0l8n+moI0j5hmDZy3sR0wkr6MpsO/aED/3NCA8OqUtdny
drlfzunDx9M6yjd3VS6cLqBHi3BvgoYnW2SWam03JpQPTd/cwdjslm+j8YOfL9i34Dw1vdBg9rAM
JOKiYNH+nE+WwRRfOw7qKhChgiEGLO/5fP9+wNvsVRWSNLDQcCGxJDQmHjlRZVc5MOszdn9SeycB
ZK+0RPPL90HpdZxZeqtebceGdfvvR80ndDJfQfOhPj58vmrjK5qTDDMIVLGgVhjYoVg7j8r5WUxh
9zIl1EFcGO2sSTMeRjtdAQffHjqOmd+8Sq0MbSrFv2xk+Ve0FP/XzWXPt5L90C5U/ttliCDEUkS8
a6niZ6VpJZ8UaOGzmr1jeKoVKQQ4oT0o+yda5i5B9dzKTSpChsENJSRudspxYL3TwxK6IRKpx7uw
cbKKNUzcBgJybwkipYTeR9B6PELEn94dEWWVOYfOc8kDcsmlKqgybqp7bx49ASY9qiS+NRmFChsF
KiL7dNA4Pcu4pEU1n64KRh/tX7dsQn7Xrm/ljj6HLPX3m2IJ7K3ZKaX4DoT+BLX0tC/MtC08Uq3t
dySp9UE8eTwP4dhNezGwZj9r0omNqyWIw60j7L8UwOtlFPHMbKYUTs5egbt5G9h0Xqs60FiIfl1p
HV3qrvInMECuueQKQINaqv1uu+KlYInL7JsDAxS0ujIH1xlhyyl5v5R0aeINJCv0L8esCTdNQk4/
89zeLDYn6z5AvFONPN/Cw6gl0NU8MgY8AjmJUaby7Z/sHOuoVkL/8+5Fl4j1oXX266sISY2YJKUa
2bfYq17WfQb+nixfoPzJKYVgN54E9lFCkPzyY02+OUWM5CgLwZ9elsRuokw8zp/RzNlsz61zdU8S
/kgXdnq5mUATtGi0j9mb7MxFqEnhPS8fVq5ILSBYhzq3HY893FBcuuoNZaFjDer0X1wgqmpiJsl1
Wi6HTSDcUPWfNyH0LoccO5/ioBczrGzoZjEAEKrJdtLnKnvVjxnTF5NZ90o6X7tqZuTqOdXc0qP1
wdvS9Om60m4jYb4djA7svl7enL5EPOgjggdBvuP6CslMImWDDpEt6s/EHyzVuB8f8LObn1QoH5MR
A0/IWvT0ueRZhAJbw5X8Fw5nvxbSk0IfLi3WLmj3r9u03Ll5+Cx6ZJOt5m/iftXkrqE/wiZQBMbG
w+hUfuMKrkRLnDBvhsI8uziHCq79F+vDYYNH/S9T+KyNVV2YZrk5RaDH8X+QePoi+jI6p0wJINVK
PyzL5XtzSMOKxoCRMwAf9Rg0bxDPa2F5yQXPeTS7W6iwVVRobwY+87nXO0Xji8GKgS4oS1y8d8bt
TU3avJcG1OfEc9OfEhc7/vTF7M66ucmGKth+Vx73eC/pnnPSKsukSo781/1bl4Umffc6G3vJNM2B
hm7UZhd2G9UUIFbNvM7MQ54jO9gPoA419AaD1YDNkns9NciL2/GEH6+BLaexBZvgpZ+54ulIEgAY
MQGZ51TlynzAfnR3Zj4mPJ4Hi+eIh7hTx41ofbfHP4ZetzTYVHHpPNJxPcVkAcAnQupXsX/4Z8cO
n29PllACOXHvGNW4loshUUxfCCqSisNRm9IaSeto0+P/Vfl0nKy8cDOXG/joibrJxm69kpXFr0OG
f1RAG2fMvJ0tjo+lcbKXRZYZERC63ouJATGFrBxRCeQZ9TW6zcV9IotTHVZBYg5K8YgwjvZMCYKY
xp4zhW92Sshfs+144tRyIsW2zHFKGnmxEdidHIrPPKstyJxq+jXwRAoYfZGhBFuXTST5pMWI/D1I
6ctMQ2IwlNzOr2Nch9BNYyC7cscnUkan3qV825hYNCuJ88Hx8zVaSftIWRntltxaJwdSJLyIeJOA
FeMllbvxCmFyLIlQ+KU5Up1AngNKkh/tqzgyi+lPDLOwOTFv59VkA+SOOTuskIeOOifxHIcMui6+
EjiGfbAvQ1kwKtxaoxgSpqeCjz+X/szr+52FW9x5j9fPUGLycLqdWmwkC8vIHevCYwEPBKZ6qZ37
CY8DF51dgvPUSzhOC5N5hqy9kKP7PY49lxbEUCtd+NknlqY1X4AxlOu5xqHdDuNwRkgia7xqKmuq
FKKzzov0dOmOOnavUuxcE45JvT3dF6ROJMc6hJOET8HaUJyTc2uwVxPRnDW6FN4UjavI8fuonOA0
7WHV3l+7UtHI+YLnL2SZPhsbA1HVTevcWfDga1OqTj843zf6pRcxf+JG5+sWljd9ca9MWcca0Dij
2RWyh8HuU+6iUp/mjmB6SZRbNvhTxI0As+uaKUbe+V50k/GDsXJWrxw/nSQZoKuhSUAlErOpW4Yh
rvWIl/V/YVQFMIO8GSlpbEfhHn8bR7hvi1VjlV6a3qL/gU3LjuvTKq1ktq0mPY+y17niWx7Lw4vX
U54SpyKl7AKLdH5iz1lob9+UzkGsX87eqO4DkXHlF5a4heUxAjeMFptMmgCeyAKIy3OlVpPNLb47
2uUrpSkYtvjhYGB59m1K+baAZpo6gmj96ex0Wudc9MtCOP5+RbpPEMxESkqAduwoaH7Q9+cVZaBf
JKdHi843K1nBG1XCeg/PRCV9bnrXy/cskoUC6SD1xpfpKf1zIODBqVIble8EAqqcJyE1xScuqzde
wLK6OjinzO+vt47vh9BHPSLGAHOwKzVdmmEqc8V0zRa01HRTr0Y+aNDQ3fH1GflhWbCwGHxUXxxX
6BrYQNAH5XPqROXStQjBgHdCZ51HaITcH1MW78l+QKgpBe07iyCN+0Y6AmMZlZ9ah/Lf0BmqDha3
VqufYM/H4MfYDtb7rMXXYUwLNBi7ootokmPYos8362CiMN5H6afb5gQvYhvtJ7BdN1plu8d2Vfok
DQCV0xbjvIEV35Fl4Ase5Bxcn+b34rKqjXwQHvP4XLfuJzysWXN4z0aM5K5Fi+UaJdDwxFpQccT9
ORFdg21joS3XAp94R9qpOJlWd/nwzJJslcNHAlQ8Wvx0R/1l4+/zJBmZL87CmcIEvmZecTi7qmmZ
e0tjHhPxIj0LSEvkFzxg+SND56WMWUClAs6i2wAbn3d/5ACv/hCYrXYDdORa69iCz9K0cXIFXmDv
ySQ8sBdhr5hJ1g9FodBFqceHW+qMjJjQrNZlw/1fBbfhWyJlQ9cf0nluZMLbIB2E3omVyYzo/205
5gDSEi0XsVs0x0eHTR05oNzi2gB5B0hvhWSJKcZwwi8+MteqiyS/cqbobML4VBoO806GaiRl++3b
jgVNoF23qTX3h8XpOxYeYYtrAAtfNt9ijT/jUacF/++mQDp2YCLCpzBH6CIgzxv5WN/SdBBUnnvM
vpBJZvtL27+ncEdARXcfb+dLgRpv2+o2QGZdcdwELsHM247DDzzZ9afcnxCMYr85cZ62jdCudetu
qA4/x8CPe8Ujli958Krv9yl4s5DcI3bp0wfT8mRJ4cYJ9vBrAFCPUT+GtIQB51Mx9M94/rXduUFT
tSdnFnE7kxrFnNUC5MHT4exwRfZll5lmiOGe6uIhJFMSG9ARki9rLZ59JY3POOumc+TPSQ//z/HH
1Thv3XEEfFy5LbYvbE61aaUArYlrEqGQj/H9LeNNAjl1Z6eyCReVzvri8chcX8fZG5q4AkTywoRR
hrT5Nu/17m2aoNXRaR4i09VrwJymzfZ/0p/Ai7n0TBvfRJNHhn5F7b6F0hC7PpJazZ6xLOpS+AA0
bf+tCJBI4HkY0ehjmCdVf26TMygwMNjOV4ooO5iW4o1f7ATRFoJP8+p6GTFtltVoJofsDBaNcEUp
yshkz7Ym+DZNH/WMo8OkAuOlMtId/0bBSjjstQClylTrLaOIa3effyOYRhtRxzjfWVhJi8SBpKA3
kbTkhwhk+WQq4Uu3auCV0unznE7U/VP3dw7AASWa1fz6opl7lQGZn7XBrpSiL7uIGQp8fkVZe4sr
CjD9yCV4ClxTqJCAMDDuTuBvlS9R6evzLLHhUWktyqaiweKX68vuLN3L5y1RhOCuFQyKsk8lOEON
r8ZG7OFOEIoXN1gH+0evfHmA/84Vn6kO5T/yNyYvMAndI70OwsVffCeEgZRuAFdqdC3ScE93MEPq
v7pcsxGFAXrsa8MdDNoYoFC5FxUYN6zFyFENWv/MA/3jbtnr8BKL/hXoWNH4mxiYYWfBCSESIlpl
moSvg4Lh2atTZa4gxkYHVfuJAr2K/oyduBb8YnC0u84ZG6+5g5/rISJ6l4VvmPYhSXqK4HfWmbrt
0EaqPUIfW+WNRJoKUeV1ZcuKNkGvK198gzX7CNOHg4xxPtLdcpXjLXGJE7btwxoD/4slxWbyU9d0
//CkxpX2zVPWAHTyDv5Fjkrp0QZhy2l4GOWjlNVSMS9Dlza9Fzn1Pmb5C3CrWorP5cJ2Hz/pVixB
CbgvSCaQiazmN3zjNl0DuHmPIWaqoD0/no+teDwmg6ctogpm2y8h0ZMPwI8/e6Lphwp/oddKpken
712Id1N8g0fgZCBCA2GhaQ7Rqs9pnp89lMke5Ca1A5E4dHgMWTPXZxtcJUkbaR4K9HS2WUdmeUdq
wLXJZCO/ccJ0e8oG5QmOQ22iQezCxw0/pvDZ7Q3WwH2sS+6aSsP/i1O2Y0RCgbiY+rF0vrWOXz8P
h/WWnviDLSo041+/gcrvUnmutrjf1iB5oQdI3Zy0Sabsoe84qcGtXgXsq0f3Evf19fciAFsMkgzE
J8UX23C0amR6moINncRqYlcP78DwOK5xlS3QaRjxx5XCTPkst0cQlG4AM3EbxL03xBp85jpi9ekA
fOtabWJVNrPaoNs/YW4y7WZ2/sddpMtqiZ28pu1ivKxD08zLzf1ZWNXD2w6EChuWwwmApCFk4h1r
kHqWlkdmgeNU49bc2+6WAm2IQANxUVBifFfptq2VX4e5AjuqS56JxF5jN5LjM9FUc3r/Y1zMJFv4
W7tRtvQENJhP/+VflWDKgrxW4uR24comsOxWKb9QoBDfClfxvs54bzIjm2MQ9mAcqItPNGgwFeFm
Amh9D9J2eh65VVjT6Bvs1xmVuozG6BWAd+sg+lMIFOt7PBv+FTZdlC3xwitc5Oh+N1oAnnAe+vfz
7Q3Z915lmUlKSTBSEFxWhOINraxfSAXLkoMBOCZ+RkBE2Bw1OjJspvluBf470MiRAfmTYu5PssiY
U05Qmxx8k6mmgf8yWkU/VJgfmKBOx7hMZnNECVu7DlamW8AErO3owauJ8HUC6tLGOo5Ge4iBJszk
1/ViiN7nr4KdbLY9Xhu9cjVnlJpvuOw0Is7JTp9zEHilg0J/DDIxyWi1cfoIBmAzeZOI0mQ5Uk36
F6M8Eklf1n6HRASL8RneDP+GxFIn4Enb4zOCyUIBfyqo0TYtiuUdqldZz1BSicCZ3S/M/0+8stHJ
dDsiczsmRUXtwzMw31igNMl0yX0xvw+An1zcJ6I5YQebVbe131m8i7YjFfZDGCCbV6LiBidf0e2C
rBLMK9sxQyl5rhlB2lWNykjW4zEwBdd3QbCtedKgyIqBytCjJTUUl60HelhHh3YZ88IEBYyuY+ol
8XTHygyPI0PGEr8UIQkaVBa71d9UMLUfkmyf4BHeszCKW1di77sm9XmX+0n0E8bRwvOkCmbWXJNL
8mbcT/0d6ZzAKpOvEgeUEzcCB8rbQA1iNxrrdpOJtr5FVq+rRQ+6P1jpBtmRsTvbkZQ0BAv4RZrR
DCQUlmeRxlestCYFs4XYqdx2ky3SnXnigZm7QGf8D+4b77u2kmoB+ca+qR6YwxKYGhkZdJWUUjX4
ucSH82/R5rEztqJItsEYhVZsFU3mBng+CK++0laLZHPuE0h/hEu9ovStvKhK+dDxp13OUHDZndPU
rmLdlii5MAAZFuzJi655trjln+3ADZbgZeSb3jqhpnq+tglaS9Q6Sf3/idyddbgO0p4/w0uoUX3m
lbl5vKS3JtJVPYNGkWW01UIo6nvOF443ogI7hq2KrhRGNcl4oVQgGnG56shA3VQrykDvSQrNJ33M
OBhikHJ0G4/5itHFgRt6rMSV4TDBqD1LfLdFZiCPqIwxq3oCrkVZZRw1SAJ7FZ9jGKGWCxMj22tV
LcOZBqdVDrVxeqSqGpUxo2W8NGZHciLchGfclKBxDQuDSDcwMKDIV4R00HgPPB1kHb3nPFpJy+YK
NaTczSzwjdY/DnUT88cpmi07g3tum64xkviU1pbVHDdSbxii/RHqECgC76IKNJJT9mqrgH7lYJxp
9AvzMHSICQ7ZryOliaGHp8WSCW6cA7GAdHBIL8VxHDKuzkRJNEVnMkhtCWbirY9qqHkG5biwwVcr
ey56pgMeLKyJ+XsJ5wS26SJXiYz6lq++1npluMGNOWLN0oaUUeUhcaH/m49OpCSx2ruUVP/exRl+
6TVUFLvvqsDtyIsbxKxGEGi/AzN9e9dRuS1UksahzJOREAHf4h6XKfQPfutGTwe0I5HuyzxpFRK4
O0G/k5FbeibCtFOlXVZlVXyJNHJgpMOVuBXmXb9y5ha1ofxbjSb491lTmdcI+2K5B3zPsWoArJyx
45U8SGmTozcFEqIRIegYMJq0d/ow/XoQFJPIkLxeLNwN5+7t1QGt21Yo8SypGFdijzesN/CAxbJm
LAS0Te4qhbOfnZYTrasdlOhvsuFdH838dJMVzderkz9xV9Hh33u6/nBQ0geba5rCQWfEd3NCUYNS
VcvTG4jpd+XGjoXsSXVL2eFiGiZMB8WkLpDVmm4McBc+zx1OqjekQU3bFmx40ndxCF6nhaj4eqyi
WWvm9Gz4JLOvLzpXnW4r22AWdq0ITeshMtNdIS93EXCWBbqSYMZFLzqbeeBJxYbSNeR9kzseb9g+
sBtClF8OT0Qcz/L6Lih3BNIgmg9kRpfXp0sLLHYuP+jDhFAcLSRihTJzWebt+vzz7dOyJrWoXUr2
NCmpl7o+zVgwRIUMHosELkezSyD8mJGlmXob+Fxpb2JuogX23HeHyPOzFX5xqBVtbNyo1qMJyqzA
b49Tp4Z6avThChDWdkh7joCeH609Tul0vtj7f0PCpI1p/XFykVGBqaoTgBmawFEFSJSqkXdFmj3p
CPa3UqHK5MP5TL6ThEdMYQ96N1z/FygNUAilBybrgk9edxGA+eEiLnidzMemoFlRpa4saYuLcuTY
W0rtS0oPpqGcFr2GXA9r2c1z7rRsGBYWiUElpnzeEvMMd2q+7LPD6BlcWdEWpfenF4hzc+jPrVSu
o/zNFICExMuwQ33X7/DNTI2+vUI6+aBQMHJSTCGLEAZXfiZE+wz/aETxOQfpbKph001+MJHwAycc
rH8DlZF1MAAAn06KkQ5wRWNiOtkbWoPSi4NQyluPzwkx5RbCv1S1cg3l5qFdalohmmwWxbMpCnVo
rYtAItv4mKeHoYYZAjkJnebenJmWRE7qqAPNkc2aPObgyjJeWCphyd8OvYRNBp5D8jX9WqZHwBIG
U3GGFX6jagJGOVMq/kBrOmVJC9wj1yaJLMXvxEwyd21dExpxHnPNdtQUEepSukjRKb8N81q6ZWji
1CxFwA7AD5SG4TEzhF9++UiFXzogCiOF6xYkWH0eDAtSx9I/LBH+2QctMRhfEvfzFLjAknuNpPzk
ZfC6plYkCz/u/v7giSXG2+vnxhCdUrC+m4DFxHQ4G2wF1J/2yPJIBN7n6qB24rOCJ/OwMqj0O4Xd
JTdGvpmFiN4xD6Z6cSNOuvvywN/NRP9yr0NfzBb/De2WSe0cIL0Ok8QVEuj8wpo7k5WPwbvjgaGD
1Td5qcod9EPix6RbsPD1Oi/3vBqt1wBL5+KDLRUz7nlCgTForntDmJXdDFMvb+QEAylTsk+n22Lw
B6qYIJ6Fr5Ne9AHNQnBqhCbDpZlW8LzcuzMR9tYfWEWcmOBwTXC4kjepqJ170DRYmIEfOSvOiexU
cMB0YpG/8n5vVJqDgYXX052iX5ZbT/EnUUq6uWsdh7x5Z8rTVe19A55az156G2AVRuS8l4zarusN
cBktYpRvokwz98s59sharuEcaPeAVgB+34jYh/sSubcR6DKE2bqhsaLG26SZAbKi9y9VZoelZ9Db
0gNgRs3bsRhSvO19pBUH254ih0ED/RSr+wTnFpKGiaoqvRdVIWD1QMMzxL8EJk7O2D0Z9Po15cNa
VMAs9I7OOsk42qXKk5TG9VHoG2pbwfaYn8FVGhcgfK5M22mxcaEiVZHiA97DPzAD5Y2RpKk6dqOV
4bbimz4kPXtCcWGRU7b0OLccxeE4NlUc0+CpEsWcpeq6dmY0K+JdoAJPntLOC0eb2LrE8DyFj7aC
6n5Q6fuSW158ay1NTan/J/GTpCgkr/6bjX4tlg4r2VUDwlgw4Ejs+Mz8SHG9iuAVNWZUZllR+EqM
O4diNavfGrkD0fHhrlIsWfKTgtOQM3M/iz6KflDX1mqQPXmuZub4H8NMwdDwEWyh95ErxB9vaVs5
Hp49cD1uH8iTgmuMWgmPf52c9Iu98JEnvwHiaZS+xx6u5V2zKStnK/OquRa/gv4ZjD3D9Ry+q4hI
yq+OzvVKPmSKkKXH41sTipv2zCk6hJ6Vf2ADClP7jTPo77cFweF5yrCINVuaN5fhWx602Rm2BOaF
n82vKyss+K7ew/mXVgBtDGlZjpKFAp5mGK0fSVEW6DDcQAwVKtrATszzFsS4n6M1I6Etpv7U0J23
JeUEwFwWMVT5dWp3ht+nUo//ysz8RNLzGqD6YNL+XJH0zoN/8ffdUA5niR0GZ3Ewi9qXdpr0MFX+
cCEMdOoa6OcpUTfRve4/NITbXGggvlJxnACTGx+ybs0pXiJm7rKPf8E6l1tUyXz868Y8idn/jd9q
6mc4bRhRe2ay+r2xEGCkJW4bS9ahYF9Sl7VqUoiqEyyfoPQbSz5zqeHxhwwhikLMNykVw6ZeL6h/
gbfvhnltB1De037ip9gecwYU2sG60DdLSXVyChBz/ugEWdsL2YHHXVR72K6Oad2mWkjlj33563IB
V7/p+yeJCZjnAenMEQ+8rDVZa8hZKCso9XlNCJiF05yBWXqzOUJoak0jq5B4BJniN7QUUXp5W/ut
cwoyF34R80NvQNYxgdUL9D+pMdx2wmHzYtoM44rNXiYLtscFk1COMLY7MveMeDglLp1pvJca+Fum
bU0luc34V0RBbUpX+Xw+yKKxeUcc3dj1cvWC4+weEKTgj1IBDhqDV1LUg/5dep8q3qa/AAxS6AY2
oUMxRbTfv7tO9GbT62nBDd3Vx3LmsMr1h+wqUNn2TZrGMlYvGqL68yt55oqrVk3k7iJ6VDpuMt1O
X6cUfva/TyTL+cgzxaOEiNNjNHpAZaNX7MmtELKD80D2pKrRAMZMuRssvxv/DlE+aPVlbozQPeiM
nORupLPJV2GNcgo+Y5quwA5Wwx/NeVtZIc5tdyHz3CA48DXK/ZO2CPohS4vmuFJ+uAoJnx8IJPdo
EHbGvrSjE2K/K34euj3LlHTLelpKiO/gWUQiNr5n2pcA+fbb8+n1fQ/THiMJOapGitDi8+ofLLjs
HU3aY5TcNF5kwJex/KIiveu/D9FkHruOVLZyT1x36pFPKZwZkDEbYwvvlBlZXtPpBL9NnhCz0i2i
Gaa/VKPJ0hJHsUZLVD7nwpEsqrFcNSjDJCWlkSslbGCDUnSHXdZxwx+4jtasLR63Tf+VI96su2hl
zFGtBLfj+bAy7VbamUOEKcc4TuxpFnEINHEdAbKsLYiNxPHItpk0XgzqIK7zpm9YP1EJpVPZf0pa
KK3FfUidzvmBSpWGw2OQ7PGLZhOTlarZL6neJyOQhJX4kvxk1HqEL6rPsdqNIq+GDNfpr3zSwiHE
oUgB6T30uvBH9BaKGMsBVI+7r0D6IGxnHNT7hY0r70Sw/q8Hs0WTLNf4FegjwiF2EQ6DtrDd04Jo
BhLTS/Dvyh7ye8M647QmVy1h3+GzQFVl2Ts0dZHFsxHvCilwPY7OfZQllveul05OiE4wZaC5joxO
P3ebrDAFJdwtQojIICC7XV3IxUdv+l717KUKIgKlyzHhppVfOWjcxJc9XT9ZS/X/yhUHoGLitIRI
iVahX//RCTBW3wmCdGyLmy3yH1rKhcYP9nWzfeJnFtRJqApT9yAF0LWpCA7uJ2j8wBcAnj44GRxh
kwZtRx+kAy7bHcS0epFbuc212TwPzkV+aklXInIq95LSLXb5eaYrjGKsqobgkaP/5E6jX6H3jv/x
pLPftNdUdaLh3kQy7MhI+fh6KE2WpGMOvhydU4X5ii/GY0yrkQyKsa7+EAunvQ42K1CO+amgsL6V
FOWGvNviYus52eRgfqjOOpNXX3qMe+FRTvvvnEf9+vVxywo8R0huSV8TZSafWMoSiBuzCIc8/Rhc
dP/hpSejIXMigDPGfoClgIueWq2pwtPI+hziL2DdLsyS0slBfcmqPcR1cGR6ubeMQBq2j//UiJAS
TFQDfAbOthTk9ueXKa3RvSPBELiqgcEbr6dNdwV48PrdxPbwIQJKMnNL/y5AiF8mPDAGzFNoBgAY
xkGD9YRZUctpuEHciXiNw27m1hK09JCFJg9ABL5L2X/8uY9KBO9Q6ez3mO9bw6Zu2sdzKXNBesCp
SxyqiH/rDWmy7FLlpCNfJj+0vVEWlHCMSy6qAOv5SkGmZhcK5ULGz3uDntMy7JALVM/+7bsYDwNy
msfd+eZwW8RbsIH1kobACOhKXHxoQERNOs+oy0oqYJgZbkQjt7WiQ8KZQ4nDlZl/yOpXEcWEdEXv
m9A7lTy42S+FtKw+6hVNN44tqmSRCHjwX1Fz1XgiAt6l6Dpr5Dx1YSLXTefJbf6kEAcPgwZFpkHb
5BsTTSSWLWJBsQSkSkJUZRxJgBnUTTYIaoHGrsz012nQsENACfEOzPsogLYD4VxIYZx6ui15VD0F
CWh6t8htrI2H1je4Yokus5pgmvnJ+DWmZW4/yh5xZrTs58h0Yb2M3S7RhEBMfn3uEAWAeTPgkpVA
CL8j/rX6TzBi/5VLIfizTZJ0s/XmeiyCLuCB5I8fwFucSnumReKzkceskeSfNP/8eOmZnknQyZNw
iFH90nEdPqpYuF7kBeaNdaWv//x3Xbofq7+H6M320heiIJJaSd1yiCXAzT6psGdZtQI2bth2nm7W
uUrhGPqdQH4MByhxLxmrb9KW7IUttPZdKob5IQ/lXJhTQquVFBVkvGFdXoTGzRpZOoqBmZVxw8GT
CFBXTYGBg+h42XnxhMJ1Vq7RfP3UV0oFDHuZoVvSSt2LiyMj+tc6U0SD7LSkB+rhY/Xzy7PJXv5U
h1CGsUipp7v/L3h2/e86FlhU8NNGihuFQItgy7txHxLihD/aNbqmiCzxBfm0k7nXPypXw1B5D2/m
gh89g3o2xzwWBAnzS8DLqC2FNyIgL6pXmm/upkEdIIG90VFI4b5cOYOYB1PwLmAyFbrHN12o1m6G
anYOMEF4Z3Jg5Il2FBiLyI5Pi0Z1bEjtxnyi7/DeaLumdHhTI+gWAmQk31DhyogwXenNX7qQlGCW
7Uw8DIT/2A/5ER2GT+eQuV4gGqyBYDmL+eGLFKQjM4Q6AaGpTP362RfcgnXKKMFX3gC/mHpIngti
4ZWE9PYcpLuWcwhllhvSKElSGpYCRN6D4C7lUCDn+yIKJ9O+J+d33TXctp2jCB1HiD3XBRq3Y/3D
O58rbdibU6pJG31VsP4axg/H0xh8D5fwVA1HdUsGCwPExLRSrIuWYupZwcXyPy6geSsPaT0PneM2
7GAnVc4z+h0QM6/QOXrdQMntEfvCPNOktzi70UdNHOWrbyNQ+xgwgTqMOoa4JLDrsFcKopt+LhIm
DNnjNGPMUsHRO7IrEfXDOvFs1dL325b3y8sBWQUwQt9IBOzG1Sx4JBKm+0AdV/Duj+ENVciK9IEf
myMdv3XbbTwArPg2clvGeZyPpttrSJIwpCTOQSt59T/K+ZWgShNmhiBg18txSHgskCqhszGPBgEH
2rbXY2D8PbosMa++sOXzeh7lHFhynnk/au5q+j3WP6lpKiQdnfpF/5sHGdxhCmmqMlOmBnONh9T6
1Pu00EGzKxweNJQ+pc5hkPY7tqZIIic23irA4Qg+mIVnkIX15fcPM9lPyJZ3LeW7WgltALqA0mLE
61pQoMaTw5sE2ZdN4NF1JKhot0Wup0GXotkccBd291RGsKhJ5VakMI3CzysrURTIdJVBAExrHCAm
sMmQmI3wLmg23MAnZlXyEXQumWBOVJ0eqdBLMSywC+1wyc1u+DSMkDlpO1Oij7nRGpYkDihW187z
GU7yi0yePMdWSwprvfjauznwvN2i8MVM3e8YxBnsXWeaketdQFhlZcBZkcv+N4xc6rFmRXpodieL
tLW6+/x9xVyjSnp6dB5aaYxu0WL++/TZcJDeIstfIjCDZaVH7zP34NW/IwhFwHLdpeKnQQB9bquH
uTQWcYC9jiOrcVIC3EH4FqS3D5lSagN7THHt4HrF4juVeGsdAxxB1wd8w4/j9qBC9wQrV+FxvNej
AYSNdX7VC8VM9nZBTbQYofOpsG7tPmuwES+d30SqO0BAheMaWTefelH8tAJkQsOvwxqcB84y9BZZ
ajH2VcsmxMJULFOFsTALkdMHxwnks9IcWaqAp3kTb++YXDr284kjtFULJshXWMOSQzyXZ3mDIjss
0ce61CYFiM4A9mo/oii0I6KX7uKa8PCvZeXEY1z6NwL/Goy78YqJysA1oHPVp4oWczIAiHdbCut+
8asyb3nipKtoDnq6vzAatWjOCweedezleKrTle/vVJnusrgQ06JND1+pDqogLtvgmNDgVkPWY4Wd
+r11IoOJ+YS1SrMbXoijyQkZTyCr1lSRpRNeJ7PpiHupI6NB4ZkRROdCgN7kk1/FpxKjGa96QP4l
gZS3nnFWH6L9IltWj9z9+bQwJbqo3kOkcozG4S+OBMxAGhDFdTsEkOHy0FgnBRbh1MvsnpG21IHN
dv5oYRYHI9osPk5g7V6wkiBZxg4kM9a1h38TyNS/8igzTWzv5e/N5Bd6tqMV++CXfgcVn0jt5F68
4BcALA/L1ifNmTIuCXZaTD0dSiDTT3rmCTF2Vgc/c5si1WLqoA8LtH+JvYWZCivyki3J9wODm8by
W8zpBwZpnFYfRrUd37C2wCR8UD21q+hIZVwAqgHQZfBmKHBDBOBT+ngy0PszXkxDlZsWpuppp8Bl
6RNOWH6zjt/6klhYk1jzwKj9d0kv9zz4siNKmb8qI+Rsx1DWUvyIkIHpDTVNz4PCE/hXWlnGQtO2
yQIXBkM/k51gJKuhTnt+/gSlFUQ8NdJrk5WKr445RWc3rbT0Y9FL1uDpM2CU9RLOfTx5cNci6hFm
r+/AV9rV9eADB+rEXyPFCDP/0RGg9tH8OHDZloKO0CcmRNZPVF+dkEHSOG2jP5I9VeTKOznHlIco
kgUgbEcj0mizWU2xHjLp0ssQ2G3hrHz3fVxp/KXTaKIYKg/tJaH5cLo/ATCbAyHOawoxSalpSvMz
/IqfaT9G0DWgHLPGb1qi1BqLx9TAQqdTQQTKmnXYx1dG54NA/VljfMboadZBMAJMiKVuvI6t2weP
PtjFXZG5fG3rerC/PvUwttKic81Q769H9ncxkLKXMl1gAh4cFquINH2YYcNyZQ3C6YT0qyBDnNOp
QkqJ42V+HRb5BXYlOMhhOyXbeRbaF20elXGKB2KTh5ClPclnTrQfvJEV5camLI+UFVB2ig/b9yNW
MPpPIF5r/cFKGDo7T1FGJruD00ZaLfzRDpWDEICIyWIrPG59hbFROnvlecENp/Z6O9iPJrpdUVxj
udQ4nzduLJlviZfELNPtr/0VUxD7IRTf6phuqPIVJEzylS0wSTdYz1mjpe9MrHcZ0fBrQEktrSv+
9q/MzCuFdEBTQvhXZ2VgC1itjbnHSL0rs0vSecR31nP0QS6YpI0kZs7tWCw82y1VJjSmDQLVOdRI
B7/xIsqVTFJxEZaXBTjQ+PvgoWEcrMs2+mg/06lnF3AtK7CHeVmNrVlt5Dt7XqEJBEv3aOthi5sB
yfBemAXrTmhSxTTfSXeBZbrRBoS3r7cTPFOUf1W1ITAPvtv1SpWcdBmB+7/T8Uek6mnEW4sjXNcQ
v88QyixCHbWQLahFavtduJx0hzeoJj6NIBvdpd+lBZZG7WKNyDYI+kBcdw0oHvrFJY2oszvxxYQR
d9AGPl6/SKFpbLOLKzCw9r1b9YzH3RRZ6zyLMqoFHHNi+8L9JOTM8r2V4zONmI73Rlvo4zptW/cB
7ofhtX0iGvaljxi3fYeuXBkf53MmY1RK4tFilWlVJ12EAFAczGYabL7WB7MlDQC8hEHIiYAVfYXI
h22NLrESwXMjAH82mXKg2ftm7tircM7+sbKgoSdhmttzQLdiP1FNXY8q9xlI1z4xQqic7lASOMNI
xEyn13M2pTGYyqeAMNHKfbY7CpWt00RuPpDrYYsgGTHIFPKnECiWkOIcuJ3fHX6OZq38/jK7PeLS
mVGF7vxDyy5/NY7jAfmZMoTV1ZZW3TjffbKRq6MalJF0DiDSqKvaj64RWLOc0dB32BAKYrIBl0e5
FFVX4dsDwBHI11UNbHbbtLmGOaqx/C20K3ImRB56I8wUt7uEcELc9AmaGCwlWT08GGdj7RFJBQ1o
p7dOBzYqgA9wvPkk0CMVeTnf5ZERY/GkmbD0plrY8GmqGeIJMQqvH+BtsmvKcg2kV4pGJ/bXk/dM
hZrpcdOyMGgW7Vr/Yz9ZRlogSfb13wCoUvpbGnSAdj7lKzgF951pKRktDDHCPk/GZHvSxyBgngNV
hYsjrMgOBDEetbK7Wsafi/8rBUi93c2DDQuVChNfiYLH8q961sfu8e22D/LlZ867ms1aHJb/cgud
aqxmFkInLVllH8lDkrsVml5LeT502QwZDD42+y3aLv2+Xo9uWZKuWWQM8c0CJhR7y74zepAB4CCE
WvF2gdvolrFxkWByBfdpXn31z4evf6k1gJz4BRJIkbZ5dwQRbzk7RRJczUHrfkYyNB1i5me/kvss
jDsH4H1GW4jPaih/rP/e42iKgk1pDS8Jg2UqZZ3dBNkkCv6fYoY1dimEECvOInkjiCbth6X6kP0J
HZdQOOjpjRWBypSdwW+IB2JE8553jbAsT9MtlfuLfw8p6baRn9lPIoHyq3YN1P2m8j6TG2WbHErU
amBkLGGTBveM+V3RIHY/cPbbkE2p5kEC+ZPMXObeR3Hjud+u3TxApNgHtu19f4unnI2PtIxhdouB
J45jPtreP7k/fgEis6Mt9PnzHnQYP53OtvikiVqXmc1vxMk8Mp+cFqkPDqtqlxp1NChGyLV5clgl
zTajWRS1UBgHMU4SD1vqfC8NNA0Ja6M2RZ295jSSl4X6QvDca6Te+L8X0QQmPRRMvQoWK9fEfXav
VqSGccZU46ks+c6CllR6b3fzcqfJUFwmtR1nd9CZPWiT4YRKRQp5AalhjWratlKNYyNBehyq3wgI
Z1ue+WAJWz/hMRgUCg8YnROxMsmvg+3DehgqSZAC1LpPKnAeOTiO14v3SNYNuMz+ZrwIdhT7n9Va
DYy4zv8gUObWSmBXIKraNKkb24b6ok8R+XavVLidOqbmz6EUqjwgnf2amWELJpCaY9xZlJj8UdLk
Xt8lWPlvy8unAPPTeFJ14nw5ABgwEe6YxuVgUNywOP4B0SI0aaOX7n1EGXH8pNEmmpUE8p2Z0pU8
U/+kt2Ba9tNWg9vkxtY4iHDsoH9kiO19NTaxkgU2wym32yVjnV/DZbF3zDJ3rzobnQt9jOwN2Nep
v9azkXgxHPEHvlf8oRBo2lksmLKuPme6Fp49Lx3ShH1mfjaBRtuMdz92dWuv22XHA3+drkQX3wbm
HY+kod39R/TWQfMSiTuwzASBZl7YpVAWCTdmfi9tQ0O6fHaOD27gn+hyvKhoL04TwOB7cmBKZWpR
TZu5T7Y4I9GxL9g4NA9PcUQiy1CFJ0S26GW2tgPdVN0Nj9hlDZYjkuiXnGCeOo7SJGp+t9fF4Ptv
Lcsj0YiLjZuy0R6alnGKCO6372X77MU2RooZ3eBeMAT6NYfrPEWQXRn7zf/2IwcdPePn2C0swBlS
ldXHG0LD6C/J1O0MizJoVJSMvC0GeympM5YjmCWLOLLNM9GkajrFDOeq2jNUciH8wwuGDUR3RDch
L0XyDiVZZRPrQGKSTm+JEejW89638GZS13WeRiy85w5tsrP3cAJe2ETzceDgxVQFP2LfIFFi6kVl
qo7+S2yP6lHGlMfY1vND6GKsNfdSN9dFF1oQlNpP68OtktvJpnu6iEFLfqktVT4DbaskKBpCa7LI
4eWQSmA5kcgTTz6OMV/Ag1boHaXDt9XFWS7EYD9FONIrv/quPxBVS/mWvDgLRqniAqelEK/Nb1Be
XpBlzCCauOmT1wVDP3T5qtY15waY+eMqBzk6zsmEeZchlB+R3oe5Amhq89vM54eyD1wXHXrUOmsH
QwjwLbhsKsTLYgXBZPaBMv3QScKQXXWGRh9JDYI0bRNIyqiUQam22smOglFRlk5MTcQ48TQo5EOk
HOlQ+v8cqdHICSkHumns+Nib5Um0HNMHto/grSD0MvxtEP/SG01MbFXY7q0CgybUh5VMV45+ESil
pAPnXYoHFhblfbBc6NoGKgXaaL2g5qPN6rnQ1irkZEyFna/lLO/49zXP0nhUUowqEO8cxN7JlnR5
2s8Z7kRo6giplsnqskhQ8ztCoJ/hmuO7xqWaOFhiiGshtaD7+bYnQYqwikEhHuf1APjI3oTY/tRS
eclwZlooEVv6OTy8caK0M3purSdpzqD5rGyCnGmyq7YVRZI9NG5cdsK0UlUfj24XVwssFjjz8JZL
L5DOy3fO0EVVUsTAEOJxBWMFUHBCNMwINYOoynKTQRoaV/pVoR7Dd2nGA/1+U2HTYym+wn7nZAiO
lAdC8/GydZXMq4gC4wawQw+aDA4U3kRCqoM9JxP81uyLO+NJ/2iMG7TwRircOrKEqCHcamVcTiIk
ApZZBkv+V74nIh2iXF7R/ieZTKcUK1AHFy4crLTkm34/Zyu8veaTLJTuHL+jMCMEDCViflERMCId
2GnxcauSRzyUGixkycs373eYBhEkFAKavR7L5lrCIlL/vzXWPrU3R60d5rPtF/j4L8nProxxVlac
0RRWwRGFj09SeRQG+eZoQf1P993EjWGkud290IdwADP/Vy1c0srRESM8NAxMP7wq76VMZ3D2mjIl
8X4qyloHuJQlvWAGUdcCKCyRafDuD+qxBLRxWq9yj5yVWvZ2Ce6ASSbkGwa4leXJ/vG63HHD8VWX
Aevt5dcRsbI9lLzl8OvkrmYOJN0M2mRkT/QGbpAfE8ATeZQjx/oX8EoePZkhjtQXCmQMiSFj3bO1
xzP7GXdCDjaumvL8F7MQQDMOGBmhzYwZxzyv9kWcOHY392007KEVYzIlV8xAz5QaA4UyADi+IO4E
k0/1KzeZryrQjbqI3JpkUGx5bm0bFLDFclsylT76YsFqONBUoH/jSPW0A9jjpxiciqBpWoy1su42
vtevAj8KqPffoLBlWcbmYTSpU9OmC3JpCDkul5eEkBekjbTyaetkt/yWoj1NRyLu5IZXwDFH4wUS
PJxZ/HLRYY3dq3PpwwZNpQP6vycZeWPNukamQBKxbKtCAnpe+PFghtAWMl+3GXxBQx7QXzyvtIHn
A6IWnItqN++Dzk/TP0VCjiro36Z+1jILNd5PUCS2eNHEr4BAcKnIZcu0oeOUzHmVcf+G/m2VXvH3
YuEt47baue2y1UB+PwEsR8xeHKzTk2qvbOyrJUGd2B5nAkRyphIh87Re9oIkJJ1iipDaI3WX0vWo
GRtPd/sArvWy7M4BMLZweQRC3hcrUCKn8vC2JNVmwMp7bl0wPew0r+S0ikV3HQmXs161RPrl2qKA
6n0DETNn1TFSUDRtahswJQe4EX1DMftjeuJQJI/EEdSb6B3ztiEwdMVDoXy8putWetDypI08LfdL
ml8+z2gsQSFr4tq7bGNvTFlKecifUrwVAq68eOd5oz3CDgs4PWwHgmBqlU5Wfd2lFJfoFykL3aFV
an64DOZJh3JxO2R63umNnTlAzZvQBCiE/KscTICOIu8nmtZow17YydQnmHIDJU+mUQIVU8nbB80S
8M1zpJ9yfCy/zy+LDa+W553cU0OkyReplg0Fc02Y0S2MEZkfBprwg9jAebbrTg+LO2lgZtFzZ16r
YambIJ8sNSW1F2p6KCGF5bjGfdRl3u1ffWfbZa5fiJCD317ANsfy7nAbcfUmP20n2C79IW1rglUp
IdwMiI9+neEKH05aiOlYKzh16y2bfJKP6GFP9Dchj6oeXtGouYslOIEVYsqPXIXoP+m7J/omyWG8
ptkLqQccwSe1UNPVEHNj30a2HjsHVDG8NHljUeI/22yGAE2NAOr8priiMsksBHOzoaZtMTc+Q73q
NM651O7ESkVyhaSncGM0WvIJsJ/E7AS+AihVXhTycg6szfm/CAkff1bc5UaSuUHSa6Wo9OL9TfTr
rL6XIYM6yNP0Qva7GsGIeT7F+qsycvi8dP1ZWEqVJj9IVGhCO1+31Mb1V//9mA2FqzKv2Jh2klYl
ZvvKzBynOskxdpoScrLuCLkgC/KWgqmfMsSqfTsphO5LNnyj54Li6o5iUFGPkCbTQE94yBo79G05
vBbLJ1Ns8tnPuyZ9I9+fDHpdMJGzBRaa5nHKv6PPiZxIUdOqbxMhHH7Vtxt8eIqcAAsLcIWfhnBp
6g0nGQWsdGKv6LwdhzbilRyTSunOt2ZrbnWwVJM1prbp55NgZcuGi7QLJfWICSI1KaxOoVuMlGcq
olt3O3HW7U6xf0qD2382PZOtNeG8Tr2NmGcczfaK4SWTppqqs3ARJSlL6knQ/o7yVLtI+QNtlhV7
/cU+j6ZNOPApWUv+VecffPCSAFGq4mYtvLGTqHKuFt7+CWvwMs4o6w5HOnjHdH+CCNtSaN/dh806
1I7qTIgE7rA0SHmwigoCxiZeWGZAqUy0Ajl/mWZo0+dDzPNSnA9DMsKjRpRKqLTQ1dnx3G9Or6uY
AQXAUsBKY/zwvmIBmvifyMjAM/jdJiC/MnIsNqJpr89crpSIEb8wSH36ng2T73ERn4gA8BRuRmpj
y+if2GAan8BujzvvM2EeSF5TqyQeo6qRGSErbOFhDJlU1EcxDXBDBvPrQfHJjgADW8lcme+aGA4A
PVrnVo0sPTtmsrhE642eNlDj3hEHAWPYUsv/acbKGVAke9A+HlZPnbK+uTu5Ej4biqwIKJQiFF4j
qUemG3NQkdIqX1tVPxeo1SyN+CzUIq+cKwNpGLckvOJSxQeFm1Z0hKJ+F0VCF/PnjuLPYKTtADMG
Zt9GuIoE4WWDC6gDss14u1pONO+rsl80SXHwaq0eme3d5WEKyUy1SR8dPk92kHsMf8oSMnpdOgpw
Am6PZWMVYtjKg91yyi8C/H6JdGd1GFcNliV/J3qT27m8jZnrXdJYibzZTDZynm+ucywNPPtWG9rL
bR411kW09NB70/g7CsDCcydQCi6lNZ937yXddB9hdFkfp+fAGRqXLaHm8Ymxl4CAwznPafqOPpre
0aKiUVC2BOSZFzinx2Sq/pt/jZ2uPdCNY5jGPoUIloD/wPjrV76NxjQ6DxVbAYTn+bWtyxmAAq7t
Xxnk6OrH7UNFDNBHzB43D9A5E/bLysOocfr3CnkWfBRHVYAaXZgFzq4IAAsW+96DQZD9Lb1dK0SI
u3xzTBnd64Yk3NA8ze/LoNx4yV/exvPTJqKuFdnRZYwR5vnvCzOruEEsiCp13lxIYJe33mj5BiYn
Pv1vmJ88fNqgm1UuKp2iQYF76ZkCcIVxgvy3XEnUpP4UeDhJC/a6Rc77mjJlHNiYmm0KUsYW97gr
im+Bpc9sJegN7MeqLp9acDHw5OUlRP51Q+q97RfQ32XzrY5kt7Tfqqe0nhPVu8WsFxYwVQpbpT55
8OtG3tx5lmJJr4I+vO8W0Ildb2yJDObGkdGLSSmyR+Fc9+arZDRwTuuPuGckLS4f5DWCbOWSepNe
Rt7lcpSNhpvwiXxCVcIJScoIDZlps0UXD/Gv95fkqJBvGqr8DAC5mDXKQX1PRnf2nLHkRcJorjXZ
zooNSmsVMY0C5qhb08pWLgeUbF9MbxJChEwqi7Kjqh/nQS3A63alhj+3cTNpmzrFvP4vf9pfibni
V7UskyERVu7HqHk0tngkynb2AjJqP7hU3n044HzQXqKWc1INamLuzjEX2tqBKoPttX5aPgvsaqbu
mULveWD9MZeNQpJVVT3zRVKG4ykPfIZB9kkPWzry0E+hn/aNRZYvdaP5wDbFfc9J+77MY9+hiwdS
3Ok6r84wjcOVyXWnqJ6Ifqo1I8gybwTQpga/BBvl7siXARzHqocxDKB0vRMG4wZQ2E1cUnBhN3Y7
/MEuCoJuEitPqRPLxPh+LL9REANrB1SLRWoAZdpUeEZ18cKZ667oF0wAktiegbsTzQ8fuXVlq8BS
fQhW3S7OM5kfNSKkKiy+GvwceZAkweEUww4bUuVBpsqfpFZWMluPu6Z+sz73AmW4s7ghoZJgnHVe
h5LY38d7PLrJdfjsg5n0mXeFN5dsE4luPIF5WBMJZTnc9bAGgk3yjUmIy34zjruadxoMvHbYUJWK
/VbUt/FCqvi8MOxzA7yX6mcs0uW2Uk1C1+K80eqTwkKJlsIV3cUYBNvXGOFuW79dO4VzfX4ocoPA
OxUfSTmFH4ybFFCJ9zcOmxeGrGmV44RdQCWFGZYdO6GtcXnbb8uZ827t1oIRb7QGOg2PYlz77ZjG
yUlCCIAS2Qxq0Bw47PFH12gIsCHIcqu8QYjdL248HvSLxb5U87DIaEttN9h4mc0V07G77NLLuP1H
ze9jmJRPyNVTmeB4wUcofvgfDyVngfbum5thvilxpaf7m7w7ap9lYNl9x8SDIOj09Y+VLzb/Y9c5
AbudRV5kuLFWWUKlFcei5KdctJW+L2UFiP4S/6yrqIz9am+Sf8gGVNyVQfEqyv6VlmitzoHjpEs0
0xShQdYd0nfmewW51UkpNz+24iCLl5p0wEzNeL+cPB/fyZz9l0e1i5AVCoJuMdD03gX1Wxukegoc
Hy+eizk1tFYs+eg0f6je3e6ZSdC7Kk0iu5pneqCrB5ljxNvHpxyhRY0f7vyohLJ77J021nkdBESz
SyjMqUOYnrqGERImQDHRpvZKMEKrME3M42Pn7Q/ZJ6IzdstwnmYueSvURH2/ywjT0k7BPUG1FRH3
bjvJXNiU9NjgNBZBytc2mSOLXV4xowE6Uys6xzOJ8/48aCECOmrWdVcjsz95D/wRsOP7RpppGhm+
dVhGFj7qnzWRYY6IjMP2dcnRNy023LWV9QxLtdiE0GhjFJSYMXrIjuNIW1fiBXlrNZPHAu8vim57
P/lJZDlx0AtSnAEldW/KT97Vcv9CXXPic/d4A3JJUbWJ+ytEG2ZWF26cwmDeznE55dqnfoc3diPN
4bE93ltAX+9wnF0jynKfATAyCGvR92GGSm4bHL/dGEE5Oi+Cbl9oupTJytvfurheVORB+w+KPomi
ZvvVrus44Qd6H/oz7SrQ8wTKuraVnHoquUyim+c4NLalqzfj/3iboujbhzMyvlABoux46+r0k0uk
ccfyZwu8z6GzlEXJW5bKhhV+9LtwkeVrZqRAYBv60V/89Whf1gReni+UhkgrHvIKku6HAF4aofCV
yraPjcCJL6vupvsNUmcWMDN8FF+8+E74MHKfzXPp5RpoyPwlCS0xXfnJL6kmDIrtN9iV6Vy3Nqo5
Y8gs5Mtd9X8CvD0nEq70sLUnJjoFI23iR7/DOmbYHUEL8stapEn7ZNgFAqoxkLxw6enlerw2RyCO
ziN2mqEbyETyDLVfEl09BD+SqvJLjMhW7hkBK/OsiNpqa1Mqx8XWbHxHbBHKGv/adyr6UexKqR/D
YDW3woMwU73F6ZLolqJYuI0GmP58vFFyQ9T2zpBOlog69GklEIpP1I+2KhFxBOOOFyllhmP4v8Jd
+ve7Ruskb8yXAcbhKCfP+9DMaTjfyjYIpzefQ4A9eC2x8lEEPShGT4fKmHiA5l43uNcnjHfxGMsP
h161gldVvHuu8liy+wtr0+hh/SgOUJBatlg9Bk03L30qw8VrMVPF/x4y+gSdVaSJnR/huo3CzDNs
XupOnd1ym2cvLpOtGxXEZcTMZCa4n/DN35qBImv6IQpnPHn3BvAMWNzLy3UzEfRY7x/W74DaSLsV
coY+hWQemozpWjMzyd5xcjVtj5X7Rt6IYFjl/gDeffvLDTqO2t6lJkpRYjbDaBBXdLj5r1hWiU+h
FiUEWJzShFahU4WzIKdbf5gNsen1auIy9gBeIt9Nw281NhJRfLaMtwxBLQkoNjrzuUsHji97N6gw
5Q3FPPC4HYL9uP9cNj6ICc5GQlU8kyNq4TLc08lVJmT9CnugtGqTRUBQIszjfIuGzqLvB8QrVaG1
ZGdwhHqDN69DoG5pPnJCrqR+BjrX8kr0+yq9mAkuLrrpe1vOLLU/Axslj4ekE7r4PqchXZAPlKVW
mvFA4ksUq9EjEA9RhCsOE7/6/CFT36mk8pTIWUf2m20xExgNY+SAj7uKLpxow4qvH2AGj55hlVxn
sEloacc6ThflxIaKJMKfAmAbzqn9BH7KaPJLniLntvItm4xypXPhxHMiX/6ZDonP9Ba+YVRvzxdx
tCe4p6sqQNdHcz05VDqjc7NmqgAroAnk9AwHPnmvU8lETHlWv06HjWz7vD0U4JaMSbLa+dptWhga
155ZLGSdwyvI67sTVvyVQktD4iO/+byf5qpQVchKOpxCHieI6t3Id5kAsLJ89JVIuRZEXaTtcVwQ
7AZhGeTuai0iUAPqpom3XkPCdVbExmFGyuIqQzSWLONw6d+rqMq1rNYqp5nnkQ6/LFvP8LywHK9v
Hh8BSMFq/paXdLsKXGUEGvP6A+IRPP4//wV/G0SU3wdXN5122sDgDcUFlklivZ5tNqrHGyN8llJR
nLZocbYHXsVaL20msFVigGWZjMtLGudDsn44UB4FeKR1Vsr/NjL45z6bqLGVH9A3avk4/OQDr/WM
8cDtlR+qklxDekiJlwmf9xmX4hV5nrUYmQZMjiVvZ5g7S0h4dsue5bqr0pAI2p/3YOktTtqruW5k
fLEwXuzFAkskiuJWOW8aQybhlpblt4KcTS3z1zE/MRwsgFp4JJrMnWfJpnoyXR/stsRC9IjHff56
GSOULIJPUHuXf6tTjPC+v+5TTsEU3y92GMCmQu3v+w1qVdwu9bBLFqu/bo3vTykgfbq6uyXwYnhA
gLAS+i52udVdjy6ZR/lGlneEZcuKprgSxFTe+BLfo6FOogRmqAGUhwBUkmdzgriIHbtyz4cHtOUv
Q4YidfnnOdQ7yj0banvHmRsZ2/oK7G9L5W56Z3r7Iio79M4XsMdZxkqjVpNo+bVKj08qHv0g7ZGw
wdGzG4RPTSjsZwrYqR4iDxu+EUcYinfAd1t+WJlKSqoSBaTDONKcWVgCTc3oH89606tDdTzUufro
zimQwqsFXm5Y/tT+kZR1cGeBDs8jP2ETw2/2pR+kT6856gDW6+Uctsl0PgtGN819ufCzH82z5ySu
hQrU/H8k0IpkUyuBkTyerqoHEzHkOF1x+aSguQk+AiaoMxYHkn0Yd3LSvAMMxGi/ytUixZK/c++w
6waa/BvTf7UlUzUbJS4+6PrwwpLwOxYcJShr7qL6DTyk0IgYs35K9APqgUMW7YN0w+0ezYSaZi9X
Ixi3cHmZyYuzCOKrNLS2WEbVsnNhJpi2h/eH1FqWLfyGxExek2lqx5Iwto3m+vIjdeOwLC27hJor
wfdG2kuNG/ImafQmDNw/ATP5tx+Nnl/WfXMvCJ1S8PcMZU54uWDiQN6G4X9HPfQobtiXngM5MhMz
SweaiNAsKwlz2hzL+WQTqJQstiy26HsaLKASu9AXk7EQ1GeB2XcQHVY7GuLRSp4+HqGbxhfSY7v3
NzBbpt5m2zVSHBx6yU1Z5j2uNgs3x6ea0GIQ110ovyLR3piFT+Ni9RHCjQCKs5Z9Gj/caLQjEoIU
TsMwP19UQKloTMcRrpmiGlLr2weu8IZ6Ajz92yIgreUkvjtGlmC4Un+qBuLKVrYRgMxDlIBIVkbW
mRlIXOdW6vIvyzPtz8u1LCg5zk9ku7XLX5FvwGbcjmKbFYXtzzoqVlyh6K7N/U+XQVPt1nk6nDQr
n5kdtoal914K79CWNZO3qHm91tQqj6zELmAeasOVnHaAHX9C8zW8Oe8q3uYtjU3IHEUcF1GkRO5d
rRgQABCA3w8gmZkZsJptlrslrF6sMZcvUojGykPyguvc+RmB4rG5cWyiqfdkkHT3AeazKhmvUqc6
JP18oQF3ywDFxJm54OGFklqOKA/S8EJ5bcAZS9btrjpcZzt18WYB/6U40h+egwMdrc5NckYcX/RO
kuGWjKxg6ecZugwSTgr6M68eAKxpX6dN2nDh4NWpH5sRAShQhqBUpv1GiDy0YcKpHMlt9qMJL2q9
Zi8PZsCOhaGt5v2aipY/E3CHMlyEAoYDoAZqcQdj924LzTLL8K8DPSYjxXAN8Uh2bTtuXCEUH8kN
RqPjJCnp9AxAKVz7EB4ExgAkeyTatmtXBnpRZhx4KY1gaPGoFP8hWbTRAeMJpWXHhiJXPFVGxFnT
thYq1Ut8Ff9s8nx+IezW66LFO+IYMqBMKeosN/FMH/IY1usvovioibyVUYdOYBLFva+4E5jI8rVU
3MwbIZ8n1EzPyM2fCqBb8FbRXgw53DNEnlcYCfGL9ah5Dtz6v9WJk4Um2qsM3BbgvD5oKL77SI95
rPVNWVMY6dGU6Ot6WYew5tqmLwMtWOpiaoJfQi4x1FLZpd33dd54RSBex3vYBIOjAlDP+2XevSNc
Rb9cQ6LQgPq1ec575CoXt4Y15XsTF3qELPEQ8YITHISZy87x3pXKDS/djG9eAgd1bueNRJuB4c/H
oXgSnim8kGXSFIuxwgLfKHWfSmyRds0dV8S/UYd1H49ylC71STwUBajGtDWpY2DTo6DjtpkhBFNs
W9bRRxeSJ1CrM/k54Rw9UEB3w1fth1/6K2ysOOZfVZ4JHzQkZMJf5p3e0Ul/f7qvxPmxRr2f/4se
taAZFjBHzm6QDwq3mvB+CfZF+nm8JRw61PfchJ2YNND0hnNbKSQ/fKaZU90mzHh7ZEPIOBlzxyHw
mW9myg0dYXFWRR0fLQAaBvjLuro9ebtWT+hmhClOz2aRnkuG94OG9ZMjK/9IZwbYWyMOlNThOPJK
d9UB3w3Jd792sNTi9JHrviQ5I3CWkAvJ2cq+36kDyPBt6LDxX0E46Mor3i24GB6mPiVdygV+gce7
EdmS5iTdfP60BNzrxkD8n6hMLWhSmSUcJVDoOdbh+sZdvshe+nkl8HdSOi7lWG3Dm/tojdFnDQsF
3jfJhD8r0CNn8TV775wU3OL/coN4PdmJiWT++56Te2ty1Kd1xQ5J8vMGL5zLz0Rk47nbFMg+csvC
09GpQGKjVXGL0roYJ8nfdM60Rx/kW6TlEIGCXhvjS7l3gXEMwjTiWCIGC4IfRNhur4RLXMgXtJiP
LatSJGZzThbwouMVYUJcDAlF3C0FQAmE1gXUaOtG2WLzp+Bw9zBpCmRMQB+zKOB8PD9XdLUNkdG7
ZFdmiSfuI1WucZGb9clUOYk5V951D97a7GNWCX8xVEd4CRcHANRz05Uc17T9qvX3WORjA+P0ENax
si0NoyY06psIV7Dvnh0IGEUWklE38Gja+kOCsyfPBOJlEpIdGrzrtC+MZYScuEBV3g+nhleI98Ov
t5BymhISON8DVFUWgP4bqUJvbsAbCHSeh/qte+H+HBuz0ZtUP7bTXrwPCg8ZtPPCoUKssDBVjn9X
ISGKRkmPDOdOTECVGo8C0tg/Dt9+FZXKoRZPtwgv6aSQRSVyDRkZYeedUAYvAFcElhh+igDz3/Kf
5qxaMJWAmfF0wqvRwjJBI23Su+mdvPjb4pvAwlNpSqrbi6DO6FBW5G+qRNAYERUgfamVEdo3pDIl
fobaTwlX7OWn+Hzp/Ebzv7C9mwv+lPT3LBJwQhoQU9ee8WfDNwb7U8mjineQiG/REGAyj6Q8p1dE
TJyLeICKCiXTNAja8DH2evrnzH0YakEssd6ITWjMbV96OW9LLit8dxjiOrXog6MQ5j2jbq2ACKFw
AzFpx8wF2dOHgq+pwLLjDgS+hckxMzlrcKVdcEiU1CGYuY1Hqp4swL3c7fOjJreG8604ixa6C/7H
AlPx3Hdx+XA55UI1Td1FuJ1jmd0XaAe3Ax0du3jUvwEj8ec84k+z1gbbLl61vj/OwY4ZYi5oySF/
uEyvjTLP1so7i9uvDD1bs+D56PgCa16kIXfCi/bc2Z64K3/AB6pXrC3kFUyaCA0OdNuPMRas0ix/
94XuhTN4/CC2elSeCqsxV7f2ndJt3sm66Iz3+Aqfj1nbaaNhLNPQQn4zOjYo95Qf997tojTVd7tz
d6Tw3rzkpTXb0ZLRTR8TmpSH1swiLMgapj2xPK4+KW0regNx739HB/vnvV9bTCQsqfETZ7C0FJXk
RbyGPrcNXeGaq5l6mCuk2/bdzczehuTHSQf2lJ1YEGAb4/cZDN1nLNIsFR/0BbcQUwZxMB12AHJN
S8IZPYGwZ+m6nadaDTIQEvJRSn+i/H+NwrbYOJwUZv86uiBd+oWWjeE5nN8STnUgsa1TVw9UrW35
ACQ85PkIQVpPkZF8UJgWH8iIsHUrnCvfW3JGrYE9tWbd+oHprd8aSmVSq48Z5JPlMR196UpCEXQ+
bMHBgvJvdIlUyQU7O81GjzLlQ/xnSa1I0zoqMB5tu/SNuf+qX3lIXXvCoSL93EWlYwsVASvXq3Co
GSL/2VoeY5+fm/cofaYrLmzRubl54fLfJYc3wd8u3/pYJubxDGDqrN181bMUuh+BYO75DdYwn+JX
syq+EHxlr24NeE0uYF4upFoXv1t/2S4ZwPleP03AS1PRPT3bGJ2dkuxMKFQsyFvlT421MIGUWJXy
1c1Pg+surn3+T+rqLVgmE4FhRlWcUGPrt9FY5Vs9V3bI9bYs5p9a2PB0Ro7lmZalp1l9xaQe2FZ7
SRTpbKUu4ZVTcQNsRDL1K4jerbVWt98zxW8h/NI+k+tJ33CrKNecCcvvCwHJeGwPqwaXqahhIaG0
3wR4mJBdIsNmCmMAK6HTfkEhW6tTylLcBh1beFceTVJ93JV0bsYJTWEugS4MX4U9ctHKL8dmNyMJ
JqJ6xHzAuE9e15LIN5OX3rIenHbpXjjK8E40WIQC84OxP5EktpZTxlD1cyNZ6qIdHRAJTrJNj5+R
w+FdRxexJacWzdacJeYBAXuvmsm7lf17uI8KjqdO+aBO6V9BRjvCGmAZd0XIy94YW6ZK2aS6Q6lD
VB++YCSuwf48mSwGodWen65CDOPyuaVPu8UBBDdtS29VXGS9/doqjMDZ+f0rudzEEGfSeKck7QBX
tjUZNoxMO20qwH9F63JhqwfkWSYUNpTz9j2CoLTAXAWmo4jhlctfNunrYyPaB2Lgiebfp/WR50Px
qv+xwySQuAii0vnxsoWw6lWuzkHr7byO8V0layLuzRB8rWPld9sfT2phZ+YYZB+9j64meDaJwZhx
6DfJhLh5tgweBeMzV0MLkhiJutITl68QVMMawC2uLGNxRh+dNSfKyoQVQuueRxFFiYrA50v/uZx/
7/G4qAiyp7OsOLgq7IyfALMpn/BXrOdBopvJRR0DE49rwvevnbwkLNy7ZJiSl6Jg5ThQORaU0amf
EzJIoBiIeGtFMfjbcwfa40Y9MVMHN3eVSt2wMJQJ1hGJAtSIeHAWn4uT9gGugrhdUIDCJ3bhUtmv
SRWRU15UEfwP5YghYbPLhgfBiI9sCTDBvIkJBd7agAqsTq0DECag3gLLcXUypZbr7MtqfSZP1RrD
t3IBNzKsWS/W8y0V6/IQM9uv3MJV09pk5Zj0b3+AoMupbeslYs9XpW2joR59U8fjEWx+t7aquuOB
uv+zI+FqD71q83PqXanwjSUxs5dvXFJFm6fmeJBQMFRAWXlSvGLIMIP/tToNOHaYxmGw9kejVQHj
xCqK+18cWShm9nTeDR/Gjleg0JfFPdSLfOGVYVW6ySDkqf+pq00sokrEmcby8dnOKa1uAQzVWed9
w03+e8mLXfVIoztZLTYmDgow9buUDVdz57IWjATxl9Y/0M0gdXf8zO94BkU+KrO6jxtJgRo8N7YE
KpETt4hVO9Id7TzNH32DKAKKRBaOKipcrimANEo6endSRXaRCXcfN5QdCZPwPGKEJnn1YkU82JKL
ZbmUL+Ed8faFeG9jzKzcEKheBCYPVva3tbMbu7Ad8Cz6cuVe4kw7Vji6oXolyekHvNGuUA01leRD
yNrl7OPzFuUbwE1gBNkztS8UyWt4Lg7hWuEeOwrff+j2Dwn/dOTAMZjLzblibZIPnX6rniPQKGxA
fbtqSD9YDsDoNra2RK8ri7zj8BlSXR3wciXFf9XNRuD9wZ7y4YlLwvKYkwMSeCphwsAgAj9zFQmZ
QZvQyIJt5ces+UFgBaGk81WLR3nH5MP9zGN8IEJ1w+mVKUSF3TayRsIzs3K1SfVqIRLIfqsFWENm
bs5wWHKT3KRyOgtZhBWRL/L+ZIKafIBVqe6F/bk5QRXEuAeHLG0dOiKU5s4szlBSdhryrchykGqL
jxV/r15T3j9FcVki5ueILd0LfZKx2nqzqBw55b11DHfKAzaRQkLdMRWGRPgepS1yLfEJzNlTv2oX
2ZkxBppKTskfcyGFk2KEP+38itrFGolhGGpluUOUESlbyHcpcSxKwbligwXCLgsoSOBQyZXU6g8+
bdssBEvpnx2/XoIKmNT/UVlipaY1tjGAsM1UYu8/OUZbhsoEF+4eTmbU30MqaDHetlw6h4HeA1Uh
bIAO9EW2gmtANBHkHR5PTE4ejrRa9qgU0ggNuOKCys41Dflf1YuKwGJ6NZ8gxNHWOi1x24xdWeYw
hwDDBUt038F0XazdMnlm90dSJri+EU0DXqWUg7VgTbBwdVBUUjcJMBIdBCuhfjq1m1zdFFo6ckBW
iADJSIrKwJzFkKYJ97K9e9WZNa2acsvhxE3GQzkPdWpCL1pVshYoIZGQY3Y5yJOxgRqN+OGfJZGa
Vo+sYf7LPlrfsWMU9dgo8z/oev2ivqfzkk+969FtYtrv76GizTLMSSjJW0CQTjXgGAplS2+j4np3
tUz+Cv6WeHJ+TOEIdfmuafGEhcmbYcVinu6DwcUsf69GN/0PrScUGMOCLZ+fcR5GSedC0FzJMthW
SZ4crlijrqQC0una6MZL8d/jOLX3GMOb8L1pqBwn4jUaJhWSzFTwTBRVgaCw3DcptEpcaghmANKd
cpqy9GGPePhrKIJopqaeJ9GZrEUUg9a5xGZ+SVP+HIzge6jNnGyMbd3uQKNPnOBcLUCuM+T/lQ3W
5u/fWovXpW7kgTucEkrVZUHXfTajTIwaAkwBvPR4km4IW5891WQCNAJdajm7ofFKmB+kAeo2YYja
A3Y11VMv4MnTiUnUqbdE1YZr5owq9XwdnbEwYoJNHBlK+M0HqWlv5PCkAETRpQiOD7cG4xBtYwt8
3zWcfJ3u9g+CJTm69v8fD03NwBjdURZYFV9hx/5fRhWSioskZSrZ4oHm9ldw2lPwvNDDNK77Lwpk
3bPZQDDBqXnHt9ZiM3ebCJan4cl7lKPqVXLoteEGBbkzNdmzAHnHcmeioi5xnLDe2CAidCcJ97x5
5Xvw/ANqE6/9fGp8MJIRRCgaXSWAYtQA/XTTbDWfC9rT/4IoBjkTAzqFRf0lqslSQRalooPMUY33
KpD/cYZZ1cjGJ5QE3kgnoDiHhqeU9ffDF0mYNETGP1baCLF+DhYMngWMQoppoTmsd6NboNz7G3dN
1JwcaCtFkt9Tx6dUHOKKJ+0Gg9Ks09AWj/Lb5e039rfUGXRAcnEtN+OelOVVJQN7gCbqDXc0Ccul
E5ggzAa8p233v2P0K6zPE5mlIr3DaGzUeALtFMlv8dPxbp3oKmxpL53cDNrMjcibwcGQ1BrhpqG5
UEIeFwyMRzPoF1JYiq63R4DPlEV0B9ZvRCGwQ/RbrwugNof8r0Ndpp3gLAbRyyr4ILnnywMxE9aM
JF4g36lYh2eG1yblIpVFunRR1TaJv0v5B++enkck6SHhLn9lVwdKL1BcdkqJi51UwwWxSv71guif
UDaFLcji7FQmjGTkaOyOtw6ccQaqPOzHhidEkL1yKdVxie6eQj++rMwop8K0G+ovZhiBqRQ7z7wK
Q2SuDRGhQDi6X/cFH1eRwZ+8clT9agF7/ebLzwU/kpKgm/PaTzbVvrHSiVEP4mxOTn8rPn8v7am+
U8wRsAf7FidBsAKFvOMyLRa5BxW8xYkmkR9LSxZwIT0AvzFNcb/xhwjmRF52WaGJJVYV+Xdnxvb3
O//hXS1nxZMv0JOKobm8G677s5qfaxv9m8bVndtHW/YfxTbJcG4+5oX/m5rRvYhTFWqCQKs1ABwb
kj2ubO7IPxUPxY+SBkq1BfGT7mARrxRrzqx33rthpE1HNIMDr4fmtQJNrkzf21KyJMNaEt3D81hP
FhyVRcqkxFe1JKlDzMz9uzkyxIPexTnOUjuizK8CnFTDKfXS60Mv27ik/1hOv1KOtxa9dSdKAVsl
3KmlKPvM3ThsBWSGc13bcYMfg23t/F0a+GHGfRJnvO6ASEKaixnCYu0g1fwH/g3ilrALU71xK001
kRtniwM2FwJKRkT3pryguSwh9lYWcnReyoq4G2tCTtQWHXvqv96MWs/rZm7GcFvCNhcHPAjbT9iN
i4o8gr6po4LuEp3XVBDoOncCvPlv2RjUdDpYTDORze2i1ov0no5Rd3dYN+HfsJ9lL36Ia6PTA5S8
SwgCVDiom+iVTK1Ft7fqvDlzCTKuNSA9WV0OLakZ0yiQrk5rk+nk4jWaaKP/mvEvtRJ/iqc84UQM
c2lKfLsViqF3V8eE8VKGwyQg46Ky6hsOk/KRgMb07Qu3OsaC2OuVbz/PDVSPpk+AdsPVo6XBkCh5
Ob+wQsxMiy2ZeuIySYkoHFjhd1eWhmehpgvEWn//yAisyn0lShlhaakETLURun8hdL0p3+B2tTxz
NlSKl8hIZC/n3wvjTjj+AKZZ3IPNZ3rmUY0JLxEjnfzjrxLAwxrB4Rc4DEJhY5O3HbYOtOZfsaUK
nX7WAxtAeFxYeqMbnoRu/sw0KkgU74Eqi9i8bCVhTF6hwP/whKBNm1xGnJQi0MyAdlyRBZgMvAlH
WTHKKOqift1kwrHuWvGIcpIglQXCD526k9JPtPQMK//0Jcug7SP0flGaUQZLyufLmrChZURYzbIo
3IKSEFAx8tr4RB/6lPCwuazW42SRycnWCCpI1iLq3DINJ4Ajs4MV7hXuh08I237Yyd1TmgvFQD6s
UG/eoDtJ4fq25SpJ5qn/7UdypoxiHw2P0VkY0nkRjwn2zjrq26/4zuMWWg6OqyjzYT4H1R9nzQQL
7Yx2wlf4yN5kBfOstEx0Wx+tNHN94Mqe1TAQtkNQPZZFreu0oDp8kifdgyUe/ZhYaGFJuoliNoiG
FVojtL+e/OkjzoWR7dVnRTtFLKrcYY4EwRXdFJF4/nWeg5cRGBDBojV4Ma2EbCwI5ChQM/ZPd7ZZ
VPkzS6H6NKfROx0xBQJi1f6gLBFhlKdJ0Z2wNZAZ9nSefh+HRPoHzlg0twOiWpK09pNM4JS3qUOA
9+MppKIhDPqeyezWwGhWXlOZSfO3wXZqIdHUUu6SA0ken5l97ZrV9qJLbqKGCwlbMYEBjFu+M65G
F3fqhMPZBBhTlFlrWK2bifvu4kGGkeVOR/+NXrvrXPktdQxWQKb+MbFvrBqybAQaVEdKLiU3IcPY
DKkxktNDQUyGM/VsUHJpFmdvKscrbBf5wg6Yj5fZh+P+txHMiAY9LkeckNHvtZmlT5G8jHbziI/D
AAS6H9N0S4A/ns+CNGS8I5VkO4bFSeuSgEY1dGDk7EgINUVJRSCK7BbkESu3Ct8ikHnCIp/kT6fB
RiVMehp+oAym18Tx5woWFC1TQU/Ce6x6Rt4N8c0DutIynFgBZYjFr/P/a/KLxs2dbubIG03IStiY
QkPUsHKJS3y6qbD/4cJIN5UjzrDdXnWfFqGaPv4rfcTITXpUnGBpvMCTdzudapbRtfHq9++vRlEh
7r03mWqNQyMeKK2eNjQ3vSC8/7GNp0kF4st7H6FrtMUnA+fZl+e4TNJzAdNtojJoa8nhlSkvcCDP
4eX1dxxR4Syv8TIhZuUKn6lKx3uYmpp52FO13rEaTUS9omrF2ZguGaw6PJIb5Xvqz3ZXB1HIcDDw
t+jWVkQ5c3tOZtjENQywiKAX/XZ1dsSC9NvuXCD2wPB6apCti8Y7mUFDwRCskXx2yETN+DNxrZUU
qHr1y+xHMGm69LJfHyluTmEA5JpQDIwM+mr3t4m9Ax7eJbLkYhDAllXXTVt2jK3UyVCRH8Z/byvk
fAqGRtU+k9PXdkhwKKcErlIKnxSF+7D/0OCBUu60dEXuum0N/HiqKvv9sGkDImovXO1nxHch02RM
V9AmqmGav12h9zKzLkGstNMgzP4S/1lIH9W+o45WtXMmjt+M4iLW42mZRs4tgv2aeE7DB//h51hJ
pGtWBG3cWw6xk1QBUKyjH3+bHT/aOX0EbYzK8obp9aGvFDoLXBK4AtTpmuMLVPmQCv74i4Lbs4oR
oYSPWIGn8sKomqR1NJk4MZIjSMacb7fHjDsGbPYrlZB6B4A7hOrodiaZQ/r6mGoBqMtEqNq89KKh
zw+5nk47efLIc4nSShlpRT4oPRbCXfq5+RMHe0W3gSP7/dAGK528TcUvr8ksNfhJbXWXJxsp9xvF
gyoilacb5+oidiF6LJXmQGnsl0MUqq9O9la1hmLthGw/5AgZH7BOwlUUaLt6O1nxN/GffvqpR9oK
uboe8r92Eqawg4uz4lVv/y3mxQDW54xR+eCmFBOQjdnJ6tYyQ9T+37kvViK1Ep/1h6MV7pu9yuBv
3xXoO5UUWrP/EhI9ZZKs3wuq7K7HY3NzdIodlehsMVP4nBuQ+0EJGK2MVa3Xdnbkilat3hWGecmM
/fG+T3FQbCd6FP+G+zZuEFsLISHtY+wyLW90NWD+YXGsrEeyioU6xPARib1YqP3fkKa90KuGcLf9
GXPNnCkKvEVOzhgv+UJ7Vn+HgfwbVoH5x+VfWFs8FnDSiz4hlmhRTMWEZB1JFau7Hw0hEwJW49Bj
ztjkyTuPZ2/vPfHZUNMNz6NcWmRmbsTiGruTPSbLO/qZusJKQ1a81QAQ7Xt8se1B9+fva4KP95CA
jWSNHlUvXPxhyHtLxsXSTNZ2uilTj2Y+TfHRuYqFhlLl8nVOZ1W3J1gBxKjzhefak4yPvkzfzort
1Tj4CTmjsKDVBUuGDV70yp558aR6f6dhUlpCjsFqXobWE0ThxOuX/g5BfkLKc1KBFYCgYSFZ/ROE
iczyJPoULo9+M5wfExuUyONFlf1O/BC7xqDcz7pAPZ4yWhRJ26jEBpF320mkXtfqBFn7nefhtpsz
ETydn55WVuJILtKNaxUzy03f7lM5pNe+K2R0A37z1xIToeOW0s1QS+12KUfw51qRVvvDhwAfDbk/
NUc6g/Nfta36pCR5D5ePf2IEkOmkWdP56AKiVMrthb2vtgw99Ac5pr4961idFjYGSExghZg5VrG5
IEzC1mHyMi+HCvLsxjwVoWFEmz594anTBnQFZHC2FWK+AZVs6x+CedtqC0OGl7DMyElb1L+96mXx
/3Bug5wNjfbUzsaWXyMsKoZNIA3oKSmdMZqoiWKa5rpm+6yFJeafYLKtxPy4oiQ8vje3GcssXeQX
BEIwzKKTmgqMbCHMf5vVyxpv6x19TtJUf+D79RLiX8sBhl4iije2Gab5kJFWsmlkUP2L+Hije8iG
kwxYUIreV08cgrOf2y37LCivbEwg42LDC8rk6RIZtaNV1url+LYL+gyIjkOQPYHMoQSQwRDpIYPz
/fbDC1IG+vIxQJQITnRqSLFOEPOIW5GXxzenIu0gnd51vIHuD42S7nzjm3cnFIF0dfTqIwTotIvs
WUPkh7YqlDhScwQ7lHnmqGDOIy8beU0ZQUcNn7bavLtJ6+ijem0lqmi9ODXF1WMZma4qfFU2+RSB
QYUcJkgaYgJJXBTqTaUluHRYqe8qyJu6bEg13rDrj5cF2jzk1+fvo+MtQeJkZHTkk/V9F2Cvj4ED
GCe1Rt6x2pGSXRN09ZIzruVDF08FZFIl7mwrk4fzJ/Ux8OeXh+rPVgWPG3u4Idj1NDFJ1xR4Ipup
4QWpbwdNAnDncDsWx2uELN9BLsJh0NdEs7IPGeZKLcQ2vU4eGFw34jwWJHOO1xE/6S5JI3qUbQcv
l68HJk675TjyyqBqE36KUto7pfKXY+JlSrD5D0b5XxDnOaAME+3NLeYfoWbs65H0jYywz7KtYR4u
xPlqkjauToysW5C5WV3kHyw9a53pHv/IIPnNuEUtooYkSlrvqlP4K/gMigfpy52IPpJbzW7sf0xx
Xq4tZ44oYR77oT1WIQkXahBiAbBkaztlo1oKH4iDpIUTzFW4ojKxINljgLTFsXFk7oyKk+sBYE/9
0xb49VU2Vpg5WYlAJHoz09qTeSTnVJc2T679PEQopsbedE3w1c9y3X9uklG6h22EqbA9SeJ0zPdE
XSZOSypiwFITeeToUrV3YCQ04EpKCSM38KKf1a/hgHsitofAaIo8CnbGdzmVNe03BvW1nwIdmV/9
ODdEf0Yco3I42nJ3z6i/8rDmqArbQ35syp8ul6K/W+HjOJnw4jujNrNNMOobcVfM+Z61Puj3pk56
asQhT8KAk4sy/M4dKOtl0E2UMsAvMaz4PwVZJHxbtnH4RfknmGUPIangs4Py5FqVXk5nMMxcpopZ
SjVld0EMJCIxzkG0ztIWAJohZAaQCDsYa+ecaz9Fm0i/etlq7K0eAyFn+kNfnMZ7bVAlDWYdhbcd
hpSjP6QFzPsB8AExQfF/kC2XTleh7A8LbYJC92L+10SrzAdxeWcMbrTdR5a9H20Xmt1mdBg+cSQv
YouvnTfaJdpLoSlwYIyRGY+LGndeiM2zddIGKLDXNwvDDql7DqhIBJX6NBlfHE2Lyuie2cCW0ybW
Y/S0jkrKTbq+bhgYCs+N9I66Naj8GwgkI05BvGjvlfGzhJrI2KhrMclyUp+7Oyp5ZzFVEDHEt6E/
odrhgE2TX5Fwv2JgVPa528t4bKnkx9UNXmWFaXZMAVgsDNqT5ZX9XmoFQJ/ISe+j3EzRKviXOOzg
iLVIMI+iuwEGkJuZKOCLKuK4ovLCZuRzCqsNvgYq6Hd/irhsmDiIaInm9g71AsvmuAnT98zxSK3q
4hFOL8z4PDq9u0XYkAAmH2jyH5zNUc/juAazE9ehsL/HpUuEeIY9Ger1iALnLRmorPXSikaz5p6W
ijnhpW7cokfiQzsRCQ9z5YgY0OGVwNg2aNGKK7/IGgbAYC6EVlCVJszPmL+fB9XOar9zveosE5eX
V9x9S4s3RksCc5Z52niziLwi3/l7sDyBCVdYzeC/OYSxiwSogkhckT0C7lZg/pJ1jvtW4o+XIs65
E4zaXxrX7e+VnwMCr8Q+DdSpCCG0mWvnFn83FVXKTXxHY37PrsfZVfJ+IKjyVEgEinXclGWeRNiL
Lm2Bg20GsdeLSffYG0zlquP4eHOczggtRoGrMFRZqgU7Ig1ile4nm2X0KWsQRvDhltM+1WSLxx6t
oIAZIyhwPrv9TV5suhAhRFe7mGnYpT3tdkx8vytGpejdLmYp1XL+0K8V9FxIajNCdNAy3ozm4wEG
xvsS8cB9O+YZTudxtTCUcRPij6LJcyVukWfQPCBF3KSLrfA96wLqZf5J80YcXyQ6EOutM4FIOxhq
u0B5N1Eat8INJj7ocSyhKW+c651dXllE+4Vj9wIOx04hgL+haPUaixTk9Pq1GYeHMf+sr0zjm9ud
e7T+s1MBMp14vwuElSzcliHMjXeJNsQHoxWrshTHR4+jJq19WVYn2OVUB0EbRxs8xr5TkinMG2xQ
cT++PFdwVi7xhcuChD1Sma02YViOR6FLWTo0f+W+Y4In3hHyuVujgGLcgWp4cdpkdE5/9N8x3+DM
NFwxGFViyg0Q3QqJmaVzGwjfkr7slJxf2AC4L4st9KhikTnt19KZvS+x2kfI+Ynzuioazt8BSgSW
tevA/+BwTp42can5iLAYJkK9lgHjMaFpjXZ0b/e48dr14qZtO3AJFSjtJa9TQk40qBAhgwi/TROy
UYk4NMYfxA3xMeb/jLyfszeJrX2qntWa+R31w3l98M+3CB2aHTBlqqyNvTxVvub45+bBx90ueygW
BrUCrC+MBLRdEUoqwD9VHTMXVSv+7wXXlxV1YBWmolc+XO7/ZDKcA++A4whWA5BdlP98oWA5Vne2
IUc48h77zdT6EJeL+Z+zxNVuorXI8Y1po9xn1rgTLA8rtAsLWONynPd7k3IybhvCaodma4ww956M
ymZkQyHyOBLkb38HuG0VtaU82vzZEb+R3sg18N1c+PR21WfTwCHFhX3++lVRwzWI/KYyoPa/wUP2
3x4hLkOWBIVI2H5KsBfFsfdNonSuo7MLoNWpv3IhWSOiOe3s+ZA4z24NBXsi2zs8JJkJs0cWuiuZ
Fusw4xqrZl42Vmh0w7B8emy2zRqCRoRCtqE+d7Ui2zIZfsWfTdPaxaSA16xuYj0pjMw7c/HvLf1+
55ejogO0JYlURwFsmTrCPr7nHKEy8K6giaKClYMqA4uIGXUyrW2wwBdrSgHY6BCnwJMqCe+Met2Z
jCAyK+ukneewH3nyv5rmdgNla1IId59UqohYXTlIhH+xOjNHoiiOrKMW85PRda/MhkUCvPH6Wxc3
eZT4iXKx7w0vOPcoXvfgyFM+EAtLnOEnw0HElzkclQgMHaizmDiCg2eSccZ3H12vBkt7wXE0JNF1
vuCTMML5kPOOIJ4sSxGSAYRNP+qEImisDfGsgRlAllSsA2OOH1sRN5RhKS/NHOlTZhGG/GfqRas4
+CTt23tWhkYm03mpaKZzd2bB7C0TmM6E8X3jZVe0PeV+JX5UkAu6inqHhOPVIGsfr3WR/98Up/pa
ScoumMQ3RxHIh8AEzSy5FpDw48UsSsrV9/JlyALxn8dtMbMSkmC8zkzg4m1/g8eSrHMtljP5/TeB
+dP+rDpvuu77b68h7f7KMgajLj0QqZ6NnuwcqiQhLw8pYpFChyeQaEC1/sR6AGpqQK6oHoXt8Vm6
vvSE89FyvKvVuaOJMpKyp2BPyF7yfxb5e8+vmuuCuaqx7siSlLX2/jR7ihVgdxMs0coM1iWxh5fQ
9BlNmZ/1qTIdzHx3Npl7d65jZ8lMm0NrjNdkfuqdH4Fi4LugKGvJ/Q91FcnYgrihWSAeJ+vjHL2g
nCd67mAAHHtNxGlkg1I74Q8pstpyG9Jn9B8Wgi0qLgzQHSaOdMxS9+PVy415t3wh3e88li9d5NWK
2utPn2BDRwApn7UsHi7SC47F8Y68ZXQSVjQQfdLeHtzAGZmvPdQ/gLGJ/ThvoUe2jBfhuX8D1PXH
WtWxCMh0/5NT/x4vWISIpbva+5GXmxeDXNjRXuBURiUEmDX66fZ/0WUGKVsjCpScp+21RJ4DqKW7
2Vo53N1KWZDl8P/ZEl4vXqgMCoGZh1dYOCviEhw15rkQ5vXDJmjmzwpB7i1iGdke4hYudKY1x72X
r1YL1gqTBWQJ9QxyYnnAP2o/OhSSw9+Uf0x9V4wZMpcIIDIICdP/tqhS7vwVpvxzNL/m6wgeUcd7
4nKapA10jpMWGRiLisuFQMb2VwnwRaqaohBVbqfkhcLD1N2DfvhLcqDFIpQjvYbov2pJgKT9NJU7
L4HvbqOBqYNsn9psMPC7v16yhtSIN0KLMCouN5M8sQwoZtzvizfrdpehD0Fie0uP1z+LlsPZaFWV
zu6TzckwxLlHkmH+s6H59aHAZJcaRfY2xnRfwycaAC1YzTeWwgXZv1OGCC29aRbgkfg39SD9qb08
VH4EUY2H1M+wSmpsxY15cyIBTWXgCYG5lVeFPPKoz72ZYg0PYUCGBBk8v/NCm8wCyxFxbdjs0L3w
1cnYyH+93Q6wepwlsgy2/B3vAfZuXt4N3s6jDcbMMiQ2s01T+qMA4bwxQhHNOKk8w8u7rWTfxkiD
5pZGkOaWz6h0XMzWndCxZHfWmiF2FniVt97ygyekBZf9DDdSdCuWNRDg9GY8fxy3Z9kxZEIPbIRn
Ev9Juc40e7zPbsgGjeFxnxdv61FcowXc7izzE+oyckJPGm+/utlaTKOuoIlTinoAscKBL4ba5ywY
eGYrP2g0Fdbs9IjtW47ECiK2OM+38pJsnR5gBgjert1bSEiofYUSPOpLEOy7ijcBqmX/8b1GyQfH
YxzRGuCPr7yhK8Cbl6tN0lRpWaV9nws0d36s3eVQY3gXLj2ArSRhz9LBiZoKb0KYparJtID1vB1f
gwWR1EjzSbik1kucaqTSFryy8L3oPFUBqS1CDquJOR7dIHqr5CuXjKG+JxAgwD5fyFe80GOOsPdN
lfikt6u+pEDOKUYIA82twCR09TvVKfE+UNgJVm7gwtSnAPNMQ3vQJLKF2PLm35H4PYUlw8HTvKf5
eESrF2v76rUTWDSRSveg7dYZ6a1ULk8p/JmJy5YZylyiRWAuGT/aCHCell7SOpcYoJhlHgCN7UCs
RNTHmLkZTzpMWZIlId2vZa/cmqznYBqxmRGAypl5FVxRiCSqGFrSzVKgBefUihDJvLQvJNBSyv+N
P57mdWovTSOy+/NoEWn5FFf+RGedwZscV29Akq6TtPLUK+4TP5eiVcxYQbFXUGR7QtvicvmENs0L
d1jPd/7A6lC6Ww6iq/FfWUQKSR5fSUzXmE4+NFfoftQ+kUxe1ZZHtxrtEDziIQNZ393LpL3omihU
wA/8kP5MA3Szl+wzeFRh5PjMjeVWoEmCN4njCu8Qal/jrzCb8yglqN+oaAy1PTXrnaI4EGsrO6GN
2bPsU2LRF5CuYm6+TVfDyI6rRE5DnN4R2gYo1jHO6SHCB2XDb1oRyu3IjSiibx6lvP8HLpNIvRC8
OgSdPoE29/Pg7ocMsWdyzVGaamoSx24LXzkKYZCTaryYEy/AZrGWBHYcCJCA81At5X926U3iZE8h
LOBUNHlDGJabz1KA6d6UpyOaXMZVp/wIkRjj3BOHqF55qKLFzO5EARiOd9NnQ+XdoeaT2eeArAoY
LfnP081MQZjHzkcgoyaLuIXSjR1q3fT0Bzv9I4TFLMrHupgAXVB5FNJ4kMs43OT/g+S2R2wvLNZa
Zmfbn9QHaerxBDB1E+5+IcJ4WVrkJOitzzqshrGfPmAOJrqSFlu5xMd2tr1fVojeyg1DVzKBWdFb
3FpWjQLLbU81redLukjGNzWvEHLoMCCiYU1KKVcNmW3vi9ZMzEGliTku6kpgxW68eW8R+sQzeMSY
It3Sc0ky2ogVYOH4xWvubaYAO87PxLVIy0cbuD1UMOk4xeJmzQjrl3d9fAB5O6PITpYLKxna4aVA
QzgUdhiA5c5IT8bP1VNPOFtE8B+qtQJmbu7c/B31EAeTnmLd62flftQ5wCb5EnvJ/fUEz5ONz3QL
Ii4tzKlvnBY4ArJ8thyxpYb6099RSZvXKRI0LaH4YZ0iwEZbZrSj9lU0BhJbx/v9fipCemdvdMbO
K+FBBShcoxH8iHo7vMRxhroFgfm6GBTHEbaiiJtOMfpFOaloLPbyhxwQMMuSV5ViBfJtbVgYC3F5
Bcu65pQwCWkG0Zy9duxR3nM2rCpiT+u3NxuM7c2cBsFtLKDhYFvwr04kuD6yvZRv7LyAGSPXAwej
z+4wysdI+s6XKt3IYot2oJfPphVhsVzmNIFk67QguYErEZu2e5RnvY4J5vC+MUmq55WyDA/BIuLx
Njiovevg1QMFTWH990eIoI3K2eVsXzoXZpAaoTE4Vhco6CDlUR8tBDR2npfnlln+/5nwBTRhd6Hs
LbQ/SimsQraVpJv6kNODw5hjbpI9YU1ZH1Eea+DiF7J2EXsRPZr1PqQeXOOWJaXAdGBkekV3Hqgy
BN5z5xDWZ8KyXS7GGbzpbKlASUG/mg2Amiv+i86qKZGU2ZaHSgts4YCTzuFIX4F5kLjTH1BnFuvU
rIw5+fdACF2rc4FP/raG7nDNeSWG3SHTwfBIZoF5OC+bTe22yT5n99LFVAk9i6wHT1lM35auyLYT
BZr67U5FHNg6XYpSa+OGwLvV4nE2YKBizvKZyww0ikuFi6XQGZW9mV2OM/xs3DrshenoIK1wgHRU
vYrtj+ZIreqkca99Z1SakcrRjsqCpkMR6nL4DWnjZe/dbYY4xbARKBhcaDpLfZrQevvoBc+874m0
UwRbU9wD55osS7VEv7GsEAjO2VgnlbDst6xfWALuzAkaqtP3RnzDV3u/XLIJSo+F+DZO9qtOMNDt
BlQZssj9MSXAReYL0/CbGKWDFf8174WMfwI8T67OTi3jtsstywUJ2KWePo2wniaKg2hel8SnEzAG
LaudLNYbeZev2z7YFVOqzT/oDrPZNSovxgn7DGKH/ISeG7VnDKfwgU62J23EBQ+GIY/hsVC/ijl6
ZZVMP37WCvubwAiBHXCDQG/sH08VB5hlSsDjYkn+2L/dC+DywD5HcKKX0TYo3n3Ib+5pPwkBxtjD
ncT8I+rFvzgBEYHmNvTC3QMWlyLN7iRsbNRY19nyV0h7pah8ThHt8e0Dbo77RQ8SA+7LLJpvmSZl
NfbuMDEg1ItL1fTbA80/CrNgEb6ycANvyyxrbba5UQj1o7IwfsiAdy7VTDWHXAqGRtxS6FMk7Tdu
LwrYrpYdfbC+M0s1jK8KF6MLPOPtLbHhJiHnK8lTVZEast3nD0AzzK5zFAMXQE6J9WGMXIHlgvMM
8iVHy5OoLXkh89Vnetmooxk4KT0UnggZzaYRlF+9whPbTwI6qxD8jHdA53rnLp00EhC+HI10EEBp
FzJM+Rj6ZLir50vWFT8ptKbODoXJUCUSTTy60Meql71pBb7vfR5+J3KDp+09HaQcZDbJ3uSFfUNH
L3PatDUJHkXFldTdYAOj+b+YDU2fSjiBFhkZKkcyvbQzhYKWqIXOhOW35AYLORogT1N4fxJZvWM/
8jrDu27Phi4Po66fHoPgMXX9NhZIFgdhem4tSHh//e/U/E+icqF/ayRXC6S21udZBsQzJJMxMxLW
ynKYWQQielzU9hTasJgHTrurCe+XYlwmT7e6UfMnZqQzrppBOimnEX5dI0UsL2o533dRe8EIU2De
rpZG1Lssiz/6z0Z8ziWTEHIXwRrTDwC2GI/Fr7qb4aSe28Q0leCXbT3szhb3XIGCMthUAtf5FvPz
vaWhWLBR3yW5uq3W7rzTpNEPINftRso+JWAYGt+jh5ajdY+F0goJHtkuWp23jesCqk77PUXfkxdO
XEw61AR0n3f6yNbkDSxa2B2EB1Mkc5gR21RnFLCT7gtQw7937kHpIT4D7aJwy1YChgFz4RJq2/E9
RfZBXQOm4PGieB4tXYBhHuc9t4c1HqXtsrbf/iqbF+YQt5cltjRDbnlj3XYSYl+GmyNgGxHSWymT
U8gD9kR36CNop19JbQ3oT2Mi/st01jcVpjyGPt/BcpMQtzekV6c/UUrMEaqCa0RDNMB/xkaJANVu
+12ZYhrjuNb+t7ocE4J4S07v63RZdqc8/99h4kfKy18vwuZ2+eJE1T3Pm6g2ju7V/QTL+NnqaciT
yqNWCwGaGnJGG3TR3Pw5kL0Q5cRoJHfOk0yCUvORugDcd2VZphLLh3/PeQ07bV7/UGvhKP6mPAy8
UcAyyvHhCw6jYZaP6gbc/ROkstfrzfD2wiZR8S2SBGd3FI/JD79afCM5f8X5+JzdDq7qt2tyudus
XSLIGuWUjth6w/Z1NNuI+ZE2iI6RZz/DjsWrGFqLF7ESuEe/tbLG+ZUTl3o4+IQa5h7TtX6lZ//8
0Vw5avCALegF83V1y0bHfhe67Eho7Pb8VOj1p+v8CxZlyfDE/QSHo2ajqZGVPpzd12p8jJP+BHG/
V9XSXvev6BWM6bu01a/6ogQr5P82N/ef8zUgHJQqerYknkDhIDZwHQyh3halA5CeSVR/XKNjsazQ
zcuU52g0K60JsplthBGF9Mhz0TmhL9MXU4CqD0b8M39TzYYBlHEIyqSzGM3Z7Yimw0I+fKL6gNOU
r3iyWbNYBYDxe7Iy8aEpPDVmbtPEi9N/qQ+CJkclp9EcKS55NGBbznu+OQsFbpgAFy92yB3RsxP6
Rj/oI7edJDZAajxraAA/iNUNjcq6NxeUi/dsWhak069BRtP8AQv7cgNGyNDNb2ipQENnkuSt//27
VFnb2b1Bxy/9y01Xdr9Qm210kIBPm4CuMv7+z9LufADLsgwZpWl9D99aROOU/T0oYCut3M26ZjSa
tQ0ZUomWV2IEJfWLX+4dN5fQR96/px3jso7CPetWLb4FLmF5SvV9kgsYk4pQ1GfYU2+BY8KEfptr
DKsQxKq8mxwrvrKuNymlsHqVdFiopWYr4o4EUlebAu8yoi+sgEYJ16Wm8O+2ig8PgS8wqAAqjlwv
hI3p9/l4raNaTE0vC8oubKpCGdIe+f1tZdCQzx5lDGH7AMes1Q02yaB6P/SJFhrItQW+7uVL2gAN
LNyeBzZJdEVMgleTJImcHt0sK2q7elfkVsWWULWsehnBI07w+CVz9HILuKIIp31iALVfEA6Drk4S
aQQ6KU+VkupBu8uzGxGue2CphNAZrM7kNxFKYKn/GgSVqGBhXs923gKyIkw0fr65oeH081QGMI18
+/w9R/oV3u78YjABSaR8RILbvDsl4Ftdk5PLWkYl5CYhgIS6sjueJu/vaBgFPD+4qhsbWG0/mTMC
pXQ5Fi353alrmtBrRkZ/PBNVph4YE8VjAD03BZRdL4tzsAiefkmbsVWRzochXp6GZzemKmkxLW9Y
YxLfZIKkmN7DuF5tzSxws9xRj7xJjJfekczcFXAdM0YEUtVeash3OCzCPZwdjkTBXbbBo5MuDuBc
46oRvsY4AAhv9bT319g9/hPVwJ8BAm2HEXlXlOpeRME8jWHnDHSNfVz1hNthGpYZK54lkiHrtvgz
WE5C6h57P/NqfEa67+flbzsmBU/ORJV1u0O2n7vSHi4z75m6WDcwaGE9WaUrk/eLAjkgQdpteaJa
fhmtmY/ZjmvDDb/4Z9iJ1Kjn/YDq3k4U5mIJWKAlc5fnjRE1+5BJv4mDOklgjGuMWEGr01ISdtko
BluxFbt6PrVZ7WH19scjhRjtEtn4qQSmnbZzl77BKwkwHRrhxp95KzMBIZQyjWz0KF+y2JiitIrT
IQI69uL8YU5gk9SpA4iR5UEycKsbdifq8FFFqOp2nvnTgEzGPddmIJBgiTOZZ1oPRYgLc3uIsYk/
QzMENSYgLfiWcehVr9RQkDcOBAADrWYjgIPKsxAGNdallaWvKlbAHV27pytKHGJrgVl7xl345sP6
1vr59zQIwLSdv7nrKKaiePHrG4rQjNdqITd690R+Ckekv7YBDjiLSUoqmKKB2VoTTJuSRNiYQzga
uaGXcUBtP6HN5Li2r9R0KBEsdKGLfd2DhUFMFsd5dxrN7lrrr6Ep/80dfgz+rlsXyoTWJ2UggV7x
CHJNSPZPBdpMg6itY1nLGkh7z3Ebpoag2uXT8lS613uEAohCGXVs+RMyfrQy/SJoCSUjeOZmdZvH
VE7nWYg95L28upCpeWSR3tDi7Db+feW1SW4joCofwZ3qQ6wAijsr1bLjF1WLQA7QJzCxf+S0+pcI
AZVNTm7ItINMyF917agxhMMsMW+SLU5t8DmZKkzgmTmnoG7JLfXiMMf3mZXSl98fE5RYo5oyhBOF
y14AFvrSqgHPID9DkixqtgRPxB5xvnkrH39o6XJCcKtpACB/FIlKDDGLyFDmrsCDHoEh6fmoAnid
7UnqVtkdYMj2eafgTyck90lIy+yr/C6p2IG1GHqPI5oVRQT8rt+rqBkg34jws1EhzEklfUEb8o+3
xow9iCX4l1Qu7OgFbpDgAwbO0qzjRArOxMLZzfyoKYCMeG2F75lJVsqaYWoJAQpjicj77NKJIBmP
JNMsYGmqzxwuSK5gLxdYZBGiGiqCx818f1qGgfPCxSLVgDeyKZmwRCg8hMtqoxjvCAjHc9VwCctF
l5nvsI0p9k6U9HVuxwLmQTVC1yLO1UhCtdOOCrY7Vt7DTtQhxoFHA6rz+lEyHvcwQEepr0yW4RRP
q2Nckk+FTfT5q5MLIS6pmC/bfYxlDxF6rRyB5z7t2JVJY/kdsFF1tAVW3kNA+Crq7rxiEW+4SQgw
nfZ4qOOwVT75FBOl3F6bzmCmEOJD9YpTvXWvsz4A45ONAOUnsUw6YV2akmKwiX1IMq3rsKbWrAHt
FgMMreaTNw503hlfpWZ0iqsaor51GYOB9FzaS6asid5pmm2Is7DLwTNyXaY+vN5Sm5Pgv4sHXXLA
dkbVO4DqlEbu8T0yj6awjhqKa8vCXEouoWtPkwEAjrXhXmFtNgwf4YgohKQMSMcrV33uisqntmUr
JLis/VHWmzT85fQWtEwH/GZHOIMzJOMzD2QPjdhFTT6KNXSCvlh4PvU6tnSitd1XweWBohc3JQLB
L4OtlREh/I5avNzM6CerUa/hGqGgny8OKxiRYw6N1ET/n5ZbUqCfvy5OoGhZWQJJedLXx/hek6Hw
yt3unomnYZo+vrxWCBrKlQBGO3AT6uvSihpkm9U0njC8lJqdmSXkc2JNPLEFyXGeHGZGIOqB1Nr4
IoMvHZXD3B0MpIAoaubcqLCTTI4tKSZ+eExEBBL3Q9awd7027j+UU93k6TAtYF6oVzuL2pbOlc9M
2MsGfN0/YUQE/mZP5hoXdxb/CoNscgOyN65Vebk6DuJL+wGvBgjHrr41J/QrC6GPJVMZMk/uOQF5
gYn34UWFHUH7gmnjr2+meCK5PgmKILOGwtvoz4ATQLzuCqAOcQ8+QcyJI9OatJTFpWvY+0fjNQo3
MEl2AVPt8sU3c1pl7wIcTnnb+BlZgu0m6ilXvA9qvIlx0JABWvsEggxWEl1H7JJCJCqfm7Fq1Jpb
a80Dhn0t0Y2lVAM00Yj92A5PXvUV7zl6yRC7ykTYZhN32Jgw7IVZkiAA4rXXyRVSl5RMXZG519uJ
LEdIS3WCz5CW1VWHQ9G64Hpk1Thc/SFnMStQIJ2tNxJgewOyW3w1Pcn+dS6JlnVKYNPutBL03p57
O6dij50ku8opym2vGowyNybcCkUbWAQJIroxSMqHv2bbaesFhlyGjvTTRRmU17X6YakGp9Bx7ecR
oq+j5HTeoBUrXZKs/zzewcFsXXyDw0AhulGGW14M4yMnQwsSF1srM1rcYFkebAixEu9+mhDhmJ0g
IA04OIIcK0IF9Iy/5gPN1UW6t9klM8VYVCPbYA/UWz11H3ZG9l+3bAzjjWeq6vaAAI6peiHRfWoy
jz3aEpQwlLZ/LjABrTy3agd+ye9gBWq5e5/SthBKMijzM49V+SKXUDTioREsUlFXJ3OsS050KFVF
fSIj37E9m/yDGnJLIdpYh2NdHsarzvFmHIVQbAFelEh6kYsXi+CSB4HyNCq6pkrQl9qZqQGfqiMa
dOwfBFr8X0WO/o6sVMO0aG+NZU278t+6P83aG+1AY43s5/GuLD1YqZiYnuCBCBWJrHe0pv2QX/lk
ALVCu4ybCHNFabqgQl0MnfZB9ssxlwTJUjGXoo1awCuMw0ZQ2DUxLSrzK5RvVd4eDNRCIj34RseL
v08D9jdBFFkGvWGheYNHEahkrHcTs/uJaDjbJK2MIwWMPugy7JC0lH3muSe0GlGl+hIdB1MA9Mcw
+x8dIOJtpEK9bsct8gz0pyptyPlxOh/Tivmx+tzw8SI8dnrRG3rvBjz7LqBELGVLbm7FcuI+QZzG
rVCuAB5biHYrHz0tMlW0l575yEyTYyAUdz3mcRvK5HKAQhkcohPYIEXQaNWVCJTyroMNGF/pS0y5
39y8WyXuf7NJaUCn3kCxjo8D9yjuJVOc7jigtE1RXur4e9rvpT+JNCedRaL+cdEVlSXksLMHi8Rg
VYwogv88ElvOxIhvfiL5SiCcLA9G6m59AAfoYPM8msNFy77OUPibaDEOLdD0rH4x+8Ny0cMYcxKf
QAcUcJ8GDx7E/qVJLHEfzUy06bVeYJkd13MrVW6BL29HEKjXW/nJlATyICCwzpMjxE1MuRl3yLrw
D2zOREtEGsk++u643ro0R9Tixz/ge+xHqZxRfsJ8HD+/D3Nf1AcWX8JIhjdSO22IuCSdF5mD4XrA
mSMJ9vVINNhatzK05yjTi7bSNWG26hQF8YYmcKyhjBLRNvjsuJJSGxMuzPTc0kd2iN6wKKUk2tYO
208F1mAciUn0SI5O6+AObOuAZB6mBbTV69DNon0Uqwc/fSIGksaaoMgOcA7VMNcPwno+9XSTQpaE
ywN7NuxqHhHyP/MqHA6BXQzsmeJsDaH21GuZgdt6vLZOX46XWuSb5mvV52mRumXHvWIWURhvlq7T
Fq4PzJJ4l2sF9buh6I/Hg1C2Js1wkpRK/7vvZSPHo6nfMpu4h27RNxA9ImHU/BKxQ7qPrJ+aos+E
60Z97k4/otp9cD6bDMjV3Q9DRyLF35LfgWSOjemcE+KyqYaSHn2AB/IOReADOGIVOdV+UNvZLbCs
6thfR0Y0KwxgWdhmOIPb/IReyeroPr/3DFNcS8qrlNSnaHwMPHZ7F6nG4Zng7tuOSUXodsJJF6Is
aeTkfn4eE7nQN6Jnf7VLiy6jh86SOTPRjKwHaUZsyWDyyAb7UfsqAF8l6I/iOsDrkzM+aZYzEaxp
scIp2WwP+6g17auCbCBd3BKb607QDgPTQrIQN3FHzW1Hg7YW4OxmefKVwsDfAHEmAeTgrH1w/sDt
20JHt/ltXfeWxipLAgMLsw5jjArucB01/eATjTQxUR/+fDy4pKqiBB6066e2Isnh2ZJyOaY9hq4l
j9mArwKq+y3Vfjf5UssW6w0YWR1oCYyz9xtCTMuYvcs+RQC8rIG71Tj11pmt4HVkwZRtCHmqakK9
U0fC9frqEQhD8bvDshsMzc8gV07JmSBly+C+5c6px5wnkKz/4RXiRWNFaoyJEPs7x5FlV2Jzxdq8
tIwDNeAzDHxXZT2c8IXbWWJjLRTQKDbYyfdrD0UPxT5h1AylMRaW0cLBP8jSpZawTsYju50c9nzJ
U+GXq/ZplSfVA7QzwUDKPCtl7QQ7ZVu531yDCahJKCZhO8koQ1yErDl+eFpxhtNMAPqnpF4DMZ42
e/hc8AoFtCv8h9nxw2S3t/I9TdOvTPppGGPLJd9d1xQLc73hQZz0vvyaYPbPnLLD0usYXtyVxt7s
WEEDFHCrBLb7mW78zDmFQwH89KtyoNPq/SwOZ6QKaJQlFuS/l/a068lPmMcIKMT6E2K0T6okN5aL
IO+CYpVG47QivNVaBDlqhtKQCQik0gBasErBJnmzKuvb63dF2UQOHGvIJnarJSoer31vQgwVNNw4
RKPt3pD+tW4MXoKRepGmoyM1RBWdHrLokF0W4+Tn4ynCo1gRCxzV7P2bMhMCLNSutgGYa4DP6y2O
SQagnWOMu/llGIqQwfKJ92gYP7tiqJ9AaG5wX9XdG3oTO/dqD1jdJAZGB2jAisbTyj1P82/AhdkT
iQsfeTY5VGA4djkKFXD5IRcprwzrs0aZ2eLq46Rgz21pnEQrKkkFw3gYlA2cakbeqZg3WhdvmTxY
WHmHkLI1Cxk2C1Z607SVIbJNS4EB/6fA8uASmpMxq9vnGTxaQlcETu9KbSblMkm2mawiI/YJ7oh0
qz7pUZor9oInjKCkVlBsLqnyThIfuC1CN/RylKKYRg8MvCdM0/tqlSJ1IfsYXasGRnh7UX/ZfucV
pwyWNjELqxAkyQKTRNZoghDsQ29Wf6JVOTWJ8QLsBZfuDgjuWPBANOFhGSZMa0LtEa6rHsNUyfB3
f7qmp4fPk7El829V0ge1lrz1wFVkzc3Rlm22jFIv5dlXK+aQoGx6KYrLtuN9UmOAkpPgEh9YtJXS
eF+x4aaJy1wp2h8M8KzffUYtHdC+TWseDtrsdvOVNFZwaIxQWIPLIQZHgkTJ6mD4/X5suQiLIzjC
Mw6gjYw0YitAcwybxkJ026bawIKl5VugvTE8/kQJvTEoduG34ROuNHgboD2Sf86WmhumcpMBzB16
rCbdYTdFGvmjSQ4Oe+ZM/wAnhzAWylw6S3UV8Vp2LBmGFm99IFRx1sPNSafCQw4AISkkbQWXyFSW
S2P95Ak4JASb0Mr4CbPPHUDYrq3Acnk30wdp6UhoXQ70+RYBXO9c22QgRnV1T74PCF9W74VWldTm
IyqyrNJY8ZiXn4xGf5i7nJ/RuPTDMquAuDN/vXwJK9PwYpxxXWfwXn68kt5578PUcnKXvMfvLdeW
dd/+Nk+fJzpIecTDFGRV0s7GxhJdBxfQb7/KzU2EDHlbILL1q4wlR449E9HOblSbVrXyWXk3hOYk
IEJywsQdM0gSJxaQo86aWVORy7jF8zKJ7cG+2M6Qdffshq94rd61DIk8lmnXXHHsSrHKlXHMwJQ4
aZWhvBuNOId+5ExgFfOUmpFR0puCA6N6V+1Phi7o33JYzjbgn0ZJw1k1LbJECdCtRQRs8c5nRBp5
iFel7cJuQV6DwCiRoEZkAHwN30bYIuy7TbHYwgxJpbi9hVmJSrzxm7cPT2kfD5nYYb6YDkhI4LdS
miUwDwMFeN4KEsqpoMKXFLPh1rSe7nQrSCw+yGlWqK5rHjlNnPD0bmlFxEQ43ZAIDT+Tw0RbAsUr
juFj6WjZzh969gX1aCR80fNkZBgVEZyAW7J2VfQKHZXLaPZE1kVuQDtK9Pp0KW0McKkTZkRQl1Cw
9lx2XOsgtRjpDdDJT/fiiMxwplE1mrs2QaeNbU0TI/z2iIjkvZm6FlRlhSPchPh1ojJ3asGbHfF3
XXraSqyBOUuL6Y9h4DPEaZI1zy07RpvgsXMHQ/heUzhPS9m58YYKuW8M4QRSGPlqBPDpVDb/bq0i
JuyKWgG4zx3MaqwQuGkWQz7PCckkmGQUW2srjcGi++zqAWM/D1OMNM6cGFNLb19k0+J/uh8AG8Ex
DD5eURGUtIhh+I/1FXEDluPWlQJDAIZ8IgQbgHYUlx0HTU3omMQVFFt5MrM8r1t7q8g4vsLB+9Bp
WRg9bRrmihW4w+6fTB2I0uRSAqDCmDbfFO/HgjdpC6Be4ACrSB44IIDC4DzeyC4u0uM/8XsDLR25
o8Tp0iakSIwYutdDQxagJl3Kl52GfuHXeek/5Wo2b8q1QpKA42KFiwfTVi6n0xbBq0mJrzOlZFZ7
3Q+SbbVyHVDUlZJ5t8vZMSWhtndv16HXiXYCURp2jJuU4MiTM/uNYjalClSyF9t7GMrqZVMUoxrU
uguDBdlm7L0DfMcUY7BrWhmasz/MptRSKntkq2q1PndseSei5XUyrRahCobp17+YhfvAgfkhkjle
nDmBwV4wkDZqeln9nYvBqS6F4Y2heYKdDHDuKkE++FeEosMyE6TVnjfDElf+3pcb6e12j5mVcHUl
vQTfkKSgzmKmj2b/CIknqoLad4tLHIkVbPjkxkbKobya74231fVqYaP6ZOLWsLMxhJD+mFQIHYAy
FDthqs5BKp7SH4gRIMiJxFKCz4fdGoxOsMiPb5v23uTgVB5lW4PXf6bL3td6gN4oQle2Ic8OWSgH
zOFn2H/T127HH+MBy4dyESPmP0JeBcCrWUmB6OYtCCG/fYrdbmJ1LIKY1kwassXvyqp5O0rC8gzw
6i9l5bYDI6znvwsyGKQNULNr1CXvdNbp/MWBPxtR5XjO4fKzDjcA8hBKrdP3qQigyX/g9bX3wXEe
YsiZuMjLshHkefTAKcfs3T8+j6YWvFbh70MXnZ062xvo/bRp6ryGJrjJ1RVy2WDQkaubOEV3ijqU
+K3fBeQqK80js4EIfxPh+5nUthoEObM63sxoiOmqsKfxXVPzE7/+rSZLVOPCMyi8bEN/Yelm201B
3k3jc4LhG7WwMQfh5DhFGX+6gOeaHMlGA9CwitEHeqC9JZcRECmYU1BSiTkRbt1ayJIFLpRMUNWS
icK5nHNs06Gx64fvUWcfpWyYyAcamKEpZs59gNk6ffAycyDuHRQypqlcg/b5xIGPyoEScrOMtO5i
tOF8vWHJJwRJSROTH2yy3Awloe5U6G2VLFdD1rSDLJiMQecxI959IWAX8Fag/nlPZlwkxN6XNQCE
ZkIH/kKDohlXLzDsMvDn8dlQwIyv0v1sgPn7AQ+oD2BajUST2qGgjc9ZEQBoxr2w+t9eH0suztN2
u0swwvXYt8/srJXM+OCeMmowqlDzG1DzK9aFJHSQgZl4KmFXf0q4v7iMa+4/jhWDkC7cpPcVXor1
CKLl/Bd7k2V3Fm/lpgGI29fUXIrQJbbRKe0M/6r7h3Cy9ptDTRMHmeCTeTkDpcEaQKGn8IDmuX1b
Y3LRMWD51VxTbmGFkrfL80In7+7xypv/yCKgr2jMNCyT9PHNMQKbmPMtatbfYF/Hv2QnxRMnmYB1
Lhc422Kzr7HXAoxJ+0AJxxEtbk7Ub+7MINe6Wq3+yIqunAr3R9UKg0L97px3zVaqWJ6UpYOwmgkx
JBaHMQDPrCYPdwOvQMeuvnW3pogMd4+A29hdOwywNu5EgAOxpy9nMIktZRn7++rf6BmjfZCAzScZ
eTJCJ+jLWlsKFJvyMcBdBh6VAyBsgADYNgo/E1eIeM3eqexzXyyR9XGoOdhRy/5yqpdDwTJQAPuI
AYzY1DoKHPxSNlVpaK1SVev+JBtXsaAm5tQzP094Ybqkv1/EPbHZHnkVXQo60ekusCao4mF8gmHn
edLOb4EqbnY/rzfzrXvxnoehVp0FhFUReNmFlxzHGY4VGEO73/vpXyROVGa4MjlAgjEAv28UWVuY
gk1bp6bBYUg0iJwx/spUlof+u/taplNWLhsKjxTtwdPqaBBASotgb8d2DqKTd4u7T7qG2CdN0PaQ
MPWGS/HwItDLjSb5zt2LKRb5sUjfLcavltmapDIylfxN5D0OFRlklCK1zB5XexHqRcbjbfB0nZ0K
fYPxMMm7e+CaZbrg6Zqm4OHaKUbAW9uX9cXnMhPdNvJC0A4V0o1kkjHVJWFFounhH9wqK+JckwnZ
kAGhHW/nlEvxqgJ8iaZD399eDsjKV34c48MQX10/3TXH898+DjoHQs8huVaLJ2hvcyElIex1Z60T
ptFKZumdMqnVDjEDGYFOsnWueNLXiu2begQId6/W5ZKpik/Ohsv4oKN7VIXXz78c2SXgdQ0Xi484
LMGbbRxOGgeAeYRL9RPuiCF5ePc3APnEkX6AEdwquGb6GCZOzNRTSlNTT8U8bU59nq/XHMg5RbQM
kH2n/ZSpHoisj2wygqgipxrelAHn74U6x3P1GrbnLmzX4ufCq7zbCN7GQ16h9c3yVLUOP0TZD0mD
q8MrnVMHWbQKDs6hCha/FvKcPSsMUok2uXgq4KUwHpOb6zROi34YfhFEt1z9Pyp2Qs8VKfgUu9/9
tq2LMlx/dK7EeD+fFOjUBCIS3RpxqfeoU4Pr81jiwwTkK5x0sbDVvpDAK8cfBOJ3R3Xi2jQ9/Vkc
rTa/LMiVo9jzlcHAX/1wNEqTdVKHlMdEZAlxBMhe7P6aSU90IhYDgYPBcDPyLMB5gJs1/h5LzH6z
zWMX8WTJX6MiebIrSjAn58ORRXr/OWLdoSa3aKo2eP7lvxKWvcRWm3N31KydQPGRpRfvavF7VJ5K
ZM2Ov8vor3OMPFAwthnxpjwAcQLN+Uth/e/g4UGcVkaT65cQpt1uYd2/tC6EqOcvnLSRVn+73S22
iavKfIqRSGk0S/uG7iRhT4Vk6utNEGIwh5AMBhpbGDFDTtFHlN0jgc6Qg6MdYdRN1KRNUBJeLH5u
zj+P8UGq32ab0CMKcrKocIcOqasfEastDOrN1ebQ5KvgPfL35J8F3MvBrG5s1wZxFJg8X3a6Df/H
RPmttn6AVsi8kztIidZ6X6pq/pbn8wbAmE9+Lufe9Jqs/80/cm2Hp18g98pz/YHmXI0A7ZPYSJoY
6knFHq4DbaODrYz4icIu9e6mHQgTwEeDR/nEGZnLfnhbjyXnH4voWgB8w8NitPmmwfUKIWxZKmO5
5zno/71pIkPcnvBRHVh0zK6KSzGs3rMQZ5bfNQ0zqy7MsUPVUCRIEG6KqwlW1sBccFBpqWxudYcO
2TAb7IRRxdIv5c09w1qepEMBc50iZ1VCXiEYt48RHQyL7KspPRCuKx7OhvFJOGKct/Z83ejojDKP
9ZDSapB0AAXWb0PhKh9ozscy268Yo681eVW4aSp2DrmGM2/G78YZd/sVOPAtqCTl6bg+GOeNQ5Vd
NzeEt+4w+FoVsHYazUIXr4wSwaCXviLFdOjkLm2tDn3RpCfiu286vensdHmOVxqNnJgOjT4pIRom
vNkMHHRCK1yz/qXgSZULxSCef2lQ9hV20NPqHpmcb57FcT25nYbNHgGtmjtrAbxSMXmsm0R7Yhv+
R6X4E1epk+AG2LnItyQW/B719kCI7RFVFUDmOFeHQ/+IbwXSP3Kd5e8k1bA0rSw6m7diuFD+BO2L
Oiki4ToO8XINmMv73dTQ3Q3Wqrnfc/RAKXhlKItKqTQMsPeAdW611D6sTNxAfm6KWYcKynViA/1n
Lfrv8niJkyDrvF0vowMSVrkiYVWY1ck0oPiTyHkeWcdEzdLH7HePnqoKx3kGdo+WWIb0NR2lxKhx
BKtrqiCD8L4zywNa5YCXbtGCTuXXUqwXLLmr43MnIK9xHwSnwU7trNt9r6w6nORovh7XwMnwwV2N
f0xtovVnWjkjym7Y6IHsxfC3Ap2gS+TWw2WzlD7eJbcxFpwHMbdGnFBExn+ZkcbpQkQvKn7wI4Co
JorRvwei1EGjTrE+/fDesWHAAfTaRL6/qH5Y1hUq37ztmZ9Pgd554t6STP9FbOoTcLKCK0ObNSKa
Q2P80AO5cLeZ9cRG2YoJRImMgdvhajzM518sjl9rO2WHvPwx9Ma0NNdTVrLVkP1vjV48lRePVi6M
RkSTnn059ez11a8U4AVGfgJhNIkbOn/l7Ch8Iauix/5SfJCE5aJao/SIt3pnPI359SaKLCa9YDYS
8zXe+Jwg3JxdI4bA7GuslUJEiW+lzEVz4+vwnzZUpPAJgcOVzIaTioQzMujbyHquA112PmoX8lW9
8wNCnvd+YGvGQFgLHy5ZEWLDaVVLWnUHX7c9ywejCg86UCIacjJJcX+D/T7TRaBAEUs5mADowU0g
4mM57pHfR2GHV2VP0BbVtLXLHJSbqoPsiETtTGaN5SG+yvTNulqDNjnzokLGXHu+yOXJrhzSA/vY
JI7SZxcpM+nNG+faHeArJxemk3nQKmu1im8Zt7sKYqFZw2bixufxxJjH+ynmVqz328P69O+yfh1Z
eX4aMADcEw2xblETVhIWQv2qx5rZRLDzTIGBhBnvjgjTb+v0vT/c8tEHUy1uw46TXqJVOJhV7HVF
UTlt8V5baJH2KFsWv4++pxvMCEEqGv+PZjGjDOUQ7Int0SlGogh9gJseZo7EBniw/wK8aBL2LPkm
WqalIOtK8R1AArhTmv4dwScOD5ue/4POLBVkViUL37svDBJR/1EaMwE03+5+IkRqbKoza0QAPgvk
JiK3Lsln7uxbl8wVPUqFdHlXdda0FocMJlwQSRe0lRr/X+L8BSo+FKOJ76GNzIRLmNtG5f2JdeK4
Aor/Sou1//JRke3ikWIum7RlfWbyh5s82bKKkbpa3R9WDQq22eB+XohYApJVfLUWwjyeSOrNq1Mo
zzWAkHSlBuDVFz8HZAE9A6KUAfirHiTw+0p7QhSvq3j9kC7Nb3RcitVVA8TnOj/y4n1k1RNXCkCB
6Bc+J1R4r8rHCx9pzzI7UW1tD/5UAk9532mYrF6pSjO5OK7QVb4RCXWE0uRLHyXs0Hm+U79viQNu
KEVb/fhVU1aMW3v8qFNnud5S9GlUizm33woKlnxPbf5icBP3i3ju6BdGewABvRuRNekP4kJ/6e1t
n3M+gTjjsoGmsj0xy1xqkjEF/eFiVDLfPzkLhnhBCseaL2LtTgE1+Z1uRfpkmTYtIJYyYscZUw/F
AZWCvOlG8A+8Bka+j0pINvRECszUJfKRdcaXj3So3Gu+TF97Edoli9aSGgDo++dvMTC3/RzbMc4n
hZPsJXv6+LtYvSxDwe+NB3eFJ1lfPM8f1+kXn2bcFo3xEXzm4PyOyNZOOUSwYK705jXXwRp/5STm
PfqZEdAke6MLCAei3/ch3cxHtH2Cm41l65MI04TDVB8lW9oXRKDrk7L4lxDEC2jbuF4rldLHboBu
k19U4Sh+7LUezVUU+gRKbnzv3FFbYlHA7yIuiNXKV1Uu0OCdIrcwHkydXO3boy26CdSJTRpQ+gou
EMy+UOHgp+xoG8ZjGK+4tOCukgUILIRN8LYMPaglUqpaIMDk2rA/40kKQ1u8Xb8Zhtoqv9Aoxgnd
zETB/xPPF3q3ErjCsPkslOTO7Nc234/JK1hTx/SaIQbrPTcMrX4IV2Sjr4Bepk7aotznrsQQmnzh
Wy57qpyjBeHblStkpfE9K6W+0sOEHVv8N8omH5pKslKzMahmWxTK2BcZYZC2QrL997/vOAApGoMz
sfCLjFErALkRqt4cy1mpyx/1iMVJBvkycjNYbiMzYxnzLFljsHe2ljNAGcWIxJSo8tGLfAeoNglt
Phi7fdkiM8Nuzbt9SQUXdo4efccU3dHlBZ7vlbaYwirD6YvoS2RJjHfB+vjlNQ28n3SC6prV1ymY
9QUlHqm0wigvdPk3yy3IWR0++5uTXWizEPdBdkF5wkMR/CfErwfvZWT/cu+Z+gw0CPtSvBTNerCQ
BV8RAJPz6wQhmbgn3auWDmaKH4U+WVW3VWVJMEmXBZ1DnNC3BhF942eQxu90/oBk4tIrVHjmZ9Lw
73W9sumUGnyFXzzD+ti3aBd7Ithx53nVbVZTJihpAD3Q1retHtM+nVbeJvBf4Wyd8XXOgUZSq/SQ
0NOMxeT0ydwGeUfLYbJ9euN5XRMpUD+c7R8OBMeAhc910O38Bllrzm63cbdihATScD+xkXKkdDLU
MLIgGWX72pn/TPZNeuyw9TLs9sys185Ni+VbkLC5wwr/EilGy8/PJrzlXJ44wlcrRb/KgXXiuBU5
rReRxbiFGHyR7ERKJ3zWIqwL1dyauek6DcEfEW0dXpyj8FPfvvimTBPtgGzZ5fcd3Hczuk0EciuF
l7Q2heQrqApkhEf5gQFZahyThzibacunf4AIHiApTVLXQSU18+xCxoAEKIVeuqu4OTdbrWlvKUZE
FGaCefFn9wlWkJNHwzrZ2ycMakR/aTDu7qi1opgKe90rChsTH3iIO69Ny8hBIRJ+acZixLom2js8
qI4efcUZQ8GKzEJElxX2IGDOC2m419cdoADsAuftbWQvXIBWVfd6Ipuor8K3ZxixE3J+DiNEV5Y3
fQybI1ByJmndjHrGzJFZNJ3f5oNNifHBifu4vJ8P8umdriSgIMXjhb3NFGTGPjaHw9+cj3Fr60ZH
vNXZa0h0NvRZ24Xw+nIAlb4U2sjDNl+gFUkgudkYbFmGRxe1qj7nsEttqNzty+IGoypq1dz2L8sC
9jgpMqOuvEPbIMM5A4pZQQ8M5WdKpE3UT4iom/9cKvrvw7Xl1btCow0xyIUpn9mBY00L8XnHguuM
wyUqJn+uaMCWJ8YrF0e5ai2KKZHcti4S1OEWAadoQYDHNqrzGyR6yZDNH+8/SggUuHbeBZdPflKF
JE44KbdxHZNBvoEc1HvupRLtHvWFNKFWBQRZerC7YUu+9ME0SRm7l86oLO/ogfSVM4bBUDX1lj0r
H3IWFwUvVWvqiIL87xTiHj1ne0TTWfB4BOD5DTCIF+WBfYksUfz8RFMq3sHP5MwFcuyRjEiE0xeS
do5pAmrHl2N0ooqAzLakeAASWeNQ1r7xpkwi2nQWEvT+vSBXZHr4tMFzPz70SzeaNBYe2kW4cBb5
bRBBImz1WcX9Fy2abWu05jsiPSejYlgd2lB+r1EppXxt0HSBPehZoab40sgyajo015qOcIcLd31T
lACWD5q5C8hTHXlQQFi6lrNdkgAk5wUUyVqRwaLlVh0UB8G8+YZuicMvKocrCJhiSzDL7kC5bdnt
lmXC3Nsmkuvw5hKaJEpGQSMHUrrXgj4JSJLtluYMFP35VEzwTCVj3OCyLCpU7ekUe9TfytcUe4Mw
soyj/Jid//iAoiYM5vghLLm4fEdCyskyEngdxa6dBOYqR40rASjzy+ys8WnZk3xDIsXkwSxPKutC
LAnbCutUwFl582jba2o6cA3qbTez6D7nI/CiCJLrkkczz0lfcasrGzHABaMU5mHrh9uNnWfJM9/+
ycAjZzdhrl9fqGHYCwsYcYzMGBqNBNihVkE9MMeyjFVs6slSpamlfXqEwkpIIy33PmHCJGB5ZJE9
MjrTheLZVnX5LRIMCKybAzCPHURZOr+a/tul+r2D/UFZxKqE9C5A0uEtYHb1v9mf/QftS8OGDi2h
p0iiMkIxcaQ131MhUVZ70jz+FNIxnlYRgN1EFLUIQe7+bPxZJGvt/PcVVgQBgxG9R8weFehsO4JY
iRimk4sm/4tKuGqTRc/vWfanaONuGvJ6HC/lJT57gQR3eCR2cIEp8j5fsmzxow1GJzSeaVaJKYBf
wYbGjrAZdfijNVSXvydr5o1Q2dj3bzS1UNDPoXG+46UVDXCGhmQdaN1f84Zfsl7XEv47UoCZKxTe
mdSv7aT2XNcCJwxZoTVrUMFF4ABd+AV+J+y09GGfcbT7NxSQp71LxdwCJyuJ9Vs3TBUfk3zDyyBS
So46wDnNuvFcm4jcKsHL/F3uNGnuulvzo9Pe6Fqnildy7yLWNMZ/MHk7JBD/d9ElCw5z0BLizrAh
mFihX0M8ekf8+7G+BUVkbxCPmLoz/h09TdxpMEhvQVLfGz1JZ1+6TXrmoZuUVdzqIbVtJwkEye2O
nycROzpOvaIuzUrDSzojkLT92b19YqudnvHvTM9zGIfLwSY38EKX8zFQnvHdLprakjEsWqmL6uXw
GzSWr542dFdZjgycyo4K8S/vlCVA7KwXL8j/WvnEDhww3p58UXHE4QXS2IXcWyQIrAAU8S/6YfdJ
UzQ2oeeGde0eyu1vk5XQ0KANz3tEWIwH6fBlaXhxKToJX0FXEPzlQgv2CgFfOaJKPqeoc2oNFzI6
OQ4LV5PtTlYBCefCdu+JqQRbIFUe0cAqOZUegViIZxlcxLA8p/JvM/HjpcvFswLQsZ0RXbNsN2vc
Yvs3JY9Zg2/kv7qpnQ4TazQQyBcxg2HG/84f1yTI76MYLTyEt+u6ABn8Lcl81VdBbnGXNHVFreB9
CidEEahhOMZEWaa5/vaRrCoBLYjVbYvahD93kz0MWj3CSLMkm0HSIitC0Rb5gLjPuEOEXk9eL9EB
T23BQyHaxgqVZ5TAZZ8I6grDkoRkPHSNw+RzYl7Ss10Guw96gYluwELidlk4rK9I25V/qeaKQchP
4p0XBjMMhNkMH0M+Ad5kV3BJPh2+vJPf1qi3TgGNVcK9M7giuTevKX7GTrpwugBde5JhNNDUyEFw
W/WO9yyhFKEgmXkuj6yKGsq4/5piMdsiLVWy9gBHfkk53eryKo+OobXTX+5ub443fdGXkczkDnG+
h1SycTaSXCqfuQbQqOOKcjedFD2EGuj+QC0YDBE8QDmcAFu+xRvbE6xC7iST8FHrUzbfZg9DtEI8
9x6GGd0nJnYHwxupAPAxt9WPwBpd+Cqk74knYzFMluFY7fhypK4fPGBRyO3Usp7My8nu/+lDbxz5
PITuZs+qiKgGKqSYcVvVZeQRhMgfHbVTdFb9EmM7IAolUeWk4Zb4Ij6E12JDfj6MkpcwrVD4QDVm
Gv1+D3DbOxX6EqKBUlyST6JWTE8BS50wYk03W481XlkTmB7jDg2/0rzM1KFrhF3/OTXm0yrvmZz7
g2bDGL5dDgM/IjYDtPTtHHhJLJ0QIDstMO68TXJzj4CeTvlMgPCo1rMXQo5ye2x9h46QBvbBMh0l
S79DX9f/ANi0KqIHKZnvGNQHfTx8zzDR4oBRIViTLmbW2RPaGXDJ9aOC1jwG/ulu02O2e7QdthD2
hbphhGURCzehZLFkdlMqZblnS1I18fIpQXajIEEBGBlutvOaGH9fZUf+zWStoMxJkpFQLiz34ugB
pnjskNk2ZkaaMlrVDz5n6nNFgv6b7M96VPXsANsxm8zXAR8xp1pC4+++nKofAHTDUbUfrGVQePqO
ThUR3QYvHd4f37tHcM/B1ahC+agc/4djThXjnpCGu80ZlWyqCuMfqBycHNrZ5SiNXtUMpx0suu0m
ducJRt19FdwVyjB2vuGD7Co0qO43v51vFO9wkFQQp5EO936CwWzK2dj37FWZ00GWCTnRcNT9+YIO
qpQ+HpVgibUNFBcBT+KyD5oBpubxOjBdgHkXl08Gk3PpNDQ0rLxulqNipfDb4NYgXgjcYu1JFUr/
lixyETuY7/ps6IVTt9ikiWIPTkK1OnzV/QsktUpVPBh9pAa2fImY8WQvxjWum8yJ5uC6tSdPElOF
kvHE8Ty4iJICqNkLT3ID/+L46fyjJw3Yfm9KQbGYxFpEiyZMcb4xlbwG7eMtuy/gb1hv6noa/rR0
IykaGfZ6TF9Tp+uabTGVKMYbkokOLoz1o5m8Jhr2ZEZAyMEi2EITp3bkEuX5GYRRpVf30hulf2qJ
TlSovfl0BbN5Bv2kv9SbwSs1gMo93JiqtwQIlaSsIXCHUCkdUX+FWEnQiRiYnLwUehKGYBz/uQHc
GP7LJ+kVMXsjbomlguSXDbMK71bAGtvzyL9xTLxI12x9q+7wak2W9HlV0Oni3/02C9y2LsBOy4Vq
IoPvivM2py+2K8ZbrmE8JtOO254xtOnWjh76K1kKTMPt47Nzrj9FXyM6sBzhdPGAYE5hid4lt9qS
EkaFC4GEAA5MLAqD2BwRZej+sQHXBqXe7DuaEdfELTI37UHeOIS9Yl5yKv3+2aEYW1eUkK6x6i6x
WAhPqeIpS+4Ho39uq7SGxYiTxYwGy1OBGDTnQ26R6qEhcWqu/AZbqloyUOmIygXUbK5FRlLXUBf1
HtSe5U9l57rICNI3lrNWHGs7UcDungC8GVyGj3CaPtjpf38hrn9m62GpHlnabPr2H3f0vy9BKHaO
o1v8D8Xs0SfsHpAQXN/jOC1V+5xN0zAj/OavGsfs5mve0FWDVeySPHbwOa3HEDsKFlwXGxdwCpXg
nDzGn8xj02FMfBF4bU1p6yrR1ZkqWRQatH1LuERoKLhy1aI5msZ3lGGUUt6UyFcZwOAXkdFb3n8V
MxLYZtOq0rI73jCk44DiXCRjvYq8Cr7G8T90OLpM18HTTp57SgAvj+Erkm+N2y91EBf+nxBuqk/p
nqTb7rURiicZxEgwI4X9t0kh6YNXrmgsfzCy8bsBfzXMdl2SdXGcAsNqsxzl14yw6QByUnCs0Dqf
xXuZMKDE/nkQTQyictxA0+xzxsOavLIkIyWMhcqPnMtcXcyJqNLKZtwDf8z64AA536V7bo8LEy/1
hSvZnCHWHU1dbX6BMRYrt1WVeRTNHOD7soVZNO16FrGgk68cUrPMv6LdSoWZGSOyTXui6G7cz/pu
qU6bXhJ8pLrbuqR9hvjXsV3AvKD8v+qG4J7fDq2soZSGDdEIeed3hxwegc6cyb+hrf635clciBWk
jrqDQjmOBQwVU9cqHaJqv321wixUbj/QELONlma3KmBs5aXZvD5wXIrlhzOvxCDqW2AdiB0cfj2i
5f9dhTjXzXQThpGMRonIsdosH6/jROU+GRr94ZBggqa67xD10Neg+Go14Bt2zuPQ6aast9xgLLzR
F+6LCH6D0C3BH4XnDZjWBfzvf40g4EP3X7j8SkqKccckwnTsK2olsrXFM2KfL1IPyKHuuDbYCrU9
W1iHQk6Zrm3SqD7wAkCyOWG6aVUkHn8id+PEo7/6bKgbcsm2I1rvwu1FRZ28o11afDGfsqs1wCio
ebm6Gs1G5h/neffxNtqik0B1tK9wCbN+uVca3Yq1Ii4+FlD4AlgxKGs4I/wM3S8EM1M6557gjF+r
SrMcnMTV/q733rZhsgA1dvyMqVzmfurYctKcDQvpijHxQ+2Q7EWRCgyw01aq2hFG9vHoUy6PQE8J
LoZ+VtuUMwzXX6un82wcz7giaiFykZgcbRXmu00epdhsMcebpw2qcBfNI8VzUsl0akobEPdaMeTh
xKnrQSniZRBrSHzVMiA9bkBkMNi9yHgtE0GBqnf9quCJfLp6agnqwRKkIMbAbSrNZc6apH3icTCb
p5cevbwKnTZH77Zz+L32qXXlnea7NlDdts/mNblsWqeRyyhPxgUZavmYwSoyY5t0EhQO93c1KX9x
N8mEhtFL1oFR3exPx1QH2MgCZoV6D/vIg4Eiqwan6br5toyw+JiRhTpariPPRRbmVYHdwu/UPBBN
iKyjxaejgRLDFFlUIeoukIeD/7Gwa3Ky+355INer1DD4im3v5F6A4sGblUzpM74yXekP/BOU8+0l
5BdTXnmDr+vCF1G42gX3XXqVQWEcjJNFdgze5QqAzc5RJoPSYV2lIlHGKejF22EoSOElwv5MFtWl
S+gfsWL74N+rYr8GGnHdQD16IiGwF+hJxyrjvFw24LQa9zozVGKBdVII5ewZ4ldc8j1SZgfklP6c
Uw6bNhqFYnKM9TjYfglE0XswU6lvjC1qIEm2+NyAfuklrtNtnI9OigX/bRjn41Smfi9KPvBGylxd
Cyj8t0UWHVS6INBCQ7qbEJ7j0WOK1miglhsJgX0pS70jJ6VzwiWShwqPP4kLj7N4dRFIhPq6VMOc
mGz7YWPXQoCB4FHtpxtcJFU8q93meGg66fM4vNd/TACQu2yPIMTCsZBfAUbuDN60K7AtGiMePodX
xUHY/joLgd5qZY0C+b02QEN3W6OX46XWgKppb1A1Vt65qfHS0XiUl+DQqPivuT0YP5LlmU3SZstx
uywcFF4snkpWByRYBMwF2lO5JB/qHoHgMeNhANyVU6S3H1VAxG5HXa9HbdO6vDZe5Hyp+QLFH34M
0i79QTsbXRPpniggBuNgHxTgZQ+nqIkJC7qpBPBZfcB9HXXlDHMdmV5ZvNNTfmdhvEEkDvKV8Ek/
+jQxnM7ltYAkvo3lgpYlq8qzj44d+Cyr39Nc6+PfOYe2M+ciw6cYvcBFWRBxDIMXIgNpzWhyurSE
yKXSPpJ9ZsjSzhKyaZNH7XD7GvRyFPJ0QboNsdAD1M6sGdUi0KRibch0MIQ5uW1i25CGKzD8fga+
TK9nMdGnfzVFB4JLJbcNcX84n4WDvjWxWJlivuJxNuxa57bm/VQwDQ7fHJVAnb22QthQXUJ7fyPP
IfackgZHI1cflPw3cOXNsIthXAm+T6ZpY6BF4dRKtOpS3Fsep1Rsi3Ki+T/RobfTAuom+u8FhsdS
A8mDtmUN/xziPrCJVedOprAUEMGlde3OEGZWHlxiigvDJCXd63WRO49PwwefIHtNW6rW3NsSUvhP
CK26nL38WUY3bg+xlrXyjkEw8b7wXIykEf0taZzeiBAH/R5YNNhP07yQMR0KoBt/6xZo1O2Gv/9Y
0JML6Z+C19SvgNy8xNNF24jMa3F6GavqXslUEhlmCz7lN781MrA+eZnIwcIbLa8fqTgQzb+SpzZC
mD2QPELQ1WSRtdX9E2KVW1dlIUYItREC9PFlXabh2BXZVqAj3oUiOhujOj2qYZbc0ZSIsR9wmwGB
SpMCC6DMypf2ziiXSc6NJwBEW2t9rEkjRqRQkY/3C0sD2l+DowYykfZ2/+CTeLKeKTSTI3nwCSZs
g3GOTqI0kv3g9TOxmXOBmBFni+yr3hiXH0Pd28aoWZWOm7G30Js6SBfpLUe7rMUqSZxxJBtvM62z
DPYcfkGL7htkNUY9t35Ht28fem6lhe/aQMmX2p1b6C+rbM4/eZIK81kaPbG2NlS3nvrNlnD84NXj
Kq6sn/+TfTcE8XKh0lq+5mUegwOR/RAaqDonJ0eVg0vP2WfC4Pmn7GOe5ty3omEZsv4MC0CKqQPQ
anLCi1X/RDbERsWhJpHfREGO4RN3TNkLg0GiCM4pjlo8+1INfQcCUEXZWgdnwjJthjwEedKDy8RN
b9ZQccRnfrcVPZreuxzMWccwmU8qtq21U5fB9Q8SZOUxjuhqwV7Rx7kixNVHpCXuB0x/byRBuMWr
d86MJlLEZ6WjdJcUeRGlVmOumASP8Z94R8rKD4j+8kOjB8UYz6SuC9pngTdCBKY7ZwWjoFgax9xa
dYM0hljlrD3BAjx36YTjeZcmfZkjdGOOQofxxcM+gXCzQmtp4oaOJFRlVQlCU5TjqpBShlvUaGvV
kZcZCMF7gPzRkArXmoFYFhLf9CRN0wV9rZ8zOAW7aVykVUt98Z9gAvIYVaNG833K6/P4r8G70DRJ
YkSxPIpVc4udWClGQiBqWQhO823OtX31aFYl9ZlT1hzGFVHq0d1bYz+IqLwtV9h1Rtvvd77y+nSD
doLqQcyY0GK5V7aXwHfYLyU8eSQ38wb/c2Km51GHMt+5TcnoEisZFTpI7G6JDnqZsq/p5YY4h3n3
ofXKUuzpjajxMknLW6cgJYzRZFzMNCjraE7GIvnzX3dMsGNForuLJ9yB3G2jdTWiwTmxM9090KZ9
6BBGaEimQ5ABbvF7Zr8dscro7D+UutBfuMGQsdRhc6TYnKHRw30VlGKSO9S4ZeD5fyR+iA5fvWwF
x4HYL/7TjNXzKKmXyc0YXZ+W/U0LuYkhhAxLBDgLJ6Pdxz0NLths2Qtybc8kITwuE7RYUq3CChqZ
1cP74R7ZpAJfPo802oDY30xjGEDWirRYsWaDcQPmrpsksN3ijIqewpUd1OGsOJVrJ75xOqWXQ/QE
pA28fTra2nSrRWfq2h27Nxn/bMbiI/ZU33y21wlFPmBv7cFiVOCXs/6A9+84Rwy4AMGCcddy9y1M
L0NORuZ20IiW5jY2XkSOlGkK7/a8h2056gd5TU2OHaxzMTINJVc7CJPNxL4rkpcMksVNDKGRDEsj
3+TsLUHm5UTkF9bwomjZK57htSrR6atCu/oyqjoC6DsHxwU0vmlYPm9RwtaxbbzPRu2S6MSuYGGf
5HNAtJ+SQQtj0tolIno6TQ58oVWkyHZjuyPNePn16Q6wZNeoig3JbX/qvkMCwzeEpDFEyjevb9Uj
oSlf5SkCmx/iCK4+MrRsyCtlZkkfEobL0qpGyLNG2opmW7rfXOyxOZSwHqJdL7PXHhX/J6jXEMUz
N6qDQhHvT85EtMla41N4+D1ex98F4FJhqOapDUYCAsxuQtb9xXX4bgZEdmvrhdqulSPUoYNtlNfZ
a1HY+vRGy/RKpMbuD//QNSwtZj5sUlO7C+MmeeA1/F9s1zQKXCJoQuGXkAfB7fTYRbsZbDANwr3E
/mzyC+Tv+IVwlRgWb7y73AHDq1CD/mvMhflmAU3dIsZuBgwVdQAmDIgj8HVx8pDXthX9ZfB67ZT1
077jT9KgTwLNYDejk8jDaSxwte5+y2F/JnMTHYbw6PAtWYd8YQowHGM37YDEcOQljlcDxCyOKlg5
HQUK9S34QRmhwyc6JnKbP3zosu7y7Zka638ACYNdiCvwGC2z1Tt4msGIW/g9FoMFkx4UUY25B1Zh
NAj2D/QNV4G8xlAZHncMc1BvQnzTOydoGqoZFNZ/lnBjaxGz+4egGQt9m4DnhHCdoW/MYCabK5KE
XY1+Zw0N7gersAzsh5Jy41bdGQhfZxfjZ3rx97SRxCJPcjkgU1cdwqla1DyYfmo3s14FrHuB89+o
8ZJbxbsF9Qx5gxffRHO/sogJLKT7r6eR+CJnYxRoQl2BQpETHNgXI1JUdJUiIsT4C4Wkb30StxWO
yew5hdZvdk6CRwaiHlG/I1eOIcdCNLHRCqRel7+K3yetn2+gx4sn4JXAoeqikxxKdKPRw/nlRmKF
owHwgRfIyN6XGkGoG99ZLe/Z9VkBE/GC5l5STOQ5t7JqqmW7xAJJWP+4bHYbNlYjaDoyfy8jl5D0
g/vYQA/AZzyg+onBrEJAtnexu1WRiJVzZtrXlaS+Uc348R3bpzeLrWcLHnVKkBVAzyWqQJHkYBj7
0FanzaU2ta4KgG3XIYVzlFQs3JfmM8AG1r4YecttQ0C81whOBvOs4elvmOJnN048b1tflNUFvdNi
ZyitRFBQFaFx8tznWF0HrvLpyN+vsFNxvjFWhL8XecwJLtsYSksRFbff08EozDD3F/mLk+c+BSal
Yex4vz3MeVLtOcEOUGVs1yV8sWj9409zl5Y5ftWWT8zVzUHEczJJxk/khEjpAX+8JLCfCaO4Iz9N
pSjmm7geeaOeoAZ4t1VHMxN4Izf36gVC2nbu5eck+S0Zy6aq/Nh4QsxdePqyJ8qgz7IQtYvQ991H
1tQwHCKnzyUZE7zqptNAr5tcf1+dFM76SuxobyinCRdQqiZwxbpysxdmtD0mk0mwzud7TlAx4SH5
Ilfn7am4z2EbmfN0OdMwaAo3CiMk6k9J7uFLQUa8bFH88XPchuYUT7/6ZMQpJHex8DWu1mtr2rsd
fccAVXMXxYuEtnLJRI+oTkh3S89WIp7JqPWxEBNaEaNi2rI5qsN+BXD0vfjzGciFMJNcUhjMgcqR
/yozIQU1UpR6qc3LogDbRPvsqayEFz1r4De48WvybgW6eR6iu4iH/df5P+RsLVmZ9Rwo47DVSdhH
31gF4lajnRGuHLDFQ8ta1HlTI/ZBhiZ5NM0Y3Np3J+3/ZGzC35Tux52qxJFMkQjSLVajonupj51R
yZWB38f2bNlnKD3Bjq1h3EwKQqMC1ybFGDqwWqmHiAs99gr/zIvaU4q2fCDHwqkk9nOtF2cFHzp8
IxwiCMugFHgHONnCTn2Yn3rIckIa2jEatcrqPE0/bpXRwrnqIzqO6EK0ezQDh+qWgeGUmQwgtkT0
5WOuqOjaYci75sGOyGrVDbJJckJXHC1CfYTeaQEPlu0CuA/63tZ+k60HvGSWEezehbhr2aX/InKE
5TkMmUN4k5JoAWMNv+n+I6PepJU6MWStp+/DMgPjMc5hZlmfqrOqhITCzMOXXWhCsmRssBG5JKKr
VRdXEqwwptdXogXMWtFgyG9WmKmhz+NitEWt3yVddFZLv6/3RXoD0sfNlvpDzEwL0SFJreZ+RFx8
YLFjhTpZ33kd2bUnwtXyNujnC0M9E0MI51G97B00POp/XZrR0SDWKMUa4tYY9BHqTJS4OTjbE1t8
yEmA0TWSVBCJsIvntZhfafuZIQFwymS1NPxVlgMmnz4QqCDJEKB4drQT1vKLJWCpTyQhQOEOqR/I
IIiRU9veVNTlcHoAJmcHNXJmf23QJQY9zC6rOXcDIJ/OuSJmHUEEBbekAyhr21p/Q68RNJHjk3My
tUwpcu0hLCkFRVum+6T+B5gIe1WfeNmWgAixldqKAqiwY+qDFnpt0V92YBRhs9Q5xk1/E5hjnKQo
/ee22iheoW0w3ND5oQj5MhB1iWPV43dPuD0hi/M3E2n4QWRWN5PgL3iaMLaWCrWMOuqaTbBQod5l
GJE122D8iCWxNgzzZe1PHCCu/LmZITeI1KGETRbor9ep7tWpkmZ+2uOr8jC6fLq2AgWEie/yCrXS
8Ga4RaSRQeAanvJSYMKa/VJ9yhzpsUJIz2tSXXFpdRRiXWBZx810IVMXh7n1X3DBd3upAyJsHlkc
Z6ob1JwtXzxQ5wm8r4kH45iJYS74fwQMm6pGuHt9MKn/KOz1T64m8v9b44BvTwAJwjLDT13tGwcx
Pewe5+ptLP6mqiT08HYWV3XhE8UXkCZ15rtG0vNMUy+7/LuJEkDoryNkYoUTbWISACkzJOPH/AdS
5X+XgyYX4GcbeSThI6N/IMCQQIyQyN1Kst10V6TdlI7F72Iq7YhkUZG8/4HqoP7re6/QRZ8X9Nf/
4DfXBPSwxxHzTauKY/emUkByQ6v2LLNosKHvz8dXBXlrwwEyV/AxCfBZXQd423EeVqv+hfbUX20m
Vu2VgkjICM4woqep5KVEpleXt3w7cc7y3a6vMzVnNIA/wAsVBoX7EvX9nk2BH33ngK6VPUowxYfB
EjmOwijkK5KVp+dcXw/NnvO8yKx4eBtZrBYQZRA9GRgUbQpdLm2UlZ74rXyRumFR8K1OX8kmUK+p
3UIEfLXOxiXmm3ODDZYbGjz54jaW77xUZ3gh6K76extXk/C8/1fa5GBw+Hr9uz9R/qRiig5JtRyl
brmEoGnA5Mr8yGRwGJM1XX7bt/OrQP89QgDVPE+bnMTX6mPU2SGJBWNpuUgVePOXc7uRmhiK+pZ8
wWRMXCfqXd9VB9UUwBS0c0UEbtqRU2RgDcf/0zyF88c+GcQkNUSI7aHx6PBwvaOIJ0oSuLL+xQao
deF9NGO75zye3pn88xZL+6hyXxtDnI63LsrZnSZqflcTQxVAmjOn0QPLyMwlFcu30ZaFCgCsybhB
pBLjFG51sDylgPHVGsY/NOKXfJUqcifqfOiDjcptNdtfMletVBxtuU/MvrJIWjxirQgRjxB1MeRf
LghHFTjLW1gHw/ORALuNktJXtmt1hmWtbYP0ZphfxICNFN6QoRKXqfIXNLal6LmHryKG5XArCV0T
EyN0Wk0lDBYjPgnPReSrF4dIALdxrK0PyRng1Mc23ok/+qfB5zTOGGi7wHAGnMaZJ1wVEMG0VMJ0
7FbT9ZgUGyQIE0SHsd5hINzYof8oDObicQYZzyTvq6lLitD3Mqs5Mcqd8mZQ1FDaQnYWjMvf+hou
D2wTVP4P5hpRvzGr40JPTb56WDHoMhb8mDIYm9bwyzXNZH42GL22f5wDHeTLgtfo8hKrMGFmo6Jq
dKPFFe+I/ugEj6uCRHXNYKOmN+VGXSyoDeMDNcWgUpJE4fEgHP/j+xJlwas/Vr2ZrZSsaDsIZ3Z8
7WLQN74A1oqCGVVvsBEoDz7W18f/wdB/eBVp138Iglo0ECLbiNf5ywuM5QZ+/lO8rgEz8c1VAykv
KS2P/USvUJY4iR1tJD0+j+aypavKVL7zSFeZBsQFgfbnH5FJz07phwGBCl8J23wFw8ejxqdK71wy
tcvF+HJLKVlJM9sCy9SRAkMbTzP5is2vlbjcpaUR6s6+WV4iHiMx/5oLL2DXvoqZDMt7Wv2HsEFu
QHYw71/NX2ebjTJ6swxCDMvVdQnmkFznsjjDfF1vMNjpWJGD0upTmxLliRTSvw7Ibv3r4QLZnWU+
KwFZhOqlfq/lyjJpgJbcMXp5WhHCdG4gv4nNhrpqtE5Wg2UY1ewiJNlRDos8rqRa5IdItEnTF9c9
P3N2QPnyrZYtaVwY0ZBAVzxatC8V4ppOM2n16smumksDfTkhJNKvkDSb7BrXvsZ/AY3pOHecdNzT
88MeHNfnrWY8p5IBxvpUJ7KOqEVcx89dPFHUS9ACNEriMkNqeRhlTCkyMjlhXriKeMayzy78ElO2
HQ45fZDwdcju9Q5AMaGKe0H4XRh5IWkKXvb72oZ7iXN+kVC0pp2sV6c5PuBwkQ21eGp1O9qm0wgA
UDKjU+I1Y2Bzu0Ylo+7gP7TIvIEi2slodnGSSQx5JOBCh9h5jaH4t/0qLis69kTAn/NRgEODbQWx
oi5p8PMCGSf0TtLAJHy+sTgmnyu5zWqG6hrOp6M1dSXkJfxS8EdI9bX1bMOkJMLtdDxbjgL59R3F
5RIL1pPS1hsSy8tHPtpcOmL35VubnupQRQ3oG1/74tbjzNfviV4eaKvTIHUKiueLBqEqaufd3t09
eUJ4MIWyFujbJE0LohayPV4C0wa/j0v3OJOigV5Y8ygXGMCFPRKbrb288YC9DKjvMu2/hyxPYPFW
MXYAIid+6QIcLvKQPLLjs9b1uoqizpIDaJrQBdxep7Q2aSS0HMJKwjKAsND9WFr9xcZ178PnRNqF
AARmJjGvHCJAXKZDNy/oq9aBAfTudUj4jdG2xrsohUUzB8CyB5LI2m3GqfOuygToSZaqBk8V5UsZ
rkNtksBSjKQ43R2AD5HHfp01cy/z/VyzFRrmHIq8h8cRZreUai6B23/nXW0linAKQC65CfCPw3MQ
HlBuCP4myMeFFmNQKGet+wOuSYgQc6Qv1bFWxy2yueLuZ6ugWoNtC0KPevFNzSW9kSa8Rc9WsdG6
XOnWmHyFWDUy+ZiUzyaBf9xOQaVm8XXS9otAgWYmHMHBriuh1eOZIiohkey+ac/vuIUSjFLoAsJ0
5QEAtzy9Gjmm2xp3L7PZRIgzCOwTRlLJqSy+0SUsknmhwPOiuEb81sc/vtNYmLIdUcsDAdVbrryB
ecBAZ+ZC4iE33N+QUB9B+Rkxsm1g0piWWMvGXdqF26qcmKJbWPVs4UtEjYRZdvx52S5TI4BSq2i0
5c4cb2hX0f7ORnzWyjg4/KmzwB8EUNigDXuZGiSeFvdQ31NXaTxvl40GMihH7X3ffmo8U9Xfthz/
BQhZ9Xvg6VrNAMv7SGfBi/UzHr9nfciYB1sxAlaPxSrOvpBzaR5JooNp5vaPgKftkr0zXHPQMHLf
J050xSqNzUbIMyHwW6s7+IVVLb0KbkX9bQDIr+Mtrcxi9r4w9xO5xqdH0eo3OSrhcIrihAxk20zW
0afMxv8Hu0o/yGddNZrPEGE7dLhQsrV9W9panJ6jbHuv6V0Q8hwSRonxg4Hur7wmO+o14j8ISFLI
yuGsYg1Ykj9TknttY1g/UNHVs388aGgGZyiplwT5fZ0R25v2c21zvEtMYALRpaHa4VTZK7Y0C0rh
xeo3E0VaJAAocGYol89bs00A3BA6SuFOicrKdmFu+iFkmRzyjTI7xeK1mVDJJgkcUSikteiBhdWn
Fb12WbTh1oiOzYSoN4oabFNxGTU9HInMjSI4mTb9o58LughNQ3jMJxmAtNhW0zsJfXBMdcww/ULJ
nsQJ34LI2VXR/PhFwAuHoHRnnSCI4EaeyHH0FLlWtWASgv4MtU4lGRjWczWi/qBIS8A3Nwn0MCZm
I8MvJ6xg0S6YhA4vFZ7HcWlo+/T3c0ljbyKbeDQYpuqNLRDwYv8rSqU7xDZHFULQ9Wkst4Qj8Dvs
vtFlw29JT9L0i3eBuFHLWLjGVFmjIK5tKeRN6AgfXrq3aHBhyWoLTkiWT5xGwbAVbvaNT4YSpkkg
8IEnQcBdgCR20r9ykGqc5ayxcKJXYr7ZtHPoCpQ3rbabmaD0tHDIb5Gnx42yHUrS1GvW9sjRVJ8T
QoQrDFsKquWvl6Yen2Re7Dz09DjRubOV5jnIpZJnTTgQ6aAzubZORcnXGcpvFNcMwmjyJW/Yk+5b
LhZuFYD1z/Q1TOFJH7ofysbaJlUFVmZ5nP5Vpk2cPQIPvrEvJCS/+UZUsJf1biN3iia4KAvJJCTI
Fme43rV+wYvtvGNDW+skpFHIeWQbHpsJjjNbyTjM1YEuyKmh/SgLZ2VLo4KpBZEJMgwJCpMRROC0
quqmZ9RZCjScoWMogu4Q8gBi2ZyvZkyttFLvcRjMg50gbcUnjUeW45MOoR3cjWs+I7j1txUiyVNq
7Ks7apTD+tvzPwWRs5aRbpC0Sd5DduD260GMyx1PLw4qPqYbOG2DMx/3H6Kcqi7ThxJaZRfmNB0W
VB9qSO4HagnFq/Xf2geE2kUtqAtNWe8PWn2bTz3JLDgv1P9FrCGQAb+gS2hF+wDJ14AUbU6/VdaS
4HZS9klR3ZYNmACfVTVzt08L/clGYHkc50CxKRag2kSmPneqa1lAJGak20OL4tOBIETTJyCg4NTb
z4qfX4tOeXgLwg6GzW8w7DZx4oEyB+1ZyAcjrGG5kucPhywWRu1Jh1a9HiVo5YyVnaQ+VFPvB7DZ
T59d87DzEV1uF3ltVnn7LToeGXoQH70zFXhT2w+FuaGAd/Sgo1ECvc7iz0VbNI5U3qM54+1A3m/k
W4rWuAr/8v2+JVmREb+1Jqper3LEMghumwJ/owGhT7v0kOAYBmy9/hyd+ovUrN4t3+p5lu67lMYs
Jm773BYbYnltyW5sitw25mGPObPcwXWoHXfbwXZUBt6c7u0efoaxkhDq3n86uhAorvjTH3VJTfh0
g4ToWWiv7YP9DKJvl/MqVKF8JhJ5qPUaISCH472vvCewkH30sWFhVBQCfj8j/R0jO4k8+2QfBsqd
qO1ZfaXlsj2DhFG7UnTQ8NMJxT8dITBFec8LpwkQwFv6QPKqaFmiabZMUDo0oNqxQ9gVsNmflJP7
x1uojVUJs0qHb5mMs/7seCdc5paUw/BFxnMasul5QUS3rsUZ5K9+W7DLY5XrxvnCKpsdStFuvCby
6m+3XH/CMKL6zYiwvZMrFqlMLqYcuK2C9IDGgKDLzgj3LTqWLAHRfOqKMA8C796rTFV9GvbN+ut/
lNkdldZ0N0hpyzRQh7Gttj8PTkmT6Lzo6BzljVTHWuRD1/UwkzTxaUtcB2z/DNsF6b7d3+3IAF+C
cF1yLpLwXodYPsmko1Ru91IoBX4B3I/zeRWu12out7zg+V1reS14Hfu9uS+6LQNIZZqIk2mA34qd
CCweQXzw/8kfQrWGLI3bwPguSnn1AWvduqM/nMhpppVeWia2q2ggsJMfMK8LFNS8o9gJ/EGqj/Sg
jsrV7IzMYaCyc0LbNoANbp+C39kVI804olZEDigHBsB2KjhWJZVpFt3Y4FpexAl9mE+Qamr+sGu2
H/SUPjvbBJKpqoTtO2RrDFoODHSxZRYWZHjTCnAW0D2qVGNKMIDS/N6U9BhEgJM+C9oaQjJQEBll
1MK9mkazE7Xe6SbnVVDMwtaelXrrPQqzBHuWFBAfd9gawLS/IwQOTgAe/wXKXtzWm9UboPC1x/7z
VGoIKAuKEPvJsGanO6gV5yQOpZFriFWygnI0ndJVV0kRQPxXYRFmiUeszYuXKBITILQF7ozk8jQB
QvwzL9xtlwFD1s+oKZiQrruuXe/l4ss6jARJ5qgtdOpwMgBAkrg363gK7lNX51ErgjfCf+KY1oXb
Y35uIoloZ4Eg4aOvaSYTch7uy2JSm/iMEQPiCwwppT+FFJDZaxke6vei9zBlQJAsjtJv1Y81Wli1
GxVGdkuOhOH/rYc0HR0UWqPHeETGWJzV6f34yhzKBX1toR7rYzUcKWAkZUH+cWN7tMI4/tLlNZAQ
cvYPqmKeM3XS1WQhdKCMlTmgIOCneRE1c5nN92qGPFofCaR13EuwlK0JYtec/kpBOoSx+/iFA35k
C6luTX6Pyz6zfakvGIDlZwyyBOS1wFPk+I0eBaUA+0P3KazN+pYKYOaxNNlcH46mEY9Pc/hT/zm5
sQFYTGt9wJWlCpdiboDxWvQKh1kKptlcnsp3iGCwzYhOBfCDl0qysvwO7peAuouDG3o3zi7PB6SU
Fv2L+zMSsUITO/qQSiu+xpi6WEhKovay34yZkFiN5T2MZRZhuM8bo1JSBMo+Ix8JkeH5uDlu8X1N
ox45yJd+B2895aDm7nf+q2fr0ZlRCmT6pzIjYqtNvCzfjWstanlC2QRdKw39SBmDZVmPfsuMEnIR
0MbYjNNYS47nF3iwoV4jRjQ6jZCyjWVQr5XnOzm/wIPZfixnIzPq3nI7SUKazzDd8AORu6B6zeFR
EVIEwIdtrLHfMBtpCDqlaM3yP/g1lh/fxB+EikrSZ9sAmEGUR3C6OwDHTW1OuvIiALYSTHFsjFNc
iITN2vwATku34Iix+HddoojYNKX1lHzRtYXp6fM/vfEuZrDIHlJX91xotObg48S82nCLJJw2hrXd
i5BmUe4yMRtu+9Fbj8b/o0W4QwKXDjle5UjH2wPqpgK6Hs3p1ScWyQMNFL+zDFQIaOctfHaMKQgc
dbBtSGcSlJn5ldQj3xwB5VUHWekWLX25IfFqdqgHW7KeOEW0+HfFWUvM+1OtYezusR5hX86RPF0s
bA8dxQcsExste3skYybEMDHdwETBhbKk12Zetw87v7vSJZHM8NkL6xc94CRjmNETaubRdhLd2/5O
H6QoiYBEnroK5YdRjrDLzHhCzexUpfJte8z+74WQGBjTbISk4BA3PXpv86ee7CFX5M1cYiAGyXPg
kRUAFHgpihQ+F2cm1ztotnMTNwR+LIJRRQl+S1R8QTSZrxzPtc8lA9BwkDX7i3oqF85Wunj4SVAd
2Q7TuMkVwWHOZsrUb7kDjYprYppEF4+zpTQgv61PVFwI1eOccBnFXTMC6ukKeoRq/uW1HLcocERF
Xh0TPoEZeGzwaZmieLCZ+aixrI3FmMxGi/B4+dYhU/Sb+p74AL2wLUffEyKK9eQ9QZLoraBDvb36
Uk9AZtAYuH8FtludwBYV2gQ1O6ZhX8COT0AxRFUUq6VG5Lx9VzXvKDIj5DcmFR2ijI6umaq8dGNJ
z6qh7+hX6lSH5rjNcR2H2VslaYtawgnFTerhDkJ3rtKqR3yrr2MslYFmrNP23yJMTgRjzU3FZnb8
qmG2I7jQB7YutrEB2BjrnSnFfQGa7PLHU0IKIZPfXp3KO9p/AoD5ybxLe1TbLT0A6WbfoXBlzdJ/
M8S1ZYSe4BzIdJafab2gGnOof3iBubuQsNNxbFVmU/v3Vm+Tgl+c+daBUel0Ay0Mcqau71la3G5n
maHzyuNCIfqhfWt54ztVKLgIgkYVWFTBeqao9DrmSr23P8Z80b865o85eiAPUOVF7ZhyjJ+PS1ND
COKY15QZXJNqfBaXSvDAxhYu+GafkNGQEKDMqyaCM1GhV1iT0B9TICYAUvAR2CGgvykicgMDgelV
/d15zxar+J76pP+XI0pHW7L+VX3bxmvP6aNGAsunpgxpwK0aRm6xS/Xl6bZJlr7Xu6jorg3mwzyS
8sbPS9OHv2E53g91NOUyNZ3+FLRKQNl+Lc0liRnOjTM8/RLEEw0K9Fzz4IjNhsv1aOdP12QGct+7
C3QnLi0oS68LuINhscfcjh6BmCtb6gqIMadRTJlVyfZASRa+0DV/LP/ANHixzIeYfvJvwAMAk/VY
bjLdGFOkAdvD/xNICJXTsRuFyWMLEuAAzZmjTmsJ/6r+ghCiIDpZtMhWhgf1hZZtPRqWgkcmDBJw
9gbV70dPMfjVnYSnQONXhU9kf7+9AuDIHjyC30yu/+71TxjeoRmBq/Dx1kw41tfexVv8eUR3ergD
hup+nGWAg0i8P6FGraJGRkKNYNbtzQITXF+kKzs4ThA/S+XK1QiAPohrMdxUn2mk/hoWpQoxyVxB
hx3dZJA27uQ+r8MzDYt962TEiPC2xcT0O6uh/Cv0hgwK5JQd+Kzaj/HhqfwE/KINnaJ9UI5HtFlD
oZPxK+PNN3BEbRt5/hgVUmA6Hh09ERjnfu6fQFwfgzCEtxuC/c3R//fu9lvlrrE/zvr/kKvT46/l
LS77sS5/hoIdPbDXDErEGfYqeSjI3N3Dztl5pCZfjjphI4UgtFWSYUwTdiA4ZAxdrUd5a1RmQ3mo
37LdM7Qz4wPuNMj29igXCI/eFUJqXWuIEXk2MxJTM+l/cm09hyEO7I7nIDaDIjkomJ4BratthHi7
Dd8cUftEAamd+QM4y3meVdjTh6At1IC5KgTZY71+V6L7mD0VgUsWXBnHek0JJ7bNZf9Ry99rJrzl
RGv2tkt5ZJHPL8uOIj4ybFpOz1bTpDcENHKz6PMnUU1w2h/MP37xu2jDeG5jE1k/Kv71KgfQpDKh
TuyY5AKbuNtcDQU8GYieR2wEZx9m9ia8sPEc9tfyH5jkDfjcX+2wQLiEwt3YUbYypH6Gxo4Ul7v4
i8CayuQ7U1t5N4oCRYP+Sb+qNPUUbXb3KynC0SiFQZD71GIFzbxYiqklW5rlIi62kkumUT1PZes/
NiZ9fnhw4xh1JsfQgc9QnxB4kdwoCzEF1sRsrUQRN1ybwuE3xZ5ij07xN6RSxlDdQUVDnDw/CgZh
yBTdIwxrP6iqqmlOkYNRThChZupzmvJJcHf26zu5mOH/JTVY35ydY58pB66anPEWxzHP6QP/Nxe+
DstOQVpNBoCWBapFP4JJsqJMEqAwDBy1qaQE7QvzA+F5Q/uaY/V2sL5qB7Gq3hxY28lvFfwgfxkB
MeQJIdysac7dKPtTfB4AjPZYP5d8XbQg2MGWz47lGRARJDsMkbR/r9T3x+9F6H4505dk6cGnpTBe
MTzqkLOKeoMkB+AKdkIMhUnZQR7TXOxhVyrwwsia6heBVxZN5AEpfhtfvIXwt94L+Xdczillawmi
iHbgu9yXSHDZ7C2tvo6Gl2V8lQUDjl8yI9xdcPp6n//6wNQFrKH0pyMPLlefiv8eIvOyBkHAcoj8
nkaQbVcP/CfAyMiJ5zujyOI/Br1ycug8xQfhx5EIlIWxHk+tm6amgox8WDaPBcJHb3Y9MbQFDHeZ
FiN7JbidCVO5eVdNYs8ApSaoErECLCNLDKBjTlecno3/5/3qUT7Ot3R7yEecvHdtOGAE5sG+ttwD
5kXGWZYOsp/ule2xIveJF1FfOUB3pofYwIqcMCqYrgSCYm2C3xpRVkiAgQjpQcBq7Uws2s9MyyxO
AfUu2+s634/FBBO1jWHq+4cEjwFeZfuDjWvN0IWHXeNvrzjV/4X+3be91gAfQ9ttNCyuLpmf0eHU
Bp6FuzB6bheJUgejR/RndZGtl6M+bpgU2JnWzzHOf1tV2FSKZsD/oDuYjFDcEjSF0zXxTYgzB1cC
Z3/SEL2evdBnnBo7zcb+Ag5oT3M5dxGlNFM7Seq+Eg2SeFJs4snXQO1odAt8+iUg2l9HgM6LigJZ
F9opoLqecqYdJfHgr4yXggpuleQVbzMXR3X8cO+qbD0aY9qPAW5aLEo8itEw5fJud2kaH15asbCC
THSMfJYg4Hkcb/iKPMm/goDh7z9wNjvQkq6jZYaKZCO9uA2AJ1RR5/AZM7Hmgxp0RL/sbiTtXjfn
rFLUtO5hd/Wp8sHK90O3jCAWCJXW8aet0LPtcLq+f6fzJTo0D6SvPxQvyYLsWfKqlQ+7UvjVcbJu
CSMEO9LfjCdpvxvhMpaOp+cYimS/P+QfcG6CASxlMEd9CnRzsyT0cQzVXcyoe2VG0aJzTZe/ANpU
IMDZpz0RRML7FNIGKYmh4RHAoYqAtldN4lPOEHmA3IB1XI5oYBbkgTiUO1E0FWpbCUK1y9oOpDc1
Zx7tTUT1Q4Ucrj+2MT5ArtDdeT4/vQhqS3/IercZxsZVyXphlGQRdb89fwubj3lAllqDILLtjvCS
G0snbRMa1akb0acvYWCMdISCdiBqmQHb/W31cbpm7BRzY8id+C/EOt4yd39tT7fDT3KaRq5pSuK2
G+er7j1wqsb3Xg3ZnYPxVJK6TGo36CZBjhJ8UHbG39+18CsCOvozZsy84jqtGik2iRkW4qLwKL2d
BhZi2EFz1ImLUDclt+4666O/3ZHArTHEIo0DeYx4h2bAniKbDR5ylKjxQIeSMPgOmDiOssIC6dqW
Ni6O7XzwXuuKnVc9rKiBMofrepGTUMjnIzzLQQ5o6jIazPJFGmetXlciE+VS/0C2Z0NO2ctUaQ1F
rKJGS5dApSQgHA3+bjX/kBZjRbby60xCu2S4jXYiJqNb5nyyocSipqFJTG0o/l0ZdAAwvojf/txf
L1Bm9zLP5AWip0kl6SJXdZfy98BTSWCrLKctV/AIABewa6cg6p8xey2JZ/F589uY2JYuVYySBKpU
WK6aBRIGopFGGr/oNz2s4nY1rWvRUaHjZb5MUFfoc4z73VnWyn1o768XJsrWn0Pwv5HDDfdY8LZo
/uSdkaLHCA6Ijl6w8C5uKtiipnPl8donZLigEF4kdrSO9jBNyX2HErFJNCNzq4cOwOn4Iqj6MUJp
fYKRp1XohrAqpZmND1E8MWoCrSNZPmBrRiY5CPdG9on4blTl2j2VNtWqTe7omySP9tkGHbp5c1S8
jgJcKBFYR1EQgxumJHiVCF/y3Q3Y7p+X+TqL9s5ScU15ts+Tj5SBS8G4mqiMqe4azx3iH9tdKz1S
FB8MC/hSJmNeZRQqbYpO2L4VK2mQpqnS8arLz0HZBVMKoc4kOZ0F86082NfAw8zuCGfdUj7r2C8i
PPRL7cLImo5XZg+IUxXT6pNdpbHSY3p3DzA6Yo9XYNeJUwQYQBGGA8EVCrHUTw+D0mpA2qz++E5U
JF4gpGLA5VJqbIyWoSMrOAHH5u16HiMGlIHcRqCEcW+snjSnfQPs/Ro62+soDl1WEKNI6V7QGsJr
aHsWsOWiddcODjP60nqMSg60n6unpfsrDQgaBXCQF8H3lRrdCDDAiZeIYVSl86T51Fv/n6WWqg+d
hARaq8sYei0ubo4xNjPNDa2xQkVXY1UjLNpEFh8kJUHQdc6vxbY1KpT7S3wGkL00j1vn7zqv4Dup
7XWalhbDMD4RKOMfrn1r4+FdJdg8mbdZIi6+nB9fXwzefMAMBwNY1XoqqXTEjEdOv3zpP1CmrTlQ
smR+UOVy1vDX1gWV/qTWw0AeXBehhIe75nGbrAfOaYVHuah2CMza48g4pSdDTsoHax0KqV5p0qvk
ohxssiIYt3a3nW6eCplM7mLQRvrnNnPfNXbBwASZcFnX+A7RCQufFzKLP3F8DvLTY2oqevwnOe5x
LxmAljnxssKeA1AyRQSplrM5dTGEbNLKuUW0nclOfeDiSuHA1t1zu9Wx+n14s49MeHOaT04xfc4N
ul8dvK1JUuq9FapX54aoL6r4fwr9MiZDJEZ5iH5jWmOhPHWvubJxqUTUnLk5Otr4Z0cMusI7+CBu
6xiEG40kdi8disADmYOMB5AxTtuSW2GXt+9ojzKzOr4r9TYVgmduWdBSuHKvJwOIq7979FRQau+l
w4UoTUKMnsoyg4ywUNtQboB5MQEVcr45847X6d0mpYNEQJgXkZlAHHRr+sXQT8F0cf+b6orzmyA1
LOkDqYwClEiQy3i5NdF+ovdcKdYwJxd7DJ/+zKQ6iBzkYvq1Tigr9radSLgJkhjdnku0IOJuyvtC
dv92XgowFVinzIyf63MKFtY96zQSUzrNvxiO91ZIfDuiXmDEQwpgpvHm53cGhxVj49ONB7nNVyOJ
2EUengCISRPCQPcZJAcBvpEnisIlNhBhy4LqAWXLEumUIjzDO5rNyMhApLgThMCfkfufUyP5ncCf
UAKNMpAjnRNl+cdvYxzY8lNpsGv4kyEN4eY7vrkDhTrzut9ClrMiUCua/Ry1NEav8YBrNtZ4q3fZ
sngmFmgiPo/eLEQ7p8XqU0Qtxju8xaLCT+PXmCKn26uJETzFwDbEFKNAnrc847wxT/VoJxWLDMk7
LAViVULzzTlcih9qEXNbUXpmvLnovz7p8MXrzen9GCdyDrVx9ODPjMLQ+sRjwEW8X4uLMkdVLILJ
IyMEm2axXxFAr7RWCUxrRuF5Am8u8PSzHOf1JZ3+U0wxl8NKuic69FdB74ekq5WRV/IqhchpqgCp
g5+hcROseeDU7SS92zK4kzJpSlKTSa38tTIBf3Xvi3zrfv+ezlfcQBw8uflMql7z/b2dOinmlybx
RGOOlCtgoCU7CpXfU/OKTtTlQw52k1/cskReg7z1Yqv/NZee0GJwfLzI5xjcnQ7mjWRp1PDRXwOT
EnBmnKyiEC/54ROqVsmah4kzGBjRMl8Oz+iblH1gJCUGyx4pWgkCLd4NVkW0bMEu5Uzv9fXIjaRa
VuSbWfTxOYvnWgnfHT90Uemelxkh7S/39VG65A1tRLlNG+F1MfDOM+Yoa7Td5zhExo+H3P8bXX5R
H4xtXg2n9Z95mKZ5opE0yqiSxT2y8PEuLSXyhmjf1E4l1FgB5SKl6eglsUuRNRNR/DMhlspOC8L+
Gaxq7wrVvh/9jf3YObMmtmZ38rw1Y5rndvE+6642UZ333sexLMxPuhnQvKg4S4xJXnkbqmFbeVJL
/R0YqazNVDzkHAJ31E2H4miPHCSI5lgkFERjYW0s/lYX6u2x8Q+iZbITh877+RiJ5kAxlb8Zzx3d
iSPVCUlpqP9tzIx2Vo3ik+eOvR7V4HxFGMXL0baZG/PZHO71HrUFCoStynST/YSQNtNB4mjqHiqH
pvEDtYNj3GohuPC0SrGBP0yKxSYFXc3qojMWkjf/jokwv8I54yUMI8VFNv7LCLKtbsGGF1vuGilF
FLqcGsc8aWvYBerGeP0788TSeKhHAYR5bNUm+er/Tk62TnniKUMg6C8gu+zveyDoa+1hHXrf4mpQ
9+KhgB43w6jn/jBrkqPHTuLD7AS1Cfw3/ju3YNuE0RdbRJhsaOXkUDQ56isaWGoFxDqYsc8yDlYO
gjD6988SqsO81Np0eH7k/ebGkJh7gML1AOLguYlt2PiVSPq6hiCDvE8z8BI6LkrCM0fGo1v2sV09
4fLJ6Abc+wFKPzbXwridWjwTjEaEtVJLBzl/wyYKGVeTXv+e+qrniovdoxBjv05jb0hCispLRCxi
6TUJkcG1SD2L+cubUJtGqIXQxCr9dttEPdMaatLopLAtZz3mFVFL6BDK/VpIX0CZwOIIVmO8nq5q
Ntd/qQzDf987SX9KWuiSZFwp4R74sfxgPU2M0iXpwIi/mQCPe+9RlSjGLYN4DBnEeLEW2zSyJPQm
gZzXa0hYpSfcxRljS0tG2bMKgg2NR6a87SsBH/b/ZRVgFiPYSGI6fkCdcTxF760pItkA4Aa6TbC5
UClm1ziO5UFpdoE5nhTvL6WiZcxXpRoFVhF1NolzIJOBIV76opQlVCg9wnR7Hm0/+72LGPIsNH+t
X+TEjQBRqJ2MRwi4lTYogKw1mUXGp7qJHzFdA0Sl8KJUHOSCHGKQ/3+kgvQZZLtaEwI5mwsW1Scw
/GiKPl7MO64b6/42x26F+qatTjrcWnoZSSD60RdY7bQGvhOLc7UqdQMYiZM15xQxEuVl6jXxfL3y
oXJXkGS9vr/nrQBopuBrUGU7j7+dGcBdSHl6DoyFmS5iKKhTM4iNKiQ++Pd2D8f3oBKVVMcKvFTW
dhfvEJztJcQe3R1uH3Yca6CDF6X6Kur8OQ4ctiO6TvjLf8tHBW2fGSXVcYGml4Xz4Y259B1aMUAP
rJpfrMTkG4xyeH3+xg1aFaGhTw6UPxtyyzE9S+B0d6MujKiorD3/yuTxb4eY/1XljpyslrakgmOV
JrQMpcmPwALKZrAdns58pLfa1JrYX3eQdSBwRuVY/ghvGDLuyElO6aHnZ5b6AjFx9CGw3SOKfdN1
vkkzkaeDzE26cJvmkwp3mGt/NGcgBFM90tLUZIDwpZ6z3o/XQtriY7uqQhUenIT5UQ2ycVVZkYTl
/pLHgFRIpuShiCyL64AC+cx5Nzer20ulhsdGsmChtE+grffYyeb2yIU8dsEiC0vD8/KaHXihnziW
pifkeDrjsxfb5gN7KkiL0kDkdKsC4FLIqmBqny1Vc5XMrGFvtk6FJ3FJBn8HNBs02LJSH3hSgQFe
TfIJeZIjpeZaY/A29Z/cxta7uKGt0R4WDJ7v6E5gX75XAlvXe9xQ0Y/2XIF5GpUmvgRcFR9kYaKs
xqHIlYAl+0yZUW2nCHUIX94JljV674miQcnCLRPFOneVDIwF+BAH0N74wfksBp85DV5UMGzlQplm
mS7pTmZxgB9ix/IqzXP5vPsXPMSTsHAV+6HW76IXlilw8wtgHJabqZspqd+mhzUQHUhl+1Za76UO
+UgveWhKEKvGRUDTJl9Wn0XUy4o+5pODTO6At3X/81udGeHZn00eA5WyCU3yCP4bD6wG9Lp6ovwV
zNHAY8pax0l9JwrWH35ck4lyDUZTwkwJbCXm4yu4BkS8jrk6dcMM4CH1MjjVSrSYd8mF7OsNghO3
s2Ow3ku9Py6e81XIWprakqVgWMQ4Xe4Dhvwl70cwlWzup5eMRrYqFeKKLfuDfvLPPHKkXHBkHqTm
+JV6DSGILHwvm4YUTZH5QJyHO4/yqu1smZqy0EjMJoV/kyT7groKK0YnkF+m84o71f4M+VGf7pX4
SzghFSX+NoY+YqyLPk50KnpZB5vLs+Txiw9k/YnxFcotHFHABI7WmKSVvyb+6qhRRPByZ29jp1+R
a+TjQjAr/o2rQlbQxlR2SkpnTabJDaXxW+TX97l8PBmFRut2lXF8PkqqxI5YjDwg/ojiDOQket5Y
XoHTpq7UdC0QZkbrQnLhmJZ1Cav/bJfRfb3LTBIy2CfQ7RhYe1huRoXN9TCcjpQFuy3Uji5ftHHK
CQXqPpMfcwKhTXnj//ETpudGEuM6fPyXDkHfTecymEjpZuom1sqEBoVSm8QdMSc52dL8CsTa7wMa
l1mbHTRGrjY47QR4/5U3c1dzWE3983blAa+jrJw0qg/r4kcHS499CxkDbP7nAz5g959HiQC3PwKe
Lw2w7ZZHog6mNhjZSAzD+qpWeTdLEy42P1yQy0OwB0cpeQfC1A9cBLLyoMWqbyIGfVHnbd8QfyE5
LTMIXTCs+RbFmUNle30hYTDTH4KELIQHWPdLHMgFoDm+m3QJuzEj+IIPNaUFqh36URHcae9BV8lE
ERR/sDguwbAc8pUaGZcWP7MbfvjzK8AZz2SnqL4oQZtK9j7kgd9ZKuiJJUYMD++8p39ekyplBhLI
zB4jkQee7b+YjCcWblJ/jA7h9GnaGJkNkgAQyoAnDB1CeO5kzWECgfwhLs1x4dVZqTcy/Ff+ymof
VnPekqR8WZAsQcLhqNMt2lXcjfAz51DR+OECa5XB4ZhPr7zjmRT+xQLIMGgl5rSVSj96B2EeZGW1
SRgpfgxc0vuBa9LijZEWTknDhVt7RHzGahheoe3PnkoAclRJ4zPcldLpBCHYwjRQn8YpmEx2eonW
O1RfOhjf2bH23b4ol/iYFgJwRxCPZmLZTNIVX45KNn71ApHniEczw/On8vd7HbqbjjjW3aqv1vuf
qrtGVAnK4ZrP7A29hTGx7l6qT54Sf39sK3/2rwiMEE4TrBLJQVp+gWW1T+l63B1YZ87JBn8OeLa8
q4iLZZzEjwM32rJXaZgTxV3SmnKSYGFA/ha2Q/r169ulkGBUXllpl9wjNXGeDEDkp4X0DxaPT4b9
12BsvRnKC4mJbps3o+8HlCEvlMj/UjcpIEdsxJxKB/gb+JFlCWPpfJLsO0k00D+DjLsmGMl3LMAj
U3YWnPTJIgcV/bK3+pfuB95qmaQB4CNlMAllR1FKmdWuBVM2WxMnzjcT7XA/TA7z6La8FbgYCwNJ
MuyJY9v4PuRF/L3v4G8ZJjDE8GljjUELm6oFGdqoRyuTgCSbwAOz6Si6HXGe5d/hsxzGFPCC+Fqv
ZTQ8LtoxqgtRgjGwg1dIxLDip4IDkTNq2holPlM6tl15FzRXQjEnxsWnvnxA+65wGc/NUgcpp9mz
lKnZCihHlnKYSwP/XOI7+/BQrdB2C4gz95RlrPQ8JYHUb3jXiQ2C/gByVmMAG3xMxf3k4tMjATF+
ZfisIPtGIj1iw22UkwEj88cRUBTXkw7ZW5wROqwrlFx7bY2+wIaTjH2/uplxDFyt6PVlvx2vvboG
wiuIr1KidQHzSSoWGE51BF+hgjxwtY/XJkgEOUXKVSJ+yvNKU9LQRJWkpg2VhuyY2YFs10XCIuBE
28exGS0cbCXWM6w4nrrwnNSj4seANYCOfGf/CGY7+khZWmAcBcsxr/SFasGXeiVom3x5Bj9rCteX
H95yy3KSShy9bteCcQ6GrmPxtaipaMh3IEnJaImORGUZVjTGyyEnyvxfd8890NPBgkJsZ5c+8WtW
I7dplZtkJj4sJvV1eQpPzz5X4fAZ+vGJFnBXe2+S0P8VlAhw4D23c8N1hzXKK7U/Q7Vi2NGzX/nV
IMdokmD2/sympSV/qxEQoxic/YDnDdLnSSO2JCAaepjsKaiU2+fDrelnSyO91mmpnUgMAX+QGnqW
Qg90FF9UayjsvcbpgsEEQonIIIuDkCV5cBBuL9MaFeuurwQ01ho4CuG1WNuPWYayL1PPQp35oxPk
cTKVd10cOjD9tZrKx1pib25NmtnOcozjS/yC5bz0BTAmll9aBp/kzxktmSaThftGAKkSHzmRAR9b
zHS5BvIIWVZP8hb8frgqYXrxG8PWMFXqWKAugXW1xzEujOJEFmakctN9R9BPWG8HCyhqVBA0y3bN
bShY+TJa0B6YfHiButYznQdlWjgp400a30H8Cc4huM8xSfbpdLnfWrKOsfES2bPo/7x0jx6llOxo
Aymkg+9mPKXPeDWaYl8xAaO9reWud7p//eIBoHTQgXYsTjbApb5iq7gcsRAwVEIn2o5WlJ+L21lU
b+h45PALUHe1kvQ+muX+qy5FkUQQ21Qdb0xODXBBV+OzHN3z4C9gUrDbgYrYvM4TQLaUwLuMyKJi
YR0698KEfuAR1JcyEwPLvFsVY73fd/pVMS8jk5H/c5T3mLum7Vb7xDxTf+986nt9sEUfVsGSo+0i
2kY5iQrTtGjYEQ0Z1Vh9ReNBCe0OP2mScUOxmTfOSODe5Z+ayxgMWGkhH7XtvmscjZqiju4OezPC
br+kY5jj+KI1XRwGkMk7sdZCi6FrFFeMkxhI3DbwaHRJtg/CF6mcJdxG8VV1iCMVALBUNxl8aS03
siqVzl+hRLD1oW2Na+2gWQ6DILJmTqk1CMxdtXHIQSEEWUONyiFob8hfllpgXZPpq1HYR5GUL19d
dvqIRGCRzUnVkLGVQ4LM0+soXiR+igFHlPTS6EPqMHWtEe58EmMbk8R7Fcbft1aPTiXhNupSB1mf
3KffHoj8XceAHKJeRT9wb/WKHFbgAW1+AweDI3OZ74vWSKWpgCYiJo89UT6RJBso46rrtYZP4Ghz
oMUMKxvx6e6l0ARpfrQSa7c/ozwd7aBT0++4FfUFYa9Q4oUCsKDUT0XeS/dE7qmGyK1ikqwhwWND
go3jU/hWHg2EUCm0ojdWhsNu+gmdQWZFE5sA9jTA15EJDb856S5+fhhpeOm5G+yMuGakxgs/D/0k
yTKA+OS2JQ245x6a5vKMe31U3cKhsZ9TQq5FeDZncvMouuinU14HkpTVMzrYfB+irZnObPR2blLi
/zL72I+15fdRt8C19jckyfLcOmFiwHJZvhr8SdUtg4AOl+4EnBvnAOuejInwfUcUvXXJdXgl6rZf
acPhAZj1Gw6ExUTFAag+7flIaLtJb+junymH5LE/TQDjpzRrXHUTrLeF0+wEHLg/NQvKKWiucaPz
h/PUQJV/gtCcCSPH3paIsOQOracPKBBQgKfZlgfciYTMo4NsMMD2ragefj1qHOix1Z2Y0Ax1vkvd
91W6AB+eYFxEeyaXNv4T861mqzJxQ4q7D+/n8GG8AyXJFJHzkmLx1drlWVwzzEa67J7bvY9dzIUG
yYgy9ZX+q0mhhl7a8417LWTjS/f3fGWC+a6p0sk1yiFJBMrmJk3R2H3QPXzfh743wfFZITFn6uoT
oGS5MqsCNxaNgjFIjyckHF4OPWyy38QweKaWpcRJL0F5+f1I6Uc/Zmiri3RrVG3wLCzF/4UXpj/D
eAjkB1dQdWqzKwvGSQi9o0mvoUiTVz1H1VEW+Ad7COm7ENvASQjBA+gTBSjxoepRJuFhXxzzoRP7
8v1a6UTJ7Z/G50ROtU5O4jKCYXgjEgTM67ppJjOxBcyUZwWR6l2qJHV2U3Umn8HrYgXuCHqJezmZ
K8u6z6UtAT4eYGQX2Tdr3KwN5EXmd2hZCTTL8n+tUhlZoM7UpOAEtNrpMSfDrK7LhtSNeM6wZ5pi
Ob3R2k4ZZTmVP+qPz3Ktf6HUqOPSRnNfX94c7n73nE+IhVZHbdK2Td3XSoNFHVJxLQG5NRor6XDa
WgFtrSjwOGWvu5jqGxg/iTKQy8k74vx9xu3fjPs1sgMX/X/EQe3kZW8J4/ajaDFpTrMVHjf9wX6W
ceJ9t28/9ZtjwNVoyQ3bBDLBCNHoBW3HD4CEuo5RWCUeKhkJpCStYAou1qNMRxRDjnUE4Fm8xI7Z
TvDr8FD5OLlRiRd3NRgAEKvqEVjVDsPtubwh4bOfo3DR/kJ/4sehpaQJcv6nzazQwHPxU45REO/v
r5oZ/Hp/nPLoVNs6zrOpsMm9FdZ6/iOtapBv+ONwQdaUWO2LoBzEJhf/ShQiUB6AObh2A3IS6r+6
kujFGE5bLLyoKoYihqRFfJhAw9r6uBlsv6O2DKFeXCAMPuuS8ka7LsshfQr5Hwu9ueLmN6VWVwfT
IEvgBW9mP1XZWefSojWw1Z94mWHcCoFD3b93Q53sWdF5LJKEtmen1JyvmJvE3xsNNNdvrl4kU8kt
gXzhn/5iBV8EENKqvWiE/8UNBertkATVoO/FvPcVMGVPYu6o6i0UBk3E6I1tyPh0KkZjv08osy9B
8woc4R38TgFEOcy23euxEnzClrTHHe5ao5toH5gSiwH4l4v3+9mwh+Hk/aaLC2rLLGMShtb/5sh8
BKuSmrMnWBDHcuA6FZsMUz5/MRS5GUaXqXMLvZR+/HaG0+QfAmvxvsLe2wIKREJ2n0efaQRO1li5
BzmXk1IbiLi0vIa+3X8SAkBVSj9AiehVo+yWf0vSy9yxlNXEOnsl525IARxzEorz9f+Xz8l2PthX
eODSHVlbSjNQtyld+4WcQfWddzBRrRiHfDRT64L9IkeCV9RwuhrCE3fRk/ZKvfHg5YVIcautsIcA
2e3ne+BjbxRX8CDMmZGLEpqhL3sy9J4uS7BYjvZIjyKVK7Uc+QFMKJ6jpEc1lTqRYY0DdsdeceVJ
+abW2exdbFrNZhdEeo6T7eUdPu0EsTV6dvUe+R3l9zrmcjPA7cBK19j7naHEZAP3E39zKbDwQu0n
UhrnqvOIVsdMCdb3MElVe1n+BNuBvro9L/LhmJFqEU9aGVBWzNMpceMFU2KKLR6XhUmutU60+7Tb
3cwPpp/zfMueP6GSOgcZFHCaIdZeGLrCSvaQ5YY9yeSG4raidn1NWK5dnjpZJosZSzWbF7+sPA2s
nuJp7dnRqK6ZhJ7vqW1DRldf2fc+nDK1eRAfHYAWyXddMlpeQtO3AHh5wDpFrPddz+0U+Xv0DNN1
lG93+aGtFoZ3Kr86zlWAlcnWwYoynR7wc1tbESoscFHZ171fimfJ9LtxMzDybp/QXmOq+hZbjeu2
IyIv4BD5cQptCUXHHmPV3IGF2K7MG95UrTj/nSQVMAyZlPPPIgJyMdpd0vrjl+gU1YfgdMWJ7vIH
izuUaYg0CokzkMOHkg/8jsZP8pPW8adAf0dI9xb5f7PTHGxl+VHeL2OQWqEkHfDVc4DcQ8d2BL7T
kfhxuKfPQ5fKAwAgyEb5y5eIkmu3deK35m17u1PXgubwDBkZicO3fys17lPKamkY3804FRMZHeq9
vU3cV9A/AqpSVzii+N879JCMEjDEZmOT0TBRfZDeGlyHXETz4wLCQTA5svbVN04TMi84VDAjmVux
WWZ3gvp8VtzBSANorz3mFOSCZXCgXXDeSD94+G0sc5KJgNqkKeWtf5WgrAwjHB87nn35GuR1upvr
xVE6IX7m+M4c3FlMZcisMjfQiNd2fvSDR8wQWenp8sx4RyaOI8e4nn/cL0W4KGH227GCC7tT0TSD
NywPCk1o4IROc/9tFYmRYJAt5x8URkTitcQJv2EWIN1hpiem3w3oMrCKuJKzrz40GKffb1pPd0Ut
HZt8FWdL0P16Kjllzx/pwY+FEGOoTZh3CE0TNK9GxaOek21zkl0sf06FZw9cC/85MAZOKih/NL5I
/8ZkX8Yt4XqKK5Y34tS6nE4w25PFkHO+8ZUfzeRc8C8+dsyYXYRxtg8t6W4A0NDIm8sjzfzxgIZ4
sObWuyhzsINhzBbvSPO7ySkkYolSE4EA0cMVl1Ywz+Ns8QivX2LzPbLDK6md0TEn8O7dZA9YcC0I
1278+dna8uNSjlbp8chvan1iSLRzuetaqalYp3u/4HKRHifkZZS8l0nAvBz9uInkEXEtRP1tdRLo
rVmu5kDzYMV93W0AACs75bagA5MZVUgrJOXSp//fprNFS/IQdwPgpUge+J2q0N5CuGfVknMVNPOO
RbSKu2t/SSHV0SeRIc9um5uuvlePOVVwwjqjY77nZuKZ4fDZZXZ5YDokc95f/H4ArZ3BUls5Fxpk
s1hrd5A9Cv2KruvAETzs/VxU/rO07fx1PwyJSXwVe/l8ViX+1z9hS5MyHEbmnu8GWSHAGMEkl/cl
Kmpxd6DPFDxNDpHR/8k/R8RJt4GmPa5eo1QqGWwIuJQiyG6oMssWfqFw36otowlYcG4vcegiDufE
vR3Xso3/JyhUh1+uDj1fJCd33OJd7GG+ko18tbmpnhnBn/jW88M89S5WqaZUB31gq8ei51gkrpRd
aTog7aP1Q0dBSTscB2YDBpgcyIydt3wmBGIqsrnOjOoD2hzSVHYcw/UhnPItiBQjeq0P3yQuhH5I
4o9SjIi2j8a7H50nly1YV/+Szu4WYw97qRQ76y4xwVDiZRz/7tazPFtxAgnIDQxomny+bvTREQS6
Xsp+hAux/pxsU4r2QPiM1vy7FHw2G5o10tbi/GDEYQilnYB1gK0d084RLWpiWNeLAztge7rHP5Ir
2byYLmxTcshAV1ww5nPeOWR8T31MVKm5gx6+4ZvwwPMYgkAcqpedrQokQtnVRRlvVbbSRYThKkvv
yIsUpGwLKi4whl09h/YSQXfsM9ubJ5BaZGXpGsQ9lSOvfSrj3iztLpEVnOh3qEGMs49C3MzIxyV2
3U9dWjdAXYTrNJhhsWtDYMRDcRDvNni+cmr5DhD4qlVo6veCrypWODR3o1IweMxZGBXZ1spxYXoJ
dg26dVrobS4VeQK4GE+LWhZBjEa2vQPbMjhumoi/aJB8NaGuZ+R4Eembzu2rnEWajMfESOdUQ4A+
8aVoV2ePz89mOH19+kBDmMcLgIRZFMLGfCD5M+wSweBpZEeI9Um1P0jViEr0g1JTpVUEVjmKP4x5
flLsI0ZzNk6B/KQsJ4RjJaCWpmUWnnW+ebgNhAY6Zc+bUxRB33sCUnKpouWfNcXPE/ZuEpz6FqQg
CighM+jWG2RL0XmbXarzrOOscyvZhXAsJjTuHGBrIpAukM3+4u8c+FKkZiIfc3yaCAKiwDNO4Bp0
sZn4GLBRpKDNSyOLnlf08v5eLJR7K8Dfq7Cd9Rh/hEk81TqaxX5MKDk29iKsQcQhW6WOEi8W6QLU
b0O67SadyeQD3g3+dkZZa6knfuslDccGkBsm9MOUU0OOK5/xRQ7VqLIAy/eX2NmBDBfUvjEkwE9b
784T13WTg6LjuWRBMDTsRCUqGZ5pw5WrL+xxUXTKvmT8HA8wxObk3aNrRo5b9aurHVTSP1efYRn/
+sjdPoetIR4pJ8rzWSrnxKV78T7dXxkOmtclo9bBHX3Z9Gef17mY0CxOP3CC+wT4h2BPVxaoCowJ
WlowCPh9qx0ctVIWrnrg3UYq6Mbkm/bYursCDc7/Go22SDapEj9af+WSuJ2ro6ssof5Bap+4zw9H
gFm+XGddFREJ6Fz0jrwUQONeb5E7hFvmuy/q5vVhxkwa8ZN6MqvfTMG5g5lVEaGiIAxHTY3c6yvx
WNEB2y8eJzAFi2xIxV5NGL4BDkPQMjhy4OmybXoSRCyskYIQUkeE0divhKqOgn2SedP5e+9zWw5S
hFucagzZTXvo5xacFPl3XReRqea9OmBGQ9u5AhXgCevJgp24oiN1Sedj6pLH3nNmvVv0Fkoiez3m
QmeuujNNuFdxa710D4mbbjEGDMZwy7xYRG7u77DdMDdNkOH+3LQgAaNSmQcFqZmew00FXLtoXXYm
1nLZAenEon+c3DRkGxW+qiqaF9OmRBel+o6kZdXUmY23RG/GiGEvuY8g5XhO6HrvV+OlZZx7jMiD
twG/QpUaesAl+q3RiU+P5+yaR8aL+JiU1ZMWqGi3x+kvhhkvGkeXPqb+aiX9bLAzRzJSxj5MwiXh
sbuHWoC7NAk3s4/lVm6KNcShv2wVp7u2TQIp8BGSOGb+jAscrQ4Ag/Ex3EYHlyiEIc2/G66jS/pW
jeHLbxg/HP+MdZPZxbgRkngu2RlWDsH19p1QKubHNdOZthltAZPcB75KWNcr9p76j20KHPX+ImeN
zwbhf54vL4nCGNM8SxhIcZeJhLpDrFUxsRFzEVeWyphwiWEp/dwkIOfImQFqxYMz4jQV7a+hrSDj
YYuOs4feWq7NXxmzk14rR/zdZDLDx67TVhWBMSRKBvktSd7zezgcwP5YrnRoX9UCviBzoduku7Sv
lH2jcn/ZKhIHWNNEWSeoStBcks2C6ipVQ63vvi7kojb9NdK3J4BYgZQGOmMzK2pCw0UlqmISM7FG
pIwDYBXdePOjwnx3zN23hmkyZHvP9n74SD8tG2iRIzqB3lRv+3z6JmVxktCHnB+g5pbkquB9+tbD
1DFCwK5ON3/u1CS/68I8kBIoVS2Ji4J1pmivyX4LQexH2fCaAsmfQRsZhN09FmzjwNkFG8xePLFY
XI+mewXObgnZdLIGqlfPhA7Rx/dV8YEhKAjl1Xih1zKXQAjSEd+reYsfxho0tLDssSfW87jTSk6e
+wBdv1CrweZQancfhi9UVLx5kbK1vBsLWdFFvOuLM+ldhFUNHV6vExzDrw4YWmZQTtVlJHCu1rtn
B7C0O5S7cx//5fOlP/3Yv4sFcQBtbOn6I3xdEstkWLAuYSQTjEKCuC9Ab6s28PK4mrYZXVqQm4E6
L51kpXfAM8+tNUXTLqDlj/L5cZvC/aYUec4WWFxruhnbz2goqDtMzB9mp4Udt0c9jAscgFxpg9kC
sPp6Y4/gW2PlW0Ag/WHWT1x7zx6bLqna3b4ifUon9bc2ejM7mrUpmlLD7fjWP+XLGkewlBnW92sp
jQJn9RRsKy4pZ4mGOunwjaSCKmeF+6RlCER7tkQ+c7GUqaS3xCzjETHGxMWrdy32AZA5kFwO9wGx
GovNaqXnx9VD0d9g62dcH0oPE8szQWrI0D6rko4Xx2da9HloUwl9uUstTK85TXiGsSwk5eNEdO4w
eZAUXxncq3t7a61FJLOfslIFPdw9NESjxQwhXTEuUC+DOcqXq2q50eAVoOmNrq9aZ0cM/kbpNaQG
Myo1/aH0pCNSkIeooWLYR0feYLwhHJihjZwRT+GjX3o19Gd2pR2ew0l19tHzetHRTV7+B8VTYSYn
ckVAde8B2bjbF5SgmzyA9VvRBXCrgqRyboMw6pza+0vIxR7mVjKYSJdzkjRz2Ko1Lj1TwTcdu0pL
CrAo4t3gBTuCMQ5fesfzZ4Cf360XeF8R5MP9ppb7x9/ihaQnaoKejfnFiPxB2or+r1TXIGzHruks
w8VRUhHed/AFKDBkx8jSmZlLN6//P+1JFs8R4Ec6+5PJEeejq4YUpFh8EaXNE2ba653zAI5XkENo
IxRILA9moMyS5CKPXykuGXOYpRZJ8cRUfg/0FLLDcoWhFL9D0NhUIe9oTxSaLgBxVzW0vuqp+vbj
Xf6W3mluL/wRsF35qwD4r4OQ+L/PNqLItUu2Xn0kGZIY75+1FX8Lv8DptUDdhJuS+2IIwKbuh+IK
VdS9O7zTetmR3sGHH+lCl7Ida+g5jy1ucguxkj2ve3I+UGfQbtx+QiMNg6uld6zgBe9npaUgoEeM
vNuZqqDw363HgOx07scs+Yba0QR4niti0sIdTDO6dDTXYENGTqgPVKcpUx0VDvyqGLJJDG23rIcI
LiZpFXMIYLw5euVrbWRcgG/MqZuvpsBYZuy5sJ4/I3IpvotmYopEgmCTjDrQFZ1Npm/nEn7+pr0D
oCnqyoQE1Jdb3eFw/vwoZb02vI8mp16FjdFT6j6F96piGsmVgxVeK30l5SCRkF7engs37vPQjk9i
FcUw1FzRZ8eMQAlNjofbYVm7kI23jgdVF5DdNpMtLEn6Clp1oi2dcfcJ8jHnFD4AxEAHjcteZdM6
+UHd9z5Uy2WNOCSegfrfx8WJB/8TTiF1qUBiX1RLh/4UNYuzq1zOsPCmYgntK8WIp+NVHJ+atIIb
XpH4asq3xIedhMxfKNmIhDPe0U27w48DoH4CZ2WsHfW3HZylXn9zPTiWl3K3Qeo8ky07no+3nMtP
iju5YLRuN/6ILMvltWrvkyS6ZEL1N9/Xdt8QbqrAUZHOZsOeMKnbnXnIN2XzeH2GYu2DJYj8Gv4K
6X/hJAxCTKGST8F8TAus095pUo1XQNCkeMuYwvqVXbNznGgfevjQlHrudaxT2Mad/g+pJagm5BZa
B5glBoP6sL5cSz0+/5loTd0X1rU2oubaOm2Ot2p4m8bqrTsvKpu6l8/9PbuPZipxdtJeYtUyWnAd
Uyv34eam68eTR8DMWC0r1C0YGRYlJeswC8cNTqyvyqXZxE/3A+Fq7BDV2tSYltXm3G9pTY2/SmAN
xAIStw+PU501KRORZuCynrS/iGlMkFRngEl28vwxk0TK/EQZ6nUfTdcjgoW8l8huSeVqBaNsXG0T
QoGdLQBGbT+wECDor4NAToffEr7Qu3D5WWOgJa41KpXnBRn7alS79DEzHYgU80ZFZuU1pfEKgTGo
p8+GNZBModblEUHI1iGkL4kg3o8LNLaMuzEuRwgQEtZKjIXQfFJ/XHRfcYbHEDHQtPVarUzEGTjA
82fk3zuGOf5VZi2cehx/pPGTlfAPfr/9dv9iHMtcrQcskJ05r5C3VJtR8PlhabYNVSBSyXzJkKJS
oGJw3JizsD3+QOoHyfYlu7mpG+7DzOrq+pGmVPJVysvGjQJZ0fwm4lONh1vvxjRUKFT9KVwppGBK
1H6bMGi+4ySt+qX4/r2N20xkwpu3utojEZJNJDtDlvHvDx+StNfGUgMndQz8Ajebak9ZXlsRhI0/
/JR53+LDKBSNd87NxOmBtcfESXW1SKUSf2ZcN/3bR0e5su+8B2DxpPp5k38NOVNMAEW7GPDsNDKX
w/NQ7YiYm/gUxjDMrCXqpfA9IS7jzn4IfTodoGWjUsRK0bnPdfMpJ7vLpHZkxrZgsTZFEAGEVOWg
Lh2PzAu8zr2P4nan4U81aHOMajnI5y+61epnteAaQ4amrCG6dTQgyKtSetk3reNR6nGe4ebEUvip
/3PO0fGDOAu4k5ZzORepuf0JZroD393EmoRvvpr+BRsQBy9e3cFDgtW7G2UJZNVtBD+yqV5svJSK
XuhmphxueFI7QVmdFssVZU34cGsXNKfqjPWN6ZEo4zxmA0j1CSes7P6cFH0V+PuyiZEMWIlQ+/5v
BUuYkwsnk/x4BpvDjrQpYxqnZWaLmmc409Z3fLbZ46VFdsy2ZJeWpUUB7YeGBo8nM8mVFQ4mAyOZ
YK40VMOAKq8pIMhACxiEbj9n+16Qg2pZ+xdSpyseSDRAJIxgJHvxOP4d9dZgaxKLsDqLOuyzV5n7
KxTdAmnsC4Peayo1T+ThzJtsa4KIUmsLhfMu5UEMx3auA4xN/T90E0Ybjmb2Jo0amFFyocbukobP
S8BnObHQcYvA5IfRn7g5zq3Zi/LNwWX4Jm6OqdqmPiWLJrin0Z4UiBURfXKueGP/WG6DxG0hTs9u
7JDBZCWKOQzJoFqn1Cs0rmqgGtE/Mrb+qoEAn3YnMP6iysMlBKaAinx7JJHXAatn11qyP2cqYzDD
X/GYY9beKeQMCoFiRrjTlR+CCBOkpzizv4OgiYQroVN7T2XnHIlsfwxGeBB/nJoKs4uql6skTUx0
SL1mq/68W2KKE5wkZDXL0TATckAW1344VylGzhlYU1XpXzeImHblrBZwVs0sMf7CbW3wSYiybvmd
ZWcbRgdfuZLixgNbWXDLn3uJcz8kpIbQ37TjD3l23bcta+ftn8ookCZq1e2EAJ2AOML0X6PnTg30
rSRECmU00oEXmxrGFdcrbgjttL1w+dy+cUfrGEkpQ6SoR7e7s3eMMuas8u4dRCB1prXeZPnhXugh
h6AkYEw5g8Xuhrc72pKsDm2W1+NH2iP8zXf79KrQhyTb+e/3Rbajq5WfLDuAXBgfjlgu6rfGEA38
S0vkVUyjTCl2BbVqncthpsbgGyw3oNe1KUrO5RxTniJ30nbsZVARP+86lskJIaZFbJH3G55F7DMz
3+sI6hfuuYrZCDMl0W9LMVRM3Uozj8+RKVN/i0TEElFcHhWKRgv8FyN+zrnazyol4sAHq/imzo55
X3Ld35ihTk+Hz5MNLKzDLqGxA6zlA/0Y42GP0aXWeON/OPNgsjbyvyvT3v6EEynYqZQxLmfrABKg
HjEcopWr9T05eG30mmmA4kHZmaLRkNdf5pINfcrmgCsVJi/AYWIw0VR2zwLkS1SOvK/SCThisMG/
jmf9ICE9RB9GI7n8nnzTB+NWG+1ywf/NUvd75rfhAXrEz2WjjyPq67M63PHA/d0v9ukmCENN12I8
T9CKxBfX/3/4U1OsyFNsy6fmPDl9vARqMoX8EpYg1Y5Un27sCv98r4OXX+lXPYmQEpibqfgCVK+p
ZNG+mT6Phsigjv0gH16Y3/FO+ZCFMEBeJ07gtHtdbpBvNLqmfyQT362uJmsxR0ip4LZsiGfp6rrS
pd8WgPav6fNDOODXWFb4E4Fn6IU6m4OanoOE/L4YWZmXZw8tiqUX0KKhn4Hsldulrj0+SiU3k9Bp
CRrVfuv2Q06dTDxXG1ZTR6dOxYDQt8R2aYmDa06HQOV51n9zkyx+jSU8o5/T7nV1KqA71YLeCd7c
nhMFxAmqgHfZZdBTzucUMVzwMMEDvct/MG7p8iWM6U5XwTfRpJMUY9HsRPCrcUzgDEot6mLkUlci
2Yrpjw1cgU3EVask/fjORsQc4nzl+1TPZH+sD1Tgn1uT92Usyfs2AigN6+IxF7V9TMXKzvuar1si
wcObjuxU4P82bdOc+ZGqzB0UXV5olkWNiAHuC7pkMbYoO6r0rwgNXMC8g0cRDXZ9LL0uMCOGWMkJ
hTmjcl565vItrPremusMLfFHRAkvm5j1Kw6ohrhkyxELvp07yg27cQdDj8zb0DvciEBfYrAuBasS
aBEspcgCw9ekhHpd3rJsKafKE0ng836FbpMWUrPIlweMCmVPREuBtZPYSNSCxpzCNQaWeH52SfH0
0mG84onEEKzEs0ezvpNXbZyMxudrE4K9CUh0g8z4AxEhyvCMHSTxatO7DXhLV4MulaO023/6WZc6
B6YZpl6OJBEhdkJmh6WgPkfpkZdIpHLQTaZJJjdSH7cSYPgXPgl1IZ0bw8ScIatu8ukXUs9VaycD
l3xIjUUD6BcLKM2bL8aYa/eF45UYQyZ3//jXRgduqF3+057tPNgHaN/3jMTULpCEd6djDR69M08X
Q2xBecIE7FEabAqAhiM+31xGtdBpITKIzTo1RIKGQF4MNTz4TlgrcUe6KfsGb/rnB5vH6gYqc0av
LebAcKuEapWFZaFDEU/MCjgYaq40Ty0gn1Gxh3RazoNR77g7yKhl5yitLHDthdhBf6AY/ysUqwbu
Gp0lAmWLSREsuNaF+VgjbO1TOaFVFkZ53jvIhLfiniJj10kE8Bsrxpm4VFaDgW8VqzSjtYVeIDQl
/jr+e0a7oFK5707z+zPoy3/9nXI6Sy6Hsjn+eUkGhwNXlWJVj48qX1ri92U53J9R4g8yu2OVg+Ut
H5lBf0U4jwYY718nI97Vqag8675LSu4Pjh7727Nk42LfA+AVxqGyiuybuGHxbwFEaPO1GIhLpKHy
qivuK3whI32WSaE2W3w+24OMrl0/YgAvzsrb8FLGQTsd744qmfUYraNH+lTgQGV5WhAUN7iVdPjC
UNFjiuyMswkDPm+DdQjFopnafPVyySdD9iV9PyqKt3+w9dGvMUoSzJewYW8YegNzoSyjUvlkI5/Z
j3wFSP0CPkGImxkzBy9Hz2e3SqYezoATsj2mqtGnmDsEg1R+riP7SkrI+IzdiAg26GD5Jtda1pFK
MGAUU7RcGnPehUTnYzizOhnYld6tmGLFj83dGacBz2RxxieqQUrDmlNglEIQgDnrMVwql/Dg+TWN
7LLpChkyu3cCHhLjanJaF+pr4oU0LJGaHJyNThE5U80NlX+uBGxp1+Z2L+WDgT6MC3SnlugDCLVq
t22wHRvugjKjqHkMr/cpByIIDWuYclq8M1f+BbNNtTz+zo2MQQMrAqiz5PrUI7Pe9IJ36gyDYl0P
odcnqnWT8mOFjLqWuk7PzT201WNvJk1r4m6t4jOsIyqySroaAvR62UJL0hvd91rMG0FHnqhQgjAf
l4yl3qXasuAOTAoeKuiN2Nu94m48g4Vlgx7ozGU9YpJwqMYPDI5FwDgwHghLSRXWMn9M9FA0ct2I
W9Wp72twLaDdTL1SO+iTZNMyRTBRNsM2rL1BhTx8Nzgrvb2ZY6N4CsVXPj/CAjeka+Z+zZn6uoY/
ABBmTSRcY0nnyw/zA43w4rHl1sqNWQcjcGZGl/oDOwANotrKWadMNNps5pFZQoYo3MWKPE2wPn7p
D8IT2SPqKYR22/7pGkU64ZzMaThB11yjZDvNpdIVy3zVYMwGDbD7qB1w2NQz4nRxXRHAgHNe/Ioz
7Jt1bWdfHowRKaBCoB7hVcHwzEC/bgo0mIGgDVDwisV/ZUAqwvT8WhPxtURA0jzhCW98bOUNJGab
/zGGYZMdTP84lmugmdESsQC5Mdw37EZGqbNlSPDwHnqogVl/IG3o77zMrTD5eD67suZEqSPH+RW3
MGSKGVMS95sWIddSnmANvxmoWlMQVPtGcCz92oZx9E95GLrvtK260ybf/usq+crvPIfDNoaC3Yiw
aXManRnM+zgLCd/qufos4JSxnVehIq9qL9Mkwpt0oWaN1HmRkbH3ygi+HIKcPW/2UsP9M0l7rh4N
IyYofg1e5sO6QkymnpguIFId+k8svsvBLefu6Rsc0ZKilnghvvivi/LU0bcUmTweRh0QQX6+bccS
AXwIlIf1k7xx1fyRYyAuFj3evEL04cBFmAnW6Blz4xlp2/wLMnS1STKFXQj6wWNsypepinF0OERF
6TQh42RreXRDhMXZ6g46gh0WGbHWsXlnrLQbVU/yBm4K0O1mpbxChgJZOgNM5wtXnCckVxAiFNax
swurH9Jf4nvVAyNAbdm8KcKp5su2/lJR/ro+gQJmrlz6FykYjN8FAjFP8TL6NoP2j0J/Kklm5e3J
S3235514S2wFPwGOq4MYLNaRxRml5T81CBxgC+X8Q7DBhpcqiihvpCSt8pNx1kdj5lxBH229AyWp
vxx4yqjYlD/NDota7iLHDw0iHwsUjbt78eo3885mpp+Ik59c4NntOXN92tcnDQ/UJ5RvCDBDgksi
M3iRSM8aZLJzmpaZ6EgRShJ6AaOA8Hh3QcnCmXqzP76Bw5cAsh4X7ZgmrjqFp6jneF3HC3nTK2OA
uC8VkPCZ0fiIc+0zcGsiN5xYXY06bflfd5zz6U8d35Brv/fnbNxt46mqxHB7FOP9AGI1K7v19en2
TJqKSvRzcLYLb8C19SgV5rZ3TmBIATGCrNv095Bf+JUs3OggoqpSTuqxuQsDgOXrr/QLmSsiMIpn
haqXEPAL3HrTgFy+GohdjWd5Nzf3/NvnO9cRmN+qUjRm2LnTJtdELcd1J2PwlmzzyJ8YhX+mWR/8
Jt+Pb1C1ugqXW9zGxSHkML7BqDZEqSinWFf+Ni9gfWFOmIAp/vUfYQrxqKiYwUyH3iD+NP4m11pp
TQv3SLQGiTbhdyI+SBtBUFJ4B6VPODd7Mtm7Hx+90ds3ka2WOvtVpCo3fyEFr7uNLrI2IyOUM9Gp
9Ujdl+YeZbCIukyQQWdoddKJsPka99/q5tMMp9tUwcnpoeRIgCtelha8vKV9Ovitf2sFHlSWZdPr
bL7L3/Y+5E253YooC97NN/dgyquOvbNAW7co2b1lMMuUHdC/AJP76zHxZXuWXcKld4/Vfb5zhe/M
fnuVATTHNUP2BXUw4CPMgOLHp9h+8tij2g5MCU+S1pW0nFdDovU+gTU+gEEgPtjbp4tirQiFpe27
bHpsBZVr54DUvaBI9Egbwflw4cDssMRsGRmphnojlCIxF+COdcjFbh3fapu3KPStUcc6Cw071HhW
osDA51OdnsiNkE7u2jqb4+polaQdwjyVCSLOeOK2cEs6jwIOz8Gg/dfYE+uWM1QV1KGnB80s/iHN
hZY/0PY6UjFbzBjU+dA0HHALX+cf8nwNOJFthjovuCrOfDOLI1PZyaH3pUVvr8DRGkHkUsmmhqBb
GRsOhkDYAIBzG8EH8ibuSyMNKrVSa3YEbJPYVOR01dFAF9eRtEOFQKaZ6z37GMx1OCoJ2QoxKLTA
Tln8YMC4gg9ymswSiqi95sDgPJvmxz+7wytGeNSUDz3rcNZRqvDzkKkNAMSFD7uMEXd5OkoEwSao
i4UJnbsAskBA2511YYrQFeTunAT5dJjQ75jv9AVBvsDTMJB3FQBl9UvgHcIO2zLnukfoAqRQHQ/m
k4fSL+yq9AOx/icOlULPJnIICJNGd7lB1NgMWtxDQU3wmaPssylG7idHFAbB0cTY/G32wWfSwKej
+FWjF0Hv5y5MUPJVV6yMEN89KArg/TbkFU+Y+PHZ4TVmlspkki6Lw7uAiR19sBjoLgzT5AzqQMAI
tDJZYL9wWzi5nUuE3kQqT2FRsR5gr6d8mylWkCdDE6QStq1Ta5iFFihoBkjIFr122KWKoSgrjMAp
0xfLrVylRceG5g/QesTWrASGeG1Iic8AjuFR4QRpZtmuHxjLAN6m/d1dOjcqgWq01w1w0MGhp7iz
HKyCbS4txGC9/cbg01Pf659nerK/ebsJ+e1n4YLBccT1ChPxo0OYNr11q4JBslpTriXf+4ZbK74Q
h4mLiva3xXgXeKQ8cldGOHUkOEP96CHQGMZzyaJFE2AG/LP+W+TwqhosLzA62NQ1BPYHwBIOS4+/
w55PpLyRKU7tL9Cle8dBid6SZ1kuB6WmwKj7v+TA0E1vaQFIJ/GI4irjF/RkjvaM8iVlLwPHn/tQ
XRBkIhEEqVxPrlA+UwPngkXwB7DXzoZkxKM7SzEw9lxjAvMOZkrKzwAMFad/Bj5e1LQFrImKY+7A
ieIRjlkLYa72mk+m5gG1GGro5N1ADD8feJe/3GB+wnt/ki6CHzbu7HWBV2bqIFxhk7YibjgOECwF
VWY21NQ/U4c8bpSpCDlfpgCPwhZVH4ea1ntBwLl2O5j0Ym6AMjjw2geFZRexofBnDZZt7U7Qcx2R
7g0SIbeXRaDQuqcxlHs9rUzGGjFF+OpvrNeQZn8rBPVSsAvkSPInFrpnbrD9rQAXPBe4LXxp/O5p
tnKJzZT6qmtSPB8VB2hCi5lCflt64I8lQQGzZNNL8x9N63qZbQC+fOj8jmgdUPgfb+LzaELwCKpE
Z1RuShiaDFXiaP9FrO8gb1k5g+w5Mag73I//+2++ECLuNpr6d3rNYrvY7913tbXJWBJvU/QQnPZ2
gXXfXjMOI3dMY/+chwWR21QYzp35ItzrywW0NwFXhWvn/tANu8dm/9ZZlYXwmQA6Yioyyl5x0kaB
DbDbYwlGybfqAwBqaBQgDPH66R82Q14Ao/8qR0d3fvFW/9uRjypOSnahl7msVDgWIZQ34PahKOan
IYuktu1Zx3f+k44o1fuiE1UWPpN3+23wu3de9mgfKcHhLuiKmD5EdoQprN4DKUGjZDEt1DUkFCgG
/xUlOxzOgdVlDtHph67HHVfj7dwbi1THaaZU7VtOsRre6b6yp2ugWgH85AAKxUV09Bw3L13GFQaN
5Bt4RFl82h9qKmUs2LANg3P6V6IpJO0fouqQoO1ldSlmP5hfZn3ptP4AVlI5SDLs/P3xAyT0kFsG
En8eGP1unSoDeTdgBQ+txqdyL0lMvlb8zbq++t1aQKXrZWtFusN3khuUUeD8Ofpv1KIVOpx4b1se
WNtUQf74JK4xGxVAUkhQoy7Mq0ngg8+tfDAsdw9+fJyW6EU4TZrQe0eebi56WQx6G2sJIopLWeaE
D25UrGUinc8E5ay3nHIWnJ7bF9VAOoEeyDnv12Pxulgj1gPyLVuEFZtOLYagofkaBByPR2nCBu66
Sh5hcNLsdw2ZUEWv8h1r1y2fC7mnNqktsocfOXJe0tzXR4uwCZiCzQeNCiH+37xC60zg3M1uHuDi
s4VrkCDrL+uy8nIWAqPI+HFhCXWqjmjD7daqtqstu+JOTZgM3jjshghTilTOTKTtVYdnLgUlPz/C
7NjNZQRbQujvzxAMbaQainEEPV4O90A54rSxuo4lhwCnQr3MJwGDfFvOT8sCH5b489TFINNiZwl5
l/hHBkJ46xRI0DZ2y87MShIE7IIduF2kJzQLy0GhWYN5ompmaUfrH/df/A3INxnyDKu/e9/y8W2g
sqS0bfBHhsbOvwsmyZFSNQhTJO7qg1V8+qS9Pm4As6UyW+NZp7/hOf/AmAEirCPHe01ZHttu0ukq
eZD1EjqWp1BfFNEEmg0d0LCbBurkGca+cO/NKudY/uDl6LtMh/WWWPKgdl+mZ4p1wAMOLHoOcABr
Yt5brSI+UQ3y4fE4A4KaKz2G8Hnow7G6kEqgLJUExKmJzkKPusgtx6obgoGgSNAxePfrNhja+YN4
catMuNcLKDcMj3iSCD69duHjppfkv0bjAIU/9Axq8tCk/2bHSyhKHbUteURudUL4nyi4ZBPE5cjE
O5xT2ZZ7+wLWbovzvsCM4Th0lFZPvOZC9oMyEN7t5kXNnVJTTUptljUlchpN16d+9909gzAJ4Z2l
SrTWXATCHR9IG8JOrh9mrJL/ZkH9QYKER0Wtwd6kHpDwiE9ZAi8HCrQm8bEy7snP/CAZO8vQNNIg
TfkURTfUAJwXCAr1KnbfsD0C3EsAqZL1OLaVIKgPQh6omjapb1HCvMFnna0sSaRCd/1ffIPxBK70
zVTj5XQWGDDfZVirFqwjucHC4gT9pgPw8prKIhyZIXQDiua8prQ0K6MwMEu1g0R6zAgY1tMqcXi6
sS1bNjaXv7jSLGqKfOiX91u2A2a+JwWkPZWN+rr0dpvxDGclaqYxrZUNzaZ9Ul4b9sESD6xAe/z8
jvc0R3SrTUsdYCQt/6wSIfPj0zwmBvC8NUenr4uSlQl9Tw38EiAJ0Emhh0Z+Oefig+v6AkfkUQI4
gKF1SOqnEdpPUHcICtlbs5vu5Cuke2AwQRomJm/mkfxTXDXjtUELNpcRZCGceTWYZN3/Eor0V2Lu
XdEjQCfqarlwYEeyozzT5FBJ1n7DVtJ1zNVgGEyQj8SaX4/xwSPpe+kBeSIXUWdnHhdIBITGR23c
cCEFjX1K2dgNvYEbYTeHOf3j3+UYETv3aiNxYZ/c0M5CuLsNF8SwJywPRJW4+kYaTKB2UB/5RZeE
mfaEGH3EA+axm7kFu0/H8HqENlCyRt9ep3eDPacrCwPnP8hQDZu0jrsELxdF4CmuMfl+yHFK6Lsp
YoRDyrNCAmtr3qgHzDLbk0zt0W4r9faQ6RfZncLqQIVlF+c1ClO5IHJLb1UALEae6pTMIh0tWNKq
3uvyW6IBxV4s5rDAp+5xnY1rY8869bxp/VnfgOqmeLTBO7bmsucC5tmLgCuVVWhgQMvt02lyJ5XR
laZ27MCNcGvOM/p1kOWV8++owvOc5FWXxFsDX4rheldjfVCWwydUk3Ff24k0jmXLwrqH0d5LYC7r
QOmk6mIbMnO4z61bXsgxtZbmfq2jxOgzb7nWUy7e79629uapWf7CbXomGJmU4Nj/iDM4Rnc5zpEt
d5dvWd1DBy6vwNTXKLXiNnelFyCorH8kKtioUg0tv1Bq1O/NolI8sz502elaFhKoCYdlvlZ8+r0l
KKOwQklDsBkbTssAgQvBgKEt+rSmXLUhSt5qDw8AfRJYCkxGqm903pcVDPvAa7q4bbN9WONc2zRV
ndqiLl+5urOZdPsyLSLd74eEMcNZVgfQDmcwUyHLPEaV6OzsFluI4xpcgcCf/foDFVf6XpapKRoV
hFiYfA0aC/oR3VDvcIXUO7B3FNdgMb6vOeB2dXL6yzQdPmiJkGZwn9gRvnNpt8/3byphDsION0UZ
GzU+DOu2j7aaPhnbE2VNt0xyy6M9FSt6L5+58P1bpvswePH9HrX98H9OHREnaSk5RZ1/hIblaxsT
yBleQeXBw1iBDW5a6PGsz7dfHxVFDIA6dT+gf2fGKwlj+ZEXWZGXiz1JdeLroHZ8ZZRQRagJhFo2
3JiGYQS3uVS2ieozXdnu4bYuo8pAEnLGTWN2Qcv/fUC+iMXr+cqiuBT9IWJUBdfquUC40o411vyd
zwpSJlYQNoeTojHaYFX8vqPTabquJBOb10/oFRI+hrqYB72XbgHEbSGqTi4eb1Nge07BcQDvrpFu
qwDCAwxVbH/yoQ4piGQZYojnxWzHO3H/HQ3z3k7f096yI6oQodovjds5adDq0xzgqWPuf9QnEZ+S
qaqlayquvCLFZ8SYz8bhSgIRz42XZHNCXy0QZOHaGAqGfUomh+BRA4m4sCRNGqiDOa5VsiX2Y1uI
98yjxOnUdJ46tr5cXcvEJNHe68+5vdFMjzQndt2ROoL0oXljXB6V0R7n4ORC0Y3urySX4ta7LJC2
0a55QHGygA4r6UGpmSd72bQtkr2k+k+feH3+n1KxGjMKAw92GNqOYU9ao61HEkJzf4VAYhVhJpoW
Z70v1dYaYoB0lbu4NKa+5K8XqQVBVlWy7EO/7/nLSphbekBhygAggxNCUDL57vUy/S4ftUPYVhhd
HBhfaOx9SEtITrFO9z+NyZEKyjJg6dmLwfRrryTKuDy0oRCxEPGjLQqij36byL8j4FKhaTmLhUuQ
Oh//M6PxkUhzwLCEzNUWbjuvT8WZEVzBAnqyVVFhJtL69iZYJ/88cERRM1dRvupxxrEJN4WBbdma
kakZNbyzbFGdXjpoBN2WpW3wMX2zC67kaplKf14gI31msVGgVr8cVA0qg8Kkw7LZX+cD1fEjzxb0
yGOBcNJcBSKDu4a0RJft3dS8AhnNwyWViQJoFu4tQ4ShEfcBBE8OEmyeCdu7q/gKrmlq6QExkXe8
xSKs+i/MNGWMxrRQkqsIkuHTDybDHCAzEH/bs09LTrujrnFidjbCjT5EELtlNVvtXvoJcqsmpFzu
f1COKYYj5C1YYo0QEIc7jQYixUIjuH89rJou1sK4aW9LDnD/r4UBf8Vvw41S8hM0lALIosJ6K1UZ
3C/nkrnU8xOnWqkrLHOY5tPDYTqdW1ZSr/0TUSKLrE8D6xJPvT8Uud6LT6qsaGxEkNAdK4qlxf5V
CA/NJPfxtrRn+RkEs60S83jgKb4xXpf96eNGOoXyaQsOhKUKex5YMagqsNEiV8cQBtNRCkewcIID
p6A1owa15hzkKMnWoACDSM05YYL1x1x4Z88K6jmwWLAqyuezuUjTwgsY6niEnEKSHs1tYrjvgqzR
O1iVm0ILQr1YYCIT4Wu5zOdR7jDUcOar6Xks2XbomkKeBnYsKk9mAEZxBd+BPmlAcCf5hS98kj5w
vnLm3t+kel8CfASe2nJwTwryu3v3bKUt6//lh5ZRPoYGPPD5QUacDQ1vtQlIlIreN+v6qrY01wUk
B+mIQPEzHwMJKpvomJ8+Rd/Ydbu66sO6YI3nFSZxrvKNfrT7xzomUUKUfkcHhU9dZoBnI2uCL+tb
1tEWU3MxzNiLLHSbfHoU/yP7A1sMcwnq9vZI6gKPGpRYtCGW8qCu6FZcLwPwcH9q+Co8G1zyAZg4
MocQz3AcGbrHSwildcX0cpyU02TAaF42G3Ooq+EWWRpeEiyGoTDagFFKUI5sntcCUcrgI58lVieM
pnfSzOnk4/G6Un5GoULaNna8VGcVcQZEMozTH4oFdo2I6Cyt3WmMv0/nas2gkChyqtKE0jtcjD5U
oUvP30Izkh+kvTd7xWZTB128mugme3uguXfTe9Y39h6KyQ3pN+oJv3byv520NpBBJfsubpGshyOP
/3EERR1pqJCs4BeCiYuRWUDaMW4wEggEPWIKO5cH6W8qdnINketdXUTbuLhZv0uiPRAhNxfroQrr
S7eL/52g4SZvrbH9z7mFuG7v2mgnoHQ4LF7pjKNMvaW48u+kJJcff0PlWB7IPCcQIDoahPVDdjKd
ngds82Q8cRJifxXsSTOmBlVXZdhAHlyLIanS92XP8s3+RMlwlsF6P05MGYdvFk2pyXquGGW2Zgka
B7P9u/brdgL7SxtIghnTHuqCvnCYhVOchqvmRSvWEz0PvOXGro91r5P/s7LXWLtCbtk44uuPxnf0
1/dFUMbj8k8o0xwH95sDXHyrsmYpiilSEGHz24CG/uKan4chy7mC/4UYtti138TU4twF283u4VS2
hGAUa5QC7S7zAgUoT7p2NCyL0Xs3Cow0jzWEPVLecjRsqhRLVhZQrO8r0WKTCOYFSKiiE5apjzJh
Tt1uJma5NXV4N1ts52UH44afqGAGwjiJ5XPozj1Aim8K8VUj6qBB8AbZJPjnPhR21cizp5G77IGD
dNLz2E0oLmXwyAfLkeYL5NZ9mBXtQOT1yhlFF7UaCxKMOqDL/9eG7oowR92KOo47wTDpboz1cCpG
KQvBQHTawleJnFEHHzgQdpJpQbMQ6jkdh/i2M5Xx44bQoM63s6ej2YX4B4GYkrKuVSpj0jf9DrSn
BmeIhhCTk113f43+DPRCBnEG3Y/BkowkHbRRwTtIIDwtVJz8o3hxeF8cDVNpQH6eZcgI2eJvy8Fo
EGJG3aNKDjrcRnTAvZkoO0Jmyovr1xgF9TR0d4hXkH5ok2qQ6pZcIdvgYXFoMw4V8eoM+8ur51w+
z/Q2T5zmnCtJjSkYcdAfKike0OcPv5GNlI6D7twwnL05T1QxxsvO8SM4D/Okzg1DgXy2gZs0ifue
Xv3HDZ78k5i+ZcgGQPMSSLhUs8uahBAKoHypWr8lM/R8SGZipr3TIxjZZLqtMS0QFYPRVc3qVLKf
Y5FhbAgs1CeCO4+KWMWcqffsiP3Hv9tapSx7Krf0JhREkBX6dgpkNSxtVrMkwca/uRFzZWj010ht
CNdN7A5FCW4R9IH4WjYZMLT2mHK27bt5zFOaN32EjduJFxL4LkvJuIBetTsqxB/tMv/vFzze78CR
lkw3M4NFRvbJYidRaFVPNix25AWEsdKdM9C/829CAkveHFIoPmnaFVREfiXrgCwOTjjiVwa84JN7
9Bp8pNAyId5PbPl3Gdt9WywOM7xPdFyNKwPBwIn1PeF4Xqivs4/iRkGKn53zCGvfFeIS7M2Hq+jU
L/GVxGHqUNXWA0cGMzrkkpJDvNJCSDbNlu4FFM+a08277haFGUZlmXnlu4je/TP1sA4Of2d6CO+F
9xeKUW7gcnKNglyIk6GFaPtOMyJjWg1W6siwksu4L2L9wU2UNsqbIdWU69qbI7Ry5b33c1J1K2QM
rh0jYXh55/8y/pk9Q66AtPKNP9MgTIlzKans1VKQKSG07+VhszNl51I5JICC/B9T6z8mzVPadLdR
Ss4d3qQDXqUZKsaByVi+eW/mDNa/yYeIqmkRFZj2qv8yDhEFZHE+Fkl1v8mxFcB7wPCiWJ7P3E4a
zIabwd3q0efSWjLXHMfIp94qOOIg3PfkTwLtr2cPsbjGjZKVMMUKLZE1YtUBqv3NKxntLaW6peh7
bz27bZNovj+Z9vljNz3yFEih+dM6Xyn92W7OyViEllZBf15P2+ukEqw2ZMJhEG/LsdS/xm84VwYb
xta/Au8UuRZfLYZ72OKwGk4WFok7pc9e6WNvrxIxFZPBAbHHQ+FoPbb01nrVVYcSCh7yN6Zy7X2f
/3JlrZtM38uOMfI5Vtxuc+V20+mja+/XtQyMzo0J+jajN38V81gF4/rLSWV/Hwn1m3r5Lh7nDL/b
Q9dqvBpXGYJcoF1o1xEt4KgBUd3tdzSFbGijApyTJ/kryf5xfRm7DJy8BXN6QIpw8mNOacYq13Pv
t4wfYzhvjEUkXELV4eLYGVmOAR1Ubu6EBcGArmC2JjcYC2Aky08wjwdbZJDG+myjbOlbDQ8vU2+T
/qV1NauzCdty/vY/DGMXm/h2qiL/ZDr2vC7oiP/Bg2rHz0w1fKrejjFZwjfV/LYC54I2kP22QZnk
ITEUQ06WbFtp6FnWW1oaa3d+LiQ4eklLPrW2a+XpdBBeTIxtv31t9FC+fyBTnnlHx/zHV73C14X0
x3zzlgmbxc1WD7+ufhMlR6q5FrZHGm2LdLzcVkqLfOfEUPQrQ7VZLE9iqmqF3M+Hhf3QCH7H7q6K
7arpl9ncXCmMwqwX3IdUHEzfc4iAoalUhyppj7MAsuugPOSHrtnYRC4neovhvoikwEr4ngUz/OyC
HfbthISbT5KvrSStLkzfICCSkQB3a1eDKogfNWoaf408Oz1qNXLH1y/SDGKAfAU4cqGrdGwTw6Ay
Y3x/XkbEwFk7TodhpbPYWQCY20ZXpOur1l1Qf/ohAP++VUz6X3htfqb0X/V7CAGKi9Ir9NtHAdzK
fsgmlVQWwOsd9sknBk8ea5aQqYqOoYAUzr5iSIJPb8285ysllgyFZ1tUCGWVR2w+wWFJDVqrAZQn
hn5FBtARUK0E2iSefWHX6r6wWP9jlWUarVvOmHrdGIudpl06/rfSSf1PKU0bZ3I+xZAmV3JQtzs+
Xd5FqDI7RXOFWKo0cnRj833lk7hvFXO7ooWLRCMe2WiLXJ4bw5s48H7SclLG/BSgxnSKzPU9KGb5
BXmJ0/xHF/xuGYtMChRC1aBHP54pi0MwGpl4MIZ9t6JeMZYQVm+JV4b+GZTs2GI4BTC8LL/+GVSN
LWl9FgZ7bSZ01wO/cn9R1mVcsnnHiaxBfQpYLetv2mjC+vaDJYe4gbOxh7IZn5xyZerZLCF/Lap1
nlKfvixqmYDVWG/V0lJE1NYqjL+3WsJ/9JzPDNczb259qGmYbPkCoOvqhmymH1x2dkegkxQFrZfy
rVe46FkvdOweHugPhOjk8JPf5K32S4YNYKkgpNE02HBxwYmRmmzHcJhnJCkJa8YTUH47LERO4AjH
Foh0HsmKjMFSzZh9ga6ohLdoKxBQWGHbD6Z83RbeWerxit5AGXFbR6z7/QDWvByh6+yLQuGSfgh1
XTJq3aBtDXB6M9EXthG2Fk4cVfMnpC7Sf24kBVuBHbdmyKPPxbZUOcTXrTMKWHv08CmV3/eo5+xY
QxRPL8lWB8Bj+CM0WX4ggOrbGIKYmDmNRcY1IVjNPczg4kcsK1nWmecUT8q4CyGHZZJ1eZX4IVcI
aZFzRRNQ8EUAkP7HgEh6U7ebTpyYJ6UgKsd9T4phmKiW6f5MobH05w14YD8eH0cWZCljYk4YDSyo
wdZgLD6TUy7Cf415Y3+KpUHQtbaEqlLrbA9FhFa01B7JSicQ86x0SQqIwqdpdLtGVqS33oFS5ZM4
9OWVwqHHpvPgXZ8+to8L86FWHJ8md/sa3aIevslEFRIhCtSk2jTLJTVtKwKCfe9MXhoXTBhCmXjF
jMtbjYNGsh8z3KY0Adx4DVsCkO4iM6rBq/zEPzzEOJ1wI47dl2oX6Kc442KW26MurY/LfIJpySGi
Bw2JGzTfPqlZx+FDADoYmaqrsUnbfMsg6slrBK543c1J7CnFyybgjdVIJgvf1FmLuRKm6VwiOEQj
9vtxEb9Y+AKOCV/2Bk3qHVqp3nQu2Z0qe0xcnU+jLCxOcnakFHiI239UpiOnbBJFKkAmtKjEDxb+
98Nw+E1apC+fPeUfCukEQLe6w9yU7FFS58pafy82icADJWJtY7CH8ilipDMpjbBRbNNY87oGgfPe
/7TiEojutrQJZAooMtNawcpb88/IGEiLEp1mF852F9/WABqpK9E7tOjRG7akxMqbU2A3Em/BULjE
GhCIq/Nq26rEDsnP8nrAjL0GtuX09ctQm1vfd7jY87nemLp2bhX1AhanmCEC2yw52o6yJt9t9rn8
biiUgwM5Kf/si1MPAcYXlyo6RFQaZoc1/AqQ402ShE2m/TbjwQVLdRaa8piYMZug/5SrYynLivmg
tS6POKV5FwE3ex8koydtA1oFqYf9qt223qCevpe5L22mBNZ8TDzB9THZFxkybl+dnsSdhp6xsDn+
urNbOtIDWQaNz/nhcdXaut3yremcUwASrnDL0t2uranMo5Dk4/aqc1cKO6d6hpprd18KzdENp1cY
PRVnNhflK+ZdYrdS7GNFXqnhvC6BdYwpcLiAtqKPfZ9z84KmcvVnsC1RaXf6Sca6Fv6jjV7Oo6HB
fYrWTfC75cJbzM/NUgeUJJWIbvaCpcpDioXKk+PhWD1UZhSCyqIGzn6W+eofvY1fAegqkBu6rmHt
Yf6vdw7Q0tzGL4vYD8knvX9TJPGFZcf+WQHBN15CRiF41fwvveGWYP4d8ltvn28OSQThBirW5sCs
xtCLsXnAwmaaFkIkxqdWT23k7gFkVLZDK/ZFivvYgG00WkrxRgooP2P1VRe7bVfv32+J1J610QvJ
lRg7o2TkvqOEiUw0HaV/c46nJv9PPsGT1Ng4efydHcbOUTH6r+Z4dMKNQwN5QMiX1yVNNGCLKpPE
b2b1fZ/lxmHZbT/LSdXM7Nk0MuEkEVKvmRYnvcPbrUVdqoqqq+So/dHATA9O5DH3DX4Lt5nqyi/Y
7HCX0uAsJNPnXn8TCSzmMrEJoXjOAOU2ldy+LeP8eQAHLatGrJqMbPNQnmEtYnbZFSgOxWIbH2yT
QI/MOR9IMVpo0b2ammwj25Ec+ojMUlQN+vVEkRI734rguNfcssafImMZ/gzUCxWSNXrCXXj9CkwL
jSXs+OFNPqZmpian9QW0gW52KO1TcGGlNjM8ktDmOLfHbLO31sZfozCNKXNgaYNoIVtpJAB5XuQa
FosY7rKAlzlY6cTquAhu0bHfc4RU0o54UgzLQQTsEm0PMH8k/bFSORs0JpIjA5S1vutRpEsKtKGk
ZCmpQJEVWUILOkYCAWlUDdatRKErdVv2kbvHEbYaNTd4zLEgB0Rk7hVYMkqF1IPvV5/iQnXs1MvQ
IMrn5yei20QrZokCWOXh2WIrmzYejEOSxFY84TMIqCaDCPqJ6X6aSZs0P0ne3QjCVq1tktVjL0uj
bWsMA2Bspe3eCkqQscNJWryP0ermuno14bpaFuOoALZsGrggzKjWroeQoM3kWYoZ+AjJ7jq6ZyH6
0E8vXVcFyvZ/SMJ/ScQvIaFoEBJk+Jq5shlmChbNc0DJU4xZrEQlE75sMmJJmMcxzM+EWEPk3ppV
Ud9xP4znuJ4hDdE8WNz+9ftLQC8gKlRMF2rlTdulnyghXmImKq2rhTj+b1bjx3m6tre1tog/jI+c
Lx6KZFSbAa38bGGdpUKeTtUQnuEOWdJ4cShvO9nWIC1Vs1fVB9HpjLGzVqpdJZJ5aWvg9g77+vyY
VPxHaLx5t/na7LNlaN7VdxnlL434DFU1yMtZokR5XA7fyfT9E2f5GjH2vErFYxv6zFDu2x4XreuR
fOLqv1+bdfUh7GfpniuXj3taRLYnE5zBP2QPs1yAq+R0vTy0zIflzCypdBl0QTj8cpNYb64X0CEM
8RS9leSmmEds4K1IHhSNgCkwms2+EB/evgYxh/UjbUcM1E5Dd41Qkml/2L3XgMW5Up5S6cefHWK4
MVCE+JWDEdFQjpPCiydRya3K1vGIu+KCrb5WGCXSZ2axk/ObWrM11Rnmnn9ZX/zRLhCEp2zWXuIs
T7d3ZrdzOY4BQv0/Z2NWR4IoWD6pCQ1SECGbbQ/CFySVl9DFYGn+gwiNaAnKMSr/5xf4iqbsIjmL
1Vqn36jbB1lKYstGHgNp/rsD01RB1OygpN6Q42AFEPi9wGDfs74xz3UE5E7+us1RcfEuyZlLdko4
5TtYErbaCyavoTEGd5LDQNpP6UI5NM6AGNubi6g2+7vRYRH8yatMK7eNA4Xt8FR/EVsKfL2erwzN
mS9YNy/hLgUbdwNGg++gGE+29KHTxreX0Pz1BJyAKlS2wYpi5lQUkO2WP8JYcNOW6z3V3gqpAVPM
CwTN6QCWiXdh3WklGxVE1Mrz+a+t25+gKGe5H5Sl2D9/j8uoV7Bs1Ypn/shNkgrbirYa91AisWQJ
dLTp+8keLkS0AaXsTb7bT3mQSO8nARHbcitBCA8Ud0IW3DAioGgPSPw7+dnd2q7Oemi1gaxYS/Bd
N93M36XLPczEkGvd59DfGlIRjTZHclnIx4kEGNOxSbQG4doTlHaf8QAq6LV2WnbAAtN9WBqIiAhv
e5XMykX7Sb32k2DS7Q7Dqb2al71XSZWOUgEEkwgGRmRpFyjdqzzSkjzvyk9e2I7NzJ17XW7Q4BAs
xBMe6zRuct2IOkjQOJZ2FtrHUEhasxYdFngRYtoJjUP5trFoRIJw5PlgGce0J8X80VxAuPjazEj5
btcpkP2zXDadq2zu6dQwa3UDVZfNzhThf81Gj0nu3OfW/wUXWAwb1fQlR39hHi7rSFYE1jTLuWfx
hCkZVtT7YvMWhY04COBpmIyTUwlhxBFvqxVo50yHOlRo1xbT997fN9itmYhWyK1h+cxIUKQfq4uY
C7QDX/K7SzbiBw+bDj/i7jgI7XQQgni8JX7FEBamC27o1KQca5iNPuAgT9lyu/Wdkpn58vlNhHty
I2T2fylAOHxh4TN7eONfCbaMSdKyxVmGB7jAZHRwj8V2VlE4E1kdcVU6JJJrBSYEwtD4SwTrVAhQ
BvGYdqluNy7YeQzPqAixVwd+k5jmV9hYrI1EcT7cKD/5agn5aiuT302CeZsSiRQrd0Rd05bFSKrG
WtnW+IyaCO+xlDHL1Y0IgEd1I2nBwh64FAQgvCx2TwJTWorV/WrdprvEGio0ElXPqVnTgArujjbn
z0eKrBLRLsA03lhJxibUua3wwef8ajB12NC1aAd4L1z1oTey4U5722jtXS9TiVYSbSH88n8vew6a
U0EBZ1f7yJ5TZngQ3+vzkByMKclmtu6vAGETq/E0FtUh3a25O0SVBaHRufcKnG079PFvI3c2TEN2
KFhIs/v8zq05bLpDPKGA4Qr6OExj8I9VP/TyJZXyLXCsG6gC94P1rf/4UeZKNT5p4SHS9ZC7y2dN
eh0c/ZuarB1MBBtqTJs7C5FmCSpxsZ77+f+Ew/4dTMRMv0gSjgz0Wyw3HlVeCsOvdzpRrh8ttink
82MAreBTEdYJUtfcOjzaRPNE7HzbGu/TguM7loGV5MS8LXrEs6JmG3Lo+NcOxtFrcyVVx0dUP7eg
oWqGsRvki63BFZBpPv5n9hjMGYke2R/htgbyyCQGaMEEbafLLjqDbaattp7EjcC3tq7kfk4+8YlI
d8sXcxEvW52xDyp9zY3Dj4dxWAmWaw5v9ciFkdktlWRmTa6WBxzDOg+Yp7sy4tJ77wHtudn80Kc+
5hn+5FaP5q/XOEEWGA0/nhhEmih5Q0I5yuuFKebDS5QaztT+yFqGCPneWbEuRTIXAJTAUPWI9tZj
Cd2Zzn+VtiZ2IEmHJukT0DthQXALGVrR3keOmWdyX880yu/1E36wKaWpmJmDtealP5mPZFgnWy3M
3mJ+TRZv69v8wk88XRpblcviZQilw2m426N77i8Ge1P+jrSJUAfYVM8pbLaIMtlPl3tdrENziFET
hBSMC6cynnYnyszImlNowRb/hWGdUDJn3vet/VexYqDaXZuGQ+HVpUYTlLD1v4MhsA/wO57T7I2r
5kqXU2wJhaVzBJmDPay6PFZVF70zrRc1/YmmU4wUVOw1hBFgqLA4NPKIUcl0AZ9bkdRWgjJk2hH0
y6VE+/ifALFDUW6Lw7FnEwGbvvnEpNwRnG+ElPX54iEgQiLJ9tsQHn99o8go4+rzP8t0xh7ZtOAf
M0GLnwOHjYIbs0xrhIxQflYQ30H9+/N8mr7eDCnuvtWaedC9fnqv4/BBcCkOB/DRn7bFMm06YM6J
/FkeSNPG92TCFESHFKtH755m7vhFLo55B/HO5nfa5XQ796OhaUHrNuCU526+C4AmlRUEFUj4U8sx
pXOGUu3v0OqJgSdH77ACFNRHUK3a6z41bo1VhBL3f6qHZBH46C7XIZNijEwnFZmp9BYJV+gI00Hx
AS7Y3aiZo3tzR9ausRMfmokljSTqfhtX1ZO5lNQtd6014TyeMaOQ/jsgrUceAAQGpksMx43Ufqa2
4z5g8WQVN9NuL5zNWY2VodXY1Vy0/GnLYRszmU6pFleZz9Cl7TQv56bUsTo9Tgvaagmay4riPNd2
kMJAyedraRJNkTaIYK4ADOPDFTB13Aftl9KCx9wKyr9h0mFrEyqXkR5u4GqlKlRodG5C9MARAX2k
OszJSnoFwVDB5dDxNTxFUrcNS9i+QsP4/Slm7MEF3t5WRiWI8SpKGMVrIryORukwZOn9LYqaZkqB
CV7mI9omx/rfVwc07J9GiL8SLbjg/srNiv4VBd3Vst7OISoW3yvD0DCXOmWwLb8agbecit0UCb93
ML8tDNHoTA42D1MWZmaF1zF7bF7Vqi/aXSjfq6+21XFx7TfXTKenMizaWJ8hdRp1mvL5yUhDtDfP
+NWy1XBhSYGS6paTolPtB9r2gHTKtPra2HvWzBw/t1ibys6TuAnuOf+i705R7RqB+YYJY2stl60U
iRXkqUs1SremY6RD+hrTtEISEAPe9AU9ZAUqlPDFiagLCy/oHEQW+C5J52Gp4Vbhh9kElGUN2VgA
O09/kIdqy+4JxkRWd5Wd/WPDF+Y+zaS2JXXefLLxvEuX+hhRu7tSmhd469pR5y16yhl0nl8Y1RBF
Z+76F1/pZ8yk1FMuaSWlrcUD/dtbBAebm/nBkdTC2ZmP8ztbLw6XiQBORvFwjdVIRMPZqmk7XlGI
3Cwi0N9MkNy110tCEsXit/zxi6fJTIBO8i99eugjsnIlYaps7gqU/g0WdsprsDPwtIyo18mgPNJa
e2GvzC4yzYBYfngeOO6o1KVMjSj3tR0AsMpyDSNnTOdITCdxOItnP/nWVkgxOY66i4sOLyTkKt7B
N5LWevp7LHj1G+RxRz3sejiGsdRP7gI+arM3LmYU0NYuXPpAt3ttgx2qsSly3ennWpf0spg5lQH6
YAPJvNWK4kZC4GvGXfWu4/863LxBTqFvB7PP5nOsTqz2L1kVwqmlGTp5+052sNu//Wy5THooOlW2
94fe7RlFsNCF0WjBC0ZxGWTHLQLTmfOoQB/q2TZLssvQ54V/rNNyOw3rRrnrGDz+ng7K4RxUdhfN
klTfrncvNoPqD99y8BIpFD4z5d+UEXtbmtKfBWxwKvqP38z8m3w4HAYkmKGWr0mochV3ZNBNO4qh
3FMAK2el+4hJl06p+0L54WrWLY66mP+nhbuVHlpc8oboWZNnUufuf+fOPqZTgxdIsa6387gLQSFO
0tywK/ZP8y565a8oS04aKOiVY1s0vSDEfHjFpIXs6rVkMYJ8l53qawbkgD8EY0XvYDdaDAK6s36G
yeYwFgi0LwzzhqhAjCvWuCWqNrkPMckBiz3kI9WMBn38iXw3NHQt0ZM2M3RLZFfYseHhxuMt8gRF
R0sGiWUkYB/60xSOnWubfz9ZQdAQsI9ghbLozRqWRZ42Q5fnbw+LyTkoihtgoqnJJ1iexMpBWk48
GG2uFTjvd0Usvi5SSqc5pUzE8a0jWJxJWl7N3wvSQ5I4oyTsjeH4Bniqw/yjWy0szpcTFe0k5AgI
Svps8Z6sW1vZvXxyNhls7wOPEIzUetGQIB+05tJMmiPBPmwas+u1uq33T5jEtpxoAexfnCyOWtgK
cDhvxd6cBguzN61J0Xs2+34roCh7NmrFCCT1QY3kfCBcaBNuafNhbMD0os2bX1bb98WtTddYMMiL
iXLg+pDyZLLcq/iuLYUlvB5FXA175EFEvp4MRGQrFYP5AQtJUc+00YOm7CPEnj14ku32nwRdI1/T
K3W72B4cFbLbMcy29nslOvck1N+v3pJ8F7H6vcpkXbUFjfQBq1mVsoshKztK6GegU6hC4PgIADHh
Y+fSNSbNwKQTeavSJbm71gSN1gtmTv/3Glr1m5viNYmGsLEAuPfIBYvSJAVG8ImXlYgjgAfIjQdK
3aheZQSaTGQcFHRg6FVaeCPnGuGljrjRldQj3k3Zm92lUSo5hzeTJzKJxChJVwCUxaFy5nG7AxA0
+fUO1E9mE49KXgybkeAgSU+pGwIXqG7abCEXN/8XvPRTj3naApvXwoERqj1RSidf1prYMBeeFw/0
pW1VGH21+dj8SZrc8sWbOaPT7KipqF3+racnR/VoE2ARuCruDOTt4PiBeArrNFZBcuKGAETi1x0m
ly5SIK5yjyFWE5AHXAkXZdwX8qNiygs1DDCa2d8k/RY5M26PEU75b+xGk2CTVMoAv2k0nDUnjiT7
J2sob8mWEopNAu2Gg7aaa7Zhjpwc4SHshP3lbHHKIx/2ph2++mQEBXMUh3KVW+L55hW9bQZZj0f2
LQ5HizurX9eztt3badScV83bfvk58MBkTAVTaV6g5sVFE2aThI3ZsmqSECOKwjHx6JEcAaXuz2ce
l+GVoGxqADIlqspumrozNPIlnvD60RttDwpchi4by7blmH13Ie5Ku0UFJc1ZqMrTS/g9ac/FOotT
taB0NJGsRGd3+wbH/OL1FnzB0I6kcOTnpYc/Flfy6SCb/BJ6EpSCh/I9TAdjyC98pD++ON/wRAwO
hN7a/euUILWFR8SI1tix2smc/kzX0d6YUYTQ1R3kk/diGCD6+at6iIRXqTFiP0j95Vfo3z5IWcdt
i0XgBqaTVA75ikdEJWdyCkPHEUGnjBwjRk1is0F0q6XyXa4xJu6H3LhTXk99UDhhcorhxWHK4DQw
KY555244fp0BH45X9WYCJMjBDNEvFxBCDsWe0QP7DNoNpz6cdUZDViVSESAXyVBvML2ywsOukl3c
gD9EXutdkIe5lkmIvWUM640u+MwYF/vc9FaUV6H/FCLs3O/m5u4796n+xCWZnCqe5AJGbsU0FSTr
rvlwZ3DmFAdWskj822RCPXVBw+jq1zUBpOrgW7sCL6i1wMUc5vyNtCjSeHdwWoh0W+k2SA7muTWS
LwT0+gTUE3wsWaI2XN9i8GadO8rra/q1P9nEM4mGHqkNR0GwR8gQCN+CBN0j7on5LFNHo70ioNBP
A3XjB3KaTaVwNCEzF58GS2GZOaiVM0QxpZTQwvjRt6wPwiUnMLBV7NaWZ6FaVhx5zTCCX6UP+bAk
eoGKIwV4UJXOJ2In9uizSG1COCj8MZP9cPk5evPDRI5NE0pb1OKyBHIjvOoveupd6MErVkbM2uOJ
bePHDP2jaFc4VkysMS+3oRBuq3G8rcP3cOVnIDQt2kz8KM61KoHB5736XVMnZZMGotWs5WAQ9bJT
mLIKuQmox+LkLI0sxmtcoDeX89SYFTE8fmypyamC38iq2+NBHdq7gSwLBBoJgGaRfXWsJkscqLRp
7kx5YtBEgoZ6+lGhYHe9te4aqiNsKZFCwrNIB7u7bJAz5haUw1LEA+qoddcPg3/e6wueCI3wkZLQ
uTO8dwjWy7eWUsibIqazTJAU21A8/dpqnnyvOKTbePAmtuzO2jGcXArwmdhwqpKZtBzLyI6LGsvI
i1ITdsLj1xiik0ugN9wEUeQOn/3WlBWmHysyQlAkF52aAVmnzz2g7KJmXBlR8kJ1Xv93aVm/Vn0e
RSrYcBJoofiN7pgzxfJHjoIthaKHbZ/ICH5kYK1xoCRNUTFn1P2N5kzRWTQkZ4IOXWHoKoLHyBOR
EyYBPHs58UWz+DLAjwg7s0Me5cYBUABT1p+LiOZjKrdGcEZUEoPWTnDF7Rea360fe6hI0SwCMsBg
fOw7l0vD9gElLkdO/L1ZpOwS1RuLQSLLBHKdpohbkHrsklaAI9w7bgZfrG4yHYaZmt3eH003ykzo
pbhHqTe4ojLm+F3zmwyAv88R6fvyiu6e/isE4+NaOkN7ugFUYEdLrMiXQ+s2tqSi0JXbVqLN9akx
QtAqbk9yCIvkKnaDk4GwVypD8gnwob3Geoompa9FULFXGtHkGZB2RQmMjkKrEYFWfvfvhbl1WWV8
boL49pWBWTJ7+kCosx4Mb21gd4EW2PKdcyk2t4FGDko1DTxq3IU8E+/HuKs3hy1ImKs4DWSu8O6t
7MHBVlKU5A3hlsdWwlTpn8D066FnWpSBKZWGRQ+fSC3ojxosNXvy0X6/AV63yFJCJwWtAHmRewt1
Vf4Qcst7zISZ8E6nGZeBE4Q95LKO9kaVyvnj8/ISL1JXT82zluJAfN/n2HShXNlcG/nssILwnpH3
cnYzy1VdROZIMajLfRUNhneIf4TdiO/F6BaBxQCFjx2s1FNm0AGbLOgWA5hBjXClw04HuXVzvuIl
pB9i6hT0yQgmpvl1pMnT12WAVe/7AhCYBWE3hU+GzRUw19T6F9tqsKYr4TIm2OtabNTtoqwSmqZx
mId82L8MJtzupQgUO9uN8luGJhpQYzlkkvQxTRMf0Bmh7ZxNo4pv9aqeflY11byTLBQS4yH4Z5V9
UBpQkMFZfDK/sfYP9iAM4xJNSqxPWBEbnhu0qUeSwHgkpngBLeKsYDtrGyv8KPV2u+ugIKAOyZs1
Hgg2fsqn953kNWwN/MIRuBELq7Z8A9f9i1HKl1FCWAKV8sUZfDMgNsuG2STnanyI/MJJCdQ4M4A6
T3WpUmgE4nX9BOeNOEMaH/T8LvTaZtlJQphILhNGGLDVSYpnNcb8ypfR5/DjqeKq0fSPxlrqi/QX
tDC4WrmuFNzZrKhbCXhFmpuzIzDLCelJ9yJQfPctmTUJBevGV9WeARHluPkXeGU8JmysUCEOHkGj
nZ2YfeJMNSwOl1kMebQ5Q+QAuccSKI+CoA35tgtEXCbVVble6UXkpy8fUhbdsCFK3r6shYd/nVVr
YeApUWHpQIwI5BZ3pM3jtsMEa3q46BbSkyyRV3PTHoAKR6dCR0ZtlOUkw/O0FPjx5oElq3idaLNI
JggMBAeUitwzL6P1R6bnYeFGwkHSdy2NJyGWFb25kTc3XiqQloAKPtW+T6YiRja1n7I4rSD83duy
S12nOtX1vnCZbIn2pFgJofGCFzElz41kOmpz6in6gznUwDMCzx7g3iptBM8v5ovyK6UGgWG8X0wp
S/OTI23Z064yEwT7H3RCGRSrvDrqc3p4jnZVStA3cZ8lH2/cDXmaWGhJpUfN+9UtdP1BnxGm+Ja7
9e04Dzb8X0KGxkKA8reQnHh1B8GbAWc1xGXKrM16rs7okgOhHQ3saows721MinC6z+NXDziW4Hg6
2VAY4KN1XWE3kVo2QTHaSdAsCe8W2OT3hJUEYzy1acmsjW2KypC2EuDYIviCYPsBOT4+uyGTckdK
a5Cyn7vFOvL1iaNA3kobPL8JfMLngtqCwiplYdmNOBBVatE3TxLm9my1XkYlUNXIShR9qiCOP5o8
B1Vmkd/+PZp3Y0GgAgNHFbbcDN/eE7BYhXkZVKK/GXDvTaN8xZWvwfXfEyXX5YhlvypYqCDtzQpV
rIpG3XoRgkydWdhdxwK8SyCb9yjRiXTUu/3gA/q5bNbNPBMT3bSbYYstz+QATqTrY4wYZ4sX2hqw
meWAy7/XipEM8WLXRAJbGmtqytPcxvr1DkQXXlG9FzAH3ItmTkNIP6Nqzs/CFgug+BHmhXPiIqab
Xyg6aVan691hBrUFVKc3JmG8kf3c2vWJWS6HPi/BjnUwA97rrU4uS9XeJHxbUxT8MRjEvqj7oQAP
Ez8SdOVKGFbc0CoOYwoaLUcDnKcBYLIW0SksKBHKOIu4lGsyVXJGzoTUoYJKBppzIHxtYWgUl+WZ
/AmOLFVhO0LdIvlb5r6zIR/yWnZvipRQfGz1yofwSJwHnzZO7RdYFbY7HeeRcOaJPHnGAUqUWlUM
SgWn/Mml1QSzvOulWiS4GCZKb7b6EhW1jujjtIDZdOnT+hUj5xUo4KXiXC2SFEHfwwra7+zMqhC/
BTBnVHOgB4Y1J5X2Ff0jnQJyusNfAfD6vZdR+7d0UfuxY8pXuwhEFAgyekmz9eV2e6qEps47am3I
uSZmbUlt3cVzAPYfE5OU31csChcHel8mun6FybB+xA22xR56VRF9QToL/xZoEYcF8+Y0U8oTN6Lx
xdoPVJVHXSXIZUMeaLXzg1xTTrg3BZkADx274vdEz07uUJdVF0f6zjzdEBqm1S3fS6/wNDi4KO+X
XISvucPVTwcJ49A211yqsnP3PvdrvmaS2AeCzIBek1WzYcNuEcyBwP0CPJpwVaguzOD/Wpi7oI9t
HpXgivr95L75kEa0X9IHfovo/MG6xnxLr02w0P8u4IxmQ20S0D2wx2JQ63VT1SOacY+o7Ur+G2oT
ZSqowL7sA+BctZTYXyLe67DJTKM4TW1HbNCUYdDxJ82vutfK5EP/poFBDpAlsPbUY9B7tf/Rfj4Y
30D7MXcg1pLJKR+cQd/FiCgUQzNxjkxTythd12x9Mh07OuGteGxoizZd36J6LyIn4nofS0fYmetl
LOHCPBNGVVo30XHtUoSrepHTAZio8Adq39o8x7yMK6DAWk9YW/F5O28ZMWUOFE3Q3vBKogZ64Bz8
7pGkg5KCwwiEPUvq9xEzIQ4u0KyQA8B0zhTqGxJc9rORBs8q1BDODKzPNK55P2JHz/C5NUzeI/zw
J/4Z+Q0m2A4qevZUqvzqpvQzOXaYDTbLl3RR6w4Yvu+jQDO0cCJIVDOrwb3G8DdMu42outO46Hpm
JK41o+Lr6YHChZ/hMtUSd9gq0e4qDH7Zqf5VKkwn6icC9P549viIwnAI/xFO1W+lNUnIIEDHO8vr
MmY77aToXR6uc9qLIj17r7L08jxO3pf3k1TnrCpSCQjRkIpxtuyIfXzmtV1wbESJ32L/9gURMFxX
NLp5Ao0ANJTy8Dyj26hF0P8pV1jqnEgMAhtclkXmzkDuapxGgEFnLLLFXqJBS2FRWur4lQjm+Gj9
ZXKoE6lemyXedm8WiMP2VUdf6kfHqLhhoWrvlVxaSKa8+Du4fm31yY13Cd42g/DhgnYeyUNVyKr2
kQBvpBjrOzShdyHKD/0T8W7NcNIfDI0fsfrdQnwmjFsuttIu4NUvweksFCSbs99a1MzkNjMBWHoW
Lkwgp4hzQzECvBPRXl4fsNyJYnlk1hMA+jfNzXZ/+btZxkaB/oxSb8PfuKQ5WTN5ng4fkU8f03Uu
lqRb4HA8EO7daA9n654FBG0QD883s05pL/uVdTHz4qzKQqLqMfXw37W28xfOp/g0/KfrV+1lKcRF
tRlXUjgV5R8JNLzvO6qkUAHdOFYsOYNA/RerTZQ56FQCqM48RuIYKyvzbzqbvxCK6SQQ0SXtp9BG
uooDGB/YWyEb+KFWap4zRJd9ir2zBvwkwwrEbC3TU7dP4F6KvEQgqXb0uak01iJXPLQ5kqO9RSF8
m8RciDoT/KYhin2jl8pus93xBxK1+1kVXk9j7ccQT5+9XE3cEXZfrXCymmssb7I0w1POC7zLLKlu
urlHDXRrCHoWKG6zRdPOAazGRhCqXQ4U+0DOtnkEf0Kyuq6dXd65f1Iefd1oBTNqbdJmC4olUjEl
0MaKyKoXVJTLHY31G1c6QNQVnS2vOxTrFDJ4E3OJoiqnm4Lvv1hs6qGveLbWSVTiCuYWzLeX1Rxd
syE+C95JK/MV3lXcffalHpexgX+TOzvfLWxwVOD70k20c1zHRZPDKXHI6Jx088paTgQGyn5KZNEm
/kySjxs/wD9GLrAMGd1da0Vw+CdDuMiYfANc0NYNJhMlSxJPbVgicpifPiZL1cQmTtoy3LyGg847
d33qJQ+vft86yWm029Fe/BCsE7FgZhR8iNHhGtlCcZqWsK9a+S9i22IuXbcXYWc0XpBZLOBGnOqL
ipC0rotJ0r15TuSnXcWtobmfYT9vNJxje9M7+aygNjkHYg+zVSw9qco0TLkyVfS/VxcwhADR3+3N
a+/kGAfb/yxaQKbtxm0jlP84QSFbanmlqyq2uwPeDeJLtzgRG24V4BecDh8O4n2xw/tem+f0SODF
LO2D56MKZFJ2FPa/Wn8av+uhqNcJxCyjXkCvuJoHA+KH8H9t+bDvU/T3SloTrWiIv62/Fw5bxjDB
pfoo0FMcjg9jNrm5vtXyf9mGr9xRgAXoKQqO0fCzUsGQDAPwtBqqWw9xSKFKiJ12L6GSibAgnlJj
naoq57vLEoewA9B5R0GU+rJA0/gXeQZwqYPO0wAamzCM6/unexiNFvQ4PYjQ7AJdtqJE/qlQCKYT
/tAxFo0G8AnrBE05JvQHtCu1P7pSuxZgr3i2zYR5bJHJzRt7YtZiRIou9E8prTViEyQT1IGvzTb7
kYax/5dLy3CHlLuuZKLHpiETe8gzkDix2orCRID8gwPv5bHc5xUy9xLuIFHJVNwcg/9pwb/ekSar
oDAuZdiFvwlm61LnXutTNVHHtsnqwFpJbR5DMIC2kKIgKwq93XZEGFNi+UPYbxxRzJtXH+K4LV4f
VMOdC99sL/9nSWBUPTZ0a4VYZ7SrHA/VniAdTpK8xOxBbn0yytH9vIS456lib0K5IPtbpa+IZHIy
se6OYQ5I5WHWoHtT8oILnoTlanCoEW58Ju7tgaUoDHXur1CmRmUun8jWM9GCujPfUE2MiU2BC3j7
+rwFQeLLln3bA+fv/KMZsOZ/yCFRAGrB2ofk4ZxdyozVxczvCyBNDuF/zUec1yNHmC3yk4ZD07td
3mgjKg8RvQ3KcDkO0LXKonlttb5xbBHGC8fZ4Soyw3QYDuZqXSJZBbMRIMkF7WG7tJJqNHVpVAjv
UnzmeqsuRcaVPDHXkzO0ZplyDq+3piZhVh09GhWOHUj9W4H9/QqELfviKjzpEDaeRi2DLDE81Qm7
WAG+nY3zSRegoKTu5Sw7ha+rUZVlOdEpCZOS2kQPpuBArVoL04o7RRSUSEk/w8ef4UfflEB27E0+
Qxefz+bvnewlVGpDmzTYxXqLtP+re7tgmSgC0x8dZdx7ffSlvYKF0YE/j09MaEhmPCMyqcWzQJGM
6UDocd5zd+CtqzNiSqMo8c13FR6tABxHG8rMQs5H5NJo/+T2lpWvyurkNaoe2wPXwSPJm1dWmTEB
qccoDLI0HNZu5jPRg+mBtwGeiB4cQ0NgaYxaGlG8lmeyeVEpkd6+4u73ue4FGKZkqXXpnOytjeKX
EXZRgYqOjZQDy08IRNeIgbogZAQ/RpvHM9zchksu+KxcQolSnCr598A5hQujg7zfvUQ5eCPcqMcV
BNacOR2DHvzJ7Jd/BHaLqk9kf1jDXTCM58aqA3/vOmRqrAWy2pLMwEgWj/KW1aoaDDg43tNF0aNa
/Mq4surqHZJtyxVmxGr9azN+SE76o0/YBnUMdle+VgeMEqDlq/eJEZl6ma1loDD72NF333TdeUp1
4Sgw5c51vaY0r9JgmiIkGqLFMRDlpsKzwe8nJ70L0wrC/RbRCVMLwUP/Ja/zrC/16mK1gQUs9YXj
DGXle2PT9aKjV5ce2L5czsRYnjD0GCPxucrqOtwGKSZMAu8klRL9OBA7Aq4puCZ+lP0t9r6AuOWh
+jGHV2DNPJDLESec6uaWQRztF4osV7+hp0G0GTgZz2M8HtvSbMPNtt64z7p3Twnbmrf+bg1eF37J
Lt+9tRrUmUv+EfiUhKsY2raOJWZ6AJdrYwgpru0RjsCLkWgwP9PDGzuOoXVNiEopcJiyAzCMVF9V
pvfw4jbn//qWiEvazxjXgRZf3AdTqeXn/JBm0z+a+Rwsv8SznyW13Q/1hRmS+gfY+J3kpUbrXst6
GeshpecTlyGrVVBeuFV7yaUk/LnT+dG2d20mjpYV8dy+oQxBIvVFPemAKUJDH1/ukQu1+WPriYta
IBAvtCIA8Rm5BL/BdjtyruXErAoQXseXgcjWc53A5SWPGwkFki8I5/9U+0+m4DOzJGrhSSZ7/qou
OgW1Cbi03JyAM11s2hox+F2ft5GniCW+EjwCFFR8Rj+knplC9TP/WurBIdZ7m4TZJcBK+dLpJFU3
pbhSmDc/uuWg0pB2cz78g5iIPkESo8jmdjuSJG8NETLsVyu2q5c+YIcTIoHy3+RZtcxBeCDpAbZ9
GLRoSzrmyiKBkAJnOr1wTntp0H3DP70Axb9mTbKntNU9NclBIFGmLOFEhyCZ51L5jCGk4ADkj+y3
8qQitHcg75Z0IjU2QR85CG7exGk6mpNA3lYscpcK9d5YaQclDXkZYyprGb+FkCwBvh4ZrYpJ97RJ
4aL2s+JNmzVWl8DS8STCOX5ezMTBGPJZjVwZLucJi96/PoYivTjbelv67aqMo5lkFZYVdGCyXrFy
kEnP0eoCMnkszxqEzY/g15+MKKhseXB3+SN15LG22whKmSF1JWA8UKqTWIzUfKs+t/0geHTf9vye
AdI4vp/x+GewLsMhoVQKIGEqr6r96NT8HbNfbNEFzu5hm2THVFrWE2ZB/6uYuiPhqwUGxCtWkKDf
lKUusMOmi1kOWQxECQ9szGBvANs42JxwAugohKF8XweMnci07Mx73aHmbzpZAKgzmLvCanaA/LDs
RH7s5o8qUm/6wnd+75tC8D3y4rpFQcuFDnxopXCseDq2BXJ38g8ms/yqnXjf2iiYA8Ug/HtOzB2H
1EDSSKrDRX0ycFggHodztwvMLwXqy4tKFhffe9BpvbulJkgRvfPZ2fGcc0aY4U7/RE6ym5SjT+uQ
Wa9USrEGWzAAwsbLwewUxXCvvYbrYf7YJV0q0/UlPAF7j6sdxiqgZr58BvO2L/qnRRq3M4HGkNl2
1uZp+L5KMwf7d7EzBThnj8OYAboAAyGcEcJ9cX05jqcF7h2/DrLo0A6thP3ZVF1gRqPOI2RGtS7F
d70dDyYI7qV5QaLf+BiGcDQ07DKrGGwXkdMG0jeVHVUXkaRHevW+iK7r5WLkdDNux8tjCj+c02f5
znYh8LVk6KjJY49zXSMpjG0z8rj6gGyPD0IpeZIk168nsJb/oOQaY80LA8w0sQECZa9ZRB2D36EC
7/1FcplBsAmDxzqHAJmFNK0F4ztm3SmNs5oB1Q+xSOrh6opKYYMI7czcC6lTeHOJZVfmDFCGLEeS
/mW9818jmqJqDdJU0Csv5DPreXI+7sA5hrMwT6fUo0GCzUp8G8D+ObFFfTmVKc2z0wOzqcnRelvN
YKuh7Xm2KqyItYHcqPIbTQdF9lsG5YcjSQ/hPswevLZVeusb/I9Fh+3c7+whuUjPIEdddrgYqHvp
bBQlSVQBAhIb/LhPgETBJsuKWss5VOrd6pBDadBL7Qe5ufzL7AcJUvbaGoYseCI21mDxT1PC5gta
WFBCRGe5bWHGkmLulAxK3GFgCHHOHGRa8Q7AJ+8XJ+vvcQRt7SEjsHjpjcQQOIgZL4YPdj4C5NDW
ZlxA/JtAnyAOncdVmwtO2gDjIIjtdrz9MwTZkGkhLtBi2iC2e7tU33hTeRWMefi1FIEqwo/RM57x
OvUwMdlwkP6rUbmpVUYAd4PIfM6UKn/fHQWrpPCXzbrjw4XZzvvaYdD29/r+Ym2Z7QkIljxW0+u7
RXCAZrHp/f1PeBsAES28UnTtepbtViOKqztmk4+LGc0GGFazRgXQxDeD/VbYxEdvMq6a9rTN2+6e
iPIQLG9ab6HCNT/XfdA1tIYIN/CnuAlHmVHvnLf2ua9uoBfV9lZWjjdZNOOLFwMLLetXvRir6ktT
WIp5mN6p66wUObsysrwD8OvBMI51A7IHuBhWn8LbzpO4m+XP2zd8U8t69TWPEjIp++8JkMbHiva+
RINokcEoBGClKh33FobT6E4786CMoTJ22Yw5E3HByW7bbPFJz6B2AgrC/NHhEESqXGbJzzfY+gHR
hvP2qQ4QwsGdUy9VIAKm/BrwbzWij1oX83hHO6QLxZ2mV7ZBavKlxRRdMpPF0kII1YRLQg6fM4Zc
pYTbvynU4QaW5roJjUHc4onebG+PpK6uSLm/QfPqoNxhXz/Yj8QZRMh7mQpjwjzG/bHOMVkJJEBG
hSRShUSyomE1goUS5Zcdz1zgDQ8ZBwUOF53oOKuimSmdjhxFrT9tzFvbiV+WkE/ypsCE5k2kWPBq
guJ+3yhmNIrxlE+Rit91QwJ260lk/zXqRHhu6u4/fq/AS0HE2jnZ/0DgxRl9FgDAx0E7I+MMG+ir
2QyQIAUfS75Gmi8GSDuG0l21WqP8+h94LcMMStJQF6rNWLeLVvdAFdeBnKQt+0IayJnHhsU5Nj5X
4F/Zj3kkDuh3DmbAkBy3HwbSUYWtqxKJsIozJ8XPgGm7kTGZbAr5z8yms5cDaNthLtuS6k4t26SV
mzKuT5ruMPuNgfxGpasHLA0iQZgYv2qSmwHFQ3RQyu9BIJFLSZcKUNZ6ecV0RxmDBMidI6jI6B/w
UZyl3sAZzqns+dwpJlb3eFikioZt+YqQWX8rCtd/L7qlYV40YRvzyyQUcopscSfVYl0TowiAtGl3
R+4NyFNma5qOa7nI5cs2iJ4emlvg/duvbPC2cJgoKVzn9FE2BSmBa1tdtA8h4XVHuxPfQJPnBNuA
HuQjVhfFUsgquSDrLTSP5AhEjCVX8wRhZai/LApZe2/pG7j0KaI1AlLwZ3nNFwGAsLrbEy/Cw9Aq
HqPmZhv1DL5nPeN2MAmsbr+HChCWOqFXrHIq0QniUmCLfmrAgzmzur65sPEH52SoDdyeUOByUP5P
Yn9AIAXis7BJT2Lwzl+aO9JwwOxouhQmyVasw5c5Y7KWHQCMi6nJ+WBdiSNr8irVn6GQd9wsS97U
jNmkVBsvSLJQnRXMEz9CuAVEpKBEukKQ+AC41T4mWCnjwmJjzmASuzgG9JD2GBQ/+dgO+8gVjQfv
pJmf0SYuwahNHJNzsYQ1pFkMQfZhiR12HHkaSfwDSnz+OUUHJM+Cw+XtdjYXATzIQWcEaZJFZvUZ
mkHlYtJdHg88Cg4pHF3DTlyg2+6ABu0yq402FyvFv62fsEvqpAlRDg1fsG+dp8cAVN6PQqkuzr5j
WiQ6i8sReJSreqEe1Le/zFDK8oDkGgVfCPPdisNwEbcZc/iAX5yUdr8/G292U3NVxzXzrPelw9qu
lNQa+9GAPlc6bh/Yat11C9W5yDT6LuHOfMeldd4mTkAARqxgsatLqfk7z5kpDEWfAARo8XgoSXro
9IwKqb9mZX7ffaJXoNypqRYomt5ch9gtoUg52douUJPP8On/AezH0dujf/0i1nGi0boGaaKHuRK/
BbwUsJ8akiMWl8tKBHwKXtuGgBw027NQiUmDEFis3AKIEp0ODQN//1E3PaA5X8+NnfxkLGCj/VsM
A/xM8AA2d63fzKtI3rCMkBr5VuDqd8K8rdv/q0frzZOY9m+nj+8Y1YQs54EFfBqsZBfP6b9WwewS
+xClAbjWt4/fUFWND16wany2L73eG7qlAc4njmZHM0N90kG+zRml4V331nGxpX7gQDg7N52hyHHz
+VtowIJC6LDF/ZacaDMyDgBMGfIqaTlZaJjAqDJmlBIAfbF+i5YTEgHXZj54aWWCOi+/9b2qeD+v
wj97fYwTqIm3TvNBJoEPpwxPxqCAzfxOwBUxsCaHhF6eoNvR62yUBI/7CRCSDHkZeZ1nFUxN6pgx
DZBdxLuvhxOl3c0mAkqCMjf8m8ooTsEHdOeR1iOQQKX37e9WY1S6BDqR6s6vaT48J6ftP/URrEw/
s5bEiNWC2pOz24YsoIxLmBfg4tT8dBBcC7Rk3xZ3eP/7NneC5zYgI7xZtNc6HsADPjirpR7Jd88F
tflbUfLlYEzJyN67IcIzbUjCI7KNn28lO7Om/nYdQvsy3kWi/LXuXnEYKB4RW/99Wz33ZwY2R8Px
WGvAbFXe4nwpfcUmMrDIQN6kDa/sAii7c1utwZHd5q3LcEaDsqdK7acSSEIdFF9C5iTK5O+CgMr+
XgQdOEoFtqfzqVvBpiF8Cyr+TZb0RJFJ7XJvHvYO4tPU/GxeMRwXHE6Pr1he57fGkjq53uvMhSXl
XaAMoqpabQsPQyWX8/QhnoQDGSh1UJRMPo4eLOmN9VH4gKDKzWCZ02fqMODNgyJOn0iFYYqY7RXC
9NMp6bSMWUsV4lsIzq0+kN6rTrOcIUOs//aISYcLss6yvMlm+2wTu7/LBJF1dtZq64k84VN91tMj
UNxT4DuKu1wpOjC03yBRXmh023pzknEw2aN0HDplPCfou0VLN2udgxB+ULHssTg78dSbEjJjGLUs
6BOoGx1cIxVCNT6Vi/eDsx2DxRwSOYTXOVgQk6T7wxBMa2jCh8E/XbKmaybvnFJYtbS2XTcHof/u
yYOuw7xEKP5r0jheOEIBjHhqdu9KytI9Z0H8G4CHBNzHh9V7q2jRgNl9uzSfIKkEn25vHjbvWBwi
01/lWj1lu+QNRZ2xVgwbBZ903inXAz4vFtkJFq7xfg/PQNZEltPtV4L7jhgv2+PKPRNaJceEvrzo
EuGov4mihu7yH/F6IhEhdZ/lcO7YcDOPbSXXayv6xqIaG2cShI+er3FuWZxXVwx90yMSHam5M8QB
LnpdkdnJWbIeKviPwUShROqIX79SCbcbKZ4aUej6+9v2NzDEiJHioEzZn9tehaOdJyvy0UopVZq4
RIzWebQjsZUp1ENtS4lrwBBPnFmw9tvpRH9z2HO8DR3UmE+QeoleGwJ+J2jA+6mDVqRi/g4cbRw3
zW50eSuuGZOXbH7ZeuBL2hhtOQcVnk4bizfIsah+H0nKpHqnQ/8cOqE6hpdekB8yMRyAo0GNT/94
+wz2ije6AxPb4lJMMRAhrHIk9Dh4YzJLqhUm4fqaJhign/oTxOn3eR3y58vhtzLiUWJpdLv24l8f
bnJqvA37PfygO9azFnhSvN7xfSZtAE+FWEbFZ23ULCOoAP7QrqTM5KisMSipjW4gPVZf0f+tL1gZ
NF0rmKor2r52i46aRmdMtRy1vSgXL42jzxAFCgylUlDBRZ6Yz6RAVWmH41QbmfQk7sWQQvKIkNRV
hI8NxHs9ULneQ2i/7ugvDCEylI2nScK55yVAmYcr7lJAnKtX8xF9CBDAPHMHdCKEnDj+GOGJUFF+
ByHZEm3/rexdfuDc/bnZngPWxkYy8KHFDRArP2LwZJgIsYrrnYkr/s8fwIlrUAey0ASOfz52VhFU
YqPwHk/gRBCntRo+puZ+KRqb8DN9j8bNrX0GP+kauWXhsCNaDx2oLjnOURhH+UXfVXKw7vXi5Tyu
8Txtxz6b/I7HGcqCPm9sEZewtJG7aQKK3XQbThAcGeV/4IYSWsKPvy85SY6wq7hb6BjJZTSaG7ZF
PwWsQik2T/XKQ99z4l5Ob2QbPH/PPJe7+ZeOjuIEKqBywubHJUNsixzuxM6R6tepicP9iJu3DAhB
e0zvCCR/7oycu4/+esT1GCTebLh9/Plrb/fpVNJao/K6pmtz/AXSdHXiNal2EHzuadmJdyDLVUVu
gHjksKeuH72Ctej6jkpjYOe+vOOqqDG5+b6+Zscf+uCcqSU6L5D80qtzHvbF0DmAnbdFGd7NG2In
bcvalt5eMhwYLWW3sWl7dP7e+HZXdwglZJD9V5sTyRNasjPb80uFcK/mGlMUobKK1YbO+zn+4eLP
LgX/UayMqWp/1QNJA0tOUF3SNCsN6jtoLPnqpFbB5uqOBWH1HLekQzQe+WPyej+J3uQvKB+mhOx8
LlPKSkjQczif1GGr+rJ04Pu67basUOlRlzCRUo88hIYclFgLK48zWziPxsVshM44fOEEKRFuDRkh
aTfP7AgRa9CQ+5N8t5JutcZ/RBVWXrewefQUPVg/062B02m6Y/Bha/OD+lprKrl2DydRmtvoRo/p
CTVdmswUJCuNx5vZuzPuPFErytROPDUQWXf4sKMM7FktKU8/bCIvudM6FLlRtnQ9PTTU+Uy1uUVR
e5ZliNouwtMt0TDFjhH/TiiYJaP/s7683gWpNaguqcHPX+PKVUALbfPjODsWnzCZ9HjO5MY+4yHi
EUPlwSme0A0+xapa1y0O+PV3ouysDMgQ7EzGgfLmSFEvC5p6TTQf/UJWfHsjnY94vCFi3sWqRnUL
ZJ1eiDyxebgFDo2KhSm2HkmHck5ZEMO2D3RbJTO+1C7yhtDxGevyPDuHg2WOuf4/uVLR512u8w98
FPIDfbiBlr46VyxeBmrXcdjws6iCm6fc3fxqjbZdC7A65cX/MLXXRQivzgb+fiv6ta4Rq7LFS95j
m5+Fo00k6OEKpnyPZqI+0JXE8pCkq7QI8WbkiT/RkZ6HmFXW/9MAU2SxLKwwbItNaGvSe2a8c4Ly
/ZKU2C/QnY5Q8XhcVcQdYW9MXufNvBzkBG2Mv+eXGzocb+RunWNi2KsjZfNSnpKAU05LGQTNB0I6
JNoPU36rO1RRO+5gZD6cWyoR6YmJRnIQVD0aQpocMzB9StnIK9ErCEso5AZ3NRlGQjXEfepEoez/
hqZC6d/kHbeFE67ld/mXKYIk7wDiHCXIsi5pua8zGgWsf3rs5seCXlG7GybE/YimdYnOfAlS7aaM
6uQJ60kpfwQ3KFEBTr93iZnBhVnp3aPRSOOXXjCU7ajSSCXFCRuKBhkRRoRQ9Ly4se91Xb5hYrwC
4IXwHDQeqh26PdrBFxWbrdI1TQjTutW40Px+ufdOyGWDvBOXXPj8rwYdb0mL7+MkmjrbaP6yfe0u
QrNgyIgi8PzKqqnpjFY2f0Zs+DfIrZQNSihkxWnAyr2ju6ZeSRHD7vyAbPhGcHy/xpexanSY5/PC
w5p7oJpmL6RCWaIlDRCSv+1CoNdlOpKxJtAvHqcVJ1/D+fwkfj5OoN3G1+ZlOZYi1T2gCX2tAQWm
PnlOI/VoMuBKxw9LqrdelrjoNygXPBIdEpzP50w/t0aApRaLvomCei6wxfLKAu+OT+gEPBlk6MnF
gowLr2FsD7roY7bcOsq/StUGIvKpaYAgRBo7c7iqCuIpbAWR0L7xT+P+FO9tA5ZDDfK3Th8+taI8
dR482JaVhHE0ctFJCcN9v0snXJQ23nbTLamlcYv176OXGcgS2fiINLZiXFiK7rrjsgoDBtDcKRta
AXRQ3c4yzGnjPUb3AGEQn2OP5s04mat7qdOk77VN6h0v1X+TKh1h6A05KzfA1vw88Sahq0Zqhq3C
hULns4yLYy7KKyWc+xZsQnSej63vMyNUkJSO+q4U8u/W/TDEYtkcPqNWOZIwk2tS7bNwNApBhu9Q
/b67z3KWGK6CSFbRfu96NMYYIIdkidIkdrwlHZDqSxrt9H1hjaBiqE0x2KL0mPiqQijYVr1QQUPX
h49pjBMuaHx4ZCc6jiGfkl4sVpjPZE/xIt62ujz4HFaIzkpGz+AAWmK6eMD56rKVMmyYiRLo0NR7
7IggtGELFoSEgcBpyYRzsBnnXhCLQSqYaJJ3HFvZD2/ppjHwJpx8+ilYDaliEdPVYCyamLVhXrlt
AqLj6eTAXTuhnM2b6aHohUFsnieKMDLaocSJCdae7yKYBbVP2LbSiDVJZB9R9FM470oF2cL4BTOy
TKb071vXj3cifv4Vq87DqDVND4JzCsvawTkqYYTa/zX1RItBFmiw/UCqVBlEzWMBREzVNr8hWNAv
NwNUQUuc00puOullx5BjUjylJ2zbVcdh5C7cuCpEttQHSeMv+DU0725t/X8OJrvjRb/csSI03UjV
dTFAgvz/5HPPLof15QiVRYF5l5UugoqVUMczY1XlAojQhecPjaKLjuBwfw5Hr9cvZkpwR3xaxnA+
rvI+qPn6IvPkehcvDipgnfkNWgGCCAGDAMcgVZ1tvCn1+liKNjJULmmRzyLdp7m4P8J8WBrhrhvA
Nbp+QQ7gmc7Uq5LaWdCFxvFrCUy9GqKT6glfuTB61mg0PEqW3IxG9e9V8Dayc1KTHHIT2U0ey8yh
BUpT3AM7Z6oKBB9JTXqfc3ZnXZJNEi1ZMtmAq8m3xs+YRyMzngBRXkJP6oe13tOvE+LJDax/zPRi
ZBFpnkhJL2j9azE1ATY0gWIvNUAKAcNjMtuOGx9lzsf10kn4Uj4b9JJE8qz03Og0qx2D7RThxvLZ
9ZigcMTfLUxVAYR/Oqk8LBppFyjodn+HuoSOS7icdAVqPe+HBcwsWqdTugQUmH0NxhBR4sXC+Yy0
dBmb7e//udUrTXGZKHricUgXV0MIhJjQrG72l8DHEPYEqRb3mGsgLGlQMbYpmzowwn++6vgwU5bf
mGRzgomrrmWn+ELIQvYCiRdIEvyTlL7uPypteJ+vWmfmTwtTYy/6hUR3ujFMG9SVB5J3LiEmP6WX
5JMwQWwDDBFc4I4EcnTD4FEYZ08yTkxuoYeG/u3OjUa7a4BhilJ0MnJ0rjRKvMdnjwvAtM/u+x1T
kEnfDKsZCzP/qfcg2GC2g2uEjGJl+bgf40Iu9a8DBXeLRqijjiRC588lLEQ0xG8GLycjWupF9pMT
88uE0GVZjQ11lyqcmYzaJ+iyWIklJIWpXumtP03fHwIl6q3XNSyQ8zJzj4I4Bsa9+3hJ4WUKWLQT
SEikDrHmMRv7WFsXaesleYx/ThyDMY5f1lEL1fCHEISSqUpRi/fRUaFY7xLInd8Wj2/rTs4I1Fpa
YLb+hoMgJ/gOzrwPv9FMKfc6/6ySmADGXBaCfJ/ZqNw7odWNR/Du5uRDuvURrxR7exdDyh/Z+rXh
TzswU/+CFuB3cOO9mtQJDEvgGM/41Wx6XiUsO6Vb6CzQ91k8krvz40GChxE8XEVwvumNoAB0I+6T
ByNbR5zvga6xzQy3fCNMUzg1qz8wv60BpTGUqGRexnPUSRQ8dEDfWzyujemTDU2YY0GlYHqjOgVQ
nS+bauIkMesRL3mkCwz4wAykGdEfW0fMFtKzi2VrxfujZUO2c2f5Wb0J8UJesAFI6xNplS2Magx/
OWKFDlod46QRKbqa3B43ylqAHPeLZ3y1FhQXBMyOT/b4BswUp1ijFsp6ikg5nPcJZPLtgD0HZQLr
F+jC11AlIdqb08iIZymGSNQb8SrpX43n8wU3lXXHQL43iNU7X3gxfiMH0YdZzohSDLDW5UR/eWdo
MZRdpabVcBx62srbCFax4ObqRKm7u/8lzjt3iSPSAT2at0sDsmr5wt+5KYKT+Ok2mB92TLmCRE8t
nSz7Dvxsjgx3AjtMu5D2ojTbBuRMWCk1wroiRK+DsUYpOW5W0BeWeBlFHdT8BZvB6hjCdmmAa0MC
CjI1VfdtO1I1eRcuW9iFFa7nJIiXHQYsR1B5UsaYRLmg+c5Rf+O50XxFR3KwHsIRDUKkpSKhW6Nn
IhPetNVlYSSprHcra/ccMdm/vEtge7W3vZECF2Ql5iMMGn0ZcqK7PfQAMht/t5J4CW3th6he8pUm
hkvcF9vwjhruHoLWESXLLZQnK2qBTh8KeeHkpKrWMmP5pk12vPCPGS+HZlIHqNWAt3oysiZsVN6Z
EZE0Ar00MRcGZOXeYC0sufqVRQ3BjO3SZkXxq4O5/g1nPOXV8HlLAzkUM1eq35tctuOmzvN2ECF4
qJp9r9BDOMdFWBLgle1H73jWElSbg37u+IKwRGioDFs3LlBFWj2vN6JJeDg2eNmqclweduQmpaU8
4yFtzbZaqKO6MU+4L0xjhOL+VWfXBfCFEOlBtV1ZZbVqDLRF/UciM9BRUJzu4dXr0eNGWPLx6Y/8
iQxFntkNdyUlJDtN4zMEOjGuVM69WXTb8xhlw9NR45fV6NZrAZCmcivGGIkAqXWaNigPt4XmZcZq
qmIBC9CdTw64naLF1OF6ohbG3/OC7sOmRNGML/r0xLhTrt8eBOw8DBx57u2N5dqZuMS42LnUSR+N
WZbrqzPSlvoJYLTPag1eqcuEVCrgMUGdBuJ2kUCmN+ds758phTbMNzGbK1orW3C+oXczE4fDLX8l
Z8AcoRRBBh/clTdc5C2Mmu2bGtq3/LUPf4nzJe8UCqfVkhthqtbosibE4apkhei1e/mx4/FyoYfx
YZYZUTVhRUxajylzve4djSLhhTWFuYHBvnkgtYvwM4SlK0120zfql1F8m2nNirAljyvSF7rlM+CL
Aw/HQymgGUcfdT9Qb6o2yeqWaau70K28l2ZjoAmSyXwTIIYHltX5Hg3OIpJcxldKWNac57u1raan
gOFQ2TXwD287qqX8qjLAXrfjHywi2UViieVI8zyrWtzlgwh28QGKmCI+UMdBRESDcoyOc0ni7buq
nPpGcxSlFIFQ5lIahqKcyc8Pcq/jGc6fSyVWQQRb5B8lq6pmi7mYyRt6cEECWzheEaY3nqcqdbvp
P8VTGCkcUdRGlyhKggQD97yrYLG7wDHXZQbvEvmaTeUQ8R2bj6XB6tDOxl/7RRH7qf7tWtYiyD2H
cohrjmbJMaialR6U8etf8tkXyD0+fA3RELzKwOUHERVNiw30BeUfxb+2HDAy1d/fAsJ5IbC/XpHi
TrGXFtmZpBIYWTGdfZeFwyuLHgeykuyLn9cXGL7Y7qIa7CR8orAV2ZPu/DK1RQGPV5JlFG3tU6An
OF1Of7qsQalIBE6D058/OYon4WWzjDQCKrl97OPJUgh6xcKjxBgEC7+F31hvOWrzC5xVVXtLQhIa
P88vkojeNllq++rSgZS1a/pdQq9IqX+RY1D8Eqfd0cb7WbaKal609Wu36AM3gJlHdYMQ4NY5+B9o
QONGHkQlLM+ElhtkSqAVRQxa+A2ffQhVx9ssR9VUCM9gjid5h2pjty/P7cU+HJ1U0WzFFiFnK/AR
LcSud4JAXzqaw0Dbzf2ZqRKL0QqSB4uM8IvYUHtRpbs1rzGZH9S7+RXshzS+MLvK7L1v0h2j74Xu
mlyQoMUQKck7begSrSar8bQ4+qP+Xdgrwzl6vmV2wBjy5PalyXZDfnN3zjv5rqiyXQZB9Ffia+cq
kE/fBbJFzRckz2H4qb7PaG4D0Wzn8fLP7m+d27wh8jlDKELWgvAsp/Da0jBIht61P4ONHmCVvqns
4xVojd25CrvAO/LoY9Mtu5KxG2L3wXXQNH/YBEhDJWuSA1Jr0RxV8NnHmiqiPNzftV6IugB7y3hE
KebbpJNqbDZ8VuiSbYoMPIW7aJ27Xb4wzgna5vdC2StsitL5KrNE3LW+/JGOX8G63ynu9/c4Iy2W
Yj1F/nFDJtnY/G66ewUUM1+hxc+/0kTWakMjUZjqgKOclD1dwZb1IgCFTBptmJ+GEs2NnKNAmg5L
ysngFvUOqhdHhxTYwDN7S1cTg4HVuIDTAJ4CxrUYJFj6ALY83J2i+bk7MpEZG8mGS0tXjtq4nJPC
VagMFjpS8alXomNyEpi0AQXpPbnT0bhuwBGYlpUlpcoV69arpn0Vcvz+ODRHpPfX715d4qbfRQ/+
UGRM8ikhXTNAsrmXX3h2XaWR/KVUA9vzn/4EhcrM//LP+9QKT+c+2LILjfnFC6vP/CtO1H5Lu2wc
7cNO8vDxJKKpzMVAkUdLPTN4hDIGfLbS32BLTlCFrNr91c2581mPrKCaVMtg55NXBYQqxI28mAjH
hrCygej2/EWf+/x0Zlh7eSGmgKkfW8YW3sBwkVQN5R/UfPwzvs9MFBFNul9Neotcv80dmK274C+d
MqUTTgb8gEmHYmcxe6sRE3d0Ardk3rNRyjoIc0zME5cKnCqvJXqWho+LfwHIWmyV5QkGsynCdSuW
xavTs02BOAHokCzagS+yE+YDk63Gcm18TsJMJI3KjSeQGbHnXKnJt74leygaFypJdAaEvIgHi9dj
pbka+b0SHaAIizKhSyr19zLx3KJYkbdu92fdmwSMG3neLFS+n8xta4DuRY6GCEjp6zzXsQcvKrBN
mfr8634T6lCY+JvAlnvCmvQV1mWvM34DiyhRwXlJpdzmwME5BQChou2E+Pc5HatspJHKQu/3EtxQ
Rp5I1A5GWlWXu8wBOL8Q3Kz2m2f1oFQDgLFd9r7Sp9VeY5ea1OcESuCtgveOV4e8yk8Rvh/al7VG
0QDnexm9Iwz+6gaEcXd3UqGAWBg1Zp0HAyJXBafEbIYJDn3NdoaWnEKp35DIHW/nW1curlnpeFAl
D8ymy/ML3MYWjqjczf0TOT9HEtioryg35pnb5LDq8n9lQQFtv/ObLerRjvzhvLDuGKKAEsbVOw5H
0AMUpAMeKl8a7NIcJ0UTa09xgFi7rk7bmpKUTbAVrl/djZwwkVq4AwqkSkOX91xgVkbE9G2+Uroq
IRrN/AlzVTNxtvkGdt7o6pCXDDdKP3zQhMaZR1ELMXf8MhG8QjBz1ZzF8VdUXgNTl1MxQBGeQBQh
iHOnrz+2m2HXGf4bHNLar1nTg05+8PSCns1zMldQzMdZVcanBvPWoKavDgNo7gsznL/KZ1svoKKj
jjbR3rxUc9MXLg5Qs4EGcL8R73NYM460XOsAebP61E/CnurYsTNOqERPS1Su0adf7tccCB8oFwHH
s5fgi6ABSGzw14tC961qroaTAq1nGeUNvDU5Mmdc0cHJm907mjpSgDGxL0wkR+wGWUWbU6s9ughX
lBNIc+ltDWllZWawe9hGESPn03HMfMqQCOoUweYfUS2SYyjDyCI+cj2QkAW73XLcIEEJ0SkvCP7Q
uHA56elPardzdMGKJ+xZVaffeFlQ9DiqLU28v2p4miWPqqeQzcfnOjGb3sJonW7oF/dz/2vYqAGe
BJTcqYam2CHcmG+zP1C79vhdZaxm+mFslylhxu3ZQ0FBUv7ac0MhAZOjAPwsY0M6Gi8eb4AY8KV6
4rBGIWsH1yKz1r/OPUrB6BzFI1K819cVLf0AnuA/WDgeUMShnOtAKUrz8A6m0Psu/ld+tOSPJ6xd
RrG/7uoL27V7h5Gvi8ZxuLnvtmHkAaJUF+ytOmhY8sKA/OPCwtnP3OO42pqdV5BFz7fsHRJYYH56
1nXD5DnU7biw3U+TTV9WPjnVnLEypdPgav407ZbH1POFzXUnVWSmxMd9qDB8iavIz1130DypmoDo
GwIFa38WmG4XmO7aaMOEmV7HorSpEjosHhFFr91OqxpoOc+LXVpuh0Dg5UYe+zurYC/o+8Y81oMc
i9yeLiXpp7f3dNKPZYpU2d1bNQZ/DvLbx9TBf+yYD8su80Hf/40vhNefIY09jKP7w9kEzTUo7MEX
wQRjxMLxIWxRbS63db+723speMZfgdUSS5bQ9BBuYOcTRZ4eVJR48MaXP89kk/G/hLcCqhYATW0J
8d82J1coev5MWFvjYdbF8mP11EzQAiuGwM6+hPWvewxF0VHsghcNZ8WPOnididJbCJQqFjaq4j44
Gkgp/DKkg9YlbtiXSLdyEqiTfXx4j6C9HACU2koM1e67pKhr7qRTETWyvoO/ccs3xdd5vym9024H
jwUEGVXDdC6sgIZ0WwHwS13m4VjH2Bx04rRlurDiV1NFmdG5rTNJEcGZ2InOTXBVTVaVb4q0not4
sqtrng1wHr9TPwzgf/Di8c06kPcjtRHhWdp8Hl6p7JDug1ogcvpuw4Z9XlmKhBZfPKbV4LWs4Tkb
yzvgMXYzqQNeWmSxGhIwXJGJHUNpazb1Wz4lBCL0c1de2WSOb1UnA2m8/cpcWeSgQoLyyEqCUbjT
PhHTVKSk2/gsmEVt/K1963fsoGptaPV2tcE7baklUty9aeam0rqLceE7gHv9sBJbwgx2huOmXdp1
zpTfRrcc5IflMfHlao9PzpZ+jrMSdE06BiA6l8mvccN6fUDuJsGny+yDWAvLLCocysY0OtUbrTaI
TJPt1I2G9x2KDrcMCeAf34MKNYmkK/Fz4nva22FA9WAwVjPFSLpSAPv/zmg6RhTxAAAjes+aZbpM
AJuv/PpKPHafnwWvML9pY0X/plj8hnXy6r/i4RSmt/VdPGdlYPtBM9hkukIbtTmx9+lPV5ZJsV8z
lTH7MpLY1Qo4XMm2j2E41sP3VyHXAGAeGDulwDPBxFib65M/2P4jPs2TkUIp3H8ZVMZxb10PLFf2
zWkxaEamAFnvtIdyqXD1xKm5ZzDthKXu9UeWGdfKFFPnPnZVqs3EMh50mr1ZaLamykahOUMhTFPi
XXrDkNTUukTOKIUGWBauZFOwmImia5xQbSycfsrhEtqdre8gNtJuWOtM6zbZAoaSXqrKphSmpmap
sBGVuUU8eFmPvNZeGyrM4VzMxarJreP74i0Eici+kyOvMOcZGnQIxb0BWx2i5p324zb9Bpugb1vh
l08Z2Vu8MFEv9F25mZWCoNCMIw2hkGHSH+pPnRS3PObtfojymQ7bCB4KYzwH08gIMl3C8aCGIC+p
wyZy0YZPowrLPFW3DTw3sYZukwZb1Q96jh+z2OQ2k1XoGbGqUqco7AxC9vif5fXMblHgP2whfDBi
FXYVVMbFtor0sQxgr62lX9TkVisI1tXKYLc8PkzbWTEUplOxd1FcCxeq80DitQcLMmLrUb3uOpRa
MPmk45MtQNHpPJ29OC5qP107TOljeRAgXdhM6UWtL619EhcUBxS0eIZsnQP3B0DkeSu9LJRV0QIS
+Fth/7mAIlW4HAi0j5zeX4Ww6OtVa37e4ZDQdwq079yc7k9CEaws5Uz6qhOlFVtYMAAOTBaDBnW4
yYZqRPE+o2eZp+q5ILDKfITJmmOONx6XQnFrziA4TdRFZNhwBjpWtT8zGjogl86yxGL5wrqssCXP
6u8vsxRE8tIMVAppRaL20Gd+9zoNHSJg8hAK30RowoWN0E+quqXEmGegdytcqIQdIykd+ZmCO8qI
E1RGkQuMFVZ8NoAssNFJjr+FPjpQx6NjWdKhYLLesDCzKGqmSmNTsIKlgt2u/39hSXJtVICdHTE9
kMwhPflOmbY/igULrYch8CJzzPILq0jGD0BsCMC38r8hyth66LKC86kmXJk+Qq4RoeJur+Iz1ViJ
GYPd+FfbM/7Pe+hgiB+Egp17c5lagkzgj4Hkh774os0TVNWKBx60wRhn1yz4CaiqbpHDzILx7ShH
kfczZKNaqdd5tnXKj2ZyQZFY9d0znZ8J4IZhT/5mfl3WqKGsCBnYokqAviWehRHdgg8m+F1aR86E
veKDNHAJNrDeAB0bJWo38fKLZCYgmgPXpLRYHNAE2gt2FTFDs+Id7+svXCjGiVTavO/X9DYRnm4v
6IjK64iXcLugv9KM7Qe7niUEFBQmFRqfP6APSUvunQqUaZMCwcQ61umrAlJzSTzw6pLmt3b9Olkb
5UUlLWQ8AlNSu/2qqckuJAVy6k1wrpjQGPEg4ZfjoazUq46YXRy9rILqW5Q03z494fwaIeeark/v
iaKrINFfc5rfpJmR7MtH5PmoB5jZj6kt3Dg09qfehT6VAObNRwhHho6u5MHSsOWQsMVO+2kRnjBi
VVSDU9WjIvE2q1Of90Bm7yoegZq/bJAubY3JN91YR56DtsbsF5+ebgf7HQyp2jtpoNjBuC+xYS8l
Z1R/NJufxWITaV8CejRg46wCfcEn1VoDtIGqRY0H8YJYPAa0gs441YDtwBXL2rfHDtH4IAvX6HKV
E2oihs4wraNR6IuMABJbMdxWv/CzIIMnuqijDqmykZoHYK13lngkD2b8uIxT950R3vUMsZaR53UB
e+rxESgY43isGdfpgwPZS3axqS7r8gkwa3VNJ98LktmyY2IelXUPDXnAGDC3TEjV0o42P83L0vI+
JN+pOTLblt+FsDn5wfnR3AbfEB+997VrX2E81sV3pDYkw+gK2ePUefJ3ZWb3+g5F7M+s3qw9/8cX
fQh0qYYF0CLpHnEDhnUlUvSS0lxZN+tPw0ygqEn94PDq/rJov/GzU3WKMz2ojNhs6SztYiYSHrvK
Eda87YviwVxM0KcAur4SjGDRtkJSn6m78Ta3u0RUVQKlt6yuxnt7PUNixvDa7pEA2PZmC/slFI6z
RrIBv4HB5j036sFJbhYUK8sFxG0P8sfPBe2xM4fXRtSABL65KMMNRsg8hKGDLTEMSM5C4fu1uIq0
tZUmgAKVVykLt35cP7UkvJmTCWBTgcgE6pUe0X90aA6n9tPjUENXJNizJPcXRAOyhlk2bZWidVcQ
qaUWtWWRmeHoDxE7LCSbG1N+e6x3/VUbn/sPk3kjv8XskwdYyhoNntzIW3E5qXFRtniSqqfW76iF
cTj5UOGq22fR8UVKujEm4dm+kq1wFMuLLHnjt5W1L44xBa0uiC0lkpqeWmGXi7SbDOFpX+dQB1Hj
uF7eP+pA1tlmon1owGZf4qHqLt8XpMaIHF4gY2Pzi3JbwVp8ET9/w1fI2FVAF+79Y1sawcVnMbdN
ZFSquwzP7sQD3xPRG6KH4A4efCG0xaB8LyuL5aeSC69gFVjZ5dPvxqn1Sg/jGDY560uuvUH9Zjzu
lX14NvywsLdByB3alSVMoFCQR0lK8ezcCs9XzkUiGv93xUw1u0G5ERqgYwZkbkoWtOK9KRZ4724F
nj5nvT9SQvjXJyNAgEuyqcBo/sz9UzVc8fuc7miTK4AWt55gyuMCGzFACCpdVMLCPB6gIBHuXYMg
RmkWoGccCtQ4q7bqsmJeThFHDztmRcknAgqvdT3rvenVjWcPjJ1gHZxP3sAFkbK9ii5EMOUqr4Vv
GdXou0mtXYhyvF0+a/VFDTenqbV314Xzoh1qQ9cP5wFT0ZyiCnhYAb9YgTfltMFbPTLTG0l8uKP8
L2s7qhrYk638jby0VAEV8pIU58ENCRclV5pxU81XL58vvkksIv5rbm31VX1QbgealwAOnrFpBCRp
mhnJ3zYZD+AUFq1+N/QBNggMFtGTm5lwQlkZJwjAXLSqhRtnBVeZ60Kr6Pm/BJrNX2Bj3VaRvn6K
8DIu2Ssy8D26C23WIPAGhVjxT60c5zZWQpAXfDeICEStsuztMTSPe1kh/DPsOa6Y32QfvFn0D5nL
EmVvkBJTs2Q6kUOzIT9Wd9Wlu1c8JBR/OF0xdWt7ffmnnBU/hb/Ed5mVoKxcq2poE8MP9wojxk32
vOZ3mZ08L7JKllIskl/OwTkZEE1ZGVyWe1h9/TQrECtqv36V5GH1wlMkkrAcvHXbLxgsjvGqxaPd
+adU+WNkBg650JXuA9nNghOthIMtRBrDm8+lXxrUuXSZVDI0O25svFDldB+AmhiTs5/RmB6HQSv4
pBTps6tZ8VWJlRobng8SvZWgzMWw0UHJrPaEFIU2F6zYnfF8j+C7EAas55REcw2mgpQUvSz4Q1lW
jKN41sbKlzm2Vvz7vgnDvTqA8icgUpJ4bmmvjTLsty2OGlroc+qvEwlKyby2/5qTQED9AuOpZIMU
ltrJgyarqEbRP5GwBOoYaRJhvLPFtI8bx2W1K53enuhLEMag5qZWIbzg4EB1ky0HZ7CTJAehuvZP
rXom4R+N3yWwKu5cKjnJ5ksbL08AlZHLQ0R/TeKwtVEh1W5f5zrE7dAOOQ4a9vaq25WO/0fnWKqk
a+NZ7+FVd+zgT9ZN+gcGcSs6UBxzH7/ucKs0Yi4F6O1krKKij5+TBfrkIyZL9aicwJz8YV95wAHa
e/YJQMPIUd3GZdeMR9f1M+gpVqWCIuNNPUu3fQ/srw/CGvB6WWQ+ta7YaROy7z19cdypvXhwL3CK
srzXSPea/BmTNgUQjKlp/1vDRyF6+ppVoDrOJt61h3YtRmfqF4cMiYdoiZt62du1BOIWQ/sk2N5H
he2D56XvDF/mRwr1mTsp6QxNeO+XDfeRRIr55Fl5pHx5jGWCWD/KHcnG2kIAvIExvKqDhxa7LjfZ
pI9q3z4Otzp+BEtHWbGy98WtR7xcBMdgE3THObX+EsPPsLca6rHjWmw8qH2mWHm4UziHAG1YKAdh
23jrsjcuCAzL9BngsggD6EqTshJ7nliyqeXYnSKDu5PfBKEfkGNuDvMswmm8ELWDrpPtwueyaqjC
AfRm4s3cVLu/23K9VSj1z8PXvfR1POHblWD1Ap4fvySnUvjr9m6YK+SFcIu5BzbynPj0922v+GTE
pCUdJSKhYNa3L7gS+pNpM74Z3o4ng8jg8Rgq96lp7Zx6vcI3YPJ8/6zQNHWPins0tJj1BQ2fFrdq
AQBe1YpreOZLCQUXOvZXcidPDWsf+TYtNzDbtv2M/Y1ENzR4/su2z+j9mi1ddQqcbiDOEjvAp+EO
iLNnwupY5+WQjimnLwHPqM8R6RtT9V3SMCR00UNzz/hescrCVmp7L41goG5+A5RuyDdB+3nV+p1y
gxTRBsgF7QockmH+CMtptz0wIAcIiGgWqSUp39zlGKwEzPpDDp0BTj6yE7Ym0WqU12O4tZkZTBMe
QV5DGyGzGfLKS0ZX8XFJb6e4iproACppCRaZUWQ9Z2ABCLX9JjPAi6VCOGnFMaIg6XrBRFzQmIaX
BAct9qN2pQd1AWj4CQgmOdXXnJlbgl1oWrWjFz9mH10TGYvdiiNvDbVRLzxQfFAiCOYRJJejb8pY
sHulRWYBeWZEf8KJNhi9E+F1qRhhk+7j7qTVCYiH0QkqhXU1Q966d44ju4ZzjKI59LZno6aH9kvw
IbDJb4wt8uaygi0IEgShlirmadSJ7UFBocfyY/3UuvBfhJtSKXHo9PK1tj8K3Tm9US3Zi0ZtZYAs
66Bsn49sFtNoFTWHsrELktBBJtOrGPycn/Aig5UoUMqmOmH5JrWjVcQsHImTs+Px0tpee/GP0A60
yHQQzXqnREq3Z90KTPNF+5qccUQCY/Fv3TtR0jBH0MOEHXDiPtRAkMSvfydjS5c1Q9TMndyFkutr
8Qt3BL0k3OVRIHAJ9BV6BHCEAvCnMXQqyEh+KVNShvELTjShp3vAbDDOg/KZ27eikiUGlsZoCzPb
myzcNcls88iMYZBzxYOnMG3lonQ+Y1XlIhmWwBTRQjfowG2yM5ec72TvLsj6c1JQb0K7b/Kdrdja
0epwNDpEeI5JKA23IFvaMXez7kC/5nqdKtH3yRildafo/waG3bdf+VwjGQc6xePL/xo/jo9A30i1
k3FFglc7qcm1okQpap3FwCzsY1tRbG88RzEaUQPOk1nDciUwRa7JlAS2YySN/+wjNt+kX4axWDXq
6RBIWZbPLl+ShlbE8S3NtqNg+aG/Npg5fnD0zf7tkcZvdLjeps3oq4Dj4sxFQDwZWQ0uSf+6hVtX
GqTtxi0WB4/yxbW1HbRQxSMCC0HmrwGvnG5Y06OLOYLnXCX69v21zyC04CeRzqKQDJphce5l9VN4
9mHLFY83ohLkeNugjOfRZoIsqXWsDu0Lgk3+GAAm22wgrW251phPgFEAeCSLP5xEpPBieZ6j2myK
AEfu/gZAI6EPDUWWng5SZCi4c5WA+tc99TO2u1KBVRHXAhbg0q4uP2EhpbiXNDbXgpTEW2nftNiu
pYqsMx/G3bfUg8U8vogG524K1Q1EGwHlO8rrHgxNhqTVNZsogS6+1emHbxZXAFj0moHIrwDqyCfW
h7CHzydUildRoTKJv08EmrXIeLjlszJnXEmO4fJAZMjg18/xRKSClnilseT3AOqkm+y+WeedX/FP
5NyOvIimDwRsZJ9b+Nv1fap3FiASW4C/i+MHRxarppkn2QGrnc5Qj0WAz33v4wopoZAJ/auQX0xp
lAjaSEDvFAs5NRKX5iXt4DXhmjDnr19mbV4Tu9z9Q1Exzy8/5HyynHSWspWwsA/V9BFbFW1ZAdgO
iP8ZB5BNmKOYMkXTS0BHTHs3LN8l4f3+qIYEP5wDLFiSTunMcZthwRAl80W1HoBDL6tvTvHhQtsK
OkhYWZbwr/nhheHxoQbpOhL99obbozrXJIw+/dbKQnzwEn6TbxlG7VN+1mbu/FBxEZw/cIqHJhBW
H3Wsmp8WiLSLXjhEhiIeMJTczVmCjpgR4U2pHbxoiGD+Z/yhktGyOf+kQrh1jo/K6NzxnwDEezOM
ehbQl4Yx0tRWACPSgBuiNBSjwp/LkJ93uq5pVg6MvvIgmQ5iaLhsck0O0/k+jgYJDDGxFruE4XH3
+tCK3ApuD5QxKqIYolslmduEa908CEgC3rQnuB9MS66Jwmhddz+6gmJ5lMK8OMe+AkOZ/OSy+4VH
3fPMQDgGye+OwYqqIQh2fop9dW4A+ub0o+dmVq6wJpZ+1mjwT8UnLeWXMEPIcqO9sNZCEWCMt66N
A6V3FBZV/RKsnwSJx43PvG7+p3KtSZP9M0knjCb9FTUrPY2Hp71XT05y7MAMoxr04BhtoX4oJ29H
CpIKq7d9vYhWzqt1lcOvVJwuuh1FI8CikKvoUJvrAj6bGLvY2HhX8p5k8K77TrHXY0DOYnHLMzSW
Fg0tFfcnRcYG0z4RfsolK6g9r1P9fPqMuohyB7hKrduFw9YJc1JX9IVo7aJwIE4x/Px5W/fSGYW0
Dg8j4RdOzmikk8AeD/ytEw2daisFpnJEA85Z63AZkRmt9LjqZi/GQeq6H/Zz8O4UorbiDLVmvl/W
hveTbR/C1/oUYiYws6ey3+4PU8gY+24x8nUIx71JEU7CAozz4oBrmb2suS3aOMEXxyZ6qiv2mejG
D1pCeH+aLCaJHKIsMGy4HeN9L/7fDd4JvnFQIY8pMNBGvxkI4Le7GDcxLQtfYXXSF/S+JVmXC0me
I8ZnA6Q56gBB1Q9ZYY2uhMTINi/FSeD81ScCAeTjWNiUfsLHv1Ga4iG6rQUSCSwuav7zv46CYqPk
WUnW2lIa8ahwXtaA5utznZhE/5vnardq8/PbUgYe/QKYbRETNtVkicl97mXbHvyXIDf3Khtw1V3K
Hn3DAbTm2JynopaYCcrKGbZyxaZ0W31TqVkK0GGVZLYozcbhPa+KDMBr/h6foVIKeXR19gQbL/nI
zl2AQoU+yL2lgtA/6Lt5BZP6NTA5dBW4Cih6QfjLnmSqjdCf2gMVNDfFT8dSLtlWvb9LP7hsAvbZ
7a+/rOkPj+vt1KnelZMVjCse2mCZcgP6x7KHf6Y563c+PSefj8P0RGaSGh7/M22G0dUUGO0mwMRl
adaFhltAMMnbQLq4mNT1aLgi/C+zcG8bsvc3fth1WaxXwLpY8ncH5GRTxzrpvQHAnXJhReWw+rK4
JCIPRaArawN5knoDHdLFUwY1MAw9No3lqWCBxv0DLp/mvX/zh1UIgPUjmwYTpWOtvvYCWXboB5FW
cK3Ib2kc4UaIuj2TfbB6QJVhHhsXkrsePUWPm2JggnSPhZu1p+dZqx2y8wqfkg/Q0FD6dwl+FZQr
cXJrstyJwOG0GM+gVR9snNGYcX9RvZDSXQ6ii838LDT/MBdRbL688bsvWj57HItIf/lmr5KL2WJw
I71AwE6asUzQ7nmu7y1x4jAH4VUK2N36XR1PO2y0o/pHVGmXfLQvjuZiOBGwZQDdR7V063gSvHzc
XQdoENnOjQvcqrA//4OSWmpaM3+b2MSYVErbgP5Ei5FurXwBWHrL4h3tYosDBRiOWhtB/ckRX+tK
9SIUtmz5BhMoPYmisFDind3jPqkghunnWWljctlQmvCTrrvcvzxFUNT8tLFrzfd9kBw2va/DFOfO
pWor7/NTyKKBfOrm7roSxZXtN+UBnWQwyjqgZp5YSTbmGGrXqUqckYZSDd+oKHgFgtAp+drhwIAi
g+VMw/FcA7lTRZuf3OtRd27qEbjJHwfCcZ77bEWMkpVcjtLH1hKw4vcNxYZSq/k15NQWhImFX8PG
/FN+hhZpGNvLoRnSMiw0PlpMJyPZxQQiUisDHKyZDgIQSEPaFQOuCW1/zmOzMMRct9bq4pmInG8n
mBVuh0W1GHz51CcvMjqHEz0IsAZApuM/02XXLAL7gG4TouOuU3cNnWMgX2dYL2Z1LITAIP/lY9wF
Va+R88tx/nnFgIuWibNQMw1fZDJJflQ7rTDaOno9kfG6HaQ2vB2ECifIdQFhvFtj7X+stXggitUp
KP1ivclf0dcjys55dAw52iXd9wFBJp5SYB5UCPrmf6w34JMLvrSvDewUbDCF1r+aiUVu4F/Wo0mw
8NXuu3gbtN2BuA3K0zQnzqo7u7w/Yd44iyQsEC3C7iIly2nQ0nLsFpgtRYM3C38uJY5WFho+QG0b
9ZA6MyTKPBNwl2lHFYV5k08wVSBx1Mpkew0p64y7mYL5VEJ3ih9SyMGpcBaGWEel9DCfMAbijEYI
wi7LvQARR8UKIpCZFpGMp510L+StQD1VsJZxMAeGT2nOaQxQMBGjJpi+rSV0E+KEAm6O8UUN68Nb
64vNRIHM7yc9wTb8kjIebd06le1Exya9L7Is5x2s59bzn+jaEhXP5E9OWuOu/nA0tCN21IIuOXsH
upF6WvSifrSzxJmHZdgesuQcmsyp2B1xShhvIkgnyeoSnlY7M8F7dbL1oF4rZ+c+RndKu9djwf/h
cUTe8SRUwnQ3YDiHrBvwXe2PXxEqPQ4xZn36HkO28912vGZPuLKzT2zGWLnl8GPXaSlw3kj3pBQj
0VUiiTpQnuIuVCmZOzUFtA3jFvYZCVg9HSnmQC2K++OdNM24fliRRP+r8EVbs8btSKV3q04mwFgu
gRQfPd1qWC1rT6PI4HX04Znia1LTKq3N9mc3uNyL799yDHoMF19orgAfyD8WXBIWu5ypva8tkfW1
05s715cADbxYpxx1a/3nFyBzCoIsYkPQ8I3mw5q7Cd71zgBdxaM0z/RoV1CyVMIHwo4xQQ7/F36g
arLSlPgxlPniy8XYpLG40nrc2kL4ugTwoz5MYlppGbNzlFnb5M8CgL3ySMVEkLUFeQRivEHwMvD0
2iBiR2J8RLV7EChcrGkVVOB6GxQvpwAFPseVmJ5XyQE1+KGrdd/cdNCgRBkVxznhzqXfd8VxmYBj
d9kOMWEWZyG19MCTCSBGYLadX58s56XDvy6vONZPiHjDr25pJg59jue7YiiR279rEHBWIdiUSs/e
YNoPx/jcfbspWX7dFO7ZLePVw85ZYk3cDC5bLVVPevg8X8KQbo0MkG2H1iA3GXm1ZNNWMeT/TPwC
DBAII83pfvnjwpLLO0tlLBlYMBngX9DR68oDUvoRgdjPtfKpEMtRPY8WBX1JRgIBh3FNlts+JlbZ
GAcSmUhRldj1OuA3hiy4g+mOYOveQrkYKnxuBvSGW0/LzHKIyo7bqDVsxGNfB3+UumD+rVloO5dr
J49TP6gmDb/1nHrxEZwgK4t4JVJrSBNJCBitsl6G64BaXek2WVgBQXK4SnOxiLcwVTMo6ya7wE2p
G5hhXFdyVF58U7Cvg2sv5C8e6m1PKZO8q1FqCPXBoeiU4bTtPLTr9riOW2O8fnsNBn4PNF7a/FT7
QrKESK2vMPpDvyNcUFwfBB34wEqvDaVhhUCxca7dylrew06g+kqfVmq16Lj2VIk/dGtTrgvFbv6V
brNMFg6wfhP8HWH+kCqJCivyQ5lhS5Q5yeb+I8M4Nz5Y357vB1pP9ziTVV9zS53wEjmeYpAO2+DD
oiajkdcsuhqvUNhzPgsk0lZYx6Afo/mLoTER3ifVhA2a1lKLX2w52SeeMRwqS85CwamqEozlZJB5
BmNEee4fO/NI8QZYN1GwNQmKKg05/F9KAaW84gbQw75dQK/3wdibXcneAwpn96FAEFvxMpUF8VPv
GGG2hCT2ypf2S6HRMlbjccVwBWY0ZnybWwBcFEiNINXjauz1cHPtKi4s++qZ8C4LfULk4XzZSvTM
BG4xnUvkG+6UsZNzGXCuvmFxTYcAsK6yPVHg2r0a0jKVRSEipHgmVEORcZibZP1Xsu1tEdLFrBof
06b5xP2I7mfIlhNWh0NsesfUHp9OGEw9UPbpOUEfJCDVTNJfUA/YL0KPMt0lfDnSdkuTGQPQOaKQ
VxTYUXxcyBk6aqipwDXRtDZKYRbwsPpRp3KEYwnjLi3PSZWqsTS5IY5OqlKK1cE8K27HjO2ZLdiZ
AMfYKsbdgBXDxKM8AOkpDjkZprkHhmY04adIYuqhMgQ2FlT32luUxJzlogL2It0bgRRD1lGH1Elc
CPQ8ES/b8QtlK7XyAyw8pOwquBxBiH76Po3RP1uL9wZUceOu9wsOXpZuElsU7+/oY6X1DB1gE8kK
78eLY+CHDgkpNexEmtoxeBUTKPw/C2HCsOlNXz5pqHiR3mv6MLxyEG+8Jj3WZQRUSDakqj42D42U
hzXs54bhcWZMuRD76xmSv4lSG4oM/FdcP7lIRJr9ek5hz+FEQT97596iXzSwuRqrWsnO18JpP95M
KO5Z6YkpvMaVhYo6vYzTuonsAdHDVZq1dBzXVVipkqIEGNdoFKLPp32PUN76bWrHvaBEQ0PS5eFo
0QBJXt1cjBa+39AXaiPxo7Wvnv/OcrJ8NSpW9tdEw0MqsGp3pRGyyAe8tpt3YKhw8DiUSye33moV
b2LeVYoxKsDtaMuEuPta7/hEmeuT6v9XmZk7D9/u5WCuJ9OIoI/cuFrLNjSnuqhvKiOYb3ecKQE9
DQf9306LSi9BaggqX//BxjT2PNEK7jXP6uzE/4qRh7ZDmFRPJEmkNtkPtZN7SB364AGRtUUA9ec7
VUY0eDBrNjrRkeODyo2ayAykQUeqMIN8d+QwQOWT3LXACbb8JRLumeIfHfCEb6OWdDg+lyezoAPp
lXRj02e+5//zrBrAv60j+PTwUHp07E7VRRgF3xewJ1C3JhFQi6gR50uYSXLcwT39k6jxKIfKN8EE
lI5Ek6VwdWgyjFjXTxQNwdLVbFZriIy3369/Bw7n3lfWlV4yRKYsm0eHQ7hZUO1hmxTfgB5cQ3Nt
/qPiBM45K8yWIc/mINa8hOEtQdgeIf16jw5PpkyGSXUtaDb166/0a/KG1k6znxiemMB0jL/IHjnV
Evaz9ZVB9723xNmov1cMwrEHJE2U/zPo7hcsvL8+EKT4sqHNB8YufhOimtioMKKjA93FkGs6SUM7
JdhKlNnXk09yTqTVLHwt7GBsvyFpTq5IzMKjyMeU4Zrw/JSmRxaevClB3oyak6zMTSTi5EAJDNPr
S+nTYP9PHXQMJ2kna6X1WaSBhxrGsZqwdrmi6wlp9gleXWKFvqQC4mnhqV57Pieg0343aArceIvg
ogsxNihAonjeseVnAMVAlaICOEZ0JoNYNYFFxbJHoc5Uq+lS6epbXuhA8LvZrENVhP7Wycn36ZiD
y86WieA8lFXyHXiCIFSzcqKhW/7mpd8bzUm6FvTYJaK+GJxriXC8FMuA5r3Xb/3+WfyusxwykpMD
p4peKwHjb5dpEIeF3y1HueXU7G+ClT8dcQEqR7VOuqxH77zqupOl7gI3b+T5A1Gkf12wQXk9Ck1j
JIGdnR1BN7Z1cuALU5U8gY46uzgYtiL4tC9HRr9Q09oYEfbGixwToKzebYo8g/0K9u/C1KkefvUs
AG0F5VExsnL0T1QW2NruIAS2EnnKRjDclfG8NgDtVVsfkgUvlTVtrgFtMSa5mWmCN7mtwDeODdf0
ng21yfFlfoa0cw6AANbksz1zjP3UO4DY1FFEujQEE6cjRRJaMVTMzfkX3PJjEGf8Ey7I3QpcFi5y
t6DkexuJ3gf02Jd++s+wxouCw/PAF3Y1ey0kw3yenKNfYVhBycsVgkUsHNfXu2y2GEwORwlKL7c/
dFHUMrl1S/dVseInP+ahlyMdbLnejJ/SzxEi/wP/TiEXODRxnKSaewy96/a+pNXQ+klvPxLn1TLK
lYJHPsEM/9Eh98e0Q3lQ3me7sFQUXXsYDIwPy883aleNyJXm6zJTyebNVMK45dFcgaRhUl5RwksU
8RuJSjlg8FCVAMEA8beOxulyRhTzju20Hxg/wr9FAuYPKBVeKUMO0SB9+9KMa92riiO4DIfhZvFk
N8PsCpbhnxmm5gfmn4AK7QqqeKX9xrpxkDkufo/4P2PXJ8RsFZz/4VpnWvo3ixpSedoaiVxwaINL
33MMx+1iCmQsnOTgf0vKJwmVKiQx+HAkq07Sdd71m04OOfUazJWDMV+A8aWKOzjQXOkIl9wqBFvz
EqhdZDd8wNL+EuVyZ9YkeXalsA+Et6q12PmgM6QneKvd1unedPGlhS2ljq6YM/UQEK6NmfqBVSfj
ZkkTlXmjMYBNdEEd0atA5A5pImRRU3hM4ew9ffMO2BPc7avDF5kN1xOMKiFFa7T24OWnEcFKKyYX
2c+Z7rQYICd4xgqfY+FD/jh+ULZ0sbriW7/qnjT3TGaBDwhz+1SZEcCVhNX8YswSHpDlU/uZc4im
pkj3nnj4zn5fx7x1v7gn407xBWxa7pdrlqUnMF4aYFfy02vKscy9++9btpez4LuNCOk/SRfAfybg
VBZj15C7Gag8B+yx8QmdZJrhVbEgX+N5f8G6fzP8dN3Fh/3tmkLKGHfbPws9bzGUHTsaYNNQA/Uj
LVE6Tdri1g7OfHu1AvdY5jGN/w7RkktwsJyJPNuxpctN2fvGD9TJtKFUAe8fBpQ9r/Kn3KaYmyOQ
zVtjx7RPFcUbQORtU0/2gL344A3DuB/diqcixWEy3mOO/e/f9fjQh7I35vil88sOFn6w31V3+i99
E47825frd5dnHGVUHUUGFxn/jJh+sUOCgmst6L9D7zru3cPjalHfhM55cBqxjFbMrhB8mbPSO0TM
N2jMj5Xa7BpT9haeaNB0hOoyoG7kSzexv9894SFgGO7T+Siv00SaCW0sgCVOh5Jb0Job3AI09Xpu
uOCnyeArQE5qqzXJfHoM/gNYtkTvF4wUSYv/kkPXYQexbHX74Jx5B3g4mUv6P9YVnjhU1XUj4UO9
MilVZtjHcOo6xNQejbRiezO3NwebJYj5e5uoYwcK2/d3P2ppeCjJRADpjpcsLHqMtVwUbwhmeOu4
LJCgBbg+IgJqKoq5ZpD2E68LhNnmmOidy+/5McKPaTdWie86v8iylRLuSphfsMZ1DaInj1QAnGYw
JfA8eH0emWStMkpEbKCRM9072azm8CfbqcMfG7G9I/J39/AqQmtLzYSbZK+h4ucS2qlia9Br0Efs
QS0FN3h1Q33uYIf+bvBsRjgfODQECJAN/a4eDjIO4CIyF7z6J0T87fK1mdfZILyhCMAxW1deTXqc
/LGADaQ1vn4DasExb7xLaneQqxocnqcpI0g5WD7BH9CrtQ8H/7JfBhpYWqLT65y/KYvlAugdgD33
tqzXQA0wjXskO+psSNkIJYr3cQl6oljYk2DcGnLSXqD8A0/vm3DttsPedxXPlOR/xNV888EBmZLh
oErZNQXNCiHkA2jevLJXbALUUp3VlODcYKLJorbKR2m/fhH7623k7rkOKmHK3WEZT9GHy1e0A5r3
97lNiI6r6eohf35CUSXkXfB2PSYvQvcsK3Yce+DGt2S6TSJTQ5PJVM6oxawEdNWnddjRA2EEPDZn
OwbR5chDtXIQmLITgL6wYbJekGYdmi9/g08q27WV7FGmO1gMttX7RIEUZ2OtGcXCXrMZ7HrMdfWs
0OUirIRzqez0x6DOnIGCVOBTqHAgJRLmCysyrbpda5N7ipOL98F5no73usgJxBc3mC7HQrWajrYS
nF/NGtXjXCFtsFIvteHdfIKn0Pi73Be5H1rXYdFAlTyClsU9xbCS1AYYQJid4F9RZClrbWb80o+G
JGMnrMxomltDT+nMQTIAeStkNJY55pzwUwuZ8b3S7nI0BRyYaIy1jf8IiBYCNay88dz+LlPVqDf4
wEo9UY1AZZ7X1L1uOsfQGYke0ww6xAfRMxkt11ql/IlpoJWP3HNgmr3i0W/oZgU3da/gwqfQWBCL
1+0qhdblPfsf22++EHb/YsLjPOioURwY2zlvonmSSn5/ObXOhmpFMLkqL+GfAAsLnDpY6hZ9lyRE
ejiaBgDYP+B8nfrdfEjQPBQO4QEJQyri5mgcflIWIDgA/qgV0kFgBAanLbaGA71qTJ7DCwWzyMZL
32fbHI5/7wA0lJxvdMwsiUupWaycYgFWaN8LUz4ZViE4TnLN09pJ0tB0efM3L2dgl7LNwtkmiRGJ
+rdGAzAzkKeWa8s+7Kt0hAepAo1bDihtDfo/2PgM4+l/BD37sRUNlZkGKfO2H09HWDz/FSVlr8tR
Z1wUPEPKNnv3pPJNvNuBSwy59DqHKpKxuQw27Q+hSE6r+/FWyfa/Ri/IWXpGtWznbl/Hx2Mvu8QA
kVAN0P5HLMFZpQeXgKtSk+oL/HkVIcGoDYf1ivtsb3UnDs6U8akcq+amkJLFuDn6C9qSrztJynx7
36u3wdx/BtrA+Y5MhCth1SC6hfvNV9tz/tJoWv9EOLHjfzcuMfrY4Ww3JBt/JTWcBuLJws2JfYAK
nsJP/V27V1aBWcEJBHfyIqKshI1Ua0FQ2LVwv78NNSCgBZ2DJB4F7GSLk0VmDr6SEM10HUiR9g2K
6UN+17B7b2BdCLj/10EtCSHHcsQtapFrQA9j1Mo6gewE46Pv3Ylo4wW1vzceOriSBXZtUsIhM+m1
6rcsYw3judaew0oORzZdXLiIiYTTkzaZFs8MYb5dYDuCcSmnxGYPvP8bRp+aphTcUkNV27Rw5z2/
DtKAm/Wyb4spOddN/nvDPGmUmiaJKpS5FZC8yn7ENZyOwZNTrfV1Cgpd2tUbW6+bFU+MW38LH5KJ
oJhEte06f+1yPS7GtmOyHwRWKLdEXXlx/56njAUriD+I3sCRZknEkgk8PhCtVAX+vU1gKnfbKOuS
Na2+83wdNKKVKfZeAYit/18VQipG++dL/S1OdcYsVA1SGEEeQI4FSC80bU035cv0P6XJiFi9oBNi
/azR15U8kjXnBW62dY8vXcUk7S+4OjBSAseId6OrRma5+o/jweqgjmgGqQESLgrc7Mzb/zSsQ1D/
Gtw8E5tOH3Fn0MFVwSo0SmH0YGiy9BhjCy2oI2gbqaQXEbq1ZY59g8SD217Xi1L3G5hSjO0/jKML
kOACd632oVgwud8DSF3d8V8ZE1gsxHXi02G8nEam15neJ+VXrSul8s/968/k+qxSFse9fRiJyHsS
FIBMy2CmC0Zs4eQY41jHpShIuJs+fkzMaZ8s8Ho/YfMELGNmJPq7kxxREEhoyd7+qgDzn39P/kHA
L3GeRo7/JJzR8GtlET4PrAqEy/w1CtPIcj4TxqLU85+VP2JcI5pJm3jRVtkYfGhB1JMf4a8MhK/Z
eB3giDlquO8E7Rm0KI7dUM0jRfAZQ/uLmrqyv+EWV+tcyKcNPXY7b/OeiqEbnmlVxaKy9cYUdyda
Y2jz9dvBFhQw+FQ3xJ4NzHYB8r/HH/bbD2d16eoNEIorvuT5LGmscSQJu/jYJviHMb9OlXvSSd9f
Lnid39vaSHny4quOPdPg9C9GYwKP2q4kipz1QUKdi/l9fvxW9ViKDZKI/Zzcw+rG3M8B2Hu963HE
NKgGjw0+gvC6u14swHSh8imgUKwJ7ffQKZLi8bE3PCJkJ0E81HwHNVNBib+3Rg3FAiQy9PP8oqTC
wSHNHIGR5TgfD7nE6m+BYyejokrvbjgdcYor6EF1v87Bc5DlYFxpjRsxOhgeYMm4oEbizCk7zD9a
6AKIciVsWL9rRUdpcUKi3IzUi44OJ5DBP/oyrVuibBZjkwTC5iPIJZgFGmyBWtOzotLdqt4m2gii
Wn/EUa8mZHqtDVh69wG2Rk8z8RM0drrIm68gvNPJhrOvK101Whs3PwfJyAU2a7MDF6sVVc+/0sX8
Uuj/TJft6x3k70sgVJjaZy1G+3k42FxW9RkgN01RKXGeezErDUx4JS0jkIjpE7XUG9SnBE3sn8oa
WCmb1c5mSK9Uk31MbZvMmMz9aYdzTP/w8UUgXLBYBtpdug+YHLv3Kez9jJIMJr22QDk4tV7Sw3Eq
+F9ryo9woGP4Frie4dUn4+9iRNVJWBkVdFt1HnF8uW1noJGLAVCfITJwmHDIyzX5qZYyWO8gU0+5
O2HH8+lqc8URv8AK8FJHgT3JLrCxNfobaYGFegIki84R5dhhLzR8UpWY5ekYV7rM8N7CkCrsV1GD
tEutPl54T3LLyXb0D2sxPEqS5o/PtJj804xcwCd8vefh54SmJc90G9BuIW9jT0Atz4zAdcgX/AAK
X74EYotRDL7pYJ/4y/0swWx+wSPTGSD8Q3NItwdMT+r/C9eI2BuswfaDcm7vOyPJ33mvRu6W2J9G
qxyw1bZY1U5QPPz0R9Yre89aGUfHVF9H65std5pEfXVz40S7sipb7fcn+jqHryyX6IDZcXhjY2BX
oSkpiQ0KahrEuqI1bXdNfgntQdsPbTbG3mqCz3+vCC2vZFt3zvsN3ofivvDr8AYGDddgch0NI72r
oCPTzEmogl035ZMvGGKZIqOLMZQWb+xEPeabl0b8GNgPmUjr1nDZsdARr/JlHMcr1c3mSx015sdD
zKKI12jpEeR5bzhbfrm6BTB8ThjK4P3utzO+ZEzhsAWVKfXV+DFvOjuSiQ2D39iChh9+SBfPLGoJ
nWmm5BS9yMvPdEu6m71eBe4usoRltyBeBidbT6P6qvZzVlj1JqgvqoOe2HxV/B+pBKIY37YkGhEX
G/hPCIVa1H8Wp2FQLArskKhteJkzVdm6/6JoDF8khsbMLu0jlDF1e0nLVwvISo9BrOd+u/tdJt1n
92sv7IaDgPSazD7NQCcylaIKw0apCKpiZgpCFg9/hWhw+9VG9nzeQw8gFB2LcqqoUbXKTe4WSWT0
dg5ZbWd0+BadGdUdJMNiKoY2Z9G1/zpI8ViCfYhzyTevxhKFvnvPgLuzwckarsZA2wSAGZeFn/s8
lnkDn4lVpQqFGgX7Zo60TM+saVRh+Dy8JxpL5qaSvEWhyj3nYj3KZFtnijlX8nqMPsoTYrF1ewZI
Nav4Eqe8aRb090BQhfoQMcQdzJDeImwKbBoeei9J1pqVD5uUA6AIadG4NvrnW6qrwY20fPbMRBbn
VTRJM14n4R/9i71T/0TozLDOrhwhWyIM7mnJtmSFJoNyPqJzjAx7+7chUmqc9zQXyD4uuAyJXAI2
nK2iYa9TTEdKaotRltruuHxWHtxh950+v8+5tRjOn1slI+rtu0Tm57wc5/7yT7b9SzrGFp1pAXLV
tbKOxGdrC56MroG2lFebnFmTf8plS7hGGFZUe7yxAMHJZ8zj7q113/sW4V+GZCK2LpS7H6kFq1gU
6cWTnbUlH+jmmSjI8aIAp+DpLiV69bE/tnRmjtHcQqZf/fwXo42ZZMX2ItQURjjlmPxGf7RaJrbW
uOtF2/GDutS2cC39LYuT4DcijnV/WQwP0dn4lJlNQa6p03F6tSnkYE6y2Vsx+GmELPwZU3cgsN1y
sk4WzXoFLwyhkKD6765u+Y8CLIHQ3QaGBiY0G3e2ffwwR12+N6eX2D14n1N616JcRcLIGOaaf++c
S1XJAkOYvSEtTyhbgUVveaEUdMRQFLB5U2dYRw/v+FTk2JbgBQf9BBN1fufm4TIiWRQl7VVvhjtM
nV1JJkEiwCSeZs6ExQfKkIYo67pTqLiWZhmdziRcWhLijoGSQcz8EMwGhOQCNE4yTxYzPcQGHFSU
x/fjXVknwq1ev7Vfkcnbwe0NNktMzbZBIBorhKzw47t+A3QX7x6GAgpSrq02Y6wRRMwbwMqkyZux
RV17MMsfGDv73SQWhPdDfNeoLJ9yBo49SyZxy7OrPlUnkOmoD7r6GFhTKTVobkoi6WqReq3OtxIQ
/lQ+FdTDZkkeZ+Fje4ER1usl6tD+ZsOvqTlZIyl3q4x5CkmHnLZ4YJJAqiOShfuo0IqeVEjQc66P
aGkaZZX+u5lPwBjicUBDcp5imgnvSHDmHO/boLEEKX46riQidTFf8s/W1FM7vBMj0O8H2jYRR5NA
QVjLGfxfRRX3a5Yg/qIGgFviX/NltfP6wt23NYNQbhCj3+hG1qIlSoCz56rbVW337a+kNFuWy2BB
CdIfK3dqrRl+KVfSOGXaq3QY4q1aPznTjf/negsyrKWFSl+iG+kVj/a4eY+lKEAKQrFUTYHh1ubd
qTIOkykxWBuju3k2hRzaLO/AkgY0oJDzlcnjMpch5vEkpnUSRA9aYWR19XGWvJEXKHENWFTMNjn+
syF6Knb6ryZ68+l6uZBrpuXCQrUuP/OE61KXkzOVaAMUZnHuO51klt3rrdM75ZcKxB5bw44XONG6
mCNWmPUaFOfy9fsUCWosBHJ1VjDhGx97/yBKD0X6nYyJwU3qv/OHcipwHJ+/Rbwc5Gnw5wVsCZ9x
AfvnhtHmCYwyaR1ANF0NQF3MrFgkG8EgXEfLhRLfRfhqv3HJewjRJRauEIcfdxp+uk+pBBHnKi84
AOqq5hOS+vZ7vqvzxRUz+BHn2MWQ/sSZjH+wR1a7grQHBbDEkrxLJWVFuOobSeaOMbjzgUm/+n9U
FxRLhjJI2OakQeN3tkQkVpVJYNUEkhdViI/wPyAaL1Rb8lsZn4wbyjPX6UmDYQMheasXh8vpDUWm
ac5YPiGTNoKHyqvO9hiHvPmMW0I4cE6piTbYrLl/EJoo2tpUMoa9hPEv3zGXqqO2Re33t9cltaNo
cuNHxCQd6yAnupdfZD96FQh+LdGZy0Kd3m/txksPSca0r4DSc4ihRsIWPmh4X9OaL69vC7eBN+PJ
yYWGDX4HDq/0wHTy+HfJ/Fp5lga2mHdVJrRVew1Ag38Hr/B0C5WSc1tBAWs0du8+2IMHqKBgVPrd
KPOzhQV0EDV2W0Nkjhy5VslxZjV27Ide1W69KcbEL3xvhqxq+TPUrwwgO1aowl9nnB3cvpTbBReW
f1UGr5mxKKlV+zv7BCBVmEW1KPQkBfYHV5Or7IEJpII0MEVrKWdlkG9TachtWWRhJ+2ndkfJAnm8
kO61B5uhPdU4eS0NphflImzcmUqeWG+7ABEyjBj3XmnSMmSo1H9aipdImjo1PF1DyFxeQaUVmyCU
wrAH/Xv80fX4KZbVbA4Il3p1qoZ3fOi2kgosGvbAMMJ9hVlYSsYFT5tdRIJZQn/xxPVXVr3dURQM
/mJ8YmkrOojBWOioFX+XF9keooICGUYOZp3OqV5BnzTrA4QPX4PXBJGvBIpEXf47uYnITvs5nlK9
k86PQiij9drli+jT3Kj36VrGNuLZKMXROBfXwF+2R+8UWqbQAGJeg1704WFkT6rnuJ0DyvnLZvHV
UhvmS7TLts7HWs5aAec7vhs+X+5320LWsMzZZKWHItvQcHUFJUwyM9SM52jbzp3rWAPgIs0isig7
oq1L7ovRaVwTI8jvRRVkU01k3ZJWTaFgK7j3C7MSL1lM4BA9SjB2rGSGOdZCrjMP3aBi8pNf9Xup
jg7CG7gWhMKDRewnAc/gPQFDQhXwTbkAkPZY7oKMnxx+BzQU4yh007SAj94wLpBX6NFrkmj/c2hw
g0g0YYR4K+/0oz59CscKSnicaWoqSskXi7/Vw6jno88oicVM3neLdsEgpWtlpP3YG862/zck1KJe
p28LH+k82WMMfAPHulR+IFuB1IuYobFI7GOSREC9+zw0HgMt1pVNZWQ5koAbCrfo9ikSkOpPRIx4
ePuKeN78g5SP4dxMyqcveFiXNqXBe1kB+0J6csnu8TEg0mFmIwNflyGof4mPT0uHlmG7LFf5wZZH
7j4qTAtpsB2VZm9ZxQcUHKTh8TJlYKMimyAdT4BwttaLkO0W0T55zxmSH3Jo0dymYKzhf3J6gloV
JKlI8TODm9St3ghwMAahhaQxi0VQSq1Y4SO6KqOG5DT8I9YI+nMZXKdvSwUZIj9s0XggSxTvZuV6
kbBOE+27UsKT3Sme2iUj5RSSnF45seuxuCZaXnpBxG02bNB+uEkuGlqTilwcX1hNDVZ7TXhKGwrC
Al5/ytSrPu6uhpzmVLfxvILGinnaJKFjfumAei5D7v19hY+dIv4UQQ+hECJKs5XV9aiQpVkcHkWQ
+72MV9lgVU3lklEvwoUU89YJYbd/hujnzNHHbqmOdpNS0dYqgYImQjxA2Emaqgrve8C+9cVlf1Rx
QmAjNMt0vvtMuehgaMKF0GksCpzNbuevS64hu0povOVO6lMKm1JItHf6qzVM/KKyAtxhCUbO6wbp
QX5WNNZekcKG5CVHg747HemDz9qXeqIKgHf4JdGSkoSmCTOJyEOJnY5OHUdJpGoyVdPqSaDk24h+
bwe+eZKhXJgtJjlIfK0pdp9hTPCZETyh3JMyI2O4/UWHDGzLif9uWDiyPZf1PdmiTwgf9tWeTZBo
xQ+kdlSMHjEx+kyAtI5XJxY9/VB/rAeCNC+dIqrdlp+Hr3dNhL9kELbQ4SQISt2J5UvVi/F6ecil
JEAol7vKTDIzAd7YKpopy/UqubwPDxtWUUIuY5PAXw2dkvfIpeAVrxT5fzrrIgo6dG9hrs9MkX1C
WAwcXUoY/78LIUXmQSmRzmw4eYmmklZaEWm/pwVR+CAM3g7VTehtte3riyG5G/tglcA3L6olNQxP
2C3v9f7iIfS9iFFzoXvIwtkxGqbVYYjJVY83sjMcRJnTz1UeEgROKgdb1p3j9jPPMHhkWgQf8cAt
hPrYDOd01oOTdkpxDilrJ+xahgNHo69Sb6JYxtufNltWHNp4iKuy1Dv6mR5QkQQ8aE6OChK70QaM
Q5lX0TpC+zKdnGIN2ZHpilsxRBXJaXvm5VIO4ShFEKl7SlsFNZ3focD6tgfV2PMQ92blHS3vBGxG
DPGUO42pm34eKpnNWCzzAo2g6LLLvR1PE4LDYSZm6I25waVg/VLmxitiCg0v8M7GON9/7mH6CDqi
M4xpzT+u9hZf9I2Q998gcnr4S/jjD46j0rMCta9HmTj4o26+438+fQjodAszNPK2pHm6e4jLgYZ9
WMeo0svBXipn9/DoVpmurpSsh+DDTX5Hvo1MrU1ttrWygp5YAnkkH+0PqbXDSUTVuezxKQoz2FvN
E4WTQnl7M3Cgbc92dTPGiFrSjcdx7jHR1rKDtb4D1BwHNpwNBadaa1VGQ9WjG/zX7GTAQq1bDjxF
Czw+ARNiv4eS7576AXWq7YUFrfG+R5NUmKHvWQBBcx1lch+qVnEz/9XHmH+ozXDhFEpPeNDXnSnL
gBlNSDNqEkEc0hISo8RRtmqAHZ5U8DEIINbZkAaLgqyVhDsGS7WSHqeuXmFNkDVxxi9AUrrLTFas
XRH2exm3leC4EAtTZXQehLIAXuQZtxXCKpp9wMn6fQ/c6lbadlpHd/wGCuyeO+/EOacxY4NPG+n2
vVPk1lFL4nFJSRtkWnZf/AnnR/Bo5/qriijO2PZQwwjXOZDUR66JnMiPfzcxVvLr6YVGzFRsfOoM
ELqkmHIawgJx7sNhSRuPwsdiAM3myKImSp02eQE7PUgVqzUcNW/f540q9CrP2VfSnlkRYNJ2vywA
vbaOaOIlxquc5zVYDiCt98IcifaqEZ0vVhWkddBvSKIaQTzCQadqawh8qK7JSqYZjjxv5bEGBXma
OHGzaGZiUhsVfz7LY8GRmov6W10zaKLW76p8OGgSe/3vsxNMK5+0Xein+JGPlDtC6gKNPrxVu9uK
niXJMX0s7dWGFRj7KoLZxrOteF29xlCvn8PUzKFJ+nMrSKyvRYbUH4riVUggzZfhNW9fzoAetIKT
cXhqe8HD+jT6OGpfTZn/61zs1XRhB46XjWl0xQCC2L1hdS4mTqQv8DvaZT4R/p0334yEeJK4ooYb
/p7q8k1rby8doVXlizuI+fcQEaiv3sxEgFh1iSjA28Fiv3Xw0weFLow/YJ9WYrClNPYBHGHUM0xP
dHLzh+R/1r7JbCRPr+MwlNnQdqyGOkHi9d9C8XBx2VtZg9rTeOONWzHpb+eLvUDLbNMGd8CkXaCR
bR8wz8BD7oSkbE7qbdlPmubhnf4phYZFS1fGjkRLN6O9Tz7r/QpVtntM72V4egtsJWd4a/wBgruH
AQDQNLg7lTHsmJ29n9jxCOOKGHudXQA2LIvuVfDxrgzAh6Mx3MtqUd8/NuF11ze99MDcFUqOX9Ga
Np3oqozEFSQZ8QWqkSf/A15qmjZ1ZBCTWNBHi3dMAEmxRCW5lfsW8I9pT0IPTT6DE254v2T5VHSy
0uZ3gK8Vo7Yex2s1jOJ7kCLrkArKBAFfkVKbbD3GHVns65rFQ+hiuCHtnaPWxoILroPoUZKg8n98
laDfSv1XaZdFTQEx969O+MHButbvBuf3zV3rx7W4YjrY4E4B9Ch8iVD76Kj2MDzOlqUUzE+vdWWP
TPEqOjw3OcE684XzjIuZn8U8kh39s0N4uug+5wetQWpXKcBpZUhotdRWDirPTAmKEkmOBY4cJwoE
h9YrcvbrZVSGQ/c0S/MHFJtWMDuQhkYkWE3xTrOsaX2G8TTBuRFhEk4qd/DlHble6qP2usVfbPvr
Jh+qHiQyLqFKE53QcfUEAc5gx/gCF2fANJVdNvoZlQuY46NSZgEuOoqnNXMmRrv/wPsPy4kx1NDu
uQQveuN3iLSbd2NFmBYRskhtI7LvJ2cDvS+mGuPvfhZ9HrV1U/SjwIIS6KmOshliE0S1F9tZp7yX
c8BzyblTuitkhHSgpYWfQpVAJjW8qe0icx0w/JWlebxQW5g8c52XRA3GgPDNzhy6zuJHAo3e2ypp
yoCuJAGfJqDD2gjzoK5Hl8RWaA1zuqIZ2bEw41lo7L1flprbv65JCiIpGMpgClQPMn2kRltMUi1S
2bLm19BWBAn9A/hfrWwCDpXt3nKQbOHs8xjcZ4RlFAqOAbRoDrN2l+IDc47JaJg5MPnuyDUXtSbS
bhkBlpf71SsbaxZX1QfBdfQyow10kcyH22yQczF1U2Ft7HmcoLXloik23mVFBJSjo2j59p7sIAry
WGuyP0hgqzRqx7akVKjyRJNfSiDyDg2YTM/oUv3cQMC2YDeueRbX7/bvJT4LP5Wy6LIvlNfFHii5
exrn1Kz96WLH+h6NThvJ78eW0NE8zKGqm5zpXqfxFFKE5CbAAFaaBP8TB2YSaCi2zIDT873JwQM3
qUIz0flRquhuDOYjWZGklWEIKzo1SkgthcGNKHDK2bBIZ7sedHtsjAJT1VR0BzwtWcoryhHCGOer
PlxYDPjMdJqBPErxMdUGtvCBTxoGb6pC/57xQcvOo7r5DS4yN7XsHpaP7gg8GyjQpNKmbJ9LP3aW
z+vX5iQZ3VPHRdg988PpqoyydiKf/Tl4iqN9xzHOwiRXJfy3aDruGl+cZOHX6M1ja7t5GqHeJ93C
w4uRkHaqFB0pjmzQJ9kWTCnZzBCgFGYyldw4ON7fRQEu0TjsN7cuuX/dYVjpothYjzPRXOwFcjBQ
eki9oqSwLvHyuxdpaoxXOAorRwUXflyoKhn3xMgaIYTAtJquySLBslOopU8eOZ5ZRuu5M3qkhZJ9
9XLWWwTTPTArDlWrcfH/7IgmG8x7qV4iUfh2S6mC/1pfTf/XscU2a17UDeg4y24CeiUzSXil7dfr
ssy6emPdztZ7h8IZAl33ExHb1aVjOi0LT2SqxwUjQuPKyHx/FQGpzleG+fRRgJoYzT7B9o35Bxbj
mHgvGNUGPRmBVYXOfie3db206sqLa4FsL3NOVMimX/i4S4X3emmUlzfdbXG2h/RdWDImP6pzMyDa
l5c4Xm34HMyXbOAcPilPtMyeY3xmoquUl4RHiP/ofJvgN1APRZpKqRbt7M5jeQXv5bfobOIh4qdH
zuQ8Q7MmvBdBivWIlim2Ml1mGhkNBx/iKktPJKy4NeszXlaTw42+Ywa1Gm23jBlb4U4CpXhAJ5Dx
G3yg9jwV+Elv2zMbZ0FobUGw2jjcXr159+cZ59P/eHMdPOVQmxfi8xdrFFA32kusDzqKPUrxFcQZ
v5GRzUCSDgTf8C8Wl2z/9MA0aQYf+YL6S+2ybXz/B4q82skBb6hLaaTpVLjFcZ3+7r9RthNDQ3Yq
5JJHwQonclikOATsfGi6tXZlg8P5UwEIxUMfLoJYEf3VCQB6pd3gZqgHe6sF5YVXYyrls/fo+rIp
EQKqq/Dc14p7VBVIo735m/+cbcdZ5wdAjwyHBPi0/ADpPSP9PzACi7ZZhe2qNH78Nb6LddVHRVoS
FO2XDtRPjXphFaI79bfDG2IOTTb1M44aSaAwypueAQUxCwCTL/SPS92ir6DWr5JZXz4kF1I7K/oN
CrEhSdhi4JpCgufiS+kPt2VRi15ZhGL+4P72EhVhLXLqqfmonN6Zr8UpzkWKf75lmZrYNO+ZrB4F
5luk3nfjLQ0w0nl/dWvdM+ZFmLaAxOYvO5ZYx93qyD3j+StQ6B+Jt6WGyWuRi3TU0ll5Hii3i1nh
rwNNSlLqRJOMnzbTOHSE9+YRYLWcpOb/j6Ca+53lTADXATbVD1KfYYn9cwCVn1jX24JhpLCcFgqd
M47HSt2kyp7YQwgVuPf1Vd/ypLyu6rw4OaJsaJ4VUY2/MsHVzkNA36k7Xm0fBdEy57QcnfcxfLXn
78y1hzqM2RtTQmSez0un0Cct+RLSgjWmslQ9V4pkb0Gz/bf9VAxsUj9Fn8bd0TLQhj1unyJol+ze
Z+C5UteInEIwE9vg3W+2mo6nknpjKPC/IZrws2ODOtiiVC6eKDvFi/U6c/pXbt1HGc8K0F+cHawn
XXu9yoWTou0tErVtIQYjSk78Te1OKjLncyOymH95OK5t8Vtq6yIv/3sHQ0bOimhczWfqKPnhySOZ
eJLEzXXUQAnB6YvE363xvvZvKAmU4EY5nPyNevvO7d/BI1n++SLUkYW/engZqDwySFW5pNlKge61
nPk6HbxnjVJiAYU9uRKAWytfJ8W/yIUronRGXu1Z+It7P/jMusTxyU+DzJ5XEwQzqX9yjFXhUf48
cnJZNzo35YRHfzkN2CY1FNdKVK1qcYqdKBXH/GZUyWXV93qQKejBJ8Fb6Pe+9F/Du84xCuWBJUm/
fQvr8/52YGFIWOI8QhsjWfB3+kiE3SBSn7j96WmH+ZEDXYkSHNiKIuytlVhzOHvySvGpvCOgy9xk
nEUMq/wdrDvgJO9gl44s8cssNAeovYKaxBS66FvpK0acVZSq8PHdBe0ZeHhpI1N4HuBVw9LvR+Z3
6WElfs9+ZpmSUlW6UM99jzBhdToK+ZVMzhdC7W6BIivV5mbjo0TrqnRBFnTRf8TheqLHWQFBjzb9
nFh4R1BD/tW25QMpou1hr834rq2joG09TIDTwDgrUorLKdNWD2e7ZaNgoX0TeYJ8TYmmjRuHV4zK
HeHKzS5qQ3Yr3jnwXdeK/1p2RKUM3CkyPTlU91JKYB5FNyzmFPXYrnXcy7V8C7uwiEB6wyHogfY5
MRLI7YZkHsOz1psA0JtghZcx2Uoa2v2lWB9oaNpP/JktpdukYN3Mj62pOLCnh4no8KZiA4okIk7L
BJWvJ7RHbRA9ihc5mWNj+rGFWNb8f9AIq/8VGaHOu4krWhIENd0lkGi4gPyCG27HNQLFKN3cy1E8
IIMoyYmsFkirBQLiIUIYmHk8dJimCukuP12e4wkxv0jh6ycYKRimmDuPOVVEzFxGIoD4Wyuw19w1
DzoCyJQHN3+UylGn+AgpUCNGb+//2z2gu09Q8gmSaxgzXkZrIAnu73D2azUuXgBWZ4AxNLPDzoPx
z4FGClEPtjZI87bawKSoxmdGpL89uGl++/P2pdKminwyEYy4xbBlM5o78VbVEcy/55mWGGwLpXCX
SbTmiPO/4M5cT+IPIZ3T7p4ASUw8LvJvSMiIsST5od0niOpYYVkwvjk3TCFCUcJQehZ6DymFx9Qe
TSGEl2BQiZFR1kbIKSJo0Kvbf/3bSlzNJwNT1P6asNba7c43bnwh7xxuPEg8dC4sWy2lLZFllkEZ
N8RZvl+ynqzm0XwVAvAIfHfwMxNs9rPCY0TZw6/kUbsiFc7NzKco1x0vgYSP1bbqoQqATwFMlixs
BPBhbwsnAXuLRpfbprYJI5rP+yOxKJonOPJNZCY984Mb4kGHGGQqrYao3Cho+rQuzr+0E/JN3LbN
iez0VK4q1B9iM+jLaO8kmPqBNU7f8jF78Uo+oH6tDFJEtdNmEfy+Tqjb82iOtIvIxM/yLQj7/vaG
XhRBAdexq/2wxyTsY1sjep2Tddp1gyeVZ4I0Weaj6Zi+J4aienehrFU2KpnteKGjrxRl/iCQaJjq
fymML+qL5rQ0Za1fatHd8m0tgBQBGzYBhTUIWcoW0aQBSk7hkteuWIppDffZx/FM1HqkfczkE/ba
G9KFMTBTUUaeJUBvEraELDu9WBp98ctghqWJ3GSp2a4rvSdfc4c0B3KJD0qMYvvH88sByf1y28tT
dSPiucJN2yXIORj1ogPhsYWtomJYuRy0IrlENR0+MUScswk5F5cbhaJV29I6N0qfM+7IGQ+zdbvQ
B/BL+e7FR2wM0BgjtDMdmQ4xzTGWIr1sRFo3jIqHiwE6cfFUCvBOiKPUxbt5mDBhdnADTf2y1dQ2
x0YIRGQ7tlf7vL3Sw7r0zgayPIZdOEGksE4qN9cOcjrmjLsv7ODF0cNvV2f/p6rDV7nxGVUBWnuw
1cNYpOMNZJqbtU+Z9vC5t9HNIBGdlV4v/eNyiK2I8KV2kPX2L9uuYEnpz1W6jHVU6R7n9NltoYcC
W8BGDYj2HI+FJJr9r+EItP4SJIQ3p5+VTHJk9LddDIkWSXJzvmoF+9Nl1VikAwso3r7sn9pBzXgG
no7HUuhJlrqteC1YOQmjpnCAXhuSLsjIw9L3kwy+BO8uw3UCjLmkfcdlJrWv90AKYxA4mRnrTxAI
xZnEJ5uTcYM5aXF8XTQ568rtvsVhHRbGFxIp7/JVJIAzdeiXhmdgxF/R7kD2GozAcTs6GJrtOs7s
fCtFVC4bnMXX6Y4O0nhEGpGENlQXAQyCxvGa8/iH7P7gvBNBTaX/ULJ2yEeM0mb7PkhMnAaCBpqQ
lYMQGkAtsxf7qSektQmhRdVMZvdFCNGizo21rjfzJmXFp2/4ZGt3IsEASk5IvI+u61NEjlET+EyY
XJP1wwPP/i6zGIRNuu60Ay8Nm1NPwNq+DrFAFUdedWcJVUr9I/+zMK1n3Z8ICdVAp3KQ6CWFBd/9
rvIX3uVi0U3nwCo1I8jiWu+a/OwZ/Jg+tVKMek8C9qqlRQVlZ7sd3IsGqWjChmj8GnFjt2HihAl/
KuOVxorHGTyChT9sa5zU3B7EJS3MtULQG42k7nO4lv0F8yoByerbrZQ+cxfpC9B31BZro8dWJjVq
o+wedn1xf7RJRp5bI+g24ccWUycdALejITYsNF/dsRwUzbRn3W2AZebHuYIEaqTOZT9dYredQygx
ndRK/eSp4MzlypVk+61MfPnHTaqSRsIQTGmKBJkO2YILUgx6awIfXEpJ4ywJKinvbg/g2TcVaCNn
s3laexGeWHVm3KbSC6Nzl5ZCfgMBsnhMPLOqJ0JvoEGyAwkVhPzw0V4E1T5zEr4wweEE8859qC6s
rvbtnTu/hUW6kdN8sVkCfMV4Sag4rYn2Jsg+/CTXBvCjSHpl0Hn9w+pbeacCWGJawm8SexLgRoui
JO2JtDaDsZJtMZ4g1bXbZR/Shihhqo/vVBow3We2aOVr7v32DW94pGrJ7SCGX2Hb9oIOUxOQrKlx
Fz+qaU6034nk5eE3AHqqJzWi0svDi4gwvhIuRrwtGtAb1MiD/wz2FlQeURp0uWPRZ3mlO+4KTK0Z
FZNLpKhEKPofrpmNYYmV/wDXIlxlZmDsJP4w3NBnyQfmdNUedr8EPzmSj/EBP+7i9y9vNwIQtSVv
cPjp/77dEAWEY3hfhTbOk8zzp52pHzZOE7Y98ETjsQX1QBn8PUuNwe+NiOV9CUy2lLr+Q9oMiCCF
01Jnvd7lVCBE0tGvhl2s07YszSgaDLqFFTLO6nzR/+hF4VJ2uWQYtGqwVlYSky0AzbkZjUVcY5/q
0NJYEJn0ru4ho2lAhX607oQY/q13IRE5wOvHs1OPA41MpjS5efV2pZ6XU3BxErtshIfOOAFK4/rQ
2Tv2jSvi0TOTw/vwwZvgEUHyNlv/pU0jEkrqThwBa7rKOmEUfNcV8XvX5KNTJk6GKMhTccH86sS4
hIPgXgZ8fKafBDY3tkTRGl7VYqYMLcMvKKRjAEiwtAipyUuTjzukOpJr1AuY/mmGBXh78QG7EjB6
Ip2jKMKR96PPGmZVaR5qfqdvJ1zAMaOsg3Yc1Yjj5R/i6ItmlPxJiBysOGvl7NsDilY/W6kQSU0v
xilruYGgF0SKy2qDh95gEoJEHgt0yImPHC3/iG3+9TCL+nwyYYGN54BPVoyPz7Q+aAgTAvqdyQV1
pqEklwjFyo8z0sjJnU8L141juBmyRAr6g9VYk+XNnX7L9ywXAuwzrnLVCu4kppkiuI/ztP9wyd5k
SHDDXYLscy2HxSvo3/omSQpZfl9c6SwvL53oSjYBPaOq1EmSRcM3TMuJY461kjEBCyRhLWgTE9z1
vZ2ichYnlM+53llFkWkh95+3qilOReftaZqR5PELiHgJHPfZzalbvi3kbXWRaCX+Z/SDHNmkCwR5
Fcqt9v4fWRGwBqWqZRMBmvJCTlSPdVIkh37eA+f53q+Tv8mz48LJH4Ke738erXDjkYHdltFaBdR2
Cjs8quLfNjsazArQcC+qlUma1XyVC49uZIqlwS88kwP8cPKpi8DKWEDhS6/vUjyss76sd3v/Vl48
J2YR2UR7S8d0axINjl8mOkqO+0+RjSHSm50frP8YB7yXwTHvobrcBunUQCLDDBJDFG5AEb7Gnb7V
bwz/7k7Yf5dS1UaWsmGlrqxcWWawS5FTFe1l/ykLkrKPpgSBjtYl+dwzMVif8U/Rj2Ymh+XZoGY/
LvYktMapc/VL04zORO4DhQTjBA1bYjm7VWh7EL5gbacQmMEC54n69hjIqTcY1Q+FS7Z5xffvP0JC
AAKs85VshqAWcbU1zoApdNf0dAJPzf/bbKKV8qhYSWN2R6FdsLpL3M3fiGpXfPSEhygFqBs4vHQ4
khvs0H8Si3Hh87eNGDiS2kAn69+KdZAY/jXXv+hAkrZIxiAM7pYveqwB7auyGz18IO8vcjhG42gs
7dNtKM0VfkUag23F0u2nTqRVfZSvtGzSUBw6FRaKhI0epoVbhYSL555t4oZxWRuMerUZV3zmwIEZ
1krXQwayCvxQYwKcINDhMRGXnd6yWhMUSmNI8EO6GNTlqZ78NMl7bb7tFuHp0RdGvm7Qrd7xv6QW
0atNsbiSpzapCe7vSw6ZT5AvR+T0WkY1rA3erW1J1wLpmwTDZeo29UExNPvbvDnCS5/RLrmLfcwD
eUYrkgGgtqF2w3PvfAnVaH9N/qhx7E2gKYZXFibsBKsDVBhhspuAyJFm0FUcYGhx2adUTHB7PIiN
xT7q8OjGmoh/jismY7AYiLCQ/W6nmwS1d95eY+rpuzQhRZoCqZrZxNHeB0wx9xNO0UuF8u0vS7qY
4qZUC1gVK0oL2sJpFgpacZ/gS6eN4cMZxQ+6C7zjAnhO0e7Eqk84YTwjYac8X1I0w5ueMKStUgCt
2KG1h/+LWwhcnnC8XM8krryssohmlloI87Il+5/vYtRvuS0AWNm2TLmJsSTSif7dg8ePjcGKoVpx
0XDyGjvk5GZIuvmCKDhGO+zQOupwY8uJZtoI8N1pbZPmVoVyIu6YN/h4VAoXgkZuYJpvjSQ/cKMQ
MtpE079+ElyoEychB2PpC+35lQuZTugNpwImanKo7ijrSTlScCkv1snmH60a5wMpqMw9sNVZP1Js
HWLifxfReRHhPboJAxlWe/oKr4kcgM1CY+Zu7LfV4xwN496/UZ9PGu7aQu3IZ0QkKa5cFsUDFbkJ
6pU6GLRJFJ8nuAiD+om0nfbGS6KZmufuMmqee1nTcNb96BeIKuDMGx/fhGct4J2LlGZjxlQvyOYp
/47LixmQGUSKj9C9MuEH69bhZ1NdnTy/LKcUnhGjHyJg6sQCs865MGsiBcEQ05YeWI4h98NDF41X
tlTVMYctn4fFzSVhWpzBZLpnM+19wE6cmlzgaA3jZgIyk6a0owbWkgn5ujFohXTFaXPFVlGepSaj
dzqmh4KGAwQSCvleGN5EGH/C215lX9f6lYZS0ja6QjVoOhtsAmL/ngHVSt8gd0+CcHD/WITdzAHD
EvMJEE1GI7kIDRgFJuSCPPoql4GJPtsbXMCfMnPTt3D+np7/N+WZK0KhpnUC+8eYjeVEFKFwZsKd
SoUzfGbw5LxaBLeGULU7GOKYIN0Y+9AU2zmwZY3qv5OEyK3BsI8GYqih/M1/kWos3ubRZx6DmX0q
5dR/ryG1oL8RjcKAXX/EbWpwf45FuxlcX3QdsZ16GF1rRxjaZpHH3Cq9US0qvGk3P8spBeGeaAae
DZoHi4JRGIcaaGAAUcWvfC8hAHueoR/wd+MWnPkQEuFxUQePJVhhJ+Wh6nFv1vO3xlvnypyIqenn
xUmkf5igY+TYbOdtVzyfdHUvBMg2lVP+lsD2a1wJoh8RjMfMW67Wb3nvS4JKYwrhegMCqMQKEfw2
Y6ytZyWctY9MgnmeUzRtm/KsCLZmwP61BxvIs7U0nDhUQYG9qdqTjyQJ4cksKSY2FWnKmrWV3lFw
L/zbdsCBH6zYyNp7TclgabGQQeCYoJvkvw3KH0w+tVzyJF0t7m7Owiqvp9FmN7IMHLcpEqy1M/02
+QoCf/bWG66dOZ012I7eGFv1gVp9XQJF6x67I0925uyQNkCemJ5NMJJQcT7+UofyhXXgzS8szyhZ
tJ2QCUG/4mCI658T01/aqZRh9Mj+pdJHVnnluFJTjQWCBZzloJ3Z58AwcxXXZjzJiJWx7OjwvGfH
gM/VBihsvWXKPnVL0Fjw6N0O8WZhzW8Qi9Cb6s6QeKNDnEr9mTjX5aftcPXSlEE9yEay2ZdKyBvo
dNf5MsgPNlRYHMMkij2HnzC8JHRRN0AIjlkP4xVLkpBcEop06GY6fdV0ndcdOaYHqM+JBUTh8zYS
SiNBGwtZuRodEXCeUx+UXMRYSxWCJB8jtsiaqAo8o7p7QLLvbFZV4v7pt0LF+0QqSppfYpu3OwHV
CTmESzB7xJGFBLpjdrXz+nwDUTmsOyoHlirvoCjOJc5z51QerOrcr/YB+pI28Io2L8KfQlYVwwgk
tHu1G7wq5rPLVUehWX90ImcI338Qts4rEwXUwia8/rMp0GTTX5ANWMEpTNAW3mSC6Zq1KSkE2gPq
UW+CaPxHlYnCHb03wGWjeNhyATBdcr1bvR47glPHg1wTIIntKnYEd/QSkuNuclNjgjfzNNuS9Zog
ypiICex8ZG4wDx2vwjuaHam79ltHH30B+o8lpAO625LymJOa68bgmxcRnaOt05JbtZO7Eaei7voT
78eO/vthE8qUdae8Q3Pi52acSMgnE+ocD2NsJd1S/hPUIlodERJBDVXRO/u3Knk4A01vltgYEuH5
k+CFWQd2jfwHOFmkR4R2XmiIfJTfizegCI/tcqIwxw4MlalbkD0i1tTdwExeV1r4T4zbNjxH6fdK
yEa07+NExP1W2ADjdYh7U9cALfxgv8+YuQw7+Kykqjn+cBFcDf53TZs3+rso8Mn0+mXDj19lyL2F
61pGhYEawkV1QbNaE6rxAhFh/APXFGpGy5t7xl9jiPZzxw8I/c8+IWIPfb79y78nMDFqVTVoVgb/
Tb3rDnaxJilIgSsaiYiu6FBTdo8avwaxHd/2+B250WIAPXSY1MswBxYBIEr6bDddUuYF6PzT0/7t
IIhWEj9ElpVAQhuyUraWeqXn20Z46wHQpN/UZyMGbBw5ZiHgKvdwznyD1/7h+dB4JwVhSek2tdyA
ZDZFz/ym/Bq8AY0a4YAg3wvZwSMhNHTEv6Nf+nBdT0A6k3IUJ+6SUo/IgAeRLVG/etfh4ftzIzOj
vEA8vWedmUooS3s6h0VFvY9mn2H1KZgJWwK5T3NMuG2HgdVkQa5otfIrSBN44LC1BUun779UpZo7
Qpl1SotzgWP3YC28p7tDvEd369HBiIcGhskRPm4/wT89yLAoNsD98GueYsc8Rdq8Ayj3xCCd+Vax
XOxE6d92lELc1QBCYN7qyZRoSD7q6yJQGY3e+gmSk5xXASnQVTKp++N5n7YT1ecLZBfUAVAs+vVH
6BdTedW+dSbRcE1Ov+jSO8ODcP/NbYCsQjzokWHshEhzB7hU/uGvBD0Wx5DjFnwIG0xBalv6suOS
V7DmmLBW74aSMM4wqUdB4kEwktL21djTcNMdsHoPizO+NdiLbW9uZpCqv0z79Ywmr0u9X+AqhllI
W1Pq8zw+fkg4vE6khdlOu2dGEp52o8qJc4/bgSJBM9s+Hp5ejtVT1QyMiYe4F3MZuwugh2tCSvR4
szh6sRRHD4qyjThvxb6YdMKv6pM3ebUonxz+tzcCPOGb0KyYDCwYAGdmehqci54QSxpWXT3D0TUn
lnO+Hwxe/B6TMdt1UbvqsUzkzoXHMHHPaNguAOltr01N+Ubb/aEe+8Jv+7/pu2FuAuBqF7NInpMH
qlkcYTh/wPkZ3HXH5AYXwi/pWtUNAwKyakCfRkMjc9xZHUCYDqh4g9M7RtcPC+Cn4dvc4x1hlV5w
jVxqZQenMBNqz62/n2MMVrlJWXbmwWyyxLR7BRirHU+DAZNe6T3m9W7S1BelTw9OMXlP1Gx2SBkv
iNN89IFO9UOq/26552CdK4LPwl8gfhaXxOBXfBDrhK5zxsoNiS2KGgea02DPVfBSo5G7JXRWA6YQ
HaJ5+dG0Fjldh2sWENA+sXr00Ern18H+HIEMK831uLwdLTUSZ4NTrrbTsx/kNV7NpLhrO38pbEjr
bSz2FpxYOueCEt5xZWD6Q4jsS34hVWL6E/4w0KUXdEp8+j18O3m8q744yusNkJiRJdx69B2L9heC
YJPhEMHuGKEtUmVrobDEYTwjeSWngLpPACXzStKuH4z2Jc+PVYsMoOBHpxzgruVzKIkRMSbVju3W
dnqgBVHtQukT1bRjNpEi6FxNCAVvAOMUYDszQ27+iZBwinLEweLl3LwFv2fEgL09YVfff2Nr3VG1
NX6BDftWNw0RFVK7s4S2iHTN4Q2b0fmCFITUWw4zS514GHuZqKZeLLP8UP+rnbcLxIiADm6RjZBW
tD+GZ2iqu3ZFmt1f4h7DodlQxIA4HMOgbyjPavJvDfMYAemjemJyb1rshtiDA1VhSl/vR/gj4HpG
UMZwWNaw32DmM59gay6DbY1LvnhVy/rqi0l3Dqe0QHsVx/OuRlEzo2BWVHVqhXcPYGU9TCG14c6u
eX6e6MeJi1rgNUBVbsVa1yQujZUyY+GzQcFL3ZhNhkaAt7sR2OBpYgqT25XAjbTCEEy10cLCITNo
b7XHPuXPFZe+doFJ9wR02MANGtB9aVCuy0djWNH/GSRpHcxK1xBs25l92MDOga0mGAxl6nTtLC/3
sWgSpJHw4clyfPcCcaDmmgyVI1HJqTTdgr4gXf5e3dLzKSDjCCTkhzHvVZ76I7icwGyfZJvSOawN
n7EUsfckJDmY/rnwUtuCSiFW89FDdT5q66MrXzio1TL3AYGiuC8zYg1WnCMPi/ecQTQjkyGZ3EU/
rAeSd2qEmc1yHzyxvzOVTvYNHX54t65dD0TrAx/7Ve1Ri2IbMCQmfQ654WYWK7P4kpdLHU/9uvy2
OuYGHYaQ4CIYhFzOM6M1HDwfa7L8f8jQZUf5z3BC7UoV+YWtDJwK41SP/2BskEfSOqvZEv8GKrvT
nAFFPYcojk6xEmKFc+9pS8m4bv10Dp4kxeptY7geB50xPfVPV/0ydSR3Gy7JTYdUtarcjU49F+p1
XLRTJYQXxagdAyW3uyBYnNbvS8TZwCFu8oMFCXTKfiJ0ULTSEd2RY8l6wiqvJfTtSC7qv4wwYu7t
QYUdfG7nZ431kod+mMml9THQnfBQ4aiPb/psjx/bpIM8WDP41wnzLzCkq+c5Q2oMonobgJFH+j4V
2XW5dkE/q/ZDy2MRFN1qR59UwKnun+WB8Q5ZjETImpfPcuN04w7Ec4KkwY+//jwsAO/SiOVRLxlE
X1WXje0Hlh7oGg6qKIviLBR9sZU6g1PNgfTqNxXL+aAjSr3osJU5DnnF+UEnB5Q27wV6JqjcLYJ2
ACXwlj9YvnhoCkA+Evq0u/YRMpvhbm5A3/MV8aPKhXgZIkGOIM3TE/lkvWKLU7iI5le6PuR4Tgey
zkJaS9K4dw+RR8V2c/Mg8AaiFq/npC9EZnxhDj+uJfKQHI/qwH5RSJNTESm8RHSDQeoiVL5O9pj5
6F34cbDhcO+xVCfbIf9bTmH9dSyg7smN6EWz18busKOuCy4Sqf5TfeHoc3GEZpZepaDVK2VRklI6
S8VYhaMQ9T0G36eYvBvOgMkJcKVgcEUHwohDZv/lxwv/Sm314maVab7JyrnIVhIKgUtkTofD5TCi
y7X0e68LIxswUtDX8tLz1AJeQHAXyoAhyoohckZsTa+qipPnnN0ATxgQxQUYOcd8Pd8ZLTzTXSVw
Vp3OVKsO49EgxibsgBR8RJeCzCykhBHvnhinJp4pvxn07nRhM+NCWNk3GBP5U1xgUI9ESPbppfTq
jmHy2v2enJ4sLso5o+EzVtZBKR/9qLKzZuIpD+FXI2bSPPHFESyeXyp4uMlmxTMl0EpDBP82vtgg
UL/J1MuWSmR3M4ulWkK5EbFENJ982+JXMNCJCdOcmJ9ZkLEUFRI3Xd78tefWK+zhmEH+AF2XiBTL
C7NpWR8YWAdIpp84oT//PelwKoeKuCj0QSDwmNoktqTL/BuuAgqZ7YYIQe56Np/uD2p89QPfQYpg
xHQ6negGkHJYBYZOrX+QlYA0fYqTCZVtMKKmH3k1w+1a/dL1gTzMEAwHZXVF8XUAtURlOPLgyTOu
Uh5I4tx9lioSNDD9KasQCV3S66jLqcKORUawv2NoDFw4rCXxQx5I+cgmDJ6hDEVFGqpgLDPmHmmc
iqud+do+0MYfl2HIqMH5w1Zdq7NMshThfxFpzd+n8iCvIAKRw7hMtRyL7LHYj4wpfZh9A5wunN3V
xtZ5LWvUc0zkw4CXkqPH6Zbzixcv032yOI9lSIwyOimv5sKjjiYnUqqDWZJ6aVmUz8i5OUN0aLPu
LeBZuHZNo5F5aXGUkVx6vuSFv/8ItN6wsv0Giqocg2/k3xlLM32hPclNSb08zTMyZSIh/rvjUCjs
OJC2uaEI50UM4/WnE9pRujKxxu5zBLG2KD6dkOSt3/letYfj2tc4VrrBnVp2lH5nY9Eaif9ZHH1k
Lj0IIsiFXyJjmFkm5onw11IISecIWL7Y07Lc9UszRKS6c+PSatzvkLPPJgbbSDroAB59yKEPxNkT
6F/ib/DXIEGVPi4Vt3BPicPCv3u8Nn96IdkmbF3QTWV8ZyHjzVpOHnWOL8cIZUSD2nkFCizw++Xm
IbRjOd5k4Xcz1fm/nIKtf4PGx49B14dMIk9U0GL7/pJyQ+gayM7S6rE2ZZb0Iy14Ky/+apT82sRP
wLcCC0hPDALKrenISIYthGccE9V+Kdc7y9jbFBcNEyVY+b0dqJcpLnuoyJpk2w9jMdwF2UBAiDgv
h9r1q1XyU0fN0RSXHzFgbujXTmN4Vfxcu8n5Ifx0QH2JkWDorBWNx2BkBefqxkONbOPB7xCirQNB
ybQyjKHDZUS6BJnamYhUKcdni+OMV2U/HeB9X1VklIGGFF5IDtwddrfN7DbIyjjznNuXfruSQN2M
dVvNqwakBRUqa6Mfle0hTOPnLPkZ0szo70nSHYTW3TutnbXwGFVQs7MNNGBqXmL03big4yy3O6QF
Ny5Z1rxYo2Ni+gbwIBMyDY36+3Wo9OEUMQYwIquShgRX4iS50QEsQV3fSjB/wnjGa+77ab1dPSgE
Q6+TuFYxuQ6bh9buFp9VIDvZXdJqCPTRoNIk+K4KKigcmBjj0/KNnIWpu9mtGIf9ynqr1Leq5N11
gAZqvk/vtgnhuLvkab2Ir8u3EehG5c6U3CqwvwMzFY30Upab0vIly36munGa5ydLLkBRlGk9PbP2
Os/XNHc6cKRQPZkNVrfGm28deL4lh7bnbu4J57XC4PWZB5ZtTvltzfpiOE0yJIITihbxKWeR6VOa
HQbqh2OymXsSGc4rOrfOsugaiph8Vk81ykQ439AmvBVEgpEI/rMQxuhM+0NOnIT64pTWefSV5z3F
+nz3t+1LYp+/t5XYB+zADipXsh3fbsrzJaPcSgH/Jk4GMNqMGgKJhrUEwPdXoWxUQVKg+CJygOM3
u8IwAQkOQW89pruob/GK6QZHu57MXTkxPwwOvVV9gQUyb+p3M/ebxbFCDil3uDj3ghqWGnxOfnVY
SJbuM01Iv3WuOLMZJyqQ6Yeolz6V0zpEYRWcxWETqrlSjndAAFdZRJsrO1fPjfwaC7zvon6m4LeH
JgdyyYccmBCGvNpTXoysfIfrWkA2o3i7l+KXSQfeF8/bb0W8yrSy5/XcLIx/EVc8TLyK5VTJ0c0O
9Zp+04GfSAIHYus4RhwrblpFLIzqMXVCIdsXndDHyUrbs4bkBvBMeUWx3ogM/lwhTT7//bMkZ8WZ
lNyX3dtcIoI17F/cr5Uh4QkEU3VUvCZV0lhWfQd3aburc4bn/ALC3ZB5SXfr0DcTDQckVc914ERc
WZjyrXR8Fx0C+mpCCOARBXcYtnrF3V/A0HM/HxaCH2oCGHwqQUoTrBFGVn/cUiQVgEgLzHf5HJ6l
2vDMqomdgfxV8Vj+fgaQaSqiQ815F5pxMSE+YU3doHRMO0kmMFJoBCQdFsMdY3Qd2wrvYLpZIXgX
Nd4JzZConSOIWaSuOWi/gmmJ6blo0GZ0wjPOWDBEHu1HPm9f2zr/snXoiUDQrspjtvt0Po31WIEI
xhhwBA4P8Y3D3jkIc7ze113YKzw5uqBUzB4TspIutBOFV7gSScPtNgIyfLaU8Iyc6ykYv+1kEH2v
oLW3u60ggS23yRCpKgY2GhuHtA+pj8LLyIxUUYbOS/ZAA69c6PTT6zlRrxC0tMsHvkP+R82C7Smx
mnKEJrffLsp7ri0taUz+IODO/gc+D37pERn3V27j6Jh0SFY8oFUKnD+4OT+zVMrLLVJKXbVl02+7
h/jN9wTnqWMRx9520AVg1N+v90twfcm0Seyvw9hGQj7Cn15IZfq2+E1AhTTYWz7OGhzxOzNmYB5L
53VfEOHGsLowcFTHu2njdK/6auSkA0HD2gT1SkvHy0B6rFyDmWSRV9fegSLK2cTM4hokyEPchW0q
CswwKFBv/HingLAEPjTUMsyEQNOA+RzJqUrpU/aCQfvX2BTu5xx0hDaZx259lVIoUklpbaC+GFZY
p4JcN81t1kR0N02A5ZyEo0NM3mLs+07cewx+F9fgWbbOgCSjO9ACVErAm8sX6xDDjzWADBc2P4mH
LD/ViUvUdaOnCZSaijaZuvwHT1CzApgbgZ6oyk/JgI5okcQiYAbk1jXCYBdzLRmv45UL1TkCT6A4
lNIxddVEzVh3G7dZpq2+reo4LI9UAx5qtCWKPrfYHUArhk9BxGapUUmsUkCZh7nhc5f3T3TfuX1Z
drddxjwRwW+Tz6Cp5jqjDcSOuv7vuULNRrhMfAd4RvyP48vJMANKp8UX3vuodZvrsHY8ak00pwNc
rCPmyf8SfkMc5+fPHhFMHgIkw9HazWkrjbP7Hrw/d3ytkfldzFWU8e6j3sBM4QbSY/8N+MVglaNK
XemviWgEFY8THvAxrOi34Mg8RIUGxOvnjInkjC46FV6ioVM/2Kv82BeFgiJxUpEMafbJfqOpA6Sv
b7TR9hX9shH0kFmMOxVJ43LJ+OzMt2JhRbfN7ISFIoQxqzZPsCRTR/toOKjnHP1yXywgp7gekTR+
BNHs49X1KgwLSd2v17uA33W3TulPY/Hsl0O05FocPZlayH2lQYcOLufJqCmW+Hjxk+LwvX2cbP59
h1PwSQhmKG55WqZZHDANaaWPFXU2vo68sEkifVbyBRskyOMvXiU17D0zX41FYNBECTE54xhSC5yO
95pIfHQEImcRGt1IPBxa0dp8CwIh1oRFk3U+uul2Z7NjwvaAeap33uM9E4WR5ksKklnz4ziHhVMs
7osLwfoYdDPsIgTaa/CLK2ZdrpzLS0AGdBkmgpHedJqmz4refbGB3Ml1jBMu4LsNhYLYThJDSUJw
Zc6xAZlaQOKy+wWebnRNQy3PCJKDkFazJEJrBXHKy1zIyVNG4Bd0IM6cT+iKOeNfQOzMllq1iMvl
3SPzcyAnjUCfBtDAxgU6VTdv5z3timgJOfqkWrg+etByPRVU5yIJsZ2O46r2LhVeuvpraC9fUFg5
WAIAug0GFG73VtCXsbfX25seS3kAXkyH8qSY3d9Jah0faNnU790pSlAvymvW1bE9KlH8e6Ai1aRn
wEj1tNAj4EvzKX68cmeH1X+XDy+pAvu8Inrs0qFu2qP/CLY6fuXu1f+YRkQZXCFZ1a5Tj1WQbymI
4NnYvawLgt3tAZHWuFc8EuwXQONJLjnAv8JkrupHyMxdXaxlnkHuAWsDY9t5W05n4dVltkibEfcD
ySEvGbNNr5AI0iioIrwnXcNAQv4mFBMlE8i358F3fKSpxcMJxBVegRG+WPkWDM5pMXKH2XPhnRZF
hCkW6v+Yorf5LwSSjG0J20PTQIK1/iN50Ss56ICaYepDZiWcxkyRX8shpHmOv5c3WIHRdKFz+7dz
pl+Asg6Xs/SjKSVyHZQxF80SnedIY1dZjMZYJU74hEzjqq6fMtrEhGbjyf7JkGW9/HHUTTVk9L6y
aDy56w7nuLUi6F3Hb8RrpINZ1SND/Y5eB+z8JegfMJMN/5f1qak7IfDkEkw7FWB+DKXG3usjayt6
4ICmF/ppNvk1e0xxjDwPARKxob0V3wi6G8oBmcAf18VBCoPk7Pj7cR9mlH+L2yIZyUHcyIbxFcvg
PSKtkpxTFNwtuqcEhHiFZ07uvl6xc5tndTT8HYIDG+EQ58ZarXOf1n5r2ATdk+BAzfTKWdSf/A4n
MfEnmgf2M59tLWQHT6HkNrdKnetpvk8KIANG6dKi2YH3ggc2DbWiR2LC1zhyG/w8RiOfaO4tHapB
sCzRgyIDRRi1StQmGdr6RgiLlf7BTf2NFRdqPvldm3oBjvjkIpeX0hA2PsNBetPptjCEqoFrlYZ0
12+i31Vy4gG06aKJvxtgrYSTy7nvhpAzj2XOoeJY6AOHZb50D+meeo6maMu6BhK8+wBIYHKC3SGf
peUSk+LMlyJr+ARsL0fisRg57qj4x+AfKFpmI+MfdAdXcd2LvrNA6rToWquQmi07Qfbj4B+lhpF0
Hj6ljPUS1S0Qgio7rsA07zAx+RHBkKuHg/l7L60XqKPsa78I381owy9jYljs8VUuFwuSshrg+48I
TaTp3nQdlTjF9zDHS/lC+nswnLrKv5QML5OoGJMWNm8xgnSW9Mn2jD/hMjwGUbTJuy+EmONuNO+8
xRS+kEcxnJ6Y6tl5oMY4JBpozxpop5twR9gfZAkdh8N3WCv2Ld+VlotJRzuFy92VtHbUDJHRZZTL
WmlpC/UWqJKUTseNDKiAw1Qv6Yk3rHC3EubCf11d6cxCvvHbxrVVXctBP83dI8XEKGRm/xsnkZNi
Vd9f88DmQs+05E9kRPjQNZpOmk35Xqxf8Alw7rbRomg8WsN/euHeHzOeAGoIztBOfJQ8u12hh3lc
N8zre3aL2jkmp3wvhs0elcWxRyUy/gJmaIFLYGfkDtVU1B7hGZPlvs0jtmQinLyzIdhMGIi4JLad
9aXypTjFezEkQ7K3SZm8Vfgdm33RVkzi6owqg2w0CBt+mT5GPQpm9Rgn+xmUaJuJFaG7ZVHPovIJ
iWvF6uy2FetOfkHn1l0F7sCOqOIvtvK++tF1d7IONh76OWNBbYCo6veo7X97lfxancOQTEKhfFR3
kIwYiDEs2xESW0XBjiIvpd5jGVrY4sUaj44TyGQNeh5DGvQDfYR1xXdA6pTMGuEgiHf4Dd/5wFoa
Id5h1r6NWVg1r5XIR1zBa8PEA+OZtnLU9Kt2c3R2fdKan4nd9daIKQDAgVaPi2ppBro/FnOqyM20
V7YHoulZye4IiZQZe/kD9mv/QAQwN7AghNFqmfv1EmFtNQBT/rL12LZOW1Mt89X4iXBnO1L4lTHk
f9WtVMiLfJQ4n4V/tPDqdZ9Kfs3xk+RBQoC4DRrqk+7VyEvaj2HlEc4kbJJ2acQTDEmXXA4f0YXl
15n777O/UOfRKJ3mMrtUGbuW1KEN2b4f4psc0UfiCxH5muwEqJu83yshatqMFk4sTytZ6MPdFhAz
PBSJ0nfiIsPEPhMHKIwdgDAuVpQx8ApodDcu6qKQlIEadOal2rw+OdH24yS0XnOpOkJO0HaagND2
ANc4tflgkD9NpKUfmqH6+a4PaeUAFUkfQwxUoDHzv1c3ugrTVngeWuBD4FwvXE41Pzz5kulfIton
aZCS9t/8DXAUm8HWO3v/3mVThEjco12Cjf/jYpZanSrkMaQy8D2VmdzdlaBeCfFRjqNc2CN7aPOq
GiqLkzSORnNCBmmt4/J94G9akzHYn8qeWXN7lkABqng82eJ9SspVygd56g8o/IpMDqerw3g3vamA
evmhDBbDNYEK+8CxBT4y5BjEAwQaSvOnPChtUgZl+rnBlheFagFrpUtKRmeLsnC1hRN+8RKzCaTY
5EHUIGWpjL6g8OfPnppwDwfqX68wfNlYLnl6A+PIW0QJ9LMyDvgfc1OOcUVMuKv1IEf7mzvxq6rF
Oas6/pTK2Vh1/QwWqYsU64at8bZkPborjuiyxrWmnc27846Xa+pMPqRN9kFN00X9ZDtWqySzC2Ue
wPU6sOYB4Cq9p1qOxG0VKR7ZR4v1slAJnPvpJs7p0F/LjabDGK4DjPLTDiobTcWhASsdOPwZoIxK
7HcuwHEUBxCE2Q4OhfpzSZ6lrUbLVFaUnWq/HPFF02sz2ihghzB54oa08Vp2Wpc98waYRTxcjd4O
/1pWtYcPnlllrDKZQAeU4a0D1tx9EanjA0spXRZSAXe3v4ujLxH2k2YT1yUxMhTsF2Cr1//xaw/U
1WEun3/9mUkrOgdorPwzaCt9jfhCVpQJ/GLhN37WSZ87HJYpwnGpBAWo2SFdrYfQ54PaZY1/QVZy
MBRZgp1aCCcdZWU6HUkcFcfVn540vfQtrqr10cOEyxPbm4Xv/c5Txm+UnlmTtPNBpb5AchD7wo3a
EJTXndNONzEm0OM1OZg00QtI+iykb7POlqNByk/y3Qh0SQUhgoSfObbZjpxstF2aduZENpqUgjFt
VFeSKYoUyKPQgcqBGbn8CsIHNFpolamVJRHYzJhYJHGWEpz6I1utTJaY/N3phUUYILUYvatX6U6O
J0aRKqtvmxObPtdMr39EctrtnImScQHErR5TlGuh+Kn9YkutIYBtyVp3f9rb/CBphQAj5Vdqq7Ed
FklHp78GHnAAkh7hzsYKHOLDi7mCUSX2SICAnlF4Ui1ZV/xXr6OrxqiRwzAWU8gTzZg2GOaEY6ZE
gnRfFgRw8jPo3uLOdqtdRwTJiZV36j11qTjuTpt8dEDjOkbjtxI34XgPQ3X/7wJX40Q2oE1eiO1j
mIheH9ot44FQidO+4kggrAtaXDr19BlBBFOfLviIPpZemm37TZ5MU8j29PvCFj84iXHZeSX8RLna
JN6V6gYHZGHZrBr5mnOEZzVPhp7eSNbGYaZKTagrndVsg1PVj0CgAierdHlA36QkyxYc2OBnJRR0
X1WyPuCqHc932BctZwMngwgmMR+0NPy2/XgDvYeeiHO6fOWoBXtn7dnhsSEn3Kt6321JUxn5h5Gq
8QX/jkJqeXBWLOKLtM2LL2PDbj3l/nmkwsmgQ7ukDY+NRieqw3MMQaH3Z1gmHp6ZJoefu0FZvqDQ
h26WRqvz560CLMem+Tr/pIztGtUfdcGig830ajuOF31TsJIMzj7R/rz/np/M1PmEEoRKpj3QfLdG
ZhLe4sO956knJpGdGU9cchncpAnQQoZ/6WV8w/du4Sc+Ion/tvsNFh3EEzhFVvGB5bpkoYYYDYSQ
BQaCtF+3zshKRgjkDhm/vPIlmbeAIFBPTzeJ9KYjDbhlZp/aJ5lQ/I1gT4nZLpz8SnWGXlGWaNNo
8I/rXCnNsogAvEbbclh5NRFQmkJG6qwLzeZafugsd7CIQg3XnuBvgskexhIfOog5W3lvWxXjja95
1WvKqm/hOPvyz57YFpKKToOldXdnpYJ8H10TzX44MsgVubeihNbqCNCDzOKLme2vQPAEZ3SgQzbI
JSdQKJTbBF89tcej+Ju5e8B5PgAXMfPRZys8+Xgqa81zFJzyuCEE2AcwThPUOfuKUk0NMjisiGZ0
m6+uEDkopcX4QjaxZdDYSUkS8fAgo5x3ZxXLUk3vNpL1wQLMrLETHXswCAWSBD4EJ3ZSuE+9hKkn
IuNLYbyTmpzm9qbdpKSkpgf+y/vl7ZZJedxP0J3/YFFvS8s585v6hzupJwD76N65yfCDAQChPmQ3
Bq+UxuPXE4M7Rj81OKtudzF4a9z5tjbAl5qMdaZv7epTKUoRyEfJv1K1flBaSjC1lTpSXhdF1/mu
3DsvP2lCgqtvmsSbOKuaXtt2AkQssZq9KyVF3w41iakkypU0tdMCkHUKJSR/DUZlRIKTUr7P5eoJ
4FskKA7gHcFwbAX3fHpYac713dowSHJPjopfdLUkU5Te4f0EWKqy0s56lMfDZawsr12l/W6yh3Ws
BU2Lmt5DBuCuqeSFl5O/4t02QKKNAar4sRdiEons0PHcu+eyj4IL3WXdkuUV++xY7o8aTvCUdrBe
JgjsgUoS+lzLnz+rygci7DcTDjnNX44dBbbO0FCGqkFE0quGtqwBP2CBAU+pc1yYEfPbkJld81OP
sPqsXXKbG6FQU85Cj6cajBqALPii0rqD9N2iHtaMAG73MKA37oyGQlD3/saIh9vqUVGZPLyJHwCs
y3sGsGcb7FYhNN7auj85FQ4b22UOlu+i8O8p6nG/7v+CVrdhG1qyHhe4TMnz5WpnFyGlMykmYtWR
GcOituBId+YlmB0bFXQ+y+lKKXjrscooU4KF4YrEgj+Od5ANZjGcZ93KiXXI8gwMJHFnJ9hbcwOc
DQZKvRF3qxzpwNvqO45/99hj5FyEqFNKpdh1LhFrnMe+WxmlKJO/jnoCSWhdwOScbEm9EHQmBkjC
zkYyqqVQf+wgg2yJCCwPDFmyVhUt6TH0CecexOEDR04gZ37Zu4FK41EgT+4RjKyjhYnRLPuPDbOZ
kU4eBMUpRO6PpgZ/PKJdmgaQW28kmCCDxsXrBpmoFBusQ+lpUWSiFR8rYALYUg5Hfj7kLjcwCtxZ
QM7t5saIwyh8p0jDbIbseX0YaAf3+x9CwuF/G/Nk5+8VfCqO8HBh8mApDIi7QGbXVtbWZJ9BvoxM
9qazD2B497NHRnCRSdHWb4AMJOu+h4pLzgEFiU8bP+aobA5BButca4OXNw4TH0Qwn+fx3wAZscNB
o8A/xucjP2OWI5oD4YGYQW8Kuc8c0IrMaQSQsQZfsfwgwOPPAMsBwWiFZmbZQWa3+nvcj1C4KMUM
fGZFiJzaWq7tlh4Qd8o3vAJ8u06vJPN6mrHTBSJfevlftPpZ9fPRZn5DATtP6f+lbEbzLoTwxviv
0tOcTtlB2HX0WelEelcUYuIB14+ARUv4mriuFxRX9vfqGRszBKuEzGHxY2pwIHeYckJhR/sV6fFG
oEiJOl0UdCAXjhxa3+Rqc5x1ZPE5Ccyue9LOt1t5axHFLruHC38aLwVyaH5fBdflEWINL/oNeO7R
SFs/+YSVayyktbKIa57CLsthwDSp4nz4S6vTHEN9Dm5oo3hkK6wr4grIFjXFrUV2e/Fr5jm0AMPv
AVHpox9M+QyDI4syTCrtP6L0AHNPj3fxspsOo4rpBdwgiySimT6p8p2CeG7f095YVUQUS9C8kaFq
pWtSZl/dLKZUn3ZtFBuUeKS3+mIdF2eLJ3Y4QNNYLB77ArgN0UbIS+E+hZz7LqPwwfgo/pxC4jzT
OUmHhg9CdXDpaxIlOak/ZlDEzdKyf9sDVSJK15fdet8sL7Enx0T2dNTuDUDWj6tohxXNLV/csgUa
OMyzHwv9LWYbukzPyfhGNFagn2VCO5uhdDXj21J8bOxFKFXHj9pywGvkT0vIBRZnPgCLdlUgHXO4
eeEaYE5rUYdvdTaPEGdlPSxGT65ClIZIEvnkK0EbdMbp1cV1UqxxZwM9RkBuyghvS4Oe0mLn/IVH
W4J8JiwRlDqcsXVhnkZmwfuzvabE7eECVYflmh4kqCemAOeKtWYm/2W17h631X8pbIMUiFLxCKQJ
bQwLp8dAE+CPcoDkYWS1KF/ThTV5D8fpGmR1ikTPvnuU/Pafb+fiIb5tDfuLk6J9HGsG1kYEhGFO
KZcJTMCkStiIggJPFRb8hBmmiO7GxzczoFZn6Y0wpycn21UspGChVXWFhxd82b6bvxPN6E/1FTe7
jrKQu1gXVR9RNc63J+Z7x6A2qtxaeinsGPpgitBrOXvI0pKONNymCJkJ58e/cIUKWOepdE8yxqAt
eFy+xLlIjoR86eQ/CaLYE14HIhg2j4fxPtIMU3GYy8pbrIkoXjCpFYqCnRrIdiVhPwRZl/cNoSbt
dfezZjXfGGUcs2jLN0G5cwRK0iV3rskOd45/YlOqC0/3eVEdSqBxqhDWjMFn5mkacfL+jikGLceN
T5XZWWF58yOFNJJqRioc/TVeKgOPfnqepL6N45UXimUWFQFQWqE4k9LEeRJJFVY1wQNnKiZF8BiZ
zkKRI9I4Mc1tyKSsTxgJOM9gkWl6TszLC0hIhnTp827BQ23K8UmSLR4I8M93K7ahB1FY3MKKvTF9
NfDrvLpTYgLz8tOC+yTrZHAy9L15PF2rXMLgcfWp1l2MIj3pmOpYkIjH5Ogi2g1gnKSWXQxZ/wCr
SlBXpeb7nQVznrjyCCKa1I8IKhbLeUaELTSM9Oy2aQ/bjHR4Q9JvnICzdxorGnXWo8fkP99kDZWw
W4OBGOSZFjjXuRsT8jKzRlxinClFEQ79x1GCAkwAz74pRGjtGqoUbV8JIrog7uQTN6cU22hl3uJ9
kN9+Kvc0y1k3Cfxpx4wVmWFmKGaL1tNKvFo1oyv5os5GOP4BEvZk9pfAPjBRi1jN9slIftRA9Xh8
5g7S3o4yieaADrI8mzrromEPTEiNxu5ZUWj6azVe6ddDyL9rNfbXHuAs/ZcGNb8AxvhuepCQyVN6
UQO1OKFibhsx6JYF90zlURy0k7e++68U1fuknkl0cwezPjZt8UMlQJgnYX0PvRxIlkxNqNkrgS1i
o8kzJ6QWqCJ4TmawH84z+TG39FapOn+QGX9ab9gL1WsbrCcayd2la/TLvrrj0BDZvK/uWIf5MWqw
Ih8tc1mYh80ugJvrFT1dpx9YfTQMScURY6wv/93Nr03BA/gDJxzqnDAa/+MmoY5xQXDUHwlS59cv
ghAQsQiOGV+eJ8HnQzg7KrNzxepkXNWOpjlP4g/tcE5fiM0QJrrzJpuj5Em92t40xsUM+V8x2mLl
dx3Y9iMlNO5BxrYhXkFYKVVXqY06tjCKqr7Fy5mPn6aZt+Mq7/uqMnrldRpfP58godagfGYT6AeO
pfG0QnNCfI89izZL+pmI2PnnUOG+ANB7JwFc9ZUGhPp8btKlohaHwX7y7vZQ5khZDeC3myau+R+X
2Jw37NwwKSn9IDycR9YlGZY+74/Zwg+VoQj0Os/j9zKhdwMtYmF5oUQO29BDnps26zKslrGuG3J2
5ZqTgh2nJURUWTgBNaBkE6s7lup+C89Boa9Tsi7CCReWYaEkUvreQfaRNLoiMLvzAQz2Um0MdUjX
vM3mnOZrz+/Bbmm3aRy7RZBdZBo8WIyhdTANMs/YTrhONO9n6zbjDJaAH4fVs/ytwDWwMH+xVhVE
tVyrI6ndDRQ2wb1NEOslnf8Hih1hBWHe5S+cbqK98OG0q62oIoJIEydHfQUko/8hJy2KXIavmSxE
l+jBVFJmg2yXj5xw3nb7lW2ubUD0KSkp7Qz5Gfa80Qs1NMoO0MhX+zYjxcDO2vaSelwPcK8X7LW/
jZcSLfcu6Gc2FFxGgURIdClex6xfhmUre04o5Z/yDnkwmxE3GsI7xWQ04AxPN5i2vAYlSzHgCJet
m7zZR8CHV86HJoImA1BayeHwK9w0y4+4uS8486sPi2b36wC7nLGXChJZ1OzH0xKql+vF4KW2sn/O
wKT5M1+3ofQXblL5CYN/aEderdASaN+REuYNdnNen0eLrLn2Q9w/5h4ZLGJofEw2aFV422lgWEWR
M0yUp7MmxEtNW8Zz1YpDfmMxM67KAhntifCZNihEvrJ2VHfK+SmkdBhoKk6SqslDlOepXy8IdpcC
gzMQgGLKQzErC992pOrOri7+WufnILx7rRaQfxm8WQK91WX5NF9CmNFecThEQXH1exyeMhAEdD73
IvkcsehYTUVSAwojNPemYJlNNXYOvziJH111DXneS83IiRo0IYPwjAFFbsAqps9xVD/pxz+siBUC
IcXTnIH0Cgmt1LvmIXF9qMhJn8IUNpHIlDrkkZcyYVFpLuSzOgn903JyC8FujglrNKTJ0916Anku
9IVwGghlD1XTmHxn6xmg6IsHjWx4FFKALAgIoILWFBTmz1b8ND8STIvqH3oA3GkUbGcxiYMSmytw
NU3RBFykYAS61/HFr7W2fpkJbR2uvXdKbaHByJjZYEZTYGfJI5R34t86kZJVpTUK7G3TpW69plY4
Oh/I0GFgST6IBd5LqXH3kQueNjFZevMTWRCCnM3amUT4wYaHGSFIisExVt1Y1vUVUKwc2dA+p/br
1aNlve5dnmIgMrakwSRv5bkTYE5po5H+j+GT2F4Zp14ebcGnhWR/JuoM3QVq5ak/4Fb+ffhSGlCN
MNlMjDNljYDw+X18lkgSihG2QWWhaxKCwsXS7ZIP7FwaUr4ac68MDUJRbPfGFRcSgmokQzg3V98r
hTcxTUyaruO4FnlKG+o+obnb7F/wq7/R2aDgq7ipGb7Ex7RQ9mlm0GEykllB7znZ0TRC8oEUyfto
Jj3Ze7zR31i61cTDFNWsXME5WUDVpKGtTPTcdpxq/xIKJg1N7v239uElF7rHMJ5c6paNx8iAxLj4
t6JOoS2FNOPkXJ5H1rw2UajyeJM7KDozFiw8K1Nz6PteR6/yC1ZC5Vds+/2WeSoy8W5eWWEU1hvF
OEaGzRONpe0tz1D9epJoz8mr0ZcdDR36RXskWznoxGK6hV0i/r2JvzFIkaf6EZyi2bhLtSeoSiY1
ejW2dr2PWKT664oO4EKjAzs88/4v4PrVpkUs6lG9YlVEVEbW+XsrViWF/QQUehOmvZ4rcRVx8S6P
97tInSFGb3QIK+VdjsX+NL0DvWgRlgQ1NfgczYQW18kMg0j/Nk+WO/XZjpX1++DuNSgYdNXdlkBj
QVSEq4ycSrJoLzl+/GUK4+ZHHphQ4ZifdVbEaOc5m0V+e+RiCaa8WPacWZHSpGNSV5ghZIzQY9fy
OrYqhTd2pvoHeBtdod/NJA1FLZg6NspJj/viD2Mu9+h0+qXVmjx6FtTYW20lXBbYpBeseGOoqi1W
LicYGtQ16ZEGNnBO82VZHBVTOxKSBJ5ZUU3ELANe/CVXHwhNJcJnH0JjaxqlZPWqG2v7E8TYMJYQ
RSq2PmR9t8Ib3UDB3OZ2aiA7Abj1rllQ9KfUt1CeqXnAkv8DwhDLnQuwfvDtxn+XBcgXTh9GCm26
M10J2LC+32RnDABTv36yi4mkjbBpi8G5nqfYPKUU5fmBXpR+WFHxI9WCLBfUvJOoHi8kgQmBFs3d
kwthRGVPZ8aXCIRTYBw07MUkNoc2VfcW9OIT+IiiL2TkscIxAEfwN0VKjF+zAk6DZuZw3xH6BTHX
KIg4qJ6lnzc5LKdOtF7MfC0H/BwZXhALyJ8kvTPn6nr4gB1zxyBUrl8oERBD/IoY6Q7l1MgaelMp
HTWYnktaOGt8qEdxaTwrOZwYpFoldaP3qzuxexWtjDOf35lrg5AQ+5cCQulTp+UaaOsmpY99xHY+
vuHPGezlaLzclGXHp8L9nIg5YrBuUjLvaatgn4XhA3FsF4uuzTXKxP/h71OzqWrb2ETAXjhW04fH
JtRMo8EjICGKescNyK9fyi3eit63nez+ZsZwe9jvyaNR3FFp3YOArCBtXSGFFXBFq4M/3F9ILY7i
tb8+/xX1F0Duvv1jcw5JM+Ow6soK7Bjin7C4CtNxzxL4JTSwJgXk5Uc2MjgTPDGK/JCHHu/51IQ5
8+qZmFHNKLueONs9QEJOr5cX7qHH3eCSHOUH+9Q1gKuFzYmKq6fOl4dLDa2+pbNg10sxNStcle4V
lES27VTmi85sTNo/B5IH8FcmeXT7F9iQqcXFpM3feVH1ycGV1oqQYJz9OgJKNR20bpXnVzktbGBu
n6wv3V26xCkPIsIuIhIg/5P/Qd8NvsxvtX53HuNmaqPQdPc7ncsrWeykaMEzdj9hAJnu5Gv+gcr7
IyhckAYIjgBQP8WwlLyfW9J3aRTomVKWxytHYwDn7NC5UGVEDKC0WjkesgTbqxq6II2sDoN2vsBN
r8leKZqs48yXdBTOMZjQhsyjMaELFh4C5uQnZ/Mjl+7AIKH6Eu3r8AcmPydQMXHktTn0iquZX1Hw
9LtaDBF+uW5CvVnDrx70zb8A3FnbPntQ6e+3TlDfktrphiqbQ+o4gVCr1Y9mr+/Wu/rNMa7qYmot
Wt3u2An+ZbpcEX7Mn9qB0uZ1LlXZBHNwClatJN9Ge4cW2Jg9LX+Oy++vcn/c9YObCzwlSxPHJZTZ
e//8p+CA+43utdNAU33AcGiuV1JfBlyAdlL3ZMo8SsPZXVKuEJKCGsCaPdb8ohupS5ydPHGxu+PN
C5W2bt/VN/HxcoPaWk6xV13onJjRzB88EbMG9Eya2a/1+iDF8aDfSnsDof0pxoNq+KLaXq2SOANx
eHfwSl0JcxToOoYRJI0YX8CAHdL8VPzEH+kLEF8l3tlxZAXqVC8ieqO2qH1f22TLuLDkz9sktZyq
gV1mtbhyYdMjXmroRmh4UIKMp1xmaqISTFN0He0JLylhTRlSaWThuk0dheyiAJX2u1B6pjPgfdR4
JYDywUPbWJ2EnE3dkRLKALIw6uQgUDUfdEduvzcK+NFIZoodU108MZMGJJEj25/2RXnrrPKoxbKL
qwAVDSgTT72MscJAVNPx0zEjT4OuJkGLR8c4ryCJRdtwM+wR29JHTD9XbGe/GKTdlc26UElWIRyW
Tq48pbtJkuVquzniDzYNZl0fB42IflYUunzvl3x5FJe9Z+gG3ka1LHNU9ui3RJ+AC4dNuU3tuc0M
MTmhwckI2+/XDOf9kB6gi28M/syBiPukIk0/kv9lOd1q7xIZTJXDMHr1FQghlS6mb1V3Rz435ox4
ASUEKwDJK5QiijiR5o5q+kyklvjBKpY4OGsUW6HxYQGj6BroqClATc2OtFmd+f1b2DRTMAbZUf1o
N7EUS6RV+/+S0XfT9blYpT2HxfWAD1NX2FzwkwkUnjB46+OiNfQFvHv8j8n1MoBki/kjqy1lhjk5
Y1tLBdrV0pWUugHNKjek96CfPt2fP6Iy56naK4ZiWTocXxzGZ02Yh0m7N5oW4EnyM2d5yJ1cDGJK
fWljxIFyRQg9cJky1oZhir+zZpU9ToWrhs5H2VvQghRuJE+5+52gjDr1JXMsrK7uGQJSKaw6Spkz
PQSfEBpPunvV8ht4eYDEPD+7QgkwxeIaBrlA5F2z+QqDFDGc8Sd9kHCmc33HkJtNP0KjKGK32aSW
UV5gm6Rb8naQrzgceJ+BAiwGKJAOFKTQpr6dbrOdoMmhhF49udFtfP/r2WeYpcXWCcGyssefzdCe
q8M3rhJnhBiG4mFyKKulG6Jy5hR9dIqeuQpQNwoJEtj6aCrU06PFq/w30np37ERcM32yncIY4aZ2
sYHa7rpJlnEtmwNQX7cLTbYyy8ZIGUnW4OSYRbMQwKCds1X33Fu6pIydECJ0FEeAWwdbVjjmPAwA
mutqDCHIJF/yfnQl1ieAh9rBE9fWw4kG2HwFhCtIfCN5vwFnE5BFrqoeRZZ73jSjmzH+Ys6VUk+M
f3cFlyXhPJOZd6hnQFQQLLk3jEKOFW4dAbItHbtGp/RcJ5ASCr3m0Y8oTHvVGyEOa0EZnIao4cFD
4GIC+RUd0cE652PNgSRsOee3toZlqqaAYaK6YnCqPQo64L6Urd72Apwt7V8jwMakGuIExHcApU+4
1Bh9IPDa2JPjma88CNvXYBiW6WYEf+rtHAOXMaRz6y9f0Wz7mTKMZBWkCCf3YDJ53gSlokqd6Vc0
UNPE4G9zNO5brwQGkkebK045N+tzGjovXRM9sqJLAHO99qa4ExT7JoIjcuDlt+/Pm031NeKFSz6V
C+w4DRbYIFyB5oe2J8n6Av4G/TjvunqppKF3Dtkqn1C1MH8cOenFBokHcDT0kFo75vuryipKTQ3q
N9puz0Ij6/7g4Pjs7v8kgB//ztG0newGf3/nFJDW9kYXWUHZRIZh/QG6CaATAVn3te1y+sNA8r6T
EZtxbIp1NRC+pGw7n3qFvFDB3kNErfhXaiYwlnBMBVzDan9/0XvNK+NKmSk2mkLAdicxxpeagrNV
H0lnjHypKBKuXqAg0R0131nhvyU74D9QwHJRUtdQ9sFnNoYxwHkD3yER8OVNK+rF4093EWsmGr4F
GoJr0Jz49RUTjK4T2xYQzrL0vUU1rmscyUBs3iC5uZkUldtVItGoONQTP/vGsmJlsF/C9Qyw/LCa
Wqup9BPYLtOHfrJxSmcRIcD2wyY+d3Yr5l/LkEVDl/NeQ3Ej5QH+E3Svns+k139YkdB4LG68GpzL
eM5wfwAEk7Dq4lQc3ftqRqLOOcsdgCZKNAR32bPZ+D1RWsvSsjSfRmviKWvI2/k7n8cUGZrouH9R
Lb1tTkuWX/b9Jn1UCRVFjbeOc0yl8gfSte/Po6DM1hM+7e2GGaMo52R9zBNYAHoXV8UoI+IQXVF/
TgF3aURDDjilrUI9t4wFH5PSmsFqK0XiH9OJCqfuc9DG9DTHcISWTg0mfwG0v5G1ITyHlJE+oMBM
v3nAyRkeNtPiC6mQrz92x5Gc0lzm2PrYoOkTqmx2lPeod4Y6aB4yHulkGfgeVOGecjpKVgWQjRD+
hCmVxSIVFk4DWnyo9MZ1+8HOHTHeOSKxjUtJa7JW3o9fuMhgjjS0Lxmv+pjhqzGCTOPJ/T2Gfr//
aFka/ogm7/nzMLLPGUN52WUnO2nCxkWw4wZdPRZvzvbx4WlN7DeDTUJTSFXTMF8J2lqhzv4f2vlT
OjrbHyDu78HtVNTdZDTe4TpvSJ0IXhUq/h+KiB2HfehrI615yCNuqmm8dh9FuUPSympHfdkrVeT+
ntzskLUqRT5cgNY2o8RxZ6Rpi3HSYSt7XcNZsbxfFIYgvqqjp7Ny2zLfAAP2Vqkspn1j30/A4av2
96bwdaycL/O29PPpKYWGT96wo1MZ8Lk3tY37cyT9zR0/0WGbgbNOM0MYIwKANRQXkqqCB+oGdHz8
cQ5Y89IwZPVMZgFdp4cuQivcZmtOwKPf7/j0tm8bx4c9oe219384mRo7aGX4Lj+5v2i7+K4GuGSy
Z/SWu6LSQeyGA2N0eZWdfXpmHziJukRi3TQE5VPrTYxQtdBMLbt4/xbBKjbugL6PINvCdXB3Aepp
Cf1B0O07dGkdCyZ+nc2n5M5rksmxHT8jkJxVzDDf8nBx2FDXyUVc831xMhuVuXVAX3m8Uopg8x0Y
cLgikIloNYHtGLjXWWeSeA5lGijdvd+G7FjhWki/AHBsD6503Wi/00uNVPTthMNdJkbagq+NuiPw
S9CFj31t7R13DSSzWEGkCKPbW+YmgWTAgOppSp02GBwSLqVnp0WMJzrJ72fphSCx+gQII8zg1Dop
8+BurlYFElQkI9YnxfCI/f43ernObExI7WkuW9iomFIGkFNemovfHkMX60GFd2DcVqHvS/mnDkAM
g9nOcuc/d+Tz4t/dFn8qm6v7owUdGETQ4aGQ/4EI36/KT+QVS5z7GYJgJJBAUFLjqTv5q8YYDY5U
I11QUg167obqy5TAQJ7XKKqdovOlMMXMxSO9cB+j2caVpThIdq5aEhQHdmruyjDXbMJcZ0vSB9nD
/dY3/RAuI4FXM1mkIh0Wjbz8wDrHU/D8HLp/y+uGzxtPSnN5t7Fimh7meWa0mL0xyohYOGsl8cd0
4AxljZaAXENyRwxt/5OzazbEHmxpk1+C2zJvVByH2JO4AHz6LmTLv3ZT7cN73HJ2lYVhqWxtH26V
m7aDD0dXuS2ZNjrGImm7UpvExm1g6bRPu7x+KhncRig7ITTvb0YISFzUR6JRrPay61P2TlxozKna
SgK1WBw2D5YBRYk+6M0kTpRx7S9LUrnbTf1SJ2D5Pj0fZNUJn5SWBfuIrVuQNUvtp5fkxJ/fRjSb
6itLf/utSP2/TbdYfEUtw9u+vN9A6IqfDdAwQrdgm7pNaed8YuJ14rziqUIMytqW4c/4roWnaHUM
OakEQbVWBCrF946o08Lcbq944h4QYs7aONu/wEWRLnvf6HPvr7rzWlZ0+r/acXMV6dMIA3t+X5xt
u6HMnjY76AMpV8/JLubleSN9VdXpkZzGGszdLwk3Pibtgyr7YiicSjoCvFEXLMGxP0hZZHGQDgOc
iboEfS4gckmQ8cLen9VXdTmxJPy9gMe5zlqwi6cW/SKIm+E/3E024W7X91hRcV5TqUgSLFBAw127
1IwqPPwK3WXZiAVYxWZEhq7BcBH+qIfRnXrJvLOHWMqFKaNtU700P7CjsyF080aEsWKqdkgLpGx/
q9TuGjL3yKTrsF/3pwiY6gOMYv2drAOql+iHX6L4fktZ1qEqmfUOTJb2TSuqDYVeDZ6aU3Hf+i4j
UkW3ZwDQpG6NPQzuzz9Rs84fP0EFUbzAY5ocIwvvhUL0/ixE/HvdKZC2UnQZ0GNAaJUAnsGgKL3D
X0rA9yuK4yYp2VHAk5r33ZzbFPpf2wtAxTjOF059tVOO95iCOAk77bgdOGtCUsHcNkWVe040w5yg
Gn2oK5aOld1RieAMfARJ4v85GQc2YxE5VtAmZZ136Y1OPu8fRQXJDdUImptvnBYNhIk12QKgRWFs
57BXHFdZxsNDR7wj6hQ6KDfRvJyolkMU4VCru7YqJsTs5fwyXHRtgjw02ToPH+8lWbTQHVr+EVnG
kHZzIxlB1DlezBlH9rgzReusqKjaUzJkNaDmO73NVSljwiOGp2U/s7Z2ecM5spSnGeWrz38kqExD
WKG7/cLTE8ySOVY0GtP3CG9E1XE1lqCii9gP0a+2IqotQD9dztUlEhDx2m4FySWJzinPbCh2Nz5P
JHCeHySbaPxd9FfKu5QSiZCW4vGPjah7pd6HDPQLOBFTXUvSPrlMRmqpQAS+LcUg2qHku2bj4rs9
r9ipL2VNcD3Ea1bZ04tK/8YB3Db8yt4WjhJcaFsPtJYVo4aY6LuwcbCGyWFNkdFyBsHO0Oe9Xfkg
7G+3WIcu6fFQTmhEDaDzpSoQTiCqcx5jKIqoddesAEaVhi0OuaIpVV+jGRTNBBwHbTkn+6fuKyzg
DBBhXb17YZIIYiQ2j/uxssU6ZGimpVKs1YoaWj79q+VrKy635AWFGqxgxd/WwOI0v9hyVKIixjIL
DSXQ7CdGuL1i8Dw4iulRkkrdDtE7DDId/G743vOXvYNN3aO50XCtGWxToMuR35c0lV6yaqllpxtD
aOHs3Vl4qCeYkveoYqfHp7qQXwp4UVbveCclhudlXZu87YxExrtlH+mcjc4F6dc9ml8pDukg9qnN
S6mrzDB4WBYeHMNV0bcDqKC/b+0IzER69Cz00OyiIvfCJL2nUpyJe3SqX0X84EP1jzmL9262DCEZ
zjsPHcEbfEPm0oMMRl4J4ITH/mDGpZgNwp09kBDHTJC2j38MUxLHkRbKPnm7VbXDbiffEHeV9fM6
fVcRanHrYYLswmZq5mxdgokYHtOwYQ1GlZn3bxZsue2f4D9IkEk1qnrCkIUIYCx3qDYjNj7xsH9B
6eQoZPmlruoxmtSISHmmAwJd9IM1A+LywupzVX1RKrG9+0VTUEKOO7tjv3k3Al9WKyaNKRGooCZG
2MadOVSeq7MWW71Vyit68FTS55F7VAX0pRsWtCj+OjnAoUvLGGcl6tI6RZmanQ6A7gsk31WIt6wQ
zeDrAODjkaS7U3hJ1py2kNAFuyWzEENdh62pqwu7yCfm6aV0aoS+9KDAo/MI+64PXjMGnJ6qGPw7
y0oti1wv1HBNXd65txzlQ0KUT2QiVaIcrychNlNCKBP391bvIiErsuj/EbZhxmTeIFQbmEIuOeSo
eP+pJokrBqcdlqGtVxdyql3FR+QxnG3OT64UW+PdvfD4QBtAnKC479gIfwHhvnl7ZjQd52TyFdun
xAjCa+cNDo0ga83dbqiRqwm4fg67O5KHGp5LVw0oqBkypbLrwdgfxgIUMdihyFfL2KYcEPGK6DmC
GbicswuIyBiApYBSpGPZNON/JYklTNV+7HrbdiA+/UIFrvzyvou9ueTksq/GLoKJzRRWuG/yo8Lm
lRYGQEE/3NqLidEdmoYHEnbnEMsDhZIvMxUVTyTaBkPBA2GyFZiNmQzXwQkUMHsBPNK5DgQoYzXV
rWgjvv2yYKRy7IrRdfPMeFAwPBYBl7/MdcXbW33fCi/3a3n85BdwCrU0zlL3XFf5ZvVHf4kQZES/
nm7uJcXVktndpJ8wOeJXIiBrNQ9fmnC/6dZZhBM/wTepZGKu4nOyWzoFtceIh8puC1a0TbSPT6i6
c4X/GpCphRqQWUqqxtU0v2JUuWs0arKkHMkdZowLa98tIglwrZtfbz2F66LLmhYqH7ohIphEnDg/
QSvxXyw0fzf8sxBFdaGNTtiV/LxUQJxzijrOWQbBDgNpOUS6fJpKj86q8wH+jyEBEeHznpCiPeZd
gc2aM0QPzYyoPS/bBfoU42vHF9KhauSfeH41KN3M8JwWXjlhTfnVCiB9F6fg6K5WZf2mNY6rRoTV
46glZdsHdZcLQGPSipluaYl4jA/4JNCobI1/6sCwRkTltG/m4mQSPoNpr7kFYSUP4r6RMGwuMACG
0XBuXYAJYZ8QdOLq/z5hghaWGVL8J7r6DS3pyO0gvCQgYqST7uom2kSORPCr1UsQBV3LtHsTw8a7
wtgVEoIVJlLTfzkpM8Hk+q++d0giSiNycvFjlqscGUbfRcaEUsB5tEAXcy2+pLGQprXGrJhagSFd
3CR+lAo5OTFD/7mvgt+HvriKQ1gaBMLAy684EklT43Z008MAKJZOcMJ3hZAyuXGDox57YWTRENzK
HPxbz7xMxWnVC8aPWiVmNM4qH4MD2g0t07T0zzkZ7WXfmibfuLV/Q3SoJ8slyMmOHstnJ4ylRcJq
w7QAD11EzC2l/AvhAUtq2qYVXN7isOgBwkp+HykUWI1SmNv5WFsgz+d5SHeKwovuanWXp6TNYBuw
MCVM4KUxH6YHfe/9GKfcW+5zfVxZ1geldh16vDkIfbLIyWt5z1U3ChyyS9G1dlmwzJImlLJn9xM1
szN7lU6Xijji1UlqgXDohzeYO1EUKKrTNCOy8XEK3acfSmCHi+hFN9PoxH61oKepT31qLkQqhxf2
tu5g3ldey5B4KbdpYDGaDiBmGDrQZbuP7X90OMKqRJbDClxtZ08ym8WxhKw/DnPbOy9ileU+I8TJ
+A2IS3bcqpVNYt1xDdGE7mjBwsWtREnUspf1EnKrFC3pifum8pAyUNHKGDELVCEB5WKn0s7KuCNt
CxOGqxxY4f65Bd3d3YDQSQYIGjGGlgFXx65x7FPiHPQ8a/PdL3BWDEvrEnZhh8Mf7XgXYmmdK3Qr
SqDGs14Ti8Cdzb54YFla4Y7dCGISZN5F9uc7AwFdJvmftc3nCiPVh85yLiZewKOlT3bVG+Qeiafh
H2PHMQoLjBgzTDAvquFVHfKMSLHKtxRgdowa10Wm5/99czeYS11vikBgENnkRmEFNqHCB5cLXe2t
olBM+vmTDfE8V622iMLzIfn87ehEyqrx27eHEvHpnZO1xVTZFHZI8NRghzInHUeYwLoZ7lAKShUK
Tf6kg7zOM/2o5gNxigdsyPhhS7wYKW4NpfTsVQ8Q4KMIST4EsO45n48uYBHnQY15lDdqqv8glfs6
dvC3aZIGF2PftV++BRo6cvBgyRYqmQD3BMVmXYb+H6uuSUb+myBipEYX8GxzcC0zyoNvleKMk+Qt
o4CJtfHOFJRmXyDh4NYuvNP5eza0OSLOXonRpd93Lr9Jk4+yZT2ahPkNuCl1f6se9AwUqLIG+CVA
mKcO92KAeg2kTIHQ6Bu8GRmLLqUS/H85F8xMQPI6ceSZBf1gY3tJ7vFJHh7A34wNZGw2te7U64kg
aQcMox4fXP3LrHSvbg5u154Y+iFaayMdTRtun1+i43o5+W99wCOcs6Aa+BKL7KrUDeob5i4fztBp
+qJNHxAY1NnxokKoeJHrERtRfrozhkW+wSVtSq6O9ytuXBZHZBrxPiw884bLSv41oky/OrcIDF2s
/kWgaLvZY3GglHhGqfcQ2YuKyyGM9KFOcsDUWh5QEkkKBCZu6dQXcC/Ohecxn+XTAQoS/91cq1yL
S+S8jvZYBuVW4d1OzAdC/nXjjt+66TYd6wqL0kTEnMchwtMSQWVnlVCf2TIIOBDKdxBV8Ro+hieR
9r24WiVgaHYUNCaYTd3YEcgXbBAhCoL6ri7vPg8bymw8YgCc153u//7vNpvi0CVV1It5fmURtV3V
ZvnQGrZry0Ny4MlgSkm27MCC0K2p15B2po3f+21M1DNZ4tgPtkrahYN9GoBkcaQi81KfC1bSAmdG
ET3IzzLX9JVZ762rTNc0q58+Dn3aCatPwzL+ibzL1qNyVKK4CW8c3Ht10nViAVIftd+ZP+lTc3tm
o3o5Jw47DJ+SdyFzqLUyinWvCdGJA9ulZHqG+onL0DT+pGFtlOYp2CKzPrHl/6bhQnifFvqkdF8a
i5hZjeCmVUutSeabFtCdxXDxK5sq1aTCqreoNWGUdG+vL9C2x4Cwp3oZgXFA8gATiRlZ9W8zGp4A
uFl5Xbe347g3/FfcJQH5w7fk2XvAaScUIWN7WUHC5sxqi9Ih6gr9SEqeS/At2JmbpvdyZnzz7Mon
Fxqa64K1khTwERu/EuMF5BsiOK+0pEkyu9YwFXGlIP0XHcsOw+hupE3Ki75VKLUpumd8CESstkL4
2WMc2NxzF8eZNLTfTcYFqtDMiiD0GBk8RYTNaN/rk6mUPNpRs3mFWXp1xRAmy6HbAS/oytcYpbM7
CDG1+aq5PGPzKRjw25kDUu6UdfRhopKqTIXhIM3x5PtywhZCvGJjLDmEI7C7xgkFKhQQLhHDBlq8
LV9Ef9ebDYUCSSUWmtBpTznlFNFoTnl2D4oT6LVmvy0YQfiReOp0tXGwBzA5g7LtYF3ZxXAdjORx
gDyF4kxr5RY6jFmU9ZLIFogieXAoaqyeArxSb8DhiLTnZqpk/H2xew4cGcLIgimXiNccYiZb8Rmr
2hus/7fA2lOE44+5hx7TWoOj9ld/qxROVUZQLD1+a9kF/baN6fgZ17ncZZQjNoVX77ZE9/f3MzKN
IHL1pc9oCBT7dnWooXK17xIEKJ+NzK3gWKzUiB9oe/auvePHwfhRxEzZpaP6y54xVT8HQQmy1173
YGyVLhO7tzKaEmQOLftAZHzrYcx1h9ElnA+CVZzf4HJJkvi2iWPXDmPq2WzGic6gQU1E3gwaGqoc
BKGwFmspo/+HWnpxdK06i5KtYq3qY85/wpNnvpwXHfT6xbFA4ill1B5HNLYi9tCuzyYCV+pFXOYQ
pyH8dJCjtsyDq+Av299bjo1PG4WANA7rtyQS9EbEwid1dGpV1UNGC6ulXzo87iOoA7LxIcEU2+QA
Es9iRUu9kVajX6TwkNvKFDtIA/7hPVLIsO0uO/YvsWUrWHWA7u7Y2AiZ2GF/2necfO882qj5nC3C
NPfLs46kGa3aiIPw3DA2ozK6OWN/79OfwaWVN65cxCmHnry5imzc5WRJdOFErqGHqAnHmH+5QjxH
qPe4AKabmHxXwKO4kG5ZCTEqCEJyZqACmNrnYZYTcWrUYUzWc8B8zJKRU9vLcIZ5woFGDG6sZ56u
Z+WUsXHDKQd+SWwPOvtv+r20Ti5SZqA5Hyudyu2QBYWiVk6DUdvKsYSvZwrv3VHJ7mgyVd7ty7no
qyq3+NKhOOfG1XaNAoujQtC9HXICY1YiCpkHYXmpHcESKXEzbc/tOQfd2f+QlL5djMBuR9HJyMGd
4xC7LeZJ3Sr8EuO1j3+FxWtIRbJ3MRFJCGOUE/WP0o7bo2DNKG0eYN10vt5i81cBYenRtMDiMgup
LTBe5aZtRmPKqx24QfTma3+PVyTW2Q5+XIb+ZBlsdKKi94fvM8RmTjqzxobhh93rMWfQzFRb9fHf
FlUMKnpnvDCdHcPz1Pj/BqzNh4RveZNsYV3IgIhcEWW71LipWRKQH/p6N8Nxtp3yM5yHcWoL+3ZE
OYKfJV75RfGnVFlKiCpEo2JqJ4tEC/PrRetPky0lqKQVji/JEz5vvQVBdlqbtowQq0pCv4tOKPXf
ynrlcjAIBEtklJAFSC1r6k/31PVMQLx+MfUeDhPnt080b8UvIEQBBs1DoPGZHVl8y8VA82uTE25L
APZqBjg8BN4dOsLv2d4MEKJuebtsvZfRYYToE04bogPBrLlpDA1eqXxBrkQ7xEZ07rwJj6llc+NE
6UdNabmZskokbsFneDqti7KpiYSiYPKFvXlwzfPs3RKBAAHub1YpNK/kRw87Emkw0nxdd85o1sqI
UM2I791AM4pMLgpr5lRyR4gi5DTe65ynV7LTN9GeelZjvsa6gmFcNS6WwiwIn6q2p5XfSkml6E4S
T5gjPOcYfMqrI1qRXwCG07ZLAU3mybOoAAcGlIqqlNeYeLoAbgXG/LOhP9fXAjU4234H4jfpIihT
U4FUQGJmGp6jjsqQolpPVJvccN1kCCp9aXPAXCIwURr8NgZrYlN5LiGqhIi556Jga3ZkMIM6X2M1
rm2y/LE2IgwYhBWFD14++zWjYJV5Wkx14jEAMjGPeYpmRvkN+K3s91qAbWtcRJOrd3+Z0vNgZjwF
yB3/PUaPs8bme0tzg1VQnkicRy7Z5THjLGVeGBuUPDHb7h3GB62ToXdONBqa45gsqFiJ9AADjoBb
krYNNQrOdFjiDGl76s+90lNRslY5OkDtVIOk5Lry4y4g2XazEBhTb4bUwlxlzNRbASODxNC9sG6m
w3DYxqH8HMQ2bRqbz2L4csPklGFWZnQz+2cAXyAHBkBr+GsrC6pcumyfRk1u7cGUjuIuKAand23E
ObzE81ImGSAf+OKlr4s3Xs87JiQSG33t4YlJXfNaJAvWi202uNwGUDjwV98R3vQCmApywEU6h5Zq
qoaIBmM/CNy+oFWUgNwmBNWNe824itwz7Kppcs04bgX2SPh/DKiPwt1cC7Sdr6D8KMd8GhI8AjN+
8uS0cyoUUXgx0Qm+8g6Rg61m8bpf0lBXz88otfpY3teG6ALaFgLzm6gTF3+aXaQ1oIaFEdWdC4Hm
5tjxbvyca0ZSyXUwiabVvKCQvoiyAifDyO14FU0so8C7wgfUkRNHHk6rMZgOHf7YJiW5/rH0TMAL
VPR2dxNt/196irfjhw7ItUL39od+c5LohdFlD5dRSKU4EBJFdYBGzRFHckcVby9ZqT9LU447PSaJ
Oi6kOuTsnyFgQUO4atgZnzBaZiDEH0N1Dr9iJFwXPUvHk7UAQRydctBJ/ip8/f708lkL1ZR8PyBW
ciqNDCcViPI7AmzLgs8XR7aaYvFSFNu1fGnLsMGZGGXktbCCiOwrQJBkvqMmzBgz96JQ/JDzRa7v
Als6nt3itCN/F/ubBEeHCeXxMrkW7HO3nQBG4VxoilckUAlT/cyeNwvohFIhcMkTCXC5FrgefB5w
1z9E3VBDCRNO16Pf5cb6upN/4SX9rQD4Fk1Dbnens571jLfeuU8M/2mxhgvisQEbn1ZXKIljcCbZ
s5bqwneBYR54z+WeWvmBGl76GtIjrP6t1wBZyssrxfc62SWxNCVMUYvnt4vp3DvHF5rJY23nfXO9
M03a6jtLNnhZZgKtt2GYUYeZHRyIemy3uhApucOKnaXGoBMkXTL9UgOsBnex7fnpEjz/kDEdrN88
/UU/hnAI7hKrVNtg3zV64IIiOoeeJI8sjBBn67QobdsIQSjWJIXoSaJ9zvApmXGoKyKAylkAk0mm
DYaa7MwXrVfT53/NShmYkWObsTiYtqUiqvclInIt4/rw5vYC/Xg6tdVRf8wT32eIZtyDiX9MFXxD
qwC9tUDFlisYUMbS3CYrC4M9jexexkvnLXfvqWF8n+lnXqrMuo7/YY8r3ilUPHadbyzpHVso+xIt
akaukcZblY2Cnp0tOhetbWt9zm4TC0gDUhQCTeKJ2E0mTR6Pd+A2dZtagGxnPced47+09xt8qx25
+iB+I9fx/rpEokeBau/MxHcMc0V62iSWFYEPntxuY1+5vvrIQXpJf8/XU0ngbdP45Ey6jj6DdVXD
SgarTpRODtFVQeXCFdsbz29fEiuF7EykMV6P7pQwGqMfdR4iOzrUeHFc0rtCjSelYhXap3ZkxezB
qZc75vMd2GMUrfqNbsNkhhisB4zKXQyJ5b/3HbsSMbCpGcFMsxNLaJG5FDkwiizMkFXZeYWFccJc
c5qCk2CFmztmMNzyBMELp/6i74tQEUnbZT/sGfaC7mmI335vbYuEiqa0mCuin6iNOgSxKdCQaPae
E7qvRPb/Hmlj12guuzIPl1N4eNbJ7t5/w0SV5FID3fTssKWxdH2bPnUOw57zJYGNfdPtlbTiDCLI
9V/JEaPOt30gG08Zl90bc8ljMob/DbtB4o+KEQV4ZJAYbzNyEbfIj8hic3in+mmIOMH+JuPae5gp
CCHaK9/k88O8ekp5P8A3s4hqDg/IFOBHWZG3w+nNhYLtyvb0yZDJAm94ku8M/tpuGGQn3EiJMfrX
uZ/1b7ZaWi8DTjKy8LCoLV3Fg6H7JUfjiKuGDBcspD3grNGEyMojRpjBzGzbcfVAnmNp1uvMF/WY
Px7I5l2mZIDg6VaLIkYwRN5pMRRbkF/1BvWq12ur051ScXV8mLyWnF0e5BMUN7kE7LhqNzotvlc1
TVaNEVZ6OtXH/n/FSdP9pUEIbmO/C+gNwQ2stLNHf+9WE1/lBRlbu2RexT4RIlxrQb2IUiffstfa
ocQHuz07A8LFuiQXmDykw0rs58K+qToJlkWCl5FRWvpU4xDRt6Rrby61gzle5RnkeiULX527dVlF
ywcTmtEFY/f8JqV20upsl0i61uOaI493qE7oi5qngl/D8KbpMDsU8pfyYgyD484N99bCZvd8s6GD
O0zsuk+nzrBOzRnWO3GHFqUlA0um799VzytOk1dnk3Ufyd+OaD3cES8Ee2HgapfvhNJo0u8yN2fC
2fxDYVvIfYeYNV7Vuib6IyWhKOJ8OBE86NdNYGpNsCTpc+fqFNAEHV9Xq2fhCsj5GWdVd4Q+9SY1
RvGJv0lH+DjllQRvGr5eyD0UMklZrBXlQKeeiDR2FDHet5jcLsdA/LdHR7mlBz7iaCEUwwDfyWw9
c/lHTNzMFOFtZYRYFr2aut3Y0zA7C/Zy6FDbNOrXOxDqUjA2RQWCJ0wyyoFZ2WJ32HmlwNKEu/Vg
kmHSy5OV+dS6ZvrdajgjMx9cMB5Mu0iye7OqtbnOIoAOnpsJRW/ZfsO3YxDZyhQQdp2czmT+/YeG
sgjNuoAsOlNSKcTIu4D2SIMl1uyMC90YK97ZKx/lEfi3RYcYqClzg+guyqGy4NUnks2Mdn76sErb
FNhjBCv/ZpssGZY6DmtYGP2biREivVKdfRcHqh8zh77sXZYWd3IqS4Q84kCAAuNiPr7lCXAMGIMh
z0a19aw/OtsRzEgZ1tVaYETj9+k8SpUuTE4lPpT/DbWe0Ow0sz9JC965O3gtWXNHmhdGBdoZUTVA
+e8Sn+NcRrBrJW7jWCtA3iPCwqMga7Cij+LhmR9f6hhIuSwyo8baGJzvDBX/QFJwOwR2pkc3tidD
PJXYKcYOtxs0DWAhSajPMe6vS6Z5KLrnBofGldV3pM9T8VISjDF72V+5IThNJbt4K4IMf+b3KME6
eRSA+7ceTnmayL7I9l4ptIvElJGE0xzyhfX52bpXwh/QwPVxRVx5N87U/QCVhmVFwQjn6YUqqjcl
hUqSGI2J6oy+RyR/4oIO6Zk2MmcFZIudOrggFymX8yenl7//1GltLta3WgmxeD59cz/DyXzf76e6
3ObYS5Q8DFxWgQSnazFvBFem7H6DJygaE7F+gSe88ZN+k7RVqZn90DCe/ptlL9AjuLx+V0oisrat
gpR23oUANssgbhpBK0E5JjyqQdc+zWJcuhTisq43Uab7/OPYo5ivL00oZJmhaTG86inDw2Evu8dj
BCwO9xKd5GmVUgFeL3WoLkIMdodWjcZFPwoxv83KmbfZHZX+LLiVLe9odfAMhZH8fp5xo3GaQr3z
EwJukX5Ko5aBnLQxqX7otk6t9MerRed134m789DgsQQtWIr97VdYGMfomb25uoUswMRES82mGrwW
PZK7MnF3Vq8VjgjRBqMtxrxnh8+zagaVujxlGMK71ie0HB/Yp2mFfp07bQRY9uI+AgEebIlnAerD
mTlYx1pF0HDXlHhifdzEgZCQG3N93P2b6i4bfxX1otcUTjg86wbUSqOqCVikFNCheHGogdVfGOLe
5V2Bl0jHAXc9OvTLkCWwdnoENvWDXnfOoLOs9Ehey9ipwKQixWL1GZGKnhVFsjK874x2ZnBp4sQ5
rAqEsF/AeeUlqLEq3itocbHu7/7AzCQaEHYlVE2jFSn9gzrwvhoCu1lkcyIlAThhnE3QEhjhsNqz
Nycf8MpwH6K4E7XHeFEbMemxhm70Al6AY0seJiX1/iV8aMyxAP64/5F7VIHmwqLkVYvtTZiB1edg
AYWeZyFOTMLMc0zgpmk9g/o3uLMgxZ2E4znexXpsMlivxL3ARN2jwBlPob/uHffdHfEus5BwNg2T
HmD45f897Io0ynIqbIYYKq74SqXHDoglDtYHcrGhKHQptyCiMhLrFh7VOwAOcATTvdi14N6ZaoNE
JAwrsI2cvKvZHbDbK0J0vuklz3W6UQdMfQAS8RisWIXBlz0d5Mj5uVTQ93LQRF8YaqwhlulyyFjy
3KOD0q+TxM64VID3BOmztzspI0YJuTiyXgegapGrIvzqfTgbdQUUEEPoY7eT7GPjtn0vJt17XJwj
VYYPGIlPCWe3hs6JOm3+1V00SK1olE4mYX/uODez1i78v2ihqiZ+KfSKKVpvv7DiZGJM6mxBTrgN
6Cqo7bnquRuxOkAgqJOjP/2lxnD+/5KevJ6P5wjCQxSyz03/VVQT3Aid5f1nookCTJ2LnJLjAlq8
ifzTmXHq+FslwrOfofyloDPg6UA8NjFti2s8qAej0/2XKz3DcfELoHOdV9ehe+IiZUp75sE/si3d
4mCkfz4h9eIEg0TcJ6Dai2RGb5TsZjJb8+80Wx3hBpkuDMVYo6SZQsx54sn0+lQk+Xn+4MjgGSQC
sRaDIHiQiNWFe6QKLTndG6Un7i5kRD2Rpo2ps389pUXY85CmCPvbDTiW4IiTe4+xk0OasLOwQLqX
nQwHafl2rwMLfDHtFQCJ2YlLqSaN1JT1JPdqSorlPxEaG61J+T8t8GlibVqxVjtAoBcC+oE8D9na
9mpYebXVdk5v1m05h5tQboGTLObla+1FmkBZv8I4t3tV5PfzrplJMOXH2BuBmIt0tvk2kq1S/hD8
GBFxQB0bY9qliwKqlAwrCi/xt4pPyJLUgiKLVsu828CNqSno6uyZ2abpuantes2zaRvhHnNbJh0M
/scTRuj8Gxc95XteDjdGD4Z962pea+6M7HfXtknWXIWsjqVIh8PmDyWFj5oX6zc2XxYELlJeEclD
hQmKA1cuckI2Psc1hK37DfgRMuHw/Cb1I8tJtm5Li6hTGVbTvWRt3ICY1IylusAEc+0wbMDKWoqO
oqkA+CGc1+r6zddE3Ee1Qrx4K6DSVNQBOFz7EN18MJV4d0gqfpfq1niEBIuODYAD+glK3f9mF+aI
SEQlcAZP/NacIhqMJu+J2ZSVRpNfcCgDWROXIdFToVXuDNxKw5mvR7apxoySIOhx4GP3WufypZlQ
2AfvhlogMfoiZ5SfbqSrftIjKyM2FoiTu5XZlSDyJUSWLtSC8Jtch2uQ0z1o5Kf0B1ZJ4cpQ3+mq
DAfFfjcoUJDB49tcFlFrmOcptymQoxDKB1lYSmQjNM1JnEUekVuTFKf++MuROXDgmAkcrgh+pfb7
z1iSq5yRWITYr78mJPDeC5pIrto3Loi3SkTpbZarzm5EfgTeSM/ylzx3fSlw2WCjCv55Zzxl7lTy
zcUoX8bzF6S/7XWpnhvGbBpvSpkvN8OkhuCgHc80N9YX+ECPA5ivM23GxY17vuC8npeW3JmE8c9u
GPHNQ9u/1PpAlj5X/PuwZvUBmnoqWLdNNn93mCB7th1ZA9/aYfVXqAD9CV1tIl2yTEqGMn6Hrd06
HUlER11XXBWK8C794cLPHLdmXZWRbai0W5X3ld46F/2nbzjO9QCggkds/2IPcS1M9eQ4kWeMxVCB
vO/t0rV9Tx+A2sLOpQJtjPqYIPUyWqB1jkAqfGrv/EYAxP5LrjiXIdb2a9/F7cRlul+gBypaQq/N
znog/Mks/iFABcTBkDxWAXlj5uVAD8afnDNDPayNab4d7q3N3pczSNSoL0Niuat+ySkDylBmOcar
9RNMCRohYdvhO/T9IeLNl1waJDJQwumoIDgGpuPWiMBHs1EdQLVrWrY5pIW30+Gpb/LPD/LN06iw
MqlnnU7OhPzngMtpwghBo1a3isVo5BmGOCFGWTFSc/q4mYWumES13LI9UABZ/b9JoD0o0UAdnG+z
XuWRGy3Xf6Vc/yF8s8mCW2vq3sLyeXWTWLmFmiFlO6SRk9NViV/PE2rPkmg7KUCWFQGuy2Uqdmuf
rCCsi9zA4O9kAp4pOiPqooafLQUVUTKoigK6j/P5K/bnv1aqyIdHIPPINxHrbesbhuYGBldB7D4o
bPNKj81NZkpAxkQx+z1jjHiJJfdZNp8APZqniZMqSqSVr46fbVv+6ETmZNmUfsQBzHACpa7cw7K1
Fi62p1+l1ghWZQfWJteIn+MB0FF61GQIE73M/7sSS0lKgYdttgBsbvKsWekNXHC3bjt5C6q8XGZy
2QCrmiNA1vnDkf49dWCj/knT9C1x3Z9rqrQ16LDGRUjPlxowC80TEYVlMHr2CSjJORzgKSUbsFTZ
YOK/sWLp9EcjJAi2pZw2I1UF+EjR6R+v/fGTYClZyU0nHMSv+XVG3RYb12rAHg4OO9gosofD/8BY
UvaLsPUgJJS+JincvMeUsmY1Lf99JtBwAe2YeEVVDA8VK9usxrSV5eyNtjm7hueEIswxK5ThePz9
6UN4VREVp39DM3tJfe8vKxXex09oxfO8Cd054HcQ1WSsJtolCN8zBj2+KB/AVSq35u4Nj6G81TlK
xpB678wXlyz74YUF+U/0UjPZkXwWn7feyol8Fw65IBmuFNPyKkGUNAl7LtQz/D2PnOUwhikBlsDk
Hz8lXAfUbbW+18CMGNRJU0ZpO3gxuxqO7KIKhVirkTw/d1PTvirFsvsAXe+VYBBsfV/CkHH4C7e4
kwP7r0Qst/xz+Y3ZJLcpChIMRhAnR1K58zP1En6LpyN3Jfw4OTTjL+KJQZlYf5Wc4iKqCeJjQdqs
UgCJoX7KEj9IZt2C7wSIkg0p0IlPgUD0SWOxGBxkDiL8U2aM4b1B7Tla9ojMvmOEzyhxDfhJ1o88
BiRnrHqsd3R/hHK3BNVd3GDLe6gU4NpfVIYomQQSfZqIcsLLWPhXf049MWWB8tRYoMSr3kfhQgeJ
Cw0w/FN+DVzYawkOTuldTxI1c3WtzTE1KIF/g7h0vDpLzKoCHLNeDuxT1nKlMpiofABloDcNHTof
JkReTth3bzth0rtd3hnsR4iMz1hx+G0XKcX59Nlo4MK74dib3Jd/lSnQASK8U2O6ITugDBT98F2o
BLCQm9oQVJj1MCTfCyjqhyCDQLeOblCy2B7NrBuVakVxgt9xYRabVTbV8kWzdAxPwUwlmSCEX02s
Ea6EYdCUzj+EfzsQ5r29IeOgrn4jNlvuTcGvQ7cDToHchIT3PiIz/EzbxkVBDGv9lHmYg6sxocgb
a7bhRLyeZ69wE+/IAFsM3WfxVz++c9HPtoI1GcLuRPIPBy4QKSPJUyBE4wMIPUfKoFdoZX2MZqzI
mFgSpima8SssTS9y/yby1GiujUwBLs27XyyhhW0xa+h9nNVzfFjZvZtMPzLkriM9M6tnxsGX+dgy
PDTbZTFlp5D6/3NdFvDvzQ1UJZ8q3+kBHkFk0W2z5TwNxiTm1W1pXyvVmJeOlHGNkbhd/Tuvb5qB
6TknA0iN0B55N1l9IY+QUFAM3ZKEqKmxrhXtPciZwrCv6yGC+WNzgA4FsP7Z3sDT+ltLnuwj8Lcu
TvIg0BEv3f7zW0B8+V8i9UHK2BifMhj4XKJjWCs28N1XFqZievPUtipkvcoqcBCWZpYy7xwmuYVO
ZKUfmjwUzrAf6+mRgwUNPPm+7tYO+fDq+wvlcsbc9bsbe0gTBS1gjuTTMkG+Ffh2ZpuVbG97Zs0g
kgcQEw2+mgkTAow1rcEjj8mhg6aGVRdDtZJydFYxTwumEN2c1dm8VPBDMayVn/pDnWmPH3AyUH0x
ipSHIN/o2sgVr0OotoV1Z/BAY9ocfBTAMx4fI4Q2BF9SDgs3hap4w3S62JBmE67GWS0MLZMDR1Vm
jTeFdr9ZzfbNOiVEfhvZuhCDRUGaPGjfHBPmsycw9U+6NlKiuXJuLiw2cDFHbbk9Dj0k87BpRC1D
mwgDqLNgEGshrhdVecMfpn5n/gAKdPIOngxDaiHC1mUH/G9sexyaDq9Goj3TZcyzlst/mNXX22y9
jbPaBhLKmHXCdxGV9QvGF3Boz1DAIWodh2K5MWgB7PCTk0xZiGCRMTq+PzX9CE0Xu9ycSpy+GRHc
x9vMUjoOQpdVZT9l4JOA7lqWeWD2aNGKeVuGsfZRDx4dWJPZrttVAbZtRT7tB/NdKe1P1eiE0jbm
UW4ugy4reCjuKythHAdJYW2ZQPKr30vhF+w48uG/Sqcg/0PQ9br5W+SxsY6hiPoOW4fu9RLduFyZ
I1uQfyiDe9ylFuR0ZxQV6QpCOOS2eXszn8Lz12ABUUXsWYq80hfu7z7IDqGQf6ySMSTtSoNoma8f
t2BK8LQ/A9heNNI3kf0E51EuuADBJnmObFfwiEVloAf+NUW8gMeQaIZDf2zUOTdyxy5RGqrt82f5
KUCFWlVEzETy6EV27MqR4MRlz8E2jtZQtlxfqEzy0qBn7ErV2VjkKYpGJX1OjlkEGe8EBA5BwgA4
FHrI72rS/56vTjr1rIIHsNNfRJ4MOYHgai8VY2wCu7NOil/q+OTslGiaev+hWPdN/VDWiN/f6/7w
SP5hSiNd1Fil4yhUMZUO1REaVZhXKQTImGzb83V2jMRAxOgibwKLH0ZC+cVyGmCK0JV66Qo5b0rQ
Q64JNKWA1IY3aMPN9Mw591F51bH8AZqlDBdBotqo6VpMilocWLyKa934+50TXR8i7/XodsKdaLDi
pErNTDgOBxRDTZLt4rsmp/m703bVO9h96M5hplQvUJ+AZpJUlE1nIRkZ7m6PEldpquD5UxqLMU0w
6guUnW9fAigHy67hlx0LpKoODV9xAZ8d7Im0v68HAc51I90yOC/PrZ8swbeg2RhHH6IkM0+GSqp6
Ox95AwUD7wZ7ORt7BiFuXqPweq8Zh2rWBSg8XJm8s8pKd42/ztZfP6SB++BkVLqqAc4MxvIUlDQO
SX5Ko50g6hGVHywac90Jb4uDNWzJ4wUT1SY9as77O8G9n2pwKBBjLgJwT7YYdoxmVkoVDiD88iRa
4+X2cOxUptCaUhn7O0oB6Z4ZrSVnBDQFmM50Wr5NvIUPcr+YMV8pJAwneAGru3essm8/34G9s9AJ
zGBC4WJ042sQMTD1+JZ5p7Jad0nU0LSJ3xCG1iief2eDOwYWnQGOg9iI8UlLwJNWkby4lL+JIZ6i
6i36rul2cz6jtopDDB6iervCIEldPtwHnWvvYs5ZwuqZtr8W7Efv93HnCVV22HTrQFGBAgciWmkr
nh6CWNmwc7JGSaY8F+9Qt13uNkYE2lXdkNzGAMdz/a/s6hdYBnPka5HqRybHd4iQQ1OpKKF7DVXn
wzT3JLTGSYal6f9tYM4jx/Tv68fWN8Gjvpd4fKuqk2naL0Kxb70rVPSLfBd+edZFKTZBSZxTMGf6
ludUJj583daZ5E8umpghwguIBFXG6nS1RymEDh3BbrFyuSPhMfaOvdB2uhUuZsu4nGoR8zSVqK2O
Xm2KzJ7Mh3coG0qUejTZFS6pV2STt4HjdIdZ7M9C4zDZLHCAYeqTHHyi1dJ5wT0T9ZztjUABztsk
6d/uXYl8+5wtqfr1uAxdpX0qmkKU2CJEBF5GfziwZn2MeewK1nst9DLhUU+pHS8u/RbIs64/bdEe
MkoFaf3IMX2eCkQKgQazsA6iY+jsuivPdwcbBph5Z7uio2jFnVlTQ37UWUss79Ddfp7PXucHRjsy
ZagDNj7FnqOmjUUxLjEyzpBKcg2ZnQB0Ln7G/dDMLNQlzOObrkfpUp7TtuBkgctjRzW+MNeTtXPU
1jc7xOI6g+/mKvgWEbr+e+0Kw4Ka3r0q5O7dg5F7joKuc7TEBlOCTz8P0UZNcTBIt6I0rvZqhnfK
GqosySxjAVEWs0f1vY8iW0NWZEOU2g2Lzxl2+BzhnPV+4obI7FALvfzGav3qdJs3ZzOt+kIKGPH6
CkddL8/RE51rcypHPanGAwwiFaO6xmNm8q4sYwFXKtN9PY+k5Vcg9Qg2/ZNgIBQ11flMxysolOL9
DJU1B6+mXBSHztapDQ7UmPprt1MqD5f8e19p/J4rtM9kOO6nW7i+4XyNZ0SLsPklwoWptxPkeCi4
DOTzbc6oKrmvJs5+PvKvrF6dbMkeXo+HyYAruyEllJ7CN+n8Zk3eTSgDwCLggqaciCYRmtOcyUC8
QFfq/J43cXpwsnGU5EUzqpeUO2TO4scbhdfF3YfqD5pcmr/Lmjq45dBBAfcx2LmyHcNzM31hhmcH
9yx71ftSRgxfWx2nqnlHZ4BluhYcvzL17g4PlGS2a817FQgyYp3jz7DN4rtwNmuRHmlpa5O/MgUj
AOVEF9ENYwU9/xpDZl5EKuI6jLI0LCJyOJVtb/xOtbwkV/IbnHs6J4qffdfvYpOqu74BBTYNZTtV
UQrCPIfAEbz34Dg89A/aK5LGoaGGdStZRMTMOeEnwOHdCKH6TP1u0aGIcUmlYQVxtUmMqT76FWIQ
cvXlEMaU1E23/wN2jYdHptb3lpq4eeB0f0mzGIvgPgUtcCN1scIAKT4VtEso7xObISz3BcvxUT5u
mIVXeHpFZAv9ByHrPeSVHIaDJgxWu23M6aD6L7K4TOjGVEsAPcpEM2iQrR8pVTA5pH2uDijuqkge
ElUHDr3K3ur9M1fcaaV6kIQdZCKSioWO1CIke5bYq01xScAFH8eQEsETCXcEBVhaoYp0MImpX3ol
Pmd29X/+hR9BmlWQjO2nKwPgf7Fm/rudP/9R+bDLiUdvvwQv/TGc2H6WwsG0pEt7f/LLysCi+BfT
RQkxv06yQ0KNan7ksr/X/PGO11pCsHRaYh3Efmrf26Emu2vccGLYmFWCnzodsFZ2YjfHGkQifbqw
CEVLySN0Cs0IA1hqIhtxhIUNHCIi0sSWYPsegjuO/giRBm8g7GH7AwrWED81zXicSMvk+l1KaKcj
ZBwz7G8yKPk60OqFuZGM1v82S9Nb1OBDZnG+SheiJ9le9BiVmEtuJiC3Rwic88NlpkGL68VDFPIz
StCnHF4nIw9KmQWAUQLc3pnXwfopGr4IeO0qlwGfua5Eidrh5kaPoZinGkTCMnVag4jwMX/jCgzY
Z/TxDm1aAvSijY6nr8TTZzg1XEqKhxQ4FEmoSThdhX6aciy1hHROTOycUmdeU2PeKnGcMI9AJjwY
JF7IdtIPXpHvs0tnLZuyWATpxNkYa5T6xCX5hWyKQ3zcglqvQOc5UL7RHIsgo/wXbUoZ+MvbbsvB
5Kwim8Qm0ndTO3nYHyXnPD0ECDZEdF0dmYGqz+YLhyX80WZdGbtO0rwPtgaIpodVYnH88UcS44n/
gLNuYhCrtgfSQFKrzRD7dHhUIhT36PCtAQ5Q6sBvURNVHsGuqyaE6IEMYOydYKc+ffPZLdXX9niJ
wbz4xQzNsMVsPbHyVLecsCUju17NGFwbH0xU3S5NWiU18sFENwbjGLEM9cqGf3vOriSp/UPZNded
WE13cPF/MHSr21NmK5U8ujEdX0r0qUghINISOG9OM3AHXi57tLEyCIVII6VY1BWRTbWsf/Wcs4t6
o9rRL8xMoKIuZn2uUYMZGS51GeO7Au7/Tc5/ASslPoSwFIbWQb5RoCg0tJyPstQfpXcfrAUebzUA
Faa3YXWX9jOaoEz+TrJH7tcK6URRMSpoGH77JfEx6DEZcAybnlGMMtygm6e138WjUPZ8X64F7AsN
Yk4JilO69Kj8QVmZG9S6HK0fec2cetnh8QxFshpQdFHbS2icmJ5CWCoNXcjA0savNcgQQto4SvLt
EL/EZj/6RTZMBDQkqIy2PaNqNWvCHtM9A1uj8VhKIB+Tau9d8X4T3ilN3t/rdGUAeBE5MZk0w/Vi
PN3PC16gV22Mvw83j/ghCVW3CIzPvyBnFkPLax0WXD7itXxFJlXHZoaP+g5VSXV5vPsCfQ5EsSb/
rsZ8lEQ5s9451WdkRxG52ryrJ0ErF/fYUzzVJCvXVTebd8QNoF/ETFRSc72k4bJycEU8cfyjqPps
dig6CXDDcmB6GrXk9JGmleK7f1WvvnYzRpZrkMk3WS7UP+LMvyfzpTGn/BDYRAXubVmhFwPijFVT
xBh4SeU8aj7jK+9vdIoa8zFJ5YZoWDWQjYhOaO/eIAlHEeuSF+mWaAuV5CNhnBf96e5OAkvAO+J6
oBqqxrTT20EpdCTbW5sBx0Z+f+cvXhuAe/p6eDO2oldwmAHWFhC2I7wBEenwKDh1dhbTX+XxNyUQ
08DEqCH4bbkVPoUKWqUZKU+PpWyxsUEi6Ys4B2bvZXsb9+S4tTXJJq3Y2PM5sWvsCTqv1HLIjRRT
jSVw31rRvYKkFzN96hNkXPsp9pClknceTDWGMNnCDjSUABmm1DSBMKXqHM42TrUULOWhAW2TfYJd
Md1IU8smIbRMAgIzsKnjFyfYfFY6xtvYId/e3uBebwf6zcTjCI+6Swstf1wu5Wyj73UeqJ9wgro8
e8TiJsSUqmSxgIkrf2haqLrwDfey1uCZm5774uCbLfNWOvRqMdPiPBmJuvEvBtoqazbETMoobVYg
woJiszEMt5IdfmzXEXOFxuHMs77Zqtz8PylR5jCfhMisUbxk7eS+4OkU130SDjWMJ/nJyVmIMVRP
SE4mOmzYivM6hwtNtJ9Yo6xC6neEMSazfmMFX1xKyTm39/B0XE9hcXduJMrnjA3BS4c5o291L9lp
tLE0K2zilk31iqW/Ypd7UqkIy+YSpCJvUZQzaUq+mek5BbKpP9vEG72oRjEN8UMCnevKTO9w+c5f
nBh6SB9oRxjG452lvqLvg5xa/+dP+s0HSP1auyQmj9erxN61WMBxzIchZdMMM50hfR7m7E7v0Y6I
OsJ80ytLtFU3hsxiJiMrFVuOquBQ3YSUwAj5uNuD5oV9OWed6AeF+jtrWjVOyWMUjFPCNtCa+Umq
35nbbLSrKzDtZqrW3YwuMPTsjZMHMJtwHg1JXqoKtmsOXd15OrHbsqXglzt7Zkjbcl7DD+pCvkD/
2O108d9n47ZBUvaPUyLrWT72Q2Eji7WwZ5GPoUv9Jj0ZdBMv8y8nyd1/RzvkSL6Nqdk1ETt+sP1N
rIyQce+qncV3lrwZH6tywoBnH4A55A8dqrf6Q/OhJRH+fEvIM311BZwKjL7apbUGzYe+0NGDPpdo
E4ar1861XOlqa3kc674PCwszvN11UhzBCoOOzl6gXKmvfwpmWYLsHkVGuCM4O4xtGuxS3HkBjKok
BD1TVdF5QQOXoBHXWpujB5G5hnNaALBRhtMXCYtQNYuduLrmwQK2JUCD7lFQL3Q7otbl+TUX3+rO
DhAi7N/kvkxav805iVwBJzlCSHdNWQ779FTPmwFzexq4Xw6cz3G4iVL68i/oQy6i3gqoHXqvBFmO
AeM7FeW+qYxbDXtBDQxYSatC2Sfl0EdOL8pduaLQ1zWlQe7oSJaMardGlPX/WCRq76sZCzw5ohuy
JFxV1z7K3+yRiYFAwoq2ZYCO7y2Rgq00uts8pAJLLUaSHgkzvlqGcZETeuuUKhBFZCcxQ443qC9D
1Llc4+2ESQULBeQ3/FD13JAQFYJybY3CfYmbvRzZgfUHyhykUJp+Q+YhUpblg8wbyOZoQS7ex4oF
mtdPYrQMRlq/OKHzqQz9LzMYk7qwFo+LcU+1JjbvfkcutgZqBQ3SiGTXpnrCqTlqKyTsPnZ3RcTO
I4+L1EYDmLE4oIQeDiVWJrLbUqNKIp1boZyd7edWDeYDBLpe+oIfFq7+Tv4KcRZJEtOvLbOH8uYQ
oKglwY6EyW4qp8HVecajyYM+OyE9gRgasYYfkQw9BNy9dz0cBu1sdrumta0lozDHg/YiRRhczG7p
GbQTe2fGvYBsr77kzSqxEldi08iQ3cWvTG2WYM/pj3mEy3GgJVfjWNXNAqTnH+zhlTMLmySFAq84
0d8jbRU9a27BbDHD+Ez4dyKT2d6BLIoQZUblwnUljvNUH1MSv1iGMl5sUQnkx6L+vahRpxlCJoUx
zO0qm0Pn3XhmspBDIC/ZE5lUnv5wnvaoTyyrnAU7z6RHMA9ifhZ4S/l+XWbj0U/q3gkX+2hKXlWC
bLK/D+SUZ971+UblMDJ5DyryeAF8WQY8QBKPeoHUp0h9ISp2/HlyaRu7KpqjFLIuZcrz+Ck8mBBD
qL0Dc/G+Z3U4EgRz+vJPQ1mvzMJupz1EqeZsvUiwnSrrDuwRlAqxMaxqpx1sUMYmeMeq1Rpf5Xlx
U6yMs/ldd0uQ8bsLsHwXaQun3I1TCvVA6i5vCnA7WXNjor2rjfH3WApmQvbdntwPa3INkkU445hh
mBvLKCAAok/2aOBwf6h0xzz5T7EqjHjnhzOVS2G5jYI01F2T7yfDvJdy4tX/rbl9q7ze2ksTJH3Q
5o8lj68o++N295oRI6sgmcMpHn/DOL1Mus0+vpDRTzI24N3+jLacJ4zPKLKMdGpGEaSJYxhYUEOs
OAPcdnGGweB+SUuj6vu4gs7F+YtdBtaOW7zzlq+Rz0oqVzreZoDKIPIMsjzOnyUAkQKddEPDFeZx
C+2BVaRM8Z8wDrzLZe+BrYu0oCFFRfJq/vm9hY6kQ7VZJZlz1BWA4GBjy17pGzVbkO6alh5zEQEu
iNDO49ej+LrOrBF5bY3rKrTRBoPc1DULE+ZclOuHVOhiND1EtvY/VuH3AYvPuSclKU7DkIYrDFr7
poT92g3fk6EpS19X6VA1E0PWJsxNbrXuBeF4WeCrIWd29+sb2eBwNHWqvjXShDaBSjeP2qw9A3AD
mV0VfVUkuvIb3L5bAOPYxglhO2Bn0a6KqDYCuYjE+ryc6GTgmBIrXaLQeByvLLh8DelwHfqLbpLy
kOaZivLFTK1HTphgblILiAArKQUraiSqwsnkA1Aw9lMfyInRUG3KTAhuAhzcL5N+7TLrgPT0Kary
v8LehcmuQ4xX0xPAnqoelKckNPX0QM2d+FUqLrwkYvMyarXFawwa6zNwKP9We3BD0GpTkk8jVAgX
osGAVPxYoD7vpVgA91nfTTZgc0hY/3IKRn8P7YpgYiXnLV4YK9gCgzdkSRwoihYqmqC4iarvfYKV
lWR6WmesX5JfNkwkoFOgIEwGpuc5Xl1fHRFcEayO/dlgJpIkVlunG26nG9GvTtXh1j8cazmQFyok
Cl4h6A1HB75BBeDvjOti8iEQvsjxTY+AOsin1iSswqqVP3rgJbN6MT5gEB6VGvo0ZE1lqBTDZQUT
GFSEgIXTky7cvuegxUhSMWTj9G7I3CmbfBJMxeDkd35qcU+hgFocWC+CDwm06uWVRs9xqPZ8eXi2
OynzNNUJJirdzPQics72esRqw/44qodpTAYot6EmqUBoPo34RrQaDrhO9fhRF+dYSOKHeLtrZAUu
Dfc+oY1otWI/UkjDb4jD3xnBqMkazxabZm99gNeXPtcbpRx/202L7fN5ab/VNhEqZTJX2MQvICxn
w+AuljnahOHX3Kph2/BIfxrb3ppTazWCaHgpFuNJBEM4+sunMzKs+vrtssbPshKrmu0S/kUU+ycp
LDBvYhQ5aDxtuz/JPJYbRL8reBB0Tx0i4LdFn7DV/lFuo5nQgzDCtHLd+Rk4F9sdD/dV9riZOsn0
dieJScTKARObLUCn1lBygDxO5M45bMAn6O8h6TptxCRhDcuZVgUNkw3UtLF8yS+DkB/FrsT6tnd4
BzclCpr7JQy5XUNAoVZSUu0wnrYOC9WXmBlSrbWIPNHUxc+cVofcuJXZbSKr/I7me6kHbQ0Rbihk
q3TLElFMhIf8xXo6naek8dlcq+kaSNMJrKOHKmBlNrHbN8uJinmjR08zTpH+XCPkWBGArHpaOQAI
O4xaE8/gvw2woGGvj8AAX+choxsfVHI4+jtNWn96nuBI1ONA34K4PQhSW7qMvuO+C7Opc2owARFd
gOIuaiBIYwT5DjcZFJmF5Z8RQRw1zRfKBhg/Jn1SXFG3Xzg2nVxOvfTHVfr/O/MutbTP+sNYod00
+pFe0gkkTIlWrxLgRv3imnDdRhQ6EVTQxJO6URSVFSRzrFZ9lpC1t5jRMX8+Two89hjBJ/G4u+MB
Q52wcZKWATMBmQeQP4kfoGrwkvgZDKQ0pIYhjCBSCyyz4yJZkatLZSRpY+FcJY4I6ezqcO9Ytt1T
6lqcwtUg5MCsN+ZWDCN0iT3+N1wSuPS5YgEO4rSVzLyYhr3wIPRfqZ2vXNYBLDpyAZ+MDbvCtNO5
YNVcXGogMzDvBw/VqEQlippp2EahqNc9yv+mFDGLSi3z2ecpjStmdwPbDCdBHW84eQRG0khPV+eG
16jDKJ0H9PqjOVf+6tUJ8fPPGeFpQd1Yf3o2kq/gul0BK8E6ODQnLK+5qDsrVX/n2eKnJ539PXI0
qCuUzWmC8zxumh9deIqI7e+mtBhjBYSCZpDKmqwQbqocTFx68BNi9QHp4E2koFZFbBroKfqGsqql
qsukGIfUEoLS9ip6DLnT2yR+nfrQbTSyiBY66FSy7C5yCqlR81Pbc/HF7/K1Tqlao6uyyjLmqW0A
lBARBYZkId7GhS5Q+pEWe35tRZKvUKccdUFevDEBlUxtfxcGiwW4fxuuwvczQMc9ePNOdDvgWcDs
rhQQ0qrwbJw0b2dtjzoZzaoH/9nYO079YvwQx9fLfPS5sDShp3qzXxbbjUFTsIv7txNL3o3DqXy7
MZlP9Tx0i5ALgUw2UrnvWeDdE/x1A0zVJH7UtTnCHNc+S0GkZbbzhoDRsdv5GjjlmViwc+vydc6m
xYKTvdBR8PA5kUjjYRNpeyZBt52QJlKQzfC4NFEFARE5ozfC4eZDg7sQGH0v2xyZ2JQFN4GaqU78
1/q7RSSuTVp1Y3vS2AKP6zIbA+LaFRDc42WtiET0le0qN/fVuPtAZJMZTCxmv/ossuhUyJS4xtdK
vVlyquWm2wEdC105GC94VoCGZnrJ+X5bPqRUpXemCJmRUKwIeN8UoqSRyeS/9ngUIbRsDJ9iZiEW
QnArNgoAHzhzWXcdLmq/oDmiYch3VzqKyRUUMSHe4XJOQwe2XPKyg7QNSAGh0SEcsdNtQBUVZD4C
YTmKoIq1zK21tNh+4cS2Xcn0CAdYJIsJ0fTP8dU2Co4lnfA7zfqkrh/7cRgUwMBUwiXC9clfxAdB
UYKHE+b/+qdcKFMin7GHNsvv329jVGvNXGvu4PNR4wf8LHvOXuW+MicqXLR50eCF+pKppLP3fxTs
xdONLlzpVotV5fHEx2yIfXoOFEErdufgqmZwoO5uluYb3u6ZhsfNIC8l/kNHmxtD8wzWnCuoOwYW
PKQPuDY29wy9YPnFfW6ZRgV/sXacn5BxaMrWhZGgLKBgYw+B+FyzwP5NBtqrXj0miND0m2VehXjf
o9quj8/p+xCoCyLHJDcARL3RErDe+1jndv75dWOnrFFOnLE3dllHzTI/ZeyxV8lQbqyTJSlxyKRa
h0b4jI4CRcF0ciGhr67tqKMP8SO1yrQx+6YBUbBBsK/e79xm9HRiLneso5ijeAbaGPr94lTbWHS0
LTDTEv+M+615pkTngVCHUhBUTSuNLT62gyo8N48/rM+dk17/ffk5DOcMv35/wXJCLaXEkkBDkUou
OPdoiQ2RgvPn+8Z69fiKJ0w54mFerj/ACYb0UZgINnGS3OkslkJChFrK5N0G//znTP5MUY0xE6eD
eV76/VvhyjaXu2uL6BdfJ8eMj/XyNs71Lja9bOzP6etFDLYpigLj/KR1qJHaQkagkmkNYTO3S4Ev
0UhkL3/uyaqrbmypME0+SmQgMPEZUhO/rM6ysZI/EP1NY3ERLwMZjukf5MNs8KJacQkELio6KIyc
4py7YVAvqYBPNyGoJ1ti7d9N0sZ4mlX+3BYept0RVn2Uof6PsKCnnHnR9U3nS2udkHieNUeQAJIX
MWVpL3xKNcTAHuSXDgNQqm6EKdbkusGShkDMblvNwbtFnbe8M8mcyC/pmQoBJu543h6rDTGoF2B+
I1SuUq2CBQlDFm6soWgVLWOczBcvb8s4YBjmcOQGcZFKjK0vaS9Q/C+rru+CyIPpC3PuSX/6fm7L
O+HxzqHojzwou6mPWrQSyvY6MaChlhINhNqIypAB3RjNKuIlrA4y6K4Azyr3Xcd5YYYgNBHy66WH
eCBNp4XM1ViX3CtP8PYpArSN9/hr1i4rD9Sc+tGysReUpWF4s/269IMcJoczZ4RDheNtYH221cAr
tBN+KoxCSAVqT8VcWtWIQvMQOIdZ5oDgNrrX35yrurhOJlgrwzJkfnfuzqTAa/nPLF63qGDD30h7
83WgyfEjzFgtgIJsSa8Xu50kkvuI/6VP2UxqrcglXPxoBTNSh3WXAsOJfj+TslfI0jJ0mUuV48Pp
a137ZJNqaeoinnMbi6c0k49ObRF0qynai9onRnOGMHqJ4cpTU7G1Eec46AcQ5nZ9Z617U/EHuniW
rXMH8Cwmh+iJXv67kpB78BodWAhZ504TEBpAnKln7dFmz3jagU+QSMiAlY6gf42Trxtpb1lYYCuK
qsfFvi8UrpSbSz80bjjowsU0L7Kv7U5zq0nSfiJR5Stg0SX2qbVpfORQxm1kJnepZDXADKI9Eo0R
xehVgO3ePYZYPQ/hMJXpDUvushSBJ15suvCBxxKwarOqY30DvbT0ueTM1P5C980D951Gi453Jc2o
qlHdkRD6EzVVMICnFHtwzRjC35kuau8rWv/BNYQ2uiUlN96AMDGZJDDEl7WkekcgZ/sr7Ol2xyCv
jW4F5PL8CXT/9mjKEB1wPbBPy45cKWsR6AoRc9gR+Mgv0UQNFh2egaBZdfIAQDyt4rRWcmR2U0Y7
8C/lg+0Rxe+StL0Fc7EOhVUprE6cyPgc1y6v7ksDSdqflMSkcm7kO1cwa1eHSQVOtKPzfKiXaSuO
BU84o181gTfxye90uXiLUdWs4tEEKOfnt1M3ZRxN+2q2G/lX8OKR0Xi8Bg5LKW927eYF2Hgi/dVB
CIOlylHy1VIg2tipRQ50oFWt9yK3Ba1RPpmyi5Foa0TcvWKGHgbLu8+nkNcyJ7HjCGmoGI79MgzP
bWrWPJfkt0xXkr2CUia7v6zGhH5ZeNfDIiL8LnLIt5QaWA9yE64Gxf7gixvN2SXaS8K99X8A/zFu
FFZEShM37o79+UmfyD03/yrpqTRbP01VlzSkNOjjv0Kaec14bsqfyzFCh9zNWwJckpk5xNXFs4mS
cU7fv0uuG8CkEe2nt7rXeqvk+0SviCyOt1a4MadIyFyAa/qoanJ7Nl5vIiZcVnuhEnyqALfD04dz
pOHOzq5I3nHEGTn4nNIZ1sO2+fnK0pNhiMVHh+fywK6YFnBWfr2cbvW6jCc+K+nurlsDSuihXftx
FBAkLf7eFIcHKW6uLVNBOl6aZxpu5LO6W1hdJX9Xi3l+SosSebv0yzWdAhrItMZ/tRiPvblOTXCs
5vs5kNVvSyFaKjuNwMgVMKGJ9vntZ0+eTQwVBIVnHrNGXZQCaKl9Ek0aIylB+wmgZK6z2X5rzJXh
x4DIjQR0F6M3+q6uObaQbeTQsqioT+XRSxts0L7CI7sj6PYooLdl85+dSyFHXeapO1MToSAQ47nO
/CL68mHGdeXahIwgBNMR8u9xLfBq8H9NPSu3tm8t0J1XhZ8mfbR/Ra3OK7fT5XI6toqbca0wZyXq
/iNFfprhiNAJP6Yz7lwNnLvAxllrpgso3pSacercfRgYVnkg38NrV/0JXjvGnbJBcrMl6qs1kB7I
/AVhpKG93h+HFUjtoApr44i4VstvVKVy5yOO4WbcqgW3QtNFay6Nja9JLT/8pRRRCezwmVTUOlmH
sCAHc3rTL1GEiNRCHVTaTqk3drWVd5BPOFzzuamlzZaXBnhIzx+MBf1T+IXcGfqiSxZDNSHcxTfp
oA9LhY97vr/FyFPajlJ1LfaureTM0+X1oB+joKsZ6D29bvt+DEfA7uI+IJLiLqvFBvPCcmkoXZen
1YvG3XH+El/AH+P6N8VhrONImygy2hRMgJ8G424z2a43lTmv4S88WvWkGEtsJVUQDUc0+i5VWsZK
AgJzFARCsK23qXgN27OXMoDHcEKakQDURIGrI5/U6L+Jz/ZV6LB2DGCZeoYvJiRf7bSFFbUI+PFF
+WEfNJ+I+27bnebLki+aRg68Tbpxa9XD27Rl0x/dgMYPQP2g2Fj+aDSaal/2+BQA9ylGtQW+K23A
xHpL/gPTRLCEGrahoIXEkhRXGW38Vhw3+EJVs6NPnOwFS//15TKd/XBInhg727G3Jmxk2EIgubUV
i5scjySzigvIc6dt+Dv6d2t1Pk41gACY+zv3uXOXCW/5y5OZACD8sKMPjR72o8VXCnltsz5NdDOM
1Zi0y7B6I0yjYsPE3T0xEzQzH6WmL8+rSk3krh8c2ctzcG6SdAnAjzDRZ4xXGp/fIe99YD2G/b5w
iOzY2wMVG24HJIadEld5BLOV0fmeipjWL3L4U3/9rrnluifsRJYu613p1TOVg2gBjB4/ByqOkHds
OygPFM7f8ijTyjYE/QbfC41eKrKBuObeNIYMykJLBUQASc47kQTDwNo/mPWFJpbHt/u6DUWzy51a
454G9aUzDYFP7JTHDAkxTsBmzNtYAMoaG2/dlrfe3wIqukBJiAO4MMnkDnba565j0oKPUK/5iD6I
M9MQzZqNLsf/hfNIKE8NHIbs8A0Q7eo8TyLC/t8Q7kXGspIuLQc29ab2tEk9GCO0gw4fTHwddkKZ
1UhU5fLeA08i3vFIA4JTDV3s5MZKymxBCl1dB+qmdt7k0DH3oAcL+1UaGakykHOK5LzOqai8J4JT
pztuZ4nMQWE8tzI5O9nn6neb+wbeoWOPC88mIqjWMmRyh9jK4U63Sm0AyUI32yjM6VrWrKOC8iny
xxYPJN0Nnj9zTPfPlg3vPQbhShk7DKoQ8TakBcyz7nlGbRjVrbHJlMDng75lAmtjI+XZitZToRNS
ghfPFOxD1UrAr0Kqj6SymZ0Mf4By6llh04TbvKDG9uTi9C5R/ZdjrMvD0//ePCuCHcxhoObIVs0M
kKQPQQmoUSF3jhaBOSGhcBewZYOnGfc6DprahqMHZiQdmy3NzhBnYLcfFKtxUOPMbsPwXv5JIVgE
SawVxz0hYHsIoThyXPXTP9m0qpDf3tigVFNMK6hI+tZI7eBIn/psRXHnYHRxXnvJgkNcK2NvEglR
hvFG0jGfnuryNMuQCHgkK15rLjMj8km9C8j6bmojxvr/5Ldt0JuISc/SwhcoqqxZf1N1E9TOz16+
QOyl++x/Ib0zXNGzdXzoSlqkU1rXydcMahS4turNFjhX/UWUtEH9+TQd/Gso9MEj1sISl/mkOnim
8Qkv1W7tTvqocNTJuZZx5NcA5aS63N4Qsy7CGEvk9bGPwCq1MGAY91NkfA8PX29QGszjx8xALdDw
siyA6K2PDJRMUT0T1niOdgLjNmddjKCkwptF9+oCSR6X/mLyNKKJEs7yVPztyypeh74DZe3xw8PG
vwjkIucyebRhMM/anw/rvMts2UN+weSmaXJwRSbCB+7HBFhgvIC9oCsApq2Xnj6HGXtZ7B0wrSth
3hEoPTCDuPwR2QeJasoW9XDkarkv1YWE82meinzlK/uagMb8d33vGy/xPUm28s8qBQm4yrWGAanL
V4KmiUqtm0S2SmIKvg10w2Lc96dqzD+qLsR/xzlmJ1Ajre5spivRj0Vtus3Y3ewGTJcAo8aRJ/ZO
jvpq/ZfZG+WKCVOHP6ww7MBX6Gt7xiiIstmubx65yi0+3+qjKbtc494Lz0t+OvNrp2KJIEuDpXTT
Up0IsLapNo2Hiho7o0XmLnch3NKg0eXmm59hNbryLokfocYeNxpcNv0dRENztryKbf72hizrBRzq
g1ReQy3pbcyzFuq+iGXg5j2MTmpP2YKt/6btdJAfnL+TW7Oe7qKOA5QF9MPXsEYBM+Rt0D/V/KCk
dSjcFvnaZFBeM7WUjiESt5uAdnoIzoBU3JfcDDC3OoLUlxoI+KHwYpleOsndULwxbn9cfF3WcRER
apsGLbYpC3ccKkkDfc230xwrt1KoAWNz+LDzYDo35SnSIzrIHkaO6lmiXODEP46BoGz20O74iVLE
VMzLLju0V6M3NzEiHOhfGtkVcOGFzZ/JV9BUhM6RI/qANv7BxauuCbyPYEoPUlM83QG1Sm3tIDnk
MWROrRb1CEVL5E+FeOLHOBVeLV929n+7oW3bWBsxT6jAyBv9ACoXN3nDWupITWzZ9XNP9xZkRP2q
rD9L3LGqVCBAD3QneC1Es6Kglvfv49wIAuWbBSJJ1SR17SukQ0xzeVGGsZ1+uosB/2k4oMmyIWMv
pWbfe8/wZyKFRf0AtZcgC1rrtvK4ZuHykQEIG4d6/WhXipaUGldkzCV9n/ehKMiUWvRl4KsLhmKd
fWt2KhdF0TUMYZNU0ytR3/Wr2xuxFA0c1LsdRXQhaQKkv1Qb55bJ2d/LnIwW+ly7CcChLuur/Wuv
Gp3gAgACnlXeF1nCXemzCk8OiV7RDLzvoTZLOJlm2UJaksJ2reDrVgV2YaCDtTCXgxjcvy44iY0f
cI0ekDjS7NEo9Dp7I7R9AjfMBn7Ztr6UTiRpTsWdAaDBxnd54m4Z3vNeZykSoGvv0tuXnCno36hU
3Jmv5CA2YIZXYgu9HFmjkAlJbPO4Dv8igzn5QyZ/aI5Qiaqxqck0zPidC/36VbXwCePMoW3y4HEr
Y3HmMabgnpJ8cY5wMNr36ltNdojfZ8IOKVoUddAShKE9DLGVTXmpwg9UKeb2mpR8Twedc1u4u5rd
tlyWIFKQLWI3x+/Rr8IWy3p7lAK0Y7vm6e7pzTCYwr7cIkN1eM4AioF7eQ90XD0tFx/YLUiaOVrj
07oQsW/QVKfp56M7Irvt4IsNNMjEy3GifUrzGNa6ubgHFccSKWrHx3LzLefmAB13TJ1F50zObDvO
6Ntby9zh2ziivSjOJ6QYHdDPSMUJ7CtdZsLvtkuZ3Sr3garWA9Jdff2ecmgD7EhyfJvKH/aZYBRX
1Mt44OMwmCqW2viNkH15riaABEKgnciZGfyJPAbx5O6ptKhM8EZraNTWO5gV/XqqYxSfg1hX4Sv6
+ZptagsEUVTIlaCs3kKB4w7b5DG3gapnQ5TjJNgHauXJ08HzfKX3VmJqNYEGj/LeK3SVRCulvHld
zxi+niTyAI1bwfqbit0T9sBsd//r1cdbdyCurMRmO6y45jzAdId+PUpnbtM+D1+Exfw+ZJmgcHs/
JE1xPFyuUTpvf5ya0v+RSuBiP5Rim6Mavsmh0O4CoVAQR8H8HPkXb/hr5RY4kN6/MsqQaXT09ylX
DZxctDIn+NQSudDnVXA7qhZKuE5xsmvbfstWcnPLCMBqtN7PwSaA6chWyZx0jWfk31vxPH8el6HB
08fX1wmxruuXQz1y3yOM8BKuRceAmLk4G8plwgk75uTb93lYorHhBWCEQ0qt4ozYZ5yAqW1hdnf8
hLs4ib3p/aKOV8kvAiHuc4GKL3sOTE56YeBEDVw3lmrPX2VMy4ON/hQWZmiCoOSkTugw7ONynM8U
VDaMovfcZnxWLFq90pSJeevZijaS4xXN2g5uiTBbvzVyv+4Ek4P7aO1H/hD6xZOa1PKldJOQQIfV
nimj49BhEnpytk+2bPuDoTZwNQm2fojavM7f+D+fCymCaeswiWvrXUDcjHJSV5cY5CcgquEYmiG1
qzvS23H5VUCj/Ep+Aozh2gzwtKV6cTdOk1waVll+tjcO/B3cG0W9vsfbl51D2N1bA3w+8XWxMBvT
rQk29VIOw8gvqVpW6ifiFQwl1JlR2RplXuNiPvXp94SDNE2jk4YlN5nug8I797t/OhPcufMzfzn3
n1u1Qi0rg7ct1yxhi4EVX169hwz5+dtYhhX89kKhn0eKoXztRHQWFwMbKb6PDHXjQ8tDWRLvqGXJ
9JkRD0qc0nwCbzwXKYjt4wHWlf3RlhDXnS2JskhYr/hdWqAsD+1ihtzwNnWTtrFYn7JMf6fUJFP/
VPwcJ3NBG31WhuFD/CXuC/ebfQtQKpIrcU5jXfcXnod7v+DeLBdmy1gypQ9nolg7GNdKM9nUW66m
mFbexilDneulhCgFAAWHSeCZjpnRgZ6O7ZLbEozT3VKbpb5MjhoWLvNqnhvV2PnoaLGLZH22QdYY
92kj2j/mSKkB2Gi+2bjfnFC1b4Z4g4lzjpo4FyshsN19XHdLEDvAuRhICPlexAC0YgZiObyqz4Mb
4G7wrmdRznxahSjnVidS3UO/kvMKho5jkImxknIiN7cMSNmc3b+bitZiBXar5Kaa4DOtdPlqtyxc
ggujhKMgxAs4oSTOF8VAEgXtm0eaJIOjlkyxgPR7EdMHEIlkApajQlT9tRg8kEalidklkmhGkmHR
RhA7PZZtX/3681gYqOwyI13hn1Q/cFP6cygo2e0DYGfqOWJSzFC+Tjqivna/N/YsL74F3Ws2uFTy
E5rJnGcUGDAJqBUkdrz0LRqT1zfDqS43xMyYI9wAoSQS87in1k7tnIPKe1SvWc5DC6G/ocXBWJ+s
9Ov7dbB3QYNl2fcqUSEsA0NfHctOwz705Xvn0+W4rSUEqI6B185UKm1HYgNdHgkVCT0KL9Fbwg4X
GGi0N6g5sqrK2Wl51qXyJErlpjbKfALgcuXJStAYO4Kxw+HAN92lzdHUhxSvwDXi2IEBuYI52xwP
+h90WAGe6sRX4QpBYXd2SIqLx4akTyIEV0p3M8qkMdpz2uSwuU08GlRsT4oFBreihMvYCBhACiXh
NzcurXpf/KZmTRSAw8SdDEhuJUp6TWdddwl0CL2heRQnVmSWhtBJXoxs1CidOPlnECV3m3DgumOH
Y/rNIRmJi+UU3GQ1KlyX//f/h8oSZCdDBmww5P0qcwqFiM/LkKhBdGqEjDxkO6VnzNt5DbW5LTEb
hdS3S0gGRT17C9Lyfg40rd6bqr6hj+UvccKTZsYE/xRZkEeKgsK9j7kDD69s+iN1dBxrTpi4c4Ba
rhRfJ8iGXkKuDTx5bJRylDRKZ15eJx6y0gJFRkS+o8iGq7TnYFAUtRXk9j9CBhZkifSKxlRnkL6B
Qi5NqVzgIWxnvipdk0BdCM5tGuy3Hf/8UUVl8+ON8rDFrqoe1ja9R5YIM6he6ZtWAQNPuq9C6hx/
+DDl8dtEqyVltlvaX81185uryDLxZi0oY1UwjWZqGieDgsJuvplX0aTCGNjLrf0Wyll0YOp821Sn
exAkaOMngrX/nUEkabIHnNudPfwMerJ4w8RLCVlk4LaVpMFwzuDfHam4ZAqXOLp2kI/vgd4DF6v6
l6cMbhvE39WPGJI7274kBZX9d7BswNYjGcMUQB7NpJWR2iOWxIPDkO4KxUVD7qYT1xr+h8Scrvhd
hiDeeMWu5PlmEv2ltkYIDnDBZkSTx/GR2EQVzv8e9XvZn9cvgXRo6gxiaUMNTtLUFSAwpFAy5VF/
SUiiGdSsJHRf/C25dcKGZredxyK4S9SuGvIVARLLobasdiQVGFmVX3n2MqGMEpCqumsp+ajkeSGg
1zbKPUeY3alyxQNNphTaIxaTCVjlhr+oFZd15msipbOfG3wM+lVSn4cIDVUyq1Gm6A2Ru1sOuLFc
Uv0R8CXeI16Kb0kh/X9yD72mCPj14Gp4FgVe7k4lZ9cebUSFiHWZu9CJhY30VaLoWH6cPjqtdZSM
O+H2CO85hyeCmzXn+GdsTt79xPDQi+veMAc17bCSQ1ppbgf/khLzIkZA2NCRMllW94vRUp3w/z90
WXk99g1/mbhDk5A09glWkLS9PiYv4S+2Cgu9RtBeM2giEl0c/dcLRrWXRS9vFc2TJFI9icEbyYBS
0b3uQsYYPvax/79g5pmqb2mtxq/CEfhlge1J2RlJimS8jFXgeZCEG7orHFothY4rxZdJ9LB8iA3p
20srQV9MPwmYRKpa5I/aD0c1XGpVNKxiBTCcKG3AO8ZphkL0gCgPcOEQBi1mct4y+jDIn+aokwyG
lCNRSlzdPn1Fp6W5ypcAKQRmHYsFNBnFjegwPqeYcGovcn0zi67PByGVNkOSmDrybmXyiOzT9oBX
8XUpj2kqf+5LWN6J4pQ3ULLYGwgO/xi5nqP0opZo0krk7SNFTD1lbshMBd26+xV6lpo3ps870Gtq
FG+KWU/oFdhD7w8dT0W9dLMRZZjvjF8a47x/x0DTXaobrxKaoi47fLYT4PMeUxoFlL8Jzrh+sSsF
liJGzYvlfBWfJL2k/OXAqpv0Jhc1UBklTzZuML5tCNnD7NbzOdPxrb3tMypo3t1S8YRF5Y1Vg5eE
+14h7/fPHN9gt+wd7Gnsl2aD3L7UIfJim80yxAH7Dm7f124/jiwaevYIr4tHrAtihwBPttIX4SBT
8OC5H2NDWZ+owCdy1mOuI1emP2TuNeQ1i2AJ7oQPZ5Lk4QMRQ78hjAzcwOQIOc4rTnN8G4jVqBh0
5cKTbVtjqQjjWopKIZ+9hSk6lECRYyDzyFdQlirxDsOjpWF5cXRwIHtN+ngNzVWV6299+l9RR47z
iI4Eqxv8Aqb6vv1t9ebkWZiJsYcS7UYsDwAUSO13Z0mieNj8D7Rx8kUKez7R3TvR1tT5fws6IvbY
vzcku3uzZMlUSBdRb55ZwnkhDB7mOC6ej5GwfPcRs4jl0+l1JcHRdqydPC/mQYCMrIxWHC7baO2P
cIEFJ6Mpp9K8eKp9mcUlrQPye7wO1pCUYqNV3JjcqSqIvbuMgSpRDX6r34iYKYiHVsHTN8mgg9Pw
J337opGyZHlOTE2oaZ4PHoK2u8ZvIHl1eJJNk7lj9MEV/akai0wHwjvIqE21Jj/av1A1EgCVP9Zc
eeYEBuHjodeQzOSN6SR8ZgMAb1i7KK9Mj/o6espVVPkREwVpyhEaq6+dd6S6LdNoCibeYqE7OjlO
1HmaHTFcjP9z7KLOHU+mfKxCI7SYsyvCJ54HepQc5MNoL1lsbR/xj/o6c0MVFQIpgA4e6lBT0DiZ
yPRL1WbAaRn6WhzdMTV5qEoFxacEzwt3Mc5Q+bu1WzqWuDfuG/QuN0txn1M7CufcxV1qnZyf9dvE
+LRa5y1jTUhhla5LFCuuiSJO31U2mmzCyTlp/Tx/7/gR/4SukHab6hFzv/VY9h8M+5rimvpxYEia
zwBxapTii+/57DA3f2gwumgQxHT4Iphtb0ooSpSemGKqJ43CIsOaPFN2zh1A2htLW/SaTcWOeYgv
wT+mCMzvZiEr60plIwKzsCrWvYtpHIh3nCClhIvT4P54u3ExD65F9UnTkJrvWvGkGopiO9YwppKl
0a+ySGFnx9edv+uWjdzfBC2xaWTw0BmrjVo4gFIRwLcHeqBdvinFnSZi5WvhZxCkAcWEvgDva2u7
NNTzY4waDlB3IgsA9b9OoPV2ECDII6Q/60bOqlYLw6fbtqqF2e2ePcmJr2aT/FeBrioKlNIEEcUR
vevI3kYojI4hs0iC1PpHGQAxuPrPrYSbCpUyEYyY65LeyDFGJqaRodorJ93IlBtMnjA7EUeJpXiH
DRNeWa75eCCowz4UUDEWUZVN74WTUsjxvR5RLoN+K9SgUbHFJjRsqsXqPN9lRcxBpuJcACW0yeOo
sudDbfghMX7RHSQrTOkgAEKoZbS3upvmMnDqucqDUiqdO4/nle1hVpmIOubYhFORSljN2+APT8IX
8mRAAy2lyq7re83SK4ujPEVtQ14bMW+LNjgf6qyiNhhHFfq4yYKr7nRLsGOxsq9NWXfXFu+CEg9J
XEcri1TpePhbFaVJyvfFLlJKC9668sADMMFvhiMKz/baiTDeJ8k6EMrJZLaaDH6e0V/u5ZlYdvJH
+VxUSti/eqqsta3Z8km/c1pWRQfxt0M8h11eLxjsZdhu+HGnIqT55s00mW+CsbbHmldg1znh1P/o
Mdf5RwW9WOqzVcPGIf/IehhCTByVPQCgEVnWJ+pCGQljlCTM06wJIZO9zI0vHYjgPvsIB/LA9uQQ
XL40NVRQu+TI/gbvNNHKQMXLI3QXbwSQ1fLZhtAaOApyfXfx2YcvMYLFdc3URmj9HVeZr1D52zQG
TbcNJfiefBhIBkSyKTsu1EmkKaPYW1dSI1Cek7pevlv032gx8/awgafYG5w0XQELTJihrbhGmh5y
WHhjDkJJOToTBKuzsisAJKGHYtn7cyX58AMqRj2nogDBE4Nw1ICX/1W3txYlKhOdcIh9PHF1zqjM
o3SVI9I4KIyYL95fMyZwogI8Bd7AW0zSfOiI42+w1/SvyQcY4LOLZ2b6roM3SDUrDk63n4B4XPux
LGYdxZs7GCd9KSrcU7cf6a6xlii0SqKjly2Q1HBj246JmopQfMkHMJetQKINkraQy/lHsfoGqRff
VlRQq0M4+jcvSPBtlPKJ5u6rskPt5LfvqtIRgb35It33BYV+bAz0yv9MjSRwBUCrZwbhXmVK8zIG
lXAFmBHPRhl9+94wknLGhJvT65R3B803d2iBX8B92JEV5zTASw2ukYo+ahp4uxVVyjQlqdcWl/PJ
IMNaKs2cc2KI5/1wqHRzcG+Ajz7FoRAi3MGTXUBPqkfSyXLM8nX2xLaJp9pql7PZ+X7jcSRVEJN4
Oy7rWB67Pm8BpWtXghMpPHvm1Cx4no3Ij23Fx8uyylTaCG++5G1mm4P0+OahlpBPuXb5v1NYFBfP
oIvJ0zt15GUQLvd+1fRnvr795VjS5njzQYx8jJQfWN0Gsao8wi1SkqvyoshVfqrnjXnFRBhSI4n2
qgJxYNzcnnR9fcP/FBdJfuAjevF3sWHWqB9XoQlaGX9wDfjJnoYYz1ydAFXcguYEHNL8pp5gtMSO
xEm8QhIyEVmez7RBd0fp2vv4M4122OLwIHMBsquhEhaF/x3r5e4Qo8a3NLUAi17Ct7iV1CWpS27E
/xyEVWdob9nBvDqUPm0dwhhfjtaNIOxXRIEBfzH6FEiMQgr/v+3w2DMQPdoTzGNKFKKHtdRepfk+
EbrGUG9BPa5TyWakOUw0/KGds5AAv1iyU1J3V97xThDHDDyZSutPmFsnRfNy4KCff8EbfOuwhaPd
GRfTfxJbvv5NrmvIqRoqzpgRG6qnbHLAYJF1uhB73jcmloE9Kgu6THqtnp6TGM+B+KkO6zdGHjiA
Kwti9D3Fg+/gGMhCXmqIqEsWabYTigNv+3xoP7qWrPe96ubl9mNldACkTfsfD3dPPVnDvGWAwP85
jl0u8NnwQ4s3dlx/WbeSaCsEm9vfYXAjW+/QBvIB8pZfrqqzXAxbPyOyxe1qtHuq90Knrx2To8gU
Ay3BKJ867/LsfQzwtbmtN0cAT1WnT37S81epXGzyZCUSc7RuycZ54RKUlCmLGGshoQVvuE2V3fAz
wN3ynSTU7VMRuTzgIR/E+NfaMwjOawnfFZZdQjP/UbGcNFa/su2Jxc712F+DCp/DZWPw483w1JYU
hRlCgtGXTeBfCSAeJZNT5NedkSRABT45zy+5VHOTfrlPJFj/Lx9RH49NfdeVTeB0zwbKO+sDwBaL
EjvAtYUQC8cwTSoHJEyPzoy118kB6IJYZt35ZN7u9B4JqhG6/rZZL4C4bfFeg8Ht39m8IB4POP2P
U1ov6vaGcbBkM2ViBJAUgfjqMn9nz1WTHZgg5N7GkLzZ/C+jZPFwKD6mw4zaOOqFl5XsVGZeNe+Q
D6vDenoSfAb6WlhAXqdR/fJJdTEb8e33ikpm2dzCHwCnZ1Nq2x/oyuBE4f7at2Cq4epqzaaxTSW3
KpIOH8UvR4gX8QDisUH9SYmWWWEFqhLK6thCns2U/GyKBm6//G3UxYq1KR6XA3E4psR8EiAcbXlY
6s/C+J+0Obxt2S4DejRMm6Gq/5SzbDVWXPSWBF6/Hea9egECUe8ZuREYoaO2r1jr+IdMvT2OQS6C
WhaYdAv+knYIQHGa9nJArPkk6hnsIqfVDlJU1uRqYtzJgYBIwijPItwpKNG2u1f8X3upSxsNh2g6
GQCVuYYX7eqoI6TdskF3NvOdK//RG/WTi2UfAZE9ELf/v5y6cJWM+jf1AqKdBuA6cueBgSvXzRZ4
yYom2t6x9En/Uob8+gxGZquB6BMI215pH/fYlBLQ080rlXgpITJxRr41y6XuJID7Ix2m+yhIgkCA
TKc3XQoW+bAQKFffGNhL0cCd2xujnxm7bVGx4U+Gnym2JBCn984Ld9Q2kVTlsJr6fSUTn0q+T3et
pa7NXfFETcCed/79f/eZ8z2fxhSCIUptPfvzfJALm3UKLkOwd4KVZXJ4relzbzMOnUKwgx3+c0GA
20D8vAySzueqC45ndqf27uFzsR4xcTgBNmPIv+b3D6kgwGlMi+iEnw7SB0CQxo1z9UrAp3KeJHJd
GwbmusI3edrVl0fHU5jC7QyKypUDIsMymtL/nbqCCzaHRwJ9NPxSZuLA2ZYTZBDXsIgqDY8CXKw/
8KEWynb/vYn4WNRuWbpUQCJ588V426lf/0ICoHVBn3VsVWShm3Wxd9PcMJxs6VBvqaOTPePQhJMK
TbU3NEfoAPgAREfBxr/fVXYOTAShGftxEUe/ymEi0SrPdNqEBAmULitVmXWChxeZN6wP56+C3fWA
sFk4puJ6ql1HtWCb0mSisrQpER79ONG8dXvq/QFqROnD+Omz/V0GqclDOvHRRQnjPpMqqJq1fsWd
6kegytK1ALlaUZ6Lwt8AIXYKxIVXNp/B8pCcfPwParBfikoGwsu8UcZmKn366rOS4MJGzUoIFqzl
YbXZZLQDP1cA8UreRPL8N6Ih1j2GgcQLAHVGvrwkZo5hUM1vj+fKR7K7X3In235baZODhOfdq7vU
mu22nuKdrUxkiE16QrZyEBy4jFUCsrqEXUiLD6UiJk6id6SVRKglFfDMX6P2UhNTTM3pw1PF8C7a
Su1gMqTK/7eya+ZDl2iY0BBpE+SGgo69SlLunOHh1183KmKrK/jMrUq4goBgXsVfNkpXeq3y+Oc5
4bx0vcpTERnA+ughDqQvrU0M/tLwYOno8EyOnckS5dWHjYKZ3xqeWP48W9oL4TakCwfyLMTpSlZH
v9vOLAgoA/vp7GzM97/LON55I5ll7zVtksQiAmnXRCvyKomAABRI5cBTikmtOfSLRSF/T5YRAMzw
cmw0ceAVzvsDI/9Gkq7Igzu/skdDsNOvM2J4vMv+CnUj/NBPb2shXZSpQkUOmpH6Y9TAc/y1WuY5
L+vrYmd+BoydNE2buu81icoYKkQVYabeyIIMyxg3+Nb7v6HY8dzNZVRavMb2rlEINiaIyk0xvYGw
Dys2ci3hOpGFQM76dJpqwCXIRaGPLZKOjX/7YmqEi3ke8k6yuSnVEUh8gW5zmysgTzINQ3Qm2/oQ
aagg6x9yPchjD9KDJsPV6g5X00m0OnY1CZwcyutjsacpIInK/9focw4DG84X9BXOyn8cFGWeLb0b
FC27mys7GUs2cYFWrI31Vh7XtqdBy/dxVX7wk2UZjqmotWNKIiGe8WF78a9lO5prhdT0+MnlXID2
lYItIo7cYPqhKfPR3PqDNDsrzYSTXMmMWb6H8fcdhxGoLsReuf7QJxiOgK+J3ZE6vb/F7lpOurhQ
tUQQvr7ODlYSYOJbttQJzAf+jqkKlNRIZL8xwVvJB6DxP7jdIeHdHdDN7NsgS5fq75b5fvPY2ozk
Htm9/Inc9KUcA8vqpblCpiCfBkBcuWGWzNeU9H9nOeWeX4OyJ6baJnX5a9bglEkK/DvC8o4RXMSP
F8Kn0jRHTeu3x8zQRex1PqOzDzlCY0zZI3pI7TD5Q9l4PTesYaAIOWz5m6VHy4vWTlV4bmfSigBj
Pg/Bh7VJ3//35rf6D2QJeDkrAVrB//N4hL1JEgP+ZQmOvJ+q2v9qluYum/+KrFtM+f/BD40f1Mkb
ixdHl0OIBXysV/o4/NYbjv4qa3ROP9MjUA/dYygb86ZhTjf1CccZRagJT/s3Mdzs+qGHSN9Fv5ek
G5/erlWcg4jIgoyQNTWeDRakQ4tNVp+fHf5WIU8eUby4HyXu4Ps0eWjsWCwQUZyouq0sqj+999OJ
4KAke7oO2PfmNZqHlG5gIP8thIB9V9py/PFreboZTVjxYy0biDxeCU9qYd9RvpOtVlQwym5qw5WU
DybP/wVoReY3+elanXUxl0M7LKjkYXzQ6U/Nt+PPiKUIlTyofvQ3KoyqUV1YcoLJMr+lkx4zzfbL
PjSGhyUtl1Ch081k5V9nc9IGmJqDjdpCODApp3XM9JZMqDZIz+HSMVqrouMTLV7tgObWO44NHCHE
dtGDYAKn5p5ovFyKvenn/kdiqTFlCvVk6q+u8RpbE0xeME0LJncOpF4I5/XOvC0oAf3O6ldb2AYu
AXidUDgEjQOGnsAiQC4GFnpUWIY3kC0pcGhQlb3j4XyrXu4IrCZHZWSGwkebsIgPw978A4Ryrc9H
CGBZPDrFKjQz2JDjdOGiQQou44w8Uq6MsgaCdnA/fE5efEX6KPZN5aHizYaLhm5JKyXVI0KUMnp7
gezko5xBZADqjptaGEt7s8g1mhpj725/L0TYCr35R8soVfgNB/qjTMMPJGW7L83pUF3aa/PjLdv5
StDfD9BZDD6rfjk+LiALtPuxyQzrswEjQlnz+yhp6xiVmRqeMWgU0YaM8ke2yn/8HqziZLqHQccg
WQUgbnDpav/AX4sDKAWGkfPDrQ9SPbAUwA5zMvZWYP1Hny4x3WGRqUpN1AaszxCaHt8ZmxOdmI3Z
pg5pKRUyccbWldR7jBJMobxmCwMV91KIocZiuro9bw0izDQwObYhlHTOBX6bsQTI2kUthDyoDrN9
8BLy55hnHfMvvdtRuIgo5XhDVxXAq/eVXjwH+8/bMct5IhtbRO6DxFrNepVJeKCs4rTIxNRqVBrb
EtH+3Za7zpjUbCwzlXsfHaKFeudyK6YK2mkfSpbdDlSh0iKoDN1zoYSWvjElBsu7JdF9YSAWvymW
+SL272G7m70NNpiCqOvNM2JnaHDVHEAea+DHXlEGBMuepT6MLfBamhVxhgJC5XKdmTNpdu94eLV0
50K/HD8JseCODSxxuCJHLagKsa9lB59MP2ZaVYpiKIXJvwpNzQQT6J02Hx63scbkbeOL9q2O2qgA
cIq/yTlLnxL3L8g5dE8o/R0vLC6BYJdEphksx+E075V1Kncpg43h+GlzsD1NSzezE3zmUcUhy3Q5
nSuKs6IVZztjUE5BKkjGOdF5MqUgbihgijcXozCex4jANUyEC2ow4aqcJGdMwOn83NS8MIv/CjCn
scuck2Ghvo1tRtFkg2M/38HqfNz+GMM6SFEuaENGB9IlaSOoNC3fcvR3TcBDExfWAFa/2L1vZQEI
EnCTBlDQrXSW2Ebc4cCvAvQ8Ixti4EtBt3io/TZ/BsCWOXg/einlrCanZrpU7G4MPjaYwzC75d+3
x8fcxGFLAV6liL5tqzv+voAPNUBvxECB2LeWeDs8ZSzXrguv2XAr+Z5deGEO3lAf9WhbY766sull
9qLBrKnKJIhzQ5JZnDowr9tg3RrU/cvczfJPoiaW2W/sCdmmAWkzIjO1sqKrNgiSAVHITmsQ3UNP
eFPzVNrN3zaccFluAmLPvrFnoqDwydqlcUZEkIrY7g602L5/eX5GL7FrbCC2QgKCBu/Eyir3Q5Jd
8rmiZFXpfq3p7ETbdrtp4qS3N0eh66VnREyKC350OXb/Sa/FqEUWa2KrkffHqpiuT1xxrqkzHeXX
L/94k2h+Q3PwIDyvY6G/JJ+ntmgLPGV/LdUZuKkd2ofjfQbt8hMIoosigOhDbnL832vZaLipR4T/
rLqEZeG/bEkjbfS8LU6thKIQlD9V4xbWqlQg3JY3Oi6B12bXTir9+JPOp0cYsJ+Fj/zwgyPWOxFF
5w7Jez+FQL6tob1vGWvH8Htf+srF/4FzziCQ7fY6mcuvtcTVPicb5/1sn5Y4r8lTzxdnMLYwuHM/
ECdlj8s1W8MdZVpulrUP3tyadgiy2+Z+1cLqU+AZb/iG+V7iCPXPn/KqWe3XfI7XEq+jbOTrSzwI
rULwAkR3k3Yerv+T2IfvfE/kjfLPwl/we6Is6euNMvluJkRY2K5gxpGuPrsODv7mgedRZf4Nk1TU
j0yfO145H7k/vL2LpanIZX6YZb09ffPm79vju2E59wgcLxv+AYy1bGOYO+56W2hD66wOEWyCu8QL
2MuMVfk/B744ZQyJNxo+5riat09DzVIBOR7v96hSmXfkk1KGNJAmwFY3hCma9NSm0+pRyfnk9oN6
O8H751A5m7mbBXaWRvUiQnQD7Fw3GvE33RlLq5QvkacM8g7hzRIMs3FziSBG32QEV63No0e/T4gu
5VUrBBhSAqLtwU7qOagV3b7UdNopccvQothoaMlJ8r7VKIO8A6SLb/5bi1meODeUWl1TMrSkhKqf
43fvXx0bR4eM3z8nHBu11LJWmxWz/+I5aWtc7RXtXGEUVAg/6guwUOKNqC8/2FE7+G3VALftq6ts
0LkAB6kA9t02QmXgaNAMQSTU+KtJ7ZtqU2Zy4yKDB8k+QQX7+4J1XjeV1oWl5Yn7Hiu5DIuqV1J/
hEnQ6mk3e0gMtHIQgBl7/++trEAOBKRqyr/RJhZlbZ6FGQAyiAe3G3vmyQxLUsYJYzswy7sz5SVj
XFq6VnX88onM/pfDD7FRAUjIb/P88ObMk8WHT9C1tSfIRB/uOmOGpjKg18JmiqL/+sWhe56sy49Z
W9UwMMOaqcs+N1d95rpNCfnwsrKe0fpo2fiJ2zHiKxDPgpThJAyoLShRZpCEebKCRT1D+zExiQXz
1dp5mfL26QKXnFC/IkwdeyVu+TycIUyjSMsqmWDRvIbrMd4HbwZBZw8um2jFDblh1G8fQTU0+cXO
X4M1hmV77qy5U8IG0TGTuBoBD2YgEkb00QkVFLRAID+5FAkJPPHK9fEko5HJqjqA8Hphx8s3PzQi
cNnX/irulHgxT0JAV7c7QAsYMmVWiafUSGJxvIwAAgberH9lw5uC//Tq6GU9/nV2sAI004q5DTfq
XRtcuFNqChLi1vYsH+w2kRP9DWlzDNM4P3CTrd4Pc5nghD+YJU+OJzVpor4ruNc2dapB6guJMoPx
bnKHnOKB+FyUZtYS3Wzey30RnCVbEZnPDPl+1oEVb1zayC8nA6XTG0Wafhiga8o5UJVhQX30qXgj
la5zPMnWbsmCB6Hkem25TzXxieAo5yeAf8+uDpuid8Os+3PLpcZtwmG/xCf0ReSfjkGw06rqr7Ai
w2K/XQ7MrEziR/zqEqxgDAor0mRdqn/+YJDd5Vucea7xcYchIYQE8oIYPEr9NfPsV34Y06dmQLUU
IrkH8ir/zFTD8LHUIsBsis5ZuZ9ZI9j3bh2T5as3/KXbCu4/61JiWNKeHbPZoBe6DKXGnf523oHc
DtPmY6bWVUju6zQodtt9Lb0v+N+4dInoBEipSKpa4v/y3pZIZ20GxTVzycJFAuRaQmm+mD+55Yua
jcnijIvcBYwj98P4bQDXW57jly+jMF4aODKOaDo0awMyQOC3hobGyflx4NAcJqLDzvRvDNjcXlpd
/JXhbO29RpdRP9c7srmAFAMDW2cSBfyWhm/wCComAVWd7C6owSB53p+Iend0gBYCvbemqtntrww+
/+rTNJG0irVNVRT8jzmSySO8m/0IsyNSxhFlvGXS6JWoJlCJhq8uC/a0c6qNK6R3XrToSp2jJtli
bXnjh8vC0ItCATcLN5oiWtASxoDlj/ckodTgcNjYmXV+Z1bwhkENE+yMjl9KjpxgqQbfiWh8c9w1
op0T9NHLzTyJArnIZt2GZnT/PGhY6uN2G3Q++O257mQ1DX6fCkcgagxL0rmuxriMSg+8KgUlcqxB
YtVnzDGH1axmNWhWI7g/7GZ6meTZ1QgDbDsRcZ/7cARWfJxQ59EQGE5Jtl3fSd7XHJMdZrZ2S0zz
qdC8e3585YADtKVJmjjeWbBnElYU2MszhHZzEcOExTYe8rn/7gHgMHMk/6IiPiAxq8MRP6DsMCpk
5alvdodl0UPSSTZUEYDngQRg3kMcrLiIFJLj783TB7KDfy538kpk+R/Q7YH6CX5/8ynoJ8tsLZ3r
4NhnQ6pWdWHXg3Hf2WgKjM7vuTV4KTvdL3Bf6z+9akpoH6TxFjYh7fRtCJkU5WfaAddv9Tj+/3d/
XnUjMkC7zHpgHdXyY6EpRasXNnC/AIIFvuTVx4quJY+/BUGcxAPeCGFun/vwhvS4bIQX1VIZNLPj
P9+I4O7aa6mxPaek3Vs2vd9lkNlVEidAKMCV7L2c3ud3VQzQHzJ+fBPrYV3j7HR3DZcZq7k+kLzy
TvGX+6zkNT5WCMMj00Oh9o33xEq8E+psSoiVp8okXAiaSZUg/+2QSCvhbqsTekCnIK2KLkJuhKeX
h0G416+tufRTOEAXWfd7c02MFViQgzGiwqHTSGUSO2WbAsWj+PPBYqQVfhmFabYQEKBOekXi30Lu
He/jI7/6dqQj4i6AZ0+LxD5BVPBH8fJSjF7QJANRVVQOAUKwjrTcqHCRHHArnOP8lhQloNNHE3Tn
pNbr+aODtecc9pjR3TZO+NTQ+5Sfdl4CRtSPT/8Z5l9ssgVITrA8I403iDoVllRLYqqCfHUPMQon
AdpCht/bdnhz4OMJKKSljHR+OD2g/v9FYvdian2iUNq7HjF0l+INdZfBlpIWRowRHKrm+ZGWAgry
xrVMj+fKNTcWqGtjQf1hbOgUrOLJPsXfWK/yuOlxdKwF0lqZZEZpiJn4Fq7oIBKiho9KiO3Gmyfw
yu9QrcUkv0Y809VQwuP1XSOUK4PFt4FPaHw8fMEZFgZWpZS5sUwzLh5rOIXPLFKj7g7U76NDxI9j
lrdW5+nxjBv9VrpCfkE+ob2KDP/1y304K2L8r98hFRIOGRRwj6EWAF5a06dxlpLhRyGwBaIW2PIe
ZQ5noQMZzb71ydMqHSaQTvLq5O9+zQUf3GwP96EOvbtmp7fMFA04/faHB0sLdhGYvmwWxzIgciXD
hT2yKmRRmTCo3uTXxYVTsJMPJTY9GmZo+RtHEL7bLyRmbagdH4do32kuYUVS8/RKZbqpclFjkNCu
mx7g3hHUMzE1uOGmEK2y0U56K/qHzpnUHcF1A/FzEC3lqrlcxGw/TVGUlnBAQBUmk7NgXiOuQXwU
3aJJlHtLPBYHSdIrfD98+FTuqTeN71Hbcc0dBRvevFjsJCwyaoC8RmBzsgrBH8gpLn83m0pPOgXs
wJPqSlNBwNoqSuErGQXtvM9U3ZyEdJUA9bMWZUhjVwUouMNrPPMVtl1drPVWhT+Ym9Tmid/W4/94
2aAr0sdiFnP4Gg42qrkTRIM1+iJWQQfnu5NtizfJXw55ggBVsStmq1RaCZvZ+svhLrvKKXsx4MgU
Ug5KhzbLYXxtFSA404kVZ+4U9HYTRBOqRIxc1piyPH6i+w0SsGd8inkT9ig9UCiO8rcttUreQKt6
ByLNJAb/7z8RDpFQTX0xzNjIfI1twz8dYYOQnjYta1TWfieF6tZPTNRLQRntKYi6RSpcfBxC6X2J
88Pw4orgiLpCUx0JsGjnz7T5uh7dbuChjZm+BJu0pk2xBdViA3jpJPNrByA1m1nzOBh7doKz8+R3
GtimgD/WVhIgXwR2xnuVMBlAfhaoDjp/wT5ASnwuq/mn9glU/VQBKbHSf28LCgYEmJMAScCJZCYw
vzIOi4MGoHpjxD8WAJ29fJPj9NkHk3hEokiqpZOwLqv7KRpwBTsuiMgUAZEOPMD4pG05Lo8rfOAe
DXg3Yh9a5bzZgkgEMscnbTLBdCX/+C48KYMHP9HUZsasiEsH/byDvIGUuOYd2t7Sj9ytojPfhmG0
Y0JCREsMPmWF/oSDxRJs87IlqRyCo0SxvHl3NhT+2+xoj91zmE1hsx48xD1ul6osJU+HEq1pGj3S
ff+wUvJy89L6QjBpYcpOkFtP2W83hRAZRbX9ZJokOQlCWPya8Phx7gbx8KcqX+uaCNajRhZs3SZg
SaLHZAla7ZRa1xSdlfL6H+NqJJICK7cn5HraLjR3f8xkqrpBWmEFk5BriNfGOjD28wid7LgVyLtX
WHOB2TQVoJWQrvpRGETH61BS39A/PNBIGQUNxCls0D4mokup3DRAYiQVHPuuQUok0z07UMr8jcon
qQ7h1kYZ4GqdKiXjFJwjjeOwBMIOAshhg4+5pvZXwoYXjtA3YT0j+Q/mpMGq3ZMrAQIgh9UGkoJT
Ua8allONf6wdk/3gFws1j9wKSGRFMUl10Ga0QoGzQXd8l8EBCjntkYhxuGE0uECzEiJgWlg9B54y
awrOAdXeV17eu01waZfu/BsOfML+1FgXVrWpN/50Escp9ynr6aDYl31qmln7J/dg16Atu6ZwktwC
lkm9jKzX6gr/5zmxE6o0Bm0HPhCaATYxqvUfkMC5vOZqziwOwFljrwWZhcQopF1xHxvyH8lC12bR
vhDB3ERjgBZk/P9UcJaf+23K9VHSIVqBURaVruU/cNPhU7KNUGHFmODjJfdi7OuRccguuoah5BqO
JTxwPYJRJFfPoNsLM3jXN7Fs0aC6Ld/HtUzoHEYesBy2N8QhzbtS/4/eR4l8kjO2C8q3YWdWeWLS
8wDjn04qXbp0FIWzR8LfOc0UF/1OvXrv3yfjVe2tVGIBP9PF4IodVQO/+cmMcFGOuJowsRCQ1hwZ
RQaLKqlQomzW8jbT8cjeQGoAoAjYlbgr6IOrb5CFBjBxkedVrG6NAPHzJd7uDM2hUWlVJ/i4ZqGM
Oe5VKniCQ2G6otYRtLx5UQgTPk9I4yJ8+MrElJ1ZY5N6dsd1HuMUBuvdpUi3MWlDdq/+hTS8TEGI
S9/BNAuOOmSz2/k5cDzVzUvaAY44oL0tUkjQciW99oEu7fSXfa0k6ZY7RfvacfNjIp4vOhhvm5+T
Rk7Y0r46EdRNbhKlVIeuqxYKiisSLoGczoryOZonvtuufv3otnNoIQ6pfob0NUXYAlNG0AxxIs+t
vUAmofHd8/9vIBmGXGIrp2XK2r535zhL4Z+grJHaF8KpL+pTeV0LfND6frtnGvRWz7S3Zk+Coysy
KkZ7s+/7IVdTjcoHxMjdNv7ysurw+QggIUoz0vgf4QRHbzV2yRNRMxgR/e2CS0CZrHKP7GUJ0RxR
1OpNjBmBL+yKYenlemN1pkNQv8fIQ8WiZ54kv7M50hILUoVYvQACvdYcIrN3QfxCRS4bLzaJ4J1y
h7Qn5Nx7GioQc0JyxzCFsuW+OB1v9fJLuPasMzUPFL5L+VYTe8NRmB3BNFS6la65RsqQ/ikX/vmF
b2QIIaQ7Fn/4G75ydZuGiSVsS2PWBuMJHW92k72PY9VkAj1Xf0PM0MC38JkQh1lxRboA2CE76sVM
NlUxCn+lGo/yjBkiRKEhgrbpWS/oL/2xs6EtatXXR+K6cJey+QsnyAdumdsCMk5YMMNfkKbg68rf
sM/3RI7KLcAputpyVu2JRvMmPkTZOcl6p2jLRooXbJW7o/2jvwLHpOBEIJ9P6wjwrPp7b3CQ+6sD
cElW8YtAaasFYaoRIbt5T0FWM8Lte1VEFixoYCVtg4ogVBdyROC8mb1FN7Qrv1FZ5LkGFv5vbF0X
JmD9GY8sc0wn8GQl2zKSEy53DtJ/kaPdPfUgarM91FdS+bQBNzTHTmXCQCmyNeofKptxkY2Ki648
8COp/oboBYzNMEDyyG5iTXopk/Nkc1zEDqzyQqmJ7CCKlQxLCpPXJBoftryoiOcXprlx3LNJzvjR
9Wni6MTNCMfMbybUMO7XVfvYJxUSgCAcgFdLfgTh5fdlRuWaarsMHRCxBPkRENoIt88lJqm3hmfH
HUzZgsxOhFctxJigO5BdDzXK6UqDDW2Km9MFDvTvmkvoztjT9qhG6k9AtGGYB+VtwMqQHWOVTgpJ
V/94s1BHpcJNvMPxGG7vtKbYRkRAFkyEn3bk7KqR68o8eeW0rwhAk4ZH8r0peW+DUwPhV7JXtBy0
mrreyIovITG8j6cAE2ndbb0CazQ1+UaSWvj9lnB6Gcr645q4wdG45tb2ZUAeXMcbq+hU9A1SQ9O8
zLpMcjeZxvODOlce9HqOfWgluChNmpj1p/KTs3KrnQ3vvfDA0m3C9xHFiVC5S+lWlhaB6QpfNsVo
gbiUuzgzq8T61ob/l2PAjUYGBwqc/XD3GO1d0chhMMHT04ujALzRLziXCFlD6+9JwT5uy22rhwda
jvSu9vBEYX0sug5bjRnkkm1xBmc4b6en9duOcw6qhF5Ct13RO65JVReQZsgaOFnKeDuqSRgUvTg9
zZJUP/0OyLYUycc8OO+1lEqXM0CTI2sokLIdKRyaJOrqrTc6ovwiyqPO/zWBtcSxIdhPnUlHTtJi
s+XQy93qYLmsZ4RTcb6iSQG5DhxPrS/K83HkmD81tjgMDb7ZkUYe6lS/4WnqQ4H42/lRqFBlro4m
HwChxkxtHT8kgSRI7lFMWdLkXMfd1ROnYVVmrki1k8TWz4rEhCia4WEOqdJfyZ+qQMGTw2pbW2wh
7/uf0Bn8SpsZPHp64+S/tTolQKlBNL+nFfZhnKtIXToyfP1TFJlEx1yO1xSS4fMiSex4HQsPKH7D
7YTAW7lJZrE5UKwUdyhNEXrElfZYwoT+rXmlY1g2gHym5XB57tqWh06QR73GJAoUipIUz+1qM6BX
5p8Rjp57kRkHjpXxr/vVEs75s9xTttSyQLR/QiF3IHDldr0vvP/Au8bhNzkwZd/Xsuu+GqbkerDG
JgoUlnG3KB7mYRusqUIWiMXTno+7sJTw6tG/QJSN3UAj3iV1y/s/1SZO3Gqvl9FEsUKmaza8gzVh
dO6Nm9vKJMHmm4s4AbFDlVg+1/F/FX/UY2sWjSFQqWEydQyUagcpydIigl7kYAVDZPLMfxn0wX0K
GjS8Nq2rJpJ0rO1dC6ua/Ft9WEKYn6Vxn2P91hIYWg+GYqy832fp6WRsibAgbQhX9jffevYYYxrX
wN4dEMl3BmTzT25Lsww3AaB67PePSvFSEpe8HVF5cuP72RsYg8L9VbAZJl8ak/lpniKJu0AsUb7e
dHWD7Ei9mTm5fIQRJWVHPlaOCqFL+hXyENapmB/xTahPpU7BkOe+Uv4ap8vhk88jVR5sBFZOu561
/Vvw33dzRO9RdxPfijJSykrRt3GnMpXBVkY4hdHSIzJep/YD9lduaetp0D22GYE6IMX04aSUdDiG
koSs4kTkueI8Za4tSRNjFbL5VbtoaETBNWz4NXtrnk+UC/K8oka8oY8IyVXIzF6P06KUng18eQ2o
A4aIa+nhzVLXie+7SCPEKCed2F/1bsLS4P8PUISOI7s07Y0OBtiqEKzjtJ/9T/CHDQ9TjWlereBB
EoP3nhzmp1OXHBcmsDSGzRbXFr7/Biw15U363xlMfDoLOZyofqJia8OobGYAZdYrrw3X3F6ibFfl
OlTAJOCiJC95fhC/RStk1iD+lows9LOtMZNeTPol37pzZDy9jbqLv/V7IUhxTfFjJxhLjGwzPbAb
y/J6xAR/JduAEjyGYaRJoZ6ZyADJb2+kOH7OsVEHfRteCThgGX9wTsUcRvINLWnGttd0HDWfTUmR
zaaj/ecyPREtmXDYdfsteubdCa8P0JKKf1RdczUBhF5j2Hm4WDtBNFlGctm5JgE7Nze0CKz2RR4w
j2oOorDpc7rHrzdM3sGO+vYUVVm/enm0KmLy/lec81NmbXKxd99KrDfCkaJF1BWu4IKDlxIKQZKx
bFbE1JS8t4eRKqfp93/0w09r1G5BuzYOEmYdRruVnGLRuXtZGbJ8W0dFbm9vzw64aplUL+OV9msU
+6p11FbXQ1ZvpI79W6EmdmreMnVhzjrOyz8vcwOwsNVCna0b4GUEMyuyvITMxMy9+ChTxEt741YH
6IbZlnBr/mePYHPLyYG4JAZtxyB8OqMlyz73XjIK8tbO4IwWHbujcvguyqsUIIz0XavlGnrm0qo5
C10BxB0yeDZwQZIgCcf5M2GR0pUYIzRiwnQEohRyYmaixx/kDeL+/CEtym3C55Ab7d2OM4mpzRTR
jjIYY49zEz8+Z5EhCdKFM0tbLm3QHdftSFDXDRFvYGKFiwDq20D/M1LLduKqHppQ8xGyLqKy4Gqr
tBFcQiVeJb+3zFOt9m9uK4UYph3pXMHKgbWeTrdyc4IPJTOgs3INtDtPOaoXUqJ5bmNLrDax1LZS
enxdIqTc6vsWhems8S3ig5KFJGweRONSHBA9S11AtVv003I69RFBDKbRiWY9Q/WgNbRJOnWeDYsv
x/3zlHQJixtHT8Z2qZrVmXF+wXEnrKFrcR9WctiVbvo02ZsNBEHD0YKW3xXS51wDwc6Otk/h6wFI
ZcoxPxDwa4Wa5FUkAX5rTMc7OMa9ha8yF0fkQXJAmZzdvU+ACEAhixPPe0j32RnzXorwXEKgf8C2
2Ot9DDIctcDrUdPUPbAJAeqfHzSKBok8P7dofjUwI2xvzcKD1MiNprA/hMIzl/El3rF45NBajz9W
7povM4jhmByCXp32js8CUF5tgV3GOcZK1UkkEGcTzVvnYedrwSycF3TK79A+QnaHRZgDEWFcNsNP
nHgrmEcxCBjaeESoaFVgNEP9IbD+ltY1L6zTXzBn+P4ol6YTHd6F7Vmrlc10A/qoyAG4G4WU3AH+
Zvh/3YxqqFa/aGYCh0xJ3DNY7XLPcSo7XSuwEmQgtrEo8wWEWVwjDIPTu8r+eixS+nmWlHZMlDHA
V9K6C35ePHezLSu0Hh/5RkGxK+kUwVRrDkLZDih2Nrdc3nR9S7w99CAlRyZyKaRFImCvgpqEGGyz
G1TqEhxOaG1LotqwpCVGmjTeWOFiOenIP01XuH3bFuvAhUw799w44uRMpVMzOmsJMsG2UUsk5+LN
pPjuAqwKQUNXFgvynU6WRDOB2JS/9o8+V5Fr/43wPrtGtWELmFtOUJOEOqGvoWeDgp2SCHdnq1ue
OlXBxsw6oQKIZwXJTJTLJuAoy4rgnzDJD0wIwRGsYoKRIiDNj11SrXCgd0yWu0ArZMGIPKv72MHO
RJhAcVH7xVgYyT7USyYKfHvKOzYtmMQ43iFefeubx4FlBErELe6rIu9hVb4w1sFyqmlMrVezTY4w
2BXUn4fc4+VA8UligWd9tesfBhgOVZlERsOw0DVbbqfp1Q+FTP9DTkaJZNZKl88e8T9PEJgxKFQI
Cy1cKTyatDD4DTUuAU6dsKWVH8k99aXOL1jD6TKjJdIAaWq7dY/V0EnLZ9t47POAkB21k4KtmjhR
/t2IWda2Lte7bbvAmZeYeb6N/1obV91Jsk45hmWB6CbZqJfWaq0HPm8xO3mLDfk2utwSAz0pMl1V
KzfN8v6YNw8wJK289c9HioK1bq+WkTlTA7C/K5LDcnziYOPQRTDlC7z1jou7gpkAplyKIXYRu7RL
fvYYC4gD8gQGaCcM+2GPu86i4ymAE1JLTX3/deJsISyeUahLsg5fqIPAqDrxaKMAnNCdT/5qsODP
z9QhF0R7aN3QxLSZu1zG5yN9rZgonTluGuIFcMatEBIqeFv+nYuoPKb/XSaR93ztuGlNL10j67Bw
2YFAbzJ9fo8sKLl1wJlxWqn/CvmkEcSAqrko421SbS19hG82gECG94XR1tWWFsWbxJomU2z0D32o
hV2mDEL66hMVyuRCTni7bvxJI3pTTn4Wb/K/qEC6JAUKq5oMePwzabMImolUkw+PSgtEiTxVIsF3
C0EhwYR4rQlgTnocQVDbdD66v0g1L9kt7QQZYwlOUz8LcBAZ61NiinPqY5uYG4gOMZL8ulVSpgPA
qMCDpv2PIjVjjbNZdJlatn0duNTwgIL+cBJdag3xJU/xrtMoQpeQSlHRRRXVUPc+x4VnWXscMbfy
D5aW+YOWJgvIBl/Y++uQN9TlnU0TM8IZ2dkYMIOPRcLzFWUZFXhzvxbhcimgcQ0/rHo5fFtNqFAW
Fo9sGO5JVsNz+Y45zL7qecr11JZcsC6YGZZtjDaBfpQ5IOemMiAgX3zv+phLXOqFFG68Z72EJVJT
1ycRBx0X+lndLC3GlJdeyDVxE7rSn88SRX5Jb5MXwQfP71l3qjQMZrFLkxyhPqJSl/rLG9jD2Mlm
AnSwejxmNwSoKxDuKPeIr+zNlG9SJJO1NOtubxPZGUCAMQEX2Xyhoqc5XVVyDiGHlQHe5pjU2Ujc
C+DSFBqHfcw35X+oNjgwW3izoHL7aTufrsYPbV56D9IhvX0fzqic1nNGNfuFm+Dzrgf+M7Xlyj8h
Z0/TNBmJkprROSqN5wu5BjCg8qP4I2CQxK8533o3UW8eo/arVd9SPjDFVrsYNOlAQXUo+RewrbQs
U6V3VQSQDldkOZgUnn2XRD6SwCwcI8Y+OddS0WUx0asgv0Qu/O88pIFZavC2yFCPqQb0AXkWggOA
bbdALw4AeVeha7rFggYb7hBzL0PM+3ue/t7GPYHLVDdtu5rLCiiRUZaGupifna5U+QbfZ4LVSjH3
oYTnLnJfM4Gs0voTkOVBPIsG3hQNGPto9SqJkSBCIeu1NJBXdp6zXpXbh5G618Tu5eu5OAS2ttZr
y22rCETjjfdo7H82dm7W8gGv6MR6w7F48GHTg9TXl46gdfm+yrpbP08qwR8eJeqttycrH0X/5OyH
IOSzR0xmnDZbzDb0Wj5OLq2klox5T/CiZjQgWL5yU8vXrL0a0tqi/vO6EP4zQNoaF8xesNas6Oiw
WiNKd9BfFiQjFr6MhEbMEDgLK3+xWUjkMSatHTffZH/cTSzwiAIgIn84+8xjyCgGbLqd8GRsVdhq
hWxqxoNEG3DvMt1ChbzQKQrEGaw+DtyfrP25SUhjNLGzwf2NQf1pRKZgXkcsBqn5Wz2O6k0DIwo8
WL/hZeEYENHaUtK56NDo1iLhefMXDJhgx/SOG1jYSGFuw6xN7Lkx4+jrskFcuKsfV1p2CczyIYFK
FftBN7vkC+1ZuXVgzdZYCHyhv7+7Ra8u3iIpWSYEr383HvURnZ7zTvcP/4T6R4Cn3F2qPyfUj769
KwJ+uFTwBb6BEKARxoHpQNacCGtLT1gp4s4T5cTrcvq8memvol4wOPCQ57KdhFlH59du94BDfvZj
iPLxB0hyxc4yJOmLGm1khlAOhz9Hsu7eLEoiQfZ1DXdixXNteWyB6kBpjwOnm48yePmVjg24x4ym
/ZvQ7V/y7tiuMWa8ZNa1yF5dohm85swqp9gaqcceqBUeQc1mlchiYM6XjkqACcHabtTsWqYvvmv7
tQvlCW+cQMvyo8PhYN6sfY4J10D0yUTTf9SXNCpw7DBuWAL93UXGOCRrQq5HlIs6l0krCVCtj81O
TVs5RoUMNRogWKjWoo+jxuF869LWJyXtnbX6sQagOgvpTZ5waBge/yKdh+dCKRys47Oh+C2d8rht
BV36KMwLw5zV+jEQWy7zqsbjAMt+fkvLsuFAiD2Mo8XSHRGXQnljeDvZsOQWUyvPKrjoerCXzDOL
Lj7GN38mwMOGO/rxoaNL2aFN0wu6REKyCTPKeRcxSeVQE517x+WBTNZ3e9J8LQNcTX6i28pHchFf
EAkGYNCv3GhFbIX7vDx1I8w+OxgL1bukmNCYBb9XOosTBfRI87W0gJ4FXkBT1IVYc9D1sv4yVOlt
HZngn6Maz7Gr2pvdC8B4wVmrFWDkI07g+nKUeupKWLZWbdkA9prqb2kMD8eb+/7WOHrocyJv+iVb
DNMUwyLmCz8JBXrKZJCFtcPvDHKR9BeyJtSY3yWwdyxk3ESM4I+ndgxdrMiYgj/EWBY/M7B0ha5D
glyLMfHDzNNEDWTABRLLslXje8cV1zutXPS6O6ixZt6UlEAIQSnSs9ogrnBXSfICtLksOep20ihT
QD8w2GLCesFq3afhvullU/mww99t5g2XvXz0A0HM/D+w5C77WUyibZacMx7CSj/X9ILJvJAXsvGb
TeysEcMp+L8+pnIy7RHwyGgCBgInMbdN6NSEtXvMb6QbStBbsUUcvUMXQFTSM95sXypz1vfMCS55
OXRpg0Xiq89X7hXYc3gwbIE484Zm9DBWsg/NBl2srFsAo7y4WVIuNEq5YVhTOQubSuSh7yQOo1xo
QhzL55z4+oHYtKUrmFCCBGG5UFFjZIrGDZr5LNR6UOVdm8H0QsZZQEC4xSA9eGypMnrtaOPcj5T5
mzpaHcOlFDASH5t880s7fKY23GE/iJIIAJJhh+Wmo7qgyWNw3XNk+KKNxPwjtkHevvo9vUr6iiT1
kfR7SKcmuL4yQHQr6xTa83EqCCvzEyCk4afrbucxutYvCd9sPRVznSZWhF/zVblzvlmuf1g7m3Tb
cz4a23IzL2Cr1Utt3hOP1L/GzpyN3zrSynkH4FOL8mrkRb+V7Qtt2aa3GR+x0QNuvB4upoXMBjVy
CIvaiHEXRPLErrmqe5PVfCMgdiGpIkNKkICa3Tf3rGlqQF2p0pyNp/TesKfa/fmSmwHtfGFsQ6BN
q19T6fO/jiJwNj8/E2uCGYaoTJARvjzOj9avB0ivqujuUFZ6ANU7/TC/g2LzGMA0XEz7I44BIVm/
v1mXPA7iHWCBKgpNDHIJAVbPeCWWt8PTvHJB8LGhfWIlE4wIrLNGmcomKE2zlSMVPgQIjrHpcfSH
kKy/X8Rpdx53MPFoihGD7Zf4//N9jdM3nxvxfq8qQzhGKGkx9cRQhFtJpci77BaM1JLNxMhax5mp
YugpCgEnfFbV8a9dN2kV7fflF/8iZ+4k3VJY7DsBARfvdC04c0kDNvp2ETrBfmhcwHZptNUhAa3w
rHKU6P7K1ylTad1aOTFR0+SWILlVzgS+sH6ile3Xq0m9mAj94k6ipSQKwPi9OhOlPEbfnpkwmjPY
A5igGd4nBb3/oO5IKg2rBrO1boeLa6Y19vWv1rqRVPF97ffZfJ+xIwPJPIgT9lJ5HCrCWr5MSBXg
aYJ68LuSoNSIEMVyC44YXjuVjb6AdSYiCWRoOUyHrOzS7DuYl7mBKEKkod6GcjFdVcRdfHqFtuJI
zZGW2iQiieQHCwOrG1W1O4dVN4F5O8jq4Ua+u0zHBzwfjApfGVDogiLsEkBMQ+0rBjI61xX1RkEN
YW4BAoJyy319QpuVFK3yun3h/xl22GrqhLsRrKRn9ndNtUJ34wueScury4Ggt/xNHKyzlx1hXBdM
fPWbZKvywCpxR2ngfWOd4DQs0NtenfI6ZhUtfadQXjlyE1r8+UqQdNMJPRe2G1f08wYnFW/6686D
A5177y/hvxwxpHEWuF9psg61rfiNOlLbd5c8xp0K2YBFlQwLmRHfOk9j8tQE7PG6OLy75jIFftGG
SdOKVYW70Cn07WFBKIVHguETscS87LiCbiqauMwdtcNnqqNZ1/SEbHRK06BgHdLM3eyepY8ZMZ8c
Lsddmnsmb4nzUJtmw9E44ZYmrtzSv2eQMnK81E4YFJ1ofG9RhTM2agUPIm1NFJbU0Nhl1LeWEh7R
3MEA1zjY04HZeAncjUSdow9e86uPaEKobita/WvPjYtdYBA6zsNksjwGjip7fhhlWQZ3tmRtla4T
wqrzzxrlxtJ2sEvGu1LWFpNNjBPrJf/RPWOiiVY+Bum0RtfHANsBsIA5gOKfAPFckvs5JgSMef/M
YlosqN2vjC/htyjMkuj0YjDldjIQU0+yENn0GggVq+HhirsVKOtUPHAElNz3JAPYyyHr2W67c38P
vyRJbNEg8e4XVzcneLXjZY5DNP41fxXVpom49ghDPHivivRdWoVFn84Zvw3S7Mb5kJ919H6JAQPG
faQXGW49XKONtg/gZ/xW5GdhNpgNcYTfUr0xCvzG9IzL7VvfN2UaqQIf1alM5wSa/YWsGTaR1CcH
BdrlauQx4c12uiMXsj/Ml47vjVJCdUbX1myiafSIauEJoZD8TzR9fsXXAgAWHO0W+7YmHlr9B9hU
2mCqFKJ4CPvyBm/aFaa+btdoUJ/AZ2CpPFIV2jej3Km0oVUyiv4pex7XjbnQc1KqXne2+FiIXUq8
03kK4AHKCffPqjERlCdFNPW9m5V7QOySVGDvz+05ywiKrWTpG1LPKLn6ZzCV3ErwZKRzGdmVVjzo
cTwbngtNLpslXrmRUU5SlrBbP0P1OmyfOgkNGhF0YKybfkzyGt8IkOKOkTnINXxHJfYJoUuaWg4h
j0DqK6R0KsUOdZTLWFK6h9DSSXRluvt/Tg1/s2x+svP8BJMUKvBUepw5LccV+6iI1sX8fvVzoTIB
TXB4rMptTRXwSJm525CFkAcEmaYlWM6VrYR3cZAw0uHHj8nwf6PBrOKG11fxb+hwQJhnF9s5rvk/
uvGu88I0h7AgkncTmxRyQL3plO8HKHew/NnhbmW1i5ERni5xQUmVE+/9dAMDLcatJ/hg3Ftboy3q
NHGW6rSJrl8e826XoRB57ZqESPZCaDn9mgPhy2xqCrwTYdX3kMl1/RL0wF4DddaRcqd8oTejuYEI
OUKd/EKq6a+yqoXADEmhZQMmMkmdvXc56sXaw9rxwz4ymDBJLWYbkKrwNcKDJc4KjGMkSmf1/LUj
MTtBE2CSX57WeQFuoOCt7wLZXYr+tyArAh57sS9HfRc79XZRZPMEtdG8GGczJEwB25KenkZHvcKf
KgG7L+EnJ4ynAJtFzIWr5eBavfU6CArgHfsqIBiRZKEW27kuuaJV50AcYPsSoT0AeVeArlUkfXde
T+aV/h7W2HmxcKXygZbLhu1UvMWta+/LoM0RUI9/pE5SdAUlm9U81o+ENJdAJWfXD4lXpG/vaxHc
ETBdferIJ90L5nbV/9RvJf/INCjoZLxjfMzwe0qhtF+gC3MTwGEIulDKf8YXYg7Jhzgjt0yVIL9a
ebOwoDFE2MkkJvw7AYkGMpuLOrlM7mRGo+z0+c2fXhSKksqD3FhzM/jeyDokwd/JdnDtn/j2m1E5
2wQMA+KEQ/Cq/9CxH6aeT5RM+cpL/n4keMMZYrU+cs1msnaremShuzWSJRE9grRSDpQXPWXyYd4m
N+zkOsYq69eY3nophgFTNm2HKaaHxoDZb16nydtFmokXQuBQ5Wb55C9dSsPlNvm2csuxRqnWND9W
BCKCJdAp6M6vju9vk0OVXBJLQFET4yVI78xXe2Hq4H7U+jqe+Ltk1NzCjAyBZHisT3VjAQYUFowb
Gt/WFKXtAVgzTNu2JLfRf8rj3uni+xiXolMxCPiBVk0EfqdIPpY5RBIlmki7ApYrYhm1oMzisDxG
ujYhsck18giakKb9yaCXUCf81kPs3Zwj6YJ/JSLwGE2bXrCYU/Zx/GNEJtkZOpIVjGhVPhkD+jE6
4GRrI4dk8B8qKA5W+sPbVUaQNYCNVP+Z2euf/new4xHW9O8BDdtZBPmxqQ8PoZ3uOj2JTr+D3eQU
NtES0nehB7Kk/UiifhSbK9LItBkv6yhqUKXqZ7ShkAjUGY8YrET80ynpMxHwZRUrZz2SA8Xr8EfB
Z8WMlo1RYz4ZAVWND39WML5mBGyQnkmGWmnJdMD8vGy3ESk2xNm6W0hM2VsuLxnxeVwkt/Iy/dA3
ZbaqB0eFPoz7MRMdXK+Sup8Hle6dlHeEVS2cec3tKbfcipiO67Lqj9fGyNkTs8043qFGR9fTJWV9
KXBIHWMQHOAN7LOwzpagRb8xVOiB6qYWHYJYcRjPJ+ZQrvVOzUXKPrEglZnn8omXPuzWfzBFaxrI
BciDYiJAYRq8Rj1i1Dupo6e6b8Dbsx0KgEvuwsyLB6ZVEAbs9jN3ABCjAPaeQ5EL9K4oKYHe18Ye
NAT4mFmxVUhSwqZbYh5Bp//rmzRmxgDLWl4DiWQTeqmCtvcC8mjqCE3BvEZToyPwJ8NCqeLvLRiw
+R5TVe5HeHtSQFAwVAoyw8B2JHIYii6eBd0jH42SM94P7Sdkonoc6PbhRnO7URhr8fmQPl0zIYNt
artxkMcpxd6Zm0BggRtdWpN8Cv+TbjEQ4ypVhPUUGkzDD3FxBEhVUcSB+FY1ZIzHAi0Cd96TqJwT
W8G3Fv4UGs11eAstVMKL7tCxezvHC/wdFhdDBYgzQWL0BVXnI7c5bicxfvbHenOD3Aa9/0z6uLcU
Xsn4WnLB01lkdR5+0IoGQnyAhAsbqaZ4maBah83J6G/+CWIxHJbWWSMLvlDNGGLBdEXBZu1K4+G2
Yyl9tlvJHx5qcDywPd1xgoGX49cd2e66SMvSD+E3OUKZnyQ9eS8iZd3w9QksxbQ0V1zx+24JDbOF
gzXjj688xBg/QEbEG+DCojC5wSKme/2NdkrIc8inqouGZ66qXcNWxRUfFZWZoS2RlQ3eu7PFsoyR
VFnqSfKAFa7cnDAOp5T9MduADjhsnYlAqtUjr/3nKc837mpJ7VA/Eal6PAyFkCBzpPLeXCHe8p+0
DoEO5Qe2HjcToN1vak0+0A7lB4MG9YizK7uoLt/lO5wmRvkOcvBjzBQkp+2WcJxtPYy2uEfKHsZ7
GWYLforqN43Drnpwo8uPo0BD8letiC1RVap49bCMYOOub/f+gIbEiyX5AsF+fGGHSbljaCFUvywn
1pZoBRCzooAK/BIYJR7BxUEA7u+15bF3iX/rF7CuKEKU0XkJ3zRFBZLUUh1wdBkqzV4IsEZu9EmI
zChMOljGU0ND0RSjICV46IY7NC4YagxYclZq8itV7zQH19Z89IblUyYvEfybCtKfKq+eH+RYhtkO
n6uMYJ+LKxLjWIg11E9kQy7csTWSqG6PlIcG3yETyBD+Wo+If83PQd2to5NkIQCgT4HdVqpdO+fc
PV15FjZ8dDH3PBrRvZCQfXWvD0C9uIWharck+dwBX5i3bYVtnyAMZHWeNqaqTADhzXXC6oewn7L+
sfgzyn6SN5ksU61u4/Jg3J2fExT4UjYLnz/mHjtw5qT+7Iiz9i+k85PdbZoUNFW4GQgUFrrZPdEE
xf6+b5YwZPmW6Nrc5iAsXI1xneZvxswE7AJtE9fyD/Ui2izElG6wte52gYSlkfTlp+Mtgrl/+zQG
tpCmjCnw9GNrDg+ZSemsHcI7II7r5KXvfOdmdh6DFWFYUslgUBdfTsyNP9wsauRmVOvTLvm6WDIE
j3wN9Nzcdle1Gq3K2na2H1i4BpXI+GTBFqUhEQBoWwccHQX56Scuw4VBGP9fQdOR7trSFKqlpjtz
wtSHPyLbQ/HZ80IFxDbbbJkle6L0E+MnDZatmV17s45f5tyCYpLv4kUdIVpn0559pQA3wBq1vB54
rKbTdRK6ihnUtkH3xNlQFDooYilKEu2hNLsLSRYdR9UlQKJ9/xueo06xDos8TPES7FexkZmEBFN7
fP2dsyqC8Zcmdo3lJiui5X6aqhvQoWpPwT2qX13eBGy/kG0ur5ygKMoXhviZbWlLf5Wo2gCdYtXu
FrBOTXTUfyVTAfU2M9zuZjnWas3bMfBeMtxK+tlrTA1aHGuiqlE3XXoX9Juzs2kF1xpSp+FAEI4L
G2M+CuDhE4jkfWpGGjYzgQNGXUxFRFCDqrMCxU4U5KeBFnmwkTshJBpdziN1fIm4zomLN/+SGVwn
0VO79ReW0TTE6ilkN7Gx4W3zsLRoHaG2+eo4hPnQ7L1CvZC7gUPa45EkS18dJ/oDA4+17lGqM/KV
+/KV5G8Z6tmgvsW15Z4RIC0bAv14Q9oFGJfApP2/zGSq9wwpmQhIsafAaGHVMSwhm29bGMk17UT1
77zN6UYdxRGsN653zi16gejxdik+JzhLfmKf39OCsEEAU4lOmr9eEw3RBCLvHMqxU4he7xbGCLZO
MpusrbJQfCIcmhclfRg+NqpYgBR/JNdP7eg847kdYst/wK+atRNspJ5UwMhoAJR0+BxIErQZGDeJ
YuYGwMVLnDwPxGx9tKK7Io8X74D1BcasKtNPnCOadzgHnVgC7EYkiuHi/TivA1pAVRUi8bHZLmBo
w8HEfpJCwV6XKxkZKgLqFELvVmhA+0NsJ/RuO8yQ/6nGOJMIVYKj89291DSCr69JGYneVzseHZtx
vDujCbmTLiZCz89HeS0DSQTIhteYCQ5Y1aGEk19xwPZby9Pna9QXHyxEMye7/AOd2OXkv3jg+bsj
8m91wVqu5U8TMoH1DNIj7an6YBnVft4ZbRwjz8XCg7b6REK923Gq8Ilj9Jm6Zkh3YEdowjlr9WNZ
N/Grh86q5Qegcd1S/syITGUfVGRv8CXeLRXIzZkRHYqsK4ytMxuiHk6t2BIue/xTztylKpYCyRBM
F9gbmEOtCE6evOc6uwiZ/g6Tf6H2zvFdvwFcQhvWZcybGwLXvA0GCaszx3sLSrDN5Jw5g11QLHk2
g//TwJYWcoSWXM7xJvzeO65kevVZR/x8SeUnGNbP7SE4JLCxX8i5dE3Kqf/tT735Je7v72x061ic
oUqXIsLNZyQ/Dfy47Obndv9EL37JaQnr4504FpIIiSSKZ+iRDB2Utc+zyurRhr2Xxm3KCreelqSt
7TbIkrY10zNnWgUJJB2iROBHr+SJxi+krwBXOwNXG0KFMU82x95rEI2mfiswcB4Rtk5M5kSzk2zu
nNdKia/2+qaHEQotwi7+ET/oip2Qf2hNqRDBDvpqin22mksCvM5BoVZ6Ni2rqFC+j43B31dqWaeP
uqcisJQdwJkP0xvHnjmBIlwOEZxwdIcpl9n8djRBvH6cX9NvWjaph68+ER/CeI/Oxx7LRPM8TqIW
LN86k5sodhZJHsyi5PkVBE/iNm4P1lP0OP4buQlC+W7ghuw8VMaYXidXLis6Elv5K1+YXfbc0ujj
2jxBA9A9X1lqvAKbaD3iniO3tL49EgYdYZ8oemS9XRmcKkb4dF/kAxj4VnVdYY87nH3JwpoTldnU
kkILkDqvwHUyG2IJQ9OrVXzLIjxrDUSSQQJARTiy0zznPpvuUr7V+C3woMcFFYvrLA3cLJWunqdN
tkO48h3o+X054KVYc8AbNAXNCWMTczdlXKu/JmB1xr7wN+yNCdl+YIsJ/pb1AQ/yymwk2YSAs9sN
4MBuPlsqoBDYfBv0NGxoz/h6AYso9HsTOICed6JeJqwMO3Je17/LOcmKDsvQvryqCLRrjrzHLSA3
xEPKm8XouJ4N9ChOEyKzLbV+4cKlm3dvTyvg5N7IGmeikUR5KoYdRj65U+0ilODK/GJoSlf0d2iW
DK6i/aCL6Bv8HAAWz7398s9GtoZaT/dQuA618bo6Yau8ULf5L3dEjBcJULd8lMao4DifZiewc46r
d/ZWlC/3naUwN4F4BCzXrOoX/m2XfURSB2JPVfaUQEjFNQJjib/5563W8fyTxEOjvTHvGjrzdtA2
pS/Kd24nft/AI4SO5AeFDG7AK3js0uFkU9v2NMiOiHHXG2iugeEJooDhKEaIHIIrAoVr/L0r/ufW
2gNqurY9E68ionLblYSAvC7qgKX0tlo+8N8bxupx02mKH6L5VSdzbbnqBGMWmuYvDrDP4F3yCdGm
hRSJPUETuEJx4wVyRjLHL8VaEIVZqtIUXxZw9uMHmjptINuxDLQT/UIY+imjlaHd2BIq9yQxztwX
m5jnfWBRt4r3TDSJ9XrBuHOLbS3gx38FfzKZ/+Nr/XW4WPyQpoFUCKYfyNeCbR6Irv0uIIh4jf0D
a0SO0kuxALfP12H1Nc32NyjD4ZvHUSOKcvkeLYRjvCbfl0bHoLqKrZm1haHeuun2HYYykSpthjYY
5OQYxN4lNA9pIVmjYAR2tYwFV7H3bsOCYAWtKliKVLRa6fzwB9wAv1MMe0k6HLG9SsEdSDwEEX/3
L3Er+YmcZO5r3QZxxl+8lw6eBZmS4gVISu5My3AdclpIK+HkE/rMi5k2qQLijIk64j7PNLpgZ2KE
dMXy/qTMUZjpo3l9EXSbG9Qb8rAbWFJPfv+3+B4jflgM352aj/oK2kVk+K5cWy80fHip1s9T4vB1
3/NV7g/ZtQr3IZrZEMUF4kcgbvP8B90CzgRuNjyTGepNEZVuU0laU0PaOPR9tU//BR1ZM9qqVVQQ
WKafVoJVi2HQICUVW5w6db9niE42SZUemT1Sm2JmTfB0NRj2ynMtBvv1Qgyud1M0rcYjP0J08TSh
Pn0QYc3WlQ1EgAenQh4SI3JxRMNJ/W0rF5LMyP3WLXm7onUnrhMFC77Ln3zhq26J7fII48czNgq+
vgh59qYP8n9HZd0+TKErI90OmsVSrwRJ6n6HB2gWylwZiSVJ1N8M7/WbaYd+ILlpFnutMxMToWkU
ShW1Xv9TEN6GDnUQWi0xp/hIzabndh4SAvMLe3HmoCRorvp4yZNOnbk9rJIzCDMVHJDuwGo91Qud
AJ2ah3g4si9wqWk+5Nlhy4x4GkdFUUmDge/uxCDSfRidDAtkZwTIEzIMR+SIVMHVYhS8rkOvJENA
Pfq7P+GkIV5m1MmLsZgor6bpT+YrEqPq05kRWu1P9Qakb4nay9qcBMtmjDqxJ9oDQcout/J2+Mr8
WHywDNyLicWLpMPtZ7syq6xYfbShQFIQ53MPQSxzkzJNLhd5StPDA8Aor2iaSvMJ6iY00KALIH7n
y9CU0z7weZf3vlPkynt4Dw8ogQcnel1N7kVCWoWTTaTX/jx+8tYOoFw0a74xdVY4BqJD7n7Wree8
TxNdNdSE3th2M0/WptNrXJc0Fby6whsguqaAridgjJPb++7pzYSiV2qEvJLPSAKAKeGDQZtxNLMR
AwIn/G+/3lh8AeVfm/fHFgdtHhywRY8maf/dm2QInppPc6RhKSym0yGm0tASjO+6Es0FHrWLwKuA
G6iuzzqzfdRVRYhNHmcrlUTX6ExVYggCOVH5hNf5aMKZoVh5YyR/5xtrS/wvCrcgOQeiubFl9WDH
e16VKiZGz+tT7WyLd6/YSnVz3nIYb9T0KA999iJ3UibUyUnlfnbWxO9UvQSn6A9zlbMfnndK431R
3h6IKxxs4p7irHPcwDGFAdDNFev5cchkibAe0MuMD+fj0DaYNhyghDsAhqyYtP3JCN4BwHGM5/Oh
Z0j0i0m3r8/4dWQOFDtbOdWoPQRc45UqP99QFhJwOMUHuuzkMPGtdtnr/oyCy6J7/vF+EMxCRkNm
bffp5BYEH7sPu4fVNSoAKB4x2poCM7e3XMi/wDltazmfyxZIgbNaqd9g8ZWvDEK8T3JehmGc2y8d
5hY/D1jJIlgdSp9NEc88A+MhvHqcIgAViP24GoLx4lTttL1YVrK9KpNaHoKxqfyUxgsQSKGX7Dyd
k6hU/W0OeNHJxB2gNR110+NJ6DSFlg7BAtnPZN174tjxq+kNI49coIb578wJvkaiRE4z6BhubEqz
wWaHv6qL2JjfuJr1N4nb3dZHJ11oSbSD7ptUzhVBseRjSEWYHxRJEWBznzyMiDpQyhOe9IURELeg
k0zVV/aL0r5v5asjmUp/c33RieIAVPqLB46xdgAiwYXCBhmDZQUm+SL17VDnUVj8YTkITOOJUMyG
q/7DbcMLbDAuXiXQzJjMQeeg40nn+LZLfq2QDKGhxdoHDd7tw/k42Mvr8+/twyS+Q4JQNPRmfItg
5OMoL761L4QgZ2TE27XjrDCoc6xR0c/SQw1S+kgw4aDp5yVCSPiTufA0Cp7+ph1nJiUCy2cJmwWb
hUYBWcZnl9tJTL9mphKKJL4Mch0Zlj0JKX5hd2/Mr4AfqhUR1RrxXS9sUJqDnV1KnQfcwikzMkLz
UryFYklG/Cagb0cLQnYZN04jtkCiHt0VFWQveXS6I85dKkXKqG3iV+dLNFgpmh2kc6mHd2PtEopL
PxUUK7ihnU4NHKMdd79jm5jmUUWYmrbmMzHHGRZPILrILK5tNCUMMwXvD3dMFXUTFZ6F9IAprBH6
tdIJKxlyiW+i2tRcge7L6InNQ0k8GTD3aH26f5J0Nx533gkUXJwYHwqjICIVw3N49KfzObCzeaHF
af7v8RIQkN6orFJQaFOX2I+YcT/fUS4n5m49+N4wuWq4P7L0zB3TzhmHztvGpagWAJWyaO+kKcmY
4e17mGM5sVcYlg/weL/aqueO/jhF+9DSOjrOmBJ9+sGWJE4SDHtwKSgxMqjqeYBSyHCnfJ0a2ddL
IUSwmMhy49ZGZJoQ5iecfDhj8Favfk4WsSygVfwtvKb7f0U/XOSYO/p6r3LL8x0JxOo7e+dbucbi
8vhayojYt87JeZyIfw+uxc6INxc3At6NICfMgtZS0AkUPIaBe2vJsBOULfzeXjUxbeNaqo+bPqcx
c5dY1xFviwtVhU5Ox4Mu8haoKQLbRk00gmPF87q752rNCLctAetR0RzH9aq84yHQUefYwccJiq7P
36EVZKnoSvKoTiYtUe9Ds+PRtNXl6eImRBVTSuYe7D8lHKmdRUeygwsV0Uo9Qw3fKCG2R74B8LYR
UeHZxBjuAG/kWkcRAT8u6aqvFeGHs7ulL4wvEzX6YUFxDeewWYuuNuzmWw0o5mlllkEzcbEPF9Vm
KL+4efvFrJIxv1GVdYpsrv87rr02x/JDBMRxlSJHu9Yu/5f6WXlCGOzGReOPx/Ufwlb5ys0X7+ck
s2V4rwGOC/pVNFxDOWQWcn+DSMCY8iyisAtbTRWMpsDWkZ3NiILqkD24Lw8ppFJdXVD96BhBz42N
lJi2kTVBD/IZ9OoipFd59TFP6hbfxbCzpkfl81hx/Qn2OxkeX9m+cwgx0NP46ph6xRRky/xUmzjI
4zpk/DkHLiLh8OoilKnVEIl/GXSRtej4yOxQ5N6Sqv1yEZB+rUOUuKAwB5Vu35em9cLO4Gb9QQYX
aQLYByL3grboLXirZqmyRuPT1J7NeOnb96jcKforiBumRXTOMPfIdR6x/hvFWPAyfQRn4PQuqCMf
pBFkZAUVry5oCGmwlOm1yx7wDbjMBxIHVsfqiR6Nm/ML+48DFtqeqGyNL9a03FSv4iVePvYBTk/z
TEPF28z4ZXHeeBam5OA+J1B3mpZEAEHQjZQ+ZSsBfuAeaIyt9EaYbHLXJjIuEy0zLbTrQK0M55dV
qdrFEJRQogmycEnL/SdQaERebSZJVjJYBeYrfIDvr5pb9JKTQlyxWfEeMKbIeHzZCMYtZIwcauXg
WPIXeythOq7RSL7Zx7iecAOAlZQBnPZO4BYdRYY/Z6yJ+Up0N4ocwui2lsR30sxnlcliLGZGzJWv
o8RXCj+eIV6Y6UUh6o8l0BWjc5sT5M1UN9aP8qxY3ntC0vMk6wvtiuttBABfeXUBI6ZH9Rngci7l
1hNfa0tRLsKgE0qHutLVx1UF4NmSGa1hRqboStK2fyzvo8jhI1WA4REz7H9ufb4fa63e3QhW0Vfe
G51Olh/D9fjnPawLOD/cdBbTUNluEKpRimpVjp+FGU/vR8BfAGMiCqycIKy8rllxii9gebwyzHT0
SRu/UhGcXL37arUoa6pjBfdLbNCY7ON3h/TKpajfVccNy2LR350182impZbqy6AFcFR8qvEsldkF
L/k+c+18F9wAebvJeo8+ScAYlMtzhH7wNzzc/wihJrfiwkQN8s0K2jIzuHiVRX7Z/6JpMwA8UrvU
3epkQ5zkpkt1NAGuOwc8orhobSF2pe8f6vnGMm4A9zIShmPrLiq0OsZP9YQxKEcvEJOOrnC+SAdv
LEzHm50N9rCgFXh6runyZj+LThKLXnAFQdtH4Bt1o+JtWQ5lFYIpSnFYZFYypPWMTKshtXyeAnoL
cjdWGwB3ybPD3M8W9ZELiA/GB8+6QB50Abvo4ZDmvRXvDhLk3Yi5vD5CCbQyIzwK2T67QVyXOFCj
oh5N9PRIvIT9rF7qj/1sOYwOD2TWZqPldwQnPxRHoX884Wbr30LqxjVNpm0mgW53hc21FQ3cquh0
fV/SPW7fDChC1i2VtC4+qV765wusjCjJtgYnVhJNUyHQGxkJTudMgK5TePg9nRA8ksOFbkyP5EAx
x9ADAoCZzIUjp2e4XdThJH18ayrCK3SWPbmvkpsaLNVBR6PmnGU0/IuOMe1XEK6rFtBLCHkp8UXB
Hn++XRRUjiGh7KPr91P99VyRDloAkoNuWQmf7ss+z9yGfT4gUzPnfxxermP7Lx3KYQGFwkU6WoRp
nWjEN9U+cwsgSftu3gOOiFhquzVD0HrmitjKmuC0vEiyUkd6snB4ZWujfgCMRqrki2GtbIqAy1v9
eP9X/fWHSLPPaq3yWnlDm6gjUSuVt+xuX9RtSHx3l9KCjBcDe6aih8M7159k9z+HA5R8I4x0Vi+Y
R9M5gbMTvahOOHneu/Xl6FSerNYCRAK1hMsNqjA4ulDQ6WPtuw6dyIvcsYvjLwcPzE3gdBu1Qe4G
V5gI3OtMXdN2TR1VBYW5luT7zPnqqJB8XarVCxDItPUi40qF0B6TWXrA0tU35Q4EK2Q2JA4WcTy2
3wtuKBmtGrL88vWz4Np4D+NYTngB5TQ1ZYgrIjzzkYqOKdeIv9Kzy8ADxemcEXUkj+/95LjpoS0v
pOlut7jkArhNH9hc7vpIfzkH5Q4xLnkjZ7lCgiEt9/1NhfF8YQHR36VA1zVADe394qHUf64idgH+
DvdRurqgothZ3IkSgnfn+BUiyMusaP8ClW4NyZU+PDDccJZ1x+TxvZst6BCb/GBf/encGLEcunZw
jr+xY0EqIc4EPnd3j62i9pzVKjeKB3Uscw7zCZX8/tcFEWjwdNaLv+Ko8kz+fOa6upAn3MsuwwXk
H3EsAUGqvhbZJdL9qqXYo5MGUiJA359jnbHSv0AMh5ngLfLp1HD0fO4zEHdZhYqhm9H2FGnMBYPT
m2wKQAxsPaUdN4aDM4wLLyaEA3t85Z52F0xJmRdaXYzghLIirvFAJu8ATRkPB1bilATwFEWhMpoF
xWbhA+8wGw2UTMICUDlvAfc0zfoOcREiCH6i2OPtPlqecABfqMq8kNUgoogl1iY+66KZB+oBnwlj
4x61dqx7zED7pPVUnddafNtlp6hbx6X6J9yWGENhNn6DhHLtefMYfs29QB7guHwvvdkmRfx1gtTy
vOlWl1TJrtpuGrDfNwmftDfQ/eC3ObAeeYH4NjwdosPsik6QelUMjotOwNJqNkep4kyDtR7jSkI1
V4AWuw+W3XN4boAMmveZhkx+RsVmi6RHdqr+9NesqA+oNSr+ui/BbITnNDeJwkB496/vUPq3yF0J
zjkFB0Il2C/bsxI98znl4mFjWDSDthQVgyRAbqeAqiDXjT/eRJtR3uGn4AiLFkk0wAddAVC0o+8o
6lCPvLZZfr24JWIfWDBIORnODX/EzrbhBnx4YpMmeWPbHPCcnYxTT7x8A5DTW8/DNR3hXyPnCmuF
XBGeu+6SUewLCY8vmN/vbQU5JBY5sO257aQrjWyqTkCTpIOfQHGrmMbPw4GtNsNe4Iv9wBBzjlE4
gVNsY0XV9NTAphNm6am/xSkDQ6xwVmOZQgqUMkj/KxfsCVGpbeD4e0NDOzepK8iCLsVSGNtGJprt
6DW/VMoy/r7Qlaa9Fx9cA77Zr+Bz3usIcgsJN5sd8naCTSodNh8ZHSklfmoR51Btri6yIRBg8H+J
M/KjpGNUhMI+3N/pQca6Iq4G4rP9dfivuxcTQFQsBFYkSOSrcvxazJQ2S4xdEVjyn3wkMk6PbeYO
282MxyF3RPo5T1S5xe+taDpruGO6v0MwuVaJGB6/FmxEJKJyevKRn1mSKL72qdHJOBiEH8htN2Gr
gu+YwSX5crCuUMIuyJX1bNLJYHJ8Q2KTugZG+3vGADiTZwew+g3JadGyRyuZCU6nBoKuPI+XDrbc
BALIjcRBhgghtmS1qbRettVYpliWLJ0IakDDYRqLvDYNvMkL8lOFx7T1LTZtDk1LjyrYPrZ9odhZ
rrbQrqBkup7IdU+oAjuNsG6s9r2mwawOiysqs9QhCXkrlOj9FOmsnDc0kVL5mqplM2/X4/zfu6PN
SIljqVdCfEkt/qLdrFrVOHHbHi1VK8a0xO47n3+tNCS8wrl+iDRrt3xs3waSx46Mq2/4EnA/ekkA
RPQyRltqz7TRs12iJQ44oLspupWXC+nDKtHyC1ihsZ6Z7Bwb2cRnKhaogql4jWejSECiWd9Iz6j3
S3MxXoaTXlWbRspWuMUzfGscSZbdZkelqbpNXD9dF1KXY0HRLx/DEBhru2FgE+1tOqFaM7YkaqsT
rOafwhGc5urWxOVcnCWWrSw2u2ip9Fa6bcdu4XFw///5Ekd9FKCff1tgtTeZ+V0/OxZEuaZcLj6G
uexWrJce4oKQsxkMFW0YrfY6Cj3JtGEe61TkIvQgWSIuSt4XAVTQjyZLfJfk3fXhK9BLM3br4fgT
lk75uI+3/5voN5ruDp0jMqiTCFbNAJpWf2GXDk2Fe0HVqvHgglStbbA62dAbIUDmOoEXbD85qEOb
GveyWIoQwkkKd3PD71R+xvuJ18SQnPX3Ry9cBEVLTftOuD5Ec98DR/9gZmrBfmwQIKvSZBEow4sa
dxifjKFrlmhA+QXvsq3hkfxxS1jvP1HG3AWADH5KBObkxLP+00UWSUNTXDf25rXLRXHUivLis1b2
NkEZ/aAe+yzJoOTKFrnHDehcXo6jWGAfZtxphvpcm49Aavb+Pqza4DiS91MHJD8ndoSGqWUapjTG
roa1UiBSsDdWOGkJthlh59PmblVKFyN7yZ3BCtgwJb4INTXLL+jPt8L5vRn/qd278k1ykWqlrgYW
g9OgH/cFha/0hi/rnI7+Syk5wP6dypG3L4HwXCCBPbDyEcLE6z69hyEaxSouUCwFpwxE4pbrrDSa
plYDBaksvl074uNsbej7EsGSyfQh0H881G7TsX+VSfia59ei9uD0HIDsPpVvu/tw75PzENKhWObH
j3AWqwIB5XAaRsCfaV+BKZcArslBYyVYB3uviKukN54yX/OfSQW3Mw8T0MEljHFQOzDh3obVfC1v
CHN3Bl5zGWXxXORf+CxWxUZkQM7aAp+LoNTmirFHFASxZaGfnPtFOXfVwJV/ULbuuVPNJ9EMka7r
VO7fPR7yIEUdRsvl7Aw5y8p0GdCT7q8jqbCiI9kKEKaaOWGClIRcg0it4m/9B0/3uTe9Y82Xf3ur
+fp9SVTc0k9N8mnqpZZO9Fqw0xiMkvZAjo3G8qux2do2IdpPNBayVgaoqadObtK5pSRvSaljI2oQ
u9U/B6vIHUVwpFIkjCB609NU+YFAcIL68+Bkq81/QiTHjtEt8P+l1BiE2HHS/yem0r+LdvVFHW7W
WpcBlkVBjs7gpW5LmCfIplw1Y2aFC5sqS94Y3A7EN/nFefopECur4KzLeGDER0r7EM0V3tubLnRn
IlvA6uVHjIpVIlHNoNiFZtBqH6d64ri7D7Qmz6wZMc3CmpaG1rzfItGVQUmqvxNSrmRgfLb5515A
j2os/N9/JJxMivPWA761NfB35ic3NBn0BpdXDDYj6i40g3ILHJuDEqSi2RREES/Jx0GRI/TpuyA1
A2yq/qJ5LjSXTE2ZLBwiTrLfREFr6bNMXfGCLHi3XEHbcOiy0chreZ/q+5FcvIwwworTtlwbCElM
RYyhNAVnTJjrRgVA27JsCMDmGw+Zv0RsuDeJZY/TzzygOXC9lB/7aIcIfPXBH+hv1QYWaZjdSn6D
/ZjvEETlaaqe5Z7jm57mErgFhMlqJ6sb18jIple1FEFXXCp3SEjYFqKLZGg6Yu2aaPBE3jfq4iFX
eG/Fd43TUT63UihlhBokz/vD8iPEOJftwQ02LZu9aUy7ZZNa2NPrRFs7SE+kBXaiqwQ9Xc+/hiWY
sl3tjH9G0/SOVCBOu1QJ15fqNbPKllZYJCKzFzMio8PnWtT3FuZuV5DBWFN+lyQ+OvvSLyjGZofv
uEIZcOjbyNGNXgzr7gb9UUfQ1TEaojC5Cj1pNUtUEcD/RKElweXop209tXyVQlvHoqKEkotb77X3
GErL8pPYItNEem6vKRki4Utj6Y1BeskpaPUS3HFi5KTRfyJofc0xOKuQ/HwRLWf09yGZWf9PRjH1
vMOkotuFKWT1lt0+GwO+K8RPbwOrJix6nt/sf4szuHmuSHy7esCn50tpqpa77Oo9uKaT1k+pANDE
pV7BEJb9F+LJh5Cj3f3mKwqO14d8feyK2QIREoCY+7kc+ebKNX/pl8+HaoeZ8cdDvoBxAIW102zp
eucMIfa9RiIX5PTdpcSLJxxC1Sidb4FaszQA9frSrPmlvWDEbB9ajnC7Y7709e3Dpaz09puIXVWJ
vY4fB6YABXF4kIBEHo7f+0hb6P7weI0IHxnZcz/PYlBglz9u3nmT61IEPJyfUpTVZsUUsdq892xn
+XIS1ZnBRehbjFjux+IFfErkb6E1XB9KLHOFbjecGKtq7GvtGAAv4V35vDZZtSzbtZ53a+3ThWaQ
3F04aGx1WGJOK/cDo6H/iCAIkQWnK4Prmr5Plf4bGDM4xV5DuNu1UbZSPqUoBFqRedkRNCLhR1oB
7s+ZxMasjxeLbHgpNlJlllTuaJHjNHYrSR0AU+uAaCyVFX2m5gk6qFYwLEJpObYdBBEiV9FvPfdE
V/B6QnHwIL9cbqwLrxKbLGMyn73JngazSdFTA1hm3b6L9wbbLuVDTIDR3SQ7d6Opexc0ef2znI5p
51n61xYtNcFOU1yZQxGV7lBWHCkJrgrwZ+cL8XJUEcv1q7VlKhXhImvpz10aaNISuQhbqUUk6X3P
mgjc3aJM0DFHyLlNOop9pRxf4baIabYVZBXbhRKa108mhIH5xlyhPECn26DMo0hqL+5aZdWKYn0i
tGDw8lYQpHaERFOpxI7qIJZZHmAVoahkmpWscU3/F5zbuoTCYjw2lGBsaMba2UICtzFgO2QsTuG0
yvTGAybaLFg67vXAUcNGizsU5wptCGe1uLQOIsvwbIUWusGgL/p8cpOCuWsoTu1BSqMGxnJeL5bl
UoNJ1vIyIyRMpTkcMAX1o9fFVss6O/757XY6C1GtYMp9F7KjMkZeD9BSJdfn51PHXcIfhpso+BXQ
UkC1Y7+CmQIRWIXB0Po4y5zaSG+ZpARanZFyGwr7aNnp/BY0pDXv2ZHaK3Oo9R0UzXAdTjcq9CB0
d/fgWhNXCiRQqmLK5q7JwgsUy5x0Kz1QVlk8dIPp/lrzdggJYxGMUT/hMUHefdm922+liAHJAFWd
tnrqxPOtgOhhE+uoeerll6wJdo2Rz1hYvmx3s1iOYBE14lKRStEKnPx9Qts4M9bSWjxMdL9nkZFw
UrPLWz8qHsNB/OGjyTdttEmgTKvgXgCh6BqvRzg6ZD/F2M2aiPGzbOXRgVMR8rQ/qeSega1GYdtA
aGhJ1Fdil6VpnWBjB88f0DF616T02hT6MGEzUEO78BXwm7ey2XXp/HOICvybHCDuoTdf0EQp4f7I
X97zyE0bkXqohzXiY8JfT41r+qZBG5JTdSGbMSVa8flz1hfkulqtTMCmC4MY9CzEoDdpqyfFsTmn
vRJmc4X/7dHePi790DFu5UHOy/Rf6EY/d+7ehKvAyeLhwxyWMGPq3spNKaz4M5PCXfL47bZMqMZ6
cuT3AR5I8kHCsClmiWNyMzy+6pIO1tEpTGelmMR2RhcRvBE8mtKxVZJ+M/N2kricsDJLVBeVo6sf
zk/Kq6KuQdfO7UcFRvWfyAbi0neqHAYKA06ucTPw9prG0472Z4Z70OJQT+OnIO+dv/hgKEFlwFZd
WeUy0CiR/6Vs7laJaUhEtDGVODNfiyihZTD5uXd+G6som5NHFt/F7fL12Yzj9hCxTOQySjCwm+na
QRdDOCm7ApPCnKjTrgSNt5qkQp9tyU1/H+040WyXotJPGQ2t1phsHDEvE5hgRHvM+bgri1x91r6K
oWhM55x0ii1fPSpK0qSSh45YUzRwPCTrZiPvOYDPIsYUFOzfQLDgisjLhdKZQCADynsW6Fdd+n7U
lDzn7+NADJzkJ2L1RH/NwJr/K5SysWHTC4yAwKIWx4wc/RTOKOoeXa81OIx9aTtpcbysYSyNi5hF
uUHU4LpjcxV57rPub6AOKqZgpa4MxOsUXkFQpWTOjkk/XjBxJsiBUpL6wXTq4/qnFcGP1Msey/EI
0IxVxhexkrHIsWOTymhLSwkwjsq+ak+hWiW5DTe5TIqEqqKeO4+PO09E+CUtDLM1b4XCB+eJBliu
OCfAic//UctDqFblIj+wVyOXdZhxirFBDpz14JdOwzHN8hWvA25l5pNUU/sUdFwmSWp1RuVRxbuz
nXQEx45eHY8HyXBCS6y/4TCRzR1DTFCNoKawyLQiJolYFjNEf+ADcNix5h9Uv2MYDWHg9G05wMlc
jt80++EgRnpAouKCfC42YNL5nixUh9n+lneARu6lhsvJpd6Ks8+5bL6Wfln/4qMJA1be9moTWi69
DXfBLASXtYAY+L8CiOByFzz0hM9BTCxuWhhKsSxiLeKtXvoFh002OLACuU3W6Qks8PbfDK6ElbHL
4ZFR7e+F9Rjs1pRFGfnq3Qev4f42hYqgERfutM3T80R6f51hhV+ILsOCY8ad9orqQYL0vMKBilNE
jca4D0um6HcBw7SFVJqkrPy5Xs2SxOQ/pVl4kguYgCrpEdDYzi0EdKVF9yo6u0FPA+NhFJcn5CgF
Wr+kb/abPr53wckTFknV6rbaWqoZAPf0bU98kQOSlzF8Lr1ZfdDVXZhIHRa6RdyoYUCI4oq1ocXl
CFyzgI6orZKE73tFjED53ME6bYyFZ6raD4fmDFduGY/9EJKEHHWd9mrFgP/mvE8kBAPdleiTv23y
tB+/9dYMQU5kNh2lkV+ahXcJkjudYoTPry9rpZ1DiPQTdln31UKqoPuIz3sKfvluimAzqbvz8rtj
N9zhTToOTF+h2AxBTL4sy2ak+s2gu438pUo6+qa5MJuuUH7CC5oHJuRXjcd0SetPHOuCkOFupdKw
/nTmK+lpt8RW3a2kGdAr64ydK6tXMEnoWvfva2C3g7VEP3OpM1lAOJA6kfFhO1mxTgxYCTUCMjLK
3ur5ZW3CvMDRT2EbJaprRwaG91kKRLyPlMorTfafEK1ASyTzjVw0DMJFRMvMtEudR8uyrHgITXik
yanQU39ghT9mLCLFR1+NeoMX5xjdxdKRxVXqaU5Gn/C2hltG/g276GWUvmJkaOjrPsf2wf5ye4hZ
o3y4RA4LDcv1D5ur1dqiPnbX3ARg8shX2DGwj/OpMsF4LbapkFLvrWyN3OIM/YEwwqRbGebe+kxi
/FcOty+892zXIgBP5WTHWLagAvyDLdD8rf0IrscSu3kRWtDCOG2qp/F8XYt+ljnwbzHQngqZw7yv
YDoP4xGz5h982YUu/3q+EBIluP2L7XY1jJg2BtV4c75s0uKTdSO834piFtoYrGc8dKaewIkPDvsF
vTHglrltj4XX2IwqMtzmVBZ7aiz50qLlbNOXOM0iJH7IP9ZKS8vrL+wwXPzredn40sOSwklPz4bU
rdPGPn5ymDLKGMK+6bIK0OMwDDJ4z6JRhgxs0qDQgXuACMu2/6OFpM+XBxzS0UZUz5/w4RmBAkcv
XjkaYeqb1neiMJllTAiiL02vmYDya1L+9QiF7luba2gpQZPdIyzUMcYkXaEuLtyq0gtlBshl+MQl
aS07jZUnRggSscvfWgZTesiP+zU7mdOOIkON5/fxxMwxafWCX+eQXnFB4anOhlskzSilcCKPkdP+
QoHRaNw8iIt4bUbYVwa+VL3VOqpAmhrQHPLqsF5rnw4f22MoJw/d4uyaXzSPxRJQI/WC4oVYIyks
+fS95wfrCLNYyYXPcnwSb8yyW9z3rau0URVd/rW6DrIbiubdMCI00qeEjLJEL/G2lwO3wEWaVb+w
lsWbQOf+6SADO6PsuzUDZWJA/TLpVLKwW3gOhDp5GCJ1ojGHPIforj6AbTFP7aL35tpyfLQXE9Gl
MjtLYc2uOjhusUgmaG4WsrNjSVh9/h3yXNKXGk8ct22yBhBfIvwp1Eq6lFtxZ3Xsn8X6m59bMylK
RF0IaRD23pgMzLWlOZH8HYPWGdL185KUu3F3o/F+up3BilrfxzbawBmyWsw7uZ2zknw+Wa4gCsEz
Xsf5SJZkOZN74hkL+IL+nGOrj9N+uImLNglmsFss72WvsGtlxMwEBk45aiG5Aj9hEYdkt2cdTcDA
7nCZYqWTMqCA+bAnyt0TcdsHcPV2LUx5Mzql+EyJmSJDk5OxIFbc+zj5PG0xlTnIRnZHqy++0LEi
FLa99fd9xQvseONYbAchtrNtBi1oxs53GA8g/VEr5FiFFnroVpJFSvyR1cnYNMimT0KevzY0FWfg
Q0qHZt1BwqvEU+gsX0wTxeOna8WRUhiLVO05/h+updz8cSy6C5KTBYwkw8beCR/Pw3nYpgcx1k7/
cnttiAVfvztgfOKgGc5NV8rmqBZ9Ol/RGLl43OIRPtJYYbVj16xT3ZUSpmEaCCoCGv9KN7YjEXJK
GUx6NnEZfBquHx2H9JwX9tX9t/sV8plI1MZvP3QCL8ng2qvvzS7/T56bycQ7PuInb7c99zkp1XJ4
izwZJPjxu0fC4uDJF7FGwiZYKscvZop0PL/pKFPDw4RbyssIBo4bFoqYqR3daplBSBl4Wyb6Umtl
5VRkf2TCqCg/mxsXVLSgEPjynv8d8oEbQRx1H3wwFkjcy5eTckfl5y6Zeh18bN0Xjj3amb0XTDs6
XKFje/JIUQjImJXOMRYAcJDgfAVlaTg9gyiYu9aqdX56zmI5b7qjY8BaM2X8n3BCRUUBtuYkeW50
rtLzez2cVKF9Nv0j2myNGOtZ8w3CYsQ9Wkg3Y8JgDacc8QQk8d5Su0FgQ1ni9svyoj0nfPJAeP+u
Y0kvi51cJTpr7cJlpk/5x0mPPtYXDvytypqWKYlg3EvgLZm/oi8iIjpPT46d2I6U7BRw7maU7aB9
vdVthBvvTuHwGPDgJUczKLgCuSlOVMPFz0Fg28437rwoEh4/sF4yvhh/pzwH9ts7cCwuRrfarETg
1/sNObO3eXYTryj6G2sGcesI9Ii9ZKDf2EbZsrqdurFnsQPmg0hzKXbzNUZNEEfDkf2Jo5Iz1xQz
Za4qZ9xa5mLDMEON+Prdefy9gw3cC3FccOryQrtFKx21JrjJK3CgY1IOqHzJUuYGgKkOWuPjciP9
vTtY5wT5xyBspt9QHRyqjaz2aD/vGqzE4UbVxfJO9LS1lBWX/DyTPt2SYxXt3s2lNibN92YYgzca
uKZuFisSoVEJK5UGAfEHcyL1jbwLUvv1mvZAxmfAoV7OPBbGHc+tuB4QA+46/uGQQO7F9kr+WF1K
/cNjhRLMmhxx3D06FdMb2frIRcwZ1DlrnqL2r1X93lApBzM9S3f/Qu4PawMaB35CJrPvX/Y879UC
W4VyK6HDig6xS6oqm5FpyPBdsaWwSeXFrJ8YT+Gg24VfEUPYUIfGuv3OyK2JZq8TV7CqyE5JomPo
wiNKkOWa9t9Pgdie6TaOAA2rc+9yWExaTkIvAoMKR+rdF2c7msFGE+x95vKhLxm+HbSl2Q0z4IhQ
72HJtEbj0KM2eFKsSKTidxcXuNBbTFl8aT5TiVcJ1Mdf1Gc2QIyp7AUBWkTxfLcIUAdcq81jVZ7J
J+y8nNOfZ2jWTGnZm2TBa+zFejHLbDIEsQDmemDNU8qwyVcdds7jItpbUVZAgAZskXQVRo5r7OgR
AdIob5avse8tEa80Uk8KhPgn408LhqsGOmsAfkn7omHKPx28BeQrESf/FmKWPngEQLaNK6ojU4uS
rHMdskNffXOU/vUq2BnRO/jQN6RuVdDkSLSdm3f+vonpY/+VBSMHAKuz+qQNg4umRsshDMvGtepV
AE3b1hpV4Nws9xPEO9RSMeeCLPWWf/mJa98HPDfzuhzkVZHn+7TnXjs68Wte33fAth8E4r9BDECT
xjpaHCYs0zUOtadg3WnixzlXg8+RzyDcYfQKHI8Kq0mGOsmTDHVty4jYU9B82RDlw+qhggLFCatW
1UA+uj7Ypv09XiypCgVqAF4+Bn6S8J9Jx5sDoVkOecAZOXl3Xe1c0qHAylxCZZZcC7PkQz7YWnln
FVG4YrE0cSxFx0YjhbI8TgInEsTrn+VDVamhJdtRuwwEgOFFw4hFZ/rRp2jzoJnl1Qws+ZqgjXk5
h8jcovXQ8+djuroNYgAKwKY8cRqTWI+gSwlqzFUYr7gEYnButaU7ABug4NJVdvd3oPrGl03pNzdE
WlfPlc+pdlxkBbNT+2bxdjWj/HJv6FWhz/HBQKeevN4O294V9pFHERA0TOvMqR7dkucVD6nwR+D3
VxAqCeEXFquLtjQOk4BkdVlV8uP9YMrM8ndeS/6rqol3gDb+giaPXbNcrQ+0Pq8dVreMGubdMDB2
YAmMUbE1rMViowvoj/tu44LYGaG/BYDVhCjSShex2BPrvlHyFcgCVOnyc0OeqJFh+bf8oX4OZTsL
6KRveoMoAFwFbtAoveO+xH//8BlRldC1KFBYKI6rQqzGV5WmBd7K3ejsRKBptkV16EeAOgEkSdIt
qyNZ4B9lFlSBEFprtjCTeoE0Uq2jeNIJr/N8M9z5CxulszQHuDc/45pm8/ieGraOQu/YFpF7pGpm
n0nJRZ/1kwo7uf1py3KlN9qlqm+ZFqPKsAtGt+xMcQZl5GCZpSlbPGF3JSP20YxE616WIsBkhdeo
hYB6egqtEax2jGrmKj9KbDugmFh+YhQQtBeCuN4pOllkfm7gocFJ7iAtXTDAmgza7zOgpxECcaY5
VXXXq1RXl+3HJoWk07e+SE6rybFS5GkC3zEsxumKVREa61slHd4/jr7LMAVkoLAaWLp9xV+FxQij
+aqkoe9Nfd4N5crM682kYO8CpFKYF0Nj2LKzL1nbCkcaSY6ndhd3vJB2HDuBElv32PO3OpVuzpKs
hJXpYBd+GRRHyi93GNaGv7s0HsFjsjpUN9hqx1cDLyArWQF7MfwWQhVXibwc8wCLhGcmtlnEqDKk
Yjn5xUPvdy5xB5wo+iKnB08Nd2LyjK+S3yFXPlcWXSk4C+bC+tVJpef12QNKs0LXDQkS4oIASn/z
42q5nygcmZEZOX1O/uUuhaqQEUerkNm4cGZOA5laXOP6Wkvfl6yF82REc5bM/8DiUU4c8Ee7AGaA
2wmXA/LtWVKdNJwb7mmzKOey6HGRYkGeALY3AQuKE8pwMKQLVK3kCARvGwwBXZJTy5RoMSFE5KLG
mb1E7ZyQWWJKk4+h+xJVGZAGUJHaBEW7w+Awl0ZvCI3pXgMNvFhmZxt2TViHIFqc/QL5JvIqxUz/
kshT5uRljN7fUc5u6VvK9Puu6HTm5hQSkt/M1nMPXy/gxQGgjSZZvgevarFKldB9cwWGy8k7JorJ
PH7UGi+5xqXO5oPskZjZRS43xr4dxhf8z73SlDcsf19fLT4q6IQORcztd/W40odz847g27tolaYt
mXy9Kb5/NkUg5P6jLvnEAUEh1xAVj+9RwO3IvRbtDeR2hzt8fNkgT2pVCbzokIPcx0qd28oYblEw
mxJ+0oikD8IYYSDkSJnKH/GS2ibZl4mj4MeLNFpNfKNo67C6qvJ5UPWzV3CIKq2V7rpm69ZwkET9
SI4Oqfva/HnJGkvxWsRd9STN34CVGWtNvDiLFBea0+oa6SE6zvBbY3vo/cju57rD53yTN3wmYWLl
HgcDALaccCT8tf8WeZbeMybmxqHEksDD4qjc6TxFthYr1BT938xLXNZfZpszpq6OXgPAhhrS1bBO
ImaSDsMhlb6ojTjs7XppnmioJmXkGDJCbPk+BqgCbjPC3ensF1e9G3i/JrwZ5pFoqQML1117TsfR
5d/oqTLo3RmkBcrJpnW6Hoo7tWbplVuP8pAmFgJK8WOeF5mGx2FFe4TyEgVGuh/Kp/2JypvWH8cO
feekA8+w0+kZjdf+LwXVKljsahiAfVSjlU2wn0obEn+Am7h1WDNupurutbBuOTUB9wdTPG1DeGpl
HENWpk6wEevTkLJ44dPX8t5JADwg/EfZjCIzPX6Yj6/hHQezhDjJe/vYAL8/knA2xPi/wQROCsGH
obPMTgg9marFjHF2QVezbnnSbIxXIAhbkwgwxzghVXbkfpFD2no2I3b5xd3AxN+cM6AH0leAHM2h
HDOIn5lmmPnzB6YgBZgLSF64Eivl3jHzBCkboZ7PDzT1xXVg+eRyiVya2+241DWb/qp30+78OW0q
/QVKfvvHR5MH/wbLr4buTkPP/ykjHxdLThbSeILZdrfmTVcYA3Q8A57gV+3ronqhIUaKw6LQCMyM
qkhOqPuq8QeLsQXQx62Lda6NPszNmqZKSm+/U13FJFBdwhfHZt7H0b+zirxcu35UWiO9uVu1MdDe
F5yAVbvzPwIWOCBqEY7EIJPAU3Gx0DPd/P/qWWlSuyV0rylWlBdt8oKFlAipDovjVP1KqdvPvc8Q
fLoVnrAkLXEiVzhwYfCQtcW0BFG8Dd5Ad2EJw9n6EA5VAsIEyUAOX5VqJ9vEaeVrD71lC/Fbr+Fr
1ritrlGvWuQaeMBbaqPSpkTpwarlklzy5nf82ZNVp+QXBZrLAfi/UxhVIdlGt4iSlT0jbDgxB6mO
6KvjF1NA8PCY5IUEb6tuEi0lK+1gtnJ1kbxd/nbxe3zOZuwDOiQhvAfCqesRfFlM5R2ilc3HcjcE
aX2/hv157oKQ8tDtxBWPPH0bif1ex9mhXB3TzYPLgj6zCw3fCRgauNkqAlLVS6bjzHksb+I5943S
tyBvmDSp3PNoN+y0JEsdUOrH+mJx70Fgw1XBcdbt4FeqqRzdUWGyJEqUohrBFKrk+kL/0kojKdI1
693K2NoL+via/WXat/ErzbpEDul6sNyPWB/SmiksUjnTqe0hbD/Djzs7CTbuIBYn4SLi/rw9FfhU
ZqPLcAWqUKoJ0JJpnUVwF1oyLenUzW4lbrC8I44DFpbz2K3V0ql0MSsWp2ZbQ2INn56FuZpiSnUf
NM5i64d5s+c8QI6ldlvgA6/flkgTpmrx/gszgB3POGJtlWwQ96L2SgKl+Vidr78ijm1uPfDgsh+X
uqpxqXO+70CrZp1tlO5nmpbwE9hw9geO1W9Rg6mw7O164akEs/N52mBTBXEekc2KfR0IBFYLb/6U
p+5Tc896b+ChIF8Q65w5VG6h1RKZn9SzBN/LHNU7BIUzdspM4OjQD6bVZgeeYSHNULcT/39MgQQM
JefZvzXNszMk6XJ40KnbufJ04ezFkzVuWz0BSBcqDsVILA+jm/krz2q9KWHccITjfM4T/39DxYSy
vdQQBzbJs9s8ZxEyQvJCEt6Ebf5vhpXigmoPJ2AOdP2vR7LvM4rB9xpeYu9ItEOQjndp8+d1w2gc
bqvD6RLOlbnIm7xlXyjb0kdWod68thH+uZnmvWOcMGaX/SfglhDLfiq0JIGqjiElmwFTfFHPip2X
jCn8S6jhx391XS/QQpra0hGlRgtGMa63KRm+1ow8Qr0EfwYXxnxgmUrba5SxgaX9NGE6JB56Fe9F
R+CXs7uaUEsxJ0N10COMEiNYqm9CvXbeYVnIHa08fpodO55OCTjPqMD6iP2Isk7rURs5NVe4dCim
ltC2awgfuIKVDnKYrHYRrxYnqWJbKGP8wzI2IGNRAuMswTXCC5egBxGT5s8meiUGkWKjiAUZbimq
fLkR1Q9lGSLuU+r/FBYgwTsn3TAESjRvPz8xjIngA4ubYPRUvGeS15SRwFmzDXLSy2v5aMYF6fWj
LeVFocHVSiqeNzgedOUG1F7bdfPLW7tkFBfXAdzeF3f6XBwIcTmA55qjowz0YhnNXwFN6lttDRNL
I4aQzZ630mVq8DwIl4qhi6McIfPZ/vS83V5vP3omZ41cw3FMXu5L6U3zkXjDNwq9dSm0nJ2wEB3g
nw5MZCtMbWirebXcsTXLZqG7E2kNy0jw5XeYaaQP6ufWwy91rkjw5GnBdXofHQqH3Jwqs6qIX8Z4
4jyzBOR0DM9bL5bS3f+NQLnvfiFf3hjYImCdSfzurRVp5liuicB+CjHHVipiecgMqwNaKAfOnCuJ
Sw+GIou96yUazbcYRlb8O9Serny8ygfq9PQtA+Cp1j1diSZk9/t9/KxzGF+wLwn0VnmiFEoUrf7z
0KUQaNxZiPPd4LWUyNbv3kL+Esg88mALnnitTWWlhPpxLBTPjiRRM4gEOJvpzCJVevRzKUtwwM3R
Qw0koznzHaGnLM+cSCiwlS0oL+NVN4w0IzinWp9HPZOZ5e1oauEmHlUfxa1RRQAnNY3IE6SzTgeR
fp10tuyvLxbIhecDiGShyAc4fotn7yGO1YaFE1ohO9o57chc31IoI9bCY1HB+gHMfdAEQM58EQ/1
HVjuVZ1QqC6bWWJLEbbMzn26ymKOM5UlSd8IJNAJ7+zpvtbd0mOF0kJPuO7s1omWu6FBEHV8EIMm
Dvhkp1Ps75IQHTUptr3odWvYUIvYVloe5sKVGxUh2mZCgVWbJmeqF4M24UGxFpNri9A1w7b5gWe4
CeuphJimc2A474y2VZxvPM+Jg17f6S1MbNdJUFIUj5jkqtqcIL96E8qG442Mm+Qty4jWmNsykSjT
dP6u9nlQPLF/JpPrYtF+zcazzfGInb8xXSx3Lo4YogF+jw/m74NRRhwoT456KqOnh4v9ZmcWeBUY
jSKWGCA7YpfKC8a6aYdMy2fB39XRgDzIVcWLKJQlIT5oZs7LVd5JvIHBLOq1fHtx78QntSbCASG5
TXrQ8gUrA9Zd1BvDS9BXpp/7kE6e1xfKOXuiirqavFKNgyC5Td+6XLvyUTY0KExYgAxPwWzxE0CK
JctOn7nqJAs015i+SwCOS4+E+UexS+qqAVHVZ6ZsQHuY06aYIP/SUruu67D8P0ZPMBVxtvv6kDWk
k3FV9mfH384awqBwNoFshyoxQjOKTucMbuPXr3GQGdNELHEtIrav49F4PsjWJZ8yISViMKE+eoNQ
5xNfDZK/pA8igH+e0Dhis3fWN7tT2MpEtSBeu/q25kAPG4wYdCrQJwnfxnhOu5HW4ub2YkwxKWb9
hZhyn6+3XomZZerpi2U3K//rI4E4nI7BvG1XiGDHc2QyacFQy7Svo3SYrMEn6Xt49Np00b2K+/ID
cKilX0SmOd7yzBM9qRnrGl7ze2HM0RUuZKsI6RDGXn+F0d0XC1fkFORLX6rvv61OFEHkuj73/aFt
b2fkSHA3u2ZJcgANSA55zX9oiJhXpY9HFt4aS/sIgkk4xVegsfNLj8grD9l3s8H5leg45ZBDGIoZ
8EbHPoG6rV2hWy636quyoBa68w7TwpsjxE3RKPl5I8c6KO7OfAyNgXP8tiA4O+i0yOFuExv+lEuN
K/v0zLiU25x9VgeD0Itb5G6/K4janMJ/oCo0z0Novvr7kS3/sWhTsL84vxI1leHNOCJ8CQTsv/NX
t20XwrElCZ9C6WAVuky9fI26USkiW74o5iXrgABkt2C07I+ak5STdvdxv7nJog1sI//kT3CZqd2x
aNReo9ePJByyAukJqY2WIjRST3L+xF/0qDEbsgBrXGasq1TKJXbTx4uxLiDICRpPx86sW1a5V9+W
JhFBLB9flOr7n7UzrFx+86Sw/YpTfQPXRGaR7ZW1pWhcZokxu2kOCGRmbZSzsXnih7DFcxwu7e/C
8CUulHoyUDuYX0L4bfa+uXT5GG/syQwJjwyfLaiqX/BFKetmt8QXVcUEScWDNe0Gzg78yCrCXtuO
AKd8GKAi6OrCoEmWOQMDt8rrYFFgRiCQErY4x8aSMH0ackOzF1ZOnpcGwqIWT7z6Of3apc3mQqCy
HjJFjZoGatHmNhLp5JJqlaRUURyrDs0x/YQoas+07Kbr0363l9IbZvusfA4+vrcmqcHDhzDAmma4
Jq3wIYao6dk6EZXDWOeqRHecDAyrbc8L7ZfKZD4YM1rI/nip985cfAFKgNVfrQ5oFV4kAR3Le9r+
LwRPA6ivl2fGCLeSG4+1ZMEME8G0alV7Ikkz1gTCU2YQA92KHCs3re9cp3JtLHmlPrliOnzELVIN
69tWKykKupFC01Jaw0IttYmsopFrf2d4bJ9H9/G5aHpjeKLVT+x8K8PMyL5falTTTen0tW68oQiH
kJrfle0qJ1dwbvxTtReizuXQ8wsnSq9oPgsCq2JZyy2p6iEtWORtgcTi4K2NEx4ySGKnXlE4eZi9
5AtQx6MVWlWjMl3Cxt4GlnvAsxTZJdJqlGJaHVQo7E9qXO+5efQcfp+Q703H+DuPPcT/HzT1h0Cn
FxrUmZr9IQLHr/py+CmfXwM2rAcSeBTifywPNYIhKA/Z4doJ6FlZogRfOAZuQhOa9v7S97Y7rNvk
jf3i5txXbyQ0zo6t1VwlFL3grbWGyYKPUoN2uW9baIXZNUE8JbaJA3M6kXctxrHa62XzBHliy0JV
aNFP5FdbWyG46QsVoXT6wxdwJba/LxhPsPrM4bOnjMGAljbHp+6TldptsJr2eaFyLP4zZNcakj+M
g4yRKkqHo2v6iexkiiuzHTMQTEp5o878cfJdrC25X5XPHEzR9eDfXzZ/3mhQfD97IYiqIo/Qb2hU
4eYmhXVc0zHqKPoW/E+PhJOV28fZHmF7Z8/gT/Z5iwA0ucFOGOPeCCuB8kXhRfQSwrJHArfDKp7X
h3c5Wsys1U2YEraYq3r7JWBtTJ/HCoH+wWvEd/A18b+e7vNwsQZprpc04J2fwr4u0gO8FoAA+D4/
hH3DjY6Mlx0qv6x08Uo4zAvCz6VKMrV9rWOT3YwDwMm+1JkZNbc5pdVaA1Iz46u0msEkuzIWrH9k
XefYz/sJbMEloYVt29hnPVeXcg+6uhFqaerq/ABAx7ZA4eljHeeBJrhsqydjAcE0J+4LjKjm1eXQ
vruYYh3K6y+ChYXFMxWX9SPO3XYc5jrBnEZZo0wL1oualqmeWGwNdwQeJRAqJV26D6VraxRjR9zS
9xRRV7DXoiuaW7aLUHq31PdPdatl4eE059dRCCaleSae6wmnLvTMAI/9OS0fhy9YsTQQi+H0CyjZ
xz/isIyUvGrpWlJuYfpCMa84khGVMW5hyUIPVD3xd4AXYHy+UFC/E6nQCG2+aJi/X77cp1FbfPVA
s39X2KUi0IXH/L+EipxJc9O67YmasrYm7OAX7+Zyy/HIHtDuJMozjnUuvzCU1O/DKvpkP8+GbwIy
+52QSv5Rlox9rNIUaiavgNSetzwvMDKktGWv1PJtRXCRmUe9kYeZUmHZRMGaBMu8Mwj9hF6oydxq
cPmCQw62SAIRSMFf3AbivQdCPNHcTYgpUE2oZL7Vg+EzAnouSg0vqsEEywtFxCdzhyUtQn2wZkoG
dB7geaDtaWxoyFNHvrcHqMQ0xuqtPuTyl1S4ZUYqJgp3vHc6dlv3q8FeAAD/EokJ+6ViPYYoVClA
xtgSmTonOr8O/jdFwrGMtTs1EWfdEQXJbXclQGC1A+JOfGGhzxnSBCvGzMWCmnNBGSRJeOPU31Kw
V9XFR43uEAykFGDpWAkmx6q/SYR2+NeFw7FSBN35tNHGaKIRa3kQyWozrEwvwgZxOMJF/0NVG7FY
CgjnA2NTE9GeiQuNafzWpaIIBkWFg4xQu46U7Xtl58fBoKfZUAqZSBBU77UpQp+zNRveEnZkC1F2
SKGoeLTQhMFlhKG0rCd/K5JmRn/BQ1UKkbG3HzTADfyRzTWpT9eFX4PWcZGS+5zjelQtJ+U6wDs8
9lniK/lPXH/KWQEpzFjKwQVa4hZsEWpEvGGYrpJ93Tq8txMk36lf4vsXdVydbOH18IxVGEbsARxi
HOcroF/0nBX/1/SwucSvNlpl2EIlGQkjMFKwOvn7apEjXT8hwoiBZNH3MEWREBh9SAVRb6m1g9en
jOmPUqJ7lCbz99lNJXVz/OfiBzL1xWvSVzAFv+Vf//r0kRwDlw9gV3yBilS4JCgRo45PhqbWmLWq
YfuJ1MdF7r9ZFnSM/brtQ2dDchl1EDKwuT4k1G/cTRjvqPQq7eqd/vDuZLP5xIPpxdIRP+ZJjKDt
MUa733pEinnx/ptcv6kMEl7fuPPss3OldKz4xej/nkD4wFA7qssbWeOWxJ7Ou1xoQhdmECKXpvoE
ZaNiob8GspNdojeLGr26E2B/fbxmuSZumWJwsjAvi3h9uGDoTJS7v70jOzN5FWf/HiUHHgz/vUDU
AVHGdl6Ea0B/Z8VyFzEjzWfCOZMT7nPz/0mnRrT+5nTyVdNFgayq1FeUTGz76oZuwTM8UmJDYReS
k9RyRJOc3CjswpOCRsHtp8w53X25X/bD58233Xpjk/AwCuKwoM8qnLotLk7QEiuBlzLGi0C7wM3G
WSu78yudniFQK4iRAdybvF1WTF0hZIUwJcyPf8RkikWpYBIbvFXANhwfywzfoaYzRnlWxHIU57mX
Roa09w+3n4k3dHswFDJwQ2IG95CIWhVJD4wjJk0dXM9J0zuca2tzPQudifJlPCHF9E4qLlsnBZCA
dgsrw6ltaj7jMP3i+oTJeUnbDTzX97vh+5ABMJ8sLLwGEsVNGvY78Rv2a0NqAuQ+POdl0bsCTdes
MZMrirvoKeZnuRdHXL5WLp3GD2JgdgD5FJVrG4AUnn5KjSAH7sjOn5ETUraRc3PFBavfdy+UOwD3
Rk/T4wcOf2aE2G2RC7bEL5nYHcdgKrw6zy14e7+VcoY2VEBjP84akHoVQNa6yTAGzv05IF6pRBZu
SvtTwvTq/L2H46QYrNiV9qWxW+Tx6Fxo1DQvSCg81uTCMHYSQcpoiPLoWVTi8evCZP6Q1H7neEC7
GIkYcfIMWHRqSccydZPtm6OxEeMo5qaPlF5B7QbEuJQhZ6Kh+ikLlE5LF9VlpMByNwAsPqPlijfx
MbqN7MQRN+2jUgT6a4wuoIIAJe9baMeD8Q0wCZaL2+14cvqec1tf9kWU3SCdz8B3GdIAGSj5ZIj/
ZKlFWLBY3OhsCyHgp55/ajNTtmGeQvGanQ2oK5BNNOpzKlZ+NBX3/Rtzj9LujAh0NGiq4EnWOAp5
f5Tr5CCztjvl+Wxc34g+Y2cs47eNTdui5TixdHZZFUqk94lSsuzzlw8bHkTsSEEQh33lP/1IvzrB
uHFF0ACFVJViEnfocxKFgUksWkGPJzRccMDTN55YeSFk3FxX21SLT0WWpwCJ9zQlqSc2RLzb6oDV
Sea965u+vcxMTNjy+EuqYdDCY7QtwqQ4q32UollKFYX1hX2L4JNduASEGpehdtiNjNz9mZ9MSWuZ
+M5qzag772sXjRcHBDY2yjWYe2CPMGmfrpGl0l03CZstzrvzlS13LUvobAwg4V58vpZrcIhPkkk5
wBHCve+3wB8fqrSOxBm5aVAv1wxOhTpmh3RyLRvfMsJiQfw/gMJvB1KsdSSPTrRfCowEd2PyNTB0
0mPh2VQ+2vLj4VgkWzGF9bJYcUa4gEfVmtC1mOWJlndxrZLOHHem1Thj4zTiFRw4YSmEYWDC5wGY
qsR0otcJ2RHpkK8a79l0tBuCwNIuMFSDGz0IQLJvLvvdMVNd45cN5bSg9mw5F2cOLTqjnEH72U8t
KvN37/0Zi4TBeAHAouPyTkfdxLZ8GCxJjUuhRqFOPhCz2vrKbhMMUsMzM17hko+ccI9nYt/bHWLr
hF9D+Vl0MTONQ2kHsdMHhtVVcRUVKPPruKulDGFbMwaDVfGZoBoBbjQQ0n8hQq9j55n77znNurtP
yrVDPntU4UGIRCUnOfJ0jEH51Jak+p7jJE3NA0aoswRk6cPCiDMn0FJ5YJuiYsdXVlVXz3NI6zrm
QldmwsLPC/AaXouHg+drmw2QEpeNRqAwazIMmr36mktBqYpEGAsZkwsJIqOnT3HbUzSFmAq88nwp
GGdWTstoV+H98Rd09P66m4T4rn6ZFUhjNHtbYQRVRb2bF985ycg6mutglhQ/buokM9VaP//rj/LS
NhPSpnhEUF3OrTEwBHxotTRA2s6Y/Zj1xKZJ7QttTh9PDjbUXMn6sVdSI3twZKw5/Iju1+L1trF+
h/IXcIiOvjjhFgrd2kQ8X3sdGyQ04bqlEUZnaUrrREhDEMPKme8sFIWjA77VXbHp6avQXTge7wlY
bZygfSSqAf57gvj+NQSN/eEbI2E9mHhhfwqxertz7l4lmvyd7XtThfhw9GY3vF/wel5vnxbK0nUM
QwkBRI6AQdCmssjnN1E1hmVAz0hO/KniOEKDl0CBQfZgAp23K6BSAOwuBR+RnC1P9CR427KUCHGK
wOIi8Lbep7r3dNlhW/xjIXJB93BudlBxGturDveE8cTVNyp0XGyGxOQdv6dv1cwD5HuQMO/XAK/+
DwMu87kxDNte1FadFc9JgeewJXI2qfv3rC46vRrF6RdlyvQugxmN16YKhzzdwRQ5KkaOYru4Q56l
Q8Mj+r0UqmMB3h6PRRPdlWwjDBBWuvj7e9hgWVjSzgg8LrfT9yiIvnlHy0ThXsIosP92CQ9nmm3M
XaifSst2152G1WNW9Kt5kDaBLvVoaWQYi4Lc7CwmEJi3haVfzAd70KV+IdTCWMIymBYyVbTF105C
RiOL2GQYE9GqdnXSIHZwsTk9yPLeKmAtAD9DWuwuYwGC0zj2gUm5s7XJ5Hl3MnNJROdhHSBziFDZ
GfMSostHy7I3ew9GHEjoNGJdj3wKyhYGlwyV8ihJ5yeYyyuPSd2s305HvQ3mAHwLUn1n3Y2+O8Zn
PNVHIYDuQdkm8uKhiCufi4oHrNlG1TNMloEuwTi0B6Kh7ATnnhtSa/o0DqlD/Mal8N0m3ImqVHXJ
ZCcf2JP/HYK619eJ1A9gk38llgCtv53FRNuSVnFWH00TpbMKmmc9EczBINMLuD0tdSePiZpBix4y
8FF54IYbDPpClKs5p6tGnZ7iAOFcPf0Lk828SMjuAIzUT9aB5h0A1iJAafGzvJezq6NkrG37sgqj
eM8VuiVxccB0+nxmNBFIRqxBEaafsEbjSefNYyhPIiF6sr52Hse9993yKQh+5eIDZTzzZDXYhjeE
IF62kJzcaakfK4dINnEBJ6EbAa1eggjCq+UeIc4Odk7Yk+uQyxqx9FLF4BgL21SigAXO43d8l7Ch
5bguRvC5Zba0ctf4J1vPRG90wWvaHTl/uS3g32wxP0bBlAO+i1Ehtcukwki1xLbs0wQlDAreTI5l
JJYxCzQ5MC3RwYbiQ7nZVnvW7fxmROZNx4AL5LfkLKgJ2tvKp3XSQQEVm93f0w2FU+HvB/bFPsBO
xwkCP6AcNI3VLgTkdrdICy+QiUtg31wFSJr2frRhEn5twHCnuFMKMkZZNATn22tsBB8b+sB5qzhZ
aZM2TfgWvm9ML1y3mSPb/16AYDocw7mBHHPr+MpjE8fM5+OPO5KnpEzMBpK86Ld4qtMOqrVlw/Di
wP5qnk3zEA7YbS64+ezUPPBtbf7SrZsI50o9V1w3ViGiVd18Nq2uqpBuebKZBh8hQZXYbwROX8RE
K6z5kY668X4xAlaG9oKtHvlUuFKGanXEymxKoW6qxJHFW3aNAz07+PwxhkNkbHszOktfUWy+Gouj
/8Ub12O2Y3dkrQNy4pUWHQVmooqLFrOpJupNIj2AAoA+/dHcysNzJVepIRragS3CInMWdCnuVY6M
BFkjdxekgecgd2ORD4u85A8f6SMLI3rmtxc2ag3uS6rNURI3PaAtorex3gMMXGdFlRYEOFgsJxsy
/HcR4CXsnD4woio7LN9voEB9RrF0M0PSzJQaBQnS5YUnGXvL4JoQ1dBzZTkoob7gewz6D3TxzbpF
i2GPOfJgjZ9uu81q/bwd31q7z/a904zdQAyRsteB9MfmuXaLCbg2dLB1PHJ/m2a3SU+JFf0f4Mc2
9cQe45Oi5T95ZOiEiwB1JJnPhLJ2gUOICCbv7aZ4GJTZI+K0ynlLu8FlwYrU7q2BmnaGvixDYNCy
pwJR203oYETahRko1X3gqQHALhv4lK3TJRfylX5mhSC4NNC0GdEsk9Mne+82zyNXYB+0c8lyNYF8
FW9lFX5enTdMS2Jnju+KogszD1vPUu+yD4OwbZQ4jlhC9+13RP0Q5F3ABgczxH1KNxCQzkZ3Jkoi
+WfVHKQUK4Y61ZyW54rLqZ4WvVpvR1mAMilT2XnmBVGn4IDefa6A19RAr5IAzsQIw8ffeIoySfz7
0HXk7dXoJU/WJNuiVWuu00+ELgydYnvGWQFriW/4An6aV1317+obAvwM9OnBMufqDoixAxaG30lL
C5r31xLTTQdU/8sFp9WBOsMKqWlrxiGjJ4b02+EErFyxHtsROEQCU1e8jw6i1UZjTX/saGxcIwUA
rjtZlFl1805rutLOksMibyPm/BKAi0Qx/MOsmgfI1JnRuWbr0qIK9ThtWgPuaNYn9ZscqysiWiQ7
AmbsTa1V0V8DjOz820a2VTjcCwfVJdQXycq+OLc+bQ8VKyCX3zHV0lAdR6wSu28FHkVXbFQ1X6dS
YKGpetspTko9MkjUvVZOVkk14XMBfdk8zLLU13P76TZ1mXCKNLH21X1LByP+VC6a94dxWr0IgaB+
Y8zuj73TPvmg/Bku03IYvDUSEHHJkbMR8kr6wR24PMb+FmfTfctEuLi0vpeR/9nqHxc4mYhklcsI
K7O2TU09IaZnmmG+XT77ebJ3FcsTbFRgKybpRpl1S4f3wdiNZzLqM9pJJUuIqoqRMnU7A2TJ/Olv
+W4+iHskj+gChxZPJuTMHIOfD2NR7tx5fhbRNi16mYKauA2iGgBHBDaAnVDXBc8l5P49gFzvrJ17
aBAxbxcbIDA2M4JRZapzs9VRK6hNPundMnV6vIdykLwTjqnqALnFUsmkhCtdJprgf9SzgxONVuBz
wy5aQ+Gjrr+sUK7OiGDtwUoRlKoKE15J3atFefWrFXcpcw+eWV8EpP1WJUsQ6mMePKdcnJlX33a9
v7vdFQX5ZsHKW0vQAPyUtodYAECmFA8bJ4JB1/ntzv+znUiYb6hoShdMEkqy4jMGSvyjL1PV0U7u
RxS5KAHIqTin7/boRE2wrzDgXTPpTm5qa545BAc+g7duORY/1UPh+QgwuuaXmThFHbMJsEoCf9aG
ETbremNcZOff1ZsOGMBgAxTCLYVXvbb0qYT1+a61Rqj9VXt7lb26Z5FIkCR0U2F2BfYp7Mowpse/
vR9EL5cWrcdmgDFWgQkErLQBMGyGJwHUgiKa4keK7CO7VjFmHFxCPqT+LmfbcwLmi7YcRo6ATVw6
8RK6uenWhtZKneNiVQeq4EtRsxhLQs45zE3/kI6SxJ8dAppqBxG8/a0zQ+yey1ws3aBQST1svBv1
qvOxSpS/w6EWIhjHI+zJ9OgjxAfT3alSzoQPvfZ6xNRxt8xyHQVXrLes7qoTCp8go9UTvMA18nOQ
axtw2ZkggsxZ1h7TNzIcP+Mz3UdPnt/iXpEgQFffS/UzXT5MmwgL7awFtwDktNAHi/feiqNhEZS3
HKZzDgUp+vwT77Ckr0W3wDWh+Jy9jRjn4mNJhaFNXKWFr16EFBCtDHwdX1SE17qkWU6Gt4c702CH
WerWZvrrQYRW+QtaTHVGz63tJZRuIsw97O6bBjh46r8pz8+gmywdEYmGmt0SEX4FaK02Enh61pUo
yWVsjEX8eCm75GA2y07WWDaIozRtJuvaeL1qcl861ATeAnLS9ayKwrAQ/8bbKxosdZE8WZ8s7BJq
Kd1XRU6cadCuihBIvkwAf7DAeDcpnbGKklgKOu1EhpDqrtjJTq6JnL/cx1w+pdAzACGCYqrIdRt+
lIDVuXV5za38XUkk5Ncf3koN5Tl3ScPvHnLCKKQfuFmi2HsxaPKTCePuvmZsVPiXZ6vO228X38ts
grUT6MMu5jdJeGm6ikPa4uUPQSvD1dBi70LOqejBopFopcGhCvMSspjjKVbofro2LHGWhq7q1uJI
FMEhNNaAYAco1SvI902PAzgjmZPfvBsA/WWa1iVmuIzU6MQM41OQqpFlfKxfHPrKUFSp2KiudLk2
0VUUtyQ5gnS6sCobDfhNKrqXW9EzvxLGmsskUKkI1bN5q5mWUe/HZWYEDQaBujbUPXijEgKfOND2
Qt4vLpHelLCnJ6P5Ik4LFJ3T1ANK1ZhFDFvfNNX8OigPDQBFkhqwvCrJw4Jw2Z5zTOdsAb80jBd7
gII35LAsOr7IJmM3xT9Jk1Ut9qPGu84ZgGQIqznLiTXVuWCztxsXihGkkhz+5lUzlOlFd6Vz01E4
oXLufvdrp2WkegtlCZZ1QnhPaiGhCv5IQ8+mrUsKMsTn/WjzxFvIomRUr1PLjC/nKWPRSWOhupZZ
eRQNGMsYkbldBQLLwO6rHybLNAUxAcDumqAtwcUOAZu9kkHRoiArrrTUNREZJqPN4SOFgLLKuAaH
vlMEVBCrUNNpdxZeI4wGCKfWbDHDo7iDiyPjp0o1cK0i2SkiH5xcH5PfBUPfL9D2il8z1hj66l2G
2fD4xufgVzTqAgZqQD3WUvS3vZJj37F7zt7ZVwV5JxlmzQbJW4Gkf/TmjVOKKEHdyRimgCuikBlh
c9CB7omEjeau/KhSU9cRC3G6A1TzVwgRKZkhaFqp/qkJS7NfrlwSn8TjTn2aDvGicxATk4tsgh+u
2nmsg6Kc7T52okLHnxODhv2er+Ud7U2IjYzX/s1eNTJpbR2lzzX9IWNA0tmN+i+e98JnVhzKZcnR
057cQy9tBNL1f2L9debQLbiguOO9Cv++QqGQnytayKRx4I5ALWgvc65yHf54wOHqiR6yWxPqM1w2
wxTXtEpUFXZiiT8xnVdjBL19fUoEaOBO1iiIaZMomQdaJ/Uk3gtJZp+CQt7YUH/672YyAT8sb/07
K2eyMNps/41z/1c+2eyOeqIGtyg7l4eN41hC9RA/JqnPRURGvDkxBQpweCa2ZEJYlqda8IRF3LLc
jZpcqaSv6Y19eov4giHEH7mNZ4OYvMdExLGzYAGvzGY7d9zY+wmtOHcZ2bOBcfZZ0Suxdw4xu2ab
SsOYScCFt5O1fguWrjbFuF5XP3mTnOtHpKI2eZLo23KEnq0LRgpRFtKXFvAqoiWb7xWE9TF609Al
W1zTxJoH8Asm1WgEJHss3xi9HwLbkliFA79Y+gWIlw5eRoKxWfWtxUAKIj7/xNd9ndVgt3LXeyGp
SYL0xeV9csit6ZMap7gL36XR9P8gEcV78msaNfSyp2mfPZJ3RJiV0gttYp6qwPlFDLs+/A1wNFla
/0PSI5gfENGegdzZaqQxgAYxEBp49HBXg4gKIZNmXTt/OuHj7UcSSI2RJbr1WvX/D+5Hkv/Qf3wx
Q3WuoIVVD9UiWO5hg7n88ASvyXuQe+y/x8BDEJn80b8jUTGv43OV/5wLHze22q9hAp+RmsR7kDZ1
tpWz08hgLlSbZ3nl3xCGAhs5ohB1WlCMGehPs5eUEmSemfCtByB8iGCRjsgsUX69YM7OmrmIUVQG
pTxF6AlZPRcf+ljL0bQnu+BcBkNg16Mv6NAbuV2NS/eqvbdPQ9hEGra7fln13iEK1OSCE7KgzYjS
xf/OWouKV0iPoVQ01q65tnRz8eTyzZFMsJlpdoF0vbOqcElIYYVhg7uQDNmeSF6gzjVKWrDiFqTm
tXnZBvLnSkU/BhrPjlEJjeNMGCrEgFJKBvmPlxRY3XRjEn0KarjBo2zvloh6BxxxCDAr9kYms3h3
/1HLdeAebnh3FGUnyZ16l2S7JSrlTrck6jtVHyjDPcTxtwK/RxHouIDxebPmbwTBQnMKs+dT3OID
Mn/9hi6UedPvVcbeAIwsqVP+2SAq2bAY9rH+srCtwhz9ANBVyd8H0i2J2LBLp5nWiQT7Y3evviyW
WQXKPym3NxWYu934iwmeXg2exmc3/BFweN7UdoPbb1U3wvYzBxN3leTzo5CI3FAypby3iudpP1dQ
518hu5YI7YLt7nvhd7o6CcMsW7UScvaeciHU6k43uICD//FtwsdMM4MtuyfjpZmieq74SFu5vI2M
WgAJVNr/QxmuBe+KmaNQD/0Ihi1x3ZYo9qMb7ldEJzgIgGq/fgjlFEbtMQZBAHDF70Pke2CCyOfH
5FZGjh1wcI/+yTZ0SoD5/lOLp4kZdg0r3j7dBNme2ghF6qWpjYtUW1mRPOSxP6uh3dNmyLp1m8zI
AQKckkr1oArDaWQIC4RNpT0Xz1W8QYZWEUz2ZoV+E0tF9QHNvb6Qnt/Kmm2k82J/DEL/HlWCI5dy
x4DVvXS5dvSXpPsdpctZXBWV2AX6eHZ4Yh8BEblDM5UWk+jZc+2KfhN0dQWHpGPLUYhkSWqemsXl
GhH6RVrmRy1+QWWpE5XqY38LGjmBlPl3X0V1RQAWuxA36cTNX0tvR8SkaaD0QxGR8ZuW9z4+4d0F
Ij+qneDX8GVlOXsKU5r59VFKpDSuGi1LK6jMzOIf+NmtGY2GSk5hG03aVbcJhsk64v8sMhpTkeSO
G+Pio2MtA8T9sMbiMp5SDiiAre1T08c3Qo9ZW8bs8xPFIvzhR30A97sTUPnlO2DRjgzrzSDYBR3H
YFitCvhA8X3ab+ghkJ8NIk02c9IeMG4qsZtirPAPkvuGdET+u45JQQpEfR/unhLJuQb4ECtAzPff
BlXpAId9Q5+ZsVYCj7Ml42RwxmEPyMfZjHPQshOhMLzwbFFWLwT/sK7fpNP8YfFTXuJUbFjCWfKs
raUPhv0qB6TlOTnC8t25lRxeRnJakK20wQVSXKiAzgjQXGaSD6SREZgn6yyQlbI3DtLOZdkY/Im/
e+rLapVkFz6DOYSrn5Ythu0Qw97LLq5xMlSD1FT9Gq6lpLWsE8Pv/76OhGgWhyvCW3C2xnmxC7Gk
uFBhfi3E8MrKUZvVLCmnxoXl3G96sXzffaIvc0G8MkxKCLqQkRoCi6ESUdWCwMEACJMuZ+vbLyld
VHb+9w1jGkACBkvzUn/Cyeq1VnbEt5EG9F7ANRz7Q7T7Owal6PlwyjAyHbWIWB1L4qiCOvfnb/NT
BV889XG0pejxVopsr8IWJ+yzXm/MuuDVGwQ7xM52VHaYNZnBVFkY5qLanqmISjNVwh+hFcNbcEEN
Ku0yYmQN8XaEqo1e3wEVu2LDm2cdkdj9Sfy1bg/zhspCUSsAjEqGptemzD44fSHbPdbP/Z3xti/m
BRTRUCMEudFBujoyRAKNW38zXDSwsObTGP28ve+0etbwxn+kHM2RsDlAkIE7X8ybBip3Pt9bvKQU
8Ckv8FJz7SsLbKPB/3lNVFroAZpo2rxWn6yXaPLxECpmLvZyGDiXoKJ7ygIT333DaKlGxWWCNG/z
wFbNNkHJYyvf7gw2DS91OcnpOgX5Nq+lxLRCfxwaxEIboOqqMPIaCyHA1R1xjLEEEddhGraqseDb
6NA+BzG4HoeOocZ8prQG/Qc0Sypk672H8s0BORjfYm33fWKbJOnAgEuXWqLcgOEeQaAy8DvNI7QY
pzrTbo+2dyTPyCodDuEyqmxR+3xUbC/HcD/w0/XtDvMfQbccGVLpCg83G0CjLUwMEls2XIYVkeJc
tNFF+lMukKKOQXJBxOWH5ycJ+4JWKy7d2d24mmI8Mfss9cvjlh4uztcln4GX79eaZ0QXCaCpDzTH
wQ7J/y0jMyIx5ueFSgWpGmyy6YYGNM58scDGvYQJdlfQoY6nfvQU0ge1BUL8BzWo9EM8zuPjDUj+
31E7ZBDl5slQ6wuKXZUhmkhxsq4X8ACJyM3y2Kt/PPOfzaRMrld3t+Huf50M1eJqx4j1yXwDC8Tv
84o+nllMN/ZOuVU5EQRqR1J0/Nkn7qWwJCge0Z2xnOx/3HgNzJpCG/7ZuG2nceIQDG/TJBhABnIg
jOHt1YsIghiZ98KmQKPiapQc7r9RXljTKdiae1Gu4y+Xo81Ihw0vPMMDY5bJiHirFeZr3yUyUDzA
QC5RYK8qSgHz9czgvxo0CFfjuEUEnFj/0jjVCXwkYHULioy+bSyOfM+fnrR95pKBgZ1/88MDmVAw
4A87z8aSVBTTiml5baoEr7FVYRbgxLgfyqogRO5detG2d0aOaov/OFZwOENKAxtCeKd6o3HRUtTL
9fU7/FzXinbu71/YnQYWwrv6TahRvudy8LxgVWKAiz62uqgjKxkJsEkxzPE9vIWdQivwnVBYVjoE
T3dKKF2i+2nQm97qldvf5qkei6RQJU28mFEb9ME78uVngJM9eJ98N1KWzgqhLav1M4Kgu/SBPBgi
Amb3Tlz/YfrryR7Le6BPMnoMriVPPE0etRYFDPfNmWqPm/oc4yA8QkA9YyX+0+00hrz3QBo8+4VT
xTgRPSW4ReC8P9sa033d6PhVknUPiHbBYvl+XYeX3Ubwwtd7qlc17MMP938zw78M6QXBePUCFuwu
RrWiwusLDzwxngEUwcC3apBYT5jVIntsTspXfowCaRf6uFi0w3jag0/POd7x+Alo6YaZnFf5YC+C
+iXzg0oy1WVm76I+6ZrkLvajSvMZulXWW1cmCLGZ1ZSq/fiigk6jTfNZ2Dyh3nvALBBhlTr5fyUY
DFvy/7/mrUHHMkVAZ1jbgP89WH+8E0+5HU8dSuV8x4SrbYHhpb64RxIfjX0wp7s+yx07m56T9iJr
sGTNs4a+dmflj5lyOVEnFYFwWbu3YHx9Xlhy/bYZlzn1HdExliUz0g81ed3cv2hTTNa5rSloR5G7
D3cFFzpw6WQiUF3CT57B4VPinbxhCmoCVzh7lOuNP7lJFiU8muLLTX56pxbixJ8ivKgBYHI0DQ47
5HFBdpAmyvWqfUKCOhbnNMaJF1kT3TRj8HvnYbhg0SUoMjbL/HkcARXlBn+Vw3Bp2b/3Ni2z+XyU
osnfN+oG/ddTbzTcIqWdJEVedPOnoAZ5NR15oZq0GCECeR9BycypczZ0IhKV05ivaeGHU3QsQi8l
PD3xCz3KM6KSxFcAjNFZZNlFvR2g0iSJvQnCpRjogFrEftp67GubWNvtLZqq2N6w/+/mYYpumjOi
dNP0IR/fkSqhdOwk32e5GcSA1N7IGWiTp2Jtv4/xuO3MLyX0o6ybzyWEQLK5h0aKMc61sBSAGzAp
FNy+sOLtY4LcTuWIA+qZSgTL7rtHeVQyIkYY8B4kbyA/lIdx53R6I2g/+9EbTptz1uU7As1bfvPe
fYVxToAQRsojJ7SCbVj+vY8vBS9FAMeWdF2nK3ZSVCsAfIBEOhBwhQ5rrvDbISPOQCL1b7vPg3fX
AD6pDLWwcLDYhuEoVmwYFtJAnCpcWM0+elWI0Df26EgvI8rkSkASMjUOGbMOZaQDIwPl5icnomDC
idstP/1qz8dWYJdxSTzst2cwVUpDfM0dtsNVqJFclecpWo1KUOI7o7pgWgwroIoXRRhBxFaRmQub
NFLRKTVmAfRDuqQUZO8D6ZtJSkIdp53Q11JYCLjjLNNtIjkgDjHN76PcdrtVIeZe7KbtKuB40Bnd
GWGv7kkFPfnuFPry7QGCt0DO5uxN5ln03adJCzHhwWY6m++ijFMjFk0PyI97azkEis7HW0P7nuhv
V7V6E6o2PV7qrtmJEhmB4vFoFUMreMcmZE7M00i9Cu7ON6QdavaOMfo1/5mtzAK9pbkx2IpIPU65
FZbl9T5qjDrz01Spjo/moeTHGoq2cHpz2X5wCWr1iKygs1LSiJIuYVh48aARcArUt8oEL/LfqyNJ
OIUpVOzPcp5XxIubTwFacYciKEYlRtFIqTvmq0RcWcF/Tiin7V+0C+IDnddHcCzITPwy371fWnvx
0IgMQYZuffJP+R7HQtvf9W0ijS60KybRFn3A6N3rQCT50/6w0rCcbilktqHPe9TMObKZwaolTLKS
J8EyYuoYWRewwfP3PkcDGIlitCLC9x1Qwh3eaB+zEm2czkAeyles1t75o2ynIn4hReo2Ie49S07E
EMrjD4y0P8IHasLGeqNuoUZAXuB4PRWz1zSH6tLiKfc4bdq88cYauelHcia01RW5Yo0TxNwtJHtN
12znoZ8nBeswQEpwry7BnRTNDvV0r6pe41mFrKZhFybpowCv5AAMt8BxO/hvJcuBPrY1x5leVaB7
iCv9C0Pvh0VFN3wsnqahDTRc/hRQ8J45fJ3i7ewOBFyzhUwwhx2SczuBgvsC58btrHkcv6VMm9E7
/iudueMXhF8LjYwb3I/g20TSrI7xwhDbU6+dOQ2ozsRX2LGa3yxvKavdYeq5FIoiYUc/JPr1WPxp
j/1sRf4S4i2lUdIgm2m6tMackk2QgWgLpxbQutV/vmDehmqNUl+uEKCP9+7uNyPxfMY2nXHXcSHm
Yq1XigmycGKLyCl4AsFQ65awV/gAr/km0JRRHT9YiSTPYIoazWEQIsKFFF38ftPGYfB4ehCeQmGo
fPONUK2iSoYFaZZVuThKuGmMrCF9y3w8F7WUQ3EhVOwQh2j5La/e80bP/cUbMSoSxzKqe/SOELsV
FxnAOg1yZA8WzKMD2jOTiHLqeC7jkVlYD4Cjyo2Wjt4fqQxCW0mVqGypAdNtGHO35kKu1IW7JNt4
kOJ/KX6+A54JmpF0Mx4BOkaWSoIuAZb0mDhbogNOuVwQX+4qTbjMjaQB72ULZMGGwmG3deLqZslz
hcNBMFya9+V3gN/6J2topyGJEMchGtO4wWHsf9t3WswFlzWRDHyaBKsekPEhgAbIMHvPSP/ufUK4
XYFoAJqHFbd793vNyyKQt9eYH4JKGFFSMBzf2sMgTcYGM9IneJDYd6/uhaGSJX2r0w++GNxhhEd3
QHIhCIjXijMsR73wfrfVcGFnN35XA2kwPeVZtpl1qL3du62jPmqtCVuvCHNcaXAkFZoEuQhgV/0o
gAQamEGmQO7CIocHR9gEw/fue0IRnBPRklbWJfybVWkxi03CN8zbkn93BGkd03nYaxnUZOarTgLr
b3xbfTdBXsRrRLmDc7A4nyU7KSNO842fOh2Hic4v9L8czTIJkxvSvd8AWYjVKcw0m+LSIHD1PFHC
SqDG/svXoPxa345NytXXRlCfLra2CsdMfnxDdATHHeafD6xfmQ3OGOpMoSbfb+zr5rCq2b6uwcKT
cmbACLAzWsNZAhzvH7kFnd3tTaCoDRPwQ5SUUgLAh7Bk3aSRWlJV92qjfW3rK2YuxVeybYPzKVjc
rNqPAq6ehyYtCmXY9Qi+ViIx24ESoO7uI4frO7s9/NRUU7ijzIvWufU66+LnXMV+o6Hr4X5kZFpt
KH1zZ7SgXrI46H/b7Dn5fznF8IcUb9smlS8CLjTYXKQttZghaaGGLCMXe5ADWwIVc/VzMoJWhs9U
2+p2pGvbCsUgs6ICNZc1rFFS0pdzZQZLdMo770waO7inRQWtDVje1RPPMQcjeJqgzs09R6lXBre2
6jN0fIhlQ4kfa9NuNsN+BhvvGUmhEHWptjPVnaHxS1X6M3XR+ekNG/ibVIsix06sQ2iWh1VR+tXd
+zw8FB/xM3XobR8QqdnYgGeffZ3f2z5Ev41EV6G2LIMEdurjFYkWzQVSd/CWjP+ixEgLp8C+JhRj
QWpwru7pZC/ftCdzl/SVPELd1JBENThcF8f6CZFWNI2lOAGuhGDlWvo9pjLUV//ozVjdkzIo5J1U
qUPgaHPrCFUGqVl+IlJtyYc+hob3iHNyY4XoXLHg+AyAYgysUaHvCm9v0Q+0ie5bv7VotemZ/s8Q
CV8shYYpijAatKObB355Z4y54YjUFV4g5oV5RddvUzoEiGp1Hi6/XnyLrEqAXypQzFj51q7l9MUd
5ioiPGYS8wOszBagsqxrScncVCxqX8XPEsks1NsbUF57FNaizSka7bHToYyxePfqyVmNmi75EXpc
IDDApeqdy9+H5lp7xu/sFKG0p9l1Lz0XHZejj2Bd8DaWtMsns3TQPvKmhIkx9BMPa0R5VH7U1c+r
f2l7r883G95rgTO5/oWGYW2riLBpsceFWSDGmkYCGMa/0aj3FSM1Xmq7iDYgHHTEUb0W97iiE4c0
SKayN8cTlzv+HldWxm8/EPXyiot1Ym3kF/GT9nJ7tWtIBjEOYlSwFpGrTslI8ZoTEl/de1+mYroa
A4ddZdHmUL1R2MUlM8J9RR6axj8cron0vnDLgWoYssth4VMwrSrH8UpZV3EuO1fdYkOmGQXwjIy4
VVoqRGGXFS3acO79iVU8OrkPi4q2b/dWoUBJiShfgCoYbT4x68Oledmp3HZkQhZPLn+5lC9qUIU6
ijEjlzpnXLJ+WkpicOsXinIw27pgCiA3SCdLOf19OZRgqQfZc2CVWtrvE2XugiUqW0p/78n5KDov
BNuC9PrEOLTx4Q7tX+H/4dw0NwNMMz9hzmig34a2AX7SvtujPGiN09qzmvbECn+OjalFwKOvqnht
kVX/F0k61HCLFpuEe+5+wwmWwQHB0jmnAijnnPuudTlF1BFIck6a++HmnVx5+QSSKOmxHKMQv0ed
NIc0TZGPhJYCbT/UlOJ4TCCaz6lHg+wkAIIdVzbq2lk/Z2Sy4+oozxfZtBZhpnhyn1omyAAfRu5A
dwjcWc2UAS3XiPpJbUB4jGM612dfpgzzdBYC6DSA5nX4pDlGh2HIycb5td/Uti7X2xM29JDjdOF0
7/THsiyJqvec4KZm5syxITt/pyrDtCjiKwAGdJ08+6DWTndZi+9ynDrEPafwVb97onNS7uzGSXmw
JmmhEdxL8zQK30ABky4bfJmHUqWvY7KUkM4MNp3TB7vhvDmJ5CU3D9HdkCgVanh8NZvx1r2ROI4t
onCBpQRD4TRJTPsvbSHr1DEAIaoLdm9NvQS2Lj0OXrx0tXbXvpx3j7SiyFLT6CGNLwWNVISE2fTA
/0p+BCXKuNH+I7tWxUVt489uUSzSNkgbBoB5vAo3eECZ4NtqC8HOI7YHvtalAvTTkdpaFi0TOMEZ
hB5WKTW7q1I6lNukCXib8A+fHTJAl30ytcAWb7Ex38jCBCsZCVS2kXGVUxSe/mpV1tvtNL0sUMd7
Hk4Fq8QQJJTIylPOIkwpbHpjyRF7eIbotR7B+AYvVpeBNuKq9tk1yIvltkSsCODJ1Udnk99bCYTj
mmHFgUwffcqibEbhLH6pJEpljWtX3Ccs3CKnMFI1qnbHQPjeXC7ymWZ5ni9mvgWypu66tlDeOY6r
F8M6AINNJh5N7pSrGYTC9V95TKOq+7H6KbfvKtYw6/xh14a0tzCpwtFbSlYoixDZzgJrll2pkH6g
nn8zM/Pl42jibLiSyu7EU9DjY4DNSsvY1I8FUvWIfvpAyBAO/mRtFtPWuxXLYDgWYyfWwzsQIFi5
BVzSSZgrXLWuwSkIPUrACS8naKKAXS2nqRp+nz/4B6I8MMuEJMgSw4cDQCj9W9zLxB8q8RO/eFwM
jnfJFZ3vqwN+qEYnw78G5/l1yYpaymWzuz3qAdhrY7p5W4bjmSsETh1Qt/VkdeWhiTn5SmmC1C81
e9179V+q0mqJvLqwa3Ncuv4SRyMhZsTVn5ECnez3M6eYQR8JAOxvgh53l/YageRe4hUUgoNBP+tY
XqGDCSNVhQLt58R5DxjDo7vzY+a1v0j1Lvzr+modhzAlUKkn9buDXOSPKpD1uVIMQB4pA7TmdjTC
+TOgEIebexK+BDeV0JuTcOol34d0W0hGN8n4iyljYvOm7CSpxr6GAls6j6y16Y/fUtX6o2iighrT
YvkkdJ+gAxknxgLN4Jb8ofTKqlLN+uipCPoXrBgL5FSh0CP/HY/ftFvLR4hzpX5zPcJAw2U4IP/l
cXh2d8or16GSwPqVPgMZf9MsZ3QJV4j5zJOxTx9X7jXn+JsI3MFGzjbB1UplM7nCagKmoEGO0nIU
9IlE3VN1kojTcCozPodgu36ZtPClMwt/C/6qPTqWc7lCi+GMs4+tMGdhJo97u/iX3QwZmMH12C8K
MIBw8CRPatkRncBOW0LSsYjFglkO1udVCJ0udhVTirBnKKDZIzHM6ssvzjki6wkCWuSwhTaE1WMU
ncTRS9RjnUQ+/SJQMFVt/bJd1ptICmd5UFjFWiKunxBx7tE1wR94e/w76rHbMyNmNp7F7HB9GXmx
YzA6ZcRhSQgJ7CRQn0LeZpwuvVtKnfB9MwDHTQpLIJlsMV8dNh2WLoCuhUrM2tyIEqiE4qVo4Bqc
Z+7uCZWoRDwict2fn/FAsfFFqzL9ZzBGiShGItDw1Pfpydf5rQBmBWtYY89cQsjKnwJA/DuXI2Nj
oRi7tvtMUF6tvyvmDApc/SUwStf+VKX9YJA2KdoFruOaPkw+K0D7NkiZto0aU3ZjFguWZvWDOfht
HC8m05KjmY8j4k66YXhikBL9VRDPHTJlFLj7scLrnmcch6wyleYfn/BOGCBMKG80hjF1PE9lVnLt
CEW6j/PaXKis2GgOOyh+zfrjFlp7Hd1+DxUxRzFviL6pkkz6JeTUvnVG+UyFxON1VI6xUBsjGL5m
ixjqQ227hhXAtf5I8r//uNisDDBcNrkok8emV7dlsBxjeFaiSBFsriup8qGaN6bFPjzoJYjynEFE
9zdqlfdilCcT6T9KdO1xbFWLaMniAdCAjhprdkq59riFzWbD2dNhCL/ECcdYm24M/AMbqBVyr4m8
4ektakyZ29B5T/BQn19OR7LyDAMy8EWSWjaxR0ngxsX2E5S2BaM6GozNTVUhb9aG4wH6BFpSng2n
obPQ85CaR+AAyiE1lyJ2dSmT5tn5LA/aFrJ6EeOs7txaACqGFQn/nKJP8bTYZlQVDSehWjrOXBXT
dO0KCkyfJrsVScIEVsCLoR36yIWoYru/ZXol2SFUP8TceatYneLDiN+ivo/En9MNsLlp9SWhTOy4
3+m2upzaAtXtXEcrQtG8MneJPqr4J3qPPQcrQJuvQ/8DX18wIeVC3tDzX0c7hSH1g6yXjcRfJSR1
XEJzjUWmydoNQExXRHWi8EhnyZMG4vkypWPXmHc1ps9l6H6NIUbMJ/DHgbPq/Sw2sS8vHwLZK0Mc
k2iV6RRT2hVPMWY00gajRWv34zI+MrzNup9To6w5YbhM3yMAecews66eLGKvXDPqf7Bw6vzvbAeh
hiAefneAm8GltBa6VxQhGFAByrsXLpQRNi82Ps/zMlDsiwtQVZPaghkMxFBHaGSUsiIbdBJTTE/e
p2H3DB2n8g78oqrXzfcc43M6e8j9cCXehAHJClMo4D3G/xeOk/jS1F9HcCC9d8GRYKsFlKp+Vmup
vFqnpAto1iKIPu4vF9QkGNuFOJjoGg1KeEvsbnXrYJQ2TP24az26f5o7r8ggqTU6TD8IYbbKaDTV
vmNov2b3koKO1tcfmxf66mmgtwSKDWu3i/0+Xg5A49+hs7o1g57MvN11g5j9wHUaHi+CDUQisiqA
VRVavf1ViV9WMa9CJ1seoKinWFWQPxVsz2xydUyE8KExvXEMzI3454u+axbqQKT6AYFw+0aYXj4c
lhpvKRvaAIEuOT/zSZxLu5+iCBJ6585xim/Bic7d0gGIyeoMzwizMzjiAs7+kxd9oRiTwXwOJRno
A10LFtaENUV/I1noAJErabdHepzSWcWvKBcfWdttNBvSffH/p5CyqKg9EBvyhZt53mVcYrhgXk04
liPGO7vwBl/wiibqvKDQ8iOO2lv6SKSh6+7ZMbEPnnju3ihJQkde6lXcDgx179GsGHgwKFeKUzwh
enAySOGc0f2BTyIWvdSU4ABNwtS/pKDkhYIpOnDE2a8OUDW8fNKW5kNMtgpMXowo8c4MI44crEtZ
w1O5vwH1A8qxZHj7tTPCvWeSMOnTW0StJnkAQg8t4liU/Km8HtcOZh8aq8+pK830+T5kDuJdoArr
WQSCJxMI1di15xPLBRFBNtAEgHyuX+kXEzYU61U8L9bJSI7WaBQprIs0Ooqd9kXawvw0z/AveUno
nWftJRNK0gDx0HOEdrpo5VKe/lMW6AfbCPDO2+QHUPz8hPrxrBgf+hK0EdtMn3wEekDRb+fjqQSq
e1JBCN8WS2jXDqkQpKbi1xkgADkwUFi4WL1Pi7EcttiwRXn7NugC1m/dLUHFyzPnIV7bc9UrcKwK
SnHQsQrkdSh4PDfWFuMkeyX8QiU63JyaTE/jeayvxeKIqjQZCAVST+D24a2Om7EB6H59xYSDi2Q2
Zl408ocIWueWXi3VWTwToaBgo1B2fcEmIeqwemFaesiSQj38nOfIoyj1LOuZufuHQEi1f2rRQ6kY
E2o2Mt6PMb613UbuS/ezXKQbwyCE1wrDhdPUT1bCKNw6H4mTol6MwQdfwqvvO/amDprwRdRWxS2F
pYbtXiVYSFWOZ5MnPSp2LASOZy/o1wkf04gjNoPJc+c1pzQ0FfsfMktiP505BHK/QjhnaYNSlEOl
EkVOjuVkhiXkKX9t07b69Fyg3WLHL9LgwRG1sDWmJpU2EQO6qODU/+/2Ugxs3ezZ+m87Sgryv9FB
V1BY+q6IEnM0+UtKR4zf6ET70/hXk/SF8MoMjewiY07f5VvQLu6H9h7sPkC/U1ciwIrwU1P/m+Kl
fH/aoSF8hNsT1l/COP6Nmq6nU2HzyWXp+LScZT3ikweB0xBKWulmAKjWcMxPgGgn+qKhnsvHQ3Mi
W+09hap6Q5dVe9JyByna2XmYW4d1xXsaekBn4x45Thn24gPaQFpWKrNgj8XL0pn8+2WEh+NpkEY2
JVFGhb2Ignv4c6ImvJH16J4AJ9qwTfva9BrBSyW+TxvGUBocsw6Y6jDIRJImjiS/bfW5GqtUrlZZ
pm1qBY2JvSeRWxMei+mV9Rexuxk2zIawXO2gLLwre4vL032uqg/pMFiMWfZBjNk7bRxJGZ8e/9Cy
sprquAbg2Hr86XeYk5bfEQ6VLQxEzlHWSVR97h2SfQnat2xKgAQYWHxyMG4DfPYMRggdlgxtwj+c
FOENM/FVdQklm/F6AZaN6Xs+NO1yzzuFWta15thu+GF65QpBOLsbUO4Dd45zhO5kNKXeL/ATnw+c
Jb64blVgcbcWyjQXx5ITI0P8UAs0y5aNHx2n1jx56rohfvNRxTOfW8J3Ig4CYsSHtY+PcLw9r6DN
mTcggpI1fmzfO77JRT7EMYht9CzPB8p50XtMep/sQcjJqF32Mmm+D9j7up8bk4AWbExCke5p/cl0
mS1fbmYyTQkjwPhPRpcR5srBbM2qUQ83WfH8PzGE0R7IwgDXYfI8DY8UPNDC1WmZy2KywpUJdlun
PxKXHFejDxoGWLIR+zxYHR1jffOcvV+1OMCSe51PKjHyUQDVx+z+zfXqaVkG6YJ0AD/vrf+yOzLS
AUv5JQI6AEd5snFLwTkaw5NwPLmrtXmubKBcnvH6CuX5Ch8Fn54VAQgatIFwPt64Neb3BUM6918B
q8UEjD/kohOCUJBg0lN67OwmW6/NdKmHkUj5TEdZzce247TktC0FUCkJnb7FGIBYWr5Up5MzyImq
n8pHafKR7jr05P6vbo3+ftTdY/jRLB688Yo8R4V1qdmA1g05rdgkkULykXmOi1g1uBh3jEJUyIj/
0eONiazTplYkQcbU0W8HR/qDWuZjYFvLE6muKlAwOdukTTTXS4Y0/jdE06i8CAWWYrZnpQ4aZx+d
edUOkR0ZeNLhwpFOD0d2UkpqLi9V6d/co8YZ2QVP2RVjayIUcDLMws75g9GqOM2Hu5Pvd6MvV66h
vpz2ooueV/gmcx43rJVSIHVqjXsvPjuI7dYRxqb/uUFi92OhkBA/gSOWrLWLNC+f3PI7i8K1fyD8
2d+SKBSCUPSlf3OFGmBoRA8wWPSbr3w7MjglWa914WC2pVn1JQdsG62J2g632gCvdydPwiVHzHUZ
lpRNqBG3mId21xzW0lPDzsb6ct5NYj8JgpBGXbT2Ukp4uNASOMRMoM2MHWlGA1tg+d6LX9uK0VMT
8aCUaavEr1oaJ7q7RkUQjSbTnO5yveqG6JjqcmDCeCBa47C25u8ft0xLzSQCmrOOPwZuMgmNLslL
46hR4gmDID2bK/ThtBpX2hC16jLJ+hABoqZjzx8auAbNk19rMvnp6ADv4erbGYrlHiD/XsImVvVw
cTXYeMLaxjTHSHLkxloQJoiMagS6MRpCqRh0nJNH45TIgrlgo/OSwWtS2jO386UjFNc1ZxBCDF2M
JAtLhBv+VdELi4uFIskk2XOZknLy/fxmSG+ea8dvdbpVRkY1KGcwjojJkw1NmoyLt+oA9S1KKX6Y
lt5+ezSDOoXem1RVL/z0CLOgLhcsaIfCrW+dOz/y6AyUJ4pSD2cgIIHyKhLs+TIGUSigkjjI/afA
TfrEsyQtplEjV+xdhtmp5nIwmzWhapTgqC9aBliHUa2fjy1LDBq0EYLqU19CZ+dmp6H1XevHoPwx
BSN83JwacuDT/PTn7oMONY/Cez1vmn+gle9QdjHQp/klhvJnBUbn3fOisooRFo8xCTEn4Bj+4k70
zM9EU20Owr2AutkPGYF/63ZeZeAIKID/QPW4zqA9iuAhpFTohZvWO3wHd9FSG48z8uB/hLjy73cl
2UPA/5mFQSnVuiqrKyG9BZEKmqjDXc+rOu4HVjLjs2/8JirBI++fTnp8CdK/ZgajQfrc4nGmMQ1Y
Pni8jB30TdrJ9hx3qti8bpMSiCkfv2vOLquCHcWV3vYjA6JPHwZD72Md7NJLt65nne58NCgaw09j
ANul/edrs86uFlWA0wlic0em/T1++/59YCzFMPqzEqe3kvSjn0XLF1I7LnZIEAv63IgAelzoicbp
97MxN15ibnD3U2jl1g0D5+1L6QRcwEe6kzfwPPbNrCwh4I68VposjRR907r+t56ktr3jWQwB1fwy
EZhXMzldHBWlvPHOTIa/u+1Yq6DQB9UvhCtHNv9s5cd9WBjzEy7atHyLtAvSMb+xJ68+UNl71te5
TIH5FY6aEg3W9SBDba13NzQM5cNMlCdonWCgHHIQ5H4v5HM+m9cJaQcTnEqC/3PKC7lWaxwCcGlE
BqHssd7IpP4umsrjx2ExedTP07LS+wcnqUAqG2SZQqVEGK56zC3w22KIHyESbSv7q3ZYhtVYtI6j
vbrXRmsCLjyDvDfxwKe8MoqZkIg+Wq6ifjpBd8F1HHhsNDKkCIQj+bg0qkKZ0GlIUf8fD9R6n5Xa
+OlBRSLQK3u3NzA1LIbGplyKQE+4EDfofGCNC4R6f/5ezJ0Idkt/GlUjPugopIXuqUavfs5GvGhJ
kmZUqjLGoMffztiwQOl1FZY2RWuozgQfUMinhSHPIm+mDt6FqlQf/zAWUEH4OhvtZDX0y4ihWEMa
e3x5megsSEMz4EbNWuFFHY/ZKBq85hMTQ3+mg2mSjpQ7sVtWgLtNb56NIaY1GruVixXDGQF4L3b4
llbI8EFg2GSYcVaQkZMnUhcbyGTgWZREg7E5omgLWcTfODsHsdJHi9UvXIzyOCx42aH6AA4Yr6rd
gZeWLe9JYeMJvBdD5nsLcvdANp3K6iyg8Q0HhBgdPNgjFCni04ERteusYsEvVbDhVcKADiwct8Jb
9/cNHzNmByBnoiKsyNG2HfmVmy9gmVUIK+yx4vk18pWDIqY1tt6t6oQmgwU0X8fa84OAS/KXtBlF
l+ikvd3yUcx05Cw67OXi3Z3oDSQtdBSU6zBPC4x6rP++RC+B7tPbvl2OiExpHSbyoJajFZyhSCSX
qjgCAu8yvjePC/CI2qCfZbyRFdLp4YPNKVr/6J5oQyrTq//PSbvRMeFn8NKC1Mk6hyyRkEMsZjlB
BPduTulCXOMtKyrnSqE2D84W0z5NUEiGjqXSW9CWKrlefwGz/QwhcKt+f1N5SpILcG/sILq6ULtC
G5/DlRfdxRj70cC9uvQpL7/Og3e2DY9VxJKfq1EvK8bJCXpL7E9nS93Ix1pW958rC34vI8MwITYe
kR4ru9xDTxXW0GsFc3lo9oxehqoFVF6FfXsNIjquaAauFJ/nNzXNC1HRJAdC3m4Wng8udZypNkQt
NyC7hlmI+dfUVuoBj+mS6Q+7FtwquSuvT+XejDMGYMK1mFynO+p8Ccye9dEvEcM7hZu7vbjvAnwP
veTmIDi82Ywhr0mhLc+mQy6tISQsgP+YDVnqKWBcmpU09LxNnn6JkrGK01JWzJvhOYIYoDJ3N8OC
1zv76mSZMzj5F+/ziJD1V5hSUHu0MxLLzycorMAQ+AEL49UgoRI6OUiGBN1vqoccn3sbbXecGcFZ
Lx6iQldZ9d5pYdxMJMi42mHheiScFbYdFX33dRcqTQ3ZIxGpXamm+fifb6UaF2IusX6Q01bMUjE2
+TPLp0ha8BH/xlZGmzV00l9iaWxAV804RoE3B3Kzh2zjyBLdRNVoISdOfDXpkaOP7AtoqzsHE/lt
VMAVFxOr+qta2KYsDCc2pRMsC0Yh/tpTDJlHSG4q8kQ1E+SNJ8vTfxJRj0DFSac6D12CdM8Mhn0X
GDSMt468RcGDkEP1Te04/6JfJPPnQnCXwE+gXUd3bGmvq7CWyGt/VOB9WbO4V6WAUE8xPrSSiqPy
KOsa/UlJXGZnTkhWYDly9x90yHuaX5jlvC4Kf2AY34M3prb6B5HHV8vScIOIx+owEAueL8YHxMAo
jhHX+oZYW1WfvenISXRFeOMkbXgJG2ZGlF4WmeZjcMhGEiFEXnxq/hGqfGkZTRhX8ELAaBRez+nH
LDsYsdVueJAWRkD1wGazzXHC3sbD6NBqgspm1A0UuaSY87WNy5O7JVLOKwWdZyYYqbngNOTbzbHL
PcNM9YERKfNhPTT5sYrdidccqH4Qyko+YSZF96kdEPuUFG+v3t/ZyLnzb+BBKTs7SNPNnV8jh0g9
DnaH8rZ9tXM3Paim6asTfvJR4acROUIwvHG/v8fLD6VM1dt9e+oDCKSKNxYng4F4OOTytuICll9B
IRlh6sKcHx84ymAOONeayYYOrnfV9675/Le7XQRrluiNpw9TVLV49ctbVBlWop51IXX5tQJNqMQw
PKB9GmJAhKXi2Jnezw8ZCBjkZv7PBMUxT4mgfY0GWiK8PgpYIUxu9XPmao56agYTvcKTAFDCuq9i
eUShOTUTUeX2zGd86UmMZuGjzBxovaWSZgcK9KnB6X7XDUl00Zns1uI+wIHeYfe7O/JM7TtfjdNu
tBW/BbFBazT4AnTqYCxs+LUMgJOAGJISdQX97wHynIyZZDSieWhthFM8kRuMPrnO2LmD/cL60U7T
oXwGn2dVqs4L5uBj9FhglxOShUb/bu3BO+BwFeH4NNP8u6OVYNyI56z3XjSXyFTt4RSsrP22UWc5
LOvJUbkMzDOVC15xQITy3xjmmQBE7JfA74YLBp8vUnM7Qp26VZbc+TnvYEo5I9HSQQ5iev8Dug3z
PL5cznuXiyO6AkXLslf2f76WS715OhB4faB04+HY9F2u/6SrViGuXLv9mY2EU+dq5mfq8i9JrsLi
q3miRLGp3lkaG2VAkLj5UJuIGU+4t22bE5ZMvWpTHe792Gq1bavc1fsq76HZ8idisPSYUD63ZMVC
hFdjwLJcot3xhRp1P9FY13SEJjcT0T5WLKeVjroo9yt0M7TCcPIbeaRv5CNHBWRvsa56jLoaLjOY
ItF/kBwAPxd/sYVgx4neWsnA3wOcFo2RzipJQFwvTezqKaoNMIs+ircASIzhMTyOQAz56glfaQ6v
qHs7cyozZfeRa5olwv4AhMKgks+ei9pwi1A0UazMSBah9J1Oes4I1kOyoVBcpvD5aVN47GZ3OsoK
jgtVRTD++mqsleYHLB3FaLmMHdbY4NtZAt6oAWYyoNZvEt0CQXzjSM4iOiAsgO2MFKADxWhUaQFU
R8wmbf5S43mHn8M40quMlH5slcJLhC/skvJ3gydTscmkGXyhHhLEsxQ1mqGcovKbwVs8+WxXyE2Z
3MF+g3l68pAhzmra9kM4TyCTAPfzQjXDp996K6Bxq0/LV2QkUMB+YF+uFIdoNI2W9IcZQCYFZ9Ab
3n3u4pXpkZzwYirvIQCFj6THFuKIhpoPRUgmTQUFjW+8ZQjh7ln4QQqT1p5rqiKyZtVeNSm3Uw/g
8H6KO4gPIraHuH3fvXlhCKa2InGg78ci/7eFXomFw839a4ip7FgQv/2q1D+JH0/iuDNM3H9iPqV+
YPxfXDA7lnYD5dr4OANkRMcsrMzeurY+7y+dUiT0wbU+wgDLDW9gtMuinW01Cf3tJ36j+7Q16HcU
YwkHfcpx/NNHg2pTQX3tSor6Pt0ePfIffluaJWTR9be04wYJja6SBSgK3/hZTBqPN2ZlxvGbtl1p
jJjpHY67y56RmLI3bL2saNNGtyAJEGANT3FMOwutofeO/oOyXzkzXx60RtC1bro19TO6J7RZldNp
tVaEjynyUuwxXFZDaLg2EGfE8t22QrPXNIHNUdEqyYjvy4gOk/phw/pgNIyyNusEELMK5dSM6dHy
p9j6eblvhms/ZygrrPOlXPgz2jxzKcKkc889CnledVXJk0yRvYEJ1r88ykVx+9wQ9JZHqDAd5f1D
b7tBoRSmP4VkZXYbno9OQEfabcyXxnadrTJhITiXoPKyx9CjA9pB29LkGkxN7YcKa5Aeum6e1Ifj
tcAygsl/UUjlqT+vvJOf3pzb/Eqd6S6usWpdZUKhvF+PCAeN3uG7T068JjgXCFu9+uFwfPDQCXbd
docRGHBa6pLfQiZo07T52O/wOpB0+kROVEjq9EADz0FaJquQZl0HrkBuvB52gHm3Wgh/F83ytAp2
4TPkFOkEoqNK86jnO/Ufu8Ox9xdZ789QRq8507Kl3WKf4dl634ODclcThDfqKl5Nr0i14dUcZ5Dz
cOr3BnozFaufxP1OjFHlgkqZ43wfLwb6g48UVz9f68MXh7FmBzRiA/nKhZRpB71LkLeJUlM/vcZs
Ekrwu2gUSujsij4Rvk+WguuJ07WZATyyyV8IWW16CUsWpsJ92p7huTUMatQMqkQNGeOsdU0MMLph
4qClGwrVUgqzhXXDadizliWySPLUve7tvWhZumffha+i65z+5Xo6JzquDjEzSymZjH3pEBSKQ1mo
suliG/iMvn9ixkT7vmQBhek1ZCPkV6vh1PZ5PZ9ZZ+1jN4Ekk0AqB2UPah6cCD8IbWfzuLBvGjaX
39fIMVuHkfygP5wQpmS7pB6ZAEWg9VgnsXQgNDG1kWfZyIuzF1IptlE97hsCKJaBNmAMab2CyQ4r
31b2bUGGnuJ6Sa93IOSs2aoKwMrcqxzJUtdk7+g+KsvvJQUvyjp8cO7DeGI3Z0Z8M8igzoONVM6U
s4BvR1KSel1enZN6gcLIFODjIzNtxqHDHGP1xQZKPMddXFbzWdWCNUAQbfJOvpscX3e+dXtf57ox
g0fFdNQbHqlJLvNKsLkg3ut28w1OJB1JE/yl1yoK9iJhRXTpjNPfcOAy6KXUEc3VqCEGsWeaDSIo
iVC/ZhXQgWkVPuFaTBcRECco+thU9KeGo0DWFA4uppCJk1ZQkvybB+A0Pdrn7hP2iSIJZ+bhV01n
I29VOWCJENTwggukkju98O4PyzpsbcJ1Ln1gKtBx3znkmSh8bispmt1yBRGBotc3N6NWtzPz72H/
s58kiJg4VRhUI2N3Z+HQxdvm5F3rln2FVRbOZl0XrW1h85RALtkHL2hjSlZwN+6uX24zTBjABNMg
iEHvCcc121Rf4nljVUV5tms5qSYVLAEjC27NBB9X8CwV+TPfVW2ZpFChK/shPwZCgNj8Jkm8BWQX
heNUfMiIncQHhuK3koiH68MkfNzhRDnHmMk9avArUJO+BNANTG9grpiOzjUr6Sl1ZdNnwdKpJq6l
Y99AsK2TTRfD7QQB5Iemx1zpgV0Ea5lMkMVYBFxdOa9lRT7bPw5m3+DU1Pm/pflV1uBqCvbqEbg3
mfuzP1tsRMRJVC6a/lvOZfDO2gw8xjPDpWbfjre1JiYJW07LXymDPHd2NNGG9laa7wUneyAAUhdj
Lus7Y/twEWxnUV2h+I1zm1e/gz19yaHowQ2UKa6gD/66J+3D5+wkhmuzzKkFahjAbNF3rlzh2khD
o6ZMH7j3Mpis7WdAiGdEJf5MY3VHB0XgFYG43lP8QnBUsO1MGjmxip/pl+DJIM5EJJC8RvXGrjf7
YdbDDy/4aj55aW4zNvGTVdz7u0ZgB70JmwbNfyfjsMmb2SnhSPOFraeBXzjlh7fz04s/MpfUXGmZ
f5X6MbdEjbcZzp1vi+RJp1Eg+GxtzBmxZf4R8QGHH5WWwGIwuwb9kP062W35vi9ymMQoysnR9+rz
OD30HV+/8UaslpV4QkNuk8pifDbbcLvrm8llXYMEgg+52Z0LpUfLckr//oJOj1uqmQ1DlyJIuji0
FBQr+I4pAvr4wbRRXIW5/Y45nGOU4MghCUB33nGEO0e4NMVV45AhgI7g9FDx7sx+Lsw9X/LtrTq2
uMsrPXrVZcdQ6YIEFLQxjwa6Zt8OB6RiDJHLZX+cR/T2jTUAYxMRGRoCS4bof4s6PXWwiR0EfbnL
nj53TLiOMGV9PICF3S04kJKo3PvDRVY40qP/3ksoj4t27w4BeoyR4DqYKbw+qcm1fJlF5A4CfDLi
tw2JxMF3rh7ilsQ4UqESWBIZJiXWjCPC3iexfkep43xNaYuMPx2SoHqHztOahUQCyVzwLHfMh/tE
mLeeRYMExrhQ7GZwvFVGXPDsYz0h3kDbc6dTsZXslsHeM1/J74/EeKonDh2DlhpjpFSCG+B1VnxP
DzOxPw6TPHeJbc85Rtoy6ugJWqrGvyjfWkapoBqvmv8+fGdP8BfnGsSsWA54KU+0rF8KmEtszRAR
xVCEF+z74RrTHKP1PzB69fdmRvtJW+0YJLf7KlUOi+ZtEAdZ/ykxccUkoesnM/miYIBJjNnc1j6u
3LMK1bFijqZYmLnOxVScM59oebA+zsGckiS0DAEXhCSKC8e1ZD80JGGtjRw8kbY7/HjaYOZQ/tYE
GyMVp1agZpsMzSTDKJ7zBoIivmDXJqfHNxKDPgy51x6UT+Dno2a6rJr4nLlZPdrl39Be0gJHXQ/L
HWdct5aA87sgCaXixYAEl1y/Jscjhnhn0rhXRvuHAEfXhQwFTQb3zD6VXgq2DTGN3BfepIfy4MYm
jdaxhiAA9LgB/90IcIk+cKAgEOi6FAHDqQieJ6pmefV9+hJOzBgbQoqXVO8Ik6QhrtZ/V4QMcktK
6eSF7ykeUt1OJVgrxjHblxqR53RVBFNgtm9J/rQT8a/wGMBb/maUcaXxfxlWZ3ruQEJgQKjYjW5a
k+bIKRfyzAVorMRwz6N6L1osEkn+q0526cSe7/rzVHdj+9XGpljG2A03giAmwebi67RuyEX+tV9A
LV8atRi9Nf/un1Swg4cUh6OMhTvIOmcEvKe56l749YPh3kASotAmAqIWV3GQ30Trjw8tezWsOmYr
J61iwGNEOJ32GWO5u1erETqi63F61/DIGXFzPO79toCBqeX8PlGkkIngjhAHoJaZeVzYyD+ENhjn
JmNa8mO5Ixb+jRQMRAcULVgMaw/+RPlPKUWab+PSvcs/mk2zNpGeUEF5bZSZPjQT+fj4LoSB96IL
mQO3qPIUO6sWPwCPFsiUAXt5RSJ7QdXBN3mU0UCi8fNjIDWJkqQcQ6BkjXXHH8SJK6BdprZg+BFd
DRgJMAgveEee8MUEIGYX5nU+J5MHR44gWNRdK3r65qoKI6mmpQ8BpeBoK/YAS0VL/VLPoBWvEuU9
BUe6zUGOlGnNkJMknkf3ADTedgbPAbIlxA74GvojHRkoBQruJsAwxsP9lL1tcRq/xDO+kpaOImpp
N/cqtivDY2g1fvgsYCtaxHO0EXKGQSqfts9fsUAjSLWfa6BtS6P1DnLlOo5kzZ94eqkgeOsFjgkg
VPPp2zZQq6nAQ7dZ/hrGRr5cUgnw/toxQ3qOHwWKSqbFKaplADtPxYPIPpvu03FdBon1iGJiubJP
ir9eGI2jseQdKLxtoSe4Kq8AJoZ5RleKdIaadit7lWGJd+jvHqKRSONYhw2AV2U93wMh4ZYNSrlQ
7lw2QRtD+lj6HKSGvoxhkvR3cbYsXpM1VMGTPxe73X14WbnWs0eIej1hSggOm37u1JUxSjX4/bF3
nbZF6zkLn8MIS9k52O/L5qfy9nHEncs+8HPjtD6jvrkNdpFvvhH5fT97ZTTky/hSrpFHjf1h9jlR
+BsNAtUBVRD0Kmn3zj4UQnmJVdECPLvcLKg8ctG1yA1P1jT6L42NZbxznAQ4MNGDuB0KTNs7S2dQ
WVmjKejg/TuwBqv1mLT5GbAHq7JuICFYhBdylp8BLjnMPtUpVfi/EiT6zPwoH3K695aZBjcj7nMa
PRE12eQ0ik1GfVisv37HAjEP43KA1OO+ZZjj8mBL93tpNDBUK6Q3091/ciEqDvj+Sr6qaiPLNQup
GZe+DfVEd92b/VPQ4xeb68zKPPDqw36kAMNRWSSQ1Oeh9BSVnJvg/batW5cB9Fy7z2GZIHxJyEKp
c8l7MpHpW7T3RjhqzOr99lbgyIFm9FoCf2DcSXsFG6h2Gpp9GiDi26wfRaGWFsljXh0xOn4GxVmm
OEdtXfWZxRV2C6n//IzTQKMx5GLJtRQPXcNIaMqYJ1Eo3YlqxFq2POGiRKAtAkHxVjYwL8Kqk0Nc
oJ2W7sBrwGoa2evfnvLulYHPxQNmaqV1bEKkxuKJP7405CHqkH3LfFP+Pw+XVMz7aQ2eIJysVLfQ
egojJe9Ag8Ri4NtQH9rbcCBgPF37Czy6op0mq3zamhiO359cGvrYFGsRCoEjxJcl5832xDN09PGY
CnT6oDNlUeQnL045rAWNMPISGct9uP7NXGrTEmyIWA9GCivfBGXlR1cQm294K3liKDTXCsR/HNx0
dTbSxiPudK4tJr0Ja55juuxNhn7onKC2pU5A4ccyTzEr9tl6ORVdm6pN4P5ZW7eqndlaTMR2luy4
HX7QzrbWFGCtm7pyC/1gB2AKGFWixULowKLDoFVJL9w9tFh/sWNUsPVx6QFyNvs0E9j9j6lKdnmg
iNgg1zj6VSyCp9mDUgYkiyntBybVFfD5YDLVPH4igWhHxo1wENDXygXzWtTKTAkOwnYLFihO7GOe
L0JlheE54LZHsMI8W7ifIEercCo65rgoJx2NNfwITuPQYw/2+2rosDD81NwPoE6d2uUiZtREYxzV
2DfKR7g1nal3kb/OVqDOb4hjVTXzMbMbsaXC8wMNor9dKb3IjkFpXHK2CIXWPcil7jpsia20c6yy
z77z/SzhzqG9sRmWOq5lSmiEBDD5ThMNc3EjSXoS5NbWs4vI+5N3Af7Y8cmwNO5jmMCBeydvrtNS
D/E4innucoVmNh6JgORTdjsxcaFjZAWuO9WP3ShayVMLWWjHjUhbtAKDVHMk9l1WwGgUP0RyK2tW
aFo4x7z0VYALDh4LSGup8Ip8O6KO4abIbUYlJniVEGil0F3uRUiSF/ky2dy/v8BnAmeQU3WlrYGw
VuYaJgrgVsOuDmWP31wZGLNHszY3bw8cpO7zGO6j9PNaOn94+grIesxiac28Jl0/HJYyohBIybhx
4e070j3wGwDgDx1xatKYpHHfVSNWKrmbHP/t7kDAUtqhQvqsieVqKcIqlKR4XLu+BGhp/sMCzyng
loJ0bLJIoNnjMBryJOCFnxOoRr94/sGDxKmvu4fjejvEu0y/XWjeMA+7jSfGRW5Y1wefWtkBb44L
VbzQb+tNlUtRfW9+VN8PYsgCOLUaLMsoIWsq2N7bvzdACNUIKpQzxPyB98cpwr58SE4c3ukTG3Vy
wC4D5iwHxARO07FzQu1/DLY6t89pA8bQcFneVaT1FaoQJTxXw9fFhYkBBImtz7SW4cNJsqeaXckR
EH+6LDGZ7I3o0UNLhfqOWO376qnH+wbBv8DwhkmCx57x/ehgNVhLBz8RzTGu80t8WbVWYzqcfOeM
V2+Ff2sjRiUC0eDL3LbJGjf0dulVofoHcMsFTxPcNEZaBvuH2L4B0iR5NFf7mgh4FASfGbEmPVG6
aWkNWCKAjxlkucbse6O07PlEdhswfu/kWHgiQ80TL/CV6324OdcvIpu/2rN8eRcZRpSjb88IAnL8
tQhTX4gkzqdlBsaxhCpjPdBbB//q0t8BHftpKt4PmgXg1GPPKUSozOzzc5rO+8hukKo1BjjmxatM
aTbGtCMuhpUDXlTg9uX7zLoyRyRwIUSmEDGERwuCFUQBzwvnAPCLwZwWdzaddYMJhLseG2lgsSi2
C8sP97VladeBah3FVz9YbkM4cBZa4AIG/0qtc4HfIgNEGXFiVyxNy4GUsTuDAAeP8ut0GQSwHfCg
4JECqzfe8sI0VRqBedboWXfFVnrVelOHshm7h+gKIWB6ApAl7S7uzz2Tz7XQBKw8SxPcy8PLyFeF
DniKQiAvd7H7gvPNdoE2EbluIpqZMFCxMLImgOTY5+ViPIp549b+t9IyHbc9rXfvWskevWBOcNhF
MlUYe/bAC/idNMus0q7TWjpi9QK6o7mzUuNorgJsqWTLfRDu8JrikprdzuokxtVuAC7ZLut97lnT
96XkI8RyVsyGOhtbA2P04gc8kPGxryeb0OZwZ0lBVPu6OkMjDj/5fFT6s7GFf//Yv0Zxjv7r+px9
ykg/oKayZ2rLYbTKSRGJPcxRfaUltYV2OCInefb5bsYZ86iArjkCz81ZIVSM6b1GJDMDLIbjuZs/
53zPqpQ+e1rdo+2pj/M7miSX9ziBmt8EqSGH6TVBnpdE2HOmlt6uQHqhuTDN/ETlLe3d9f/RINy1
jBaCWo4hAq6lnPLEN229WTuFV7GDHivB9X303aHtvk+VdxVm1syynTeKIdfuLbkJTU564UNvRWCm
ZaSa9dmbk1FF+2vLlS5vmrLX9eSQA4XHNwdUFnyzHkbgRrwjSS6vdEjteSch1aAa2D6ikgZfYd0f
iTgxV/fNBY9caVBLBZEXFRzAMwU47UTlpUwAuTMn2X/2uzij4l0tcPAmHvw/XoIF8u9Vg9/MgNd+
o2mklYqpc1X/fFxGoblyuoPoASO41Rn5Emoa++NmmhBoTzltI+8/Ggcq49v3Q8X+9Md/W6rAqoUT
3vWSgJMCUbh4honbkYLfunfVIWSfAFvLI9nEGhWYpG7QnId0rBf6602ofcgJ1NN5GBiayRLKMLTC
Hk6NPNFPh5BS9L9FD6jRtsTSDxbhjVGQkLfb8yFn222oFmJR1aG4peqCZ0A96xBu5n4GqYF3GiRV
98tVHBatGTGRmUN8OX96FWcyxX3lu7SXQ1BFiB1yGXFg5aVb1PM7CNcBn5k4CO35WFka/o35kN/X
wD7Etb3hVTeEPZtmPjTayfJ/xbKxUDp0J0ZVBnVE4f6a5TYWaaBhgBruKtv0CQ4FPQnNptY/utZd
F/uaV4T3xw2nqq9miG5LN29V1W679tl7cq7TGQq+/xhU1ZVE8NbFngtDkurHNdwvOEfhKLVqKDTg
zxn/VqVq3I8Ktzt5TaAFcb8mUZ7UiKtyM6QW2CTOakhbLktPA4YMXqVPfMytVI41DeNKv5RmPF6K
xAI6Y5xVScwm/9IeAueCgiPKV94Khprwe8OwkkSy8TN/4QXnW1BDM6CXOmSHb/3F2oCTBWPzE0Jr
jh5ujiimxohVQTmTOFxw4bL/3HuCIku+8ElNoVl9DL1fZBECX8xCZcBGzCF4dYybAOQ0mA2lnEa0
vGDYdwHo1wawxR1GgjjX0YPLN3X8E8hQSUacCRDpqDW9GMuaYr+KwqTtfPPlWNZqWsK/9JkvDVeo
yijRcHiRba7X1gu8640ajJ8WFnVeC7jvuK97j88MYhUusu1dNn3tLjXKLHCsaqJOa0DizMBHELL7
MMTMeeWB5KjLyPQxLCo/R8OUelbWgyo7bwzfZaStmptk/7dU30KIvjYp8dHlcE6ER88SimZVlSU7
dP8895eGC+dsO0Xriz21YkFdB8F4oL8CRVC8gqz20ltyHaEnn/ySFf5dg2S3bASW6XXUA//4zq4y
OG/k8TcswEnaRrihYERPA1F177HbsRp28KRJJy2aVwOGJRD5SqIKVs3dqNC4ClhFAfxcDUEgJ7Un
fasDZKQ8gZV6BY+mRxFafbw1Tmkx0xHermT0JphRPAW9YyC8WiZzd7NPMpRcBwF8qTbkuQg29Mt8
/Hvi9B7A42UPwdfUrW0ShRnHKvZAfqzzlML7BjdiPd45eXijg8MbrEia35jZo6MC6BxZm/umZHBT
so4TgpMvnJoyrw1WgsnmhBGzrHK1WpwyApCyfXhuy2VWroLrmoR9Hq9xSTUFu5Ohkoa05KBDaooD
/dqgJKeeco9BS3ti/eJbvnGXDmFh21lJ/6hXBpEEPqNEZjGcoOI3nW17DPGKJxd5QoocORhFMm5h
EXreNeQbwPWFwd76tAWDA9W3kVwq+JgkZaY7P9yOdN0d01yiADwEpmVWBDsY5vD/r41nkl1MkjZ/
TkWvrGzYy3Tge3hAfSGAhN9YaYxG7jI8172Zt34mPCxP7r5noYbDTzGIzmTvQYRPWfEnQ/8L9OBv
sfQ/VVLV6x/TSVKKPsSAW572aWTSjHNETt1qXDxfPTWcL0Yz+hmdLUnQV7XAYwIJJtexhlC4VBqg
lgmlKzYp1RLbOcn/PN1GNwrwll2ZERobMfuvUenxyih9sT7OxsP6+v3NK3ZJeBvAaZLRtwjTojw/
83fpSsFw5cysOXWYtY8JQQc524iTTYi5ffrrc/UPnalsEzHUcITmOdPhrw2eLZ0hfllOjqiXNkc3
Qlgc5IU0nUcF60j0rJG78a5TMUHJ0uoT1bGHJJZRrgZTgXZonIzDMYNuiw/fswlIe0V99Wp/0G9b
CqD693WT5GncddWoNgWIUf/SNJH0VIRvdUz8bKIL6+BW/MTJTKX9qJ8In3mUwMtcgmACky+t7ZNp
PVwO9SxGidNLRhZVUrubjS5diwDmyZAQDhwEoVRvEDZaSiXlgOnv+Oohpyv4YcvJTXZFg7VTXlyo
pBIX16p1vW5QvQ86aTDuV/kvs0tVUJYA1ZBGSMM2RKvaO+LBj5vOkyiJUD/8GA07BMvjRIBPX9Zr
uEt8Jz+lryW/A/3+WhyphTx1qpyt9DYG8/O+erfJbaTCHYzHI1pm0n+ohpEvM9w+9GjtGy8aQRjm
DWIyozIUvPKsPNrnsfE37I7B51A2fYQIUNjuUpwVNpjN+uq3g4Jn3Zg/vf2xrojVMPWGcfBlEbN3
VQn6GX/BelTaYUB7XUgJ7tsjgHYpHM8PeptJEMl7+3Uhetd2kBg3kZhopV9Q2wAed56NEBo5q8A5
rd2lCxqWOcLgVhC4RJmMandXHNy3cqhr9lprTs95XX1hlZqbLgrGMouUQAnCO9cgbu2JNQT3hPW1
uB9voXc1aa7Ykoj40vqIR8okjgA9fJ7phmINPE3N76x+RF7GZHyaWAuJfCGtUwf7UmaQT0vniLxT
9h7rvfd+o8H2eSrr8Vs2OZPGAI1Pb5R2Vgs9mqoJBfAhZnmdPQx5CXWOmQUmMsvGqYexxAd/17IW
BMKwWaShGxW6bBwZpuLX1ZEhetRBv/y4OSBgSkzlAut5rywLa5roXezF+u9d7xQvHiI/F3Vt8W+N
qVSTfRTZ5wi/vM0YQom401wtUQhgB+0es63Dftizq7d83U4az61Pnq2lQWO0PI7O29fOycCiy0Vt
98mrB88nXZ/CPBK5M0JZsJrgIV+jb2nZDHX5qXmJ7VwxHGsWGsvuKCu/NtefhjmCiB46x6c0BdtS
/SjONwCY6UX5K32+X6a2YWTM12aD3GkJBhjA9JJ1MGAwe6c9PzKxSG4NdQOfDuwwrRLyufys+zS9
JgbGYhF08HW+Lywe+YkR7OKwOoV5zsid09Rlj847dosccUZQiarF7vuM2yq3KCqmUcz9EjpxQfFE
32NDdOiWhuVO+Mm0F2NCyVbYuKoBQ1EUnN67luPGbz/fjOSW/ZVjGxnKhUTMsXGcmA/ok9WXVYxx
ybCws+IY2DHOHX72ho1pW3lDNtk4ekflJ+/ciMBNl/Ww0qdRKS6nXjiQuAsjhoKbFRRYG9vyWykU
sb3Hla4TllxLeuiNTv6BKMwTXQDtokXPkjTilYjUrwGcjrfVc88DH1pKzjo5o6SLOm9r7iZqIFnQ
NXpIuRwhV+ZrGGH5ncRJZj5RfMLF/ySsZKkZFJwUX+sAx75a8g5fRWsRBijwUklpBF96COStuK54
dfQoZ4IROPCKik7oI5srcdJ+Pbn6T6lOzxmsXCzjYhYtObSCQfecr9RRe/KFkX9W9h00QDF413ns
Hahup8PijaryPhI5K+2c4ytl6jxYl0WdkUhcJP/o8oiNaNKKOFSQg0QiIVtYn7Ys6pBJtKNjTaOW
1ul45sCBg/XruGlmMU7Dii4MTP9ufM+0vcNzDRe8ZVbN2+MGN8toYdK2TqdcZ0iY8x/s2nwjrC5W
hM3OrcgNmyoC4KM2Iv+0UPcqGcfWxFOHbd4ZPko3oNsjFE8jLbqli2x1kj76H86aqe3mRoGWGI2/
Jfr48EuauSVxqnFQG1k0Uhoqj0Y3oxWTYH4t4riPkudiDR0azoVkq85/C95AJUX/rCNRaT0L12Zj
XZpy1EXZjdyNPIhX0TWu3PA+Hbamme3fZBwIHHkigeBTylB84scdTHYuftOegoDzNDWpRNKN4xg+
jR2B1mE8W2KqxA876UEfhqEZ4casvnRHycyTXIf72SIMWB83gcsri4e0EaTqg2SvltJeasalOuxx
2oaIP40SzoESM0K0miE2hRs10Ns+o3n+y+D1jb9xWMkF/MswCkwwXMzxwWoVoRcClBUfwDPyK9vp
GFVyUPwQd5MJVttjIKs8psqpTOQUJLddlp4eQn5kvMBPmF6H0lnk1ADXhr5dL6uonjbW4uAwPix9
GdJ8UacIFmIcmdcUf2EVmSjeih/5taVdL8765Ll9KBkGoiiLEWLp1D8dWJmaaV44q0DWiL3P+LVt
JFP9BIdTYErqes3tZE2gpIaHljAorEoO7xk3x2N6EPxHQya+ZB/gkWXdb9cU6niCTFNgMndrd/Jq
A21sJUQWM/tFby+NSOXS9392MB5OE6Ss8tKE8Vz/K9NqKHHZxZrHmNVvlnvbF+n0otu7bewVsG4a
J7+uxHnKDIHtdNVl4HmomraWuIa/8H5WN9gf4+1u/Y/nU0hkhqX+4iNAMFffRzam7bIcSFc5pW7e
UBoOPN+BElhFeEUZwIg8rzOhIqriu5Wd1sEPiXVBz6KxV17LDdm9w5wsZI2Tg+usmnLFbyYYDWti
m9ljAybay9ZPTuejRYLMMTJwHIff5MijgEemS7lWw2Po269rVma2cS6vQykqXF0ENXBn0fRdWgR1
k9WM/1bfRoAw1gwLvYXvosbH6KA4kCGHGJ8Oz1FYGX2oVGnkDormU4tbpgBuD+uBYZjU4Qqf4tqm
Lq3XgCG/NMfNIlW3THyQBfpzD4TVaFJbR+fRNNbr0QDggA0nzuHEI+teLIE8FF3W/vbpOi9dLPuY
rOM2T/cNWxgj4vMg7E0utqyYfLYGbtSDOPRtpcXOGfZGD186Lrm4lNOQ0nB0f5NjZev8M8W33dl1
CzHUM1lipobTk1oWT60B/VjXtcWOrNEk9GZb4Oej9WcvrqSzoUT+yvyXtkfI6uCgxfYTfl2PGHPG
ePulond6GeY1CM8SBCj8XDBs5imOLv+wBx70DQTHiNtSgjM8PwPXOcOtFlJ5cIwEEIp3ikma6woU
etTvXLRsa6oBpd6gkqNFfjKjOa/6Whf8ax5scBfxIIsRvqBuGS0B5PMdtu+SX0D3+IIBG6udWFXB
LNk+WlaB/PlYekJ3nHLHvqF6nP+Utb3A9lu19eOMp8ntilYE95MeCg6QxYki9cnpflOD3CT7FFNE
Xl3oos4GeeNOd7NV3bEdscNe5fzmZnBBUwBucw2ORdkMjPF1pHRBDMYOkPi1B46XvN1nJsZJCanl
2uh2+EwiCQR6Nshtnuh099HlU1nJP7xbljdMkPRJCm/o4Gnpz/tJUJwWZPRD54ehjSieyBD3ory/
pObQJerlPVyIKYKLyoPDMSvz1Z027/gT/2BRlgyblNnFePnGqklZNplDPyDUAj9d9ux9Jo8lP+O4
tsK8DGjaWdj5mzOc8wGkuDht8UUyZzt5/FRWKnhR5Y466u+9WLzzPRPdxV/yeEfHQVdte3E0Zwgr
4zOWMqst1MCwN3LAfnSZc7OMyMoxrShcQddIyM9grWj7S5pCI3ibFoZqcVYPFzO87m73diFdM+tS
VTsfWmN89Mz8yRh2H6MlCzsPbwf0Q+WxMZnV4xQLMqvTZDNQhvTCVrGDYL//srlg5rCyksycnJLs
3+5/+6kq1pGvNDbQtD7UfVxHBeUcuPc7NmA0DDYSx7FiWvzYdrjYxmTkzE9mf0lcOuMf51ZxuYii
CsuGJNOw3jwVCvYDK9JQ1fgGRiun156yMuab7u+Uk4/4+g2lRQct9SG5qa5Ky3oz7LYy7BVgO0LN
idMKKnite2o+lNkwhRJjW4wb4PA/QGz3kwSaz6cjjbKyeemkLHQdHc045qrpfVNtCcp+wHcjQi+R
+fNJG6D/1QKT9ApZtYVxPibvLRja+4GP645vn1OOkcSAAoMNlZiliOsq0ViQwMhT6ElZtPkgSNTm
AD/Cpal+uQYlvSuidx4hvFCCjSqosHMpjwh82kg2UJzVycLbnfnsV/Xkjd7JLGITv4LPRgUe8S2y
qSeyoCRMOyt6Z1L9uwS8G2oKeLqDm7lYwa+EaO4H5bVMDhnJeY6Kc2jc5Uck1cC2dvVJ0/clE6JD
0LZes7Yy397oYzcWXdWCeBiLKuoU2+IT/umHiC7ZTemOKrqySXTqR6RiWaurDeKFHvnCJfOpupbW
38RAJF2P39UIIKHblSReI6a+x2Ao4Jx5P8b79+34bGE+7vlqWsN1yAYH1mgkmAeAXxNPwNd8gAmc
v2vXm4G59KuagK2dmO9jhHnPM1XWeC1BqmbdtCt+lywCD3DmmqDY4l+Nk0Pe6dh4wP0jQO3WQb1c
cNaq7XPxQKyE04Fif1vfUq1w4LqGVohcYjgJ6OK7b7UwntoBmd2xQRQ0ds5YqMaA1fNHdc/vrSMg
BssBGN+4OZJN9ArpgTGQR3KI4ZGqI8NqFpI1H6rbWy+4OfR3P6aQ5AH5mmEqXr5g13BC5kWpMg9V
qnWbPHydY3ULQxwdm+fIPdWJ0x7Uxv4FRHtQ8SxLyRViKHAWQmFoCdEYT4Eo24kkr9VzOD1gqNk3
Sbir68qkAbcB0OVCrYqk/vGTsOrYHdyVDgn4GrBGVa7Pf+PBGItzO5xUtsnpFu7tHdFCWzD3RGYf
KB9kngRPGPPVRNcGo4O2PtegPrIi4epYywxFvvHIspe7lJxXvfB3EqxIV+W4xzuPDbyeucDKBIOw
m+Un/AH+HF1zavXgEEf3rb+JL7wj7QfYehuI8ZhPeSYwHtC0TpZC/PbMjY97UmXWsAcCCWdzQCDh
mN1R223rWbrprWLiJKaenjgyNtE6CqO+X78SCgz4iggzQ3pC677W5Ae11AFUuRcyAdPamIAzlQix
oTdSQ96S19Lf+w/rfWbYupKQMH4bALK/wFJjxd4usd9hBHaBaiipD0OLhDutubimov2srUN+Q4wy
JKjoUJ7mqVYGGEUM0pF8zEewM0tdZ18lUp7k6uCUFdn6KdqW7xgwa7Rw6yXrOiFC1PnhaKnvPzlH
QtIUmGh4ff6P8SH4TKMXVPRz+FZzCXgNXA10s/acJyI8jWl/8AvFC3bXDpWbg6msy8iOwSwIMy8d
4SpNDc6wZuK2oth+nKvp6agvoHIEoIXYsq1bDrAEppXYrHEwZ9JdXUIKmTAjwaV+2cCmw4M/IOVN
2KOtn7ixNsAKTNckLsLYH7pS48njtYUbJha2UXdOqnudLecOaI3cLJX2tOXp3+xj+437JycjFGjk
hH77gtmHrL3J2T3KIp4KpCEMaWLVC0HFSUDnDiabsjwh/cYyt9u5Mocmb9bKTIDVA3WiPhKxhr+6
Ta9fyym5zdSCPr83t21m/PTgpMUh5UrqXc1nLkIcxWe3LNsb2bLP6iwq7L13MXwBQ4LZx5af4USn
fT22tP1SeosX56I/YiTLhwkEqiY42RBlt5ApGUSmSHy5cpHFCc0578X7gSED4Ko7McvgVJ9/OtC3
33EkToMQ02xbhcwPGZVr4EqrdO1LA5ATk8KoNoBvIpjzu6/r6JK8EUBZfikUIll8YNmAH0j98xtB
S1df/H/g3+OlDOuIGzyUctMsLJI29+F6WE3vHx5Xdldtk1z/xs9wopU7EIz58x6jf0qGxyBMgrgL
DnNXHdW1Mt4j6le6DSiXEedwsVr1Nt8cj8mrVwda47H471XOuL70gmpV3IkpBdlDmXRo43ge+hB+
teIktD46wIIGgL7bLN5DWfvP4nMWMXyYXKq8PTb2/ARuAoh2KfChv5KlriokSx/O3Na8m6QhfmgP
8GzPWmcidBAcwJKZlKS5PUw9ef627ghVEfAWIICIJ/wwie9HqKX5H8YKuCCUnyCfC7y/XolGF0T5
XlGGWDaewg0AhJQ3y/jJbsvjBKAmcPeWcCG9cwOxWN8Fs1ImZsp0T9IYOMGN4UVfDIeCkqnXXuMg
U+K9TywvPRuoaMLwI8EsMDMf9DwZfUpCM1Z1E3zyQcehBr3QjYNhwZFBujet/iBt6fge+6LbadAG
6m7xQX88vESfixELqryJs/jLGlkBVweg3QaY8YqLswWAYHfg47rDeuwx0lMLx9HrkmpP37d220Nm
dekjlW/Wl5HaWScp3QIpnjORMF7Sf1BDBuU37iinG/w5GEafpkWKjF05zrmw95wZrJyIJEMOh/ij
L9Y/Pl98MxtBckFmkkLcExPl7K76Ir0xU+GlTfjyTtxnMpz2lL6OBdkP71nz+rpmYNSlcv6Tvg6p
z6QxQbFqlsXa2ZLhhO5rNw5/vb/Rk+7VQVMKSBFzf0thB40hMrth9p3xF1yb03UbjvXla6ZS8dup
6O5Hm/USOHyDo6JrgBmulBoElpp7LrfcBP6dJJu8V9woaC039ZNycrR4hPghc1K0n3bSlIWYUSWm
POHcaWhVN5y0CoYI15S2w1+nebTWKU1sT4wnyxWkLk7I034O5StJI3B92/Uc8F7BsTNRXtZrgwHr
LEaum+YsJG0jQ953sWardzCic//KQ5CbN7GvMlHWNINqtNC3RvgrkKOFsBqCgBE4dwsEJc0chZxa
cQBH8nqhzXV66qa4ynaI7130T3hESK8wChAzyQfONeGI1s9071XbjXzlajAmE2Vs96sDQJAtvWCN
t9NtK+ozuzoZ57q+pxUkhRprqbYFVHOrhmuLnUkrYU2EDiuC2jebCVw7uvM2ZiHh49PSb6Sje4FI
qV0p1d7aPSRA6qnuWve5nB5YMPDFV84nlCDZdwHbkxvJvVqU/A/PYT4AT1uvOf2yLV2L67KyvVWh
fNEQRkg2Rhu2DVlL/SoBC+eITr4vLBo5yZh2YgEW1YwLgYZOVl4dcWXQGc15cwOSXDtEGBX52VG4
WYcHL8IEvcr0nt+Wj6PF0q/52cbrNXcAeTZdGv57+t54ZOddAfFkF1oTcyyI9ZF7LZ+uYT5Ux6u7
5vKQ8wyKQgJ9+G+laYcQmj4RMnFsX24JMIFi8+FhLeFb/UlxT8Nlk33JCKASKd9i65clDDe/8bhw
Wq1ZpUIjRTFHhG2Vdt7ueJUb2nNO4xPdqeadz2RTHUDXeJcksiVPPXN33ukPN8nrhysxjcyNZ/TF
tOT192wknGOfnevjzjKGZ3fYaXAM7L6cm64/neUMJ19PAu8AG0ZMR9E9S6HUQvMVHXQtk6uuZzEO
/VPlEh9Elr1NTw/CqqbLk0GPt44Sg+Oalg9gf1sWKs7m7FzzztwV0EiDKuJ4AvsnJe0BsPY83h/9
sapURQdt5cvTRA/x1xmFU+qjtK4DTCNlOppAKzGIC9O5uZcfDNQbpg4nbXXweS36A25UdSDk7Xg8
HEHpVQSnNfeQfVsCTnyYM3ZOFDQWN+Rw9DDo+xqecKZKWnUQ2gEVsWDwm+le38Y0UdLja8sWtJDc
4/IPFbfZyxp5zqgs0AF40j19zhKuJNgUTVScYXd3D/zAb3LWgIlOy2X/tvXaoHyVvq/lHK9YQKx0
Udn9bGD42QLJJvYZijoAzDoPWU+GdkNyx79bNhIrkk3O4UvUuBNYkdXl+gDNXxWSVSSXqUuOco+A
oV5u0xROB8WSy8cVelMtF6Sso8e9asaaCScfXydoqFaT+RIT6cyOXQHU7g/PFJm1NpFvwQs6+5fe
qu7+S9UhyIbZr2gsYc3noKLXzWcdEA+T0SEQRo+UcOq3dSd+gkLhIrrhZowMA5ji0Yc63jNwGJFq
v2sWlJWzFl8O614u2rjHcyud9WxSAXBM6odBHBJ5kSut29/e+RRaO4EAPzBBXpxym/8bRbNTJf33
ry6xlZ0T3bG7Nnx8swrn9qUklbD8Kskv1jtQArf6eP29OZxMbIzOymPTyZ0AiTCccRogMrrbhijg
hz1DYwpFgBcqAFmYwYb3h20BGfe8r/MgbQwz3jBt5lnvPHlBo4YR7F+U0gomwJXJ9t+NrR9DG3Tb
kC23x573w9qgJ671mznW1mzRO7zg5Zda8c/G/a8Ym7qS/7QA/4VC0uXrdj7mAz/xzOhX0kENwJI2
jjGTwq+Ud/P5N3XAeM6W04Dg6d5Z0ENDzqSsCYJCq43gaDg4meeHVjJuheGv4lEmCz9lftGGVLbc
2x1dniZCmfHS3aJo2txO5wTwD2KJCg2TXLN8+D1xVdreUKHau0gnTUP60Cnz4TU2nM6ZmL+q0PZj
ORXsyGEIfUc9ckBfsof4mHUhNacn79AcX73lnSFeu+UtEpqBrJlqJaySFogENhQBWguUfihF0Uar
AWL2VoL72u0sOKUuUsLtT7kC64AzAyjVNNOqqHLAX7kiXxkujNTImaY8n3c7sZFumHHAesSjsNVH
vBhr7wUkNQkXTrLiBqfiVa492hTutRZ+oBQ/hc91w5XVlMWPE4HSdBckzMtCLrDS00xnnw/CXUB0
3aSNqbRoQZW4ntJcomoS79oh1iinjOFAVYF30enaEktCoGwl+Db9zVNQa83QU3yLBuD/pmUVfp67
GA/uiKJ2PfdBP+XDvZ08zICDmXAr1XFqfthYmNaGGPzcyW1JLeYEMW/WXMDoxt+5MSBakwdlbeFE
RqWdjqXS0BMyrGZO7s/pnssVQioUm4Uak0o/+rS4v2eeAbXbRsU1YGkry0k63aje8BgpYiv4DOMC
a4neX5HPoE3kyzH41O0EH2gYg+3NZh2D0My1K39ImmLcW2Xw/BZ0ZZT4co9tHgzowDiP3P/L6ZXb
9Igjbrx2yMzcL6niEVleIOvRZ/iKG5AWZE6my8MGTunMd3VZ5yF8tINMzQwKIEilTbc1xrDoinBk
/JLh0pxRD0xqdk4SOrtXdbQQ1bL+ZyLzreQwEdfY1FgNbJSFfGWMXb6WBebVOdErWVK+Z1zRo6dV
NpVRUPI8nEe7Daq5yIkUCdLrqOaDaBNvpC5XtY5Fs5p0z8tQym1sk+AR/0PVxgdEFbrU3TyBWeUu
Ynhtjnl6qcoZ6NSn9gxpIcoI2zZghyRKXKfcP/4CXs9Bt5ace+zy32y9Kzf8/q7506xe9MQsGoHc
6VWK0RrTGqNuY8V7DTesSc9xM7SkUp/AGyTM1yJPSfq80GWeLv2nf3cCsX8K7+M6RZar4F9hkv9f
E5/l/FDnOK4/Glem7Jqgh3wosr5/96B4GVrceaAQdlgSbPtyO4fK3TZOyDBk7ilZgKiaiNkTWlUQ
NmvYtXgobaEtRY6esPyMMqxhEFISUp2Cdo/kIcFvzux50PWmfHWilu0EbmVsZfpDlXdaDkHhwtM3
+E0PwUTuAWTbDrizPrbqz/c4PbMdDbZaMZyi54/lBJAg3iTzMwYRvjxFOBSJHGCxTgMFXYBoXpSi
ySS6fVOhsd3uIL8DI9qY0lTwch5Jp0VfmXQOb92ny8j1TaJ1tjLcgJ4hP1BURgt+xogEIPF6Rn9/
elkq/OMGSKXAEhKyDsUxkhJ/7LqL9IyTrfFl/3y5/3LCKn3peo3ipPYios/n6Xu86ob9UOW4m9dr
mNkoiCpAnk1AU866DvLK6o7KlmAxylCHQsxMuQM/yPWI5zabKVP0nlZgEW+rHUoFUkp6WdGqbz08
kzVrTKCCLK/gS9PpF34eTE1TuS20taZc3JJv1BpalXoD7/0uWfCt6xshv3Qp2JbbeReEWl5RKPft
aAE/eDiR2WA59HbGlegqZN7yIo1HP7wNgUvdA7Wdo93Xuuc9q/vKp9DXyNoL19s5Lkh70hmhOBCD
Rq2T2MqbOEGSGJj+LdxxZykBcBxh3DQ/dIGg+CpOo0DqB7ZZw1D+b1NQKfzlweowXMB7Uh4VzjeF
hXBuoqXut5QMg6czj69010t2bFMOFa+8rQR47FjmIMkKFtwHS0wQxgxNC+ymtnqOK0SXY44pBGJG
weVvSGvs3ZtKzG6ORgLEouXFqoIGz+2nvYXQBLKdSLqiUFSpFhqLf+DsCKSsIymSOPXSjoQ08IXb
tk+m8g/kK2df653PkebfQuUuUntBmtjHUHq37s8uEaXSYNnj8phtjpE6w5NXI/VynqUAgtsNFTJK
rOTMz/yGSuDT9PXpPf0neiNRMR7JMCO08mumYq11m6/G6qVnZ8pIr/wt1i/VJOuVJMK8AO4wsQQo
rt0+9MYUDmNNSfZo9H7LrB6uhz0QacsrQbkRBsJJvNow251mN/fclz+cWS/jDMNd7FQ1xm74GDXT
yvTSkt6F4ssGCto8f9rzH7dC3nRg9dqI8SI/yYlKQsZe9JycCDztBBALW7rOWeoWKEzvRyeZ0DEV
ejopJN026vCuQYUevDxCm57QDLTNF76SME597yZYJbVgkT6ZSsOtrvRZbdqkqgCHcwuaaYZa5gur
QntyryXJ/aqtVsRi//KjFtNhYaE0eqjp17Lh0dkAoLgyLTjN0Eg5b2s/lz82SXPT1TpK13narOBw
WY7BQGp1yrDeA1iCGsszrVdGq1HgmVMMMEShO/CLZ+WhKhhPuDpbAu5SNeH5jv/WF+GuHnuiKHF/
Tu1lniVUhAIvgNBCA9kH1sZr1McXTYDqVHkt4YPpuRyonu81+2eaAqWmlF5yFW9jQpBbXvwVYgfg
VeA4FZ+nlfPsPOf/WdmHea7aX6ff8/wbsDH1G71HYIH7wHmTKRk93t8NBueFUrIoV9dNsxFbo/uT
wqnn13dPUVPZzmXIMrbYU/UZFaWLKNjbBnOgFF1//rF4l6Oqrdrrj1sryb4FWyAwHM0diOcn5dhq
lfzznJAuxjTxC57MNnkWYVAVSBHwk46HUjban0uT7Sq5Ezaf6XBkS3s+sBm9k44d0PUY/M++ZaUi
o0498qqBFQTMtg6BrfDKBfu0282NrMycxvv8UGELF+Ut7SbE4R32rx//UPLxDNoQFgk6HNklaJ1+
J9yP7+qruBwlIUEt3+l/hBHPc3ZvoADqYyfCGX6J8HwNeJhJZ+UNpOKpi9vmADaofQ/FDxnIC2H1
CYChpPGpmy3SvDE2/Fl1EGYpHfEX5elYkOf6kvSiO3awcG1HMQE7JlWs76lwA0i9f2ETeuDSh0O+
tb7kaJ+2rlxeagCBvoeeQg3L+Z3boMldxl+qS0buBaKtlVp2lNybMSPvQuWsDcdqrjctzu20VfD9
lX4/JGftjlSSjquIt4rRI9dfPLdTzgCD4EbihQkccQErVIa2tRVLQIpnQa7T+kqcZ1XYoc/xBSt4
r39N87/RGHvEsCpj8SLAho73xkLqV23kxrHJriIrb94p44vXOz99HoZ9Bad/sX3m9b2BqHNWiBfj
UGMqqHrYcmZJwIG5v3qhV9piPZRKIVELG5x/h3/CxYgEuZIKpbgmWHrzf9+rPFWlhMwlAzjOnX2C
Q01XUgz8vfdI7JPQ2htnaq5fVrkoakEc5miVlc4Ymjp5j6joZE1DKDwZ/NG01bPUnKcT5+RB48GB
bHmaP0xhNIOuBrazrvGmAIYuW+RjAiBagkOT/HNsUh0UmGjHRpC10HTUIGdEOYZudaeaF5gxD52S
5bCsiOoyp6ISWmqesPc6zvQ6rSne3+CPGWxPuYYRKEEdlcHAi48y5z3xGRh6ngNOF7pw2hJ3TN6b
S9smCz1cGmqvQNWQUFIZcDdAL8n85UMTP47Lg4K4r8CtZjobtI8OmNiexh8yuL6WXsUeNX+PX5oU
AtvVNSAebQdjB1NSSBKriSkZDD43iGLZwBz1GyAwQHiNrfDN5Uogzer9Nu7blH9Mh7lzfrWKc343
SFk4ZQ0XyW6g7frPq7sJXYcZJTC3ujJXI24z9L8P60w+G8mp5uFHDKT1/ChVMsxSxyEyFNey5UBV
jBGO1uHOQZkx/ntnjwhHQWQeMwk3E74gCMAHyuv2blY0e7vWFrLKsZ7lOmwAcTsuHJxO5AwTxjOr
xi6beN2T4F+V2E0pgIJOdT9A/IiKE6yYsCII9sD7xMvru340YcMb7E//Sy3Ud+timcKl3SHyDnvx
utQWZagp3jbBBdfXvylYNJp1jubPT2kXyT8bO+RLVJRleCFlZaat0j+txsQHSdun7w6ts3XJtE4f
L+TsKBZZqYOtJ/LuLfyt6aZ1kWPNBfM/T7UeGztBY9+g7p11yEt8OoP/nAzPLaOqufZjkixIFFpR
fNqW4J4q5oILlpvqDxLgIauHrYC6oVPRIROLuu88j9Mxp+LtrcBX5N8SDG6GOZuLXLTMMBbQ9LK1
2lvFYoYE7mpAgxYEd00e4z3ItFY3sx//+tlsSFA37oTXrc+GvNsohnnQ2z2s04Wik7k1Y9fu1aO9
zGK1DduWuIOVhIJ4UzKkn2N/nB1ntu43lFGul+GZvtsUi1cVCg55C0pioU646+RRaXsP+laMR+7K
3eJ8Jc1rcDM4sWvhZCH+/WFlapnkuVY4Et56NhsM4YR1qWg3wvy86cWRl6oCQbD1fM1C/HbaVZFQ
ymUgCPHSEnvnvOXgW1CqnLoCi69+/TpSEOZ5N/GH7DRp5JKSutWp9HwalkBOB8uWMsXNBLqCM0pt
39iCmsGB2RDHPJ7+Rwuh85HyAt0tSMhb/8b9JlgSiV5Ajv/qsH6uKDcUr5wImJlL3f/0P2twk6nb
gK9QilnUYVSFrxzErLkEPUBySP2LigZvC3S3nwfdvNg6Soo9Hqicia9bTt9JDC9d81rXPnpE0k9G
t6sRBjFAYfw3alVLKKseJ10excw84jb6091U+aIfB88m0d4ZDtNKSDLkhCfp72EtakoNtxkU1TpU
55WmalhYGa0IHINOOIFOTP3anteSpIbwqYmBMA4d+TvK2LRq31zOp7teoa2F6l+okamGnmJTZgiR
YHqgpuEQDFkr+KhfmdEq78ZvG+0CTwGqpqc9ItJEJqm/XbTC1u5jBYptrzdhqCix39xGoDtkwdlT
Rez70tRHVsyGLabHXa2p0CEh0+gzBK6vYq0eWtlEn/NUnFmwiw9ScnoLAG/Og6B7QvFkCBgqu4u4
2Z87MoJwAU83hr0v3+5x7JERros05+4OKGMVGHxdjL0raI0nKoP00EXsZZ54OcxBcq/L+RU1MEON
TeFCXF2MUcJXWtBgsZSzufnEmECek+SG0zglI7qrxyBjUULpjdXtyU5e7qZgFn4aljywELEUKucy
np/6Q6m3DI2xJnFmrILXh5S0UoiQd4TU54BCJ3YMqdsr5o7TE6mzVXlgEigT582kx7uCbESnfR3z
FozOwtzvs6nc4RF1JHVJF7o8bSPqzhjEnW7oxwJKOQDDGFnkcJS50BfvLCnigSM0XpS7GwhBNd5i
+87IEO3YhBFapcG34gfbYb4iaCJ/5UtK4LtyB/+HR8AupAIu9bXNUgSDa6tHziN+jwoh01+U3Sz3
BGhjau/WcUqJu7HJEhg5rnRgDD0Yn5Lj4FS6fSXwOV7YFdqxCJZW+/AWLzWHs2HgFvsJfPBPhyZW
Bmdh6hT3w59NZbuMqVyruOgHeOlTHKMFOtaOL2ntH5MHQ8Td4+DYMwDDeblY9WpGQg2gVSb2lcJy
BHCq68uGR9qtcjPVGyayaxp6Gmarzf8YUw09npEQoitGdY013jwhsEirnhLPgKnEm5XW7jUQMlK6
PBGMC8aILTNU5f4s/f0S6vPZ1i5ke4cffQO4suc5nTitZ/+DrP+0KVRLl6Kn4zch9VIDaIxgzFKd
8mtUZvR+ENTniRgi93tawqZXa5UHltE6f6W3FPv7pTEUZAjJ7skqeCHYwD1ngbiX1CoZCClT0jol
0YxjrVPMHKFe2NBBMazcGf9wtm/rSDHgUQPSACgLiyd2nfeDHgcdyIW6qe+8HmoygiBDZ/VCHsl4
sbOEiKY6Ku330fagFkOwqoo3UE4VMiUO9N0oB+xx6h/EjBvri77FhmStR8053V8DK2c1Mq09pu3h
5Ry6kxHfQ4GnRszSBhVsgDxjgS9+adDAk3wO4axwP0IU+ZSDzy1c8MsY9jyEBOjaq4eLOWqwU5lo
5bKYqCr1WM/bLE4zbFVKMxf+h8kLK6mSbEPs7S4DmsxyEYXdKd1N3ALVGGhtB10RMPnDR2xU0yhW
wvMbxe4jKXjc33IFGRl0i0YZXQ8byXbCGcROrlmArecHGYyGG8mSt2xaM2uIH3BZOagASPVq7jB5
ee/dCpR2/He0Jp/oWtD+glcizBoWmkvf1U6eXK9onNVPB8jHppbSSKvQgm8B8NgfQKOX4yZJNHmV
frSVaUuPs91u77dV8dj0V9kE/ZV8p0w7MA0sAqcWR3DOZIfp43MiJQOreXQbN5Z//SaG6Sz2RI4U
RDBiyX1ZH4kG2tlNERCkQDrEyxoqy34JzUxTKMJmeCTc0KPL0R48DcNi59YN2BCZAc/M1NZtnqnD
2m9Yn6dCQzdR7CMUAFyBfldpJUGD/jARtY8UAUVtYz+3qgCeR+srFuNd3HYV9k050CYkqTGHOtyi
4CW3Hp1Z/vQFIAd0JLWBF6JvMCPXj2RSxA5UVix70G5AlxKsDs6gqHDjcwWyzx9FiGpI70e5SUMX
V31JL1ThFP7HJWjUhTXJp4f18QDnxSg17MH3ZCWaWATCx5Z3CzBlTNmfuFKDu7hYrt9BesG8norl
M9Vd1Mz/4GiwZrW8h1rNv/SEhMm35d3D66heQk6ngTRRYbaHEH41NgZ2BdHyKlZC0TRLMgJKlpwV
MNYeuc+6aPAgzMNOVjROdXYZb290GUu6kIa2OW6GOjYgMLO3pgEfBqTzMxVrO3OlN6iaMHD4ybr3
DTA0aN3tJ5TLIFxdD+0cbLUrWh+T40oPt8Y/H4sdceOPvNShk3JFtuMmtTgKpi5lLeJooRUavMzT
N1PfRYtg7eDV2LWu2L8wJQVPWBc9P+WEcLSkQjeEZPrtmLcsXb+tRJntkBWoaR61DnsT7vGsLaWl
5krYddhD/owViZFptSp03YdvfUYnLBtUJknIhM/t/oynC9lrvbeh6qUIlmtMeh4+uZlW6WhPGw/N
goGs5zGs/pIXdWeldRK9Z9wS40DVrRkcjdPmiv/TtzZceLWP3iGccEnDHJwltb5Uo+XWf2bDZE7P
OsGbQrAmVdQ+qqfE/N37kevu6oetQVAwaKwhwrMof5rO14gsATo/O4ERfCOFCzESsAwzyJu2vaIr
l3DKSib1OO+pZwNlgcf+cfy3Ei8jG+GDISZvQP2bR5aJWnEiR+DnQ4J8bZzNGGqBNUwx6W73+/6d
249OPWklSLnC91YAI6+4UBD3RR6VuN4svY2AoTZwBfSjvj6ZOtfJwTlkcXvZsTGhkoQliOD19HTC
TEOdHxerYP+IG5OSXW82i0D2l4LKtGNayI4b5wj1Au9gNdrtIpKB0Ea4u+0MKUIevltvU+0Hbfh/
Juhr6pVZg2LHdmU9o5yyNx1ALyaV/l+l1Uif9K0tEr92goy+tfnUG0Bilq7UmWKp+40vj2J9O9HV
D03l2lDf26I2QEg1bEY7sryQJexq8gS9wNc91f117y/fHIhaszay1UwpffuICzZazdGBaT+OaJCV
vigzG/WiMUCK8+yjGsyOpY4Z2H0I/9BYGTHd6bqy8GO/lxTGiGNLQ/aviy2exoVcnZDALsoaeVP9
sNpnSodx3N7jt8OKXDMKFcKCHJiRdVtHpm389Zy62I6amgbSHqRmGvy6+yOAtXUXYwxY+heQmHo+
8yHqNFsklNXnGZ5IZfZ7hfvBWEBy8JZoiIJWYj8NxA9C+iKI8U7iWlD/2ZRxLFTUWih/aDZqYqVx
4IrM3kPcpWnlB5+SkkIp/L6kC1zh1b/PVmDPOtHyAqwtdIq/JZvGnLOzCg/UTG48mzZ1AigHwXxZ
CylYoX92qDLkMIw2P/JzO1Pz4jR+pPkgLC25mtFL7j7vgLGvMmMp0kCOET9rmTaHh8aHAHU2sZAv
gkAqoikK+f9tvjtL5Lcy0UPPvTSaBj0hC8bXR0pRVPqGwafTYHDS6Vg3CG0dXAXhSUoeJhu1D+mO
3qGEU20n3jPk/A/C3574ICUqkJKqh5hi/iq1U02vGxNTvmjVaWuB+z4CiKGqIofEvq80aNeV2kr/
J523igTKbScV/Mu+VNWiKm9ri9y/ixl8OxmugtF9tj0ZtETYlbSgI/6UyPhyjon5KFupr/f87Y8B
0cSd4iSvk+vEBfeInD557fZGtd4pv+oYXep8D03HODGNEkfD9utdFKcKC7kEbGTrzTGsBSYb0Zyh
F/0PyE1bQ+Z2FYcPLR+cjjyGF/V66XZCUQqZLYUV5tO9OhMn7QAVBcao2NOghi2c/1Qvya85tjZ4
Yr6NNsutSwkZfQ7y9DmHsV1EfTNX3/SNyL8jDxBcYBNC8/T1pKn5pvbV2hF0EqvMbzi08v2zvs/j
jVrawly6Ay7X34TCzOCqJ63WFsHap3OXfuymxL8wKm8XOnRRpTcJirMrrIsTQoREISwDH/DM8s9M
j8u9pajc29bsmDbdJyHWMw8uMnuwx5H+PoAvNP610Azc7m/3+97/sA1tRpvdJTMGwe2MkzUO3W20
w1KlWnCrXzfvgXB0eNWRVljWvKfxddnoNMb1ZYGWy7QJdzj0fv84/K6cph6GgCNch9UOgM1NE4cN
qtukcECuXDMZmE1cEyVKHwzlAiO1AzHNbb5OSplEHa5t6lLC435uc74+xhJdSifi4hQ9n3Anyip9
dtgqOD9jASStVnFe7hBX/qAcT+JwXznAoZrUDcP7WUNvwSOtF0evLa+UcClV20qTDHY3Q0XeDbiH
oXqZHlxh+s0DnEU3NxguAi83NszaziJdimfK4qrOsaXAJpa2BDOcJymUXJqrYi6c8pWPnEMKItMD
1WEO/68iNkZddNJFDAJyty/l5htkQWTp2sVExzWFjZJgE/L41Zs568ZxWDRHLn4YrJv467M1JpIp
kiM6CV3h8zW+NHDoZe/VKMMG+Qnd1NwXLKKvKLJE7Tpi4myrDFTze4gPZqUyOrvOy5rc3lMu+I3h
NVngWhJhQq9/KEReM+KDroNz/Sq9Ms074ejNFvqDCnStNc93+zz38n9Ghz9ZmDuJEgbOoIUitfdI
cOYVx1hH/G4c0QmlQzDQ9ivRplf5QOPcwUGadvMTdhjiUpARa9/2ZnX79v5W9+5KVeoXIpKUghd5
MB9+mVDIb8YZjYxBYoJHKSrWhhuGS6E437Zywi7lTIEmNqta318z0rOCFFtwE5mw0hlpURyUKqhW
7QrXM+TeLtgX5Lr9DxGleX1aGiFcCbCAGDsncBS0tU8TpY01XcLXPTVaNhdSCcZ2Z3AkNYogYP5O
qJgLDKBii6HRCaFpQy5SQaSSPUFnmc8D2gZyZe1JkN0XIc21HrVqmUHNSEjvQIHAvTUXrYwPQNq9
piyStf4JW+zkkYGF1wsNx81nWkwVQIBevXH9Pn5lUa9oY6mPaOJE7A3snDGBCnPHdFTXfJop5X6w
wUdtPc8rGmvr+Xn8YI+PD5c10wgCwaR371iebpq90bQt6G8itx3AQ4fPzCf7o/peTbwPFaV0EPkN
b1zIR24s/aqyF5r+SYzyq7ooQjb60IgOca9PSP5fjH3JjkzIoBhp2tMloM5TVzk9bu3kW9Z0DmH9
GEcLVO91LXKPKkAJX5Rm23Kz5zoAJjpLQJkX8rrRfyZfgdl7Mw3CDFWZ0YPG/143Vectn/JjF8ZW
Wbu0MUC6EYny8bzpYQeBQOcxbveUudC5v6+F6HuU4nK0cfBwPM8vGRXVPfunpSey35yf+60RnPie
qcgGrfM/8GSQ8ZH5hLJXNBeQNud3NofrKwIvrIVXGCe5yede5RW3gPmG3H8gWzN0fwsnGTH55w22
1rfChZIwtQkYpjqGPw5spQFk6TB/yA8zzhe631UHQcvYJdAMPeQwkdP130Cb4L9hB2f7OgBuoqXP
53dg6etADO62BRkfAb9Z/yhO9uV44mo+ynpEv4i2oqUmYaIdPvR3Yr/wBJrrgFLGvUjInFmar2Me
I8fJIZKqN8QWxa5+DxUdR963RvqjqZ57Qs9yKjtmHdzcxnM8DLTErY+QOQEr0hCoWpnMIsmf7R0x
bTgsi9HjhPLG+0MiBeK307F6sK3erDM+86LTJO6wai7QxTcwcjqeRS3iV2tCfAtIoz/ehO3tdMmg
61BNrynBj9vvR/h4rBTBJ9dMIfiTIrM5nGUZfBtfQivS7CPS64f8emlYW1DoKHPXKZJXZAheu4Ic
MELLb8N3y6I0b7fWrAEiRj3M3N+amIVOpzqkV20pDGvmyQl9ldtmgl9RLdQR1Pd2M21i9WpH0O0n
XQeTxQROzQKIGf2uJhapLfTfOni8zHu0Z+LuPdsAg6Z7j4CXJHGTLpYmv4d4GmtHg6v6+j62ECPD
+GSo/HdlTBxT2dACiHM7+ovw5lrjxTmPP+29wjdcEe2MH3HrXf5p3+2KwTsru7HBvuxB56zeu1Ym
d72OjjBh7f7t92Q8h9G30CtVnhTkmcDK+Fmt3JFTf8pTRnlsaikH2QU84IFFvNgGRLZSSwCFK18G
aY+CspRciZIrWSXXURSAnDq2GxRc3fOLAnA0rh/ksKit6b5Xcuv15j0FZEBPJOuhpukjo18Bi1Fi
4CqZJhulg8Xhnyy/5EIBueed7WZRR9jn7CokdUs44PzKV4kT3VjtRq31S5Pfr8MBO5116CBpyLKJ
5AodECpocBtbo5VlmunlaV5H1ZG72Am/WtE8PGbHdRi8arc/lHnEYnUJV5keQ6ggvhXOC9mO/GOs
K5IyDpPv9n5uo8Jg95OxvnYqf5PljrK49REinTRotk+s1kG0yqWMpwlgfKru4Oo3GcxbCFncIHxX
SizLdUtTByzstwWerPsMh/wih0KJuYikbAlqQ2OqFZzKzUMZrajBzuuD59e3SXPyPyfdPHDIg9M6
yTWp5ZQbYXI6bq/f/QyRg7yQHpm/2O9UWXVN+UYUyQJrpo0vEplP71sfxeB94YZ97xeY1IxgvAM4
Lf0GdnC3qQFX0Jxse/uttxojtH2WekI8ZKEOOkOZcfntmBruYD8OKGw+nd8yqDbgtSdQvZyabXeT
znhFrSHVolSo8VKRhupV4HG8px1VyS7WpFrRLj7uYlxC8lJ6dYI/Qw4/1EKw2RQrgSwZW8qkDZ/u
cq0TDxR9UqRrthOyQFE34QeYlakx44BFav/LNaVk+vk4P8Y5Z23ELUln3e7uu1jbBUQYxGpkul4Y
Nn1Dym92Mvs5RrZXPE3d7AEAYql5+LRmZjaL8wAcspWHTUr/qsBBcAfmF3y6/AlToeL9fGYDtNw4
o/GZGaUibzmTcDLYO6cqk/0WXnpK8e2FGUNiiNJF8SH7XjjTXuBuEYci3vnZA/XM/x8unwTFVb51
nPxVza0p7OPo3LeR0e4gf4/c3zBLEUlwjpfVT9blV2F6vlFMd1LKGgVhPRByl+AQJ8ZuZgZQSmTY
GjWSaP84c7IFE9MST5TMWKHct1mUPaAWPzBs0T/M+/L5P3JD3IRm9d/qu8d4W8qiAmyz78qpDPIu
VqTaZQkOjsRcIRHdRlUAQNEXD53S3PbBs+xPsND5Rt+yljsJBS++jublsiLcWyb9LkXODAC5RPHG
qdspdazwgjR8S6TWYbAk1iUShHXKuzw7/sG2dQ4SI+1I5jMmRXaJwityloy08QVY/S8MSVFXpDuM
ycMYi/Bc+71dAL+KmMP/RUcakFeiKWYXZunQWwhM33N1KcuBW72wgO4Dskss5CeC5pPqqnQWjvgu
7jq9c5yxAG/8Gd//gokWOG5cSsssSbGovZnfdHAhXlTyf+2gKwcUchApxo8wsb0VFr9dSc/sJjAK
bldpCO1EHag7LskxSzRtlmmKdJmJLSA6YB+g77AiHT2Z4lD36CAGsQIh03i/Bjs4otUYjvsHwp5D
iPSo7gdQ7xKCNJfAyNwa+yH7x1RkJYZjU522JA+kzjcnZA7y5JZaP6jp0d6JS4aBi7Z490Aeof4h
UUlT/EZNs/U8mco0An1J7mH1AM5WTLWyi/1thjz3OR08QE/Ce+tkODY3RNOhgryl2vdyKB5FYFEU
HUVC/FxhcW6b6t1z3Jac+7G6oIMAMPOuSxLts6otpi+P6B8MbZ1hTFXa7pQFwf8J5gFnxYcev63a
+5Dkhk8866nfzYRnzYSXYUqIRYo72wxRb8v4dNooAXTz1cSOfTb6WCZWbJinUH+/8F3Cje4HhlsS
PCWP7Y+pCYE6DR8ID4xcb/mQP89LgHHCnWeJjD+Rg6ez6CnOs+1qjCiSGJPj3yLydduuJir8N6WS
x6kWkhrI5AtbHXaLYLLZnupYop5WcGjjADzZLt/Bm2W58q08WbDfNKqbDazhGgIuDvCEK1OyFdcC
k0ql2mKTS9ZaC3SXIuQWx+B0A7JYgkSDSKPj0ndX7RUyppk5O8Z21zEzsYFQOs/jJ3O90xvGmgZI
L4eXc5dHlDTs7ODvxjot3iE7AUM1tKb2Yhj/MwwGCvkaTKxzArPTXl/kg3G05tEbTO33Zp1CLg8l
qHyUk4c9tz3+Kq1RAD6zwPKC7alPaS+HlvfH1QYscqYzRP/34OpirPF8ybWZMAixajrM278sDVZ3
Bc8PwGzpkQ0DEN+YzFgcwQQjWZyBF+vAhAi6/On3mtfrhZv3bUIaDycW4TmlLmNctLtUGBk8uG9U
/RQPZCNDmEbEl3GQOKgsoJytlkAdhcvYXu/dt7vyb4XJL2NIGtxAn7ejGswgK43h2o2YISH4tThT
ojlSMCgWOHyEZcRFXn5oOPN/fYVRrIvQumpCBykjmtGuIxEHyOtnSgxhobfBy3ezWRthmXegHeqQ
h5QzR+FezbqEgOoquinhUlfcRAhboCk7bCR9NW3KNQSVkYtdpE6HRyyGuqIFY3+cxtnSSx2w7/pC
j6/Jw74S9W6VemHjgoExRPNlrSwatqmb50TbzQo4QDaG0QC8evO7vubWVB/OrjT+Ygl4P2RymvKB
0z0y+eTTYsfYuxhY2Xqqvcubx7nyVR/DkXGNmDN13tNUPfhe069+dATpl0qFGB+SCeCF0CO6Ji/0
hV78+l9QT8UtuSL0Nl+D9aID/6wCUa5l3uDt8Oq72hAJGAsyc01y1Fgz0ZFAY0EXn6EUvVGZm1Ty
P+KaCKDgvJhdXz2v3YaCfEa8O+/0aknmKThBZ5IJpCjgOsmEZXE2YcSH2i3W4X6x8Xmhht1GJNle
7v/QnY65lrWSVjv9Q5cRZLPxR0eFo+2zwTwQ9X5m5euPPFP1TBO6RRDJUvI1yN190cv48L3tgYb4
xp+BXyb92LJlp8h8SjJdsbRc1/7vb9rFbTWm0a347FwaQVWlsFWZCJHGHFI2oCNR7TsbSoBnd5DJ
Coo5CiBI/us62D9KZ3rl1wdnIOVe3w5lVYK2Xw0iY0nouVThb1u4Pt3GbVtuh5n9YDp+QmTan1m0
CmkWvo6UIEBPqX0S+DAzs1MQpCXXEGg4NFdjknMFXrZd+PQ5VKP5W//msktRkTMJnUsGBhXxGGzE
Mg9ScWF/RnXlAsojQPKroNFCYCFZDQWtJShZUo6oEFDcKABwJfpPeANj4qVtUdvNfZMnMrP+74zG
I2gOdyAYD69E1Utfp3hLD+aCzj61TZ6+vLQBw7Vg8wire6/d4KrbXsXojSEF/fvx5IpPHbNcZAbz
mTz7Gcxd0MiBKLJrmhWHPaC6ndlON/PxfArpMBYrxFqve90vsez21/9KqmTpgCCdSFXwyYMFMkNs
VxdsgQammCq9eMYlrwW7RQXh5hCtAttux529ZD02Cfh6IjCVNYfQFDCak/8qhAOMq9FFq+h0dqCH
W++KEJSSkVfqwTN8vLGXzubznWcFLR/6BEPV/A5hVKdtxqfnehq0efI5eiTtOYLLgy5ekJLY0D2c
GFdsfSrPsR5iRF4EQl5VMLUPunPT0sgHhdnxbAqM1/dwDdcJ7fI7GmgOjnbnS8pFpUxo/M2OUUKQ
Zg+pooVZ3V+bzJMkGSTqTsSEFbMd9GWVbektNfiKRb4bQfuq9jX+UDLQbxglDSUEvzwNhNw+b5bk
Q20C7xpjF0Y5GseaZqjkEhJF3vR+xuM5UKg8hHEfwi4SN5wbt+HvEgqnBPmcNjvsIWtVmjiyNpRH
GjVOsSRjPx5MCE0NbXtVlEBCtJt8FWJW/4QDq/dzLLzHv+Caa3pe28YcV1n/Q3ryqk6ANYbF8U88
CjK2VdleZcz2AhXyNlxIoeek1+wyqMbZllfNRm1EG0U6GFp5wmIhjtWUSq0r0v5TTyyg3pFRbKsc
/Wi9ClfPqQg/om9sjAymjPl1rvkcAo7XHExYD0l4hJnrhCHr+DnxlaiUzJDoGauokuRH/5CccdfX
75aVm5GCD8kWYv8skd/ZhDJ56ukXpMPLrcrGOqpsCpM0F1nbtoMJCXs36uwC5HZaYYiknhUsVdcp
LV66zVZWTE9W1zUFHrUr0OhBNMlU+f9n1uQLwyxgMmze+D5fnz1l1rxRUbhux3G4u/XC/VDtYhOR
zI0HmyOoo8vj6g3vmPsHO1nEevrMFKX0Sk/38Y6Md7tSoqrx+Hghnj5iLSizjfW3McMeDHVp0ckM
GHKvL0vGEOHkHO6SkyY7+oG0Llw7guOqFtKEYTGvhz6C+bFBJ1zX/mNOz2OfdmAA1lE8ZgWajFeS
ETiSglIPKMhwHqgqCUherw8A80PEMu+tYUticq2+6Y8NiN47oeU44v14jTqYB+lZo0cSTMJQajtP
JBW3r7iTijzW4XpMoZ2SqdmCl2fEFc7voi7dtcbZJmuEZnEXMhQoVGIwIMAfsMKx8Wi6XAJVsA86
BKhLc6Y+f4lTATcPhSz144zG7BgiMde9RmPWSB73SfDtNQYflD/4xvFj0mjlFlE72aSfVOFWs0CM
JVn2Ivk/iGod9MDxxOjQz867t5nECfFqtz3vKqdQl1anzBsYZyEwutvM9RQ/XecLTI+OlZUQ6Kzs
J23Uriist4yUFPEowuh9nwLQ8X6ZsfEYL8eRgAsnk3/Lg72rBPOPeFjqt3im2AR8yEoEfX14ndw8
qWz+GAzuP3Mjj+kme03/3eYsE3FXkVRVJaaCOEA0fIG+7uzQjJcbYmjnOI3tgd4BIziysv4mII0J
6yNBQBzAltY8Y5ODN/pvPQ+XPuEYs6W9PGuYC2b3htb0fEbq6L69L4x8hRciPkZu8nJohIAor/Ar
GGYe+PhYX2OvC5EX/AeYZnhMRZh2GbvsbWvGNV6XCeV3pJeYjx4jqRjhlKheLP6xzEWLIxsfmTD1
j7L2lTIy8Af2aIovG1nlLF8QXBquX4OxbeNsL+22RJCiNzAJjvkWlXUM+ikrepGB5u08zNbqak1O
Owml6pI6AkpMKB80R4RcHVnMw+mCxTz9wDruNdg+EFZyciEw6257xq0EvBuIDzSkzi6InGEjj2lJ
7g6Ygb0wre5mapryUrUxYsdG7gdQxRXNIF4K+QpPcdn5nGglxxAEfa+kCd00EShlC/z3dEZoSRN+
74kh8s7lTK+f91Z8tUjPHERGvM/el+aXdGhR9rofaUzlF2n3sl8RJF+unbpP9qXbh7NxzUCWuzmB
tHYJOjW6ZGR46W7DFaQK8LVdOUeSLqwLvyxm/DB2wwXQTygFkruECYdHVUhGtNQDrzvK28uBZQRM
z4UCblcVv4TDdQywM3jps+CId5EhURxBSmHIYA+dDHSbYWbIfQIGyxzl/txFwk53G+9xld7AEMy4
CRQmD0djB4n9S55T3SGsJTO/kvzNRLovD384+DqMGmx7yMr4ihoVMTMttlBzKyNjWGtJYnhJydLu
DYIRy5mXT2WvBhlFra1bJZqntEYkCSXe3Vr2vP2Uc0I4NzxEyYJS6BCYKRFp7ZcMJUZh/ZGPdvxL
inKP/MOfNljha5UP4/6RCQ9Wk5tmXmfxRnnTZDI0CpHVacQuScXsKoc14Bk/xHorAM9gpIhB0++o
5uwVGJc/myt7+cdF6OZ2UdYcObsJAP7fkOwNezzxBHHbY6AmRS8RKvuqufK0xYRxm8DMMprjlKou
V6jIlorSFdPxnV+saxBSETN3TPcDF9jKs04hBgEec5vHvHZzNyxrEJ0z0H9l2WAkxNomPd37VI0l
xSwzurA/39qQ8yKljRoSb3kYicw4MUH9UZByR+cBxaOoFP7RA1c/QkCrRmr7uF4Dbzf79N/JkaQR
GgRvWjJ+dwriUPE4H3M1QGF5lGKh74i0jSQ7TiwfJw/NhwiFMmQfkUkP7zyrKW2urDcqzDw5o0TJ
xQjRjjnIqtaJDCVs85bSO6KEPrtB60cFOV+lDhEmc1a5ZCnwMY2Dn90h0Dl8sn/S24hmqJy/lx4O
mvhPDwrX3+6Q1ohcJCSbBUgvz0Qbnf8KRIL0V6VO+dyQ+/7L+XgR5lGKXUL05SoXQF76y7eh2djc
MPTOaW7lgsBt81GAD1TGSgS1nsYBDOTXtK2179Eakqng64ylaSCHXlEk5Fy+QuV8Rj6o0jWNX0od
0nq9GwxdMJRNsZvNz6vcG7YFwSLXSHWQakFzkOlqbIG8dRqIIMjfDwMIy7rXVIysLBI6kRWjpvUg
Oz48DxSed7XNhn8NT2kAJmJm7aj21uQzABB19oAuaWDRXFpQbiqyDTD/4VN3/6au6Sw5vePISNBl
vnS5cb00FMiGgUbHnSI0vd+87eruQy3hrnbdtflq5yBoyKq1w+fSdJJFHFOwHEV+2Fe4qoUqaRue
pNi225Cpyh8bU2NUxNccNnHDll253wsCA548S2wCKYG1uasbpddSDxtzQJ0NRZVrZo+6mi/NTxkW
uFh1gVE+BzlV0EJ7cFZ1oINLD7pP5U8hOXcEoQl+qxkzAGCBz0PCbeSubjNGs0H7iX9CQ8oZJ+T6
Ky4XHoH95Xyndu/xqywYeRGyWy1xHPywKIf2lObIGKR7V/lZEH8o8vVWvCFnbMmSSsm5kIZWg2Sm
e9MvbXoL9BFQ6mDAjnoW7u0vGLE8uNINslv3AXFeSjeDlO70YpfB21NvH6onDNID0aMfI9QqdLN0
pBwPG+ul/JkjiOcrY4wNgM/if4u+A2ehtiFJVK24vlN96DPXif72gWXH2qfjkDDMhL9WQGOPd41U
ZzaiG3msebvLrqFr5xQmRHyP7Hl6h2yKDzGNeU5dofj42ItjDIAqcfZ98Qu4i++eKq77wnf+wkRd
xzQy85my3VJtr98CDG6yBrcYdxJLyHQRVgtTxQLqCtcoiSEZ3Hhwrk68KuMPWnD+AyFSkyKpSsWU
01xc5v7ycf020NsdY7RQEFqHLFjsoZ2AKodnH7KmpJ5Nm4YdvTym7aJZ+9KYR27MyTenPG6ZbHd9
mHdF45tUjqykZF9AiZOZyAud1gjAkF88qg/3glevdQeB2tpVdUkrcByvo9NUcwkKFoK7xIIJpmlW
j+S3y8gC8V6EV3q54852cKVwwalE6PgBu3S3gA3Xiu2t20OSX30lwiG41kGcwXSSg3PUSa3sk93c
pRWRRYuPbhrw+GG2Su/er3FjFyNAyeVTe8NOdDO+hR+zgeOkTSawpB/45yTfa8jGDLFpmJ+H3Em1
DC9MkgzvgNAVEShDM6pMphqTmHISU6URia/gK8zyQprNzqv3Z1mcCZJt/4r9E9Wau8AnKoFCwGvj
7P8Ag+qUOg64O1GE1rvp+NTOeTuJcGXJsIKv+nmre6idq9a5/V+OvPLj2+SoJVeYrdK/CtEkBqei
de5YFJKbVOUos36W4tnl+yDwvs63hk4Pkfi0NxUde2vRsrMM+XfN2F7fGpCaMOa0E7WpXOYuMShW
rcJaB1hNZOIY4e75ZizRCa6YcY/+yclspiG5ikMGLFY6EZG3y5Ng8GFlDclAsdNZpy2poYesjmfo
EX+7xxbkNWs0wT4JIf/2HobOrbLvCXWeDXFuDijxuPvqlAjDVtDJ4bZ0Ovh9MA04TkQh4VrWfO1i
Jf1PnLwHEX4CeHI7HPuLbZvDxqIEbwJUrYi3VlsXhGHRX2az0WpYrBTOQjDObmOvYJCN64WLwwMm
pr/qhA6fhyk9zdjpW7UQriee21KWURrN4PrKj/G41ZS3zVkbTau1o7MUjJZuhDJdaNjdm5DPXhzA
d9RrCzYomkQUz44qpbSceAJ/ld8+8CX5ISWQ/IBdsWOU8IErVpvcEAXT0ADXMQWh3BO5BG+FlLZM
hE/i9WziKj2/PAO7c/+7yoZTOT2s/nDCiYMoIUNdqZHNj7voEFK3NpyByFSJE4pB2XFcchFKnmcT
041E0A+BM7ig98o5YDh/0euVKYrlu7/Bw6CzpYj/0jOsQe54J6yNkwHnP2kScfQlwXzcrWqdrVUd
gqSh33tb9YWYDD6HvbYSdxV53dICkrGCeytBGk74LhQxBQTjrHtYVWLUw6O8QGhvRJjhiuAXM4s2
IfpotbPqmOJkoPceRqwMNeDYV+JHmDxHDin+PERlMbYFLrzb0hU11OkBg4kOlMI/I5FNMyfuczDt
tYrPaNEqVUVjxpvNZZ7e+ZacxB2Q4y4hYuk+xPMxnR/SmA6mJGJxKbQswrpcWE5Ajjq/gNtzZ36E
9Z8q5q5z2oHqe+L0FuOgdC8uLQhSZ7a/QoQvxyqBueF+QHyvZ5dPhZd21fqXwrxZHDdRQd9zrw2o
wHunECy6WjLLFytE1gSgODg20dpsdcjRMTbWI7tU1+8Mbyh0oesy8Lt0RQEnTjbHskZnchI3pILi
2tw42/1ARAokrsKRn9quA0ZSfag5I8qg45j3UF/Jw83nwsqY28oClmq/KXKQ0+VkRLwl9aZ9JJuB
+bU7tjZIgXeKV3h6N+ujux4+bLhukYnmB9EgKIa/NJKNKXBfJuUGCOI6qxEBC0OCoR9Q8xp2OV9U
jLUNXHxGUfIGTUaYbz4AWXRwfJowsvCrBeFgNaL9zDgunXHeLaky3mU/WfK77hSYlCTWoHrpGH6W
tyFtNqA7YpQBRN4CyssBa1Q19tjw/T5T8FlGiytjbues5SF3UKK01pLqErLW1rROLtRmDAp/DDnS
43ADDj1XffLBhRFclHnJMiR1lvhrv8rroU26goSs+/c0CxFHiQjgPmHGvg4zkuUeg7hzV1vBl7//
xOoTTq2l/B3S5ynMtmqdPdmhwFFg/3T0zY9ES933k5y1xUr+2F7w0xC1LadRnZ8VTVpq2vMKJ1jL
uagRV9UAXgbNmnpeuGEt45HTvuqC6HtiZ+EcLbrh60P3ru0DpUZkYIF9lImD/PliWHxNDFa24ENJ
A3djbhMYEunebdjywiFbpJaN/yDLP6NhYLVadEUjznRPc1aEo1rygOwpd50vhwbDDTeF8FKg+bsx
lXEjMPfh/t0LHj1zMywMGNa1QE9Y0DR2NleCUk/v0GInTg7mmmiDUKKVMrB50p3YStsmeQq8/oVa
a3KJmo7BY7TS0J8ZRTedKO2uv1+INd9KTZNCEENGQqk4JXSZ0YNJX+A5PZI9b2Rz7hNwCVxm9xiL
5d7COl91PZ3EuTK/G+9fevvlZ6dG+mMjswZoXjl56ZhYlj6BWuw0Z79XSjQrUFQW8kGvke86vFhY
rjnhsRyEnoYLxP+7En3V7ADO8iMxNHdXR/GBCAmKtEcxeXKZzXThfSQR4ljF/L6vFgI/cYCEzhDU
+4Z7bxu3IKTT2TLsDTSreJhvQS8kGqahk0H4G2D7Sh1LH03k8S+sG+FMhifIS9c/NItXpvseUgd5
LXnzBlmevTTVhPPQC6QM5c7kzCgwih5oSM607abpFKc8w24s1QdKSBEq3X4csCr35cxtfPBXSUT7
4HY3rz7DzMpB/azlm1LoPlk2ak2guWNLtiEbd49mdMKl3oCieSzqttgSVVTsJIQ3msfaFzttwI3o
8EixnivofqOQzdaTtxE0qTrkSypxb0bEFoo6bf/J45btiarmoJJjspV4/9VzoEAfwGf4j7LaGW8X
OovaRg4cgahAR8Q2xdsn8oW0P1O88MAyXBtPw+zBNqCI2I92+bo2cBJ6XT2CrnaDPXadm75lNcXy
7X74YH1UyZO4C92iS1QY16LKlvNf6v9Lz0ktLfsrARIJP7PEdHkI0WVAp83LnHVYojO7Rbs3oyrr
Ko5gfL9gRaD2ZkY2kQGJ5wi9XNz+x34exgzxWKb4zAkgNV3wG9tps97DpFFjSvQRAegJSm1kuGbB
ycLDEV61hLCNZRGUl7dAQ4vepLb7IZpxkfGYqSNYod3dklSWLrz8k3MM+m1gWm3XC6ZCJzNUyF3i
VKTfuIvNEr6Klfa/WR6skSyhArnEYQcY7fHAxm//EbwpYF+NJhZdw1Dy6hi2cjkUM60uWf7YzmgG
6uAkBVLPhnLpNlFnMlpe2Mbqw9NQ7oH4fJqLgeADCvL6fuzNxIl9S+umQVJ9SKZlU39NBv6G50Oz
bTx1e2G4ea6ACkaCoPIUdlYcICvvEWk3xoXp8F/h+OOCru7sn4tJEUWe0rJVftJBKUvcVOFl7684
YgC42PpBzvSDerE0/9+ca44FYR5NLFfWHffHlMJZaNOYgcLXze+c4fj6Uq5Z901ItdVCI+WBSeNF
lGoY6GoeTv5qJGpAiY7gk8/3EnzV/gL/mkaEwaPdxWjcjOi+g/f0tUcUjK7T++yo55q5KZbTaBzO
Tc97cIPjikSyZopLYVVhnDQR1+f8zkmEp/KyY3JzeeP70CXjmybR4emUmQ2wogLxjN903XPgCVd0
xsf/2Jo64xiENEOA90b6Y9MXrO0cBG659XvglmMHsezvKhebwSJ+l/fSBNyDTC2oSdbyJoaYVQqM
YG9ClFr+bSDaX1N79yfKMMQRc0rBNjexaLUg9Ba6GIYkrSmr2l3raIU9RHWTZnbdVJp7dWBXx9SM
cns1jD1/FUH5KSyUugrDI9OLZIoFoPY6qCPhQoSVKuLmnoddaS78up0KC7BPsgQzZT3FtfALHLPD
2Co44HkDx2Iukaxk1Z55rTtr3B9ozG7WjRNpuERKatvCwTt7fXu7u/YP/wfOzKL4Co3jRJrxhY+6
albdMczPdyVaoPQzCburvXw1SWTzpbCieSaGEfHRuVW1pg6atkDtzSzQzhiydzcYAgZU2KMuOkVw
LvKwSOxxtLrDHiSLrLXRIl8YJYXfcbX77OxcnpGd12ISsQVi3gCVqjk7yBQZxZwh52piG+bdIRg8
wWpECibmMK3qZ9N+k/PlTnJggPpmQa6c+8WDVj+n52f4rJc8DzWUZ+QG3mi9uOHxxVgHtMNe/sl5
JikdrpsUM6lZwz0VpVPL1uayDe6+B34cejiOyBKUIKMOlohhYDg3bBO6C7rNhi9eaa39FMi98E07
vxwqqhyxeYw9EWeFCp3oheTEZ3Bt5Dd4IN1sJsNauQWkffyXsjSWj1PLhQrfVZm8IjnkRmorYnIR
eyUFmXE6rgi1t71qNcMTyr4PcU2cuS72U0SyMNY7NeBmpGpnVUJVGqlbVG4BWZuSSPMWHM0RFnHK
2YkgQnlWgoxZRmatpbXKkRMVFHVe5KSdnWWG5HriKmIYnw1CVe9VsVBMVUi1lGjQFnBCjS3s8b4L
sfeV9BxR1wofLKaHJ/5CdTqAFJXT4ydns0lHyymqEwg6Uf43U1S1eGIJozIHqFz9RsCOSqOlQVGd
UbNCFfrHePG9hdyoBWJBgs9/Pf4Z6FG47Nvg/INivT4drjy5NUOIfidIBwXlYkLpVAq2J/bpjHV8
7g+f/KnhpGAZag5TgS8YHrE8GMLSjKd/T6gQHjTNvMFeTur7Bex54AXD594ZS8LXvwMBdDbLyVVa
dsR4qsyLjwT/cLCAt73k08ISeHPoC13HDy4LHG4hgL7rNM7/2QCcgDJhHqXFm5T5bhWZS5r2k/6b
P5bYWXHkt07II8pdp/+DncAmIPfSoh5C2up4RT/8efHZEG7cKO4IOfG3VdPkGnToEaxBYJeOewr7
chu2AR1Dr4wMk06ttRexgfoZFy6H4z30iQuA1xRPaiDPczvZ7D+Scos9ySFzLgdLhAUH1VYkfZSv
2uX0bLnqbiIpqNEglzMSa8vkXOUzBOFDzYtDW5BEcHJqoRk2SDrLWBWVPL+IwSjD0sIdffOwdkL8
EBqDg5xyHeBsW31TSUVLpiG2gL8vnhP04l8e4uTKLbR0WMTzpV0/Fpc9XZMewYLiwL7FG3iLC+1r
YvC2e1mIX5uKfnaA3GS/jbtGUdOg5xbVgrLCYsvQYfX84z8ffl85CO48A19HY8ZnKBc+kqsv9xFU
+BZenaKWTROB+7JQmBdoQICeWZjGiusG+mDY02tyTO3XQpIOI4sXcfMVEH2WyCFsQPFkut79MKJy
XT/9ErrHhEt2qreHI8jSaWhVLim/t3NBiNjViK5eHwIGR6ZGX3uShSNEU3L7xPsrhCBou2sORm0i
c0hGf31kmqOC+Nmuxe31iojaxExu0bSWtyaMewWV2xHd65r2YFBkRAvb8/H3Q5a5RvUvQjZmSwXh
IzcAx76iOI4HF3mqqwVoh/a2qbdhq1tLCcIRAZVL9sv+wrMn3w0HohRXCRAV9MdOP5196vT7yUkN
GWasTN4v5y0lBHsTGT2K9k3G4aG889oIYpnk7eJjYcEx9CwjHrKA2pkfPnjepPk7VuZBlB4EfLzs
H+H5RkZfw6n2su7BAx/Wx6D9HtkNYQSd3QTiENKJIc4jIwkxOSXuuoWxX/KT9xPzZhKLRHzQnYz5
fEVa/wRPi2Bu1Ci9ChZe8KQ/KKREd230jBE0dfwWh8oV5sL+lgnm7xCjC7/WjfI62djSewO0gi4e
NIg1VM6MpN+qDnFajHk4rUI4PmmQsjZji3wWA13WDzKWiFZHcVc6iIvPz2tnek+x/M1R1WFEE20a
Q7cEN9k4oqAJnXlh6pP6Vh+ECExy4jBTIODFMGc/KunBaTxWDsyU+ARPgMd3FyiEOkQQd/NdOQ57
EaLu4NdfqBvCMh69FiAikQJT5031nKg2qzzblY+fFs0/mIqqWLvUOtOw25BlyH+XwxG5XYaz7O+8
0wFmYPlPGWp9koOXj0teN5P9V7vz58QCa44Pv41Al7Myk1Hs3hqdyYUFJzgd3NCULIKByGEZmq8s
SBqA2LlQpc+Ls1mxSyhveMTnhY2NLYJS5q8WdwPgGYArhnX2SNZ6dPolNYTMvpDwchZk2zxRWYJt
GKrmX+PpntuOAOZ//RKmf71Fg3Kgzdlzf0Akt83nKXXFhh69g1spVjvQABUr2tZY1pvQy6CfccpN
vxs1+oHkx8wZuSbIUdmG/PU7U1HdtwQuNaVqPEqtt21Qhn7Azmv0U8WrZLqdL+8gbAneEIKsQNmE
QaSlTcQqQUhq+fzWnOznkn/Xcel60m/EfXnXm8x/BBdFyIRjvdHnj9E6XMQOPzmVqZDsax0CDwC7
vA5QY7to3VL1KxXqS/i8Kkq6VmKrRoQ2ysfxW5Vx4gGGmeS8hUHeMgmo4Y4Q96PIjoVcn2dY0PG5
IRQHxI/FoEOaZC1NDyhnU0MJoFVwYK3U4uLsSJjLEEc3oDOgF0uXmraE8zPBlIpRf8VF8hY1f96m
cn0nwxbYZM5zLuxwSJhwfMBASlkFI/OCyogv7LhDDC/q2M4s0ZVMpprwh0yiCnHhnPTyg0ZV2ldH
1l9DqkfN2SkiQVr/h2/0zf8qmqjNyeUCydAZJ3xQiaNZfs0evjrFpj1eA07dL6Ox/iDY0a0seSVo
2zTJ0Yp2FBY1GRd0C4GXYM1IclFue78ZTEVYPJOsI47oz10AC2s9gk1C4X/ZTv9IboKhNSgVfTXv
8iq8nZJKRGP1ycVjXO2SwEzSZVLqFLCUjhL8RRMT7jZui99T3C5q4TAIrC5SrUoa4LLtn8XZ3Tq7
VlbGSoeO0k/CAp3aJ09XrfLjoGuwBHKyjj/VvVhZgl1y4znY2iTAOhbbQ4kgNgud1SDM9YFwrMlC
mSw5Bdydyc0I/KQyTexxcUO855wQpAsURwT9c1G3z9kAbZhU41Kn+UpR9w5PN14+VGi/xbKpUMLc
ss1cKp0vyf+Vzd3PdL3cHYgKQn7uJQxcIQRuDpoBXjFXMutOTuAUIUk+AWa5mt4RlFjUqt7//7ys
+SYv0xOS01g0cvOGy8p9ZjOqrdSYcih/YcuqGM+pI2fonVm3DU1+JPTaWB1m20/L4CUnAMWENWMm
SOclq5dmgPWolM0vlPE34aCzn/OmW8xvbBL9oeShvLPINr3wRXx8+QZPd07dRSUV1tuPtifUveON
nx2JHJkDpXR9pu6fnZtXmwB+RnTaVuBtv/oEFokzqmUOo/rWWEg+KqjmhCLtXd8u81YFS29aCKG8
VhSB5V+PVWzcahQL3r55CU0C4SlygdQLaK29vjX8zMmA8epzBOfHMmOV/KzxzgXfQO8lEGeSNzOt
V0vPf47tTgruIKDAsWHPT6AiG8Lifp7byrFuIDf01Rb+t13b9wKOrT0FjZIl/JgMOYZhc08Ko2EP
THiPwR6Wk/ExkoWLXsR9Nynsw9jYCcKbuCmrf5O7L6InoaiNKRsG7+WAIg6o+qB88g2bXDlvMlbT
Jm88UuTu8i6ZO6534lIKVfLYvjeBdXy/4/zl/EpiJFMsxB9+gzNEJBPZUvAeMC0HuPUuOcZki4h2
AWWQRHAX51SsjiIa7JztQc/C5XiD3GFiI3AfEqsISw3SK8a3TUIS/gSX+e5JVdXeGNUJivB1reBA
qvyLhtEaiPWfvtP88xQeaqa8TnkKl380XTxkf3XK7SlUyhvaBPkF8WvBlN6Vo8TaVYp5inXBIAIc
KI5ufn7KLiB4HAf7yUO6Jyp6WBlj28lChT8rH6DJulFDeXg3fpozws+sztNPrTAl8n84ugYoYWcK
nJGvjLuU2lwXvbAQJO5IEzpZh+VdwO+rhUo9F+8Qxbij6n9CEvagc775t56E9Xnwrdls7BuU78Yk
+fIhHzdzoBmnu2Dd5i2hBd0aYJwjXyHW7/+vh2Ik+CsbthB9OXQ7hMKhkzqWQcGoU7VQ/MNBaTMC
MSxoqXe02nGR9LI3ObzGgjU4Ts19UPQoNGVBmQW3MlKqR0phUtfRNt9vDclyC4A+KPScybirf87u
zUko8CploTtScaBVqCZYMmD2JMLnErUOSTkZf4vTrWKtAQOOuYKYvNGJRqawdU/2ikMdocFSR0jB
SJGidFSPJEkRRf93N7XaMe9trYQ68k0CBqQ1b0N/nqvQOvIR6nXw2bz95ee/6NBgpxRMNslzZEBx
3NZnEhelp15yy+WGRk4mqlSFX5P2Ri+sAqLBtXI7VRug/foupQB4LSL+Zb+rFoOSTHrRFLf9r7Z7
7ar7OLzbx/JSWCxOQgt9GvK1RgKpK9O/fNbEPce0mr+VEi9MiT3uQueKISTwj4WybcAYSPNz9Ara
ql2DbS/f7OFCCWcqCltXut4xyQ5nUKH0mPRcA9nTakOQGsfuJrWIssJLuWwOjlctUW4+GdDn79bk
hdpqL3cuxUvASidXiXnQmaOAwF0GlgOG+qv9vpItTxGMDVbM0K5rn3pi2PTSL1BMfG/DWDbrQTJH
dgkisV+i1jDb+rv7qmci/mHLm01o6TzngBhxjdDDz5I0YExFHP90cSdMFm4TzIgT+nF97wOOk8VJ
57WAy5N8rBYor/j6pIU95lZ85hRYl3dxgB9irf9J7RfEmCulXji3RKXASwKr5i2vYFBpteWKMIAQ
hosFonwK5Y+4dNJdIJNWk0KmXPKRWTcvtwbEI9yeKwIyHOnlzJjdkw1vu/XR3gD/lS5T0VJ1+Hl4
+pl5+ZaDC7PiDkCIlUAw1B+G+4ytkGXMj6gokjVdeK9SK+RIt5xQZ2U5EijzJCt6DRYquCgYfqVM
kv4RUpYdmoHYNG+qskidqo6KXQ8hY8HaezB71HfQ7O9zIkilRvKti6mMgiKMD2wZoJA9RtxfQQOp
Wwfeec60LaVFgWmG1eL8YECbLopLEkjiFPoKlnAg9h7u2kZPW6lqwswtmD+rjjNUsxcpTiSFfHYY
blTBpoItavQ5cGv2qicTYFQXPYxMZ8+u8yQ2r/FpGtQTIVMk2xZgJh/gJUfdwETRxPZZ9XVzcrqG
pYx1zoxfzMhb6EpXPQNNV2or9Kk6fQhkpQEiQ2UOjGHp9YOGT+iUcse8LYECeB12xSpw1jrcl1rn
AcXxQeUMB2NGFCz8SV+ghdzKz731ONY4iXUDfu6sWutbBIBzfk7P6zYFa9krH2kA1QlhXjdnOKhf
vJOSuuZuXhfQH9Pdec2eSeeOX05S8g7HHD17UxK8zzRTXtc9SbkVTNELZMSayi2jRzpObJtDuXH/
LfQKSe6JCljW8263ebDNIbDrw/HaEeE3S42OOXvnlJkYONj3HXkZZaeIliWGjLyHFNyBryk2M3hF
GBkag2fh20wnbJ4d54eZxUSkt3GNugTyQUhtgrQryeKzcZhrKAbNjZ9ERt+tuW82BajST8UK+L1C
TD74Jei54nf2574+qTUHuwIRZn5rtn54rev8CmrfeaHINt0PWPEpkbPhKLvE9KUcuW5pYXm+NKV6
57X+PKoYeCQ6Sxf8yjKmBgJwLS7jT6EhuNd6xVLv7L8XClmOBfOKQ82SHMCdrGxVdpsE04cFeXhS
nCV3RPmyrODLmW/8DzqhxKOo/3P3kMBXprxS5U0a6G/Rmy7YRtjUggiMKZWx7yWtLhxgMimKNA57
tcMI0vLS+MP81ufzrAXNhq76EyqAochLD/jbnsNmFmCXw6l8AQv7nRULGDubbKq24N+qLJXh5B/g
HNMTMR5gjZFJRAA9fMWySHIHm8Zt6PRkWTSon2deKy74A2+IK1F8XslGARqEmv8eXHdwMY7UURNQ
3beg3ftwyu+DhfLL87v/yPVVl1kLMNRduUQfWJsVlJNLHvxqpQY/fY7KjQSXnu83b7la0TeXDlAL
b+oOyBsNWWxRBliN49XaibiOX5gq8PE2MqFxb6dimjkvb2fMQZOaQJf7KZ7E5zeebyWt7Fis3idl
KGAIj9MZzCiVEuQqYP30VXzB127LAOkym1aBYrsV7WOrKYSmsNgk73C7r/kEag45d/UgSurP0q95
VMRQajHFIDn1yQsFtmWiafx3vNXdpy6It06CsSRHG2AjKkseNugG6AtlaHOTNB4TjRjZdDKQcNiB
kExHPEXdq0GESMg8N+AxZvwZ1B6KYTfBgcR+d5npJzevFlMaviUvPyWEDS69gjVKvX4JS1F9uk+B
0liySsD4qn1VV7StYVfVssdakY10QGXinJ8T8Z6wkmUSI1gKf/AwWtT6f2CngLptU6u2OiYRmsRM
DYkGmLX9ZVQwKVB9KV4s899ijSlDCNqxGkuJEeWqE3UCeqA+2eC7YSGPyRpEMADSOLm5918gst3h
gk47GSeNdpMAKTcxEu3dtzPhBd/Xz3qGF4C2vTw7Kmc63Qxp1ZMo290ZhvAhYMwR14E5c4KW4eIM
7SVh/Eb7oB1EX/ExifxeBIzu8psxPOPc8QWzhE2vvkowzU5Sku4YEnQb2sfpENTeZ9rOET+nrZmg
Lxwo2kT5Y6EHLQrz5mHf43okH6/l01beOKwVGjvtQc5v2qVxWywr1sxGXDcqatNfCZxIWaQhdkwP
eGxcBM8Bsgl3Bfv5y/tDsuo8C2kSfDEPYf+Xj+jU6XaZsu3bnA+FGFTfUxMx8bUWjCBTL++OqJ+k
0iSY5ZAfCgyX9vaQLeruQLLchEt877nhkct63DsJL5MSqNYg/NvOAi/46XvhRFnHleqAyqkylwnr
i/9DTG9T9V7rscoXnTk+OlDhJj4C146uNWqjxRwst2/NknHjxnMznWbeGtwZdaN+a2a+4IaBb+YC
lnugF8E/8bPHv68fHVNJDNVkpCZsXuX7Ud4SP1baneMJZypjHClY3eWDKll9X7c4ZcG1yrP+fOfn
3yvSUrG0GoskB65k3r0eWtVard+X9qvT8sRavjYeiSf9AyQTaNMLBXoBtLoGco2GtB6PCoBy4Nri
x/M5MH5eyukZh4bT03E/Ilb1Bsblys8gVTE9JswUW2V8aU0hh5PqXI8WBgi6LYdvXag2683/xY8x
VY/buyr/JXGjy4MVyrI/aGbAqJ0ZMDR7AcEIYKq72ENHPIEmBvSq951LnCuEhhC40qtF5f78t+V5
JT6BTW357E4dqCfgQXaJRlPfqniIuu+r2YdW8b7FRux/mbu9G11Dyn89K91tdzbnVv4dqKPuGrJG
eP47FA6JUDSAXPc5d8qyPudvuTa9DtTNkwRlahW4d4C5U45eEBBIvjw7b7+iG1RbC1Qq9CfEaznu
yrAAcnpXBIU54Vsb/KltT1ph0jT0UQM9dAM2MCHIzW5fZ0mw1JZKNmB9jrE4N0b4Y/jqSXirW6vP
TncTdVEVY3HxvXuVlJ4J71wxXBCsWu1TRcO8Bn1Vw83F8sJJNaYO+I7Wn/rPV4utIORR+OheM+AG
x2rQ2CivjLYC3szED5j+MrHEcHqSgCj5WziowpIkwGilqkOZQFgYpPikZU5fl0WevoRsDiKGl1NI
oahhkZLgt7kxDtYSAZhgQl0Wqmvyb+FQbNZON+v1T2eK83ukNOwH1SaJGYCEtxSDfBoCL5bbI4DU
IStWXE6+B+C8Idpm5x+JLA8oVPbtHtuWIMnkSmMQezxGJ1N+UBg7sWomOvIdeior+jxkhyUXTLhj
9XP/CqvjzNVf3vLBG1fwTIeNP+6dZ4fcSFXQ4alDPYfQ7TRkQYB3QVnGoLK2wk4P0ZyxINAu8ojk
nqBjVVc6PW3sJP/x/diQx0uWiY5v/AIkkoF6hh3gyJefp1cJG2thi9Q7+6ptcjGJm//Yl5w/jr1d
xVlluHGjPHDVzzDgWAvttBh+Kh8PyHNPTFak9JUQ/8ldhRcNLkvXP6Vpyhzl6uNbD71TDNFQsx8E
gQsphuBiSrzisOOCFXAs57Tj9Z3pV5kQHkWqBcYRzeGa5bSP0bmHqowtyIhMg25oD5VhtraNL2Wj
Lf5DTX8h04EbTf7NFUcFY8v15ysrZ6YNFV4pwJ8nJe8NgFC3kFMf/n9iKqZnElj7+QkM/bv7jmZ4
tRA0PBOOsP1bty2Gl6s/u4OCqPD0NPcuEaqBDsriQmEulge1mqzHf0Av4iU5HFsVlo+L5WVMG3WY
pE7yDvYhsNeNRbFg430YsPZTFxlzPRxPz/D2/b53ucPmRoKDDV5IIu4HnFL3jQcjwW4w9wobnn1i
5bNhxxE2fBBoWroEH/Mx10poUP+glmnpDK3F+9e9LDoeUgz7HFnN35KQ907Wb/AaxoBXyzTmYE9l
y/36//QmdRm5kRhN28p7GdO4EeEk6WjjTEAmP2YwDphyCjIo6MWZ55jJzPt4KJfWyvZ8KDzINpvJ
pVUu/Sc3BSmY7Yr+3fl5rjrcdrx6nEBqJ4IRTp5kymxdpGOLjqPuY3/Aehkv/cHbPNO1aZjMbIDl
5vJ9h4WyHoiyJleAbP3uVPz7h5IiNknf4uPcdPe0LoiypjOLXrBEX8MTQtBmgy4dMJAWT9PwTZF4
41d6/cdDHsOtWxIauYnw8+MnK03MxPXCGbAPtoEd86JQAOO9YK4RASQOZZiw5B0p7bOAVHPZGVWm
Ue4Ogm34z4fqV01NHJAnjbPHFTZlQgNrS8pl0qH5YmFP+jd9mA3SXX8xl4NFWGP2MCTr04bE2UFr
oTtC92zieIGUR5zHhFCp+y51bVDnGG/zYNvlwT1KVHctvp0LM3+VorwP3UpQaQK2qPhrP6PCO/sf
P4+KvIZqsISIuBYiP6tERMDx8exFVEXUkZJ7DxSOi5f2qEreAMGiSKplUviMkvISxMeDpEysOgao
+7SJjOoudqhHRoOtDzlF8BxWYqeMS8lCx7r9ZbR1Qd6BROmLw1yqtqssx3oL1GK8vwQHb8SVRn6W
c8vq2pWfZptaYQG9J3qEsp5qIb7Mfg1mePdKH2f50kZVDpHBs3gxRlcD4IqqWjTFmz9E7kcLRCVH
l2j7FfKelSDfbme/NDD7JHrUL9Einv8GXftg3fvI+7Qn7838cGY987fBIN4vcADSk9LU+PqR4DhS
YMSsc3nL0uhfArOrrC6DtuVI4ExsJQP5Alq/zUbYB2grwnmN73MUVeh1LLrMYd8WcXbSCuSjGIuk
Xo8/IUAKuXLDaVTN6TebQEWpu41buRpA/M29Fh8Oyn6gcghhAQz33IxIo0eWHkJPCuJrgK9WaGht
8wARPlBohS9FF5AST/FUpejNGawx5ueW+RpzvfwIgJGurfuf8DikxFUqkkI3WEuWq+6cMvEZslfq
VN8u2puYL6oQKskJleM/ZUTQpYhDC+aeC+jO9vnD3KzZmkF5DtEOkmFwIWwYf4AsXfRUtHcOtuBH
bX0ju0czPvH5swYPnDYD308rXGPFw4r/APfcXCq3vqtBG5biKLEWQFjV+XxhqC40Tnfo2Bbdim/V
xkPQbzY9s7h2fWK2Eq5cVxcMiUI4eDXuQ0n3n8iKH6kxbLsI5y1ieUQZ+eV8pJWCyX6mF1OECApr
z0DBqBdYgV14N6uwLV9lo4zSiy7YcgtvM/01JrFYn7YrAL3npJ3wfna6hFxguSdaKTJVruUDzgZf
l31ifwcxMe6bFVWVuPKZYMpJAuR4Ye7QdNgYGwvcIUjj/m5wYM+fsfg/kIg63uvnLfaHmUbbmhJJ
6opAcjlU7SJkYQ0bJ8SUQjzn1kqKq3cAY+oCEmMj1zB478r5u3RZNjk8YzLpr62RtDXYnPhY5z80
XQ/GCf3Cc+9oVNBohKsvr6QAt/4J7l07bm2glvS5TEgrM2NZ7HhTVtylQoK4LSUMMiAo3PodIpZZ
od4Ub6tS28PqK5soDzMiwLqfohSpgpxdwq0AnOEble65sA8+oU4QtjZoFANk9lErSjZg0w+0R8hk
NiNczt32z9NkVLDtKiXj8xrMTODlg9VYC2yCIQEY6ZyziOtVo2W8P5zfkPrXZieqIeyTrJt2G+wh
N3DbE2Xl81uJAnHtOLoEtYBVgY/nb/B1ZNb/u3SCgWhfKQuSdgO3DY4ivqHNUfdG10nHenX6F/Rf
3/NeAWRSkXH/DOBAa0gNL86YWRPz6jqYXOCmVxYxfBjSS/OtDlG3Oe7okX6nVZfZHHw4z15WvU6S
FDiNZlVI8VcUEcI3TlLF/u47Fu456/qPkT3fHGibCpiz3dUDCmkoVMhWj++mJe0BBxIWNMNpX+nW
jmt9JlTZLOu2UjUU/Z4903P1bR5OJhFUdKHCOniOQhpkjnG7U3v2qHGPtVoTx6B8u/RE0J3L1kNM
Z9vB4DqxOVGxJGa1qb05ttrUTzAW9xwzeMQRb2kXlMnwBuckzafymxq16EwfEvvi9PpoEvoGbwui
5EMGkI7j2IMSFgbNFgIuJwCrdNAl5No3jz4tmlwc3pwmHm7P3C7BQkmJjVXUOdAW6sXiJ61n3g4w
agQerCkbapwRtDBOoac9KMp/HJOE0XNNoH0A4xB0OONnixwtgNdVZrJXP5lCC8QnTJKXbEbN65zE
v2FbOe/9poZpUQBJwtPNWlZ4kD346ejtyiwkbrJ4z6Rr7iSRahcwyfR00PopfkULXT8OJQG0oWfU
ZjQCRs7NLIN5MNXNVUojdbsVDC+puJp6pMMldnsIbIobbco3lCppOG2tTYAQ1f+uhvLIt5HjIl9R
2bOquk4PGCdWNE1lnzmbEKVlsor/dagxGi8VfrMzCVladgcl+7lI2gk+YUpdANzDfC+CMDP70S0R
2zahCMy8haDUHrjsksqf54ZYrPLtVricd3+G9FKcpHM+6ksw/yL6pH0sJu1rvvY2UY4MwQ2yfhcN
BqWPfrWnWul/zBHcE+mcI9EcFQBLCS+D54Z7TNFtDGnK+OLQuh2VZgP9SEof53MnXFMxk7DTdb54
RswWLdLqoSrx1WVSeLVL+kY9lRvs0Tc/WtI19f1gkT+3eHZXiJEHwST6UhUrhhIYBmyMUsMEO4vb
LvrKdmgDpop/vTAfG0iNoSLP3BLNasa6qvEfD+0OMm33qqmBJuVp2FcLct4T7aHwYY8qGUjfbqyD
e6fJCjMrmup0sJbvW5cDVJ6fjE60jFs6rV1M8tJsAO9czP7ObfnCvH8Uo3ycjC04eq+hELvI1k1k
felx7qeY9IrwOuphrgpAf4N+ntHv1Z3dubHp2QUoOU2ktrwLcjmaJNPd2Ot3xEmr3hLSd56mrdCo
swKSFNOkWbfE8mYohW5PYKGP/+RW/+OE4FAj+KgHh1nf+BM7B18nX9l1Hc176KyGkG93TPF2ocYs
dOlRVFExjHZ1tMJNDNHwsXTQx0ieGGBxqt5l0v5jUGvR2MCQcp9PS973xIYHlWwxoytor+xA1c5O
E306Mk8Ftig/5PQRdjRt00v1bah+LOE7KxiBzuxBu6r8ycpBjzbVOctdiDSk2WDmp6Zj0QXVbh3s
35bFgXU7kGzqFDh2YKbZ2xe3yocTeXdAoDGD8MwahUZY7k5ukn48RdeTXsVy3JpfmQr/x1zbQBTV
3IMxzRwVpjrtUnA3xWYz7kXZP+0oyftvr78NPZGPu1oFLbpCfSZCcy/WF8noT7uphhrzJu2AAmts
Znh3RbhnKM+NgLf+T4Hw0ykUAZxDdGAIMnSIo4JvKcmyQ2uyEB1XM2nXcezrg0ilA0GsUy6bX1+L
dVE3gTJpQTHpt06Y2G4y4EDmg0E7bi/81qt2lBTStawzO5/Ym4e2QUx09btmwaBPH0QCCoWqYrNZ
owXVKlJsC17vlzUahClEuK6emoF/K+HzdlSTycJwApWif8QnH/kvMTx+xBiNyRdl8Dj1h2rsAUu/
/HyCLy1YyTIK5OtEYqqLjcbPuJgU8jPTJVSmLCy0z51v6Wtv2RSAkGAyWSgQeZ/gsdICQRoXCdHo
J+AXqcUMUuIUp43TO7w6AofXAuoL60uk5D0vW/SCPAERvOlrZ7P92MD5PZUDNsunWJDrD/X6NbLS
iFmlHupXDA+B9gMMA4+JOsIeKNmPT79zs00TfWZAGcyUuZMb/2QgQRry3XUK5j26i6QDXTgkXfFT
ik0Xay/VzHV3eedQz0ACti760MPlhqZuAhGDpr361dWkeHYC29uMDjGAGb32d7ID6Um46iQQxeFc
V2hNKtlwNjdFoRZnOVwd28UQU+Yt8PysobBs/eP8p4VYzCKEx0uLcVqjN/5DzYsiQohXq6oZ2EUv
fjyt3lp8YEscAUpIDa5x14GqZ5zmjQ0YonfC5bcd/geekgeq+2QJGOlgsWst/vyCY8JvofjQ8+Bx
Hp5GO2vIUg8WrfkTQTjSEM6eFjfLSu1ibQVCDZtxUjqhUTkGe1Yg41YDC4u1F6GvvOBiYTs0BIge
A4RtoO/qv+uTMpkdf0PKTC3Z6rwCNth/MbJY17MdFwylPFssMLezXSPdv81/Tf9CS7ZXceacLtJz
i2Q5eU1xwJqzQ7UqtCzNEtdL93+Trl830QWIJI9xMpJJ6GA9tlK0wNH13mv4ecQRjmKR5ooAUCAK
qRM52TRgIQZDUcL3o62NdJ6kT/DsqiT9Fk1DtkmQ8q+FjIK2GKTKRPkm+Ch79WgIRz3gdwEeGrcE
HsDaDVO+BMh50LdcrpK2b6oe+c4Uqc37RUadznXIx0xdSV4i5mEOuxbywejPvrW3iSEzPpyGN2JQ
9vxRJEyN1dbLE/o9jYqAtynTosFZH7TiMI/1bBHkB+qL2bk//vwQJUw2Ur06U5GgwJQO0d/sciYF
pm+193XohzcldSLSJnvlui+Ps+D0OFwKZnf+YC1+AIMO39yHU4EfCE+KPxL6L1x/46QoNWV3kWy2
u9PzMdj/CBmCYBrktMmdrRwyejWjsGRquRBawO2Qhir5vVakyqdUGwzgGLu1IgVwIGQ/N6K9LVby
n3fVxsZpdYb5XCyPACKqivM1ucUaO710nUIbr7DjoqzBeZbB2VlA/Se7HbsIRRiD4jyYLoK+kNyv
/VWRjO6S49H523aTOp+SNPOqYx2VtjQARinCPd8NkVSYY4km5rqy9fgnDZr4KXJ0T5TUoEF8RVGv
HbY5CSf6wCVe/n+te9zLI9c/zy0aYHwYEWWn8V0BUPkjUg2N8gwLuCZGespwMNU39C4EeKmBT+yb
ZaIEZFQJHowdaM6Aknc/pd/KnXm0383lHQPzCl0v/1sFDSIkvG7MjlrFoGK2Rka/KaSZcY2+Mhrz
llgKJSTLy+F4tlmpv1DZv10JdnOpEBc2XF4P0VWfajI3oWq2OesGBvHMojK1ULqdwXjg/gWh9sEg
BYgoIKzWq4qNnrtMf4Nxc/zXD20e6JymIYbDsJxuKGQYqNEMnU+p3CEM5M3lsQWrCZilzrf20nil
qi7X/PVCDsSE32z1suXF/cL1EMtvkyEiXvksaxt5Lp3iIinX6eArXw4SPY+tiCknP7ZmQ631uJy2
ycbuqu7su7DjjfKuWOgH6UR1UV/UARzDbeIYxYjtLtQ/CPYyWUTeuRN/bsPwIQZqWVR7y/NGar11
VcoAntFSjkjC0GuZk9N9QEJr8tzs704iVC5IenmezeeVwsJDB8hZ0dSlqtqzDq1Dp7Pk/tMIhzev
PM1eLNvzr9sG7Cbaz6OIDx3DgrMVm/DjMi4X5OOBK/CvaRh50XHpxylDzpavxu0zmSlGKkyB1YO+
7f67sDcpnZhX35q/4gGh7Hjqjs3LVToezFbnPIr/GQUQVWLu0JtJtOIQPxagDo2zH3pw8dkH5ZR4
tilLaoukDQzYVs0YV4jdSy44lpQG76gwLfy22ND6/pAKXwQ99ijH7Oj4exy9W516LYmdWo5ha4O8
61fBkloHeShHsEy52vYto3A0U8eojDtOdj1Onw02VtWbe2SClcr71HnEeu+7RBz7TAsMZgoTCo3G
2oaJVGmUItXEgGMWJuP8+TCYS9N+zm/u4F/1bCp+llSn7HJjVTcXbhPKSLBdRzRmgItH71qCPkjh
lGxTY5OEQ1+37UdIAPebNd6jsFyoCDxKYbQ7eQTL2koMTO/+3aVAU7CBI6U/Shj5AyAc1c45TJA6
owG08h7eHUTVrkxzATb3PRLn593PBqVz2CWU+C3mSK9uyKNnn2IBK1P8TVM82YM0aBoVoVAbnxzl
cqGw879YbC4e27AVy1jXKp0KvYk79ADWXXDhQVhYSEP8yvSZXkpdTp22fdQo9GrbWIxdJut4t6Ry
EpAFUOi6xslILligC5SdBDlzh/1nwmP+0+xza9xA6+AKetRyxtP0ziXYI3yP32ojNS6OG+z6Hp3q
NUbvXD24FM44pahuTafKRtOGYOADMoKwb48aMcrNPHgD+vg7xCt5+Ich07E+Pbf2xnW9JArpgCY7
VnPxENQbX/KDVpaI7PLWTJkqwOeCOB1EiduVBXD/0T+Qw3T43SzxImaEnHIeNwW46oPQ4id+WNUI
wR9NnjrlXpGzAbJNeV55vpahcQ2ygrViS7fr8nF9rJxqii6kYbt7gyKnerEIpAE68s5k7KU4A4Ms
JUMLWh7MmbU71iGLpeO9rKQ69UKl3k72OkNfVbIfpbyCieL/evV7buABhqH+vVc0hsWJELn6o8yf
K/8+zZYcC/VfKe09tfMIDdFScy3Xog5j7+j9AwEmLv6bRm/AYKRvQsoEUH3xRUfQG5jfmAF5s1Cu
j74GxL5Xo6k6pl3GIWUkxR0L7+vXk00PE7BE+/TvF+To/cTcBAMisIOj1DEfgCkAC0T0tlvszecH
9FldwK45EEWxHpB98g4l/vT+wqS0EhRAAfNQm5rmLG16AKP8ewWic1RSCS9YE15VyZv7ikqI+7ll
1cNHil6qn/0anAQQgkZEBc3yvzkf2P152RTMpmcykTD+kFRGtlOQiORFA/CP3/e4lhT1YnQ0ryWw
l70cr/uCNUsT5DOBaPVLXECXqkNEwDz7xWWnBYIcW7AUZlOBuieiMi5GNrympYCE9FV6EgIYfWZW
KPzY+6/LhPrTTkXYXmGnYaUP37iSbTJPfIMzGiYWt/hOCxRsECFHj9OMM1S+63ekdIAMxaC+i0RW
so/r6yfrxknBQo5LEX2NRt6BnSAJD/pqmUD0kb7R41Xvodx8nz5OlgMqhH98WDILwiMwM3nV7X9p
MebymVOFE/DHD0ty2UOaPp5w3D1XJBJpg7Po5H1YBYC9JmXeuWNjYDRlbWa0wf07U70af/Ire4PW
ZttLlzEXhKMoQVMae7+rgTSINpAGlEn0SruTdH3MRNwBdz9ZunGf8MWkmFJwzDbQ1x3ww277nztp
3qpsVLJXDEc3EtITFgJc07yAq1dHy7/in3vkG7hU+RtGZwtRnQ9UCL3CT+aFVp94vnCuA0bmIKDN
B+JRtgH8vBzLB8O3JFW/kjS5/z9IwXAZQlGvKBAymxaf3CMsZcG+7t0G8kA0Pc3xvy3Be8u3ykKR
MqJSA7gupIL4lyvuBuV1CaFBpC2oadrdEaBVqitGeAxnBNKsTTmBE/K7x4olH87AOVMvygORSgaM
irIqWHbLWGGMkB8LFFs0FdtxkKZHf40BG6tPJtZ7nmz34IlTSdMLdIcThtVyA8RkZ5sKpPRYwWhi
otHWMzazlGr3ITHxK8XJd3Kpjnk+xkvNjUfGMPr8TE7ugqX6D9zK7A0+vmqjeVr0RU79icMqqk3m
aUZCfk+4G8tZAylrk8ZE+41iFfEoGP4iCb9ZaI9vYulH+gSN0QYE2fDxUxhDW8cevL7FuQHU4k5N
5cttFRnZbqggvVsLwkqcW2uSZoO9NBjAOUBJU260MoGN/AyfHpSISCPr14aKuryW0cpjXyx/JiYA
ZuN0ZOxtP98NBPRdvRW6jduGJIPDME7gX/g9BEbve9PsJyOCqNb1KwwVtNHBIjPW7E+T1maZD8Km
Ek2vEQj2wNvwwswOwJaNYItovnyBzNzxVi7lHfmARLbV9o1Y5trmkPEfTe0RNtsPiX5lZRfdSyD8
+/AJBLllIq9Tc5Va1OT+9oizaDzCcPbyR8yhcO06/mIF+03NkXZo4wBSkzrOuwrKVraeF8u7/rr/
EEvx1lVxfQQ4p0i7Q3PUjRmdrT9LNIgJ98H39eEDf1/6xkaWIblewWJhSslR3RQaEfEtCneKX5tg
8IhBEtEPQfjZSl8xhiYAcSCBquYWkhrL0lgI6rOX0+UznZm9A4i9lCZCVQlWjlDsk2ok25b5hSZW
bziXNoluSXa3Uvc9e70z6gkExVb9ohsVGv/w4Ln95KPgfsnbHni8+kXQy5LFFJe6pwvozMZH/4Sz
Gr3b5vQ3DgnxlpDVJKo6be0WdeovQnRByinaNx9k64Y5l6aQX4OrX7pJ2Hlj92idlc7lbvha8Q1t
n4S6HJu/esh2upZhaeowHaorx0S8Z82mGfuX8zllqrTufozGbZ7ZkUNc/PfFx8pjzY0Rt030p69V
xPKJ3HOrIuXowffHOXlYTzfup/CwAIee7h3Y95s78n+tkdNVdMU3d+0GVaEM24bOEbRo6VJ/VsbX
12DEot/i+B6CBIc3eogJThvtfatUB1R0yDm9rnO55ziIZyzKaZxNX205PfrqSfr83ScPxoV6hBhK
hesv2CWR11Kr4+kFCYtI1bPuQf591FbrLakNTO2STUTVKoFCRUzAhhWeoeLEPNkQYx6fDqQVyeg9
Qcoq1pI0u/PLqlglqMwyZlHyxwn5WDejU1SVQ2GUqnE4L0x6ANyDOmoiaSLnD8JKNeoP+BxIe0GR
VkuxhBjQ/6EhXrOBfeABF4Mq53P4Lv0XUUTzc8oinljInha60ZAR/u9rDcZcH3DWIRBK9SwVdr45
EvZzp21eUA+ktFhFlRH9YkRmh/JgwF7nvSMTu1SXdfMSk00wkohzbxAh6kZwTT7hq3W521Jggww5
i5pI/HWOwr78iQTZ0yHMXliBFN39mVWr4ng+zxUmBjFzKSv5Bepxj/nbALzWuvUNMby3qQGpCfBy
qZOWVXLUpk6YcqNF9DXdh4tZykmFBXBb1nb5GBBXmhg5MwRHcoVGItBcbPRMqYv2KMYGCKUhyaUx
Uzx5+ONQ3HF51sQbmj2X6CeUJCA2BGYkd2AJRxGnKZULYpHGo3ZqA8A2mhBzfJWoaa+mnvetK8R0
5saTbjuciB+wscLwRZEiJOAk/Gyyh0aqGwug+SY16c+EZMaBCW+u7bfH50JZ9IcgU3lBF5vC1K56
AIOupRY1c3TfUhpyjR2PQlhS3F9gkts1jrILAMt9xZ+ioEosqogGWevRw8wzbvxKzfEfhGcjUlCf
g9hT6sXtxVAAvJ7c5Hz4SakyC4JT6VtGF90Mv1ocjX/hrsUUrMUdljCE5J8+KRsNJj3eLyHnHz05
n8pbobbllz47BWbtO0QC3KWV51fqSBei8gLaUt5F5F4NKcP5GO+csRNDcILmB/dzCE3o032vjDJz
iQHdoU2gQpeVEBy4rZigeJ8l3ovRDomXiDthOfWT7oaMksgcc9khpzcSi+zyfC2/TUpPLOB+iVoz
fxpwZs3CY2ZLLajdP39ZKSyrlreEeuMB2AcE4MnwTvnICxFULtjLD+ROyipu9X5nKacWavfNF7Vg
NCIJyZnQPtKO+gkjARGiaMVhemBiufl0WtY8/5BheA/aTtlJhi5jIXZPNPfKJk4zraVh2E8hDZzJ
AphoorK6UUrgcoOi27+eEG9RSR0uBFaN/VNJzWzeajuX1MVg1Phyj9UphM21aA2QaKXPm1V8NBbJ
YYiiIG4cYCrbGd1DHTpbumvGSDQF8c44qQsb2NJWWtqeKzhkI1+zqbCP2U16c4vjIc8nfqRjsazo
j5C/2VlLTH3+Dg5tXT82kV4Ldb1riOQxTeW83Y8ps+vSiaEO0tFwE53CSKxsyt0OdKlo69X8jne4
2t7vVJvbSUPoSojCeN34H+W0R/9lgv57qGMyVIqwvOGjLFmPOEsNmK+JIQ0RJ/CBELElB81io1q4
3f9q7AYnI5T+xCSh+ISQM4rq1g2gP/3iAxsQvyLHo2LSXtDA7rKysa69soQYM99yMI6WSI8rE49D
4gzmmmCnvwMSuon8vw8gEsttw6J3k/wRQ3X2oYkusiLjCob2an4JuUGWho91XwnlIJB2kCI08ZHC
nQMp9FL0r/kE8g/egi27JFyNcnhFbTcJBuh/0X8W0u3sNRGN12AsuAbDP/brDLcdNCFBSqy5hIS9
/wGNM73I7C0uZ2IKQqp6dkaslToWFvr3S/Xu/uz1cka3dlVLnijjh1r2pcGoUxiW/F3nfAp+X3fq
uJGbhq4IqAFr1+Ra3NKDFsYFqFcP0vmZ0XmwOXKKECJG9qcfcAaEBQkeNWFniA76UDpSj43QOpjF
Fz/5gJRoxzj/D8sw378q78vdUCBRGkmmNvL6/5Dr7m6A7ZMrf7SWjapIZ0gQZgIIiyt8mISnrq9o
bPfHzUs6MEwmX6NSjpq5DrhEK26RoJGSIXaeIqDvw1gYuoUxtx30xQ6RLy4lUZAdRp/+Nh0yyQoe
Mmf+FYLZfAMDCwYbAlskMYeEkR2hu3RX1D2kaF6I6c5NsIb62h7oNquhSi0dAUMQWJlzDbYlRAXj
XE9PNOe0MKo5iM5tDlSzgsqcPWnk2/3jmAerL2Z/Y2efDd5FYxxA0sxulQzN+DeBuhiLL8Pr6yXU
8oswJhjVEC9bOxihUT9n6r5EdAkP2XaeDJnGH3qS2diBnE1OAPvYD0OSsr7rdjsUROPbhPaRBqjb
tmvIAKoVtbWbc6f6E+DWu2jfsnkifyUsuzIFnVQo1522n7ro8OZ4nxdfukVziKXtGc7sakozLmnf
bQV8rqmrhVeG7dbEngwWGwFDqZxbvJ7Qxjlb44udGrc1AZoiSth6iWm4rWsza1s6EJMBxDztQIAS
77gUaQcw6GRqfDUAHoQJ8IDV1dN2qOrDzdOk6yEJjX+I9shm5hRRXXbPCW+D1gBVCdA37R4aR8ac
os11BbHlS1tLiza7A2lqqJuY2bj4m3Sch1PpPbBAFcT91+zWyImOc/8GWxJqhyHuXxFcijJvgHn8
EWRj12ZvEwmO5nRDk4EMsPio1xt1npb/yUoNlro3bAXBj7JnsV+M1/QcCXg3kv3lJlZlDQT/yJS4
n3FCJSbezGyV9PctrkEbhoqOCwiltrAoXGml3x1pRl5jxNFhC1PL9AmEg5eZATNxlgLEQYlK6bNz
JxXGEnY3H0Z4qXb2GvuOQ6aklwBb7A6NOgMI6qda8TFsbkgEN9OEPvnRiejU7tnMJ2HElsOkxNnv
bsSG5dmZOXnCoLQMwidNnk39aSXuWQNuhYbvpv+4EsrHACg8d2iI65do0eymLa8DuOLK1HSmfQOL
s49WiROSEPrjnJtaSf7/JTFI7qMZoBg7uvOavZr7+cok0w6KDqFM1PqOUjB2WoZpc/2GCFElYIQK
PvAxQE4gqphRb77rO1iu8Nk43HMvGnB8GysmWFeyvc/BviIXZvxvWfwqkUH9QjRN9hTLnGPWSIw2
IQOYjvjAnQXSAfPaoPorVkKphHPhKgPUCUCmy9Yh4FCJ9/qIn9YQKBWM0CIU070wRc/fDjSVlhaB
IN/Oau1rgiV4tnnugDyHXCioRbxsls/nt9bADMXIV7F79bTq33KZiLJi2JVmZhpJewuqfQ7q7QcF
4EsGppI8IldLEY8NeSk4B6861/PGC4oMlIiJrCTLl7fAEqWMKtaY20T0OFji5KvUJdtQVBjYfmIE
xyWvn31sE7a06TAnJu+23Yv6lg0FfvBUSm6+QM3VoFXm/nAg/1Db2NfSTVU8hIU8WCloHPvfm3QX
GRHpaiVijNhgifC9w+X8aHZVJAawJseVXr3RKUkgdn3DgBPQfdeVk0IqAjfPYanvyl40xwtK5gPP
hTqV1my3Qt3v86yx7ekQjxknKapVoaFN1kI7W4MWTJtpX9/shsmdMoxXExIUaN2h1aQywT7K6oYL
7NtVMGKx1jWnG7mQA8JD/e6NWqExx1M2Qwa5giuiOS4kRZnQ34CCc1Kj17kMkgEBO4M0UKXLpl/L
I5yE6dNwB1qKfCg45dQIvfpf3J0bwLbNMyo2L11Q/cd7y7eV5fsjTOHL4hXy2qBXweAT3znMbxha
6enONG0yaGXFII0bdC9X2hL9WYJ69f+S/rxp/m1i56MSu2qV5sHW7avDrCwye4gHLQKqhFLExxvi
GjFkUpADFW7NmUuYDCJvCyg4X8yFWz4J8JL2A7NoZV6VCay7B/KyBr1dul3bNgouBqold6AIejhw
EBoagU2N+WZsnHQwBgIdWI1xnWRncpZbWXg9K0eWgT8V8HIZdVVDJhehZqkNkdVbRk3NRh+Of21S
vCc5IbO5gIeYZhx2j/rtD3gJXA2+zAg3wnloivhgFybwLKZBGwuT1VicEgZ5cc5rx4NaLbRKU73a
PE264RnCE3xtApkxHxb/8nuNjrld1n9QQhAOvL2joir1Ezkbb680Fz6BLS/YtELcvMnrWC+ZFty6
6sR6/GkmuLyXrgXJ1yhpzcpcNtHHNxy3rtfrnDoW24CFRj4sEmTzRytOpDup922iCMJt1Ds/kyZe
8qtEaGlsGflNrBvoERhLJm1PmZHkm+ETClhgTyO4DD7eGC8O6jY8tb0IEfyrKiayq/cbg7RrwxDt
zx1uu9XyNzkqPyDMwuejJxsdPSGdtZaB1DF4QTaDdb5Rq+J7vUgsWINn8z70qCspnhGUK2N9sIUY
tZlcGzInZ7FanjCIvnolvnQTh3sNeAPBKUHBqEo9VDrK+msVzEXT3EoybqysDze9chAo1SUZwhXP
tcFs+vfH09MwgDJ/xXHfnuPTQ8DNO91Yh2RytHBmKnqw/u4ezWIx8s1UM+MBP7IXBOWBmwzeF0xN
FhyKxjsACOhrptg2qfY0ZyTrJxYCO04iqIxcNIzPVC+tkrlA5FZQtHrMxzDI98nZ5k4TLkjIZ72E
7NZ8YkDE0mwRIeCQnEm1lKtT6UvctbegOtmVhuzeGmoKx/JDrE2Pzz9pUmb6XPD0tkTq6XJOBjaB
kwZUxYoC6sN5ISJcIpVsojUBltyxhK/Iezxi7svv5FAl6YaF9F4VCRDi94BD09A2QhUrhivEd9rz
xNnMfcWPB0cA9gPy3tF4HIj+9zrHAe/K4YELnfGo8dW7k4wmoFObo4Fr/6vQimNqwNn9fJbPb7Qp
PpkEsgem67tpH3ZbajMy+AuAjR8tb7VZld/fd17DkLZR8F5XI60W/rMj9poA3g0hpS0bfcHOIEgc
8nRUOBO0TE13BxBqnQhunpx/hACZikek7vlDzctCJb7hl9mXseVwfhUbJ1agBw97QhJrrwuUJAMz
a9zehThoFRPatn9sBxwXEe5Z99uEzg8r8u2TsscHdi8jx2n5dHtT516pmb4qZekLSoXlBR6P60TK
Df+aJPwvd+0IH4qv8SLCT9V8lEkJN6wk7CSqHgJhbEM8k2TsJyOsIVLV5hMV5zECpdA+EY5Jl2KU
KsLMVPV29A2q2fzToFEQmzo0b9vxxzdmomsvvV8Yot0E+zTsQ1UwsUgTzX7u+wUpgEtNC7RO6GSF
I8QcQlT7rvTYWZsC25wtPDaaiNDd0JWKmo+LB7X/kN0T6tvA+wpuZmaYwu47UHjaVir0jmNCLE19
GBioI50++nK7P+HBFExeoWYcM1l9aIzX1Se4H/MtzLhaiCuC9Q3b8JXeQJThZKvEZG0cp8oqWAgG
KqD4eCMJl4yabCchNX3KjEqm7W5cACkSy1cOQbg7royVVhHBYTr08pQTBJRMg7Fm5MXs3IkU3kAK
Y1jR7tzPHsQHiTR5QW3CANBQK3yr7XHtI0ne/4Xw18jBkg1zGpk9SN3WlUyMbLcDO1/jaGZo8eVj
j0a+iC4XLKZUbONGnJQOOOWFbnhTcYQYn0eA0sx5pUkPtRLTjPy7MjEqMTuNrHlGADUr9jImGLvx
zArLqNEN1BG7gRkO5EMkuK9S98NsHjIZ6yPqxaQXnMDgXzlCIEdBfqXYhm9OD+Nj3LAHHW0sXKHw
QRLf+9p/xtdqFXE5xpoqru+x3+Fj9QLHTub1UUomLL3Z3sgcJdB7PZ1JK527pGjaKkZ6hgSnz5+Y
TQO2OlXCJ8X1FTumEhbPPPQVShtueMgfNW61/3xJwYa+K4kU8Yes4B4hmsoix8sOLVQeFhXpdLJM
Cd2ctDENdEtcixDdfuVsUS5D6U+7KJm1FUOZxec40evefs0roZBm45JFB0CkqcATQhUXTT5cRlZF
v0YoTStq0JQMVqLNLjOss1C6fYBpAogVv7x40KUT4lvYxg5+1EzOnJX51IBRsJRwuMTDMkzLPzaj
KfeGVrPFk5eZO45q+bXD3GrbS0fW/M5ZIrXLfm5Ak6rUzR6zUdGcWlF3Tu88THrDHAZtCkwzy++n
l4PbpT25GBjV3x2m5/JG28Khw4Fjy2XjGQn43zs0iwRWWoBz8HVzHn3GvEiC7rGMSl8pFKGh3j5v
YbdMEJVrBt7vLj8Y/+O4Wof5nSXEbwDa3H168hvr55gGYmZ5DF9QEXHQ+pJwRRT3JfhcuqsMc7rv
gHSJKw9dDhGjQ+JU417SPaoIUH1gQ/KqZD8xMnCIxCRgkLWqnjQwBLtNG/3b5YwfZA4mr/3l7+yl
CUgY/JklPJ1vh+Yew7CApGAsBZ9r6Wu2n/L+NWVvoAwefWQXWW7G6doTUHdItpMwq4uCOFBa3UQ3
rDQrqJUMNTPYzgdIcbM40dHUbHL4vK+EAR+E2cJDZEETXexRT4LmP7IiIlGo2Nv00d0A+Mm4/hHI
Eu+O8Z0IXGp0RaaRjzH1FJi+RNQk3DI6uzqWAdTOnlN7m2td7oMOk9SEb92PpX43T+G/MuTFirR4
4Xo9/227bbCr0RBBFYGspsmEza6sN4IifVxn+FmhpYmtW1+KG/SpYW+smF/TOSWu4SBpbgfB7CTH
jCbgxus5zq/FA6gV16oc/mxFZjZcVEROfbo0Ufi6sK9CoM/l3++ajyt4gEYDNND/3n4CyM0wtero
Mth2ny9JBVJpkQxoqkNT8T9h1yPsJImxhqYlv+1zvgbswmQ/fE+5FNuBxGjhoV7XVsrlMjzF+2vC
RaV1AE4smcXiqZxo6/78uwNsyA5Mj0G3nzldM4sPklPizZbD7oC7HLbHVRs9TGTqfZME/B4fp0B3
2D5vxVGcCUF9ui1LBo8l42vmnL+5pECeVWSQahngnlu8EEe0uCjKjHZ34H7p9xjkvPOnabdj7qnq
cuB+jlbit/0gMu9zchris5dm7o3nN/7vIcbLxCGnUtjlHY21xTv3tDTD5DUlQm4cwTuHhC6EE/0f
1mSPDvqitrntYveqk0lvLCXHeTgboIx/g7e2SWATB645ewY4FgVV9pnnVrS9u2iio8/ObzIaa0A8
xPGaNHNPWof7GswAG73Dyf9E30cFuwWa8p3QD6IPJg289GnkqmWRJxaoetzj9SjEPf5THZO612yr
5NhxQ7FCKdZj+fpbFj0LpX/xmeNeZfIQFsVR8CECT+l7LHpWmkk/n57sg7JtqIcjaYqOP00yIJqI
M5PyQGgSqiy4emxSs+vXbz2rNPIQwyqPPzSQyjX/bzqliRLapqLncOUEiNzTpIWC7nEZPC8K+HTQ
76bVsCg1vx1EQ0HaftUa6A/paoyb2klewhhccIe61PVMDu/StUcdUyoxl+3xelHcWe9WtaYR4Xid
TsFOz5TmBdwnF8LXOusbmWa8+ltJjjuVyotCAs9SqZqI1prMIM1vtxECvox8UONPSN1ePHp93Y8I
BbY7mrhE7bj264xYbRg7q14AmSdx5rSzRRHaUkqlxYWAw21QXB62Y63PJqvF9il0OdLBiDKhJuLQ
9cC8e/ICiA7mPfUhLbGR7n5cHEn0xsntkm7dxzDcPHdE2iNrS0Q1JXAZsvLbmbKfprZqwyZnotI7
G6jssmXRrOglpUCDZfEyGfQCHE4+swmDSK6tVdHQ0SP2OCFX/Gv78KdcsHwnuAYppSNxwF5mIh78
hBOr20xVkfAcdvbmoBDOEJiHEbLVsarMCjsHH992lpL2m2D7ZqCGdiotg3jiEAA07SpAtV8Useel
RtO9E6Wm8Ux/sg8aEoynb0c81GdepP4TVlsOvTIj/mjMBNbMpjanynq1GfES/aWY2JzHCQjY6mfy
YMfJSraL0T27kI7eScy+TYCOI9cPhZUc1mZWoLB96KKiGiXrPaNP/mh7AsEaa/+uEVfoGANxbl0s
ctf6A+UlC7BR9vC71RNJwKIBcJO/cFC10WvGmVPgml5NCeOXiaq8gg3oIve5oouarW2ft3BKA7bo
V36C1JAUPO2NBlXUT0Ve/kPRGdF5HD4uaLm8d5b8UEXtfqgLT4w80BiNgGFJEOTLXUIMYxmjKADx
E+viSdBzC2Ih9b7ZP9NyP8bX7fdONuo3+GaRb7tBnfHWuEL3+fJKCu8+oUjfOZlq9jzLo49bvblt
xSTqYODv0cw3enY18ymIdaBW5UI2c9ZKggVsVEh8ese9zEz5xXCTms9x3a/hSxXiw3kfMhtfUPXu
eP9+1C5na04e+F5Rrz+R4Uce71uNOyt+WKmWzfDVn7LGdE3JqNV67F7JyqWwiKGX8EC0gR2Cskef
HHhhoDJJTk1Eyh8Thb/V2mSNmk/3ZbuRyi9xcrLGswumTCe1XMVq5wOtQxO/G9NmV0ad65A+fJZy
3PTUCbMHfmO27tqvsXkGfLw5mhB/WwQtJoYDBSGDwh9kewI5Ty+QciQ9LsET/Ef0B9rCJXJiflsz
n7ZpMeliwM8hSJZzUfnobeS2KNbZ2hEzBNcQOMH9js1KBrvLAs7YYzLTJael9Eb3nJ2rqRO7mhNw
Roc9mtbRI7hotrIUBYlVQ4OrUa9maL4aRwgP7QzFPTrxsl5dDE5ZqVBuSzzwh7JxMprLifd0GxsO
kxHllUoq4WqeQA4R7Rlw2VbFiwWd2g7WOl+vSUurGpdOUoHvU56A6ol/d2SkZkJ6ZZRS85aVgyUq
0sJxbkDfPkjqEPlm4JSZQH+5LnY/9wthvGzPlc/wGHzTlzNDC/Ac1g/je9zzdvF8dM4iAM2oYaQ1
IVD5itVtrssoHwRwQtgXwv58djJz1qEhPNfZw8Km507wqq4ZwV9pHKEOnR/dnk2xJCVt9s4D8B0V
qpDqY1kofMOsi46iAWeWTkPqLogE1A5mRRrwpOcGguQJo3LnO4Q3gXJKZq7G6oAlKt0ywLqJZUbS
lBncIzefNcqiiiz7lYzbJfGwKLCzZnZO8x+PjhEu5dw1AN4RV7APMqf2NDA088CRY2CnfIKRXAoU
iIFlMgpJUC0abinH5J3rV5z46/5zMBWBBy9ZKVyDKjrvPM+whRdFSfhN7r5y0OLQbwwfVnnp2M1+
IR27DfcEvV1qzpEA4SZLMJh653qLDkdfUK4JKbzIzjo+s6JGXppxIpNfbw0P0Qb3bcG7PRBm2Nxi
tf3gfkKdWw74JdhZ5JQTZVQB3wu3jBGRi5V1CPu+J1n5JEVkNI80Pcin5vVKASzK2XfQc9Ybzmp/
aaMKnts05GPmOLUPAPRxWHyvzGS9ah3c5AMhcUjUy2EI+mRUKjOvo7g3RnhBHF7pvGulIdfM0Ick
Is3jnMVnekLY2D4L20rnoj9QpVUITjR+ZbP3JI2SC7wGEr2l8+e6AAvY/fh42DTT0d74VQe/ThTN
3S1itqJD12+lnNO9a1zHMXdTmMBYhiPjzxUnmClLefniYSpgnlrVivfGvcpBkc+OFHKstt4YAWO0
ceV267VgcEcmgSqqZgimxZ4KmrcaxCwVNv8BseriiFBSASzb5fxgJ5podvQ/gKsDZcuvfZ0U5iNW
ajLw/1abXIFG1wmzcyltmxuiGcBMoIX4RWnDl0VXtdm6UGuEvhbt1PZ6RNtul1D9f+pUhIShsQcf
VAWf5S17zWt90vT6/N06Xh3JACs642NzRLw/M+tKXOWYkSdScCqKeBybZlw16zS3/g9JIpYfkzpj
ostC5IxV0r9TxtFWAU8aeaKdeloHhXzyHIdj0jCbcWGQAIQFyxopQPnJM/hMqUxmRMrCggg37zPf
PkVcvL+H70g4X0Jn8w2c5ck9qyfMDvTAt9MSb0RyIiRY2CLch85VWzQ8mx+ttLI1679KORr0fENX
ZwXfTe1zL4M5vsXbEU0s+kswGTQ8Jyj4MKh05HY2vzVnH53FUc/uUK3FlpCSOpGHz6XsECbYCqSe
yigh6mJhTKDPLnw7QJQCUk3O6TcoNjMEszq7m+XIHsHYXCv50ZX4bxw3IRMJnxeVYWcqk1lVHkzC
J7ZPBjmc1CTZ4Fdq+E93ljtrk1puYkHKDxcrYbn2xu03GhGFWMfB/2rqQNYS5Oy/IuLCytZj6xI3
Hl4H+pgmPwC3hr54yrE4pt21HMp5AoUydTh8AvGXs8L9Q63B8kWKeq8RwQQND09r8WPqg0gy60kN
9MH8XUaGITF4Qju8ahWHlQH/VPQitxHOIdhnCdZveN/omeWk6lJJnkNdTVC9S52kxSkaUuSaXDGO
XwuCiuZh9awJ6T+/crz0zg8gKJW6jwX/V2kUK/FHMzS/f8LOIMa2NRwAXNIubLPFarRJsXdaHFMU
wX5iyFrzycUmljZlJa3jaPnMTNMxC4/1WBz1fJvy/lnpY5+ZTTxLdSV6TbQbaWPqK226itgJQ/Rh
QoueIG7jR30YIq/KySKm+jjuR/wjYs8ZOp4j3GD01SPV8PjVxvo9exxG9fIxdVD86tIkELjELoak
9CWXmVPTNyiA41Z9mqXNovYiYO+QrtNl+1vEyNe2C0m9+8eLXYs5QdS1Jgv8XtL9GTnbzNSa3NJf
v9mOvbo5akF81vTqNUHNeUnrDcdpGdPkstLNM75KnfYqDAThrF02qZvqAC7s0U9oF13rIhbP03zu
kboySGgT7C8Uz2p/+lTAnm91WgJqUPZj1PFtnhk6r2lUOb5YPv+RirkYmqfUJX5eo3nEKsA4jDw8
o0tgfERDBk4yLJfkKSXWQ+gztNV8yVFyE0dcGsYNqSUnB/0jRTBl+dXqNUpQlzy1MdNwo2gNXBLC
PEk8mcLIf3W8qJpBhUVFV5XtmoAwfEVP9wG6M7w82rrD7srcxxCs1U19X/GJrt2SzDYXRE3a5RVF
Jz/JmZn4A1AniyTj0kNNineyYL/ymZuT5Knr1XQXwpwAjHYyViIZVjCVTS6enPUmoGTtNZjPaaPs
gRl5klT1ViN4tu+T3nZ1g5Ro84jDT12G/8KWjWmnRBGN7y/i7m3K9fyiQXRbwfqcgsq1dXGlGEMg
s39EJIAQ44H1hS5z6Dv6MkeE7Y7vfvd0WXi3R2x79cD/EWe7f2LCCM1szngDcVsh4I/mFs9BPnHM
OyoIy6WHqC0s6TTxVU8YS1Um0amjRpnf4z0L1/Zv8ndKK35WtK1ExZCeLcC8PFI7o02WCwQ4/74Y
6KoouUMxarzP+wqb80pY+vk5Ft39QVhML69zdoWa1tPuM9nyB8BJAGnOmMsNPNUZ+EJfdP4cDKq/
Lg632yyoHFKLefjMILpkolwG0yowuuBUq5PKs+FJZWuJAkacdWFLPHzwvnK6FWKf1YgWLslJXZXt
qyGATdQYFYD7ZcPqYXSVWL/ovI782LU7Y3YLlr8D4XdCWB+ftZw2/4Se1Rjq74ZKFogawzSE7A9s
R6LrTnWdiRmN9fxzWda25ieUSbWaZnXkHBFpx0WrO07N1bYkO7fwBvEpn2psiDOcZiZvpvdzPBii
ofz/kJqNUu3nlCzPNkD/4wqBTujruokbTUJ68BmMVfJ5e6+Yw26BR0YXn0SYjSuZQkDhy65AbLRb
NqASIR9o5/cpzOKu/G3T7FRXgG6YFwrDTIQVqLgmvnq44L2hQ/uM0vrUAx/eiX9z2RKUxiEhYu4E
ip0Q5aa7oCS4CFrTI46n1R72iyBLJg6mERRi0V1826lqF0skoAGEPYC7CP4dIjILWPajFhyiBteh
v8Chh06sFcpjm4ZGY+fVVEhacU50bgw6/6fhPbXflBU3wnI/K2dWpaGkbIim9d6F5hop9FV8Yyx3
ZJvdG4ekp/9ydnXYTtWM7MVo9gqGnjQ97rqGkR9hhX17jkAqC2gN5mXL2MxcYIzN88cbnhd0jErw
2uQJi+xu5Smfh1bT2mcCTI2twTC/nrxXnpdqN3IwZHvKar3DOqeFao08gF5vqlecg7ocfyUFwMB/
KlKMKzPkYqiWycrlelBvBub0R5J+bq5Hw6kALfHi0SFs+S1t38+DZQED7NmUlambN+0XGrI90cnd
j2+3yj/NgEmLcvYmw43Yk1HAwr/iH4fowgJvKQbpdYoItdN44wmgP3CRX2ZWWHAGteVDid47rO7V
wiRR1Ho2dUTNwSl8dNofLTtGPGfgiHx44VHyIGnfHDz1kvMDeQuuzbwXXiiTtI/LAprGMUAlzZQO
h+cyF6u2kTC0xv7HeUheayoVXRBp3xhiCcolWXmQuQdiLbrDzhMLBQwLS2RJqGut8wPZXRUQtb/Z
4czxBoDxtbQB6zCiB8YpvTQVDGfBDLVZKt6gG//joynAh0vbBXiN9NIFYqLpZPDBeZWRn69mu72O
Ac13KKMaLF2Dl9Xf53QZtkpc0WC+c8/QoazHgQhUQg3s8OKnJRGJOp4bh3TNlSGeumdteVKSUTXI
S7zzrB/P+gz9xR2YWzoUPM7/L0vPpJVeki6VzL2rMAQR1LxGtYlAGUj+DgqcRPwRwU9EGbmSUobD
Ui77xjCZ0yiI3wraQjzbQV9Cfcopkli85HenDIwQtYFs23nZOd5VyiAhCfTo4MNw8VlLFElQ7TbG
iDcDfj5yZ/yvW/iM/taoa8P1f+jfg1fvuxmII5hQ/xZQiaSLA9OF2OEoMgMIV0paCOZlKyyA6NFh
2wfXeEAaRKsy64IYxS6m9FN2vtoiryRurpUuz1xHr8vIlsDe277XcDTw2qqlEfBVvyyQPg0/uu8p
9ArKmeTrVx6y3ZpBM23wP1S/zOLmFd/pUl9rM39gT95RE4cLHw4oOH10iZkUWpVBgnlHq9qsJ6QE
8xrEjfGu7LMVQaqZk96f4KhQrP2H75os4hTztCYaP9sfaAoUKvtWK+rO8vrCxeZpKtSV9SelHwGo
pWObTYe6fMOsqQrS03DDInklDDeLPwG2zApCGOeK6PEOIx4ogHJMnWDHS1MS2sMYDED//VoOeNFY
0G1/WG1/MEL34KGsXY07B9UFH6cDq9bOz8O7pTVMkTl86XowikBUW4gaw2WM6ft6EIbG4ocjpmeW
5euJCypexeFo5uPj+8ZI+78A7NyLKba67askAnlKPKkOdnat4iSNKf3QNY2Lp/bGZSRPJxTTyLdA
JULtwKgiJqusuT6GWLycdX5iB9ol64vdKmcYAkTZWzDwhU4Q7xsHLlfNClshgMi/SeVfcoyhdMkv
tl7Tt6aYPRtpayvc58fmj9+T9pBBcE1InqnjcnieBeiekFBtxV5wZ8h2IGYson2k+C9ykcE5aCKt
Qch2/QnQMOmak3rAyUPDSABDQXLXT+s9CeHYMdH9yQOqisW/D+/85f+p9Nd51hAqZlBBQQLJedN8
hO56YRPJgd8oTd9kg8PXCe3yskPQgiJgirS3RmUhaWCss9DmWRRYZDE5/4LfwNGzwDHwUwUDhZaj
o9yEIKoTRrk7h34O9MhkmTYaWq+mcQSwC+sM7ofstazIaWglRqPQTY/691bxhzYa6nGCPAYr7ec0
gSUPJvtx9uJmdNQbWT5qrKfsfC2QgF3ZETPs3QwIjqeZxovooOj/itGwNgU0vOhQ+gQSSzkMSurD
NdjyaLCfdlTEzjoM5IXCQqNN92K8QzXAZ+7AStlrg1bqshXYgiAR3q8igWuJbYto/X5Yogm06oLN
W6m666l7LtPXywlAI7Fplcuwqn+A3ogwRSa1iy9Yye89wtsb5UWtjf+D8HTSAEJRb9EIkhz6wd2h
dDrpQhRLBtIry7QdmdqZjd0spqXBHgMRoTlgcK2CzEuKAbaGCe4Um9seFkrXmfY/NFX+sicQqqIS
ftRPTQsGO2xzljXGJWeM9OpBPjLRyHVWZcwiN3NMd6uJp67SuBec5MGUH7p/YAML7Ld0FCspNMYb
+F+3kUmFhdYEHHrXu8c5XPrGzvksgSJFZmPEDhXBBHqT/nuwqtN7p1SHyZ79z96fv7M2Wx44NlGS
AeMLSGhiwNjCM7ZwN5vN0ZB0g27vfZSYBExaBu4wdx26wnwCclLIrpZ5eEqGC66BVeFwy2Mt7ZA8
hIx+WB5IVXs1TNKpBId3JoRIV1lhMzn/WKG0pFqOI2azSPNgbDcMM1y+7RhC+yodq4+jiXNja/Em
D71/6eVYJHRHSrE0SjrXAZRBm0lecqJWp3DnGzGUWmCodefOs/B1pojmgbpsl8W5gBCPKRCLvuos
fCkA/HUaSsKuwFY617m2Mg2slIS5z0MdlnyRBEw9FYIfy89/K+IEH79qJqiW+r4nl7FI8KfJ9eqj
enuQfUrnqwKs2A2ZB84Kw+PYexYCC3DLsRN4GCh2J3kzrpSPSnWJNPqzCAuZgdnH1jrQsutvLtQI
ZsZ5195cDcfqEuZGFfBM61un/K1lRGS34g4d/FKk2kgXt0g0F+QppxFJd1XabnypQRlYLC/yHyxI
bEILglGd0CohHcHmLzYdEiRPdF5jAXAxvJN3+tdBJni5wAaY5T30l1I51cPBKpslaGAwtodRuq+1
FGigDF97E3iDUX9cTpuYiGjQPEqI3Q3RAF3I2gNskTpdo8s6iVD2tk0szzg1YT4wXJv+Bl6rHFX8
3G6m46g5ZTZMWs2mCglvCvNYm3z+JwFOuruJsS4QjCZhmBu0Xl7XI9HgS1cBTb+97oyeF6Nkh+P9
MpCiXxNSTIs+0LR/rlhr3gqR3YR58jYL0FVJNsMYtWgZty2Idc3ucxgnbUk9ZmOfGnW7POoXmu6c
lIDn6bq+TV0fJMyLbi58HjOlSSyyonoGaltF/vZx/qkxbunFAT1uwZN2SacJb7uKIMiXPKE9fz0t
zvFniHOSdJpJaNs2/Xm1q+k7BjDefKJdNH+HFOxWMG9n74u2vcolY/122xi5ZvMBUVCT1BKMnrK4
obAu0dBRHEWFSTC4Azp46N9irZWdmZc6MHEKP8lFPV8XlV14Rew2TfxIcKnISjblErq/F60ylG+w
Jvs7J5IAkTY7havJiRVYavCK6QfSkwzK13aaD2S9iJ7dLARUG5iMi7bgQBqZokpGK06ja+4PwxHz
lJ/dg8R0hPPHUExOeNu6y0KQqJFf6t09odzrN8zTnJW/o827ZrT1FCAQZtdyALZ7kSWXsj8QmLaE
W9YVEtve0mjJlyyjr09hFzWFcnHwiGMLCGcRiyrVHBV0lqwmAc0JBK0pkoLVR6+Uw5wovMRO/VY1
YsGDvtiHPFq6uiDEthe2P+zBnpvPMIA81DJeADLWGKBhDRU773k5vprG3Fx7uCJItuxYz12GC++e
wEojXMfzQxOdqAhy9hddXfmnOHfBj0I6eI441mYosU6jjmGP65aozfEUAXwS/mkF1hBMtr7ClwcN
axiYeFSxA5Ewnyklg3XKnwc2tp3Z31wo/KqPlJrd7JlbnBCU89mwD8i4sfcwFYgT+WRyKjQ7N26R
/Ju0u2t+E1GGKHHmH7YcO2axR+nIlTKCCgZQ46PvQRu1FKoRjjXAz6T3tRK8lQN4OlYnFfOOMMjc
thWEJTNEToOBS5nbVTiimZVG4Cpf3eQPd9LB6ZZFxCxZ+ii7f9hV+W1gN5FrTpwiYU0o9hmizZB3
Zv6+K3+a2tnop8op0F9XFtjXPabFCbkyRvThK2el56O1d1fqI1/end+s+PvMkFYSNIOTGea3gL2Y
c2AjUKx2W4x7Strg7v9PBxf6MOYMCk7zR8EUke7NeH61NczR2n2m2dHeEwhps1O3QoBbNxMBvP70
pNR6yoiQFs9usI2qjiIWupJEDkYSjROXJ4pzXL63XBaYhqYJgd9DO1AxRxykO11XyNHHQYTS5BV7
/fgnwUj0p05JPBnQQVaOwE0F4J8w51eQDcEDo5IHZ6q0pm++4jplMNduWpOqaMQqb6kOPz3MU0qf
WpdTzgakC1VhPsglWP/7QTOw93rRBdPL9hO8KCcw9b/z/XW3YC6riTs+qRHMVXJ5UcHqcsLscgf/
brTlc2P/DzcUDkfM4oZLczicYcsxDCEyJLFWL7DAR8EyHfWsyF4GykWlYLUfLkMxTsYXxnlnQQvh
6HGckVPQpCpq7cfz7iuRgq7eJuSejRw6/Fr4Am96lHroDBWshAEp0QPaaUDieSKyfZv7jkkaG/Ju
4WqrHWnYNdxqh1fCePHoTg6lSGBGQVDRCBbIo1+FNm4H6WqmX1ZheTp7sGR7BZoJnBEYwBQTrC3t
23ngXs+a/GTSzktN6JlCbSv1MCvetY0CINQnC2VNyVnYNHNnWSdz8LQvRzmY0bHsqG9+u+uhatOl
9b5FsNMWzM8ikrNLirHh/gtrEEzT06DenHOXiNRHSD/NRSrU7kKuhHmlabjiaI8Zfl2pUw5/5PXJ
SQTIIYNrLW1eMhy291plSkbkYpWRQbysUHbZW9GgOCC8e2oAR78PbPYgAC0YIxNGgEzD14df2UBW
7t6RXvacJBQv1B9MTs0F0aN/MST9j/I4MzXBDWHeWfuOZpFAqBi6CCfHjvRB/V7w4ryWdxmUNCpH
URdhhxredIbCsmshxifAHcd90yjciXdypfw6f2PnKj/jPK5XDa457DvO+UB3uk5ZGQPu14w6n+cC
NDJT9o0y1O0tcY21Wtgkhur6Tjp9cTrZzdMwa7V+/xQxrf5Fwz0GeWvhQ6IYe2POlliu5pi3Ckyb
5B/qCNXfe0NIz4DXFhSX6sZHdDc0qcm3Cdugw7IjXZUsItaU5Cv7siAudR4HsJ2eAZVf/3FCrWE8
EnQnkwSSSgClL6YUhWAc4AJ+tBckb2PH3FowC7zAX50Cokn9TVwRM751KvY9uV5j/0Fv2KPZpCjj
8IZJux4AfGZVrh+BDz/VQmV2uhK4AM894q1fXGFGYDk1X3V8UFGKtxNiNyXm6+sEiGPzXFC9NBga
PXpySM4OPF3TOmtNp0pZl1TqknmeXNdnQujuZSJ3tcNr7Y/gG5VUnwtRk5f1yfHvmNB7bGKkOiRi
Xij4VsFAnxX0Y4He+M7kf4v8gS+pYGozjvcQcqaguBWZBkJ7SefBdG5dj0soM+6ueOWyl5CnSDXF
csbmWgyjgToselbfMDqKI5By68m4ohl0CwIEwl6Jh0DJLcbOzK2sq7aDsNdhVPhTJ6QD2N/qjI6h
daZ6CHieC7Z7w0ctPO1Xd+P7xKeI5atw4tFmD6w2Kex4rRe4jWNtA+0t1f4kV2UuEdAVp7hPMiTx
30SrmUgSMnOp8JAtL9sDi3ANDzLTDVyBZvF7sInn4XmErSmLMfkNoYVrfMnDygtIDrkm837uiDvd
69RoPHHyvUE3dKBeIBRmiO3kwfkycWwHsOy9yfe4kLkiO/CnhZfeM1nHXAFT5t3NciFG1nH4TP0b
rSuMTDSnA8+6BFTTNk8vs+ROvQCYq2ivKYEoPB2ncRrmdSfGlY4y4Z3uWns35CjD1IqIEN5CXgcw
PGi8xXnuyXr1NqGyPzOT+R7B2APWYDwMGb6mTUm93Wt1z48DqPpPm5ri7n8sP1gAwgH3Xbptc//x
/cAuEH8LTjxGGYJZYVCFZtXcF+9XV/HbzX94J20DDl6tai7rkdK7Sd13eKobpvmO754pJ3crpn0l
seCj7OV13VeCP0QIRo0ovLnaTYNumuxtPgE6dDzmekSSLWXr4B/E9YQxLyxvM0XIzAVahGYWW6l3
+FGYXDg4Mu+ocrC66dUBkd8YRbosHSNKlX0gUP7fx7pK3HFqI3SnXtChy2+BZXJhmiHhX9rqomQD
izQBrPf5vmKtLKOkJGklfssh7I7S9g+kmvP3C1JiZTCtwK9yytGnkcztsg8nAxpo+9aHKaSCE+Xo
ja+T0yuPH9E8q1sxXSOxN/KUGTGe7oan81vA7jMsODtamwRJQcUzgcOQs0/yOT5/tJFb35lgnDNr
/XB+YmvTf0xZsa4uk606tXm2LNspk+p22+o3eYaCXhYrQWM7RRjE8titUeXys6tyttc1sc/GqBwD
iYSjNSZoOpgBZNuRuC93Xde4kf8b2xRMUTMO1zKLQ24MRaE4fU0wDLAAQxFI5v6QsGRFvIdFUpAX
E+Ipx20c4ruY+pJyEJdTQrvg6ZnLl6SclQwLTwk80KDrBYnVvjNlzaewPmZlpLMAFxE1TViOTTUD
kIsDDR+rHUPj6W0x2kFAqhLMeYF+mQbjmnsnHnmgrtjaoWZyaMytCyzmqHvUDYmw9J5HKcd4F8eX
aIqNopuaJfB/FIwx/412LYvLon7TlEEsILBTdjXemkgvMlUI8pcT+ngJzWmaQZoe2rfkwKIfPk4q
3TvgFBl56OjFMpsWHa3+AUnjZEu4Zr2H0hBQ/rFjWnb1UK5JtdrMwr7EuSRgB7nQ/hz3kuupE1o4
rxVcuAuJDYWLbYXNEjKoIKBZ6NHPuvMAmNoDSIFT0jAitu2UsK5TTickoT7EVtsrhdBDiZKIuIQ5
uNv+4yUZ7F/4YVBE8gJ9Kg6bzENgevQYLBB2nqDYI1T5LCYSi7vzsUuI3nmayv4OqRKWvQQbFhQb
WK/KAWRA0eBBuOe1X8M08hA8DeqehBySzWwZp0lJPA9jfZK0XnqGyEY876Hh6WbXe2hA/7IB+1kb
1tj5XphzazvWcnHxT9+ONaxgNIegFaS3k+1w5wE0YqQp+3bmvHmFn0QzhjnB4kkhXiuPhmGRo6yu
VlKAOrF77OAiFq/iH5zz8wmmpTPR4lFZYM+d5VnvucB8n3un/E4NJ+F/4Na6kzq+WDj6cPZJcXxA
UM7YNwqYXuaKvtyu1BwzQ/Sv+LQ8elxGJGfWQPxmkH5qPWK+tRQoKErUMB+Jo7/cdU+fnn8jjTkI
ld36BS+NpyOPcuj39m/79FQZpUPduUDX/lNFjFHYUY1k3gbtC0gmqo/dO6bgXqAOsoAiDWh5Bq9b
KBKEeuDcKp1VzdMeiOme7E0ZjMzQLxYS0D8bFue651c3GofAhJgPKuc1+uqu0XuE1YjQ0923Q7WF
UOQFjAP5yiZlXXBxNvUli+3n+490hZNlZdq3hAlIzZCTvG9STIuWTpEFN3S3zjfBxKHf5KODx8GD
O0mSYEzqJn5hx1knv/KqzH4AZKcxGtZaDMnqLRCoy7UoW2i2uj8qY5x2b4GIKy9Giqq5dVfMtjGZ
LwWpGKHghIc7kR04bWfNtiRV/48xQIJYEI2uxQSj+CHgvprHPvA36U4euUjHJoOsWjvPlB/6tK9b
ViXiPAA8EUk7syn3DJRqJJtaORawRIFQ/ylk66vWOmZHWSH0RmWce4NCSEe59PdMaeoFzRxnubjL
JxLk5cMxgdq/Kn7XAxXhxcHAnahpyKQwIr/jNeuyOBLiqDbiJHf/rVBUNvoBD8D02J8ffscD6LXD
dfLJodifVrnGRjagO4ovNODIOANPzJfcIiw4NQLetfjwZzU0SAIQQ+DJ4TLCCkptlNlC4qfiO8PD
nonV6+6l1EvS2AEnrdLaZlQRXh7gmYjyinuKizaefwDlz0Gg/Xk2ByQziEoFjyrB1UGnLKV8kzLS
GrAHawc0PBBF473SEfXcpTQ8ksoH4+nc6xthtlFpNgw39Ah4MC35UuAJ38wXH6vaySKBXcQW/fvm
xnKW5kQBBPFdxq0h6HI4Ab1SULo+/UbrI20rlUjLzBiV6ge2pJFPHA9NLx/XNNOlsmq2PwmnwtfG
TINwscPjsE4tsDceNH47pI0OMM73cuIW8rc0NIRd2SPjZYZeZoJccskRyreejycqdHr97kxzQfR0
ntPONqt9GjPofkUQGXYoVUITTDRr2wxVEIuOi1vPblsakrP+aG+D9gnFvJhqhd3hVefbaZZTc5Up
CAPDEZJpjJw9N1k7MT42iydmu8FK9UkGLhj5GY2wHk8pI/OV6gt2p1793N5qAQwk6DkrFannpLRU
TZQd4Oz4RleblvuaGpJTDiobrv+4/OUC4mumLSQfL2HN+i/AOPFsCz7B1qjb+g+QG69Bo3G8yyh9
5zx1vGMps1ff4mItcrc50A8c50jVKgbJV2UZWOBhNH4GbR0MrYOUNzv+NkaqpLot1YdSzIH5fDHk
D4gDjGiSlHZ3tFUbekvq6Go582ucBzv/Ukwl0Q9rFE2v6fgok62OMKEEBbeSBcwXg8jp6TbpyZI2
vTXgHmvLvkR03RrGZG9eYYQKoEtuH2DO18vR3SgnWHvtVAdBbo+A3B1F9KPKTy+Yw9XiM8otdd0q
KOkJmAd/dU0FOO+WcXZBzM+KalsDqIYd6C9Sjn030yKWBDEC/jLin7D8hBe5TkuAFNzhis4ITqu2
JlgEYStUZm1ZZdCNvjvKRVbJSSSWCn41pQy0CqvSUc2bjAvlW24IIyZl0gBZlqBEbQfyWfjp21et
opd0leYFw57HQpbf5vRuWw/Mnnwk0IN1EjrokpmhT9qCc8EKGAk+yhfCtQW9MIMrpU0n745dtvX1
0i5/EIcsogEcWLbwDWhSFmYDOgijkKYKMqiToTHOOhGleiKAgNS2GMylu++7gdNDfBJRuIRcPeed
dhk47nrn+Kwpp2KNdMvnqI3gVHb3GCvHwObz2a9nLfexU7y2351NhoseMVHrhohHmPbhO7gOiDTD
OMHpwuqBzK7u10UgBPxKx1ax9Izkkjti+aolHszqP+9UrfDZNo+YL8dFZVnEWSfuItaHwUgKM0NA
Ja7J58TBHB4yDHyF9nsKtJULe1OSy6BsyCfFyfn9N5JUkm3gx6DB08a3ou+7dq3ACv+pWzlg4QOB
ChhF38+ISlyQXuzY4nwnFxaSEkkj+9u0hQTGr8qC1VZrwlN9VX+ph8dYM9OzeUevRrjgQxX4RfNx
9oAwcQDw/X9uRduCDqBi7wO8reFgQGVCJV8VO4DXIyuTgMfruC9cYTQQQfllGJAagqbmk+rBViT7
/THayIruxaINq4XVUC5+BonamL+F8ZrW23ogeKbURvLaGeyGRfRBvUwQMDu6wT8Q5C8183PixPFI
PbWUUXCUg6VwNwoXlu4UjtOM8KSeLy5liNEtJQQxYQ+9HGlwO401TFgzPoGumHp9AvNYRdp2RbhJ
uEvP6p3gp89UBHoDkgVAFHcFbFh3Dzfvi0cxPGXJN4ZpsEQ7iTrPvSEI2uxY0kslYsDL2cv/Plm+
ETapknD7h1KRek21PWlbpFww8B5Gp37Jk445vcX0uQhG3F+dKm+pk/LXzwKq5FsNKpQB31B2ihaY
oIkeN9qOQXrd/b22RVB9aoycGFH4gjEPpcIxFpOCJr484ExPc/qJbhH3DLUUFDyUSq5wutnKgypu
2EY1DCZV+f2wHAp8sKUaR8PT/1e2dP0IEFj+7QYbJ9MhY5JocerpxXRmAJB84WnPEHHKORVyq7Sf
bIOIjhy3cygF43CZ+edJyIn9nBcLP8xey+zs6CM8sC5CFuEhUo9k4YvdtDicvO3pSrl8pSnzEZ4A
IIwO1RctgnEY1XtlvThIq/eMxL11em1B3NDl23VMP+f0LdP9aZup81yt4KmkJyFx64rVrieH4Xhi
Lz4bcs63WbW2WSK9yANS4ilTEZRMZPPkzslrMkpa50diOs+Azv61FRvOZvtcK3rI1538HltCkmgH
eUA3QYb4S+BhbnQYQZuslY4eDrOSLdgS5LU0IG9DDMm1OFUwaa+MhHbc53TvVNjdrlWCvf8E6hdX
QU83LDLLdzORQyLYmzGyfKkWMc3n7MMUbuuzwJlAEYVJH6nadEU1Pd3fzGfaqHLd9fYybbNpW8G1
fhzIk5Gecmy7XZ1/jjqwEv6W+WfSidI63ZnJAMqB9tIs24L5RzKyRXL6sMnC77KG5iDMLd+fOIQQ
5oCLpsait0YvnVvlk8Nig1mhguZxjrePt4zyvJnhL2MZTHsot6HjKcwDN0WXYQyJNO2BbPmYhNPb
Jc/4euUH/z6vYfpphgi0CLgiQy93DhT74Wnw14cz9Ks+pgr0dxYF5pEsK11zz4DS27zJuubb4Nb7
PmJwQ3VTmptVgO+2vU8jaXx4CIqDBLZ3MSaSir3WYg78UJhPbvQq1mVGoFRXvFDoQNYVln0BQ+wU
kbm7ey1wzNYYUIcVW+MZsv3AbrAeDU6fdLIm89oVsvVpcx+W/2lNOf/Ay00w75n2rdMMxoxsRBxc
5Ay71g/Tr24reNjzu9rgMlpki2eN7/9AAM9kHaidOnDY5PoSSUXV/bMB+yRQkIYvfOKRYpi54dz1
1R5aXWYKsBMLhpVHlY3lWnaFNr44YPeCohueOc3f50xkxYWzvbSzJEIGwxjVu79MKTu17GDJ2vZ+
y/E9U7qao9SOwPFf5efSU+C/DBtfHu1l4zqpAuBL/c22oC2rvbcDf2t0xXS7Tzo7Fe/fIN2pNZQv
np1UlLIgDEZ/EqmFqsteehqnXkE3kUo54SRAIRkWG2xcKy8w9nqKsYRIskKh/Nr7y3aSnF3EjSTb
ZYyfi1CW0yWrbp3E8zVjfQayy9laF0TqEIc/oTeKj6pZaCn3Uook0+NiJem/R1L25eSwdjvePYtQ
n0xu1qWHFgFSXablgPDF0ZcUDxeo7aIK7ugEStk5DVaKBxSZLpo7GmEeZ/baMRGCUzsgZNjwpVx6
KhvkO/UGwCk/De1a/L2xOxDMUvwpRQ1zkBw04Mhh/GpcITpcRDHmkC9N3s8nbR7FURXo/La82O7g
k6srdkMOurl7QmT40Soj7gcVj4lFWYEu0hU1EpRuPcZY9GWHjMVaVgKOLXkAfm3HSZMuobT9StTS
TIlQEQUCzgzQf4WQulPyItOwbaEwy+DcuUGYlvW9esftJpcRG3g0rsfmIlOgVUAmdmv9oiByE8Ce
csRZ1w3qGAHUtUk/pH5RCTLu5UJHQVwspeUlLb0SwcTzTXdYSUstVz7XUjqPK+12Z8Jx+JE/BdfB
ISciT8bRsLntXYF5SaqCYU9DDKFVYSW2o43jykGNu+pVlphCPhJ0FUf0kMzHKsKNhnf/o6UYqJlV
7FFSf/DbIyABv1+30DdwWV/2Jf+hYkBco581XwxlQVhviUuAaV+BGv5pIYMffD2de8miOXSgaHJU
JUPgikosgGsn4+30f04qPJIwTYmI/PoSvfZV4hIsPHoRfpGP0zua7h15g0CLx2CJ9N+boVfazJJk
Mr30Q+uDrK1NgYBqxP67be/FpJ1Gut+hQHmoontVSy2mrI5s4J5A7nrs9E+uK4Q081ihN7wAhrro
OHrUnR4E/T+OF+dZguhXGn4O83I6781GGvXXkGxawV2CbE7D07Se76wu8t+II6W32xouFvE7M/2W
IuYyI3BgPRAcJANDQLktjoFug4naVm0TAP5khU0EasaSIWwIodYYZc/HsM6XbzK+CL0ixiEZDlr4
KbzdCSvIYiEM7SgIiETa7gk8ILR5fin7GwL36KaLyIyCBIC16WV0OjOPv4JaP9OokE22u+adIvsM
N6vLkw6GlHt2bU/AadjgxvkwQ/gsZgyGtxnIuclzIXji8Wksmu/lf5J2OPhOSglu00aBTBDGZzmR
rua0zMEez4dD9UzJ1a7oIlLyg/NCUx7QR5Pwre0OCCIgRPdhdXvjoOJmFyMbSu7OaDFoOVsaFn5U
DJddsbMOGeD2b4+zB9Aoz3Bwbs9YqsPFpda7BQ3glg/dk0FGB6ASz9WsRHmcJYkNsY53gEDWb2tC
BCURfwguzKHVE9f+st5OOSEc0pVVDXljFVSXHelRGJHtlShW5Jj+AZMScFgGCgbHffziXCuTVEoE
JGpfoo2FYM+wnKdp8ulbzOrkPspYBnBaJCvBqeBTvDM4b5A84p49Hzs6gTSu44MQHNoc42ceQGe4
ZdasuF8p01CdlF98E8942aXkae+/NHnWdWmfbwR0FMMhz4dcHIbfs31j/8Cn21cxmCXt0KvAzV+c
SIPdhjeugaKcHl4IgFk8wDqFg44mxtofRFTu+ZeXtUB4J6HwntgKOqA1Ffd6zqRJX3x1NIE4y6YH
rsSc3a9fMFXW2RgnGZJ1dTNxRoS9NrxFCCLeZQV0q7O0csKJ1lzanxt/LTMVoCGF58lQnGhqkih3
rjX5S4RzBkE/pQUrwpdArHVgMZGm1krxa0EkN6DxPLLBH+PaSbdQO7cRySFCnOn/j37u1XXBO87c
ABOOQ6Io3CQ9CM9xdGQ1roF2ipbtq+w1+lqBpPrvJgt6pyqbPv/cnNkvdZBh4T97wMmvpw7DCprv
0KEEci4avtMTy5IvSNBJc1rDfKBtO2kHPvu8uJBespGigTvS/V9pSQsXM1To7m7n4+GXa/2hgXpD
Xu/H7fnQmWHi0wSGndTTSclrfqQqs8UENDP+d71Fk3tY16QzRpy4I3QhDI6VVCvysav1JVtfG89S
blegCVLOPhDEybpyVqV9y//43y50Wehre1JRfMMCwNKMP6Vypsax8FkUCZ0f0u3Ngcse5WtzjtTT
h2KHye7GmdOe0r7MV2ShmkM2i0QU3lGSF2kenYKUs95R/xdKIsgzoU3D84erG65L5yELpEhhidc+
MZPntI9krv81bbHVTbwO/O500rXFPcLQ3SaRtoe8IQFv6j3ITXAhFi7YbtdadWTKe04e1vjIZ75/
Qz4Yp3rPr88WTosua/moeo6W9dwvkQE+jHe5new1nI9usFQwxct8iFJtNZ4grN4Hz+TCRgAVJYOb
fyfDzz+Y58iKUXqQOLU2IkCGmzc9zhmRN4ILMtCCOpXLbqAVrxDlzqO6nMrKkyCVKlUnsbm+DvqP
cFSSexlX/cuVZup/IOguigGylJFqaFblWk92XV3trkw+wHOZndElpkh4x75QHAWG7uEaCJuixlGX
5Umvty4JrtkVInPMQrbGhdMfbrcm1Ku0VfLxLTK+7TIVSV+jxCREA5ouLZTEYAhiC+LBbE8UHMkV
2oPQrefl9YwFi0WWY833PK8PFVNMh9h5M4yq4Xk+JFmhS6dF0CUZ8xFUVeCFAZtQblpW/DxLVHxG
XAgMfeCYPF6dObaej8UivoU5B5eCafWMNtrMColFuAjrsF8jINgNCdqGuTuUsLTgQik8Ndh8rIZA
vnzwbsHDVZ0smbs2w4uHcu9i49N2bBLsJLfwY/bNIZBIgnGeDhuA0POK3VRuAf2Yk55hXrq6nYkr
+y4d41GeL24jcieXBZ2Fda0PjZk9ZCaqn2Chd5bDSeShN1Wc+9kTteHXp+2PBpL3U6HPnb3sGNA8
FmPmXPviv2VCGXJgzeqBCgyNPoJ2+plkeMdNpmg8FIZAmWSxVFPeLV+hBvbKIyQr3KAXrYw38Mfv
eLcjnn2Qw3IPheTX64kgcQ0EBRL4WY8OYCvde0ZJjdTE7p/0L99JD4lXA2v4pI1MWHbg3jTL6Q7G
nboZlxlH1qpBfW5iyzE45csxKedLgiHzz/UOpu2WjNodjMcX5FuZfGccBgXNSIz50ErXtvogp2Nk
g+NFk/3ndalUkUnAQ0JbRAB25xCWHaljMXv2Yb4fxiVLuGlBwwrkZbL/ELW/AnchFvITuYDaayjy
lX4d1ug806C03SZmU4PXtTIYQT7b6KHImyjbR3CkyN8jns2LmS/vrUFBipqVsidiTgY0s8Z+lmZ8
Yfvl6YeteLGfIM/hPo0mRaRtnlqmlPvtSp60RGJM6u+/nocKsmc6jpEDFVtoY5ESoecuJpoGPD2k
ibW/Vj6lwzSfacQMNZ+EI803fPjG4w0a0iBBJH1TwZToYf4s7aiZ4tj9f4JMnNGNR4TCEEhvmJuL
Y8X145eYnguB/yoMvFctBywSuWdAzabFemleNhO9mbqgHGIdhGtFfG0qdgpEy6oqHKfcDZm8G8Rk
mmtPOi4qqCE7ULBag2uAkQN8gTBZ29AtNOTNYikZWUHU/TtUddmmyBpgKh8K4TXcn7iDYUcq5cO/
xdjzhCTbizBh8okLUOQaIUc2h8uY/GqHY9RrGFq3LldROMpamSqPCrbeca2+31GNXhwAA/dzvLBq
/+48R/XVKKRrgiAkiqwqBuNrkOj4B/cY6pX2xjK9lUimJnvgZxRzwxbeQXq7A+SZOrHAjZBG6fJy
6yHNS4RHc2R1eodqG5K+GTmh9cAFzoVbSoL9vn962zCzGv9YSltFPj7u4mJxfwZ8nlwkfYtXcXsU
JfCx89/n+e09UfgQuxzFJEnLz0Tpu5XtwXe23JMk33KPG2BQ38+abofe9nYflYcdq5hrPZAhLAOD
TXgjxrJEuMOljPV2P6ywo3C9iYWX0uIt9sGBN5BLajqdAG2y+2/o1A5RyBBsuVKlvb90HKweDbxB
u6p6IY4VhsyhSn2AtiHS2ETeoUwIBKdQRvI3fnc1t0qfkJNdZDfuEBfntPUkp7ko1wgdaeQullub
seKqVxFcJIANkkC+8dvVdB5miZKCvZyHWfqgGKkqBdUpEFtQZDFZ9mU1tYhufm4IrBvTZ+mvcYJu
9ZxnLIMkqJ7+/b8WUI0PxM5sbUOwMYJIcDkb56+9tKgjePTjgZdVT5PHuxnjbPNev1G8WfUD/qa8
XR07zDp3dG2sgEqM+dGEDjx7Q/mwdKImwP7XnNDLiJXgRbiDCNPh5oLrBO0v4m627/DxStbKg7qM
fx8gAhYyi2DevTnxaOhkAyUA6TR8GhR9wS8sNE3Afkvlb2ZpJ75+oyHoZ0GKVNdKcrClI94Qxd+a
cnUmNt60yym4t6w6D3KpJk9o/gGzUE35yYwQ3WzqJr4UhwAv7AWvNoUzheifSNsPovKd/qC5pSFz
8aeRe3wJRrJHIZ8vmdDWkAksYOkVh8MSdPhcgqEB4T/m3R4DVPMxdhHj+iPIsV6q8dsp86UR7PPW
8+qa//2w/xZdDWnYhmRQKXoSsUI1aSyL8ilX6KZxYyEbtu5zajH/mdHU4wYXPUhgFl0bIBXKB+T7
BYUB7Ene58/BwHkqyT8l9A5xgpZmLNrKljBZJ5ZEooQGO3cAaR3iyvq3sxbzH/bOSGU/Huu05gGk
ZhErjOugiDfb8e0aK7TJ/zKGONOrQbTYEXGBmW0ED4vOUEG+53VV16VAcpvsGm8kZUm2KGwmKUAE
c/EWL6IIjYBIm/dJkLLrkZ2WeQYDbPcWEzUAB8IJfv40qBC1rNp7iViAFXaMnsowpZTkJAd2ivka
a1A20liaRVRfnbAX8aH7fd4+8kX1bNFnphoZF670Q/C8eaDypfZe6AIvlu5w8yqvYTYeTXGYnos6
b3POJZqph+TeUYq56vFJBLKlNKunwIEr4o58knOMGQN72eRFTaIEVl7UsaS9u1j6z1TaL8ULWS+n
sfE4/d6gEn+RGarhZv9G2dMAtEcXXlgJ3RIyOLYlRe58d3YcqpcEcJuWJSwK7ELjG0ca9O5Chs2L
AsSmp/Fmiug0wZ2OwXzc5IbwD4JcFe5WRc7Zbb/SKmi/JU9MZ022lBWgvrku7bsu8sxriZRvxHY+
OTMDfRXYXZMP+RF1YsaRIEx9tkUr2zI3vWtCCYHDV9rYo5ker99JrxRDeyY7kzlrj0aUjAArFAdb
7ttKLKz+UevlZoQ8tZnuH08Os1puGY2uNIuldIyukaGiU6LZ5WjV8qCXUmgKUFBvKqcaXA58wQxu
RjMsQYJCq/QxBW3dp2b1OhiCOvXFbyVRGXoOSFfB4rnsVp3qwNyfhOcY3Irq7rlmr1y0ejOhtCOV
hrzrxwzILZct8xAb5yJ+A5YfzPSm/Lu7YYjqjDjuYD0RvxRzGSMKAAJ1xsFFxlf4ONeh6intcZzG
HwgvQN8Ev300gYeO3Nk/OR2zBJU+raprBCV6qkUR/oBBROG40xAsEBSzVAkgV7UdT22+iOy5vQzc
KjEo+HpBCyQ45sXfneagQtQXpIi+oIHNwIzjdZNxdhOAr+a/o6LgO03s8+MNNAc/kHSsNzGXDkXH
mfGjSRGkaq8XXQV+pH8jVv7pBKFPTKYmOlwybFbr6sMeD8ohJyeE6dzowKETBVf1XDOTZGMTVZdl
dxSltwC9kaEXok0MiMCDTW5Wxag8WjHrtZo8hPXuVFh3d1v0W5XRtQXYnfiD/PB+HwYff8JMmUlH
ppX+vIb7CsIv1ahAX05waSHXOFoXv8RC6LNZMiSfqwWNrvnL6szbDlDBaAEqF1GDwrEJnLyLJWAf
F9xfuoHujEljQBg/B/HiVeTRcb5ftFln2d3ypL+NaaF6GKfKVDcQkyKPeLZnoNT1p1MbFAenEfK/
ObZFtYsLe4exCkDrGXV8Hqb1y22bYYLyNpsdR6ouO0xYYDC25VLlhuhEPkVgvRGoT3eRgkWnfEW3
sAjGbIcqs5YntsdCra0tnRhXi8bt/gbMxK23v4uXYbHUWHdoRa1bPwnCWf4bqdLy/zaDPUIBewZ2
p47REYBJDt5if+d5y91b5rdpL7/ASypY3kX5B08QRJuYfa+eGrmOAja7R6nT6L0taa/i07X5wUGp
TnT4HOvb6tUt/1hE7tyrkh0wJAxom5S7bKl+YPwoNo8d+4wjvq9UzNJulWw62/n/AKM4eaeImL1+
32UkLZv+yAR6BggFc3Uoqa1aUqfMoDuUb9+R7r1m5oz3ia3jmvAcOVdA/qZyiczJ+e08XUTvnIZl
GhfN7qPp+MRWGqnMF8POdXrnr87jBELZJGE6GbAa3omo7d94DcXSGwjNA5Df17ZDBuZMIxy89/AW
suM3cFmLK40fx6PeoNaNDMB4mdgBgnaQocyyjbf1/VjGK+RnW0zI98xA2HSLqoDC1UbhB9hpIBNu
SYahi3bc38jOt5z4vKls/IxMG+aUjMAdnUiOI7h8QReljW6j0zMCCW308WWQgf93el53jV9kTXzY
6/xCLTvg/uHnEk6pDhQPQnTkXohLcD1JGgmcZYxw9XBK1U0/tfyOZzkfUIL5N2eJY2bBccZ7indj
mlymYeSl8nAvlYYYgXzYnERMUMYKHjv/Fz/oduH6BYLcLYzAiFGSHVmDwNBJmUh1fA//YcdgxRtm
zreO/y3mOUgYeYj4qYCoKOmNE7x7qaLbVPqCxG6mkD10XJZQNvS/rXmTnjkitk3qIwG97qGR8PFJ
I6wByUjo88jH+u1yYvykUGkvOMa38OLKuABR//iZtBzoM6ie1kQF+5xZECHo2LbCLsI3yHJNEDDs
P8JdFf6lxH0KFxX4yp81Fk6yCtNdaMW02anonjnhkJ1aaVvtuQb6nT1E40C1homB/Uy5BWfd9FNx
hgk3dh7B6t3GAkCcz1hX+MpHtU5GBDAU37Xc9PZH7JwRCLmQ4nSlsursKA++Hqj7ixhBNSRV+REk
sm4MFYqHCeHdOxPL10LhDRtMFSKi3ERVB/tMUq8TjvjbESU3dBximCQp/8WS8mtm85pUIsKDaAe6
mQ/yO/Odo1miMMsow1yNpc8blCEEQNBK/hQeY/Y3TGc2+umCN6+MhFBJe335kfuDKfWOEa+Cr+Tp
T7/VMBOzq9Ry7FULNDvhCRx8kWJwdi1xCfvO1aJtBrL48KLGwEbYaVJDR+0pBeJBVR4hzZljEfJF
Hnh0xhDermZwX0ygwy3C2QJCTS+Ehu8InK1IOYruBH7GkkugFhHSVg63cKXHt4zh3kuyVWcpfexx
lJnU44cjDRDvH9g2ZTevR7SGXCD+2eEWDZbgHRzl9ag4tllyhDXvRgegjJ44xYP5Ghfj9ii4V1z0
myFEKB+agQ/LhL0noJ+zOKIOH7kaP/Tk6svoIAL27LZ8DlMgdH4u+EsCrtcDkiue2oe9rM/Gkilt
TUbp16EyHu9aOCa2yRYov2rmQ2dh0LauIR2Xm+6kraZzPcGjqU7tFBFpjMxbu8bakiMFmBkKKWzl
/PxmPzYyZeGvNKT+TPbzTL3tZqmNAuqH0MoXDLLlMocvsie50dMCnUWe/ZIcbdQA/hh6hm5w6Ff3
VPb/CXjTzCVRFKWiZjdmt9gX0LdMD8iYsqzQWTwi26xTBZM2//dFnLPCGmzxWEHZpZF0yneoi1FJ
jFqw7gjX1o6xpMRajX6sGO3ieFUsuhCzV14LWfmgeuAGstDzLLtw3oUljD1yUJblXg2aJOWANeN1
JlfOsTwd4gvGdv6H+m6bsMo+uLFLy2aM8C3Ve/hr58k2bO5ZZclPzXg+6rWn8CAt1LVYZ7dnfNY7
DbkxOBtDaHTdAWiLeg/y+oi3EcGM9j+tHX9t9DHkSL1SqWLOdUNnZI9hQIb9jkud9RCg7CHOtbUn
aAuhJQ4v0Lbffc+BIyskfUCkXoqbRn8A5QdPFEiO6parGansRfOI8z4Ow4XUkCjVwmYkcBRRzJFP
w+H5cKY/X+/aokwVj1hrQoK8sbBCAqn50nhNxTUxGUk033sKdeSL33FnDobvpKOqA2mwuE3dCqUd
L6F6YH7srJm0MuDZrj/Ke6CmaMGFP5UC+sx59kYJyeM8tVM95x27Sr8VOVHOOZuipC/EhCh6kXmX
5cqdlIZUseMltTaFMzhDfu2jzUgge/0Pliu9FIEJ2r0vnC91CRqPjyJzcvOmtwuULqeqPG7rexCu
1VKd42Bz9+TG7wGoZOVIs6WbLcFWxfZjWSYXeY18pLQNrd19cSgKs2QT7SHO2gi1C0r+NVtGzcRS
Wdaus2taO0H1+WFkw+DIp5CXKvTnUPT9ZRnbl4zWrNF8oUR7P2uzJvRLetGZ9tkCgk6r4WWjBwPR
SqVnCnySZ8YJzjpCQCtUwINds0CPmQFXz3h2hxUGOUHXs6PKC4dlubA5B7V987EhOl3dvw7jz06A
AzIvEreghV8nd2hgIMpTBKfv1NMjDMnzqxRgQut+gk3FfdT2tjT5hwFiscbiwAyWoNVUb1aq6+Cz
drRnb9TiYmfRQ66YSh+6TBC5TgxMpWXeuQrW7VbRz8vQ2tY7x7blu5tsWy79BgHRe7N/xFJtMS3E
1bQcCtrZ3X7KNd0dOh2Z4F3FQlLkgRnIgR19PsS/e5ohazyX9G6Y6bgUamcn6Biw8cbONHmfvTrj
Jy1JwVNecAB/gZir5Lk4v01Ydf5pKvig3ghuQOl0wawXFnNfPrd6/TQaoKwxmn3wIP6XFYdRPFwj
8p7g0HDpdr0p+BAiXMhaGItAMZrLwYeWj+UoKuKr7K3AF4K1+9zotvN4SjPFV71W+45JqsOWASmB
groXr1+4ngcBLOt/VvGWQH6oIGftUO5oPcW4DSvU/JFiW0R/qLCycfC/d11dJnHcFBigI81EA0J+
S9ZfUdQL5IlJ8U/RUsDTqD6zHrr+atk+oQB97O+junjfpFmEl42/wQWSrQah0BEBXdFh/BuULMjx
w18ZfzkZVuJrVRAX/3jzI+rYcBrXrGgWMBE/XcUj6FBNozcJhKoIBVUABG4hH3SHrwzmT8X+q2dr
aCm9JFfOS4v4zohGHLMUKgyZ5usT/54ojUBkuGcQOrSfbsSovSFG/t9N15tmkiIJ+EsVVde+d8EN
USoSh5el/Le3641zFHX090upHoxwgKycRHZ9JlY/R5+C7+sBXKx78BRfoCk7nbR83FxfDY5uKCfj
2u8x1YEETjKoTc2imo5vksIedKIwLXmbMj+2xFFvYbMR4KK5TfelzTjR8xLscRvaG8mdMbCjN8OI
aH+2ZiAz1obX3RGYwjwd1weM6jaBhV1CFtQPFfIVSFIGKGAgaarsmu6KLxHxijc1xvIkeYDlvupz
CxbQxZQRBJQSncl9XDGUtsPLPuibSDsTjOF8qgqdjaJj1sftIF9uC3UH4l4FMQQUyvfJdd0FPVrA
9SRyq978asQ/n4bpKm3GUxHvPlrS2HY5hUdUKvWpTDfvMYAlZ0+huE4grfECxAmN3Ee6e/2l8wnx
P2c/FEvOgV74MGJJgmi0s1ciaw89Dv26xsP8a+DB7CjL/XkfW4xmYKjxUUVPt0ZpE6PA/MJlcKCf
XryxNC0WPMQAHYAPj3I5IxztuecX7E86WVfIobZ0iTxJV5GCbJOZiFYBQH6tfGt4gLmYBfoKYug7
OA/RAE+hLWSiPviovH1LlypVIfF4kX/VJuvdAxc2RCob7X1Cxk2jrzP+4ZTR6y4joGMc8BuX4W7Z
Mz0kFbnwivaxcrJM0Xa9jGXCns0ZTb/LOOEMLwT3A2XjUP+C9UUMwmf8awwJKNI+4hmUFFfTBVwC
xFFnc94T6gfaPvoAXOfat2waApiX1T9/BXsniP9mQHUnAyYZ760ucT6ZopSlJtgbIBUR0393wJ52
GgZjMNMqVsfvbCo31gfm9tvhqlaKwi6CeaiTx30cQNlax8pUQBsS7saFKcjC6LX5KWt2i/3xs46u
Qnx+53IXDLWZOWwx5ffhOpflyQhTrhGvaewNVjxsC+onf0MQ/fk1z7FdK4HHHScqKMBXcnWdhbeO
g6SkSZ3idHQ9/xIU8EoC6Nt8Aq4seQxM8xtAZ/sa3S7Bp7hnL/J19yYnBDag3hRtpC+RGjZTpWm+
iqcrmosto9e4djlm/YnAfcqj9fHOZwSSYV2YjJGl5qxz4DOAPhLlQ1R7nIV9JGnN4BgZEU3MBxfN
Hojms4waA5RatbKvXG4Jg+CVCN0khMpUmDQeeK+AG3uPCE0kt0K0+RWtPod6fk+ZW/Sf+MLuJUFx
wrk3dCz0GBA82ML/v6xdPkQHf9u/kNPO84EBaAUYjgp3FVbAc6/vnzwDIq+SyGz690CUKhiIjt6l
TFmRh0Wio2IpxvxSjrP6mAdN0fXsuMDp8HUC5zX8hAUrDhNFKVScEaUwRs3X4a5HMVmOTu44od+O
U+LnCVsRjKMYaiC8ptzSycq8veUV4mFXU1HvpBJIAM/IeQaejNMLNOHIVJOM4Sz/89xw5NIOyE6a
3xM21v4uUf2HIMcBLlOlML7UTMQQ9WeEtphF7/QX3bGlCXigQ6s15CemOTHXRUy8pTuoJ2coL4tw
uyth2pAzs2Z8IC88ACZH3tMnsKP6FqgPIIjg8CgPmYN6A7te8L1E0+HHTMqA3wtprdu3HIFRCzMH
UNIdrhj6tKZhZNB0hXAf4BYklBg4v4fCJ+sDwrJvXcl/V+oHjGF8IGMh/q92g8gjgTTF00vii0a3
h5HXDgisa7xc5PJ+wfh2FCQ0mwtsb42jAjBVYPFUMamFrJBi63CFs4y4i8zF6hOqOKntcOy8Fjsu
dKdW5m3erBri1g73QSwoXx/rByAz7SBmLjvyHg8esNSV4vn0Amcu8hPe3VHV4W5TApREjwHP7JBt
YaGRl2BziUEOgIbykIUbN3AiArBPyqlruk/rEl1KFMz1ZbVwPZI1pcFXkCJSSC7JHS49kvfdJKJw
w38O/45t+dEd4nJdV+s+Wr4sDxqFMEnArKNiNyanZw7OL7bTpvdxVRLWY8ejcHRFvdwTA/S0WguS
JeN+3NlitJNrH/ViZ3d6sR5VtJFIKExkn6TkWEO+B6vjd2VwdmtRuS22n4Kpb5L2sqJjrw06RkLj
rSQ1HGyhpUDlkMrKz+IcTHLtv2IKvoFml0nglBfB9ZvrGjwDq3v+oB0z5Itk5uymzkdmeQRd0JzH
d5PVv5wLSo9M0ZQWI26jPE2IP7ZL8v+WwZnawNeIY0b+eJgOVrpROHETi+iDmeN0Ho29zn9X6QYO
onGQiWKS+JJdBK2gPb87Jw3LTLlay8MtTVvE9DNX7m1G1qkoKu7NnGxckw2/5Nrp8JteE+VPEhaj
0gpQdXepNVwkm12hpQGiWDzCFeI8VuqLBC1nsOXN7KKOSxk2eh/GRvlAuIz6sOu7Eqg/h203IkGb
65BGGOVqM4j+FjPCbcBNX3pLsg32WqkwMfWXUZhhyyD+D83zGGqKB9+cOwcGSmEmFqHepdCZXQLe
QG+lVRl+Tdoh8vgl2I667rmEwNIfmA98Y0ezMJs7SBPrAT47AnRuBNR7wWe2v4xrBM8XXwBLyC3b
UajfKQMQkVvKN2t4xvLu5qRlApJ3Tu1K+Jk1z5r1wd8fNtIWBkMqW1s79yQiFxt0r5azDx8cC76I
/gYUUzDUBWAkI9dAXiO8ZiK9gIeQe8QSJP/oaXRZVuXyslXsKV1gQl8b5Jy4kNTDlqVKPX7rHIqi
bs9aB52cc1Fk7rHiZ5frRocQBxQB2dDt171JNkpDO/W33QtoEtmDeqFCaXhEk1H6FUraqfQDdiYM
JBGG7SZKJJv7V3YJenbv1eXpCYFwlziI33B4eRC5IC6B5EYLIQ5gItfYs2IiK3UJx41jdujQlU3N
v+bSLwvNNDlNGSPGO12G1P/4W/8E6j2+I8KrX8fBpOJUGMGauM5od212FjXk86oxNXSguS1vRrgc
MNIPywm9UtiDh6MpQnD1JUi701IfkAZ3D/SgN4J3pjyLErS7lWRffcJdjk3BQjMz1lP/R4X+B6jc
G/rVQ5G1nt5ay+WYuYPS13Z9ixtOaCyp6y/D88E9VyZlAK2lsxmhCxoUcGBlIajUwNLEHUGkIyGK
MDJfave/glRqwK+dXYfmui1uB/LlPknWTc5dEpgJguvPxjMaLWfc3FZMqAM4dFdE4u2qk6jvJRpY
kd+2859CiPFYj6QUpyZrLU36nSHc1h/64WFWsOJwj2tcxgGQh7eCKPDoriwAXB4WopLFpG41ED5d
7YhJEzI82ZASmPj73aqEk+4hsmzAfTHqvMnQhmxs3HFoURV9Yxu1XEE9+3mLXC00i2ywQZGYtLYV
fwfQx8M/oXs4M+kHOo0PBd3qTe+wB0OhC7CgsL723mYPQ95OiSZbsoneosZHeMuZ4vPko22jqmuN
sp1JQeLr5NA3SCwQmHuFQtIMwIDcPn1emsWBWFT9oqf0b+Lb/QK+KQXr62lyOw2vD5WSp8PD78xm
wtdTJJTuFRY9k8Px8ZzHR6m/Zokm0FaosxPKRGG4IDQBFF/ecHxZlGgPci4Q4IZmcxN89yfHqCrS
I//vxcQLuHuEiIdAxrU5p7Wxttz+1yv92VpkswukV3elDttf7zcN82Yt8CgZ39xLf9DW+bHmB9De
EtYnnc72gH//KMhmb54gQbXx5UcISvK9fEWy3OuVGA0t19//UKkgOlcy8gt3o50qxtal4rlvtzrW
GLElqLRS7qKUQ9w7S38zvN7KPOeT+M29r33bsGUNJdTFOJyAxevY0P5My7mWrKo/zvmhlTXVqm2j
o47GkmYDz+fK/X4Qf2IgJuwQrUbvsy8ah9NFZqSH/88pmAFlSUP90JqgHO2qlc/UjGs3yV4svpmb
SxY4tMijxCf2JXsd1KGBqAtqURbe91HR7I8QCSyhOtG1cwhjDTa1RKitwqU8EBTzcmkef4oJyCbO
Bp70KBYNSBXRZkm8qJOan5LrGdIR/jUYuL/Dx5Z20DdQIEJjb5sQs3mNXJ8IX85OY/WCAdtsrFPL
OK3lp5v8ojjbg28/+pCDKeCAEnpxh8f+krXjgexk1kIVvKpggSWC7aGO6VCdtNAjITRYGvjdtRF6
MsUjyonv+9y4vmuVzdSk8I3J//H+wsPmsa790lKCul7fhNGStERkguib5RS3kElYV04/ByJUdrqr
Pt3RKs3o2Cl9IC5kYh95q5IN9op28RnLPHl5zjvJ4jfJ16H5kKYIMQxsckxojpPwk7ByxkBzyiRJ
g+wHozE4c1gL/sU4zHRgYeQy5FWPranSBl6GpfKuxLdK8N2PZP/davGL5soDjXg5wQm9r6K6Q0C7
YrFpac8o912zfoYxMf9BczYy9a2Si1lPKTccXkHV1PH3J4qe57f8N2ZGi3GCDLrUxjNYqfL9iOAU
OLJCXwzOBL+GekYxUyfsQHFS8b45qoVts11hl/TTYtGks54ezPyOjnjJaXI4Gcle4xdAxaLXXcKW
k+fzMGszhp6AKNqbhcYIb2tfiw+AyDMfVWOywW4gzSZ8HcpE4rBTSA5uFATgFOofSlMm4Hzo3hJB
RrewcbqAfVSLuUp07+880QwA96WFR6jyukBFyHRffQ996rQXn7MDWOt37ZV2SG40qujzH6J4dJ7M
2ZXIabmOJ0LrJLIKC7bQMFYlG2TuZ01mZ8BGiepMDTcIh67h93xgQttx1QkxKoS83p89lYQxA/z4
zQCityv4wCYmuFf59gFL6Ehmwiohkf7dOlwJy31I0nur/juzQ8dZV5rDttEVLS5qeItlAs9GbGUu
ZepqDUn/J3Rd5a1xLPWGjYrBtRnYCt3ifAMIdJ3uQ+65rOzbHcZ3LhM/sO4NlBVTfaMq/Ew3emrR
pVeexywE9HgEVjo2ZG7jLthQc9jYWEH/FqemWFPI6OYReO2Lk0zItdD+vhIOQGc9VRUCs2DDOvUb
V6dcgtlTky9MSIfLAfLr+mwY80D/83kc8vnTZhmDueOZEaWckK1ePcYsqHKZJvgpYwDXAHlNkxNg
GChx3W+OxpZ3slGrZu2JAPDHgYTTmpkGrksRjYRJ2UvKWQR835XZpzti91WO6GyyhkK8PWf21f1Q
sUICiEkr7C+AdJUYHBu7i4m3sIub0ugOScmzwzN2V6TPcETcrFbUGy78D+LvHFdDuizBQv0U80o5
lXnYrLIeTgsacZDjZ/8xc45o5NDSevNcdqrGze3nXQXzCAR3fuAKw55gP+jVNizPhdzgIppNStsP
v5hFHjXgouD+BBxBs+sejejmVNo9g4fPiBnsBCn4aAgJeImPYpiBUZdwAMD61RD5K01cOQvZmFQa
ZEvmbB2lC8iuJsunWhQQyl3O4jVQoTTwWBbv8CkirR/o33TycwhhVho2CuMB+owAcXNRyAYHUthK
/NZVzdipPgJ2biai/FAaXdHjk3O8OJsGFvkOa5MF1zIvr5lC/OsO4ZenyYblXLoiK/DX+CZ1ohBR
XjI3D8JLyX4iWoAZrZHW4BsghGKe7nqUpLHqz9gapHKxoGCdeIp37DUab3TkxkyYIr1aNbylUXNl
SbhbJVHk6HeUZ202SBaTFRQ63Y6Hl63xRutEjgIV6LO7Xgfkuu1QKNN7XOYZFJLtAMntj8SmcDWQ
M/kDQummIuxnOT8SkX8trr3aNKu9AhzC2I7uJ9+ocYohD+TpXtdHH9yw6gdUZG/ME5JBQ3vCQV/6
a96646CHNI0xvq8QOl077OyZhQU4ZG5Td9kUDQ8xKVkusqcT/yRpkVOuLevtPSoVFbmWUm4R1suW
8NOBZqn6CJp2YotIL+oJyo0i5EubgFfmVQ/u7jgnC+aOd3pzBe31oubKTMSSI1W2zD9ab5rS0HST
s8dfqiQT+0erlLzogLlCQmNDpd6LvKDZtMJroaWBEiCvDPOZm4XNSft9q7SJYfVsQXACxzeLufTb
USCY2OlGBOVyda17dpZ3YHiPho9bkhexK0ZUA2HVA5KLM4bj2HN35XBJZCoiIQC62FlughE0wvoi
/iH8JOyxP/kr5PmA2AQTBTcnxjKn9rjmpG2Bd8VIDgOxmue3SsfWGuMD2XXtA0zTETXod8i/TUMw
tgenEhFPoTDpjABFfaw/8U7pLDAdh1vfkleYKMuCsFF7ujd4KchNo+ujEi12PPUyjlxRG1zxjatk
XmmdNo4ICSUhUx2ps7onVJiDKAEI4Rf2N8z75w+1PINLc9b03EeF1/pGOYfNFxJQz/OrN6cBV8FR
uf+G+zkRGGjYQb+cK66JeGtLs6qvp5128ky1TnzP3+3x3Ra4T9qCVofZBiA8NyI6/DguCBWeAonC
9cQrYm7MgZpWiVHcoP0+9vpd2OzpdhxMRj2Sxvslxr+KDYcCHdTk70UmWHFnep7S+0Coie1yMDhD
Z6+MHJE1j6GgqNLlXdqL/6vB9QOD31mYTgQpZPT6fcMH1MB7EMCi7dSn6ZFmpRUPxpYCvxKAAf67
KZZg9XHjUrRqvn0NQaJxpYr5u1uVNQ7gd30tJ95DFtTU14uewPPrONSKK3EbwHX9/RGJNmBQWil+
2k6CI6Me2kK772U0oG/YAWi+bptk1YqBauuXGt6CUuSX/+AvcqO/71LICzNB2S8yRgJGgWrMl+tN
yfnHmoAbJek8PF5aNHQR5X27RFEhb3rLcn+wcgiqVD+//nA3vcDo/Lisx7hj4ezitiO6L5HVAlBy
xLWNDpsq+tSClkunBtvBkvXzgBBQyWM648juEFiLlhEbyqoigOjdqkI+SlVwq9l1UA5/28FhQdF9
kHHTQ/VqWX8iRpa32xD1HG8lLXOB2SmaKhrs4bdxJd1bEndsQYH8/CRcJUxeMkSl5n7hkQKjtJEh
B8T4jV+/kMZHiaUIRamvbDr+zXhKvz0WhjX6gnhICE6Uw+Jqq3rPE7SYJ92cXQS0wBP8zQH95KcU
UGQO8TIb3FOtM3NAnX+KVoYX3sRzhK01vHzkengRE4mFDDQ8/0iq7KJiJhT0VNf/mFQqDeW/smmK
eDBjpyprSLz5P0uqJz8XBKH/YCOmlBertVkf9Dg0MwjYDvoRGvRjl7zk4dd8lLknnMBYnCZYx9ud
Jkj2lueC9RsB1pTi6x0cxqPBKpAVZW8Ts+K+XenMSQZHrhzZpF2Gfw7HPu9F8i4M2vk6bV44b7+A
g/Q1w1R8vO+yCWhEdZ4lFLZvFG0wsjwkZyI0KTaFjB0ubwvj8wPc4UoeRKz3Qu8bGt9qn2xXwqPE
rTpdekJeO4zIAYPnnbxkVHDoQ6WwzWc1IhSq4Mv0IbKrFRlh4v1zZH50he0V5wIcOlMhBVuPzHs9
OhW8FYKNAprEOLUZLfI0iJ8vItVAN03A1fA+Okz3S5YoJjIzymzX46c2kHr+20sgvOBS2r91u5oj
7Y3Ay5yhqY/bBLXhFEfNzYCqFBnny5h2kbUVuoRGQptZXCgIQWjFrtT88ZQ/pDhh3cllhLsS/+IC
MnxIcwweuOwfaWOJPw3DhVC0bqhz6sDOr2WiLPma+jVRRKRet6p8CIt/lA3GrP3daxVCQV3ITQNZ
uzpk/Sdy1TFcGdl+TT/rovjlm7kUd6m1/b3v6I4rlFwakD6mHAcqRUroMf3dw6ymzILkCnZ6/F3V
DoLy7xSckKH508T48NIswITTWJV2Ei9MqpYR6x5p7kiP+3g3diVFFsQyl/cjptXuSF3O3JxUNjHS
duWXwPfGAU3E8Tr+IyonSIVyX5U6Q59dSJn5mHCh5vLR9ZzWWFQV1iQn3YrJGoBvebxNftC9+JYs
tsmhnmi/G8nUM9ozprOlWIC6230d8NZ+Q7zyvB9KWXS+N3a+21a6k3QUyHFteGy+WeKYSkJR4gpj
S7Hb+5u6L3t5AhRkRZ6FOfoMyjDiYa3tfWmz5j0P6LKu8r9df4PZi/hcG3fqZCulZsQIk9YUfNQB
pWVFKMa0y9NqGE/OidW231d8geoD/dj8sy0Tck7MlOMtJ04cahJJyVqNX79Uy+AkX4DFlOWsqpAW
g6RVMwZTiuNz+9a7aGW9jo+hO5ox5P6zghE6X7lFsgNVX8E83SYKWKZRJ89AdDJWO2vivbVy8AkA
F2ksPMAozuQKMV6WgVWW3s7vX3bNOASoGN1Wtfuxscpov6LgGOT4QpvsQCF7qQxBAFA3S+HMGRJi
4nGmvdSZY5rHLPnDHzYq95cKB9CT7HUD3OQ0CFIjXYFtoT5YwlcCafI4/NUrhMOBagJkqJY9S1FF
0ayaASwAZubxPkTNRvJVk75LVveYCM3i3w0Hzi0g9PWwXOYnK46gnQpDBxrlDrKQfj6wyWed00T2
xGNxz9gyGRMoXAN+w0kuIE7DY6BJo0hMT8k4Gpu0NX32RzMqwITw8xuJbhdVujmbGpwHSeKBRDTp
9Upof1npyXZPPf2Jy0S4WPICC2v27yCZ2Wt6P0QKOkNi6J3JKbh9GnK0FchTFPmEzFx5kTiCgsOm
VCvWcGmgZ0QnbD8BR4L0DfuQKHbj5G7txWIC0S81Con7CwSixo1wTugVbkIoNz5uEkb/db298utl
3P6ul05g6/fCeiM2fKR4S3QM7upM+U07KKfRYdTeOUapfkxN3zJeYxp0hkerlrxOF2V0HEsALYtM
D14MrQsHMNHE0Oanrn6ILdfn6fJS6lA0tAo/+Ai09kBw8Tw5OWPB+P1H4XMkscitzom4a3EBAFsa
53WGX35dR8wNtXGXoPEcYu+5nX9/awQtAwE/gHEs4VqtMj2R56HXATPIHgQsRd4bO1yRC5FGrYag
rZsLeEo9HXAXqtO0zHG+gXgEydmgzxxfg3Vz+ZrW+dB7S3+ve0NiCs7pZQiH8keMVtKVW9OLk+OA
d0Wr0EDRancYEDVX031FIQfygF0k3MEqKh1AojfTBYz60YHqTt1wKzFjs7WikryudqSF15Ms4qpj
YRQvK4EM5me8pc8SlZjiy89s2i739QhnMmLQmvvL/kdCu3mgcQAchhSNvvxFhRlxB1txDDalhFGZ
8ZCks8cFotcUC3C/qTFYRdcAHoiaCmmXcGveXqAvFtMUje7kVcDdRJyhyrUegJF1KIUKcCrwhqCq
a9r5v6UeL7HYUCVKv4ZId+5hpjtTM8Q4Lg6/FG/LJRtm1Kr1tUE40UExT3yXHOtZscYh49vOohQt
dYysFuKxqtFkamvqfno3huUGD1t9yPMzC2p53vUA7be5TyBr9HZswm7oYT1VRyEXPINLYhw3wiFa
ljCiczC2ZHXWTZ+YugmJ6y9Ru16ZyP5h9C9ilKOqofApalfNf04kUr3V9eoXoY5MwzSfL7li4rkZ
Y8cYn3V1Z3J5e9rZvH8mVueilsPBSztBhYH95yEKkxpDaNrqUWDv64ZtswAS5sLx25CaU8CU1+lL
vL0VWwPalQ59xwTOBwf9zPAi6jAKMySxxb/4adg8mifx4x5kqTtKiIniANVPn0WfcSbmOBI/XX5V
Z/FEWNFouqtwA0YNV+3Aw94A6LZESnWYYiBxlpbbKd5hooQ8V3ziYCmpGwnXCrs31eIVNQflyRhe
HdAAYMi6o4HW/aqceKJDbXdyzqE/Zlz2IWD7+uPI6wJg8VdwzNZPZie5X/iEroMnVf0buFRB6vsS
nDjJLq1D/zbMdJT5+ZFhQ3N2E2/obU/3SYWTfNz05bvxTSLGgxK7NE02plQab7BIJz7ujbpjyYg0
ByAYHOY07PqZ0bQcXqwj9YxbhFyoF4+KELCNOtKhvk0VtHvJaQHNMv+IgAMz5pW9zX8g7RQ/T+Sx
cj/XlVPHZf8nuzoQ1F0ucqEh6ZcvcwZtleBKq+fOSjrrsUFwftF6mBTT/EFlCq8gK1y2Id3H9mzT
48Sm5g8e4r5Ah/6gZ/uPVhd4WnMm0gNNLtKt2/Vg43s8CFTaaF/3vtUC3x4obCAfb4INF0+5il5g
e/3MrGM4cCwUBqbnbzLNbLKDM6A2YiFyMQ0/xc27SYvhro0XTikZZ6j+nUga9xKxQCF41qp1T2HI
zqK7py0wpyM8a+0xTFjR57aN3sziorF/r/LbGfFk6AxBe3gFFxqgmzX+EO4MWiFmRIt3OMm8bQpL
Lp15PayjrOBcOphyRMf0YGXbXxEkSWBRDdh8GVf93NDQpzveeciMKIOAADobczyFL86YpuyM3pW3
HJVXxFaeDFdreT9igYzOrS5Y0y/4Qk6CxxFUFsx9Py8LW0h9LBWJ62a7WhYe3q/ROduXh/dSN6xY
hUG/uj2SbYMwfSRQlgHMsdEL6g7Q0lR3p9Go1lPDYzjzxZjsRYnQlzUxPdmSagEGa//5Hg04b220
INQ8qLzw01AeAYJLeghz8c5j3l99gP4jOP28OD0Q9v4mK83r+vZcWgHD6R8nUiZzbKPw3CjYk4Ha
wYh6AKKyR2rLQ7sDSm1Q2SFHdNFpyQkuL7kBvO4PGrIv2uue7abJGe5rr5LOoWscSmKmB2P90q+W
wXd8IHVbXZVpiWt4VMUHW/K9dZR/WQI1N2Gg4cPETYavEL4XsC7Jxa4+DUICJAfDc0Sm8koYnara
IJoREQ6zFoT1tHlCouiZrOqiLvmV6YBMw77Vyew9k26T1hgo1Ld2YGmsXgIAwrYw35lh66eh3nRn
+s9w6SfETKU4dlymsskmMBKTHazhE9yL2+NFJjSuQiTYUHwBBOEFu5xEqIJV1BfJ7rHDA+3ZQuoz
JKpXuHhTrm9GtaWmMJNGEYBzTAzoVu4PiWT8xjRkpzjtYFPThzlyVGo/Mi8fSyrZ+s0X5dM58i01
mLetPT0drFp6TecQ6HbzzvWXOPsulKU3pGXeFBQW3dc0fFXj4N5jDwTT/Be6xqLhY2cA6s8hvKa/
9r2eSHMjBCYxPRBdnOWWgVjkz+TxX56ZZJ4yzdZG4Gk4Zi3cjF1aodCTJS9jQ/QbcDuTp11auQwR
jlufgz/Wp7vlvWKrPlk8taw8PVPjwIYy7TBNy5RqnzvMA+YOcWKI7+3U2GBBHMw14z7W0HkUb6O+
HBBSKxWP90cBTH1GDJBDPKq9LTYMOwSdHNRKvI836W2unfrepbpnY7FNLrj+GJUzf6xLjYfx7KBx
DZizmOoww8N+/wpqubFKE3ZO7zATdm64e5EDvEpSTz5UCA7KJaue9mmSRsBvcWc0heXjB7X7pFRH
jaB94bkRnaUcOpkAq2YTyzYB6EJddhH/kklUsb/lRpddf4wGJ9JSlE06UsYbZl5dLhyioX9TsHeV
zhz/r03xJXFO6MIjAsahCAVCMsa4SxAn1uVlMqa3R0EjNdZ+Z86keTVPqtov44lNw6dToHqeldT/
JM+K2of9v58HOvhBl9KfgiAy1mr3tsH2zkLrNm+x9uXXFXnAO6rkM7uoyr2QKER8YmNTvmQAsFsz
e/UncC9fjEphpp4lkRbzalKQpXba+h+S/Cr3tKxEs1lXP0HplohoODiniFYFtNKL5P8oppA4v0hJ
lZl2zW92eNXThFjd2JX9Ygo+xUqAiLFj8f9bvSPCb6RYeyq84EjPzQXMLCh4LkvoJ7rmzzGCP84R
T58L9YCi8gkRpYvg+yUe3itf9L2Z/PcBBTmeQm85lVbSYTFDDQ6AKkgI9wX3vAlw0uYmA+VrYLnl
GzCBRpZ+DdgzJFmU4sO/eO2u1XeY7DQVntS/BXW5ecaG+ZWxJNL/jem3VwCUoaRCja85U+5nPaKL
hZqQR5ZE3nrCSZ15aeeNNuKJhBZnDv7vwegdKG3sIEDOXzcc7eIfq3hDZAqj1s4SjO01/Jnj6yo7
koQ3RJy/EgDYV/6r30XsBbRI+BHS1Vq+0q/IBh/JPI5YaMMCcEshVrHt3MpP4lLA4POKB9waT0vB
TcD7Nv+0WWhD6S9y7kdE9RaKTioSQ09BB005jNy9zaDmlKl57ncYXisVFTNAjYxAB9fLs5UqGJ1H
8Q7bL0zP+KQgprhM4n9mARj67Be4oMtHWLo4z0DZPGUMc+2uy1QDlYYG24lKb3IRyR4PxSDn3p70
6qaUsbE8x4fcnJ+ukTWo/l3Z7L3Z9lqyhE+An93mn3F/u3MJInZHby9kR55ig9ixdCvCAKvmB9NV
6Of64oFivw4Ic8oT70QxHiqmRwoDotib0eMdQXSOi1sboyfLOqr1BBUQu0IU+vFcyequaNftQBiw
qNL1fdupO3+EuEZ02FBlA1PdZtNihLV7zkxF0AyFtz7zMHIB2geo132qxr17tNo5Pq/AmZtwpHAc
ypxjzn7YkAuizTA1p1Lgc4XTfrR4HV6y8cRwEqQGPE4LGB8beAOyUBoh5NCiO/sQjsrczY5YGfMH
w4repSOy5a5u8zqDPBgHv1+OrOoEsoq8YfaaelDTUA9jDKmAiy2gn5m2Iad0CQOnuH7lyCO5ODSz
ozl3PNr0eDqw0lOwJfN88sJw6IKYIP/flKJBUF1KM1EJdQBmsUy9RUQw5YXhPvu9WHE8NKcoSG66
lmBrZEv758EfFnstzSB51ZuKc77mDQ1Dpq1pmIKksBKXhE9RRAI3jNQt2+3vlbageeYojbssduBY
wRlYQcenCZwOj0VgVqiDHzE6R/lUhmPcv6Uw5faBoPJITSSiyh+CIHmCU/Fa5eJJXmhzfryH4mRW
084ZCXafRAEaL6Q65DqUiK0nzyIB/5aVB3lXSSHk2IBKoWJBhTjCNYFLI/Ij/i5UdtGRq/9Icb2h
5ZuWYz0ZuSdv+SPS+CRjzeSTX+PDJiEcQfWI+L+8t87lIpTS4YjAWJoK2SGrQoVb50iZ2e69VW74
vGTfQjyBqNUHJDYFVkitnjtQEvcKcKOFhRtuev2++iuHBid2GVhHE9wfxhFfG47egldJ8J6dOhkK
MKCX0RrWHKiGkuPA1kgGvY8UDKBzBm+qz+FTd6Q96chXfHgkubHCvn2o+eFmLJHjdqhh3XEiU1O2
u42l+Ra6ENgjPKNX++QEd1par+dQc1oKQkCSBd51MAWQbhM7F37+ePvl11wHVD24r/f0UDXAFnPI
MwnmmLT3whrQsA5Wc2HZ/z5QEsYmQWSabmfl3YBO29jtxHN1gpgEZX0VDfop8/Auy52eHBed0rSz
btiHCSbW4gO+cGtVKZsnQ7Z1yFitnLZu/2v0pceBn+otfklfFU/2ZXz9YUtgyjBzSOP1BleW75CV
LphymihvloTZORxjEOTLF+9pjLhEp2kUtBJK35zZ4m5OZOdKcHMh4ryuFfESw1Ca/pXvgtLvO4yU
DlTCXryuIaAwsRd2+YTWL4HNlYR3stbGVDcDP770oNgRRnuPVQUM1i4pJwaiVsZ+R3EedLs6aLcg
2eTURhHqjHQ5W7JmYW0RHBY7ZQBpV4lGP/3fvSXD62rrH5mMXY7lBU+rSxaZX7xqqdOm3ZN8z8qw
AF1n0Vs75sYCNNG9SuV+SG8Twlq89VpLlX6kLvOsU3ABfQMRfWl8xo4U3m7zxua8VK+8VB6t4HjC
PfDKZnOIJX80wy4tWiIXSATOi3xovxxeRNoqpiDhzoRF4Rl0tJClcUJ69Qyy2dNmqhdIzYl2Kb0P
N03U5azzgcEWIfZdK5qaUinbugd90MXl3SkgCCY3c4dtn9r2gPa1ZAYlE8J3jjG8pjXJPUd/vFVb
m2TJm9AcfQXYEvY4m6GkoJ6q+MlVyH7BMUm9tRLgYR4yGtI+t6gNmZUrmn6r9Ilm+97fxDP3oGWu
wnbT0oFEAOPGGhhqJIcKTaVih2cmrP/IPyRI3n10QWCuV3J6byz5La77syI1f8/TAaHZyxSr+fJf
0gyaiahkpAG2r8Kj4/2fKZ+QcWPE3OwCdkTOcdMg0hfM9BT0HE1SCffMHNLb4Mpwin/r7hYf8NKr
APTMhWKZBnh9iJ+fHnm4bUhLVclMRcjIea2ZznlopDz9IS7BmJ9WxiHKuCXjORrFWhVV5ekMar/k
ADY4nBTyPBjQsQ4YrEzyNgogFC0t3JL6m5juvZaSwijjJp3c/cLSWb9sSQ+DU3WQPL12yeaOSu9C
I+dRMQB1MTf5fsv3/cI9XsCMEtSF5m1y8160KtfnIUobjRTJEllCILVmBszNWoVvp2tM8jvKzMWn
Tq3OujFHt34X2/QkWr0Dgwa1KFyMypocarb4WhCt2nJE4dmqtxecI691e11394+coRTw/7nJMNVk
6TJRahOZ4NbeRdpKhE+bzEHBELxRN5Gtf/PT21G9b83hOqPazLgNavBOUUHmiKVOxKho7jGlQ+Oa
obxQE2f8Ipv4iohZFk2saYgrqQc22Hph8dGZ1Av5zm1XoPRhcRlLxPmD9WeIKnkWKFO0wSHhWFlk
TgpZ0uZgB+r5ES8x3giMyWNCAPrvyBV4kU75TtcmYFRqj0/0yl6CVPN3U6IQtrJi6v6r6ukuC4Hk
hDyxgEeUKSgTnagGRprg7Xxi5p+5rhxX77G9WDsgQvDfIfA/0IYlPFhJUom1ZHwtMfeTRKpm9h7B
WyGymEZmjOqDa7NUYwion6RVaxfzR5EBTWvO/HzVTJDgORnu0AgRUghAxqIpXYHA2y4+N+3oI0Ep
jHuAuIE8K+lhiIaFlLGS273U2fX/W523aMEDsuayuBpjrQzxOwTJTP8uzD/BfDBRbmnulzctefYv
vG4c7OU7WpOvl+Ukmkrar2wXGWTn695Nps6RkCwRVuX6r8gmwCg6oju8la/OlXSELjQpzBM2EeIz
qYdfW00gnf8AURqYY/UtlGFbiLofC4OFrNcKP9eKMhZgXJGIOcO7OO6hPUyE+N6QfPPvm3ztDsj7
Nus/gbRhO4xPiYJOZ8NIamBkYyU8qVl2VXz5X5gyUC0xS8aFF4jeQI/XyfOSTkwrar+kdChVsrNF
CYruX7RNBaL7Ia8wHaNgJyZDMFTOKdzuyGGrGUxhmArRysccdx1Tslf/6E+TARozAk1CtPfT7Y4w
lShn8FeXPe2cAu1bDcEDsF4S2J7NEYMJL/TSzIXlkSkb3Z0qw6cQUj1Nz2QbIVpiNwn/qyqaZLgN
wxIX6M/c+RMevOImU9hK8k089iZl1jSscx1DEAGKKH9F3rAR/5g6gdvptTCh0LDELsD3Bs7hhpsP
kDN7VNzVZvTXGCQ3DXAWK7Q3yWZhnZqSQgtU0gW1dy/UZfQhBcwuuTkHD4tFRUCQewU9crFLCIiK
6FyZvR68h7oytbMEh+YDdkBWvz7NOzp/svJ2gItfPFcTHTCNMjHvj/F6Y8vznVjjGl0/v82AoHn7
ksB/rjw62zeSPSGtPLe2PwdLEKhIztAOhk8LF5DmapHovkUoX4my7ht/vJxxYkYEitWFqfEiglHV
qEzrbn8/mRNd+psNFvVBBsyO182KLZaLFA2ZYQmxU+fbaCw5Ea+hyRFjhKkQN265Ix2oiCU59nBL
ebJHZB44TM66BOpbmL/n3kVxqmLpeD1y/EPmbUvh21POt7kIvrHwjRpM4lOSvyvRrd6cekjAPNcn
5VFhAmH8oJAaFV4nsK3Kb1nY7F5xvC8VH48qe94CdMFDKPoKr6iWFOeu3aX8B0ZguumIVtbnKagd
Z+hTlYU4IrPts5STGJWWguil9M6EJlaPu/OqmmwJ2EYXCN8KyF+kcqRmu/GcQhBAjOMHaAK+7cJ+
e+fvhaceb7jEpyMeQ5ClIDp8Hi37Ev5cCvCAYSU/09SPgBECet9oMzaOGrTV1fvR06o+GqcCZHKz
R3jKttjVL68cmNhd3BR9Qza5UR1MRi4ZN5JMxSGy4E0EDM+3HEfZfFR74KBUC3bcx2IRIbV9nxLx
WxaxxPrFbGUC0dY0DayAlGm+ZsjA1Hs04Nwl90mnyT4Yls3nKmC4kHdCz8zrhkj8u/i0Xk8DDhpw
eJSYE2h+SsBDX0pHsPzREe+BtOrf8kV3NilbodJfQuE+3nzQK2AXn3HArQYvLIfMpnjgEmkN8JlK
YOtZe5OLuGIm8f3Mj9aX8IkmarXVwNP0FfWI8LmtcrQWD6BPem8APlwwNbq4voP7yaPTKYm5OlSP
p4uDq7dBeJzGSZynJ4ZUX8O6A1HVk1sDwKL5ceXRtV+3kSbb3vH7ljhYkLy0KGEnCuUchzA8nI/U
2Q5MSR5YKSexFrLgLjhWd1U6S9zPzH4OaPaTMh8GXrdrhgg7cRjYHZR3E40n3sHK++sFhBeO+qSN
mSdKzfZ5kVALbqJfQ3aOctylgu+7d6lOi/peGPtVue1yK2IY+dNengswViHxhqERQiUTkBLiOKUx
qEe0d+TLVNUI0SE1L5d4VJiRXry0EKb0UK7RtW2+hMZtILbNcF101aUEeAFDjrM3/9cGextE3v4b
3Fasn/TrmznU3ph/dyFa4jpYi0ROAeoiO7s5t1RCJL5d8UIseNLBwZDWzCXKzK28BCDztGBud6+3
2PVM2CVo0J0mqE75CrGC1teXECdSrsuk96V312YL/VPVH8YQnoRH8b5T37ZVogr7WIKQU/Sg2Sey
lPyhbX7n15strBT80bmmnoM7nZSr+odK2p5/pZEcm4k9aGzuVW9jsZ03Y7/0XOQdW+dYjTQrkmGc
5MlfunGeEHBJsIRs+wVDpXs/bIaZsJCJMrrstLgaOe0TQvSpovD38ys7nAafVh1wq5HIIt/Zf+Is
LqGtInTSul+8rC9H6SucbL3WI9EUMERLyExDIVMy8dmyCqYxY4En2+VxLe0creWQRYLTFZ3FYOnl
J7N9tEwmkcEPPciQSnsEDxD5RDnK/hfo/EOUA8CRI1xbzUptolH0lsY+RGxT2f+YG20NNQdd/ixI
wYySQ+oApvq7mCMvTBn1rRxosL8zQsB1YKqI5N/rgS2HJsvSI3X7ZI0l2fkrKEBsi0g77f1E9iRJ
AGnDKlwsXsrw/J/PfBDz9O6Q2niVNJ53dOeV1lwPnLKww0cjvUyEtHj/fkxyO3ff97hpdAr9RqU6
HgBDLvgN+VUHhqCuA73kHeUAHSdmUItIoULQsItJy1AbnIspXu6eVPyKOhPMVFgCk1i/NTbRDPDE
WkQHTREjOiWPsWYN61qRZQtDx14rHsCukaEx3IHTxKu5tgr9xJJoJQojQyOfF00YF3ponDaGC0bA
EGlIDdmhKuDuB2Pu0oveki5DQB7ICERf/2qjOBVi/H6kDyNYBaF2g0OnxvD2TxOGNplQ0p2BBZYj
wEofiWa0NSpaBz33VVHk7D3rD2Gt71PBQtkUIuiaBsYo7Rue109dLK6Ss6p1Kk9uS+VAQ7b7o95N
3G0CubhnH39SS3eWTUub+2sGAGZTTtAwA26l9NamSUS2xVr7T1dg/7t6RL4GoiiOzYfBT25MiSLV
luGG3XLJHpJyGhdao40+M+BhBQ8Yl9YguXc1ulXpfpjc2k3LAJZu1Lk7Dwk11MvcwP33MXyjZj11
FmDpFHXu0uhgNFDylRfZeyvMrAmGGgino21C7db50ozTc9J9QTnUlLEkAs9hc+Z2XkTkwiV09GKX
h0uzlWwm9Mbw1HnmBg4Yl8Wg4NS0Tsfjme5xAWorz6TAFXZZbL313MEufGY4F+CWsSNNVGXJSK+D
Xet6sGjrzbyoFuJ2b4VfyrHdP19knRG4djAv4NAxJymX1HHNO/2DbBkuHqzTUHAUDzEpZ4ynvuyk
5r9yx+3URZPHZrbE62Nu0vgEVFwRhwSyYcThIc1sxLJq8ZShNyvWvh1EpeqKRFpRN2h2jjT6DiHr
nj+7al3LzZigeeRPs4dmifuwXCEhmjuN2d1rSU1ub+qwPBSrN6FPmmTIdxF+1yFTjyGWcq0/WDXL
ES3rBmLp22qEgFS4MLrKtDzthht7ln3KfgqC83OY4//cK7Q8uYKDaSmvDAp1fih5Njn0hGPusJyE
5wO6o/ngLJ4y0BpPjckditSYoqFJmjECyhVM6jSkSB6XM1uBvm9jVT9oTSh3/NmvsStbfySGa+R8
yqziLaGCDZ+q4foyKhR/xvcJ65kCfE3DZBMHTNUQdUVjXl7+Jv1Hi1hMzb2xAbE9vnHDnw6SfjZE
KPyYqd2wWObG3OYA5tZLTJ2E3xZLkx5RNVtj6/EWNa+wT+jkd9ndVefAG7B7VvK3oEoz0JNDW95k
AvULf+KXQScREdXsaKlZDSxQQilSNUxCsXLOK3MmK/jzSIipdYWbfzEyNz7yNUX/ohZwkVa2dpkn
A1Gwgt6xvTUVxv5f+wP6z/gho7Z33BJTAgv+Ae09VuuZCceacPCMHSlnapeuGEDOAC7RRZgPZA3r
Ol4hfmpunlP+ZQeVldMlS5yFU0mTQJEdll6S2CPCUu25wv1s4+1UaujoLqlUu239l1XV1afV8Iem
Gttr40b15Jmrj8uNk8a1QR+IyOkBwmMtslyvXuvlPrRKmF182bNbfeMsvzI2R7wRrKSsvdxPcgkI
tbi/CHY+O63Cj4S+RFuAQr2vCRoZJOCgLZVnN/VnWY/LHqPwDWPjnhI6vvmTCLOMv9QS9SbwA3Qg
Bwps6fvlrlEqJKups1o5dD5VuYVlF2mohuTwHpSGr7q4Ieg18GXC1/KYwuQgUqY6tFAJGTBgP7Or
x4/oG72a2lAJLn6mcFczD/exXPVVRiFIEbMVOfiwNePhOdD/BMKOh4azqUgciaiGIjpX4mp5/Rc8
vy0jAUSs4RCTdRvnrO+9XpMiit+DmYAKq7A+hrfgeBhah4L35tiSA5ldZFgQkJwvS65x0LKCE7NL
jqZrmp0LThU9nsoKsOH+QuR38RxKLxW/a37P2NBFn1kFfEETzeZ3OFcdYEq+mAfdAB4hnWgG7SmJ
AeeYrDx0PndQG5fLL9ZGlGswbLNo1gYHEvTHpL3QK4FVGgDeAKVfPVksyiQfUz0R1LbWTJKr64xg
BZct+ZzfOK/GLDbTujT8tOYd7VCL/zysEqUV7kUScdShDaXSh94YN2MiZay9HGa1lYcP+BceHYR5
7/DBVq2GyGiQ04GP8jv2votMWSx5Mo0hLwakPYdrKp1DVxT5+zX9eDStgApgLGQl9VNVMPOlsKbr
VMvbdWqjX8SaDxbozlCHh+xw/ERTE2ca4C/W4deCKMvKbRIEvnXDBJPnJGEVX+NGvDAMS3oLpnRy
hCse4QT28WhOr5F2tUBgKFxZ9PMRymUedS5JHOl9fTDXxdeTkVFUzggWe7YK3XipQ5JMka5r6xx2
63bwEJ0uDEWiyAV2VeIspHT9iR2OxIJA4WwAh0xsONFDX4El2jUeijVHdK9/EAnY6fYWPwTMjdID
HD0fbk/r/kpSxnlDs2OFs8CalRFR55cCUQUsoQdwyR7kmKD969l6VuLe3IGqjWcQM6r0Mq4Bn178
a11W98kpkYHFE6ZyDXYzXWhjjEphbJ+y0XrVNAsBkTzx5Ol3lb5+2igCtvDwh6zveQsnJNZGli54
JHdv7KhtfvhZ7JQICn/Gb/yrB0TO0BSCfYCyQEum4yF3psibem4lyAJmu5M7L45bcSlf0iCy/kf3
S48tTxo+wrZYUkNypg15UaYXipBDfmxldfz5JRrkJJHiUXdEGOtPTqLisxmc23WWeRpML4zKdDUc
cAZvPzxEK5WOYkx3ThQgH+eorrMGYtHgU68bL+2zqWnUqtSv+wIgYv+Zv9ifKNuRus7PD++xFvBv
vocZyPuTUa4QQ9zOgN7ksnGrSkMQVGbEuvCoceflZkhAjA31jTDMEAe0Iqmq6v64/nzChoxGZwh7
KvgEoSqM/6XibHoVfcqeJle9CjO5OTI54ScA32DHWhqfHI4exvTnhrw2B9o5HoLe8zZDghl+/Bc/
N0i3OYOniE+06n4FL86JJQE+9nXw2cgLG+e2LEwlzk4YlS5j1Bz+VnX7Z0d0quWwXNbDYCiMB3wT
3+6MaU7weXfceSeaJgcxv+KlLt7Vz8HPIHUfJn5EW5aqQskf3D7366k69GppWJVtJOzQLo2ke8Iv
DKP03ASbtgHs7Jp9yj59WxviW/OExZU+7DJOUK651x9kQRlHSIQFlK0jTKQD0zQ/Wkcnov8DnK5P
+/vNb9QjPxQokLF28o27rDqrCc6Aqa20q0y0fWeNYBNiopNfN5qayb5i7h1E+FzBgGQTZQZkhsEV
CCyocYNnjv4RZNjKlk/GR5DCwBkzatE/PCpv4RY0NQcCuZpk4qdFiKMOJ3AhjudP4h+Zh5boCo8d
gGmCuVn9nTDoHq3xIxgkbc0UqGEFqLTQpIA9JxaAZSCRFAyZre0I5HxhLQ1BTtNpJqQlk4NAjrjC
BWJq8vQFqh4TRIgATZFbXDxReJEqfILapGWQKpeQIRp0AjFw4OsZr3LXonu8ArmKjuD9jtQ1c6Om
cpBuYzKkZAZw7S/hkJzyPZof/SvqWYtbMeTMessURAzT2pRv5L88nH0qLe1We63i2WwW7P4AV3Z0
ILH4Fkfn/LQvgSA/HEWZrDHJJ3TdfZq77tt2b2FtRdeaxfe9yQM6HUFgak1xlFFZiAZUvSilCFcT
D1jpO9P4kUX+r8zlt7nfAabDjlkK8cFOc+mCQodY4KIm4BmpG8XDA8rvAAO7aghrkZENZChPxE9J
e49Zvc2Qn1GRo6DOvRhkiGdu5SK4hatEGHbEtPot4RzWe/8xsOvqUwsde4VISQw1hqiq4OTsQO04
LpJ8+HrjvLnn5SZFbES0tllGyWokJMFGBAMdpYasBulnxtC2uIhGCryvQT/WziLK6c6+2vAsbaKj
qeHlrVo5DeIAvyTSRwbkSpctmqAjxwz0Nw4GNtQVVCpxvnGjTWftI7nsHOawyWGqm/6TsbP1vcTI
F0xz08dLppjA4yLOAOxq/fjNHc+I2sp2WAqBs1r7y0UgSLTxYdZJUdFbXx+vg7fKh49NzwCNHORF
ESPvyAoAwpWNjd+BIU4dK7ndmUIe/w9fW3Gu7iu4Ut6wvLSgkdWOoAFDSHJUF74tnwKxrYHe4ZZm
viGKUBBzYh5vZfZd8X0wasyEAVgOkh9wYy/pFfEs/XFdpXfxEKOw+OuKRP66NiyI0JoyV8XYmsX6
TRDptfTU1hurMIg/nj72r7PyZ6+PsMS9MpoCCXKchZ6caMQPDxO2yqsC11sRVFPK480k4ofZZ61W
zNo0Ylq4Z1v9jQ7DollYpo31V9BTI/2Fd7mghm+2YyoQu1WGG8n9sCyZ7jPad6zlM3c3RgobADpL
0X7PT4ewuDUVshBknZ1gY2ogicriFRpae9mVMB0MlqpolcY508ShMoM0X0OjNSdfNdMO3cyrWkx3
TD/EugHVyknVcbuQ/poSXFApYMCrn1kZ8Q9rCdH+N5LZhsxKn6sNIy8n3LD/JijEhxSeP6exzx5u
w9lAU8TlbAC/6hnuZZpATdlTM+DcvgRg2i3I1bms8AJc9CdrKLSj721n9MXJRSufuPFfFAL1Rcdm
h5YrLXIJFV/Ewx01bjjjXpqIdcAldX5bL95Vfi9h5aVUvJ2AxIssEFJVFD8LTtAT3Sd0N3jRZgqZ
eWLkvliBt7tOGubPp+7KXOKcevXgogBQsbU5/q108KFREqJZekOy9ZGvVxUi34xXNk8dlmvsPBI+
WQ4Hi7ybwd6GggAr6a1YhRckspdAYhsxaV8yOXfVAISjm92/ZFoseREM0HrMjbCfDNP/gqMX/1jH
OLdVJQCqMkafLwDeoXYo+60784B23DdZGXn430vl/j3qP17D1aP/g3svI22lAXzn0HzexvylcQjx
VJvC2tmU1kBMcVGfY4/c/wIXcAlc4LyMUNwTUJ6UxzXh+81UZgi9vjzmQIa6lZaWVT2GwbPm82G7
o0zncCfAG/P3l8oBA4Yg1dE/AzAd43YOmzBHHqENlEuL/DopurF4f8cvFcGRjc24q4ePiyAbv3+b
SfdujU9fEUSDEY+wqMenbGPDBzpEN22SASS4bEOqK/lDLZfACK/EvblNvd0pCzkJxy4r74vF4IvA
MOeq+yKa+FPW3I1aD21kDTVnXcojDQkNc3TGiSD1VuiI+8dmeMK+gftgpT3rHfDXHMu08fC0EKwM
fWMVEKP6vmZYNGP0GCYWsn2uEQmddoQwxc52ndef6vguTpjiFZiqprVxup6eTJfTm6+9Z9vEM4yX
QS8ruocqBsxp9H8wYZ7OPe76Qz1YrDrIEuRt7DozJKv92/Mti+Rr5ml4XfvGfM0mkVT/+Mi0yviX
lfEygfwEtslAZSiTNLEQjZV1I2KysBAnhtuAPb2I8CD3jrkXQfgKpw9ceGjB5zCJRyqXiCL/fdsJ
5NMobw4Z9AE4kH19ABWPzRsGi83aj3KADRNtw8DI4lDqvhk8vcs7yIIAPMVWQ7GLOD/aoT7zqoqb
IyUV6Sfxk0IMZ+22wbS0z2H2ZGKxpwFg4ISoVghLI5nAuo3YaFGOX6HYHJo5r4NVOkhd3GJxNIe4
gTBK3jr+/9FlPqbr6lIPo3MvcpAg7H2mvbe9nAMWkaeB939PRMBh+pZI4qB9WPWoHx3edKBbyIvN
b/cr/3F+B3+6YUuMhnebxO1SqafELDBm5acCBbIfQ77iHxo9o8MrPyOqD/d5Nqn5511mACMDM3Wc
xKxTXnnY3F9+yHH5SK6EeJV/esB/gguRP6opnQ9ko34JPr9B5pquS4ZqWssRejQnLLHoiAhBhfrA
ebYpmoIsKpUhbmzAche4sTv4sQk1jjXQ5i7BsENT7v6v0K3DbCsQEjODK/5PHTsNGrmljPcU9JdL
zSCfq7u361yjUDd6HV65fj/QmK5rwldha02q68UKof/xIxTY0u/li3/KOHpCXw6LEOGFUGcuLYne
ekQyJHMoGJfnzjHTKrW/7PUPQxgEYr5J52uoXGJWFfSC+lJy2suvwkJh7N6Br691BOiHf6JUpDVS
rzDSD2XN8Nx3RUKKt5mIbngxs+NuCcQKC/6irByMgrmvK0QWGm/I/zoC0oXDC6Z7P5C7jqjbS0xz
82HuEaU2eGvh79jTvPrlh5CycxcwDX19VLzrGNteEpAfVUvy7SDL03gk1A5Nc/8DoEKKT5KjomKi
TPDlNyVI6SwPVwjwTVnLSLWgQ448PQXWRkie+pHJ8paSIVgRRjs+bkeryUP4cgky+3oTprNd0TP2
DlzmJ9smL4YNfS7ezPe32E51TI/w2qPgrA4lNH/KpZLREEp7+a+z0o+vqxVV1GF0yB4nP3zJiHNU
0AKO1vEFw9FXfPSvsqEA2mwApkw8lDFdXxrJxhlWzt1uG3XrymoaCxg+bfOEoID0evEKj+wLuCGh
EjQ/TJ+NtUKewRXZwcNB1QmSpqz+oN3jq8Br/tc/UqksilMYT94OTnKsI6zYLMHNqTS5TzSwxUTH
FCqzh8R6o1/sI75dn06mp/b7oDMGlt2muAQXHjlbe4BfmfLGFsltjtXdBcIEjmUPG7mHO/ywExso
l7mJkYCcUXPk0opD/QvppJ9RUN33LqR/JtAP61/VF6AsHzav7VulSqR39sI7GyHSCVHzoBduibAs
x+k38ZJMFoZl2E+t957lRsqoj9m12D1I7a5f/bZJYz+0gt9bWAoBJv6PZdDNDbjezylELLhJiLLL
Q/ZDjC43g6E4JKaVI9c+OGo89NM0k4O/Er9VD2Yyh06KyOEnMW/AHAkB3n47+h2g9qBOgsZcglCp
vRinSktsK2kKlXuuioITEuVvsqkoQN+WcbMCdnEd0K66HLPdBeoo/+O++79AT7emOxNGeE0xTdkL
oACN4V2i1gUUJbQV1OF9iB7G896xYfEKTw73ceYHvI1blVvQ2gN4tDmDmyUI+faTK0Q+Pql+YEni
2V1fqdLfVmXAp+vSRnoVHCcwUcN3Zbqo3IbLjIUMs2Qtve8HLY6CEHK2hKza9i3bpyphD8wVovJ5
n9ZDBlzG7CFaWO4iu8Eb/EtamZz/RcyftxIVABiifE8DhYqXJV8I7YA8EaAy81OWp81vzp+PNV2d
dTKIvSFP6ASJET7MhGCqwCad05NL4VzpERJgRReJzOYJeTLGs74oOuDJgbFngNz60KQW3nR7JX1O
gokmicS3qTOroxkby8z0X21j1y0fAp7T0vPRtNqsoVUlVIciYMP+rADBPzcQpsEqJpfZrF39YPUI
5U3mPq5YpVhNUEovM40aM8ESImLZbzIFVbpCGsFh6w182AGZsSznW4rK9yvSUUvYfOD/9z4JgFOr
xiiwOf9HvQgCIYKyN3JHbSNfq9NOxIPffHq2s45Uaqf0NaBsUGNsH/pcwfnkVqGF9hOdkfI7LzUg
JoqIjJmXps1XKukjtGoHDxBWH4V2ljW14KYwIIB2iZLihoNslWXvCXAPmH86plQJbVx03S0Eay73
vWT/Vy3V3xZDeCkDydQp9xafiDvnxQXQjiZlfMAbmUDn8L1ldmAUhYs/iqt44zS2sNfp4JBBBGYl
TjVfqBxdLy632BLmJbd60sOKIU/NMybrwBLiWn6GzWswaRcg/y8FwoKpM1dehAJsb4uviCT3yQJj
GrvEmFp1zNMbtS9LEWFjTdjeautGZ0T5PXTfxAFXrsGyxUhQaBZWL0XeE4yRBd7YEnQm+UiC1dCN
/p9wGTJ91z/DyCRIfH2/yJvW/mbjjSTd+riYlRjoAiOII1Er5rKp+JrRupgBFWtffQ2RWTh5q8X5
Lkb9nVVu2ccJmBVSm4Be48B19JyKrVq8ZgMogC1ENM6/Fj2Zy7898aF7hwVggO3f3B6Wo9T6fEiZ
jD+73Sa4QFtLLEDED0ZRlcfY1BPCOwvCDYeoEtegyItxcow/JVpTUKJFME7s+P62Z5soSLk7l65u
cr7GLEur2XLWxOtVQvfA33hhAftgpN6O9vqJFA3VuiBMMbIyeAFd28ECA+NDVolhJZVp6NujV5o0
FTEh/mfUX2iQaf9/sg0PeUaXFyBqIp9aaCJa5wjtT9FRMLhJZczov8I/wda1Cb61CqVUScA9/9TW
DTgsdaT/q5qUCEuUnSHaxfVqMyPNYvKxYcavkhJ+g/sd/mQLeiewTdX/PZIQdOmb4SNF9k7HqcQB
IjNAM9L+R3Z4YQMkog0bC/+7bGBmt0h3wy9iv9WWvH+ZMaX0JGx2oHuICSJSEwaW8+aVerKWP538
1MPzP7wvw3Aq0mLwalhggdFRfW1eoK8LhqJk0qv7KexkTWLn1SLxsInOPJHis1HaJ4sIFCj2wus5
puNKEJ6PdKkPQoYYTSSBjTcnXLWqE9QwYioJuYczQBsEMTiGjJPf7LpNBaB360D9VAF7uBWQ9l36
RHUbrsVG+QFfWMFqeR2p/8x2Qb/a0ZjcuUwwQvAZk9B4wqIMxNSwKoEwCqKYv14oYVm4GswM/EkU
SxMoGZYOZP//Ot+G6O3NdZGxcWIsTvmm7GmevvSm4ULesxEBGgEogIN6lA136buLQ+PKpsp3Qwz1
sH/3oDd9bf/730P9qncZ8yfQDiUHRloOKbomEIjeOQlnZCN2TqACU6xYdjmxE+y7EN1PtqQbJM9v
Mb8DS6jb4TkC1eZtVItLUSl0A6QQ8BQW+v39eLBOv1GjDkSuVsBX4PYaYQ+kyW64FPfrbie0w5H9
7PISXqBsKdhzerr/8iukMrx9eqtxPpKb83lCJ1cpFdmkjAwpXiJ90YxT5Th/vWlLG2MYh+morJID
RKdMWkPN8L1hogTa+eaAGNKfu0mGB45dFLW3k658gPqGXyhZ0lXQMlc0MHKNLODUqaNS1LM6mBBr
SqCpKKx1lS9MvDAbmLoJcQyNYY1EOq5QDeaoZ+j99UyRau/OYXVZ1G1UayyQmHliyo3IpEicvCYY
i+DHKtyDb8w9rHBSpfg1EjcNkJm3q9s28cUw2XjUjE322D4N5A9TKVjo//FbbHZvrG/dI5C18bqJ
9vralDr5hFQ5UQvB8qJpg8Yywt3mNWTw6A7j2jskIXWlPUMd/grrizkAsI3pEsjGNUWJKZihHJ7R
xIZvoDapfzEx/GvJUFGwvqEHUviU/6VHqya7H/ranSQCT7DTvv5PlkrvtUyadSnwfWQ9nBIrqy/6
fo230OqOYbK3CYjK+7K+WeNR4lzaQy231twQAEEXS7Ma8M5qntoybufnHwYFs2VGqXTIx3qcao09
vefwD71RWMLFm01JamJaw62MBq5WQin4u4IBpZwQMR7KLhu1JbJmvObO7N+fNg/Xp+dPNSqeTmMZ
q9QmvczlpY0HsXOmNb4d06kM5PBIC6y1gP/Dh2iKPSM9J6xUXqT4Vr+Ej67E8fOQwYnmaXBdVW4C
ci7aKs6DB3DU/wRB9GVJotCTHPXC6oevfoy6pwlfWyIb09m00jphkdNB5j71bqbmMvAC8Nz0/W4B
3mhzsupNLSyHoqPDZ3eTC89UQf1zM07PZon1kJMi/ZHsgkS6oaosVBuXCTKnQnV6rn8udH9vRXMR
3tFeDeBQYAERHc6Z7/XWmvgO/ErHFHJWMbDlSqtrWOGDDHgeLQm5ZJA+cFLanoHLeHojWarSS6JB
KygCjqKx+u+s1fWijd2tmgTLDFq3GKbp+zMMh7/w0ecQhmX12nHFKb3Q2SqICD/FHuluV+g4bzSj
pOnnuifLqiYu/p1DOBt5uJ4MpvK+6SsCgiZt2nt53OmhIwEiEnlcAh0Mewdd2TwV+n+4nk9Tj5i9
9RsI61eiN8mGptFYcs3e9kNUwU0mjxJedxfVX5iK95Z2jThVOakND4gGFQNS1aRmR0/R7F+gmSW+
i94hr5+CUMMUW3lMCKM3Udm8RFRF5AxpKgyfbmmoYL8FPlX2xrsxqR3MQSOVcV8WGYrx83BgMsqg
CKcm2ZjU2oMQAcWFoeBwqrr2gUZJsCov/iNO/jddusKXymStidMOKRbPF9xYC/l20rE9CMJGhjO+
yF+3jwcFpLt7c0TjAiZEchu+yiOf+kj21QVKjD6pyJQ/un14yogjt87lX85m6jnJ9/vBzjysbBl9
EN21qYYprXqihbf8zIDJkulxOOttNC/+hDttyMfaAqr9hV3rS0D5/H5IV9rmswnOETDhE3qkT+Pr
TeJXdpA1vzdmC5mXVaeVFVq7ZAyCuW/RdkO6MTdOb9gP4RnlyFj+T+HGgWx+3vRWaexWIpChiyI1
lTC4BD51JVPiVyxTN2n5G0Ibp2EKrT5qByf3NlL+Z4hFYNoUTM7cq3gGyDYVe2RYlV2hQtcH3b0i
QktlsQPgcU6TngRootSYgMFQ5mv2CcFB7QNm/lZxHoLWs4PX3AKzKzXIKt8fFIQ6WNyCufN1wa5/
/8o6hVMJiANzmO47n62Z0S7wCkVPy/8lMhPrLZckrjtK1oKSzoEFhUUDk+/jD9lB9t5iSEZoinXy
Q0owDN/ITC2EOp4XW8S/CAcNo5g1mPGoYNubqAICOztL7uIwGozY8BwkjXgpE44OUFhzZ3GOxV4X
4hBzHT2L0m9UmhD46nBX5OlYgGKRCuvnQEvgFwoK1sfshMe/y44iwlE8wrmvNGlcpDax1M1dSQDw
FDZADcSDLSZKAub3O8je9w/eCeHvkYO2uQPX31HTuAuNG3/B9nIViZoPCEDtUjBkSxPhJ2lE9VNE
2Pn7SePSPNd+2HKPV/FdJpBAJPgc+cLUYgWKWi3vcD8KY6W+XwQnti4tQrbM21IerIX+6v0geK0Y
ALEhdvBH++/yEWk8bJUYy8ALaWLKH6gOQXkJODU+dpheV+XBjnXPFn4udxQZGYVHuclDqZdo4GqM
n51G0ylVkTJtLVjJ5lWPHAaxvHX4J0SzNgeBqobph8essdCxkO3aBV/tnR2LJjyw5dHC0abxZGLj
7kiRw6Xlkv4igUPbZn8AMH9DUwyokO/7DKkJNu6A4P2mLd/sUwsqlhW/aQnRKegXan4Sln+pc3W8
Zfn0FO8c0q3OI9BVILmthO/seS2l1uQFmcXiuSdRee2qzkp8qU5AvD5ywXTSE0DMw5NG2JgWaC4c
6GQoA8FQN0lIbCascnASKVPq+0c0243SZ6JrPHxsjcNgPALfQ5mFk36c/LPl/p147soFcj85KnNN
oV5toghkcsvJ62jKgc1vXupJ1XC2UkfEg8UMqERYODiT6cXllAbfeWPQ5iMG+QCF8GKdatFyDP35
Ipra0HIjqJZ3pVuJmTKbMIRrCqKTHzAx05S4Q7uKL7xqzCM5LXUu0OZWcnezQSxWeqHckRZquE36
wsTwbJcIPTHKfmt70QqRLk7utt3T8d0V1ZLvbuxfSNn4lj0bnfMCUgNEHqd3bzcsTL2zhTMTKrtU
G0HrntpO0wNj0/EFBfDCFkhFTnpry5ijMADkR7w+2kwxCnUCtFhOsZQDnHlEA37A0NY3mHhRX1lb
DZNHtNLw7aG9qzWKCsE8DNW+3qxTuafh4Q8YElH/UM8Oh3Xo7yiig7LOQCx4PtWY2BePRHhhv/rQ
XHZkUtkgsFMsR7AJ3hahCsflnYx4W7sFOWi0fkKarsWHRYZioFDcWqMjt088Rtk2HNLm8YcpI4pv
k9vwx+Qf2jczqWeHXmQVy2vLoKdNEO8RUdY4D6CSfMG0OHv1Lc6hu8ReV+CZA63nO74IAbhwqws7
D23BnwvNxA/PSz4uP+ZUq6xJhiaMRUrjw+fRmYzhdklT7PwGAGnylyFZ5aba9kSMObX7efHm79Vn
n3Gdnz4pH77Dweb/NNnDhMr6GPdEVoNmrT4rjHJbxn00ee1PqxI85RM4R0G1GQojDA01ldbBvUS1
aMsdk158O1MBtc8qFsiZ9iB149go7NUr3ORxx7hO2e72OireEnOjSsceQwmPiUDls10L3xyIXRcY
2oc0nuBKcLfUcvuDvEnMFMUj+Wq2BqmwKwhuFiUv0rlhHHaFCJ9bOQig5dYulQVPULZ16Z6CE9DA
hvHm+G8TbjFc38D2ufIlQp8wVqruffYbGmeAShYTXMX/USN7VQkGec8tbWJM+n28ejVbGZxeVy1o
vzSwb06zw2yFvAcRLuh9KsP3nxT3UX9gOJVfiSoAkZn3kEh3ZTmZgEHC5CAICyiw2+5XJahrj1mC
EvCyZExVrpmoCJRiJaM7hKgezoM2G2O7qfnZX9RAx9KDmGqlLglgwfoWvpfJWVnC5Xmeq1An7lKs
3ZtKm64r9cAbcgXou+gkxErJQLMg+6QvXPouS+09Ne1+gVY0ljRA4oGFHZrafH0gSAsCCEq4aIT/
wlqA5rjKZ9HG9UAjJIMbe1hpI8pHXhkOneQlN+bAmQqDTbzJok/Bnpj0Iu7qFPdUNASftlxuHidC
hP8VBaLwKjNBrbzVVGn/KDb05WUC/t/v7ravTDwGWa50W0H+F2PsIBz+iBrAIICWdRP2IVWHrCo2
IpqG9BKJZHtZeajKF8YUqTBLdA6o80JnyUQ3NAZfrhICiQRdFp0gXCc818hpZfnXa9ZQ9B4Nprj9
Wl7RB32vvjNODxuHOvGmQa+Y8gugTsOmG52g33JCmXx1Q1elKwB8FDiTz2qdHadrJxfa6sP9Gmof
tLYEGfdgkvb9xsfq7pWYGIE+d+VPFz3xlz365PeUcbD5sA2IZz7W75Iq3/p/5vgqJHJh5PYcmXAu
CESPmCyMPYVgObb9disJCWcZWKYNYdR0a5QSYH191BmNlzpRSNgwHqgq5tJD0VAK5VfZH483eZcH
Yuepb9c5uPRN4Hfxoh0PRz/ZfLcVqE1lcjO325/UBJvfrOLr6SB8fHVjf55CbqEDl7jVJQcxYH43
XDMlPvtiujIPTUIHtwZMInBCIlxW8a+VnaAJe56qmzjv99+9Lba/ReTdbGKWD1f5+n69fkPqfc9I
E4qcbypvbktjqqYmMiHuw/c8ymYSjllTU8tvsAx5eaTHAejkWeaZEtnufK1gm2sjdYYRTyg4mMwP
sP/Yu1gwaLFz12q9oxS8cZtrzA4ps9uof2aRXpPp6c6Got1L82rTl5kTG0Kzjte7z4+IC6N9bkJO
XeWMW6OnFEsZr19KdhLLkSatOwCMNPtk9MFQ1BnpYb/3sQ1EQovpmpvlmRDnRbR6yKchffJo+gf/
IkHnzsI5SYCjys0Rz6nUUg8dmhLl/6qslw/2ad5LiKOiRsxmcoHSWYZG/DeJzl5SzrfEH4cjhrAG
Uu1Rr8OMewTZ/hG3QKjojkej9akPNoD2O6eGm4vshKS45oKcEhzXf4bmeA5BJSL/FVi6D0GjmzuY
VzYlSSbDcaIjLBnP4qLqpGV/VrhsE/icPdWVpkiE4/JLaJ9h/HyjyYOUDrhQnOmdLk4I0NPnJ1zr
w8woxBvstgpMPf49l3EDQyxRdNo0YLMHhRLn731BSAHLDE1XYk8LIvuIWwWW3FHescQiOs9x8CE/
W9vVlO/Iyk69eA7Zm8aGJi/g4jVA4yWQ78UOii2CH7Vs8O6Bnj62kCujZaFQdR+/a26kuUCysU8K
vtLBUqNXvZ7hKw/Pusw87sbLHSdzLr4QSTEMIvdQascU0WQdDwopsY5N2oDg/NnqsB8OECDw61gD
6+eOGbC7xPFpqGfun8xk2jGut+6FBo48c85hfBE68HP1RIyuhEX9uLEiY8/60Iq4JZrv1MTs2zXs
N4kVPYZx8YbIJ7WSVwvUwOn3ZlWR4ywYVpd0SJUkZZlp5g8hUYsCNEnSPh4hGEB6yV2UaDO4om5j
KW5WPfYXDtt/RCaMzkFKY4UJ6t4RIXBMEjWBFgH5TNqI+GspNIA/r8F5VNM8kQGrbr1EsM6KTI8u
ehhnRWKvzKNIBZaSKquIkK6v1CbUKXuWQvxogm7+4KU/Wli5psdKQ4LmAC8su5p/AkAmLad676J+
TkOS/fK8Y0/URdervTL98ExefYdlps4fJ5DYy3m+aeYBFvPrMTh3erlrJGJL70XoAKfIWdREA7u5
jqTIIVAyA1RWvWOFlBe72V+SbCRrCEppxy+a8MVcz6Cyd/gnKb6GyFG1V5AcJ3NzsxHMR60NdaZS
iBpopjZ6ICSCzX13IhI+sWihTABcgQJgywB8cY5TxG6Ox0/Wz6g8K4hWK4WzD/Sp6whqEmWz+Zy8
54PgcyigizYlTTOJtQdZ6b+ZS2NbLe6JZqwRryCRcT0L6fIwm+qzZngCFp+XJyewNua9WHLkuFrd
4YPMXi9XZbrQggjBKCd5Ec+DJvgwOAQnlTnsqEqD64IwoV/KAzByP/d3NyNKbF8lD56isWenuf/C
1rw8FHkn2R/CUFtuqG+eYfmQkoGA3v36cgNA8644TtyYTGGNsmlKtUid+TF93U5zWSsGGV4JX8ez
b7a7+rVA36fC/J95C4ofO7/jH4IPQhsiIhAyVGZGIUdxWyiVhVGdaoRs3ucQ57yfhtShOBkimfoT
f/zEFQUpFBWMzM/xSEW3jiR/1rxXKHkOdQOVXjtB7sdMDHesZVN2sp0+89CslFvzqXcJ5RTz5Wj5
+6gDvducGVBfQZeLoVgc6nPyYzTFItpB3bsiYXLkvQ8bkDOsyLF4A89KAfNqkdOsFcsfThqaG9KJ
WzjCYVQ7nIXCmakwtCrwwHtJIBPA2X7XrFAvbAaq8lydk9GwGbvroFhcZdpuu/LGF8gNhKynHTL4
EZDqOl4Q1aw4m2f5gvm2qdDJfXfBVIHdzsGEmB/5d8Ysnil3gfItEpUYxYNboXsnmPRjFW2oqiK8
WTSZ3ULmh1oz09CQQ6Jy5o+uNOG13zvrEPMAr4Yi+/fEoZr1XqbHSYArc0TbDHjmf6AxdgMeP2ac
vc7Eu+oNjkN28VF1ntcTJsc9u6pZMLFH9oXrsG+r61ku8upvonTURzz9Paxs7Xy2lFxTiEy5Cl4m
moUKwMa9rqk6PSYFCU6vZaK97yYb6bHw2TJK5R20RqJw3xBwJwpmRfAoK+Eh0GJTraiuaaEOs+40
BvpgH/2C7yKLPAW4SVDCoW76LlrzU/BulMwDlhFiLhM+wywOVaID0crJicM4MDP0Tv/sgSc/RHBM
903lzYYdTyWv/RHo8nbGbdOjcjxFmewuWn/1VVPBxZwuKvi2CwmionpNxhBQ9ikTwwTJlaO1rfpZ
5fxW6g+uGtpilrDA659/1Eto6Koo1kFxq+AQagq642sepWjslp6lX2dHiSiomGeOiX3nOuR8A7Oq
O9iUdIWAmTCRrtzPT7SaXTIaE9oTRQypYrKjg5uG6fEv8YCSLTQWupVDvH0yT/YUwNZo5RgWxdhS
xaFgcUD+C81DYBI9QBUikVRA7/fes73wSBYwtJ93RySsp3sQ3fSa3syvjO6vLnnxtnVQjeCMIH8u
wx42+V756xNav16g9yTkNh6WRs8elEY/z1vlKyO0t//yeCHWAC1/6kl8uztYMAGCYDlRFZMJT09m
jy4IFuXd9rSGGinwS7FBtt/Kr4T56MHsiK81FwmTEEE/CWXxqsaeCpun3iPFpJQPKzlGb9O/tOnq
z8lIwOE5qMaZw2rQxLVkQ8UXCMMtfz1K1TTbUg/smFTfDPtAh0dhyA2WBc5VUOwc9RhG8FZ2jOkx
e7jp/lqUV3dyoc1qwyG0NpXQmeIs36KFZ3zrBwpIUGu+jC3gRbcuRGhjmag117PjUhgPLRKa9FhV
Y2KH5GuUQN9kRcOyc9XMCtPytcfMsegATwrLSJ8mBP2LYtMFUCbgZNwI6fMCt80XElc0IjxlFX5Z
CHRfBTwXOUnTPAxbs98exsTmRmOABlyu8RFAG6o/ZA9jfUUy+4k9xafKI7mGniZzEXA1Uk7QLUkE
cyCbv6CjJF7SeQ+ZZmwoZzpwdVp6I3ROeUvYSd/MbeGQYqnNhpB21TGQ7FiOQCzANwQuU1Gr9Cm6
9YSomdVWYs9gETkc4/saYlZYX7jaBQJZkfcDSkk45RpfaO9AE4zSVttTBGkUQbdOJoIm3bAF6U9u
6L03J4tyHkMmDeQEMthgG0N9qa9wmIpb+029QEO0WyILEQdENMpiHVNUf2PIeFhluIv8cwH7H53L
ie3r7wIL4HoI9lPaDP+8/px7cHiia0/Lvev2AQ1KXXGTi0r38CoJ1/EV1c3G8nGdEfGcMRfMmhj+
IH0Gmee5D+sm+mXkEpK5BUMKsNNETyBBJIQV/mEXFLF82p57HKYvVUiPY3gaGS6esZRyysTI0BwN
5uw/745l/ZU3Ss0vBLnzI7ZtGX9gJRDYI+0nY+IyXPtVT558Jl/XUA4JejP+nR9YYXAtrXgesYwT
kPKf/zANpQQ3pZG4ch+WMuMCGO5CjB1P3XIq+86z+db/3GzrMyCCsIJkeh7dAqvEgNQB65lOhdVo
SKLV+mIAvmU1Xesf/UMe+FdbJ5vPX3X1oyv3cTH2St6NEbTthRV70OEPtwZmY7BqctMa2k8JEe6i
UOeXC/L2RO2GvmXtB21ihicOAiKzYSXrwaowhmSxpLG0G56PDkr9Fw56aJsKhhvgNPAOi+9mAKSQ
hb5OpFXnC9nv3Psy/fVYTW0MxEzsq24kugBuaP1E9cflkGmsOzAW5famo5NNwBSJCBFVDw853G28
rNl5esgU9591fSvJHJ/Gdkv6r6ufFy7SajaW5fW1SN2TjQf8gD+cjKy0KppgeKFEjTnM3lpylSfm
pH/Lf/wEYunUTSbr5eZt8402Fn8tmYVhE3kGkGJCxLL8GnU92g6kxvI57oW3A0zp32J3NYQIlTvK
2xT//GGZKA8QESFTKqDfa0I8oOiIwv8hoU1v0NB9wtO38d8DXfwuqOQM5c/FeZODSrHbJnYN2XtX
Ibr20LuzVgWXCS8YkVn+PpZjYUuDjV1fdxlT5VKmc1EShNVyPMeKtmjQ3yHXZLLh5L/qTsbJZaZm
UX3Wy2nYlA0ylDNaDBy6jbKPBmIJH78U93D8FnjmKhvs9wzPiAjNBaodWAwGscS35ThylWtncakL
YLqt4U+f+H1FaOZZ2KMXs0gk6Xo6USf/LqVi9/eZg8ewdqfeujCbnnd13z5IKkfyi5cSBptV/A4x
0v43IyS6PnieIIPGxzAmQG+R2FJ778pC1xVZkhapvSnvfvV4gvpzaSBQFHcYJ0iV18fOier9coXA
ljP+cvqzPaNcr4TI4RDgLwoEwoxjNGE6Qf7GX0LcvAJSQB7iMQz3phjopqpuKSu8uH9MLBS5JA0y
gWLCZjcQ7xmp3OSGIKS1CAi+pGIWZA3c0fxmyh7/C7/tYccXFceIkJh1y2X8JLlTCfERQhvp/S4M
zWf1fWUFtKkJ9WLK9XE1tcgBJqaLE1ldrm5awjLpIzu+BbXnRlHMRz3PjgPd5wNVXTo60qwhb3TG
aOK7f7mVoHFYWGMt1WRG2r8myGs4dfB23m/52fN56Ynzot3uK1d/1E5UfiWHI6TNLW125cinha/X
MYlhz9irmShQOQ8uDMYXwdo17jHX+tvksZqA87mPdJAUyUrZVsoErronfYEmERy7uEooa+DNrdcf
JrJsZeE4WtDCQ9CdO0JJdTVhd6ZETgDvkyU0GYiOob7uqqj31BZqIyAPu/elHm/RpEY0Cz00KbcV
JJUj1WMWvi+TYpvjQkXIB2FrQg0HtMt/aRY5CpbeiqROTUvVS111HwEaH/lIetYCidDc43ZcSydZ
2vv17xJ0ShsT7XPipRUYcXHMz2hSLncr1HiQSO5MC5UXUBQ5sFBb9Onv23SbSmqxiEQz5+m/xBnb
6qOtO68VtzyIT2ddE4Vbo2/wwV+KkUs8EmndYBmY/w6FOATlSy+j1QXzAY0V86Qz7PZ4UvsCmpkN
/kRkizVT5KRhYbFO1USKCvm7vulxesogG7iZ+wKNnUhZacSNlbGtca98L9NMDBLVVMsdmH+WrYir
YAP0zwJeX7t8pDNQ685JjXdB3XBAJedcCZF0S8aSQ/QgQmAsUUYMsrBZO296T6RvwzpcgvH4LFxZ
bXZtz4o8KyZCwVXGO2THicCPONmnDFIjoYNiwpyZm9IIQPhGw7YD2edjLYKTbz/Xmdr7cTHjwCfF
6p7vKCjFi0/5ToXAn0aX9GqhsiQ2qeax43ei/TRcUe3kmhYjfQgnX9eqT7wOnrPJiX+aNxodJai0
dCIlpLBqJ0YgAP9dh4pmeKyIf8J7fNpc3u60ki61eRdhsU/lEGRA5llnQKDsrvJCDMyQqN+K4J8z
VtWzeTtSKnpXJTIC80NUMm/Ja9cPaji6BAEMbtUxuksWTFzSoTZOyRk7T6v31963982yV+926UZ3
Zu0wVq3LIfvHn/1WiDT84QyWkrRDV31EeWeImGSPeVW99vPe0CnPNEPlqlAP6uzTbwF2XICc7kLI
a3C6gI4igITq+MCn7xOJK0rV4VaLwcaYdxZfCOZ/uYKBHv22u6fyqzJDlEzkgfvVndQY2pSsFx2M
8Echq94xQTHRaAUfDzteDj/FtsWxGftDVdewYNDxWcSMIfnZc9EDvGBE8lj8DIuchDnzrZ4RhB7O
JIIMF+T/rteIvTiUh2s0QZiVIFGljPJSuQBLfb8y0+XYOHU+U9O9W9f+6ANpRXdykpTy6c+cZ1I6
3jrH70Ez8SohKN94CECp/koXkxGogo60iM8P1yWxojVpE9kwNtaE+iUNMeQzozBjHfq0nRKLTBaN
U/MAaxGRgMO3ohyfc3qUyLN7xr+4yqgUXl3lpNf7jVPixbqkobBPw82Ntw9lAC0x6gneNvO7L35X
sSMX7RYyHdPTpGehY3/KZnqVMp2UYAerMUBjGFdbQNGIjBFVF5qt8QQS4lmzLhm5UVDyjOhlM9zp
ruj/nEHzKTnmMIZfZ3AZArPxdNXKvYDBGje5XqAMGwzpElzT/czLUgc5U1WoDISMMeCuUoz9CIoD
+LXNA7mHkoyACFFyFY9GIAxG+0+if8/uDrwBobhjgPjajQHfsUolphgBHMj9l6TNRCVM2xkXBYQo
+CVVtxAaF1Pl8okC+FgTPu1gRbjQWLJ5+8x8DIv8QEYw8//iep2rqMf2dXcdg//cQurppvbRwnlv
49aTZyq4twKoee9lNEiQvIwpPzhkOanyh0iWCpAg0lJgsxQzmks9ooBfkpoRfSgNEnKBbWZhB/5Z
kgepH1kLaiILiqfnYur7+stlJaevFQObOtKgKjOH/ksHSjOJmXxC/yb+Xm0HqLdxErR7KAJt+Je4
ov8j0TYYpjjZJ8WSOmQ5VFr4hmHQtPyte7+tt4QdEBFfcnC/OaaxtWCjNKY2/1fvZjTdvp/10PmV
xB7RPUdyeqwuE5xm8jcyATP2rjcnhfDKRkEPmu0C9UiPUzoFYY8q4TW70ygOYPgAtc4/hjM01C53
0Xw7LJSqchX04Xmf/W2l8K1UNyMHZJ1xoSB41fP9/ZOeMfsG1tF+R8hAFRKLtovVKsoylAc53583
zWhHceF3EyEXVY3YATkRt/Odf57/7gPIDLL8JL1Mt6ksLHsIu0DEWQ0N964ZSIPpugaevRFSuf+S
Y9fXBDBmQNl3pdMtl7ZGd2/XS8ZRI7x0j2SMq7l0jc1hZe4up8T89pizoV2XNFPAARl73zVsJ676
7K2QYknQ+0jv/s9prNHVhcKzQ5yI4/bMymzLdmcyb1AHfX5syU8xyjNNt1YXvolW/vzTXPjh3wsn
X7p2yfr0mEgBziVOjGl6aMCotQLXwOC0gpjzlBQHA08pmxpM693eGIioxWrzIlcMXUxTP320+p5t
UXMP3AtAlTBNU5ducKctEByp0H5hp0BxLVxxv6d6TDVKOcp09dd2UN+eWkLbWR7TNND39Hr5DG2h
eLEVAJOz9Jf5Bre1Oz6noQSGq2Kiab+IsucWwVa48e/70QYTosY/JX2WKa9CS8Td29sFCi2mgGUa
GStw9q8XOMtN4R8SuN1S5WCJEa8XAqDUm0/SbNsNDKvHrDn2TTAC1dR8o4Uy30WyrpZMzy+Zl/dQ
K/S/PGV+6Xn/sg/c8P4Sc03a3N7au3baNI+w2QUYrQVnZpaaa40cWnFykgbcuMWAC5wnBZ8kNyB0
8FpZvmRsAI4fgd6/EvL5Nh8RsyRMTP27PMtO6ww4AZ7wj6GJm8Gxlfx63nULDD9Wpkr0umfRS+rv
Fye+3PzHTiPcFu3jPBwBtmPsjV7dsOdJQq4i4QtjsAgjzEFcX5Jc45ajQ33dVllKGN2YfbhXqyCW
avIGPx3aibACWA5rfo0YYGLcEU64Wq58iAz8c4sCq35otiQl+OMusmIriq56TlbcPn+iQngrDltX
GtdtEOTev7HV2uHj6YpVLTKL3xMZ3EoR7u3xIjAXlD9bDZBdWC2vCS9Qhf9jghyi4C3Dy4Sf8usE
ZoTmZ16lMGZY0yE3epizGrGzWxQGJxFz3wY0zCXvWd2b2vpZ6z0VAIYtj3vfytyU/db620YZWVBW
i3pa52WzwK5U6M9FsuXyJyJuyc0bHiLiRXkS78glQsPfVKZrqFbzO6s3oZG+oQB62LlOKLVmSPST
ZSDLJdekCz8Oj/6yo26O7vpXusKavPZbyBQY7KCDvVdtXgqB/BXB3/mw8k/2bQmRmL0Na3xS1VBe
vFuCHVbTdxKSV+cmIK6vDEctUasUW8PiUZCCXUVfwgN1lvkbphb7d4B/R3eX+AG7mp2Kz+3evCEs
jpS4N1g4sdXHTpE9b+221ECwDOoq6eL6YeystYvzrBMAqNO8MK59QfpdR8qx1Hpzpp9jexrPl3OF
qdMsyuAUgmSCDKokFO4UelKXjLvgQ5CSXyQ2E3xnE/cpbclR5DDXHgzfmD+R8Fxh4NyAZ1r9AN89
xrqriUSGPaI4qCUnXJOJmEY4vJZraaSnHUkC1v+jSIlKGxO+nLTpr6+DKW0oIiJ1k/TjLDzv7uik
zUfJ4WrbJxgLzdtmpCXJrBwmBmwzJzs0WWo9XIlNrR+jUXLq4eMj5zQvV+h+lJTjJe0YrXQLWnCF
nACqLRER4y+l6srFHxLuH+DhGxOWYTBeylW+X+ERRML/q+0a9MCubT5s7dargtagAABZvMGEcaER
TqOaEfOf4O1t63on3wP/9uYsar7da+nhecXlEXQGH4OajmKezb2JvPJ3Y7Nn2X3R6g/isj0fKc5Y
SRtldrlajr5OG1ZLUDsOhlOj3Nb3x5OovHt0r7Int5dMY2vi7L3w9/aIagiDurs67oMGUGtWlOEf
aum6HR9yJjXK3renSK11okANcIdeWbZh/zC6tkJd1/1gtWyuXdH6GAAn93Y6vr9w1U1sR+rNLpSd
P0tt1qsjzy/a0B58nR6myC1Y+3OSTV5eOIvrED1jywzuDA+4/4ERCT/i3RxAhe+zn31lp3IuPTtS
vUQ3EA3ZZJySoAZ/1HhpSe3BiKL/v/zg+5N99gefwcKim6/mh9Mx+vtvfi/T/Ti+AiHZAu4s10JQ
acKiCLy3s6PVzEkEaC6VL32nks3aHoDFU1QPIB+k9plEbn/4RfI9KrPCB42bEyw7dnOWp46pyPv2
aYTP4UREAcYCLsXGwu+G8+0PMRpiEskRFNZcfWXIHv8hTgtTDykO5ur8xeFFWPXU5xqZ8ddRJn0x
vpMF2v8wLLPQBnunHA7vtcruaEbZBKDihY7QFfjYCypEyGDFgOLA1zhH5T1g8Kz/+EQ5+WqPAipB
VaZUVG9QCZ2KAdEzsxvJ6VJ2/P1OEATVF10+vXKL+4hIFFKj1h+IEw/17sS64sZ9d260P+KKoi3E
zDHCVcwfJRZDlPsQHLaVJlCQ9B8YNBQ5mzVyT9yyqAEEFvqSDum0yqoCicx00EC+7FUIhQhpGF0r
zpA5ojXW8a9d0Y3/5OWhF5l52xtoONwSRdxB/VogDf2y2+LSa5FAaPxIAChHVR+DT/S7zbUUH8KK
wDtzfNmtl1GnVTsQwq3gtsHS67vZ6IBH9Moq6jqD5BwmvoqF8dRmGbZpkpQ/Qqy2GGwLynGt61Fc
3Fip6kW+THcAdoeQzBZD9ZHOZIrxNQ1dhV7wPY0O+QoseU55Exa0LHoYoz1n5PG3mTrbIabbz1YU
ZPmns/xCjQAh20FaApIOvpqe2UiaQdGVSWhAZzTLmAfngRrXWbfO/4oNsCgxX6/ArZX8TQ/MlRps
d6v+TA3EMaSbSB/ck8vYfN9CrpgKH/zhfhi0b4ximCo4L4AAef9TS6BqLl7TLAbIpk5zGi4/sYP+
JnMhhKsgAX8BzbRJJAS6L3BAxqhVx5RXaX9AWavfgDkKkh/3p7XWOjGxkbqu4CwQ41fgo26aD612
+4R7VIOwWYTdHSad8nU7GBfBYwa8VpERUS4rV19Wdj5jBLCEk12qOHtc/VSOw2qK3VF2uREQfKg5
FnbF8Yr9oEARRyD12DXWbC8F0SGe7A51O6OxRUzfNnc+xf/glSnLEEDJRda8IClwVlBkD8kCn2m3
XcUeR6Ix5Re70maKpnm70hupxbr2L4FBkvplgDAUJA7r+XHtQsYYHWEWAjxLe4noYSCYiItL8fb+
VNNZg3Efui2wSpwa+fMWwjJg/JVoBJccAA60nj50jlWGLNRmU4g2ZTz0ZYbO4s/xhLvXwzxTaVQM
E/1R/YuayH3xNojo3SZxcCPfbHfwgfPNj3VZJDdNoIxWMO5oifYng2+14tewqJqsu6blfLQkz6kc
XxVkoB9CoYAUN8oYb2Jny9wUl/lJ5k/sk1EDZEsxjX+UJuLm8AD7yS2A54YG4E91LG4so3Js+k+P
aEZpHezeZ7YM/A+mMNqRCnox9UY4AF3NukwYJsozkLR5q0tUzvJU7tATqIGXf7pnLKUVWxHSCGDR
cGx0dfSINrNELKcEiST+0wfooLFJchg6nPhOIQAzsrBW9xFQiKqoWpi0jhS9DLu7YhzM3WQRIUVO
6IG34Apf6wzKBhnoQNkz2ulcquAcmqrxQXJSjIXwJsOFdP6yi0hztyGGZnhJ4xbHlOht3yUBAm6e
8b4IZ3u+etpDPHIMuqs2DPdkuMDZEpIwxDNjqSKF+biKkMokrUFQWLPneqKCiJ9uHL/KKvyrgeEN
bmf4MUsrtjUVRfEAbDYUgwUgTqrI81dsnT21kbpDJFJ6WtDQCPT+DMoZP1Gwg2sbos+x5Fjs2xcw
HqMWSGpWNkO5NYO+Tr0hwZit7JwbE+6ASOVDA1QkTP/tPvM/VwpBf4rTmwFBhPtBIhNnJN3RXdkh
Zr5eGvsqAiRCFCQ+36lCx7Nbqut/cAPx6OR3sXzvyPWC3oLo7NAz15flnCAKTdQdVG0lETKsa2v7
EmDgpH+RXI1NYdxDZt8bbxhvqKYPc9jAueZBA8jySbSxwoDdGWWI4K8D3XA2oG0giKNboNiuTA10
Rqwel9BRW6rUhBRhH8vWBv+XjAgt9JFDKqfwGRQdYXWE5wttp5ARSRiZQ3jPNenxIrfScV+zXvqq
A8sTXVCnM3ieO9excOSrcsL7eMEYKLT3vV8Pk3P7LruLMAsLfoUs7mxWdOIPhZl4eOQH0u08pdx/
khuEFB9YkBpXReSatoXEqSslQTlQqCx5WDyLhScZKlLBzIoj+RjT3Q2PuQJn+WtsKUWMhPsEat2v
EKlW/7FzUZWJFQAFF5mMwDrt0YkBKL6MnDclriSHhR6bFkEH6wyhTIHtMuPKTLLTMlMNhXcTcIbz
kmp+03r2eMjdEf6jEhn1zbW4RC75Mrky5jemeCWh982z1AS4TnkY0+xCNw3AVviEzSWfcFBKA9kA
9+fdJZRgR+MSiT4oJcFSe10/DmF9ZzLLzu8kltEIpralA7f7M4ewH2uXErn6DsG9mMJqZi+YFzZ0
6hXrcgzn0aKAepKUEFkUbV8S939+VTyuumnAow0YydZT/nN/2SDDwgBAmMJx9shvmTNAVKLpgFE8
KCjyVb1aYOSwAkzBmJP+udIaimt7W8ZPtwQNoIJwT6HDf0g6ZeyYZ6IyuZ0ix8LztlQLWiN3FTDz
dbK/7VDX872k/qNsfBRQFaZxyy4N7049t00eDbGOqqGzvAtSIS2Cf4GlecYG0D563lRKRel+/ZK2
txnCLlG6Rs0mVJyyq6ZXoT1v2JPfRDoclhj8S7gD2axPKaWGwob96yrMklcoqPMmtdKSaOr1+9+1
5m38vkBAI7Vh60CGyVr73UTb5Hbn0g7+cgvNeWAM+JdARcckwuMyyIfLIG664JqqKBD7BjOeLHA6
SwdlL8FVRtRqqK/ahJUjBTerU1P+gZJIcbzlInYpFLiSn9h+RgxLLopWRO37j1IiSn8ibSgjRM2J
OqjwVGH2oMFz+Hkx5FxiB5VjkPgunEK84B327tgcz19XL+dfbFPnUTWrxgd2leps8vXhOITw06fN
ksCcePnw3OJDALDOlSwhPUTAznGwRYSvz0Szlp0eSPAIrG4WBcgUCY5D/52mOMBEsV48MpDcVkP9
s2BHRKq9tQ0qmtzUSvY61lBlyMFLtBAsptrcGEPt8THSFTDijcQXTdP+8z0VITRxDKlTNI9iLU74
VHVqqZk3ng84cHudnCaGJKIQ+PRGhlvWEu5Tyak9gD5Z7oUwe4mVsk3rtNchHgi24UFhmZctP7Yu
ar/FUgqdNGBGv3KcP/qsKe/rNbyAF9Bu99jMNc3aEJiqOX7EQc8rhUM0hz5JhEmv/LAfyNG56/yz
Fc/UvmibbMaLyK/jcNjgOnQsab2Yd8OYiyCwXrAu/nWy6tAAT36Ua7NiYJiUDlZXY9GuIfHQnWuv
gpxh70X8ioERQJtI0Evt4cQogENwLa7Gmp+e7adr/xTxIIxJDHwUB8fkBprJ3yvwLhQOLDLA6aTb
czp7gB93wltPsbHZeyM+oKMKPsePJCHhWVxy4TuzN3jZZCtf/cm1qvE3Vq9De//RRNPrsuUSv5lW
oRLRAbfGDHJLrqo5CxWVT4MfBeMHIguWt+9MiU5Kh97Vx+J1PgePlzJdMtIsvWzGVbNrVfQ8F/j5
VzQx7pf2VHgTUe0IdORj9E2HmFnXkcdKWlD2cqoCz4WkVAVfP2OatxDKtAGhCTK1s+xhxYjZOycy
W9AjelzlQtHbkRbHevuezHVJXvzdJ4IrqqdgUb5cdmVFKrQW9JFt0kSbHbacsAD8OykNMomDbA4d
fa+6oAiWxXgceZpDrVWTliaewqwJn6B/6mLGcmnCab3OFQBtpebGZR9aSWT1HxhtD6aym+KnhFfW
R8wW+ZXWbeuXWlR4qzgQDWWc5F2e84SEzSWJdJ+V30PSPZgvizOmelhsSgS5K3oM7EEB+EeI1Ylt
vm65xiIy5125CNabPCdHxJSecmUzd6eAdtnHIr+ouPJo9lC3tUFi5KfNhtZxNKC0dC0RyS1isPK6
e8IzXtYCiqWyTpiVmh11RXaA8GG2joHEZsql2FCmcwoTcuqIv14/PbZAaTBs2Fy5PFZnlOJ5PS0s
DgYvEUr20daHDBBfY6sOmL7B9dVdCkzLtH3McyW0NpuKrrbgNVPFE8iUibbSzORt6frBGkq1qcvM
qYvuxJEG3mLgPkEjP+jzgb4AnEwIRbp3CIIUGpQ+zVHANcX9eQMWAwnshCQegTi82VIvh/iTwvuJ
8kxeAolSFXM7uyIoSS5U6/UQLyibYBKepuks3u0QxYD+Pa7BrPkd7pOVD3I0k+wrsyZrD0/FcmS0
8bOnq4zjyzx8JMV876kuX7/JdI8AD5ortWIZWmUDZOSdxRg+aXLsJWuIe4gbuwQoGIzMGoxluQza
6jTBWEWjKuyk6J+McNAoZpwjbmzyd5Q2Tq/02eQB/c1Eus8UOg2CRJ1RbSJHiBOkLtlcMMRbvv/f
ga8Qbv4m2AGrVRk0e7NvxbvwseseOF6f9DSxmzQRrx9/7qtDpRONab/rZKqN/5DXaj2j443F3fzL
rAUKNP03p9hu/0STnknCHoZ9TbZca/koaFJ3zcepC6ZU+SeAn8v2M042RUIXWB+XT4xM/7qkuN2O
rJqxWVJ21WrLL+I56HzDPnaDiv5oq1BhwCXyUK8RggNeX4phjDr4kGXs+sCPjetyqfrPglMZZyf7
s3Yi2NVxAbTKyXxPWFw5WoYrg3qGFZngHczWWfK76JGZ8jQu1F89y1YTomeeG/IDOYQnNNVg0M2I
MX0qy1RiBqHywPISPqeg7pIbRB3aCdeP91Ol1kESgBWfMg1LKwihk2N3IfZl/6yqfCNS46GYGli8
eD78POyzSJT6HNb+s+rTZOij5XCJFO3MzG21jJa7zT+jIYu3Ru+U08HWIejPuny4K61ilgDM0I2O
kgedvGbk39NnaapDuKv6xAKgY73VzdHZviQ9I218jiLRXreGwVPvz+3oI8BgWqupY7J+7A8lYKZW
QkQ8Pe6nOFFMogP2gXFIVLBy1xWZENsPyHAItfRw/q5w+sx8SLLMGEWD0wnXhberkG9q5uuIefqr
ByK/kQkwhjOr0aoNMVpfGHB8uKurV+6Q+gggSGVYHCuciz9Y3ppuuh5R9oksx0dabWif45qvp0zj
m8ZK0FO/HM46+/pNTCWE9OalZqEalRNylUlc0f0Jp5zzl4hwa1hdJ7liz4dk1ziNQsqdd1Hwtsun
aoYQg9ZbTk6NHyHoRNtoMTASEfT5879T0dRfK1NB14zdgNxjr1CwkzF+jZi70yWgvKtHywlZnecK
hpujJqNom/d8rlvun9iaE5HtPMc2HwyIWIpV1urIeUd1pTh6XAR5vYnzO52M+FwkkJz+zJL0GvaE
QND5PXxupQfzJAy2pjJy7/qpJgU4cw8XRhyDe9rCyHpGADc03rptGXWeFuL493Kni4YgUiuRdzk7
XroQkx6C6zk0SXDBplroJXJE7MiOfXPrFs52QKTVKjJDNTLqYSb32p7rn1twZuIoblsClA67gZXk
GckPSq/41R4lCmf/3gdUxi9DUkd38cbffyQHaRpShqnUPG2kzXeYpGLeV7P/llBFcK94A3y27leA
6bPKg9gJ59Jxrsw7CZvBK/OevIf7ONFHNAFHcSYeaz5GCmizfJ5IlsVjs7hYkiUUO3g0sAGlC0nS
StfLUPtguhnizKjho7lBtFu8J9AgyeoAzrQ5TyRe43/J4QSIz8BV2VOvqW4B44qHMv/x2/sOy8fl
TOfW0ipSDAY+/AdWYksZHIvCFQLh3IyP8Xja0HfPTF//0FNpaWOE2TVacjXE2U9Vvg1UWEl1jSL4
D/A6l8hjbhxitgA0ihBjM07pYjVhdLKtAdR7iapFdVUOnG8xLnlgctxGjhq7tX4iga0fXDT6flRW
cUCHu+vZ/x3IOtEQn3uCOzq+5GfcqbZTHBSlPNslkjQOSHUNDpNpQx3OrhqP8cjtOCix0CACVObf
4M/V37+Wsb0cVZZ11sK/Xgl4hAhqf5qSWAM5C1Wgc30hYamcNIJvavlePhBkvvQz8DqHzb+4jVyk
jbse70hHzUgNzwxmxmBkub5+Z2avkhJY4lYBQnEyR9bJXjswBNBu+K52uXIr6YapIg/M7RD8wq7m
Ve9sB1lnrVsc1K/Bsl8HzCwXkgrAyn+TemaSifgS7JBCXXeGY4VgdJnVNRG+nlMTxwbcbeTrhLlS
iHvJPNcpNVWaYvR03lhJeMREExIDuPtJcxvxm+yK73pSmQi0HPc1npxfjwWOmUfFzJJFZB88NavB
BQVBaUOa1aeJsGcghDxBoYpDHpfnrDA7BEqKwVfBlaW2PttXX7bv2h8Tzm8ULvXwv1x07S9nSGWn
9oEmdmS1JcHLe3eqPQWedhKPBGu+dVwboz8dQdAB5TcDc3kyCLPLIXiJ1P42eMqbjBh8JMC50jbn
tft98PFbit38PeqJxf59QWburohbfRzZmzbgYIV9jeGvkYMnu6V14ZcdK6GLQIYu9SucYni1Cgmb
IaYYZaaYgAT176h+/rwnrhv3c06gTqHzlNJ5q4DdUCeUswKA8v44aGgjqHQ22lwOL0LNK8/wDjkc
UKeP62oBVkR0nAN802DLWhOmLYkR6+4qOlHKgZFpzzvKNWbXLqFtoBdwudHKEbESHWHr6OKRsfmr
bJPIIWAtB5V+yWb48humvtd7Q2qPIaAY02CmiqxL1Zjwgk9K0t8ZBTQYjK/wpTbnVCjKviax/sKJ
yfaT8uN0vxLWIfmWMFbOIFJU2j2n4tVMOsbBDM0B5Li9KNss1BOlfPxBqg4PBaf4FXqdQnhwkPUW
LBrJiXGVb+5MXbkdMQEOnTeTjYfQ+0niEvwjmqVvJeLkmCV9bXJgv1JlVDJYkgjh2z4L+hwYimGD
0EFJjFCtD//PaM9EL1UPA2at5WYzerReHufTU13hsnKFWxkUoEvswvZd+UViwMGNnF0RaYfYzM2p
raa/cyAvvfOXbgp/azx1JFT94fJi4c3n98mrEG9VNSExMSrjS8Y0zeEjLLy8wVEJnaEk/dhB1UH9
mm/P382KzxZbQIooz5pexfqCEYqs2KGOoqzKy54xyuylKjd+D69wjckCOfSrSuuNZHlKr1L/mePq
8YhGEXXK8cJl6UwY0bcAZJFsm3SXf9VWElIm4y2704oK+x3hncWnlFcRefQ7oJMNlBGkYdBLVPcM
Hcy+4eeIKmBJ5ig3dFPWa4+bvrgmqPZghMnOtaEiqIQsSc/+xKj9vkfOY5/fSFiMu5GRAAyMkUW1
AK4rHcDMLLglkevzz2qMoTIBkfJD/zwo5l96m3WsgUwF/dwTBZ8063F7yPxtMOewTUxsCNLv/iTQ
D0a3zeOY8soA55g/plTxkdySsouAoU4XyoRJ40R834u8YXcMLrwiCC37//xhEegD4GOdP6CRhA4I
jPu4RDmg8FQgvvte5+qFGnaSmP1Uxee1JtUb3iJiNDmsyBsqPPBZoVmTTty/+PNtFMyD7JtQfxV2
oojJ5Q01/HFtI/Ujn+Etk852moXIPT97KlciSd0Gkx5huN3ZtxQLZwcPssj9HqVsb34LgTG+oqAY
X0Nz+nAunxWoffGanLSqbpVo2wIgElyrhjASynS+BKJwGn8MA1o+AtENO1QZH2VqBQ1WfSSDH28+
++wqsTiunjRsSj1Nhg9jQUHwUfDvLkgx1FhEUOsOVkV8+L0Shmsm10XiaIMKUIKi3vTVX1jK5SWt
2zXuUJJ8vxzXdqa4hRg+vIDAJUAPgCE+EG8BDwDzTHkFEi692lN8JIiCC+pcWNJQ9HmujzYUBOjS
qbtEkrstqHD9E2/kVpG5pPDnyJRmKdSDEXm7H2trv40K+aaIbG1p1yUrwuU3a0q5jMvy2MXVeBbI
eGy9y5m8GZCuDCwSS8rd1SB91lO6haLsdRYVlM4nWcX1fjqbbBO9TZ3Sf/yhG2Or1mJS/megHa3o
Exa6uFt2xFrT89sKYJJ9BLrHg0kQ2oWHLiKmBJuVT8eZIx4wJepu8dMTnf6Blv172AXYW8iLyNdT
dytnLqGpG2W8kxlRgi+xCuEVUQw6FLOoo0phq+TljIOJE05LzHnp/CDdtrUGE4fvBX0WKlGeRQRs
4A6GcjpJx0ZGKiKsVTt2dgRicWZrnRdDi1Qlzkyd48W+SHGFqJkw2ywPoEWsKBMPV/5BFnSvqm9S
7Vha061J7MN+DeyYScFiyaO2vH8p0sU51p/OkVxjrQ/t4fevgVcZvrQh1ATItcKep5iww0HSafx5
7bhg2cdFNOg+kCuZyf1sxXEgju37Rc62Dti9Oxb0yj77UKNteKKEgFWhFUGBrNfXbW5pHCdpV+XL
+LRI5q0mbtmCVij/PSLm9+oRu5KdTYKQu1jg7xY7Nb6vz7h4O+3YoZnwt+SY+mXzO6Mvor+aPsmc
mnVjaAufk7m4kEoFDpcC1n0JK4HG4XVPxbVYIUmi+HtDNJ7QoFgKDHBGDQKQkY8M+w2RjOaoR5mG
i4St9O5u81UuXOY09bN/uG82b9+mxf9spSWkzUegyR58KsI8W2O2u4gE2o46s/ReBnFGbOMcRTuq
ry1As3jM5guBrJL3oY3m7KRDyON9yuSrjqG78a0UOTi2vaHmXS8U3HCtqTOVN9lxiKo9nOK7RDh/
Cl741y7lltI+/OoZyzUYAVTLybO1feLt9Fpob+ov4p9qaZTvygai+Th1Tw61HC07aLpFAyHIA6+x
EtsmlUo63jAA99yTjcxchVtyrot0PSSILWl29lPa8Svj7S/9Ltj9+eOeNKiUsJolADUjjSP3nxfe
FU2nk/LjlPLADfMf3tGwWZnkgXc2qw1IgypsVYcMATytvEjB6Y1pPlG6euoprVJPUaSy15boa44H
TTuNhI8JHJcetBtBW8eMNA1gqE4g2Bh2XdgPL5ENwPdk6+/qZY6k7b5XHl3R7oKCn1dVaxhDzVgM
mRhQkogu8N2/FchEy8s3jW5zvqivjYm86i7Da7677lzLrD0aYOx0SReM9jx58jcDJq3yYDknf33F
kKtNYcnYALSQxaJjWu9p6FccmqF6KsogUfdTXmS81w8WXogLBlokfc56XVZEJGKCOgr0moNgvEi5
xCfkBxqyq6Hx5bV55pqCSoMRnCBpVOYiOKJ5s30lPSoSq1A0QO4unMQ1S9cHkQ2yp258MdZKuooB
7TDhyAE47Va+tOMXqqg/B3gqG18hvZs+JhK0GmIBsImE8prV11xJaSIjHrrbi8I8Sfb84wI+pMJ9
cJrE7XzwMsJku5J70As4ky24fR2N+Tpjfe9uQkfd8nKEwfWl/VhcLxlnfV+U9Ff01IolLJVnk3N9
pErs+5frHDPGwOyGD3wdBIxQCCj13+4yKgHafQi55+nm22MHuNjJBBGkWMD9ONwwp8XcDp9geRCN
A/+uyozZre4ixiaBjC25mS+0BIai/OFa7uzhebvjANz1pzhm6ghwGIRrSCmEfIMANrQyq4XCoI4t
/0308i+Y6lW7sdYr+xYY9ktRe9f2jbwRvU4uJ3TUmHdhvJh0E2cvYh7ILVAvr+RiVED8+6X9LrTA
pBSPuHzOLXN0661boNjkv3qnLDPf4tfxJW0bCsjNntg31JOBxtrkUaPqwbeCB9SHuKLIBM+UUjGp
Q9oV/D6FELKuBs3iwl4s9qL+cSRZF5wNubcBNM/uTOU5NopIpdvZMh7zBsW2BvbFl8tZ0gEdLsWV
0kFW58cofK5zFMhT2ovQURR7cFwkwFx+vq0RgYIUymK7QwnDRyUW+jqeaAYsG0sFwknDeWpM8OJ2
J+N/LxYTITDqqHW0X+z5w5Fh6Yw1t8juJwN+iJt6jWBCaCoVJzqInD9s91Bg3uDdn8p1sLlJFio+
mBteNUUwR+8k3jzDMDu2GGr2n+YXhS3jQ+WCYHb4kFt7jbNTK/vOb0xs3AFvIuARZN2Q4JIF5A1i
KbsIOthDt5f3nVm43bzRIpXNY0TahJmLRab53SMnbtvAKKmFt8xbkZtXHSdw2WPodU0jKEA2MQ6x
IwWP5KMzmgoUZ0HlolEL90iVx+9h/ofLeJ3cNSbciUlWBEmMY/+ARzD1OswSsN1HZf6HqoQT0oHp
BzpNe+Bngcid4SlT0ET7TeZKRl5HgaO1wOCNxKg2APY8sJPUzdfG7b3AdC0EMUXLVO+cslCATbGo
scsOiUKq1VLt7BLLvksmFtq2ias/Ji8rE9vEujpIkD56yGM8u3srrcEaTk6ke89ftCZWPTia+fC/
7wG2Y55FOEdYSqyhk/ruJF4FadnstcNhG4Qed0t7j3FS8XjbcvX4u3rxtXNxZ4n/Lpe37hgDsC/b
DNdjetuVffbTEOFF+VbhktUV2puJJ6mM2FdJ0IOhW347qlRXabGjbYVxw0GbWg3u/oFWmDEVdheo
9n1Tym5l38FaZA1zrUAPfNq10MsQYhodq1sogGpTugSVm4OHTZyTN8/lQ6iYkAA7qDsqIkph1t4c
trukx3kLRYrUC59EX2okeETN8IxG3J+3RGiOFKoXPQTt+5WTq0hHSEwIBpn9EIck7RYt5t3XscdB
UWaDpvDR5tuUzxjDWOnt9eDomhaE2cWXBvAHHHhpSa4XFiDmiq2on7IfSRZEm/3rUNbiHoOHVmi5
A6cZZ7M9ZLKfckVrJoah2rTYd1Oo2wbn7tSP4VksO4jjUm2m7NmR0CoFHhr0L8zecWAW0yqUua0M
bWCYMCG24qpDVfr8wLTExBg1oAqV6BIrxVBY5y/IyPkQoHQpALVMJgBfhilicLzdV+Np+8zptj1l
f211SAkj52wCfQ8BPC/M+zHIZUVRzGeHq7kyAz/IvfZ17b2TClBda2sFqcLPE/XCEmI9/4ko9YCK
8KXVy4X7ZCi7NrELPjBW33D64C7On0ETHheZhU84X5UKNVcvQGAtkHGO4NXw1PxueDCzWHrOOsH4
iOGGo8FXJ3brUulurHgZpr/EVEBUl+nuaJ2e4IE2DLd7zmev3DfRJPHxO2koxdfR1Ye5doLU3XGW
Md8CxEygEIOCOuSqwqNAX6fKSdhn0NofzCJI+uVjO/kDswNDu9vdtcPEBmmSgvSnqnjhBBGr44lq
6E8wathZ7eW1+mo50GxpnmM80GHgbBa2mUwvUOLgsGuRna783OIHlhhdeFfiKcgK4juF2YgQl2m6
ck821zd4l0zI7ILzYVi0Gj9TiuI6sO84Ew2NMelW1omSfiqRDmKNK9W8zL/NHYoB6ZBnTDxmDF46
OYKs9yHAsOyQZga3c8vMluDIm7VXwSjltzXSh3xtaxnNxMUe2/Xk4/CfWMnbPPMIgu753p0f7ljI
p1bj/pwY96XYx2EnnGZOUWk1oJ464FLOIDI4AQg3/tcvBYB5OIwWeVnMardgyU9DfUl7AeMfP39J
VKvYkcebEWc4gPFutcfpzRXLpg8cbWcY58nW2IvMI2729y0NRxHVZVzuuj7dyjanXTw0qndgKRlh
PtNqXyRn/vLbeD+sBTwo6DVoao67jK/1YM9YEM5q0drFUhWczMnT+CkWHCFJKt/4+p8ODl9HsB0z
tgnoNFHlAR51+vsRNMjAIKmh+JkEwB17DEyGc0jNKrrnvTc+/BXAh5eQgjFaQ8YBWm7OoqudhH8M
wPrB28l0UywRbPZKHrINJQz6SLSVFx/bljHMw3x9CqV2pdslLHyW7T74V6m+NwN2sGKYJzdTPOI+
A+bPzNqCf8CFzj+agsX9Kosr+hdzXZU5S4zFNmm86nYNIMTxvtMX6NtNIE4Q2pTNeRUD0FdkJQGH
vek19fSLkhet7I49vN4Jf618h4Dp+948Prv/8/5tMzuH+GGMA2mSoCyVSa781LVxm2yZjxPfNWdP
rJxJoewo2FYFhEqskhOzw7TbfSpwCx4J7eRM5do7CmeN7fAQrhASmWlKSVUAfbCD7frA7zo4vjsD
YYWlmGqbgL3TvxBbiKjVChrO0w/DSOxjqiQffT8zz7XZR6TBS2gVDyRa6XvyUt/41YaTlAsunPoH
JB3ojO+Wk+99FjZVXMPQeXBzcF8H6XnHzEt7b1hmzNStURocdpviFM0XfnTrFVc2GEYXA5V3Z1yK
lWNCTMAPPC//kwPLmNXF6Uim6eK2tVm5CuQgn/Ongug62YVY9z8Yq2YJ36sfyWlutfDOB8B5ogW5
nn1lvQBt1dHfKD2Z4ymQB/9XCpoAwBCorNr7oFDaoHQcHwZEfizvH/SuMlgbGsb7ylMaeyhvZKIC
ei4dYR5OtR3m01ztzHHhBtFnZ+mGTanFGRNhFD9ANUDVb5VzeE5WTp56JZgxPkqMx1fGW5YLVKSm
B03tEtUiHBcJYEBReb4A7dJLgIKTmz6RTRT1llh3FmMBTc0E0WsA9mlzaA4bVSlemEu22umkNi2t
l5gKUXlzicBDC+Hxt2pOQ85PsZnx611MmfcYT2/UQnXdJ0zPv7Mi3H4iC9DKYkTia53gbi/niBB6
XmZMFBZDtqTHc0hGWgo4N4T73SvxNjv9rGXjj1HKakmxAi87gnIZNdeoMVZKzrs+8i/swhIGSPs7
EC/NsVqZ0m/VMECUaVfopbr8Gyuhs1X+mkB+3Tw18oJil7N4yvz9SgO2daXXwFe3seU0QlSmUqc6
mH9VgCDTrMFwZBsQwbqB22VSOOt+XS9gPfI43El4hUyfr6YdLIyaokDt1e3U7Le06BcgFstLLK0L
2cM1o8tJwhJqJtkxHw1Ze6PPoAXv3qJqr+sDiJK1SNlN+UwkbNWnscYPhGXD2jRBzTj8RXA/AKGa
oYrh2YBm28eu511W3cxXxLScDf1OoJG/TJtL7HZZ9CpiJLim6TX2G7bWIPAoBsNOm0BdIiVj0GXH
XIjOL6DbzvdcV0vikJEj7cvNNTxjtYuCU3VMoFUJbTbsEfEvkCMeoWyB6yCIbFQ4CrYNfyYdNXuF
x9HZxlFDNEr/vR/0vxPh/b0pCowdmI0lb7QgsVgf8Cdbw93dJcZLu59tpKKO71rxZzzn7BOywg62
RloCHsKRZG0ngOtQu7R8QA08VIOIYQHJg1yQOvGBju/IRL7jDc+n0P848tdQz/cxamXFMdpoqKHP
yBDfou0LgexRnoiKoO2D5FD7c735x2EKCxPVpY+BvViwpUN2AJ+uw6QGFW2GcSbswg+44OyDFnXu
MqCOsFccQxtjmUzygQjv/yqXFqTIizomEZpfgY1rQAqNoDPOEC8VBXIE1aymu8Bp+l78k9zC9NQK
52mt1Nvm41GG1qsw4xz37hFdi76v9WhCp0pPu3TpV3SOMj1DMdxJjNBTvco8hrXLwO7+cyWApuKK
tkZeWeFteP8UUMnV8ih3Nlf5dqqfK8MY2dIV18yY2aZ0sVpdWr0RhL/FW39iXpB7qd1EFbjECB92
qXNqhcZ8XHxBM3RsxYsCXjktwrbP8CkDeDeAEHgo1ZACi2R1N/YAF9XYqMjBuXiPw3uXfJUvNKrk
QnZ3KWGmLdU/ML6dEo8pLKvOLksO765BNboGeTMFMuZfN74E0b57Y+X+Y08Nsw2ofGGYJt0laRU8
hi2GWB0su9fHqHt64ONw0+trRe8wMFzXgdek1zw5PSqN1F1yWtqhDPgg7qOKnY4S/1/ndWU7GcLl
80RC5qkTzaayVn6Q9BZnxWLhunFofI19v3EvimOPpaaYNicLH1v3znK4mRxAna2DLbj8XHsZX3uo
kjPOfUew6djtmA02WZRsUEYAegLfXx+N53zchfPah6/vIUtv46xBuYTygAZbdOfJpTzAMaVTHs8+
XkZFLQyiHC4R4txkm+6hahxE3RvLIVkFCyRhKrXWvQ3wIuVtSqmf+IuRzlo3Es2nBEjqO6QC92Gs
OIKXnIY2rnbGLLGpe9UDrGghDVH4kDZ5rfuqEsCcsz4P1jcN7NGOQGr2fYenyTcW/PDGamPQCv0O
y2GnH4/hdATdE4Ft7YAGOczSvXmGxlXF7To1H6HmMbwpl+VagU1N4q1UXrexgadnkpCOUQVEnpc7
hSCnNEw9SCZzLr1PsLTtDUz7Np2hnluM9Hj4rtKXH7ZgIzBU/sDwrZR+sg3U53v2L0t/fuoMKSa6
VmOypWWiyi+NX+9bNCI7nXoN4SRXNEtjx3WGetIybX1k6piT748U6/4H1QTmpjXTzeBaOUIVLmlw
TNbsd79v3CftPMF0BkS9AfV4GXBjrE8FE9/c9XcDZdwvNcY3XRbtRzsWJUNEtDzhfii/4UWw3eNa
uH00S0+GxWIhlcpTLLrE4J+LUKWT5AFgzLDun5vEjHKdcX7x5lzlo1bWoiCU8Q0D1mm3j8T34cQz
2WHpq+YnzY+NtPEN6fXW80ZmvyWfZ7yme6ynAHtdywx8mYD+N8stU/bzkppkvr7OrgPChLom0HWK
x8g40rkQFFp1MlutLbVERXLZFwC7rGkg27ITUbPr/kTjr3qPE6VPZ1XNfCbFSD+AhCk5r5cQ/c3W
tPBCoa0yHcEpA03ksy+OObw1s2pqhVPwel95UGXqeWQNubQ7+8Fw8YxQgN1ou+jMubPPK9RvmKHi
rYKm4mgDvMLSVjjAhXI11NTB3qoIvDzVYIALNBCzHGIPdkVTBW821fBoDdprDzhR/lETvGLUUYWo
0D3GSiYvZpMjPRsnVmTa1s7TqIayJ8ljeMXqXO+L9mhm+70R1XcQhVF7c/CARoCJ/rXUvJPbQKJw
rtc4ZEY/7Em+2LronxJCzdn3o6vBeVjS+7tjKrr6yvJtkHF49+bSGuKlvJloOKMqBGhOXceyy8ki
23nkUk0ZgmwCR7SwH0X0/mMTC9JLpzESdseOKmA9O+5ZOvX+X9+wNCxDgQlAY2kRwQbLpRNSLhzL
fA49pqrd/kuNiu60nBWY088h5FjdVUK+AeFnmf3zMtLLAN7hDfnFiWNyKv9EjS/r1MxqLiw5fP6/
r5Vojk9oCL4WpHSDHiRIojIWpZKUHwMzjmeky9VpELtVZDSyvL/sfwxBzRpL3OWbqrIt7ZQlqKe9
3t6KAIt/hPxPDtS75jh8f3cm/JRlFIlwvg2t9YLEwh7eeNNSG6wpUWtbYpPkXyvyGEVwtvkDPMC3
9g6GsmMYY29rU+Ds+O5zRIJfCU+MqtAdwnIgo3S9JhYveXOTG8b4HFDdIcAwq8XPTCOn6sjn7Xhr
KwQfXDGRVKDwATg875FtA1tnmz78K0HVTdR7gYTJe3yy4PLVFI4TIiWJUCvbNBwdCGL0UhU0b3Gg
i9hWk5dugqX6fyy1HmHllTS6KxLhGksS6T5O4jHUp+A0pPk113FkQmp854af9NV6E5mS0f/pfD0u
u5qEgspKUGiwZQBvio0shAUCrJ6I+7YymNkk5OWKvV4yjdS167fB0pX75OPe/lN/pjn9sF/8cEbK
pwx2e50b+7HCk5o/Z5Qrfeq6CfgiMVyzThmSwJ9UXG/39BAY5hSeiAV0wRlToqpT8WgLOI/m2Qd7
yVLfBf2fPv5X6m5j5jtLR2DzltEg0Xd7GXVmi8QdN7A9z/BdrnZ0vS8UTePg4LP1fB3ezbGZQwyR
Sp8Pi24zubhySLl2xBkqy0iKX7T/mplb+HFN8HtcFHL9azLLwseTmmzsVuhC/zUK8pU2RVjtUaBD
g9sw63Sac6FIa78P1AbbiVB+G4pxQRSgeFbRomykCJysPZE0PIorhF5TAdYaaI0eFSyR+1LWnK6C
np3q32GoVo8D8B9eV2XemrGKQU9QxQ/I0jo66IwE2/PQc5EJSckVKTiQ9fxXixJjXJxGTr+vTpbs
qudvFo5xTsn+sJameQ2ixxgTg8SM2FtqYQDFuLmMvdZMJS/jRfbodubKdCH/XgAMdNiVfYD9pNSS
/kmBHOzhwKHNEPTfHxKX0346xFYioqA9hYiS4yx+kS2WttKs3TJ6oivNnH1h4rd6IthPFVIm/DeK
FJFzhwlYmduVe1V5OzLuTKpdf65RLuq3q42RDRya92lvslhp9reJ6dkdPtczydqgRSJ1rzNW//k+
fMldz8hjEiMxf1iKB7VB1hrgabtBeWcgykmGvTaFbSjxcmvaSW3Tq43WWykIrNc5FLHuC6ekDtwa
OgGw/FUxHr2H5/K4VpSXSBfmb52vADQB6V1zrW48umHVoTrt2hGzybHBCxM+Y5Z4dFVvYLLMBIh7
da4uNFxK/Dw32Nh5+muIYE8ZLzie0YHcQcC2uE2FPOpkcKsYCiCxMBkc0mNPDl4CJKn3fuCHFPYw
WXP8XNsGELB5lWREm7dnhNySpD74x/PKGSHFb1A7w0Z3ISdQj4d8Q7ldoJ4+Wo+uPypnI5uGAxBs
oSfuFR8wqvNCAnBxPIzFrKdHhrCizOb0SXJsbBwt2TXA+95TNOjstjvDtAFsMGgDWfAeU+9+kdOb
lDlCnELDrwH1Bmi2eXmoTLosITYPSmdYmb4pLJ9EJd4jTnFoZy0ZtDO3fRCsqJ8q+7y/hTtq43YX
Y/tilpN2hDrq0C4C72gFWX09ONxEi8ChwvI0YSrf4v9JaI9+5FVWoX+pWx0OG8DzPBViRU3tiOXT
0hRY3IZw+yxKe1FGDSXNkNK+shUA5YxL1f1tlA5w1NmCh2L5kfy1k7zFnShFOJw6u4hcJPn82nFU
7ticgAXiAt8XScOptxSD5Dj6ynOe8JUtQVNhIiMci3gmi7sS91qD3fJzqGaE29YqNkKPOUPP7+vu
neZ6w1YqSjXjdBxT2PfaxN4N/z/11Scg6+7ZQVxRAL5t1mFT3duUDZStv7+EdiYYBsumOvc8wz2u
kdwThdQNE0v5OfXciznvpAxVWfMiEblf6DWFxTFvX0dQBaYF+rvb+B/eDhjTFZUSrVL+FmkWm/jJ
u08Zn4/9iiFEkJdjDWwVIl+8lcfBo6D3YxeSJCu/gATO7Vy/w3YREZ4fG/yxUWWskM6jl3vXoOI7
LBip7d2aHqfh4KpMbDnXLvIkzaokDeB5SO22lcgbOUdVThXPgHfhRC+a4Nl0QP5UQ38ux8jsc+aY
DqGlpM8B5lF+gIFnIyYS7vL6qJHKQqEl0Ejuv2KjITRyot0fuvznN79wNRxGCSuMoSE7ObVuHsQr
8DWJ00LAgFtzR7/fNiLVIXwzys4OLPk2vh7LwuoELNBk5QC2iaxh8fwfvZqKZWJjeqH3rPd+BCNG
RIo8hUH6XfFk7L9uHTdWPjhLVWZWmRx2H2i+uraWD2xZPjO5KbxWbYTIIULewKRymZVD8XU9c2ct
bvHCriV7mZryregGoRmc0njeyvYN39wouk/LBJO/EjuABnXzqnqUS4FazZfbN1grvfB0L28BhaFy
aMfVpF18q2fts7x1oQ3T/lctLm4mWCHALrgDnv2vIQTCmcpcQMPqxUJBLk8bFhR+NCTH3oTuSWYc
es5+msKi8WnWcPgO0c85uIuNjPcn5NYTrK6pVD/6KfxcB14lQ3X/+EJVVa6utM/6LwcTkJYp6ef1
Qz7cfyiQJ2QlGrjFueN787XzUD3tz38KNI1bQmmJoHnQBBX/N9z5muYQcMsL8WB8yr5/BGZDo8XC
4fAh5OLY2Rv8Ru3uuTya+OsvYALjk0IoySfiONfqGsPLvez1Igdjjzy67JBB1bAEsl7ddt/TOG2F
O94ApwjHxNmplDLGL7ZHIVqbpCH3mLKBrfFB7qe+jczvm8hh58khQcesNmYignn6O1+90eTvyg5C
A2NBxdXBlLNzHrc3Xa4nVfjtj7pMIazQ9MsrKUh72PdTHvVH9Itf4eSwz2oN4m2Q5upm0iDxRbfW
8rQcT79mXHcOMub59sJcpKMHgwZnzf0ckeeTq8ZcJaplp0NFtGDfNdT/XBUsk8/lgu3JzI5CryC+
Str7/E2pDWBZOeuNbmO3vHGAR1iTx5AhvCY1XiuiJ0pREc6FkocjF9z4+LmR12ktD/0TXv9xoqjO
m2lV4YJKlYRnQU6Mqy/oMHjjjX1n9DzAzIpskkS+hUy/inCdeLh6xS39N0c/CgzHB9KXGNFsk3fW
Tu89PtfGOfd1hI8azSS2hY2bd1/o4384kkW2zXKr6aexNTq/8OHXDvmkE+JS0VhnBbmqU0sQ1yYt
yaqagt/OvSXGYsbvf9wbpnUM7oBNrFK3bpdXseyGwjJX+oQRcCG83i+meM837tKqtPw41EAmYtx2
Z8dnqN1KX1ZhZlMuX3WhOKLcYr/6ed3vRQjIthmYFi6andVBhjOAR683i00XjX5rml6r6XnP67NF
iSaySzs/OYehuzorWH3G282zC/5tPcDPceYPB6lhZppd4cHBzRQQEDAvBZ+rLlvqFtCQ0YIIZGnR
V1PqMDHBhA9KaaC/NdYXYudmLWBJjUj0k3fWdWyD5lfOQ5MAfSe42DVAfp057lS1znFpjiMISIc7
QbIxHay04P4s37KRxAupTwQM4ignVJl1HTbYsz9+kG/Bw+WFM4Q75577tTvzZqiSy7hcG/7bad3A
v+581MX+MklGTS+GUMxuCJolufBwI1vydacXSoUls3fugkx6NSHgpLSWx+73aYFHm+iAPU/oFkru
NWHdXMQifkmc6Jf5c5un2M8dRI29RZxN4INEcZ54P3cb4N7a3gBtuwKxkLvaY+UGercxO/8jw3+m
ragv3z4OtjLmfSsnruc6MSuxVVbQWJuubHlYzAlPqDV/L4sY6tpHzKgMZiqMvCFc7iyKpt7WRvgr
4wm+q7BRMpfCyzQsFUytFCk+T0Tnt5Gr6wMmRAnhQ8vqlSRKAL79jWzpnay36JXp49tVjs2PEJtK
vfeqdgQjOVzUQOPWfLx+f6Fs85DaFVyi/mksC1LvD5pDnGeAqZDYgo6jqbWNyqAFYCgh9Wdy+6gp
ygxoKt9RG1g11dOZgFFRUyzUol5hBGL6/bXESYjgX0E9tLvCJ3xUNIeA/1cfo2vIRWsG3nHLcbj5
0MpG3siMnl8rEaa0/MYe/Y/no/c/WeVZUr/z1mHteOovKSUI24o/rv2hdaPSSkbjdGD1qn4i8hPp
MLHGpFsG6LMQt8EC0IZw66C3ggT2kmckoABP7lcUrClracK7qFmxXoQpfXs6GWU+k+ERSK6F3ngE
ui5HKlXCqA1pYm1knxyMaN3UbEiynraou5KU9VMheYsL+TgwZirtGSAxpHFkY45X5k1re845l3N2
eE4+rGOUjyWBxb/Vq7X0z1OMdBrP8uVp9SWwjuW7tZnljbDu6jyFvdf8S4yR2Tzu+890z8V0o5jK
2YVzSqNEYcHqSBLe3JVKm3AL4Kh7StXooxQhZhf/jWXpXEfx3VzvPKlTmLLXD8SjlhbQrC5HDCfL
MeDeg78B9XJ7oiHu2aYkcGzKsBKPIcPkFvxRDaVK3FEy/isUDi0Mgef6zey9lOMG0kjNIMlQfXIC
f2Ofbq1QfuLOto+k0/nIpD5RhUR5kefjy+YsL9h/i2ZcC5IPAHu/IgAZkW6x6mUMVMtcDE7Ye3Lz
F6n7fzAeCO6yidq50jq5TBvdvvr+8zWn9e/ghR9YvQV+aYyxXHHmzP2aGGNis936l6ZrlZMlmw/z
HeT/jK1Ivz8duVvxj2/kjr4fi+uYOmji1vzYzhpcCbyVZIK5ME6PL3M6ZpUwHg+7Nny7Z0J2QdCp
s3QCz3OabOAFRwffZfRywpWBTCXAVLL3QaN8T7GWwC+nr/hKKWe3pcYrHqgcIGSUKb5CLV5hX3Sw
PJkudEMvr1TVko7Q0jMndsMUqeb7FrbjbOmnekdpOf1RiaaeJGyJUsDG3TRVp0HxQ4itY2P5/Iza
XCkdYLx0ulRf858dCRN8UperyxZsBx0JJA0Rv12PzvNSzmXgbQoXM2L8rqokPSs3Ysgeqc8+e6pU
ib7kqW4uWhL4h+kUXwrjJGkCpW6H6MZkdyiaouVDYJSMBUf3oe5vsvr1RKmbYtXfK0TLaKcSsHtO
Y9Iz0OxN5Ql25R61uLncNNqOvhkh2A2gg5UQvfMoQpeOq8D14Ngm7j58+sQIyC9MWgUJ6Yg0mo39
LpJ522+xt3iFeWTl5umDmWXehX2v1XUZlNap+/TxlNx0vfPeUrnxNlu+ARkWsNL1prBjZSxDwJsc
NI62n15zNKR4A8/QtuXSfwLg18MN/+lA3WQe5TNhO6HddCRpu2a1IN+/QLO4uFjffd5oGhYWA8xQ
U1/5hsRbqrHOsRwN0+/Bm2yMUQeO074wnNVSc/1Skpwc4t95vdCsznZCczb/lDscPqFND6mOoblj
0uc4wlwIc11CO6RwqdDR+KEub8z6CvPLeTWCqb0s2KQM78I/PKGE3+UzDo56cDu9J9g7sDigAwcz
O9id76pKIGA97RYGPUWRezUHoAHqe6HwU7LpcMAZZO/t1k5h9oy6cfVMYiRNjh9to9S545PJ9bkY
giGhibtEU7FxHYwCgaMqoB6tKh6b9pgfbKI3IvWOXKuhmwoW/z16/Ob9sdMgeLGFp2XNVszjdTcp
2nXGDOtQ9LcWTBfIlxgHWYyW5F8nhDQKXPnQvpDy+zuSIaTKu9hDNe3OGzHJYYyw+Xv4LAI5SKpZ
O9KGw1htuo0iysJsfejjxkYrRuGaKlajYVIcIJ+wfpm3bg5OzXPP0BYv5ZQj72oOWfYVPmzHMKVZ
YcYlmP2AapNDDeglikctv1llnEHEowj16AbqmN3E30pf9GKcU1u210LKwYDqHGAoE4+UbHeVYDny
R/Xc2nS14Nyk9aTpa/YAF8MWEtamjLtGQ99bIqFE6P6CI8T0fSj3HXn84em4ROaNZnDd1ZA5WKAH
XMyuz+5I3gi1umPvfHICIfpcpaFX6cGAuohtO60tTq/09KCaY2lqWYyVzerNXDJZ20UitjDOB5xw
Pz04xEMGk+qUbZGcu+vjGObZLZp3OzNReUG2yAxC/JfWDTKkiuUpW6bFgNm1hxNs53mhccqK0PyI
Lu0RjH+t82pG+VbYNAq1cWXiK8+iIqSWIn8TaXzGdFViTp15dZfxClIUTwWi11yWhsVDaP+npBqf
60zCbDyudqs7q45Oa4pJk/2KKo6WGy3f+gCNPNhwT04Nd4sx+0RRITy/qLM44gwpnXXRF2mnVQ38
r7rdIbII/Txn1DSfg0TV+2G+txUHuUqME9hPEHwQG068GlBJCiZeUCYEzO8Dl2V38beFRdAYX5MU
dsH5ybjIS+DXBm2Q3XlDCo7J8tH+acbjU9rp3o6ioUTmSEaiQB7YYfrUQrafdrlrHd94DnkqvzEt
BGbXTLCxkx4LqKj1+kQspKCctNR+FZy+0Xldfd+0lVh3F1SFDsMln3MfY/oSIdC9CaSN7mCO+w2N
RCkO6QLzWUDGa+/UHsZd1HNB6D3HPpOdo9WpO8692Z//+4VJxIQ95keEAVh8YtZqdjhvFSHu+cTK
7VAXAfGQMxTF5Rl4s1PC5I/QMpV/8RfZG4bvLVBNhOerlsc9H8fLvmW3A1MlspNAyqoffbbcUTfG
13/cb6NWdJPRKYJEUSJHu8zcOncoe+UxxsYnS9rvLarl3o8lI9MGvypm5zVjYJ147oT6juL5YrcM
ltkfW3+UWVdQS9nDj0R8g+JRyXuWoFrULBOB/JlWNjabTg1sKyCvSRr/zvXfp5MpnxowlbikmY3B
n34kEf1PsQjJE/UX9gxVQP1l8odc3rvs0WTQ7I0GyjKUZW+ly/uo89VY+l1g93/GtRKCxqGZj+1p
UlEaLhiQyNj6A7q2mm8ZtU5cUHkhW58U5WK6WE8G4qDc44KIe/h8OisjKJouUgzFZujFyROYh4tj
Vf/zUMxPDsFeifF3DkrIqBnnaYMhovLuX8v4yE15UT1xF8NS5bs15/Qv2ZXpq8ol+SJrV3hoXV5K
5U9X/Oy4rwxUZbNbYBAFY/pADGXy8gV/YqKd7vudgIStgVKF3R/+zS4gCM03UUgDYGHXpsmSREGg
5Pg1xRSbhU6PdFYiKH1EDS60+2S5BmadaFlGs5oVoVqbGVvvgZ5s2aKLk4miHXG4bEBJLIKDRCwk
3Is7FaABj//jB4NPMd1hqDLw/vaswrQQaipa84x3yrKCC0WOwrLh46Bydl7OSAojcLrcBOwNN1aA
jX3OpATf1t8vH77bI3axFLOU5/i8Ibv/YX6R8jI0XwHSbXa8+AWsicvnlX/9JYNILLstqIklkF5S
i6Ja913YnzRs+A7PdmvL9mW3+C5rUGNqM71Ayy8FsbBWIeKGS7O5R1B5MHxrNnFTUFg8N5Y3F0KB
+l8zHavxE6xkpf/PnBMy4LPxy7LRLno9Ok/1PhEUETf0r3etJ+NJvJTD6Sp/lC6IId5cX6202EFR
clblhK0EoDnMlDxU5y1Z0kimcHJ/0Z1g5onDmep739Wtf4ZHCRwYiwYm4StASqUvZAEkpg762l2k
tavdCEwt/oaao2D9tA52JWc8e9X3cWw9V44uifPZDG8jCadgPSVF3mhbh06rjMcB8d0GYG24ko0G
6DgBumvcc2rqmzR+T8ivydWHqQCFp4CM+CrdBOTFrlm9yCSVCaGhngP58y2YTFNU/jSkguwMugA5
QVkRpYo4TGung+NdHtH6IZ7+mqrurc5HMDPJGoG1lj/V9cntls1wH1OWZ7ytbxvRWb9epFP8/zi3
dLBhJ/21xnYfhivKqIz1Dn+sAlC32o+M/IBJCuSIkhuaYFmhRUW7/18rjDOZL79CByfrrBNYlMWq
5UsSlavA5cH0qM4m4rkddZdgS24WiPHnD3mngk8ucbASEn7W79R4D/q9yJLSw6Jedn3Yn5L0uUPR
SBbbW9kJvXM62Gc796RQt3XtHiBMAiO0v89IK1h2/Xt5/3ziw9FAEdzDjDxNpyYycl7VE3RX13WB
hgFMk+xum/REUYJQgxkqFioVrjKkf9AMPNOoeeYeUtkP6ITiq3p/rxPyPmhHcPSDVoF+nGSeRpjm
gWOb4slos69aJNCSdbmwMlEL0Sfi2f/QR+Bt/9rT0pEo3DRvVKsKfru6vegWrvn5Y2P6CJu3Le6p
7eO9nkdA96tkZYIi+7wN4fVFcDFepT9XTZNX66WuW061lTgs2E6kzas34dqK3yO8LJoPY1KK6W5I
s3DnvKo+uHy6Z03DoqPvPWV5KuEwxM+20eaPUeXtxYDc4e3iGIYB04EY5LZlaMFE6rgTx0yxd9to
uCXF0apiAe2Cht8D7wDQA1I1xCwglZ3kZVelAnARUkD0KYHlIsjLRCNAaBZDWZTfavTOXecJ+zux
FZbQAZqTO2TegaKLsa3gml3j0ONiRlncw9ZDnWcMKSNZ6airYP2KQd2YXvA8yQRAD2ywVqgGqD3h
Q29Y7ET/NcPLwTEavsTM0pRRgA8T06bFu4i5AoEJBmPpRdHsLXx1tEino1T1ofrg4sMslXaWZZJo
LfRHGBhAlF4KvCmQ/ICo8ZZiN4XoO0qs5jx/ntPz/5HWxFlWafbyi8FMEK6VstydWHpxUy0clfSm
QHBozb1KfYPp/cV931yiexsk+vnhv95KG0n5aA6WlbTj33+ZCbIJ4k3bCE/pQQ9AetqnBRbC5mHL
AxDmwRXb+X5g+eKaV9fmqNsv4xKvChfY40Bwggjmqz2yFT3Q5XBJ8DGgp8ZG6M0dMMEN5gPl1ZAB
NKtjLcds9deYpCl4LYler39V9CYVZXg7J2mRYoU8t0RUig0WkNF+Fl9l2lMb9lmE8auNrCM5Z+Dn
j0GrHUmLR+mQpffBSzVyrrFWMxu1OEIQPTIP702UMFPV9WoPE/i4zHSvEv+dpEHj47vZIkMdhSNo
c5cLV3Ctm38d1FTuhqGME8gKGIBYt545Hz9QS+OCa6GWlHWjNvDiM0i500DN0TKxOwv6SoSFkNDm
8rGQNL8zIp2/q/wTZPnsClR5JNK/CXEea9U/PTqWuHZlj+t94coaF8Eo+7+Ad/DROS1bsSeUo14Z
GL3oF48NLRJZK45M7MMWbt6b2Krf/26qWtYcVgo055tMsuHIbVQ1Zq+hGSgCC4BKIgTOY0ZmmeEI
g06SIRqFvqouVWk5fRFu4QuYeKJrslcLycbrgWWQAxxj1h8hHqtcQ82Ae7I6lSy10eqB+w5oERh2
WADBVAymWLI6Udzs8qYSSjKuzYntYYfuvPIewZsat3fWvyzx9AZtxEnA7ucD2XSYomI6y6Xf3sAU
gef5DG5km4b2FnS0OVACcTSAoUJ5VDRJt/UZ5QOlxT1J2rZOaVQcg0+aR0DM8u74Ucrf7oeAtsi1
Fr1jRths58gldNesb+cvqIqiysdgNhUYx1i2FH+nMpEHbmXo9hI8N1KSv1YfSycoJ2RC9xX/0Yki
jfLGvIGpdzX6E+w0F1HTdpHd7hI0PpQrHUbuA+3hGVm8fU/s6ued3gQuMZHHnZWCkZL0IM5IXd4k
aTrEfajuRyNWqw1ipjudLrsUSkWBjgdw450TAcERzsAVTj3VCEO6Co9SmT0DiJOb/wO4Slu4d4g0
hR2MX7gPM9d6w6Jg+RTqAR0kovJrd3Sigl5QZjoTVHppZY4sRFCbaxbCNy1mdGPx1Iady6aPn7gM
KaBpzSqPeKqg6svMRZAnqALoZqHwF3AyTwMMz7JnOGRTOuRPdivVaOAnduGcNs0FYBK+oxxegXjZ
lvCCcO6hUkMDBQ4GiHO/CN/lTPr6NL3KoU/aejctE1WJRKakcLPMJsF46NSV9s8uqtpI9iOP47M4
Z9OHqJ86HJS19tN2UfkVwsZB6ey7MEzrJhHJhruyb5cMNzR8a8feH0qdN9GxPshfwr6dggf+ueLL
U50876OMD8fzjYwoepkBwxH10yoQUQqg7cfamV01fi4xdIlu9n8bMZwc1SEYUWThwZcioXEv0P+O
zfQ0GVhb4o+/nl+wclZFJ6V4A3mW/0MwP7Usq6YlgPWxCmSSHZB/SUMjr4YSMgXSz6Eq191q14DH
pEwk10aAEbYndpFyj8wDTtNkZ89nMb6LjJe8IiDGaer3RHQd3anooOlpwW8sTUQCy7myOneaAVkI
t12WJpeLfcKh+i9kYo9rvCzcKPTRC+0Ra0B0sN0EHSTACOYWHx1CH9z8Nmtx8I6tBkSMdirIpKFl
JUjDoP0yRaGwC1aCz6tcAKwUhMhxRRfegWEr4q2UYMxCoBdnabdh9rvgVBfBeqyBpCBswVUBA3Lm
NNNFOD/8Ta8XngZD6JvF7BHXtnYrycXEWQK/sL3x3FLlkX6983fDjlpRHps7hPSlPNejRSfpZuCw
o2UNrgxv7YWNq0YyC70rDZdBx+YXnGxzinhzylizZ9xiDgce+9xgbCMqiSvIWZi7lvI+ZE6C47Rn
OYdOGluXFIr7IX4+G6sNUGE3285MSCIWHjv1heYvDFCaeI5LEllrCjyTpUBb2jp8szpArBf/Su2f
gLlwUo9j2xqnoumQlGPQYjdqo4dQB6mO7ghz3fWkMQDQ5uCwVaxvwrOc4iK8Cq1LfWCkJ5IfUuTS
OxJBujhBVSjYji7eKa1vi2ojDYu4tng7jESLRZnU8blT8kkmNfkVyzX0rJMPcUAUarB4g1RcvdW4
0vRRmJkArq2q5B1t3IZ46xXN4t+zJo45CSNz0penoEJrPOAqqShKrBCdn+0zzI9p51NJN/uVSB1e
Q7dsY9mqy9l3ZR3pPDGKJH+8B9vMepLBelzAuEnee01Aw1xT/TmT168sHbZhDcpZNmp28yhPwZCO
1rmYFI/5rNqrRJHqc+xhPexoGrGNnHCKG966XlkYww2O/tyeCz/Ff4g/bPMvtkmqkGsAcZeP/WQj
J4ACJ9jndXGASEUUO0Mvx9HggHjatheofOx8xWkrRvqyYA9G6bE3qr3CLIrmyQ//ms8CrU/XqBPj
Fe2DP6T51nrIct1GFOoxyLhI146HkY3fjApayRSUK+euIv62pcqDqsAjmcGJEKeg9efU52EFHK6o
2IevBC0ovIKQ9UGknuLbUnpMl818w1qSEqUBX3v5nexmj8lgRov5UqH15plYI2AdpvwRHNkXzME8
zKh1ow8cn9/C6hm+vulV0LtcKQEyyvAPeIlkuvdzfbiRh1CnrQat6szUzZ22bCRVbaNXuAlbm/ZF
NU2jeL9vxAgqBHh7Q3rb4d+KVPQzuuZFC4YCQ+p5Dx1fNzHg7svlBOVrObQIJPRmySif/Vo3wO1n
ooR6bjllCZ9KsNCYfifeyyhsSdxbFpNjkpDoZ4OiTXXXSg04OMeUg+6vFO3i2G8VnWMhuM8nXMth
6eG6AHCXlrud/hgTK3yD0MGWdaQwP+2zO0xAa/qRaXIA5IGYqrRHKXG4NPFpYIqEoonKBUG8bgxc
PFh82NVWOFStoxpqw4YR38K0+mzPZ5Ywvs5EM25OzXWkod9kWtBrGc4QJjtfxiVnyCKXZFIIKOPa
3sPlq3+p3JPSUBrhz5XYJyAnPxbs9HnRdaov3goxkjpzP1H8+YLkeFEBo095M/S45EbkSa+ixhOD
A7Y4FvxGaP0eOeBt4zkiMWu1K+CDGMpKDzwj+1m18UndplAEu0w0thXDBZ+Vic4R+OoXP4T5wDBO
x2ZXHYM9lk+K3vauw/dl3QFdngBGlgWfBsGMpoYopsRbHEkolXYloLDBEbqmnGikvdEjydANCli7
1XCIFGbZ5TO0upMywKe596kPFRBYXvSVjORFFrb13tkKnjsT7wNW9705YCNii+ciqLpTqSQmnhcj
jaI3awqQAWplEG4VNlF6tPOyNNBTO0G88w/cVsuwRstzp+QTHvdVwytFh/bWS+1osDAPnJWqR2KQ
34sySFPSZLjnfXNYg9/s3CZnSWp+NL60QRF5QwThqyRRfV+iEn8lB78ObFodpDZiB5/MZ/q5kuZm
wGTh33xMTNaxN0nCeCP8P1jvF912OZD0Bud1x3i2dqvKO0unPygr+LYfLL/7Q3SM2/QB3dYz5udZ
/oNN3Ceoj5SCHPvnU2Hs+tUdDynjtpWRx/HaOl3GPX1i4PHQzF5b0w9bhdL5BTvCqbtPp2BDeXgE
uSuheVBw5eYFRWHtpysodZ66q3mZtAvIPRqIrTPy8v7ipimkUIGKoh16IPDJeaREXtr9GL58iH/T
OUdkMkTkp8YnPtrz9AqIy6nAc20FxMNn8Wa/J1j93nWbIKdOI3LBnnzizus+Im/YaCmz32F/vmlZ
SCaUiJuO+w4vwwl8TMcpv+HdLB7BM+87Nwexbwb1UT9V2wD6XrSHqIFIek1GH7m08cGezSZ2C10m
ER3LRj+3o0Oxr1Ox3K6ys2muUH2Gb2mIgODg6LuR7JQIdXnB6geQr+9mwavuEwTLopTbfikBYN4D
cc93f9GFWIz7+tJmsxrAWu1QbmQjKmOtBF4AF007tCg66wWOHkCS8AY9Qfw2kmzIQKP5dQQZbhjC
SiyVxz3hfw099OvtM/FX2H5Lyh9fjtXjYdYNwmMw9LB8jrMSefxXBvJCzJhg6kF1wx0rGBZRQ9as
4uV81ZOiqWUeG0CaO0phskxwP5axFuNvdYG/RvIwh//P37yonrfRAcElxKrlsUC6ItY52KzhxIvm
okGbCiW/3fG4dvWQtOFA0AwCsnQkE80sEVHtzz8nsOfmfnuCw6b7Q6wbLys672uqAt5z5uWfBU2Z
CblK/dHu8NAy/aRZuSTMa3m/JiX9JEoGDRQ1qXpgGdTP1IIhye5Rejy6p/u6fZy25HGPdPCOcjp1
ZOkbMJb5TCA1FPC7XwzqpsneJ5XOWtoO030CYj2+igNV0XB/DrLn38Jp6SKyC9RWtFnGDEw15cqG
CNat5Yyz3Y5lRxObgKcO9YA+i617w5+j0ILpW8O0w7LeuqflVOkXE+LshcPDpTKzBwRYe5nXApXC
XUekxqmYwqjNCnkM+f6Vqu1otsvedwC5aXh9cvlzKcBlPrnALMQs6rmwIHAo2Js1b+dEXz+5clSc
+XjPEDLEBxfi5BFP9HQsoKWuOEVo56KWd49vzoyFjPrPkJ6y+4augXoRQD4slP0ScdauGAjigLiB
1gvOqOl58oAEIr05Hraa7ElSjMH1yaiq7G6lEyqlX06mBAXnVPVQ79ESLZNpVCepIwlk6Q0kFmWL
v+8a4vt27EOhT7SlCTIzYqep4XUaKpaPyVupxYYYq7/5KycWgV377tj5uFIm4+S0yV7jf1Ueh9/H
zJGMMOBAkggLIOIjjEUaYsnqk0xWtUasstpK2T1Bdnpqf+6sIOuks9E29ovU2ApGzEqp71Gp5gBr
lg0dhuZ6mSLQNDKelu+47WxiyX8p5sjTC8kOKPuEsp0W20/igDQ4JnoJFyoCSNz/Slwsn96Q89UQ
NKhh+zSrvz292aDtKtpOv3O66CzI+DdCruetS5aAr4+Lm+kEKw3u0Ix5GegHhAfMTjc01yo7vlA3
LRYlNFiI31jojGTbzhXDS7viP1wi5mSnzkj6VOATWehiHsiTUXyuWmFDElnsoJCic4ZMfDBcKxzk
YqS3dGe5xr1U/Rnw6dtv/uTMiw5/qb8+wDJzsBDkJNb7uCcHIGm3MbJAA7fZViOYc16r0Yr4b7bm
lZ9pMhVAJ9Q9BhtG/OHs3/eleHKNFLV+4HKoGz0DJ+B7aSo1IBnoOGnsYZEvK+sIORbf8BTUWYbf
Ow8WLzQoFQ2xtcIFZGIJEc6Y1KmLK7ijkmgdw4b1Gt2LkBaPNNox3ZrumgWyJl9KKGnnRWibIwgh
X/OJewDo8R3PNRmTs+YTsUyjoyQGdTVNi7XCD5l9B7NnWHZDb/ypF1imIXSpPiT7bXXxTMmocHFa
c5EtWuKcGj+UHCdPId4LfMLlEOSL25ZT+QkpNjw0feiGPQecdzmh6SSABfkDg7uSaJlWhpSzP+ME
mN4GRMuwfozjphqOEJDf/662i3Xgo4Cvk5iUIH+5CLKARZUdxsMpwPk598S9rfOSQSfzpif5hSXk
iRHBtzo6FCHaqc28tj9kZrK46ZX919ncpgLIz4kw9vr6Aqm2V3FTmyhj7lDzx82JaJ1Le0hWYHqF
GfW3TLGTlG1WojJiIAvRQe3wQhDQBq8dPpIKsV+B2DTdfaCQDJrP94SVNOffn9hk5hzdm4H4SvFV
Vohg9oJy/kadNQJi1OA+yFwN2jT93zOquaqmwwh0zlQfIKyOjCQq09Zxur/cLcZpupTe/w5tZ6pb
QxkDAvvTPL57u0HKvLguCeFDoTKwSPbCM/xb5S08Z2MLpaoooBpRH1kntA4vtTLjuv7WqekXpLTQ
h3/uqB/UyjPMpjrD0yNcsEJ++nrbsfG+GVLKdRwhAJtJ1xToAL+a2AupFt6jT2M5nQO8urGUfu18
5xlilqEy4Nhe+A/a2neC6eKvZrtFFrag6xU2+B6JI5waCI4H6lpkBVOtmCt9QDqXTmhzBFrdIcwd
pGH/rw9XnyqD87j0tXwFbmsYHBDKA7JNm8s0YtsMdps52GObFh8QIS9GWLt48V+vOSl0SvTFr+mz
VzhrgoDuVbGy7htat/+nViiQm0v/E0eVw7PxNKJ6PRcEQZIKBWEln37xWJV9j/ReGv+/2OcYYSIm
pYpEy2XfuYgugN97y1Gr9sz+gBXO/NYYEa+xReXah8HBVh8k75E9VJLXAB6LBI4Z6iL5aWaytdCe
zJM21XshuuRvMr2yLEaLmj48VS53nrtce9Wz9rKe07DtlDcmD8/WwjHwI/N08DLKaLnN1Qb1P2z3
fsyWnqRy1X2noQsSpE8vt8z8ipGitS9K8/lSFJC8x5xlQk25OeDVAIIZR43E0De50zmuj108i7ec
XWt1g+6zqWnkjtqs9ef+ChJsH+1p4y5hvWwvgb46R6aGUzfu/uEDgkUbm0zosUlympou7e0BUGYh
xIvK7PuyMTS8axemlirkAaBGVIoHh6cfTX5/gTMkEisFjaLaxxzS7cxbC27nxB/PDCVIuuqJz1ef
8nOmg3Mnl4sFydm+ELHQeglfZbVSos1QpxEtoNyNZvP4JmD99lG/Y63mAWf7kmwy5skF5c7nAl6b
GVU0VH4pd20SjpQqiLW741tyK/9QfqZQD2E+dqXl25m6oOf6jN9scUcK7ow3SRmrOFYOE31jdwnI
M0WdLkhVo8AMU+VBbU1Is0n4p4M93XCk1wMqYd2tkcGtEdRxMdhWOj83HOy76S+vJkaBz1X/DDyI
3V/+0Q6av+IaZbpKQTqYlSkMRQsyzYsk3SBPpCleLEHeyEpFAQhLwCyJgCkqmLpBRk9zQtuPIONE
JjluTyFlzVN5z5fBTSfnxkM6RY3LBMaGmed0CNOe4i/XAj7yVIBL5YA9pcfHZlcCVh34TzkrcEHc
fdLqU519NaddPxZCTvLpekcHxPKdNfCkscXpGWqMPXgChYlVi7TZrqdlIDKyvYtVbs762u7lhghQ
4rzRk8ol+BUoN+nRIeIsu9Ahxkf8qk4DjoUf6YKEP9z0J5NY/Wni4LkpUnUMuI3H/wYTpR5dpjVU
/neKrgzqKdxIrqyOGYdgfqglGvjvmVq0eTzT3Iso1MfLhaEvmeMgwQjx6WdvN+kSfy/xTLEx9dUI
MAEHQCsYyxhefEgqEcKvRcpAXGAvV0cLe3fexPUZHQrr4iOjiNpajOjoR9/qCksXmnUkeP34tkLC
pilpihvsdpc6AHtv4EWMg5UdUgEKOOb0U+P4gJ2L8b5/fxxPTsDv++1aQ5bXI9dw0NlSUamW7V28
0E5VWd8G0ptL884PvyQzUL4nh1vDEj4ie9AjGDUIOFTCP5o98VzJfAc7YvRO+GVZ46V+xOj2+GJP
yOuUscnZ58dYxAI6PyKfc4VIUXT2in7mgru1OZFIHTItQCi6HuF3FDet1UXzB4X5LMMtb5uMPsNP
JE+GAK83Cx6rr9YGyee6wI/w6odlYMmlVf8jxA9PAx0ZBvaHhMIr9k0u6UIB5bF1+mbjNqNmGkK6
R26hQE8b+iwnINURSLjtE4ggFEBgPKhTFtc6ZIuvuRyUiVevtl2JcrQMJKBj2lU+rboUxdo0fbhX
gJJfVlE6aJLeMTbQjbE1XzXhcHPS8BGaL/k5nhBw0y7k+ZulwyQgbUHI1NviR67KTaSfLnX+cjaM
qEaayQyni4nd+YdxrsOCNk3v3Apl57xhUq6DgUHismIFozXWOm2X1z3ECAe8jhy4SjQgyQI6f7zS
UG0fL6RifpY0SNSA1j0WcFmYlkaOr7JX0PshmDzgAXqNhfdmDM642U4+voVTl33QF/eGJSSUfioR
MinssQ68UJJyLiMn1pSwTOaGO8dcrwKfI1IWCJ/Cf9xtnvX6AAEKO1nbTkIHS1Cd/IiQlHb0QasX
k12Il6HiBY3u9Tf+uuIKVR+2eBq37J4bUTfz5xOAR07AmHdUYbQMG5yjJaCu4/WluWeX6pqPCyt1
QL7WpilSAG+A4A1cQjY7p3apb8gTFWmZcLtzcfh/bT7Pan9pOuRj2XBt10fgNoM/LrNKUQVb8LI8
ACvkDQ/TpIhmEENnQ3YzQCEYLkcxfhJDc9pgO4Se6sjr2bvNtkncBRytnA7y6JKSmfuR974QPuQr
84z3szztwQPFnsE4Yaz0U9IJcEqMN5QsPEL+VclfQp2kr7kdLikEhaiPSUO5muJkTZNT60gGohkK
BSoFwGP6o5jMp7HvxldGDrT1XZWthY6F2V3I/UwSQhxE7f3N6U+iNVtpNRc8NNiWUWogBZKrjnr0
MeTis+9l4e0hcTOxsm13wrNnR6/UDuJYnojQVphlgrDAILZX1rV0IUWZzLZ8JmRo40IDSLl35Wz6
1sOnUuy8VetpGYC2oz7aZz2/x+4tjhTTfw0ujTVd+1aaJjWf3sKi0PReRXVU6TvzD9sW/44b62d7
PjS1zykuVbZu9aidPvfh1kcnpNPT1KrDbKyon1y981iRzY+mabrckB8hV1zFRNhuwLT4wMLIBtdc
Hz1fMDQakQqNPuuAPHQoNhYmRnwBdASOf6k5rL5JjwnLGONe6HYmsu61Jv/WX9AebdybEC/21kRw
JfobJx+TuidJYQlzR21JszF+F4R/TvqrI7FwnHWEs4na0MhDkNhEw7U5+/OCJdquTjdKoQyt+b+9
UdzOKRnEXEpoD6MZfd0c2/QCBdXJBzQh6DMfPhe9pqKW9WOcwvEOg6fLtlZNEcJf2Cx+F2Ae0OWI
Kmx39Zu4Gt404gMPZu72orT32D2Qkb94ay1P5lEHVGlanYCpvZp48TfFzewCF0+uFRon2lILlJi/
boo5psgzhJAUu80a9ciOO6wQp8lqlfbohiCO8XDSfCpFVySLNXXzGo52SOPIBkZykIN2dQc3mBvK
KL7xDpbDxCi9RBWsT0g+ToyLj5LIUAF/C4kEG04hGNFjvBrVeVegz8+3rocbp64HLCHAi6hIjPNu
Dd/elCkle5ayg5NiLqiAJgC7zZccEVLgRE4hSvZU4vxwaKgKwBLRg7L2sIWA6KXQLeWXttndMhAD
0x/InZa0f+6Ip4Fci+fGeHgNJiTqO4IveIV9G8j4S0CtryMd+R35avf3ddF0iC0WPDv2pKm7DLmF
XbIr2t9CQKlAiSX1bnnVZ3ub1atCouZJA1ysBONK+Ma1K+2K8D+BYcET5jPZO7Mu99mVNWTZRtvj
n1MRkmPgMeDvvpOrK/SjL0Rc56Oc85jzDHELfG7t+uGxLgQ+wBt2R2/s6UrW607o1b3eKdaVCmRG
JfpDsKxJU0jujvuHUTvhP1e4y/RvuOoR+S4FSEpgqPkqs+2/UKVo137XSKI3667/gvSnSUgrH4cv
MRdMKkYJmZPxWxAAoSIqRYVoqitRU+xGuRkjdr/41RFMGZN5S5InnFK7UYVRFmT4Y0dpyala3Dyg
zNAAAU+7elRbAZLetVspMmYC1ZsCrYW2o/KyqIIhr25E8yzAfWkW+N6eYuheEG4C7mqp/eMIhffL
4X+tI1RkKSlPEoDU2CibtuMslv1i2gNSz4BzLC6Et7t6GhJrk2DdsGilu27Zhd0uvwsMGjMSiboJ
DCaEDiYBb/tBvKyjwgaKsaw10yRXDRW77jjIA5JFOzSSikSABL4YJkU8/U1nkphKCZLd1K+OLRiw
utFqocgLyIwbusvWdivBvwpHFJwd67tXqmIT3ZWGuR2TtB/wHBCLNGSoiWI8Mu93rbmXKwoyuykw
3I+CJpT1hxDQnaVo+UMRvjr8UWh6H9w86wA2iygUzAIkAqeGmneTMLpF1NM0+KIC0OQ0XQmxlDN6
d4XV79Xlj8ZJCncliv2/cnalk+tUziWZAN2qnay8alSSfC6NnMyf0cc32GmUDE9TZ6aVqofr/1BX
g3pVQO+HzwpMh36zL/WDqcOi8c9I0O9zuRi073XTmSiRkYNS68qy/Q8Q6z9mg4tP+0xeFGO6FMJm
+vb9gvy+ZGPNU/unOWYGmZvdlWfEe9RTAnmSqww8z+tqIz+KeFMcFFLfsmseyrn9Twfz//jse4vI
+IFCKhZ0RM4e5K/thU+NFOUgw/2xs3UH6V3NNmowMa6ciw2Deiz931LJwl/YDYHdZYKZYLfD/EMl
tyC8UagnmBUAgGMnufwIElqfBXwAackfuBLIOrr+XD49e/trx75VfpodDIAlsIGz+QUdGOXyG9zU
ODLCvHSjLDqxf2hsN0E8JVSm5wE/zKhQC75V6v7MhG3AQBXAgGwwBIV6dBlP5UYAMeBKBf1aiDxO
dAHGlIHFa6Ezn5m3a0k+c/MAEAjLS9uugc5PRmhLX8CuUGNx3/5hzVvpcKmam7TDH8dHcgkkYWS9
2qr28DhtfSyVsNwgY7r2V1dGvUcWwRQoh46sLCYqWWC3uw1hgOEKjOyecOg0d/eOZPMAXg+ww9oX
RKCYHe8nm97IRLLt11yHWz8UILXh0wA6/SpcZGpyhtZA++Twk2nbIzemZRb3ePv762rxM398/nCf
kN729riLyTbG07IICIPVg5WPlrUYRcwBOD3PIfJD9h9+WiJxjXUDgJRd9MqGyu8TmfIVpJMZNYqV
47Rmn+LxtakOotrs5sWixrbPpdw9AE1d29KwWfBjNaMf6DATkzaERu6TndhtkLWBFwVX6Kn9YfIo
RivXtLQRGCW209QBadC/UdFrg2NFtBIfqPUjWBL2WDkNCDg8sWsR4JSx1CQvaj+Pps6vyqbhOksf
r0Yi31uTg2VQsdnSwntiSjxKNxTixfwNMwoIuuCd9dSHCtgAilkNP7fQzqBnMLJhATVckRhummSW
rTthJgbsDQOVfYyKjrxNQKvdxZFviZuIV1uvc0D95QZ0U9YOTMY3JWkT3AeLct0dDydjPesgCCP4
5xsG06KuaD1oAiU+EFSZ+gpanb23WRbxiKtEkkV7PBXD9SX7D05/TyB110f89k6tbvSFk6hbRuMQ
asuFONprhjL+CibGlHZc+4IoyZASQ3vSygSbIXz8x/CxcD92dbeAA9qtHwhcZ9qKyVWyJ73KKDfR
Tx6Voxl+9NvtDtKL8YDgb8AycBUjwaMo9m6ILWrHk5vxCbnwDv1N+glh0gf+Oif4ms11cDw84MSr
AUYfO9r4H3hP8iy7EFdpkC9hppBFbJbs9J37dKhc4F7oMea406aYdR97mZCmbVmvXN+juasRQK0+
Ko6jbz3pTuSJn5KXYG3EZ48uD7AtAeZFmMY/De01jPCXG6R15eNojnXsXZaGiHka+enpiVV5ndDU
vkk5G9/vC28pVlKpti4yZUquDMyQhR/e6WBDhkLWSk4mLMhs+lVRh223PcPs9j2mckvw5DQc0KMB
GmFK4Wcw4KVXqqwtqZyNLWp1hoGgmuc0zYAaH9cuWpDcG5usJ4i1XTwADwGXy4UmVARhYpqQ3CF0
wk70jJNPFmiJfIUdKTVOohq3U6YHQjx5/3LOKCC0XkNc1bNfxr6lwTDBB1AKviIrld+hdLAAMQjt
rEvK7v7QPcjFyw9HvG23PbN0RI353O33MTdb0XgTSGgDA+jXenjxigcBK9lV2Fu6/ha45xdO9OO2
4iQh1kc5EfdYhbTWiluD5dFxbz/yiU7WIy1iJPBXk585TYji+1ODNeR2OHfstidR2DclLPsW/GRd
MKTluVBSCyD5jbI5n5LZFljZ6TdHom1UnYvs/6CHLfl2UskeUUmU5xhprGlmyZ8RZq9S59gFhgVU
N0I0297nIKwLzqyR4E2cn7AtmFMrzj69N8sXk6jqvhj6H5phe1MhCFYlmGLrpdLVVt2buHePH/3V
ni0ucpV7eAU5OqAr36guesbA4/xXTg6zg4werOyU4/NNrX0Bf2yvQw9CKpf42ZF1P4GrMnv3cv6W
8Ehvlc0f/JekpODYKW0YpqBP75zitLymyTu20gtdzd2jjX52PLnswfEq91SpdkOMMsfVtg2l0Tbw
Xzmv6XtDRAyL7vbFIZ2azfmrs9X2oOAslYswYvU/UcFHnDlSJ/fmBdV/gluaiWtptCDASLVWWJI6
Up7d/2JIKufx3A4446termLdB77eG1VduOlVs/EdDslMWqryd5OwqYgSSOtL8Y1703twH3v3K+YN
42umL1o1p3NbKWyLb6KR+Dpl+oSepAdYVDInDzkUV0d0rB01iisnDh6C5pUA4srtULXVpJQfiwBH
z5TPHqH3CDTXOiZzOXGPR+A3wmDA+OJgle86IWjemvkE1T5P0saZMrW/V8TR19fGdSz10EX4ZkDa
8GHegnCGWlWrHYKVcMg7IioiYXp0bNQtCZ+uzFwMkZJJhSdYV1OAakYWUFov1WohSuI88MEdeuJU
9nqLS4K7m+qsfxB2GmyrllEnM/khv5BS6JxAZIjhY0felhkYMKnL0P8Tjxqa0v0jQHPR71JEE/+x
Z/5coqEm63SMlgAf43PQWHQoBEaXtWFxbRZO9RrD6JqamxVkmp4yUxJ/8v9LjWD3VgjiD91dQ5T9
HpQgYHrdl8CulTB0wsNeaqaM4f1apmW3RGz5eQ87UPxJte6SyzQlYfu4xRpJxN/WmD463xyMPhhS
F3f2Qo/AU3rIz3Qb+LKirTQCOT9UShXQedH+rHIy2EE9YitNrTLiI5NHCPAzP2y2SwbQSyQdaI6I
asvtYcxDcoi09YEd3l46PYq95a3qx5Sgz8pkafxGQSHS8sZX17kvN6CuoOodgXNNZ3PLAjJqvvfJ
vpGbD9SZ4IpLNpz5DZDKBsjCPr1z6fZpR4OadCEKb+dhSoVsRMfij2+fhkIx3uo3y6giFW8/bN3p
vjOAEDn5oAZuqF5N3czJIiVMiClgjBwhMr1te2W/8C2KsipZ6pR3z5JMInAdpkX9Bg8Z3HIb0x9g
OVPzR4xosgUF0rGfXTr0bq2gopkqUEwhUmBMuRzDOsXfLcXyW1IYnBLJ5vXYLW44q5kibfXBnMmW
p8NHUpircoHoD3AgExbw4DMc35amd/SjM34x1OBsl12/aOTYF3UAOEV1hh0VVQdTF02GED/EC3xW
Iusw01VGicrrGEi6e4Hs17JOJ7cb2afHECNSgEILed+fhx1m9jmea34nIuqZGVjC7HzHIJkmP8f9
3M3ZhKXyLtiCJCoUfrRDc6qsRg25jRWDtKOEDaHBayKp+kcYpLEXfQuTWhmnAywghNn2oj/4mWc9
YUfJ6g52lTW19LDIyeT33pOTVGeZenXvbl3ibl1b606puGVc0FOOPuTzyaz0dKq3poEn0eKzBLxz
I9zVUbfEQonrzRaT+Z7HAOEnkwL5KfPm2oScRIfn8X6a2Jh2NlEkVn8TtvcTMkyIewddWvsIPQ5T
GHyXiTh79AsDk95imeJ/GBvdDZ7qogNJyS4qEVIVWWJo4n5V3aH4GPC9mL/QmxZSg2IxzN1M5udD
OBiGLS2xqjMIggM28Qo6vpo37Ks3dxlpJ/+9DkwKQohPuZ6bJtFyZCwsbmSz+ZEiC+Tb4JTa1IEh
rTJU/e8Q8zPxRi/eYPkGvZg5lQecVMNyVsHFIYmccthzhjIL2sroE9SnEPIsuyC1MlQoCqZYpklB
R926ujSXzSrAkRXnFYMI8YGZzXJx7kyYTzqihlw3yOIcd7o5WlEYtJglkT+I/UcfcNZ0XOQ0i/Uk
KxMtZCdvs7xzy2sRrWcxl9Fi7equVinmdz2bMfH1BhbyIUXXyzxm7Q6YMfh4OQxSTIxtD2wzOiJm
TfCwHur11eHg+8lvqazH9LylhUHIoVoO7Yx3V7fH8lcedPVlDiUUOZ5nFUPWHnpfIDGtA3rutl8I
zskOBqU7cGG5L8vWxyhphDTAsKA5NCW78uyRo+KStXJRF7+ZZvDYiNGC4niaDMW5U2204DT+XD2m
CVI13hjUAqpYPkZQmTFkgXuieh8S9GJ5HKCss/LqFvgoR2q8e0thtN41SyPai6fMBEA2fmYSEYGO
HVGuAjqkKv7EpO+E7CHEcua9zy+lv3euJeIiCB9CRigOoOdGJihfIqdVPFJ+eJDB92mDe0TGtgDG
K5NKqcyd5lSWx3g0ElcNyeZuu5DCpwEjDIC/uBcgsMolZkqYiYu1z3B/0PkrPXLx//uJ5pyPNBLb
9wya52kfk9dYdVODtv14brpWIoZu+Ryha6WSe9Vvgyv5qB97AKonisn3EVPDP2b/LvyuVtpp9rVk
oQU/PCQYK3N94sLkvQhLUJH2jyXTxQ5ZZlZj0YFYOnKQuy3nv1GSwajzc0DK2zNfc2zCan8f7rm5
ZmEQX5wA2xuyJa+Yi6hkiDYbb62ycCM0BnNJGwoiZoau2T38BofPygaBStdY2JwgfFGBE++kmmx+
3JwzoOBKS3NguGu/KsNMpU/oENNykZGL8S4p2a8Y+JHDx2IkdaH7Iz9SiXmzkeAtRfUStwqF4KQD
ssMEuhOtkbNvInYcnhwed3tE5m2FY/FmlRt39eCo1il3o7ksLPVzlAKOjCg0LgRn/QPNq9ELrjK/
s68+AmKZcAKLRW4opKHFaW/8NkgqoaR4kD7+Gzk2s2xJWaDBu51m2yUIcuCC+ENQeLGzYXqSWP84
wYVFvVGtD2IGGBzpsuf2o4Oe4R2LXMHOaJnPFzO7Ix1EL0A9wbenfw1jKDUTe3RkC/dbQ3SRsuKu
v6jdPpJnQw6oweNMGbyDKqA8gPMxaEG4+08yqeagdgloUg3zeVY2lSYBtsALyGBLRE0EIrCiaGYV
lC5IL8OP3cceALN97YCJyMLaS5x9zuEUr2IAsjET2vEnz9zQW/KdnRjsE9jTPeOCmvM9i7UWzqkg
8bdesp7quRfiqIb1hkrmgtqZ+a3skrQHzVTLDcHeVmNsTiNpS4o+4x1duir3SdtxZklf5f2+WIn6
4m2g9jZYTEUdzlpxUOr1/hp6p6jCMcLQaq5vd1jpKdFGoLDOw3LiGW8+gDCi99DWiux+T1fpizYj
EpO94lWAGIe25xxQw3MiWgGKJm8TWg8Q40g3m8oP7X6wkzc/NYpuTSvMbOVGaUHuflEIm7jzXXTD
YzdCYwibwFg6PxTyPCzalAREvxnBDXD8ARm9SwcNU+U54PL0k5A2T2RecI+dD6B0MVtUcc6dmRBK
H9J1yqka2H1Qzu+XXcowFd1cIvmHJ3031GDR1Bfvyx4HAV0+1BnB6jF7dtSu3RJlD7lxmDtqoiSG
rlw97ovHBLy0c37P9oLINurz6e2+DZ+Pmg1YhrGogxDK3EBKix6sYSgrHZ3roEdhblOfWl5e8DPV
ETHgqKw5Rirs9NZs6nNtjdpvImxOr/hXwTThwwp8XimcM77CrkiW0I+7VL88qjNTo/853tFmcJPi
HWld5evnO+WyDU2xLt0NEfq/kTdijMe8eAx1pUZ5oVCnADOnJKsgBxrg2KFPZ+EHnIVWxPSbRfK1
KiDJiQf/C35XTLEgBXR2oZZkUJg14WXrzmukVCqoOzwTYQlum7TrRU/1rPvMKL/IxBG+jAzY+04/
jGWar3R6C0s9j5hXyGulP1R3lohWa3TDT9zhT5QtMV2mP5JqBPRJ8TKvpGXjdM0z7k3bevkTNzbk
Cd0XQ6qh9nNuK144/1lJtEosUbPbi8ZECFobasd24HB0rDwqPzx8oT5QQHOKy1JqMNG+luadbjIG
tWvMl41CUydgFAqOpszvlY5rTnKSG1enuQjejHrVWe7aKqHwt74mDdF1PPkRQi4/zbuSITt3J5HP
yOdiO/FiFcFMMUS0irE+ztWotzPMH33P1OtYRh9p2edIxbRpmlIYFdQfKzfHlmQOLuNdvrKNAfls
ZE8e6C9y/899pbOxUppF0hlbNLyXzBDy2POwMUH+wxqCVt2m9NunERwZmAg9bxZCdk80xI7qlLq7
wd7nldkG0Z4P//IA/mFvr1cdNyYrp1MlQrm0Zwez1hbVZPyugAFOgJDWXtHlSCFpMHqrCeIhTlfg
CKLJAYwkAxRbakjwFEC59fli20/jxfOKIpeTJub2TkbT728GV7718NIW19Jvk5adY1fZj86CYTgD
ZzMzujqrnCyfb1cyc3cXQ2PDZdp9naA6Iyq77WTimLcMR217DsdW7zdDihDfLQVY+7pGc1VfVZne
1LezboH79Ou5LtDHA5hTHdHTxHKcZAQWHph3lMX4xCOb0rR9Zoad5yVb0Qh/P0GFvIWP9HPVRU8C
15ycTu8kIWUMjUxpc1X+rr2LgFHXY3plhL98bqPaxFlcpxq7EEkwLdUP3rYqKrEHRm66dO3PdK3M
xP1SEQ7XdwQCorHzdciMphVzuFyqTrscrs75GuJbk4rmJlV2cIqgHS8w7eRJ2ekNOt6mUp2/hmI1
7XDEurojJHTbv1x33i0KixUVLHSApe9yiVIQnw3g8sCgWXUPpeJHDP0CrYbH4xzDy4DQLb76YV9g
KlxiAJ2YYGCSYtQxEIvXba6FKH3ULMll0S7O7pauUB4XIgiDIYD8IKpFuiIWBk3ptlQ7EgQyytlZ
bxajbcWch22NwJshd2cP4PnrshLMwNSV6bgU1ruj82Di0um5T6QgvkLtu/dfwEdGs3XLsI9Rzf6O
Xwu53cslz8WOJ9dFObADTWJAz0n1WsJQosbt1izKkBHpbmjkgaRdHqI7jD7J6n5URIE7dyci6SmW
LaTCDNK9iaXLkO3n9hDoykLGhkhr4UYBhk90/sWPd8GXdVXNvKPfVHI2L82h6KgVgYHND+FpsMHB
GhInfkfgGNBdX2GuNI7iEWdBICkR/GuiWHNu984R5kN1A9gorZ5MZK5cHiSfr1p1/8II923fBS7i
KaLHKwSrkvP7MeUm/s/EwKh4d2HnnkVUS52Je7yw4aSD0dpeQ/UMYBGlGK9vIEtTUsbLkM8cmCuq
LTtBf24sv+/5g3e+D4T3YycCGBTwezTk6ZEC3K2DkNA7r/BpKUHUqzs0w3lJbGfYCRN3oclYl045
cdFdT/t40WhCn4Abr8vNKB3GYP5+/JokWfigYz5OWVpaMT9vMxM6+youb2eUm6lUUTfo9Mu4F7nE
Jx6+/N+20WaRu1oGVwyXzAcjMrCJ8Qn6blIgWHaHUnlzVC4NfK/e1AR0g6H1nNQnlG+ay7925ugl
w0S97dOAfOJZCu1oKOyobgav62p+q8XJxBN4uG/e89icmS6x4bV6iOgZYJbLhW+a+P1MipHc9mvX
Gdfq05DYQh7JWvhH+FP5kkr/r01AIaQa0xHEBy6mHp2YYu9ggQBOydMjHUyl9OzHXHk1fib9rlVG
ibgoK/OcYIfj2qKiN+fG02fqC+fbR7JVmgAFDdvKkMosXRi+TMvplX4l5sbRqg3pgNNaMaLUwPI9
Uj3KRMwf3srsWQnpXXvoLutmGLHBTojf/N8JS1Wq2DTtP+yQ37pd7VmrfMUgKMLquI4/VYoHj18U
m5iCxM0UP50egzOucRrWOmyiWakdLAn/zJZqHRYlJRnIVBqGG7c/fmqAgdaYR751yA4cN/gDwBvg
CsdSGyUDXFWOCVB8AshKVoj6HSayrEwsUPCNv2/9GdzgLgPQJk5h54UkRYsHCru2j/B8dw/RoffH
4ZcWKcxx0fQAKaVTx8hPK4uD259QyDMTiCpovmYwsPjOzzQ7tPNp4562EiCgX4/i5Nvg3PZQgXUq
V/HeXK2A3EweSTMGYm1UTwFFQZavz2hwAjxvQHXuUGa71i92SrL6Y3EGqqPd5o7XOeCNGKoHoHKh
v0oE0bV2l/a13rlojuHKzmG9VdZ4/O58zry0IRULkP6dyMpUO1fymGqa3pQvqR+6kOaoVxHYIWRe
Ikn4S9Xg59/u5U49DgFx1MtzaYL+96y5P+BczcD8vd6amkAS1jeAEb303u81qcsXw1c5nGXiSDwM
D9/kK/7ANCXR55zEp33JYEd3zxLimo2K0biwYSCXq1YWWZ3dIT5/C/Uo5rDL2j0qGsKlCWU66QKd
JM65vAHvMM38V/Dv8ooSArAgqVSZYf55pM1J46yvKxrZWz+Q70zLdomlBxwBc0uYLPlSydxetxis
C1KpLznrTCo7kLf2+LBkpoDMcWpIxdTbSpAoIqZna4X1VQ8sZ6sS328s6sR6I3JO7Z+Vrx5KSXQs
7lld6KANcYS2RA+M8A3NH0QYi+6Gc0UJ79z6RTNs5C0lVlu/l9PiIz4nUrrtTAUW9jvx9Le3y165
LKwGEEclIiPtlXGCI1ZHTWQ1ZMsdxRpVXZ7wAZiDn1TxOdaPnGazyZbyYJ/HJuahBq0uGwcKEWAe
zYDOkNP1/j1fDylRjpX+diQ/xqzV1O3MezBrnwRxjGT5X8EqKnrIdhk3Lc+eMTqWmPydr5pvn1fu
vWsXohXdiiwyT7MTLuvmq0cGbCYWYz8Lkipi+fw3SSaML8iFdXcA6azxw0oews0AoY+97tcxEIcQ
cin6geFhnTnN7ARwpf+JEtcL7dLDH7XhDzN6FQekDQg+X0bZp1e7OvTCPfwMXU/y0Yn6qK/R2cb0
PwHDoxlTEScFkT0JzZHpg2D4Jr5nQ6UbckfX/ejy28AfgnXyMwprmJZhKRXHei0aWDbN6NbcbGvM
0n3wGOx1N/lH1S6y67a4SpbnilxvPq8ZAgR3pKkUbruyms49FaIY+hIxP2ALOdI25psKknUrsjHN
3bdq6fkTQWcYaz34CsJJMFlPL06uAaVl3Y8a+rbIP1/p6q7upmWyQRiEZ32FcQJWdpGjOs5Rl7R+
/AxcMA43w2nqg9DPLNjJLkhohIg8wmNZP52Ktp5rpPxVV92fyS7iBBr7mXsYgy7n2DLLcB4728Go
3CMNUfpLY0jlV4JQufXtkSGUfcd2/laFkGw1IA85HdZDWA/gmwg/6z2wIL1bwTe+dB6z9zOdLgv5
b7FT8p1w0ev/yU/rSzEJkEfHh3X6ikY1vSdg/2e1i0Avam53/TGZ+VAfhI1nQo9LDHEL6OwsVsmg
ZIG5RTZC/js5HTCGCddKLacF2CzH/KwPGFI4QkQzQQuUypqX6Lei1BO1XDdDthqWOVG8/ccybhSz
GDs19B+yYvi4GEYXYCf77C/zGEDQJUvoMxgjs+6Q5+KSPSenODOsnENCjzOZ4dpsSPW4cSAPeqBA
LBTWwVJoN1C39xOGDqMVrpe0QPclQ/n10GIbpUPodNTqYDYik0fNGi4o8EPxgenYXcqxMWwOAJ2i
wB+Ptbd1ZsNmjpiwHuaLGYJ7H355t/wKzZab3ccDhDdxqMo6QE8kqYwLeeioRflpH8QeaJ9IpauE
ZSZTf5ERfK+d7D22rL2YPTDCafEEm5u+tLfOCzFb9XzYLJm2UxvoJV5C9kBGXVaeCOkxbRbwb0p2
n55dXzG3jzEiV7BHTExDAYkADpHLYqwzK4kkJLCw8Qi1VAlmG/XmoLEUorwl6guzvbJZQmSZ5oXP
6qy66Ml5BLs8V+DbNAH4r7EYYzIS9rZ2BBUoMZtMkpykMwp5T0vKqYR03P6Cvr284FLNm3PcIAND
1NmWhTzg/1FpK/ePcfRH+D9jM6B0lnyKAryYkYZjeMCaXDqH5oXY6o6ESqo9C/4sOp8Wk5RCKUJx
u8uie273JXvscrbhrrogoHFrRjIBfkMRhJFv8jxux9cvNyoppMYLvXc5l1d30/L//JR7uWuSV042
C7EfWvJ5anDGnGyWkU82a1j9FbnzZakgHDC+qqf+ja0QZIwxM4l5gvWTkkCyM97nPez3NPvOBo5A
5MRE9OOjeTtBbiWCha1rzowaCHjyc8/eTvrNG7bHGQHwPxf3FlCKAt72mj2r7DgCeeQ+0SRyHP07
TS4z0BcQXj4Afe1HPr6GfouH05KToHT22ifIh2MT2KzA8KB4URDuilga5zAh5Fs6IpPZvHeCuT8O
eihchgA5kcmB0BAOSxmx1Wd2JBrURa7mfSHi59oSHWCmYGjy90X3IddkuAfHGz9fqliScOJlF2AV
csqSo90chPugH3qqHOREIBahcwSvNi80vOAWfyXBpiJ8xPWSmxXlJMlsp809E1kERwSsDNh1puLU
ZT7rrqSzNQEX/u9nESytRMMtJLr7FRPNAH+VhgQcvF9JWfLj0uPrNXUYSrqwHtOGGfFwr3JW6Jb0
Nh9ufsukMkufRIaSk/U3eAVhlH8mtSa2XHVWiHrScB0KyB1+nND73W1kruybjZF5VS0RuWdUgfZw
emQhQtJKL7n/nDw4e2uUquzH0kl4OCqDZ24Pd/erouKCaiyeNI+u35EPeV2f4aoxuJzC+kMA/AQB
jKo+yPemD07ZvU4XZQ7VUYz1eDpGdeFbcY903rV98knAKWpMhZF4vVvxaPKi9dXFkUL171lDJo0F
RhUsoZQe2+RrYaGrNjNUH5JrjkZBQPd9JGDRKaQOHpFYgizPuQInQlpJezxXhiH+314h6VrXjuLr
xQqePTe14+XxNP44fRfMxY+zAIHcpvcdQnk8Z0qED7xIPBhF2rJe5bTjzt3vd2VQO40a/7ARPA2T
aj0vcCQ/hDiBu9pjf7Sin9o5pqxPKHvWAm4IGNE0J1ggv2Z6apwAfrND0zeMmuC8GIFo8c/2oJP0
pr9wEUFfxv0qhNU+bHqCtBZVTALBCUYjMr6ylTzOLDAf8w1NKS5SWIj+lHWSYEHHjblP6tzjecUs
QaM296Jwf6zXJg5WxAla3BUyHpMxlM66mvUrIz+eziDquSbgGaX95nP5ZQwNtAbTVcAXc7YED0Ml
T2rvL+ptSaMEsh4tO5oe9AJ5azA4OwS0MBBF/bUEJFnwDRdYoZDp/xNr3mR2ADgmqjQXcw68ebQa
Cm0tV4d6Q9OY3vlBbhAeAFu6ksKoCsxRgVaOpYRJ29Qo5CgT59mNNLEvI4byE5Ccnt1DwFiQf8w0
2oybP3StCcGfp7bU/dDlsfWNxye3ru49g4JenjhCGf1k3294CcrnImptV/u68qoyHlDaQUgDDHvD
VzAkgz9eStW/11HUT7Db4fVN7F8aw2uoJv6xtMrQ3K9CfqgtJMjZIzNvU6467+lvab/HxCrNudt1
vIoIyRIvSz0Yks2+TQOA3x7fDWmh5qBj3/aYuT9rOvhtRp/A3CiezoomU3pQ6SCZyqDkRrw9nME1
eGMtm2vu+3rC9Y+3nfIw/4H9M1Z/vkbwNtU7NzF7nM9c5RLUhpRseiqiDPyBH5W0209A59NrNT3r
Lu6DUk3iT+QJBX0bbdZt24KUTTjbcD3w9t63jEQ1/z9M6jKkh9EnUhloY5cvSCHxhpWIS2GCK9Q0
R3o58Dy+E1/RN/9wAUbNLTR0tyLmFG85GpylSnXMp477c3CLB51iwhKkMAIHChJL73TU0BfebgkF
GB2/LFh6PNzW/87Zk/sNtj1LRMFVqoOxHK+hqQpI8VJc0qtmLSuf+ugsw2Jf2L4fVKWTb5ls7fOR
b7mHiUMnLRwQou924joW6BK1Aevwdzi3H6BTDWaq2cYJEmkAKKx+mrw2ycRYLXN/eiKHPvpvHnwE
DEg0t/Z2hoCVSCzLQtC7oJMolsMTKnFPPA3a3KaVW5r7S9uL5nB/A1nDeQxFGFzKCY5SvadOSZsa
TVTieahiOzi/T7QVqNuD5Xq7XgWaor+QUZ5s2//00kdkHqQV3aX0DxEYYgncJvGy+myyih1oUX15
/8m+tGWkY0JdoYYNn5dJN6Paecp82GA/gTCNXSq+5U2qWGWBXxlJHGNopOt0roDmKcF0kYQuq6sQ
9kaPf+8yc30fXlrCaCsbcdjApXXA2lW0v15e2T8MnfExrhd5IZLjnQ8/9FG5vUDS/4/aoz0+hxq+
vz2wnOZhjW18SG12ywOBCIzzdjOR/E9m51xdeT02833qoiBxzQY/pwA8ZbINGcGN0BG5PiX3/Lix
i6T/1cFUv4MEdtbJqw/pK5RHeuvoGCiIrvrnxQRjnCPUb6PFUzEzUvVJn70Z2ThSdPH9rJbzuFZM
c2nLrAKTKnWOh4YRoejdh2LACP5G6uwegVUmI4AJ44RfpMifrSLWo1FH0MeY/vYEM48OQV7z0RuE
b4UIAvHczTp/XF2Xi0LIL7C/i7DnENd9KzhYIAi4qixTu0L+CWFdXBVPdurYElwnLFsFsBxNu6Q/
Om6kB4Ni0hOdrduabZ33IuGcTW7XdGhPWE2Qmm0B8UFK7X0I1pjAr1gAPrm4/b3zEJy7RUyEUScH
T3zODjBNRAn+p9gHSqyIeyk/wERc3FpCBl41Wdc4LeTk3WQT6ys5M2bd7ZpaBr7lWymEuoQnbDAK
QrYDPYE1y19VagoD851vTlGiiaDNqiWWBuuGIOHyC938TaayvUX481abOxlyrDYxVDaAZb/OxVSm
C+a60h3dbY5azhGohNedZwztojMlyidKL3S7IeyCSvlc0rqDd3nIFeLPF1tsFtPlG+wvukGiviq3
fef4AQ8IVOuzCKrWmnHBy4f9XMBqPPhM2g+iAHgDa6ruRUzl9Yw1TXHZKxjkm0JKE1bWorLfK7Pr
P6uyVReTdrVl9yZ406c3j0lzcM2fpFz6lTXhVZ2lLntuktmNJMlSkuzG3NBQK9/wZIbPMY/ANXCK
0ChBIPX1648renFc3sVo85hNavXKQUCh5WgnMshaHgXDk/+WvBHtC9QHndlCVk2zOnTh6P9tm3Fc
cOYvt9NJGeUNs6fHY24BMTbJ4wBNxFHHSBOAQwsarGeGAu33buozXJTut14AnDDqmJku7LnVXXsn
hAQMtxXCV+tBoIJNvgjciVIhVAGPu1/Ycg/3dmT2jjo6ngxiUbT2MLgLoCXip78Vp0Fe3RELrGrv
WnDCGsmRKZDFPPCkZprfXtnrMHVzmvsOQfv+aYeuzigv7oPNY5GSoFzyQdZTwv6mtEV3ofh89FIv
GaYzEmiUUtjGnNAUEysBZ1nttbx9cBuJa9l6eo3eB7plr/5/DebGSMy7fGGqMzm8OCyq3ZMyy69q
8SmwBqYiCCWmoNmUDAmJCplx7Kl2W2P38iBn21a4NCsis1FdKXrYSEOVYe23rBjzdMZxSpcBQ/AH
+SR3zLaP9S28xkfDsUNCRchi7JXPeLIcyz+3yzvYmlEbr0tcGZ50XpemrKFpCGrBfkCQeCqg5BgX
qaDr5C+frkECXcFVYm4AdwhDXuqfPFS953PS7/vYuqgbTDWbJau5f7kxFi36g28ZepmMCKSalvOr
ojx/Iar4PiR+KK0qU9inhVLLCWD2RlJKrrA1fAOaeFYOCYQ81YWmOhO1sVuaZpqUokEEdyHhcmc9
zXjqo5UopFIJSb0w0S5BZQ0JPJ5Xb5FmxO6z/mk5D5+sB2FdrsIK8ZK0Y+16OMl5yEiXuLd9wF5L
Iwy5B4wqLrn7EpCojLs5PJO15YMGsEkBUbop7BG9puE9Dg7LMT1Xs4SWg5thxO6WYlm1LfexA4hy
2QlC3B4pdQc2+z1w7C+RKlYl3rKyHUzt2OwSIE1e8SCsp1pult8xSSAtzPtL/IH1TuCdDmXIGYpz
EBS273rvDVbU3C3D8PMWpUuyFv9Zzm6dtb/ZcGgEuKFt1iZ8aYz7txCQpBfowymgOqHZztwU6opZ
Ur3tKNEOIP6itKYHBXDh+rcpz5tN2cy4iMJkoc7/gV583vBn4xM8c/LHCUZ5mxUUeeX94xTph9m/
18N5s4baWFZwpZGaWyclYa9f0IIfXQo5vdGZ7BmJqa1mJuTnxZOsyJylE6TAXSV0Y5HzVpOLYI3q
DunXac4zXriW7QytrwFxUdJuSXB5LatKZHAi0z1gb0DoXr2v/hDtWOLN1/ygabg2z0xcX6vW278/
NmVuhhrND345HJZE6jgGyWcDHfUuCWtkV7W9W1wyF5+DRlOcmqUZFhcEbWORwTMjwbabqnFzJP7j
NMtwx4bgqW5Ah1iZiz7RW/gBfyIWEwroe4w77Wy4nPZ6htNc801KmqU+zEEHi6T5xec9ujYXHt7X
c6bGi5419qfqBRUV86ds+uz10enyIvvLNgL0oikfW5Maoe+1MWfwKAvFWc9o62j6Nbl5xH64jg+o
rGxbZNDz5dQdORcbzxrnVhIjNaeXp+viSIBoaTBvgCG2TmDjT/VdBDRQyyP3XmNWo1TSZ+7VwZJd
TTE8R7JGiC4zgry4IkvmmCridi/Ib5ek9qNOXEvWsamSY1t2zLcvZS+6j94JMugsKUkI6cXbLsdx
rxrgErSgXRxujsBdReckalrEB6DMs0yxNcDhxlKVAe/vgxQvL/Zq/QvOM1K1NYalXZ9mmpc2QeUQ
hX5i7tm0gWtm26/HVkzfH+6z3R0Pz9JssJBnAap8CJc2FLfwVn1lvdzirpA0NN3GWR3LTVfWXHRt
FNBrwnbO6pH3Iuyf5U8XRAqofyzMsJb4C4u3tITVzFxgj0Zd2yZQkVqhBRuRKkNVQkReH/C6+A9q
/odq9Q5e40IctkotnhZDAe79JgJ5d3MNZgKCnwE1GhL12epyhtpG7flE+UEYhyB/8l5pwTt1hW7u
KnZXBBBAy6+l67r2LEdvm3c1RCEPBwa18iXj4qt3psWAHBpkVoKriO+7PM1tuDxqK5POVQzVcgHq
JbObJp16iTNKNifbyRmUxU7VkQuYSGS5hy7dc9T24EYRFONNF7G112f5hfTTIBM0qKKuYTorIcWp
mKJCQachPH77pFO6If5hjp+K2aqbPxepJisumfj4KS0IQ0HxNgZUzG7a0kxShJh2r3toKt99UN5V
pscGoUkohL4oif8XnBZEi8hT/pndOWgpqMRU8rOCvqxkgsVKwb6ILw8+L3QAk5OFh/ByThnCa3zd
rLu14jtxgAYsgn3aZA5UxDre6vXxDzl4fYVc4Wh4Ve0CVOwDqi78hl9BGf/DjL1YAhsMDJ0byKlu
om7O4gx4NiaR7uQCVPAxHj/58iLVnUntdaP1860yQJWMaSye+Kr8lov4YVGgXSt7pm88BOXG8L6j
QuT3r5fqfLneix6cNWahf3waLaCG3jCS5mU853sShUUNSqpf9eeXMmMlEGUrK1o6FgO2o9zqPAKz
xBzP41eD/q4XX7MBs1TCXMjmzrVAFiEYK76ZU26l8A1RPFJUbfnRzX74EBkw2RiaNu++GMxunAAf
hsZE4nwOL0cuH4O2h72IOvPp6YcvBiouxd+a8tqzgno6YLAplJiXb38gPVubUW1lJUrgcQoZpC9H
2yVBTfHCwJEWO5TeP/jcBFuU1xxRn8fQjeBdMFegmiGC622inI9NZrX04cYcCWsHGB6oILF4Sqwb
3kxI1Ugh3+t/WcXQByAQLFzRNUjRIfdDYvRP9EBwQmCvbwo7qCv1jVmhdzuQs5m6x8PdbtXNAdC+
LAS057iOrYiytLDJb8nVV1tjjtV7o8FspdHWJqz/ezCtaWLJ7ODgbBjD9cL/+hqNmqbQOOHnoMW1
o+X3fE447b1p2XV3stSrHaEA1cUhjX43WjG/AIBNo0M88TEmqDmPYfxr3+6WPntvB83X6IcTqE8s
r8nSmsdFMYFCDbT+di+Z9UZnzYVTQkjNU7fG8ZoF3A7F4DiciVUFb7fea9WghBiOKbhPY8mE5Gql
1OKotNOUmNICqxZVFPnLwzRkr6+0R2lJp+EczS2CNwPhbwdZ6lOMS3wI+vh6z4bc+1CUBRGBEMUr
JkHH0yTp0NqEcjSjeePgSSBlCPi7mvK70NhYgb3UeR7tLPHQgijOrkr0D47WnKE/dNN3ZXd7A0dy
y6hUKDJfDnrAq6cFQs/dGqFehk6Q1R6O4e2+fohycXMvrcO2xqd1nHJy6EtllCfqs568T/OEpCrs
v93rYyVKeLRFK47rbHQtFd7+/qdQS2xo5qtJy3KEAU8kVBelv49J8nS1YyJpvT3B7rBXTxpGzea7
wQmMR7dal6IsX2PvRdT1tmiMrCYbVPeSjacPS/rmoXi+wzMHtfBzrJk4m9o70GX6FBQI9Ev8lYtL
3WiHenBAmr4HDA4ix5SXaWec4Z/ewk4b+HoSQMtllQHS48n1qMUVZAuN6YVfF8/xycA4RhxvWeG6
ePPVraYZJuRnrrtOXJupwcrQODwx/Jc3JxWZ6cturlLud0mttm4CHxELScGZpLYaiZvbU5592cwj
g2JjhFsKR/aNzunTzdgzFfMMie31Nb+0v4okBD8OmQWC18LO1FO25agL6tMczjplabC5V/moAUpr
i44kLWAvdqPrPbW97KGubIAgitamQKiYzyt4KMAUEC1Jc1mH0ZdSfs/dkquqX5XtO1XtMaElyiAD
eoCPeerGBxlsNYqfbvK8kR1jJ4athA+SWgbu9A5QkiVs8Bspl83GvMvCRASJ3gBNmy2/p1JHl0M6
UZKpBzajfRdWpNH3iwtFpnh6BWjj655riTd37dTejKYRIM5Rn5w9ytwAitX/fhFVZc77ecEY70I4
0thaPO4BeX9t2JaGPFQ8FnYtuI7Ohh2ljpgGKvUluvlQwiQYMkNzc92cIfw8y/Ny1kQ7kqbIZoCM
KAAP1KBdsPAjppmRdJ0qhZeNzjT8/6mE9GPyKeIZ8qbe5omliXxZJhPQwmvE70sUl801UGVITYnc
wsP8uKrdXuE0ZWjcf7R892EccVXOsbwgs0p+8SCqfHsPD3uZ1jaXTmIwpEe+Y7rgWvPJLpY0Rf9z
373/kGY4OBBxf8556PNkLMp0BqA3eikl8WB1N0t9BDIB++euWrtKrfOK9fVCKgZRJ5ol5ABJT6xh
pji/SaUT40atoVt8IOxXYmd1KytKVZxzVGRMeLN4DKbRYIWG6KT5bOd8dGQvjF6FDGLr8UVejXdq
FLjtg9bQt0gg4TLmT3P3T019IXre9GnvdjNQWF84leVLIgKIIhRviJGjMjvd2C60OW3L2pIpM01i
phH0uViBT/rD5mYoOSyagM2ne1bCjrY9kqhUkTtqpolbrj7aCm3+FgveVIH2HJ5bmvtO27khZ2Sz
ANXt2YtbVZBvHPlMvDeftU+gQ5B4rKhxNIVG6S9SAuZsH/GV5MQYYlRLi4AVnDY827ahRtVcgJbn
mxRGEGmyEgCltheRIxL46bAB54lh6RtA6Nyn0d/JPH11JrLlLOeOZ4VszH8IaInWWqzWwVBbOU79
PQhRjOx4qNRsfs7bv+MkXNgfaFdYiP536mPX5X3Cjy6l5I893c+1yVBEmAkhNHtp59cNgJtAz4jc
JaiT4WClPPiXlgiOq42R4Z20NPKAaP5gzXnZUVoISVJtxHJxtHePghnXTRnn3qszcU32clHhCJlP
AOvEKEq4vfRWXCI8PL79cla/cma3sBALb6zn7YZ/Q9CZUxlUZj2xnPsIWT8opR8YCYR+37tWuTLA
UoBJQfsjRaHO+0RzB16fwbF7TBSSVQTfddTeoJP8CxPByfe1/TzKQf7i9Xskjs7vjG3wLUubs1wo
u3WotnG4rPlHP25l18nuP9j0w6xHx5snmyZ1QYPhwjo7mR8yJtEHsACVnf6yqAyxiTux8pohTVMt
nTUmRKKF0ttH2bsflgTGenmcy9NBTvGYRB+i/skHUigQEwcXEM8WKXYHJNXS/fXuKPWe0nR1Hjfr
F6G//fzmwBhjPQ/seH9WEkdUT1mB82TqsdrvE3YI0uUWa+1TTINn/IZuZ8Q7G/wImoeFa1GWGppY
yoWgKOQfjjv4Z+1YDLUyv1c4k0jUJi66THdRLzOhMuGfBtfmZh9jimvi+NUQkZb07WwYS1p4vlCL
IIr8OZPU2xeuhO2OfsAT+5ybUdSCQjFdkUyDIvA24Uva4HGzD7EAkHfaLoRKj2l5vD/mZTvVty6+
TrDs66vKwyCxjDvvkwyz5POyxSmtruKHPI2xAN5wTyshIplclWVxk3tmKaem5RFAIgpTwfchqK0f
HGRwYAyfUELkTlxDpDYWEGh7DGcWY6fUfUHZNp4uKSnun/8+AJgUE7O18U1t2W12FnTnoPZ90CE/
J7Q38BIlzyJC7tbjt3DQGOtn1GRVL7n4awq/KD5/nLaP/W2WuUVvtXO5MtZfTExnG3FUZc3WGc2E
OIMax8Fh5euQWIWMqNZSpTP0My51CJzJ6WAq71jsSQ2+nxMbTTWo4nxJaZQrgFqwnrtevRGk0fCa
49JPvVra+UUfYDGOrQ5TDLvnyRIbnjMwi+hvaKhS2IpK+RIAIA9kkiY3sjvr3csVuCodOCzz0XHg
bKGxoZShWKreBoF8qsYD7154zlbgK2s7ohin+03kzQctP/GD2B9qbWkHBCPyC2XLDrz4DzPw043P
MEYUX7oTYi2CNU82CWxEt6xI/jiQMOKa2P5qxgllaNj4qWER0fWRLOg+CcjbjG2ijoxhCC+QXc27
2OokTGqEvkFuPC5X1H2slkQ+/aO8/FWyOjzEbGnjHKAb0EYDNLrktkjxUBJcNdJLoONSrcBO2a2j
Cq2U+Z6V/e4qKy64oMLOHSZe4SnD7Hfx3xPWeiJDQ8CWNB2+0Rc8B1pqtl4gs4ilNaxdNd4JCFwb
qvLnyyk9QK/90jVfzsEDhdDQ+Y8/6jl6SXza2vVWqwI+jN7o1u6CaC4JunGpeoiJtgfH25gpnbKJ
qQRQqYLKiQY3ybH0R77hMd5OiAfesq5bYnw17GHWUGraeFI6rgTThjhRg9eaQwA6lVAB9ECl8sBU
A46vghDkzHy60DvGkrKhuTWN3eRAeirD5vzah702PX2cnlKFl+Xr6s5JkDhgdr0afjWZHEsWuxjc
2P3F6dgGWDpdOv63jUASOeRiCMhRQUP7hCHFYYs5HYIWONHd8QyOOJpYON12+wHqAlt2g9wLIs+C
9ppG163VxOxstIbVj1Pybck2OJs3bcy2hmnFgbKghzDY4Aqpb+1PWcBYqgUiLyuan94PcX50jk1p
eLXPRYykbPU6wJ4U+jicbkXixSN37thyyPsYGXU9XZXtPmKhuVjxZnmmr2Ws3wQ/qM6XbSmULDMs
T3Z8C6uOWrODLn3ANzWCtLtxVenTHCy/z1vLYnLr3t8ARX5ve4yuuIrJaOoKis8NvWGYI4sep0Bh
JnW1DtQcDo2+UgtnLyfY9c5aqvqX3yKtOKdzZyUSQR7ikN82WcJOTIqnJnlzoxxRnhvo7XLfL1/P
y1nil6sLJ+xowDg3es3OQPu4KsbZgh5NTZQ2MBARCKQHTxLCFc3XSvefHQ+3hh0aVOwTVAg3RbCg
kKr+1wSxoh6GQfxPi0qywtHOhoO5jAYNVyvwuPdtHgQ0Ab2wkbQnaC3VMz3pDL1DNEoueH6g0fMS
w+1tBa7RiPe9prEX6S4r+PNWAlcY3bsHGrda79s14tzjv8OUPT5lJPGb6jWZ0O3OxWFLdcNQpgQT
c/4/IPXXiU2QF2YEWlB4agR7XNDxRWyRshqWh1mjNNIeKFZa/TMbbDFOkNVrF5nT9USdyEiKS/dY
Siw6JHhZ/2GA9uHyeSyGjyWKqoA06/EIZ2O4Um7wbfi7aniE5/U7I1MFLagjykKObQVDs4TdwsKg
lLVNd8OZvyABUStRSRLNtSKuonQ48de3fnvSQYcZzIzhuxHSaX8BaNCDxxM2a6jX/PfriYe77ZCv
VvXtbg71ZApyKdz0GmYh6GwgttgQ/kOSteLrlqT+ieT6vQ3n/IDKJbvyPzHs0akOI4uBPDchYgvA
WKNVE3hySeBNA7yA3XSo5KQpPzeGtZKB8DMmfaVdVgGSvbY9022VpFbhHQ+FttszaiakzDp8jZUj
PofK1sFs6wNs/juVXqY/WY9eh/OpmDiWNd/rGW/G/x25lHGYUvtncIE1yTc2rxmIYfyGSMq0xAD0
QizZbuWIx4dRObNiOA8X9C1Ci5gdYD2o6krVu9UqkQKLpjfyrwVofOsSzldLteoiIWgcEqIKR16h
1vNYilVFXxrbP6OENLwy15GiUhBl8OEzXjrnwLpE9oT0RCszCvg1bs4DIJpWh5D2zd1BbCDhHiob
/yYFLGZ7ylq+Ox/yJB+a5WEdnvbl2HpoSuMh/1meBx0L5TVHA5+e23nlxuG6/YbzU8pLh/WocEhw
6/R+WbWqzB84g2fOgsIKjJKqD/p0zGMpmar1oqU6BNKsNhEL5Z6Yoc4RaXAokf6aZ/5gNm2f0y4Q
UDCfdke5iNWyJAwbATjVvKmgrkFlNd33obV0zBXsEy+DG2gp7rgct97cWr4fnY1JVfiBiUeroK7S
u6t6umyit5UpymqO2Uie7I6M6zqDux3snW10h9j6V6yBBYKFArYa0mhgvk8B/lt0xQCHlVpPrFXQ
GOwPQ8TuLCVqgj7c+hPCgcUEcFl4dVjtY2bFW1uJlh1GpX4SGyooeq91U+6ws5tZOQ0VXDeoeA/O
cF1nLlgnrNTA/RPeKMj/8g8T8kvmhYbA97IjSgSk7rBuCCDZUGcdq7AQnOPDNHHNR9D0uQZj3sR6
K6z2WK7mzdgtZz2aKxg29Y4u8PQWrAb34nFjpmj320ZOhbzX9A/EYchg8oaRzhRtyPmRfSs1k26h
+euyI1R6O4p+Cq6Y31vUztoJBpdNkH2VzYDqlVkoGriUr+Mglq1qwSJVH9d8RtM1RCf8F9Y6VJOS
4mmR+uK+0NB9gxPsRtuvVbWFc2ZULG+iFlzY+wVepMHhNj3a5DswA+ephiaXRu6nKMkwi1XsYHWw
62FBdhmwhvlyMkTz54o8w5mFkLmYns8GxVSWjvmwmG4hg4gdVdV4WaQujRP5bAKmH06AmjA3jWP+
+cS96WU/4wzfovpTGyYH4Sr60hHHUJC6PQQrIlbnwEfKz1kfrBu5zDUQVoffpyYTGDQNuUHenmvX
qqQ/hSiR4mclAx+6vwzcsZTsWMoB3npLFZKuUEEe1MvwI43mXiGSLiDS+Gfy19o3hST17ZDHB1eU
/MCsf+tbIkRuytENRPcju7UZ7UWoD5kx2FORdIY0cH8SS1iMUGrkOqcdRJBxcPo8n1dPR0q4f+KE
rKdcD+HgJ3om0SUuO0nM45Li4HGVsrQHG/s7QaEN2HAHdnD0nLBZ0tTG8oZwI60ufY7Tdk87i8q2
J6aCjpTA6RqThC0/YHbgs1c6qlhs2KEZfHtlkOdhy0vG5VhwPRSDjRemLb6H+XbdCCnQVu4j/IYJ
wteIeZYkvoeUl3sJ14SsfmyBUvMD9MpkouopWZZfjAesRS+XWjZJ3QBrx4Uk0Fij/oexcTkkJvYX
t8DUbwvttaDXHVz9Qs02Rq//eiK2+QfJ1MfHI6JzvvjAYLAK3xeoJjkUB/OpfUz89o0PWyWXwFcx
Rc1kVjZf2NTjZ6Q6wpWWeRhS+YtHOYUfLgIgeaS1pY1R6cmPPGn9l0PdX80Eoi8KbRfEH8dzicUV
M3ShdrJl31KPev3m8s4Uo7t/OFdqQF4U37WIKuvAyr8zCPTgJoLZtSIHQPJOa44FsCWoQLUgHfoM
3N9mqIw+3bXgvm+sogqTi2l9hykmkyfbOzlz/zpWwurj1osag5QMbki3v+yNQlV8V8HsyVH9vStK
DRq/UL8dM0rXzRkhf2g3ZxmOLxm535VCwJ5Zx/t/tDtViBnlP/0AbhI4y53y2NEEdCgpeJVF7D2E
o3IJZ4XDjEdQXtoPKKeKT/UKrXDKLijmi7ElA9HFXnR448Vez0+Vr1Q9/gMeEPNzYGJMOuEK04Eu
nvgFXkHsyz+paSQtZTN2KN9b9dUGes4mcAERHIVI5beZT2ZokuGA1eY5PmEj8HPNm6UaY5jGs1Za
Ryh40fJXf4PojM9/6Q+hysqCfwlibRmJI/Jgb4f/vcNWmoA/V5h/p0CRPQTzGtxrteHWyb91WmMS
QyCM+E61dxpeP0mio/Vuh/y0cHKWeeTaJGNa3HA9BQjmuR/kOebQU04wLIZFitBeV9miczAIhPrE
8Uv3z7p/aGGowj4IMbMPP27SPYHsBSUHoZ9ZSZYq8nBd2/QRwBszDDLnSHzGFgMmi7bUZWejOnzz
axUm7sSgyIxQHOjLrcOIZsu/CJ6VIMpC0S+ptNt4nTwPfm35R264/B1TaTE4Jl+7TG/cuHIZ/+b+
mo03gmInZVkrkv4icKdfHfUfWVaw7u6bunEAuAZiHUk140l2tcw9Rd/c3Qh5tk61N1M0KdeQFp75
hmetczd+1PFI8j8zW5o/+8Hr7tHtOpcD7V7mlkXSlhCzJjWZhD6HDXqS6iHSUgXydhifCNHL1oCa
+u3YanPKw27Rz8oVLCIbgRJHM7KE+gT8QWHRMZcCiMNBqpKqWS/5IJXr31LLQGQFkEPNMZB5t4bX
odGe3FcfXAM/AKffOev4mV5YfhpFVDGKrmWKQU+JPBRwZMIn8TOt9iUlUHTtkFpc/r3KZEikjQSV
O8GhzNGvwh8iuBLKONXVvIeKAjcQ9ZXOWsjxJGYFIPD1RHZfT/f2cHEQYg8OFzlb9qA0L89pj7Nr
GXpQaoMsQrshGmCeu6jl1hsV0XZpyZRRU2c8qcDAOxlaon0o6vF7kdIbi0FLKnd9TpqQBxdQMnnQ
zdOeQjNaKlas3ESnB46wE9pAJahncG7OvfWOxDjNYabaXXk1DIXoeGbNo45H+TEkIUsW5WKgvkoc
Y63+QxU8KNUStPyc9UPOedIfciSvrc0C6omIiboWJMT4kuttUb53FH8jpFnBwd4AuZ3W/rmTtzcK
ejTU2UBCAMf7efMtKPIH/GLXzYYCZZ+CYJxmgHcBOomsIOBCgVeZef9K2UrBPzxeD/CyhK+4X+tp
LDYSbbJxBMLo2GmllEM8kV1UHbHlKgkfSi8RYR3oTmAVUPNAZKPZ1B5TVEyjOOd4SdTZxypwPdJE
LvXxdX+BUfUUsCU7IqiyqcCJP0TNJwENSrrvOS7MduR+UEOywIR3H6vu0K7O2mlmG++EDxqFDODg
27PDKK1TewCiLE1m88T8yFy5uXKkxm8W3pNo50Q24sXT1SX1g1bx7L7ublEz/YoD+BdElPEEgxiW
G+PFZAsZDYYfDE04vAl9g8inLI5A4RINb2hp10W3rxBgd9ZXz32AMn0q5ULvdB01D0p1OIFL2Haj
Zxw3QgTqurG2BDqV0rFY7LstelJzumcw9ZA/A6C1xsQp66/iZ3FMHi5Fow8llwHu+0bBPl4oLhKQ
6J7GaEYmHGJU/fQtLRB9RPC5SZaZCGv15KPzGaWN1Z4X7odSLBJAE/crCbztAPNK3IyE2TXj3f6f
19sN40EjQanzXiF4d3yCXresT+eoWGJxPLY9t1Pvgx4Jaz5+Z+RTcXgjJS63CxO5CjMmJap6M5Tt
OlFmb7GT4yrblh2P5sjziTG9JGI1rz1rNeKFuUfKMLiXnoI/nfeppUE14LJUu2SXSOm902Nvxl/u
Heve6BRUIBUnodj7AtkaJFnbtl0yUExS1xUeLThhbRWY1B0WfIowj6LPYkag0okpERC7D63i6Usk
Uq/dqvutlbax3NElFffC3QxvXoszglc2GuoTJiNwRo5TqncxFr4tup3fuPdi5Kl4homvrDOKKDtf
Kz8dkVL83tIaygIYce1FMRJN8PiHYoxePGed/Hx5fTmpzRiTZT/4aeXznMC7gJDbNalqqcI7BSyx
zdABMSCW90rKRF4f47t0dSfHH2mlJpmk8gnIE72v/G/C9FpYr1+JExZEiiaZOQBpBPIceZG8kp5v
7eOfzVXRS0bUnjS4PNvcH1OHNJHz5VdtPcNjTL95xk3tiFIWTjHLbrCo63kocPPfMZAMyubHVDqp
ZBgGJ6X65sUTuoVAR1+YbvsQlcE55vnXOBP9vFYxCqAy9wS/Fk8BZwvdXpH2J18usE/NV0roYSkD
Iyc40f6e6ZwWfZkIYpknH9Lr2wgCqrczLd+a7kYGkwkfOrITn/c9SjEdF1mUFJtt/oVGtdgmQ4+G
9y6XsdW1ixxeKNYwcMESEMli9M3bAOnELk6kYWn8JEIm8WtWchQNBX2Ld7jE6Fhb8qMcBF7Pot1Q
9Vasm9eQs2KmMzAuPBMbTAKWzAxnmfyWR4oRNtgqiJugaOVY0c/5siGgsJhUGdLCt4DSlCNeSTgl
LGqwN6aVhlPlQu3XIpWfFJUikf1VKsiwP7uNk6fkbroZrilPb25yuYTT7IpThIhujTt8TVn6Z+g2
Zl1F1MeF0kclguGjiossrlJGNv19Pcg8q9899xriHqZKbUDux/+12t8Uhl0EfGt1EYgEPF+nXJ1r
+U1QS/7Qc/i1/REzXed1p7jsqGrM6ngKTK4vI6eopOb4otgWd3kB60fu1Ohj089W63cWQpyRB+nv
bTiCucBxomZpBBSpcegpe7OPCdjGdKTXTybEhKAaK/G/88gCbO0Crl2hCpUjGeWq7qXglHWOg4vU
Q9prAc+eRpakj1FTahiDEOvmSic7tzuxSwKpB5ZP6Gvi/VV5g2JDR1Li/XZHOSPQpooVAcI/0rxh
pBT/GAH3natC09k1MeoB6yWuKGyBOTKN1lQkXrdp/0pzwgPKpOnR26cA6ADrf5AA/BN30HPMrOQM
gcncUn2Lz0mgkZSlEv91SKSID9H+MoUdiUu6gRttB+KKp7oWXXIjXg+YhWdkjL/7HM35H4SOmNsY
xyMKNCn/WccZTcGiVPl5oMrfDXgmVOMIZm7Jt5DQ0zB2v2BbyvMciFW2xXCtD9ym378057mT5CIn
d1Nf+IBAdT3PySZjtsM6UVqD03PfcjaeRSnfjAgfifNARRkQPsM0w7v7IOOugjU4HFPTa0eMhEwd
hHMmvduHl8h1qZ5bQP8UAquyYXGQLkZMgLBikkiAMX5CBbpLjhjude7AlQqx+vMy12Cz4kd8KxQm
a1wOW4Fwa7v8tmuxqN5xT6ZrRDGxpEZJHlcyk74u1Hj9TL72cBlVbcTmDCJA1aPkdj+350uOt9Gc
Z3ZhVn4F3n5BTUajSoOh706MGdmP4vRnOCycSoswXd4YyreMxBotUeYDw8N/0wupk0W2OjDL9Elt
flUKhaEXXmIsoZOxJN5xAB0/2Wk8xk1N7l7L0Zagws5DTiNl9wOL8GVLSxBmhRsmbqVFnMcw38pd
/+97ywJW9sR9aGWxgyaO0Uf/1I4PveNvXKKW920Qp9ALvQMLOIq8uxtIRPx0FfoLa/mYKI9jYQDV
+lJ4p1DGHCwg7pQUCi1PP25/HvX6QeAnaM5O25mAgPK+uNnDqkw4jx4qA6y1aJdG5YnsXZPacAAX
KAVfmdTd6Nxt6EsggKmM3Sokqq/h1SAlsIR7NBvxAkI+411XBWcjMcMf1c9QgesYt3OqtAr+0sgj
PAivIsbapeY0uj4nZosGA3jmge/K1aWa/TB+rZbdeo929XlibmymTmBh5LNw4/YSESSEt20JiBgX
JE8mLAQdmtdifrsTkKQYagESBSgDsXF4Ml+yrrLyb0VjrB+kf41VvsYBoFZz/W24Ds5WpoXVrp+7
F9ab6gOCBVr6klJGVSyYBsv9bMZiO52hXEWElJHAVb5oWrV0vD/gWsgMQNsKDjs5EZ+0avyLn+lL
0BcGXw9KxhLwvjSzJCMT08JjlPkXYScnQACbk4e8Tzeqhcc1ndUonjyU7tgjHWLQDezcx0j/mGn0
kMYF2DfEKB4vl9HQRq3LYNdQ28pfYnxrjicQhN5gIE84w559K8e8lr/nUKQMwSQaPyyJRpOwcVsb
dmmCgsNJccEplTrsd2zMxgCPMUI4NXXRRVf5yJJ8L6jab03FhU8ggtmzZvDWKM5937R6O7QWDAUy
WcZ8eqgrKGQrNg9eT8w4JiPPGpGdH1TH0IuFdAXIAySRGSLlDp6GIQb5oCZ6VLsDGSK2ZCatuHy7
q5X5ZVpGrjC5kC3vUL5/YY0bLqNe/s406cDuxNM6VIDh+1qsk5qn3oQwNCDC9pUwLy5xPy1cDGz/
HW7jKA0nb3pOnDx19uZbmxyfqrzAD8zprC27kKQB0bFk1gEUcZHo776x4I5SD6KH1GKm02EUCkAv
a4V32VEZTrkwN4vzTjlGDOz8U/kqVYYTl0UgbJubYK/eKlwIyoRtdq/NZ9fq83Eb9n5JIsne3ogA
iapw0PWA3q07ijDpxflAze9BRCWlkxfrv9vSqYZ8TIMhit5ZUWqDXYqTYmq8YZ8v7tX8OMuqlTmH
7Int0B2qAymTTCzwk6oCW2RG3eTFPyTuuvdCLnfaBdVGzxKaFNp4Uq7aLNxGsNi34mQM+i7ET4uw
qI7J/wwLn93HDUIYDHNQo/4Lqv5zcdZXQLCIPeGHJAv5e5zUQHm9Ds6Rz8yvEWtNXB5CQ379K8Cm
BDQCkDzuvONkun7XCyUAu0AWfogrjHCf5p5JQ3dwrhGO2AA6K4oC9DXaztiBQstztwmjMpaOcyk2
a8BT37myzQXll8cU/+2oUNHSyZHYDssL202FJufXJ4vNm+FejhWy1zKlIwOJTMNCdkgJQiGfma4y
4nOTbFALbsW3kXKZMh591G8tQ6j9MlAXhmaftxT4ZznBBZqli93kew3lZTMyp6+BNAvZIGmeM7CR
lFt2ivBk+mr6OYKfW+SRNCyEijggptvI9lvlYg6B+dpaEpPQTBRxNaKVkQFlXMVzRIAPLlGPkQXx
hhk+YF34cG7Rhb07jh3AcbuT/SXlSyhnz3T1l1sWXy0VBd+hRzWVCIe6qP/+u71tj2Jiln0KxRpO
tWHTSXl76ekik9IQOMvMhgY6mzuI0bVjS2lPJ1XvNX7CqqojzZ4KJPvjc2C4IlFOq2ThJ9l7X08K
xyLNWcUOup/tk5hlqiBLRQA3zvUUXf8oTnFaJpOeksMg9rD9osBj7C1pQGes6j7PQaPNZU13HGa4
xvcoYlW+cYrcFlICdzGoISS+z6tZPwOuS7llYAY4ASDAgddsnrZ+PxFade07vKeZIewjl/FPrFQc
K69Rt/h/QF5S22F2pkmXaj6hUhigqa4+c2bXpX+jnbsdck7xDu0sdhYvwQR6vKxnKxOQMmvmVyFq
UmVWO7J1LGixS6wm8/BD/2FsY/qjlbqO2fSrH388CeGD2l5jVyb0HVFdan1BRd6zdOulg4PNuKGW
DIde7NA5xoy5pY46ZrjnLrqFX10kfomuoQZW0TBR672NIJhaDAWP+L6+Ju8XimdIWLk3i1t7D+fs
p78Ic5i9BEzLWvr44ZCNqnbPOdLiJCxh9rIGFXtPQH4bILMI8RucBa3o9ngsDK4w+z74bAZFDyZB
vJtf8Sy1MEIN52WB74GBgZeyFQR2pNXZbkMZjM1o66oZfQ6SUJTyefMYw4TWvTaNVrWk+fM6yTNa
3m095IggozeKL0qf5jdvIx54a0yEDqL0f0cmtXNqy0vL6rzQHVtxBFy8S4DngrM7eOObuzpoeb0m
IQIpA5A782nzji7vFzqDNTpc89ZHuluoVLJ+QSf/Vtc0dje5JDwelfNFljVfnFaUU5N/eoqjxEUK
I0+bKBa46/HnmtkHW4qio8OGAx7MYxGhSw0RrKS7fp7DLEMlcLTWU305vtVbuwBJ+Xvn8NX9fmRd
QUR5ru9VolaqTQuXIoBKyKbV2hkzKNv6JId7YjpcYkEciUiPycmLWgr19BrJF5L+6wkcHeUfNSit
uGe9roDnZ54+6sWXsaMyNZGs/vUUjBrYtceXa8+PqWvg+CqxUuizOqljTSAuIvU9eB8LltzIiRY9
+kANTV2f6dO1g4UJIloXnOSn7lWunELoqwPK5RHeM8YVVh2u7JFE3n9zkGPRO8R0p6md1fO+q/OR
DnkebA/r+bTAo2XUkAc08oFn2P2Rn3qRTmb8ip6YnHAODRH6AWiTJsICjfD9Gtn5xekgbiTKVZHc
dWA/7dxY+/4PZzXLTE+KcwcrybQk2aELtGgQowhKTjH7jAiOk7yryDf4ABsdNQSONXe93Om2vy3U
0dhV6SvvDuPBXKF93iu8T2A7uxvSXMLcLnmAOH2e7aSbWOs4uTX4rKNQWhdpU8TBqkrhzSXe4ODt
s2a1f95a3y1UZjAs98wvYhvuDNHkrfgP+7j22JEI/B1PI0Fms03lZxG//ZAToUYkn1/nKYuSv0Mn
eCHqaELiHSiYXUMYkP3SsgndcJOpoXCZgJHVPzXp4BYYW7lmBqBG33UWi4wdfPP1HTygq1313IfU
xTwSZhl8mIUFTuvKBOGNicIGIgkNJ2algt/QKfCtAKaSCbd1xQjScIRpDll23AJkkSSvPP1neR/X
gl3mdPn1X2TVtlQi6OxAWCSqLTDGbHSCz0J+KJ3vXfyJ47EEzaEXzBdxu7GTj1G2AEFTdjyi3rVn
bWAgQv+J3DtKSigDT2mJFl1DO4SEgeW9dS9L0EVAtvbgnW4rvTi3Y02Slbx7jC9eLR+lU0+3HaRC
dxShTodnSi9Df/1NuMExz5RDg2sWTOX0XPkFkAoQGKlP2VfE5liC8OBGQQg4aT8j+IF5GvXfFeYG
4cYhPrV5cSTEOD71ppOjY3Xa0SkZpmwJ2/kXYjjlzjSsdwSLoXfN9gF/3j0j8JlCDxJ8hBgf4A38
8lYaVVpZ6pbSlOGRZJiaezQYRiy29/5gD9Mo8Rgt5iyTrMCpysXcwIOYziKzL/tNvrJbMlmL0L+j
EGUDGakfOfPKB4Vrh+qfcA+N8s2vdFEYIfpMvek/vkSb6Q5fMD0qlE310f05STtFK6rExTKPNHeY
UyZ+FEarHXj+MtBCfkSHJ0D5wixxXlCl4+q1yy1hOQ6+C0f4Sxjyb6ow3hHXW7dqJBLvRag2nb+l
ERf8BWFwYimTlEfqpwsKZQDYL2MMfpwkC53XSemyRRj45ueObuWY+2f12mmCix3uGxILch9mWHCx
7gpl6BoJvIh0mWEK6PyVk5lzOeRH+RIR/QBNPFNYu4VViy3zEaFHB7YmpO+1/ojG5x3uWAnHhbGP
zeO3otEhZBcywbPyZTbm7QBcvcmejYlwXBQlmjfJD89R621RDYNXn9daY1zF3S3cCdYtkkh5U8Te
FR7OSAccxXICW72yaWLozXhxxLzK6KVyvsEoRISYh5yZ39IGVCyQ85Dfr7KFACqpMaoyQuYXGOYF
a13jBFhAh8Mb8mwMNi56XrzKwxPeOMp30mqXhS5S38mG6vA6KWsBW5BRygI4y1amMOCcfDkyypI5
42uWdQF1MeE8UfRY80KZcygfLVVg7WJKrA5vxvQ3m+x0+HaGlbI4D15GNz8PZZqwxJwx3u82LL+o
gBJVuJkrr/eY78wEKPY5Obo4Aj+1I+Fk/4ZfEJwMcmsuI4/UGCsciL+4mVDthGnX2nkKCXIusuMX
fQdaoBBWq0dNA0Mpr8QmY30XHTlB7omw5rF079w4de9o/TUzgRjt0anUBRcSUYQxXo4vn5uy7fTl
BZYh7wbL1o0ktirdUPmYiLyoT9/ZOwwiLEmkmCjPCNYfAB57P0tU4BdV0p76nCRP4AtaJH8VJkc+
l0fYqBrZfb32biH3g87T6c25vlaOWNkpFNTZCnqIxJKy++15/UQQbEexwAcAmNVuIe4tF7EE9L2p
G0Yp4mKJPAkkB7s1J+Lq7F+mpSp1NT4Se8GKs355X7RK5Lui0wCxm3lMIca6eiPLpoFv8g7ybVVL
MWyQxlP/J+hUPt5cqrHiI7rzhz2FSkXKXKdY5s9K+IAa0t3ZNkifangZ1JGmBG+9I/lWryH36AlJ
0YVEH2+SgnAOXww3ix+QoErFATrXQ10ISv3dDtX7FPLRfxeiaWUNhsQ9C6OgGjvWNv1rgGAAFTSh
KeYMQf5k78K5yoVnyZ+OtSG7isDF6Q6cmTbzCF0EGo9jE+dNShONOxW5Mic6LimBjoIfDyqD8lc5
DF9mbihYUxn8eVMabWOqaBr8YR4dbEBVl+8sUAsVIaiBn25QZLJq2spzrUnrrD9J2tpyONYIgcoD
YouFfjxWwEuMP7oB1XYzc2BNWwY2DKUtC8NcBCccnupxQO1NnyGxy8Put5VcsSEulFE7awVLwQBC
X9laVmxmJu+Mh1bw7rO5scBiEy0kRBx+28K+BdRLI172IIs48/+wTQPkCv5rXmhXKMzCUQWEPZae
m+bTLQ6mzqtLXNMbdOfLQNPrcjmJaz72kIF1SJFKVT22qqDY6Jel8x1/49GCqkTDAIVaxFmY6Kyz
ktFY3Op8yvL1kZ0KI2rFmBIHtbPOnXx0ggfSLBWGrstqaOvhREY/5YUVJp+ZeEFUDYnZNtfu/bv6
jDVPiP2/J/AWkx5Igp91DEQn/EYc6XlllKd5iq5oOArHT9Wdvafj9KcNpdXYep6MtaR6r1lgkgB3
hY+H+K9nv7v1osxH5bUcRnmeVL3ET3A1UPYDS24XxR/qa2zT8uPq4KKcwB9J9iTQN00vQ00Z72xK
7ZMia6/UlpEIr0fcEofwe5GJyvcTlgDKQc4m+yFfwus0tK6jffHLxEEiGCZeunqX5VG8m383jrne
q4AZo/uybYKmWQJUs4w1/pqWXWj8S8XtIN+/RmXZryvwA5+W0RW6EcGWVsYvMnjvDMv4WHC+060a
TsSdP/JBiusKfwMD/xoeD22KadEj+AJzcEgTXm2Qr7AkmPxE5Hit41Pkg4o07zGWoem3IEQHqoWa
4KUTsBfcgUKspyJS4YTUwIYDuPh55NzfFWL4VHBwUwsY5kC6P099OUlcne6zvr7qAVkrTwHxNd4o
nbmAIAi03O5X+q3gUipABDgTR9nRkfrczsj3nPubz/ruhc2ev0nlVbF3U4j8xF039OoYs0h66zoo
DumbGF7iBz/P5unW008492HBcRr6Mt5o4dlpRIyi7moaRJCQR6ZrRRcDDx88YogQVeatzvZ8htCZ
fCulzjJfAvJmzqDk3q9WXbWLqZ1Aucr8iZb6YYNhlogBB23TYdKwIYQFM5GFWPCeZEMyf67W7zhW
4PIv4WBQVX2k9xmCz8o+KO8IaNzPBbRhF3fUqRPdJcVJ2mcXxs+ari7eFEQSQNWJwQQouZOfmtX8
t9S15/2YeAU5Yq03dOU4soNyMwJUK/U9etj44MKgfbMcZ9fVALkdsI8QAZ6bNq+DpH5YOUpmjBt6
Nrmvd6kgugtPafGpB6gaY9zqmyxwMeUkatdvNLHTmrdjGBFiO3W3v1m55uMckpIIEAy3skmMilRc
LfA1TWaNj9rkQ4Ls3nvrY0gtfjjFXg/p1hYBLkRitXS5TRcYiO3+V2XAbce3njqSCZwp4+01X8h/
w0CLgzmKt4UsowmzeGMwXIadfhFwR16K+L9Tx+AzotvQUI1VMrmrvIKt89zOIy1NS1z5jed92JRD
SIErVpdw7QN+UC3dou/zLQHQ4qKEH2uWGSZP1LY1bm1W0O58yO/XeexQglyYIa/cBJzXKrIY1hxk
IGLKVXshbptLHBViRkqet9RsKpXNDiruleS15wE/Le6PADMDAN3AP0J5LM7SMm8geWoamheijPI/
MpAd3H14qXRyeyz/mye2ECo1S2Rf11ObSfkGzfxxs1GbwBnEe8H0+ymcleOw8zDZVHmTtOC3NsHQ
btgzCEr/5N2WHQdISCrsTo9AJ/uWsgpssYFAritdQ8RiwYKa7XPsPundzno8R2Cbg4GdR1r18B+9
QsgioXnAa0e8xG2g4B4aKctPboBx5woj0GHYNnKh+BZvT+K+o9596edQx5cOWLD+/Wz1qr/W9U/w
/F9LQ+Cs6lbC01VvhcgKkLsMrBZ11k2f0QB/mXQYQgxcb9ceJEe2xOF0AXLX2ArFb24J41dIZvXr
MbKG3ZhfDp3L2UYXhLlhx2Bdf9k2J49SfejthdkqYaQ1sPYXtrarxx5z6AQ6pSdUVktBeih5QeCj
YqsnK2A2zdYackADXUxHs9ddwn8gZ8mm7q/g0tRyJaGE5fiV9Eloedp2qjLsa1v7ooMj1uR+A6ds
OFpuPZzWRmW3j1Kj4xYZp/OexgoUjIvfL5SXX/fZYp8/Tq3fcAQ7Xotumywh5ne6wIB7WmAINOKT
kkIfYA9bj3jSyL+1PjF/5mKFeY+TDKzj7lNO3dnJQ0Gb1w/eS3L9/r0zH7Rq7dMdMCNnPaJX5Rte
Ow1340exovgpjF1LfSoNFa0Fe7jW/AFP4LXCM7CYc3uYDa4POt0d5JRbEmIV1eyRnmFREDH7Vc6f
sCY13SzUaijiJLGZtd+tfmrPxLi5c+ppbSYsyps0iSlVwMewHhf+e1G/ec1Nv49/RbX13F6vN/0E
L5xfarESu+bQbhQHKXvoOmxTzvyMtFY2q8JVYOc9SSO5crRTvqKHrcg0laAfV9fMsI+QTjtrOJmU
XrT/AOpccnJcHqsSpJjKdKGv8UlsE2sWj25HsnqP/feq5uOYKuyjxrdrzpKuIRF/lyXFUr85ul56
wRZBj9aSS0lz0WFymEOAa+1VQQ5pANwhikK5vEb+SW+7CDZOpGwxN8FoQuG2j/yg8jjY6UHFEgVO
hMwkDdY4qlypyOywDdBbyZ69+sysoBswzXUvKjTDPZ8DXraXimMEf1r3SvocKuuvBm+czzR1kfcy
9Pxvvx4esHeobaO9QGK50GQOw4OH62ION83+r909ziZXNgQorO2hDl227XvDMmX13B281LW8fPAS
w9Chclh/urGobzijgCK0AL+xZNJ0RDbBc6hdTopanrDVCdDhsYNHib4+5fg5Lr3Mc3YM4sOu14Td
d2NfQU291niuhK60adQg+sa+jXEX5RzJS/sK4vB3x4T5GiVBYxil1AWIsuYh5upP/QJ8qJsrcXdt
6/Zg2d8E3Xpi8UYd/Z8kImc7f1U+EWHyNBfe2PxYh4A45jJJQWAXOKti1Kg6CLAA7fa3yl8/5GL/
uQcq+1xT9ox3+PGPdyUxwUbo7WGxWTgphmE/aS30y2u0ypm8Efgp5f1bn8MGE46heP4F20QGRt5b
IxmLop8cMP86v6dv8xwppWLmIBBodaXU2966RNuh3WF7oH56xa1/Rzc2m1wRynC0MPwfPrNZvZ4/
anK+6z8SxMEQnm20Reuy497q4BjFoynkPKLl+ftLZZlVCEY/9BfnCrjfXFtWYMgq+b3tYBxaOzZ/
lxqIdcoVpW2Zxm5PRHV5H9MWOj9NmX8zwQMNFcFbvU/nm+K/tfgbIjGStyN5zPCaMMqBwOpFktL0
+5jPBCTCbiLJ4NzmjHaqymWibaGMsP18ZEHapW4wDX7xWnPWaGNTREgQ26DDt8rC1jOz94A4pugg
/WeLutxhMB8DuWnezpC2Qwx7y9fYkWwzgsTcpO7OrvPk9rzP0YKxxZJe1ddLaJt/929SHxQ1vEFW
KuI86GR2nduRuhaq783Xs9PXTpSKsPzs/KbiCtDyDrcEUGmLvlyQ+44bnG8+ANSc2zt0u1tyui8g
3a2se7VUXCRVKdbaMGUwAEYXr6mCemmxL6Krx4QKzpocuhtZRGCWa37CcwVeh7yONLa2rQ80spi8
pjZxHg4lv4S0o3YrL3F+AzkXhiFrwevuQvHZB6Wnw2v+n7/fX87W3wWzu9Cs6IVTNpbA0dAkOZVL
5ix1bwZx80+hQnssIZqklPBKposn+BGcnRYcmFnqvQFuv5lNpl2uWSpBw+UkszW4NQvV5H3knNvE
ho/iP6K8slektQYapBSz7AHL/0teyq56rNvA2IiAYoT56F7+ksq8RZ9TGgTMryqyPfxPfQUJVzds
8tskPp05rBfGWO2AiTc5dg3nnvuZhWC3oGKgLn3IOTz+Dkcp2sff1s4KsQctDfQbuZVwTneaP9UL
ZuM2P2XJ77V7dns+jyaT6dnOW02LzkKqbXTc3yiUOexbSTQvgFEyQa9AnPWm5WQdaTX6NW1R/cBF
+TkMunWSfK49LZVZ30Ey8pNgy4QM0PTO+OVpDqs894TmG0h4kC84cyC0/Av+EHDBVouTLrlfc8Pn
4M/nMKwTu5PTDRgL1kmSKbr6lOZM5Mbi3AN/D2pGlyj4d9myK4tU27xyD45HBEw2lFjpHAZDQfRP
BExyoWeh74KLSk/k7v9GKYt05LnsyB9/PrrX+Hw0UoGp+OWTUWHM36EfJEb33IEYrgtGGRpdHxrW
azb4UgLv/OIPRnY9J47EDUTmbgRHa9y7xzICxFWOY0Bkb71TRYt0bgl3wjgZgawdqa/94og2c5my
NhBMSAMKK1jcs5zkJdQBexpo9gEff1BkEllWOoHlh5OjXvGiLaJRKwRAuEchH4OzIUfL0XZ/4r7C
c5EMjBBIpHtl776PQDP90GzNuTNRMYjiTPoKCIYBsYS9kQxGip1eS0Y5lUx+Do9g1BYcvMLNRHvA
DyX/NAok6Bn94kNQ05LclrBHrXIbzHkF0BU8nEoFsV7O3VuKJyeyHlzae772uyaxRx3JCYNeOCVK
DD+P8NCWsBEVMOvmD+yUg6a1UY/XOvEscVEJtBwHM70jmfd4iV4HuwFULzohVZA/UXw55IWbBcu3
uq/7zh8yC2z07E5A126qDKO0mSyFq964Sa/UymfZCM1U+6Lc+EEQlvXyTcGyp8Y3o/RWEgcO4DJ+
K9ghMFxIacyA5Og1xIdcQOzPiN1x6ZuQfS7EzsL5CXFPsnD3Y2p1zSH08JSQ3pv+fjS0tRXT8xaJ
qYCmNvSIys+ce0/FsprpEZ9oWtJNiEA4iOtM01qh4tST9hzdmIhdKB4d4l+IpkWTMAKRqPhh6Idq
SdeG3z2nw6kdHa4kgLaU52VknNngjhZZyFMDDMnDlvDZnYvs7F3sX0tM5xa6c2gehbGom4Ps3gZN
rL7qBqtngFi5WoZQp4cya/qUwDzhT4w9vfBCbSzDFB2m9s8ueJjhvOJYsrIGNd3JMWv3KrSBeVqm
4Rw5xCyqiLr6bx8nGIA4ZDs+CyfS3ctVJ/+pcrrMl9bvd57e8tkbfExGvY0hlIxB/B8NSNED5XyD
uoXgHlbNaUttaOzazfM0cULmAx1t2p5iburuA8cQs7wk32oBamSxlT0bYK4FLmP2fCokJLivm4Rs
mOsFw7lXUwoFToRjLhm4xHQojrSXl8IVk0BgClhXwC5lrGH4PhrruputNhqoWAWPzCP0bUDrNxC/
6aiuNUTQYWG/4SuphzzNTQwXe4yNnAzULwewdhH7eCAg6WrRP9wPF4huDd9A7rsJoUmO49UqgX8V
wBteFHKxCxnhFzbTl/GkxhLx6xZXTHsWElW442tOZT6p2qP4kzbwBfWIxwIV4kjLZnt34mhB0vyt
SiHSrr00TPh7wPRcgklBZAbML19z5qjxzMGeEgbvVdPhXSDgZlyyPXxki9J+Af0ewXfgpRB5V3qk
ujNeu/vw8BHpWg5214ealM3K/tkXf/ENh6iFeufhMTAe4r9/E8W5r/pA+9TPbzNEhk+8LhOH/6eP
/Sq3sTBH1eehfqutizPR8XZl5+w5lr46PLlFF+f1lFzyKNgEQIVfDS7mimABj135HFzqzrdOzZ/C
hlCZkueaw1cD7webt6SWFZCl9VlyNaXtFwkch2t+2IKjUoGwf6tWVTbw16gt93t+HJ24qgvENEVh
7hGU6mx+JE4ms0zmYEu1EK8HN3GTm/I+40iX6rxDIWAMXQo5HJ48WAXY9mpQAoV3AlV/8Hldjncw
B7AUctx53/OYcU8bvUBVXol4Y4QrRNruDz8Uw8eujmgWWKr4esi2Q3xy+8/0XnjL6d0Y33LfyIBY
57V4Y3DdDrfWm8V3Qeujqwk06MVINplfaAidjsDwX68WQkvhbaCdixUmA2IxvsgCycTSZmJ6oFxh
haene5b86dae5ipDSimgKLNthCKj8esJgeOtCjWPlaDpkYiAkL+k/si3zDTCcvLfYkFp1lr1dKmC
nSuKq1TRuonUdoGX1qvzc1v+JnWJC5y+xFix9W7nnLNNLwAAp5qPTh1qIKG/ZhOeBxgkkguch05p
9UaDkcSHVeCobeAKFXosyy0ugQQUQ4/qe792BrhC+7Sf1hXAvM3e/BchYl/Yqm02ZL2WSsXzTIgr
E6IqXDgMjC778w9+DaEjQtP9I0dxATouCqwZFDtrQkFqPh+kPvpSPr8nZo39W6w1kMLZtMspKuzV
plX4rpazo2YP5hdYTfx6LuDTVYNqESsfPgpeIcwPCOidC5r8dxnbXS8IJbs45L5F0bnj2eFrzV9j
1AQwl4LUK+nNwqa+Yo7bYGsq9AOaXU84RNRnPbav8M/KnjMXwF5zfkxqPs7fUrhROx50SvXM0YUO
v7YdXM9KrHIdaagIaiRK6ciV5WIxUEQyxKqugoZSzLFmEncUuTgPnNDG2hxF9fstV0Z9OYZ3Fas1
E7qFDgIO4ZbLA/RcFTOf8JUFxsGLZJej+Kb1hp850jRHgmmijNCWP/0Pet2i5+U89ImoMvSIFJUU
YlvNjdQkB18pE9D13lBkBoMDvAJ87UUTUCCONl0cgaTeRTfCEAG1+YrXnQbXCFAEndT1KBaWQqqn
Bves/FFy52ljnySPoUDAQ/SaR1hZkak6r32P9sl3ulbX5ALvJgZXmGA0bQF4TeLJ1FFg/MbsC9cd
AUjpM2UWk8JLfX9Pk9Fdktfo9vePtDPDPKmJz/F1+wzQiJRuZKka367YDXJSIMekfEPrRVTvZk18
cXvK8hr6KRljmkeLx+lKpI3iFl6aVHit3zL4iJ8von72mMV+GyXV0pW5D6IlYfZW4aqkVGc+qCQ7
OaHdNCl4bRoHn8bOLWfOUkv46LgrTZQ16uA8Z0vM070fyup0nGQrYptPcH3Jp+HuPBhO3MnZTXkS
835XUANZbVuOKzRAoc+UJbAdQG7zTo3MsIK6mFwf31UuhNa5o4Rt9IJoUoMeXkW2tiq3/uqEku25
cf47ZpQ5/47dFfcCtyB3Bald0rbX0H+eskvrxEZq8GQIhEjIZ95wkLkoXJX7bYfR9kWal8IL3r2z
uE789lMsikCBwq0eMgXZw0R7VpqgoemOJbrfnAfJ4DuZQqvZE+qpoh7jV2/ztUFTgd5vXTn+0gG8
sYcxma9fL7Nh1JgB6tELso0HANvW11zhWlIS7yIZu4CErRgAwCXiNjd7Vvc80bF9bOfYWBzwrgWh
48BtNI9Y8ButfigHIVe931IAtCTNbxy+p6X3wullLWNh7Z8CMxtxZ5HzQ8sUpHR27fCjd4+Df0r2
M382z8WAvr5DABE3hgyJo9kgx4xDQFd0qni8b927r1U0bITzrg+2pHcFBlyhVDFErQTFkc/yKUlV
0yPEsu1BNvHhy3GdPJAWRn/E2mrU8Nr2MxJRR83KU7ET8z7D9uO6ZJvG7b3R517U7H3cGiBG2mfH
dm6nYIhBOLd6W/8/gFI+WJUiIWNF8E3uOvWqO0AcFu5krA7DuDVRRp4IKK6ZMZHMfOMAScUOBKeX
XFYqKIQOm43WW57jLEwM5Xz21maOgXR1YJPTy34CeOQmC7ql1wAp/zjLG06WrEMST/xHAVe+XKU1
wq2IFHTB0RMWYhudRuotOEI5uBNQRXL3gYFINReYzO1UlfEEH8kE2ZB2+4EhZoXtwHJj/lKR2Whl
zKcycwDq9UpmN+dX+5L8eSdpPVkEsnD+ldyPkG14dxCKkzDwrAOBgrwEy2vPwv1XNAqQLHso7a6W
2w1qe0lvblf78+PSPV8w1vlj4dSzW5HKQizvBcmfTT+Pyw+NfshjWQs4PaIK++ooIptJZvGQEU3f
hype1luFU6P6FNG8JKSTqHoSj4SvdsG+vTOL1U43hyL/qW4L/qFTQvb4nC8rcCWa20J/7cGtVmlb
PN+RwEyxuth8UuujKX/2Wbm/3qKth+t88cXvU/1EpHoaei0B0jT/uKoQQnrP6pv9Mwrpf76Vf5oM
nHPnvquOtvmqWD9rEdTcNqW8Z7VOmATU/ZpWOD0lQhje+OEl0qZw3GRWCpb3mRz7DNOSfdSErddY
6SVgK6mHN7YcGNw/0didXFudgrVZyj3E5vyk66Ptx5JNi1W8eJ/CPplAQwXNelYhsu5bnjs4bBtz
+SKqAw9hWAssx+YlVkGxYOZ19OS2v/6z5wVrAvRpbL3qpVsOm//5kxgeqE+oTXWjK5gCAhZ+jy64
xZ/fEv4/np82bdxsQKYZQVXXeP497PwHvyvGq5Q2vCiyuXT/CL6omJBMc5VkhK3v8Lk/d1KnCCWr
gZkn6IViVc1MSH7/wHQwb96wBTwTzYbSYzZVIVZ0FJnRBEIJ4NIwukMgHOFpLCYsw2TVwGRvG/9A
KMUsoKSeYhyjFw9gVzHzMVPmkL1T0z4XiZeSzC7HkcleN72jI0CEr4A+UNk3rf3Ag1mTszhaXt/f
dXw/HcFqtQCAqtkkOUNkIo6jOPlh2eABJOMwpTCZeS/tYXqFlg7rYHDNbCWxWBaACYzx77Np7RGX
r0dbagp3c3fXLkAe3FpQ9yLqoNHNxgayCHBfy9rmQ0XqYEp8E02PrEAsmxMVh+WRhHJZCEWnUKtj
cpx11k2UDUXYXbvg1anTvglumLqK2VzS65m/hVMJ6ndCi8X49SgFUU+M0SWlyJMUp/yA/AjVyfDE
1HKM9VazWKUVZSVmS5H2JB5KnJ0E7uqxOYB1GQIKhY9aSVAGLJs1O3eFBRp6/2ROtiY5Po2zCRz3
TLYAF1uMKY+xa60ySybMg2WIz+b44CGwP+HC1sqUeOV3UDsJ2ExRpEOxPsA9ypAxjsULQS+60I76
HDBxF0f4jfxyLku5qlzRE/kIzvs7Aqru2hMjSXEnulxC+y5Muok5Qgx4ArazV2TllhmpJU+60Wbg
rkX4HPo2YBJqbP1uytRkYO3JWurEFq202EZGn6Dt55Ehd4LHDyMcyBtYT7xN5fyMetVP1TvDFPLT
Evr5W7NKxPEy7ItWfVlyvTLgc5JQtyRLbqnICCkpxXJ0d3zhAC2rvVR/Rfffz89bAm5H/CsWk6V4
SmLiEj7oLz4FaFAtj7AIlx80UYrVZy+v3ioIK2VjcRk88SY7OemwHe8bMtt7Et8KymGy8nkeJnKd
IMMgB+nMyl7ztsiS6M6TzvkIY86PrUxEmshSr2FHfHBPkPRqOgHYdAR/o8vXI7JV10AUoa61gciF
c6tZkA4TOj5cSwA1yWLOrdreRgdYm8IXJjX6Cvf5LnBtk80nb8OFjIi1+yBSmAEOm7FnwTu9b1yf
jXX3bz/acmlA4M+xUVMTruAunznmKlCLzBnVg2G4OubfLzhsjJVZjKb7GycbUglm4pbgxGe+hNol
1Yet3XN3QTv236iuFZHfofJSgG89Wh5hTpEGhRDOPTOIco0/6JpS3XZvv+B7a56i2wAH1aRexuQY
vRr78UBXL/qfWitZSljjVvVWYVI6JnEr6tDcLsNIijzZHiFIFiRaK4dnPc7wT+QhMWifc9huvinI
ZvL4t9vae1DX1Bak9prewXHxqrCe8WmCykdnOW9rATKpP0mZWrsIeH5GNyiAoyNr/qgcr4JM+qWy
ladXRfQvntR/ewP8fbiaDu31bPbB911dxIVw+Dm/egDuWWJ811fxKX0o9ecr2D4gyueEM8Glf/XF
vdtzcAcBg0F/N5U5DQ+3nYnKgeuZ8bkfrsrZepzoS6LVVEQvnPHE8TCwv10hrfuoMipsI7/rmH70
4XPeXZbQ1XiXX9RwK1wM2Lv6R6WJoYJTEFZ2+739s9zntRHpTPGIOOGClaVSt7v8m7SMjxdDImQ6
fRtvHB0ZZoWbFb2UOwWdlCV0omszTApCs9MEyP5I4Zbnqrs0dwEvzMnxnYFuEnUtF6yLZSgBRi4N
2j2SctZ+6qwLDyGcoF4Wr1dy8thdsN/FdCQ62OYPeteIlMuBINisfa6e2Dx8Z2sgeLGFtVK8GsbT
crQlPZIy9DmGBEW0ubU7HOecasybXwRlko6p1NSsTLf7zAU/z8iDLC4hCg24nnwDPlOoJq6n0DjV
LKai6HOVGUKCqBF5fZdifcTUG7/tY6TFq6xk7aPRgHbKUQ8Q+4tJt+fd13Du9FX2SwpzMdPbIkWx
w95QDawIldFSHfJ702aH4DI8QQkjk1YJahW1DQWWNI2AMe9mzp5wx8Oti9Oc0AGvf9qWzh6BwaUt
KoNH80FWnWNv1K30K5ciwW1jYXEx00Dogv+w8pbJuprxhUsgraW0JNKPrhzHJI6p+7zJTUQcl3ad
e5RENvYl+o3G9BZWP1qunCbCUu15nw73Q3d8hbkfaDuniCEboXMvzK7yuiXMOO3Dnm7qMD1nipyl
l8VEjOJXSmVpQbYm3d7qyvHmLZqM6U5yOlxr6W/DkzN7+h2Kwy3hmNxDmYI9t3qYFJeRDSoVu9rN
hPNTKTUNxhMZp+F2uMG9NXxrlRnjo9rGw1ckEECptjXJtFn8D+8woy6OiHt/qEc0FwW8tY1UEucE
+80PZ9sKGOXMONcRa4LLbyVnbQIyT9L81uCRC7XLumgCn1hd1I41JhZI5Vi2ptNqV8Ese08lpLjk
QeUohPTuF54QHANUhvay79bVpvn7RCk0sE+z8F/qV8pk7KIA6VoIp+ue8cQOYvn0hMtp+mLVkFUe
axzc1BvAT9lSHef2UDHkQGelxmibJSGkj3/ceiwQc2mvouUOX3U6+CIz+z4knndMC95veXhAMPC5
bIzg0gfATdLc+D/VCs1C3CasoQUa7hpvhb1AUYDTFTw0iDZm4EMwLesyXIvkFmozi6bBysoDPoKx
p93H3xDpxmBY0jh2NvY/yYt1nmIyIq5oJ4UAQeKFoGW7wZpm75URgDz6PQNwcONZ3piu0JxDjp4a
45m/BdP5POk6RyAE90yoTG1cYUMmV/61Q0TcEwkoi5gDm7sPHcTxf9jYC3VGGfBWTQwZG+97BLvu
f9wIqJKZPOH3+0bH3QLw4LeE+NYufF956owNyZQahOiHtOJetSKQUKGvAWNpzNzNwjYDSndgd0Y0
wAlxSrwoKBI4mjdlG6Ap906iha8KZclCWuMWuGEAO3UakR6n4Swd/l3NnaPDqqK1QrgoGfNXil5M
Qlx/EXJnLLW09+1rCIH1p9FXaP338W9ZRqLlJ4SrmvWgIzyQMFVdJ6Y6FrAMIwhZIg8/IZLD+zyR
57WWgmM2B4fWKkzHF/rOwR1pCkKtxLkWWmmIdZzuI5t6QlUKGmHp1SF5PFv/p1pshaJJCEr1MQ9L
QhBjbTIGHVB3PBBQWnsY/e9HQMLYN/RJc2h3noTZX857+WiM/N7fIinUY/pqKTeHYebx2JfmgVlS
ysuv74HC81W3uatFRw5GTH/AkmioynO3p0sS7KhiUJXSEbu74UXanWksxQzmWr53j0TGw6KBLTXn
3UiyNtOjmO6o6p1nZ5HhsgtVMyDUu/dmln3Yc58dlMksimOQhq1742QhRv5nwLV1Ooo14r+lwSiO
QLHGhCENGEemsxVee8iOFe5RC99ELNDfv9iTPzTR4yi62KYGgQnAPTB/hnFiZf7GH/VIgi2I2S4L
+7nldFrISmaal+czv4KIltUq+SuSSSZlPaKNQ8owcE2hKED77MnVHH01z4zgBzGxXtJE5nN3nQ9h
JgGuZXoE5Dmi3kFN/vbGlJU+TdjgoiGDx01pglvTIWbmxazXZ6LM5LVUIucPbWqmIzYltLTs2H9Q
PQRkZxgHTpsIV4i0oTQb59OdMuPRD0hLNxEDB7Uq/l2O4w0rICMbIWPgMaYSknJH5EN6ApDRFBpB
7F7+2WDgdmov8Dmlf6AFJ0cBV2AgWFphhQ6rMLyAzZTIEiniQNCXT/k4tWdRNk4tqywA9AAxUd79
GS4gEPYEG+fB7iZ3zPgFAB0fMXChOFzYjTCI7pvpi56J+Ol3fBSe5v/fbAXqtDH8rFopcrxUL94y
ZgnGK151VosJ48noyuSkFQmcpQ2qKzfLEckx5+KDu6p5MofiZp836wsWZRP3+HmphZiYDDPbs6z3
BNsRKKm/jSaLlNaBc8CXIMKvJNf03yYY4luLUqQWl5nc4I63bAezFTo2xKyf/TUUnRdZcurGsRMk
icNmO4frAI/+J7UyVEEBf4zNkUJQ7ZeY/rqtQF4YCJxwj3gohAHb6MrkNCdZd7mYEbShwgTZr14N
Gx4FmpKd+AwPKfHF8j40sHVQVG6qR78nPT49JgdC1ird3al8FLdif18pN9fOiOEl7mytG6kloQOc
POqEQxeHnx+FkDh4HLcQHJAu0qxa+oc4Sh5cWBF7kbH3801D9x2e2QfnIr/UIk5AWVErmGyh/fM+
BwF0gLZx/myh0HIFBN0haFX7UTWQT0MQP2AiwhJZdr46iUdPDGB5jWoFQN1NyhzKhn5hXXYYAiFf
MDJA5jxxVK4RM3PDE3+Xk5cBV50Pnt25AO3EwyF+sGnXz1l1QOKYjwV1ox9YsVKedTU/VIePC3pw
Uzs7jlGHxnl8E8v6hSXR5KsPmc6hNHUnHXPDDuPcUDt50ZEoda+Nd+nNvnJH1odQNOxvP7iv3W9T
seO+GbC09j4tP/XyiSN9WdiTVKY3pSOGJLwEUm4I2INPtDeGZy5y5BroPbUGPgFBx+xA0f3HIGQp
nSo4X9td3+CBI+ZAS6RDNGsn82wmcJaP0mPg2B+ksX1RYbQjSpQw3Wo/6vqFM1ej1/Z9Isu5I3Td
FgrjAZr1vrYVyBeWVpmMLEMSH8ohv1FwCBUW6eHSYTr67sTpFG5+imBFJ4Kt8SKIenQRTm+EyQTa
VXIcJ3b51NpB4IlNWXY88+7Ha8Huxw+gVSbBi18ecnFmBNVn8SworOs1Rdtpx3ECA1bBExWzcd/n
fyCwK8h3LiVBwuPSeBJliH/jnUy/oRWk8gKzIulPbsJwu0Ji/RVBoHBlXW1tR0rEK9RDlWuj8RUs
HaY3ssBa7IbYrcIrcLwUB7YEAHTIXdGNyRV/kO+twHF7kJqKzC7kxafpD6DDydQBaZvTYVuTSQqJ
SWcvUdGxHMig3ZkURxqd4V8ewWHPmtSo70L8NSGwAs2CyNa74dThEtxEYiahbmBcvG8MahiFK6vR
q7ZkaQy4M2lTgkIRgNDYcgHGcH6hkUBKGOQ+jlsBD1Wul1fKEZ2X0PxB41EX/9TvfXtlB6G4GP/u
GmlfaOyc3BcfQPzGKxf5k/xpAJN74rqjtsXPNGeV9sQJiuzwbJA3capkeOOzHbl4xPGFEr7n7xt6
Cuzbjx1hLzPQ0IgWgiad2dM5DkiJg9gpneDtWnxTCh/LfgmNcKC/35+Ue6/ydQZFLm6SSuZ1wEf4
Tl6BI9UjddX/CYe5phlQHdo181SUT9+v/Yb0WOKgi6x+NUB0Hbt1qgWZhtziON0HRdQFABz+f4ax
1k+7i1JDzlD+B1DHO23dtNpE4TyTXfyPLa25oT+WxAxY489tFBcHxvocEYCl4hTiMolumopNG1uc
uMSSTE9TSZv92XVS2QQik87SumoZRQ/RxWio6MZ92lSxcyNdO++w8knwnLFxeHh+xaX+9AzjpNvj
1xCUgrumnBFlzkVoDFx4kRp5RUdIl0VlpZciTWbKPoN1m1fuIlyLs7Vbvkf+wboPHmBLuvsySLyg
OEGEfufunPvz8LL8Hnj4nD7XiOZ8TEmLr8xT7SqnUNkfm/lU7XkXJvLStAQWao5sPWnYXd4mVyom
wdbTiPZ3l5Ncp518e9FBtv8/wOAoOtRV12WJroW/M3A2xOBrqneZlwgiM5O4kOARdplH1oKP0COJ
qLcPs7AID1PUha2HNysiQLvOUTOoKRsaVEkCHQNcmlozeyZhhhO6DAYY/aqchQJ9DF+BJP4N0vcC
IQ9EiyiJfY8r0SUSSu6dyqiP2w8ROk9TCmAB73Y897dkoN+jHPd34NkUuWp4HuszWpNFZ+nfEITS
ugOtcDNfXeGHl4CYcvQWsYyTeOdOt4iSsB7a34HCM6xpMPL5PVe5xnTdkKJ521xDPZZB3BAVArNd
xsRF0HilnQJnv5HBO1fhRPgrNa46E5Yoz7WoNG7wVs3KJ6vxwbkPR5uAd4b8sgEyTjqZzMyCvu33
EbM2JTFmkyV8GmAi4igtlpvAFqlAcw5Ko4E29QVA4IPrVPpXowz/kyohqa3/HVfa8eu92sRyyY8F
K1TtIFzthKvAFuerQlmBu+DeQ32sA4zt/K4WhLmotPlGWtQi3FAD5MqpX8MUVYYMMGfD5jD08jpr
3hsVUxekOMepmhqNHbs8qxYdMIJCvZxnm3Ej0fQ5QNvmPqTed1lwRdJc3i4eonM09aimhnqJ+seG
sM9hdfRfxdqc1D1czEGv2hB+GjJUDwrrm9hlSeBEA0thCgyV92p4E4wFHHg6XfycDVvT7OaZOPm3
eOQY/kARdOoAg9X90zGwJIgc3aD3zooVhqzWoEWs8VDOYoQRQgpkUnxqmvCJPbxq8xj+qg3hDdkj
RJbGgdRssEQbEGqmD00uE2DT2I9Yqyrz0/4JB5M7c4GZl/wGDcY2NvyknjQUHgTz5ZKmx5nqYEDU
QBHfuxeNUmNyIdTJPwhz60cMubmV34riCDXnKQhQ9W+WMLTwaWaWObRYNi3qP9ANr7vw+LKGnLAu
xlPYoUIhX0z/U90DHgDfKK8cAcpYf1Ce/ExmF9mUJOF+VWIp8XSk+FBRcvSyGc0mQ0Zha+IJdEhu
kf+d2AveIegcb5sEYRHbUEFsodICXTTRq/UMQQr25fcXbKRuC6aZgqFeh/E7f9iNhcbivc8zyk8x
qUIfMAvLatBAzkLUa8+0lhsgDLOFL7flpKxIxaYjr6UEC1aHmeK/14O5wY+h6JZy9CGT+FHEkKdt
uAMS24FxJ3PQdFWcCahp2noUtTY62CdGBFxIZlh6PxHk2NTyUYSxqgKH1xRKHQnnpyfNFrFLbcMq
bfW6W3PrrC6QBWfHI7za5qD+FLbBLfu0qiIZig4WpDUxAJGMZx32Y2AFsIKhJ6zw4T94iROSVVsw
nFpDjyVKZHXi4ultN6jVE9K8PWad6NIi7egXP4x7KCAGzCY3wbHjtbRvDnCRs7QnSxvQem/5bV3O
Yjbw3tZOkc3jgQJABF6BXXgcQ1FTHd+G2Bpa2rSMM6kKIUFTT+smfh32WEj+tRQuEQECSftC0Zae
hsMsgHZrj2Sq/pYFCe99zws8GspXI8VGCsboKhbl5VuLLNucYkh3L0Zr6YCU4NhqA2h+/3fdUYg3
uUhwS+XxYajD+dYr6t80+4lsetzmWIRj8HmZVFlLg9nSK23/uvvZmrSqvuGSVPGWdvuwC4nD6/cX
1NUI7rvY+Px89aKQQf4ysMqA14gnNrxrSwW8566uLT4oTlSGViU9DnW+7ik2wn4xbdhJDKhtc/EC
dGHoQU9yUWHjdGbcUkCGwgnEYBjnnOTN18oP2M8xVJXLrdGwk5V1kRUsdD9Kw4KDJeaLW893RYM2
+7oQWOunQHtQOr4XwmF3l3fhz7GpdYosDsUT5iApge9HSCb1V/pqK3yWmCN/J63ptEbi9swdddyn
dyCbuzjQNZyE8vUfuudhHlqhKplKqAmpC0mH8t81XQW5B/aRNv1+hLqBjbpFf+kvqZ7qWfoSHGxm
vNW4ALLgD402eYfJyBd8AZlsUxlfuMmsHFnHiVKvcc3XHGprHzsDnQEJbLxaMjB7Kp5Kjf8y5XhB
zjwaOO941FnbMJbLM5gSl0otfT+005zF5LxzveikoC1CvGQAOuyiukLv4759Flpg/j7uPd0h+WKJ
x/xZUYWXZ7uG2greqyESlTEgJzi4MAp4l4aIFlu1hgbapB2IvM9/I+lNvjTfpJyfEKOJOOENQheV
kjDvEt9iTCIEcIgGoCDE5wV7zRvIL4F4wX6d52klbZHpOqyvIFu23ietRsUT2ppR7TTWP8xd7jou
ELpSfiU7b7w9SDviphpOtz0P63VFsA4YpLyOEcuC00Ie9uCTHpy2zgH99MtsDP+mGQGet3ABqcL9
hjgcmYJ+bSrCnOaoe/2Xlo4UfqyRY6UZgNAqNrXoYigCuc3Cv0eq2vWftjFGrsL3ubAIaL/d7VWM
+HZgM4R8ZZCsuSph/vyBZLgwOi39hyXAcyfyfY7DlbVviFHjZBtBW5wtVxo9rzmNIGnIAKaXsbZk
uNBbYfffSpnhK5hL9UR/AIsP8FgEUfaIreij0+gOBI2QH71wqzZw54DItApTumLp6o0c5RyENIru
CUoCy8AS0jeI7TGNCK7rv+7zy+X9Pz9KWqwk3g9BmxsXs63+Vdc+i2+0U+lk8Ctyn8Jy5gCZ0qmh
iMCeSp3dOuqP5QR2zVPlw+xybO8KbiOnzbMLqdZ0xErYKhqG2lD4Rz8+oesKlqFlaIz+rLQDBxNE
Uv6RN3AwPmp23n+GAprwjQNX84J9KUh9ITyh0ybgTIfbWYqPj+vO4MBGj48UhzRyo38u1+mG7o7P
VxpivXYwl/Yi7J2cuFb79OEuFsD5J61xLxu04yAbgZkt21LkkjqaloIkW4IuR3AK/o3Vv0AvtMV7
al5oDq5qhALQeYnqh/OY0MfX6yEm0MrHAFEbs64PlWL8Ed6WrchpgtBt/rpL26C6XLPA89ezzkfz
OrwZ07yh6Fz5dqQfzkEl3/FVm6RoEpTfzFTMZciEIVzdiU/59WG3GQLG/voNigRwXfAEjyDpkCVC
kRH5B5a53PlSK29iB8BqoWhjQyXKCJvZYRnCXCdjF40F9VRICPWMl9wzHZKxj5t/rHT54myFNvgk
8eAHgGeGBbyo+Zm6QceaLOc44cOmTB7ayAObro2ix+g29ZaH+M8vyIDoICTtFxY+zahyJUK1wJcM
EIuCoa20dVBkaCxCBL16Qd6X3ejuJRHVoRVF+j2ijr+JeBy2yZ0EVqMzI8BJW1OLJilL9u9By2J1
Z7/SeCHYovjf6VG8q3xOhbJ4EaKqKKSb9KuLyIIx0uOeDH/RvHFHSCVXXtthzJgtg2a2oAsTDlEZ
39nD9UJmlnoJRKHxhqTwvMXJQOeX7la4q9eqdE7s4AFNrkUFJ3UkzQyIAE4vkmK3di+Ek8xBO6jM
nWiI2wcVIst1ejWfV4mbIfVnt+uYBlK9E7ng2V5zck3XmCeqjhGRUO16WmRt18n2uORWrYVFFsI/
mSvFaAboLsT6ubZJH0hvTNRJAB59YypVyX9WkoKqdI7TxUkmy8v2PNGxXF5o8jdpfL7+OqYRh6d6
eXwd2RDwgN8A7p7k6J93KyVnUKmdteL7MgZIaBXoZCmJhqKkN7pdiPLuJqyZtO4asj2YPSvwcUIo
TN/2NMWeq2hmtn3M7J2ZJl3loQsiAZVNeTnZCMypgHdUZeYlBqWquzC0BOtkjgdDu9aKPXckKJrV
t2q+FHIWKA84ks+uPN0pKTjM0jeTn/d3jfHkoXDUYaEn9NdXP8S6HmtH6EHW5g/g7DOyDilFPJat
puO7HWzVZswPvRSLQGi5AvLdSu7Gp5CEn8f+Sp4dT9033l9KJoAVjwLZgn5snm8sTfSeGTyxApr1
qCVBWFSHJq+3rB8kEM2CAppfynlQB/JDzqXvGs7YugrX1ufd3cHaSq77ZLYb6LspCkC7b5z81SBU
+Ce3fcw43YG0FuGUZlZwGkZ3vbFyNU3/DxNJXGNLEk3rlujtsWB+OwGg09pYc1gHqoZ5uepIXDVF
yXKG0bzrqNGq/5XzOakvUkv11OKvyH9RnVLhm1Bg9IF24Nc6YfWgb1Hbu13Dj3MFlMvxkpyxZzmD
mTgQNTXGvQVIBWTw9qvwA1FbCcy6CIOO7YRRKmTNY3mpXLusJOa+heq1y6U6UESRnd4c0FdBBU2U
A4DwmMTdYIKWRh8rawxI7l4pvouy3ORPcBUpwzziu10qm9o19hdQkngjwGNgordxp0ZYo/0OJ9RH
lUKVdSo7pmXYxHjB6cBRSV+Pa0/8QWPY8ZL/E1FYyXElVFSvy365nmXDYHCA+jSOVa66Zr14eYq6
6fmuP52qpMsUPv299datrKQZXndjeoY0AmLQ+yQd0xUZyX1yXQY79yU5QvFK1j4g8L1gpfYjo92d
vsKTkjJlzVFO10lFjWLIPen689B74O/8dZhKnDLSNFgcq9e/lE4qfnW+4Y/DnqZ4scKd7hYc2+EH
YjM1oLTuHQp84Qf8n4LJcd80hTbwEbu5EVX6/YYY6PiGvPbITGB6/rNzBxdhFKOVKhJ+VOTlpjdG
I2qtPNYr8oyrqciam91gJrt3zL/cTjXI17U5HgxtlbmfghqRVITtCeYG49V4HXnFkQal2KX3Pf3P
sRF1TRpApTqGWF3PgsRQlAU/R5Z9Vhzaa3XdQgQDJunEO7e4tra2tUMeT6bqKlE8eGfmrDO5vof6
kwjbNVQoWvGxhFweCTLLZs2hlg9n0oteL6Sq+7RD52lAAhJO981uuhCFq06pKGF9hxauLKk3yfuR
Zq5aeI73lNsFoFqZg5Yre0nvXfOFqNv3HHIkq/+aiZq3w2SzmO4hz1CIeV2n/QkyT1m1saOR4I2t
6WApYJ+tHXrICn8+6jpZvn+Opa+eJoLkMQEYQTFxsBLwt89D5ttrml2CBsStOTOrx8CYXQS96fCx
B53N3wQ/tbOdEefnw56kirkCtgjI/MoFkfwL9VfXHpznS0NvepFfDDICm3hqpwMZnnDtyeqr83BB
UYCoytNS64d6mLIRBQ9YdA0jVn0bnmqgCCAd0cKDtc38pdtb0jMMMBh6phKXsnhY2rRr2LQ4u9we
m7lZyhlTO38FA6OKnxd7/ZgtLFDvm7uAOOQNPFay9qu0+bCoxpEWo94NUIm3aoODbRt8KFhE8cZ/
eizywfZhEeYO/DNlG57IIsZYyPfTM83UfyZeEk2oo6EbajnjXKO4NIM+Af4g4EZM0Q+wWd3EpSZP
yBXb+M5A0Qi4JwSwhaEX23svJ1bGslpkJ65MLiNplkBohV0OyiMFjCKu5o+gBvQg6VqBJtP41pKe
7tKihHG6zpvWbD3+/L2VVloBD1ZbQAKDcdxVQ9hhn7ohhOEFq/VK/0zYtsF4lCcyi/ujJT0WLoYS
YdPQ6BbXgpxpxCXynHVxKD5ghwYya97p7lnlaYmmZZfr+QCEJ8jbbJTrIcwKlVb+MR7esgvhCkCK
8IiJWdfm+yjauZsIs6652uycrsg1Sya9pXvzAG2lAfOgc7eexiHu0hjgvDUbyh0Dp4sxjzUZMXku
ghAC989ozDBA7CfHSW5gpES7NVFWdXn7BewR4jGeBw58Cnn8d+iL/z776PSqtAtvFuMS+kQ8Y17X
yzDX0PkMv75uTHer11UNDdsIdtfFz62o/wdaRwt239OjabVxkR/Pzt4IuMBMioIY53QlSOqbz3re
6j7IjnBVRrxguTYDvtVo35wfbStZflvvFCzLd+zSFcratd0oW4C+ttZpUQVuNxJpbCqsDmUAhmVF
WRV/TEMs/kO9AMw3pfa2Nj+te0CreMrosa0Ac3Wt8ZRXgNjmocCMrJC6aMd5/b6XbYfbVLcfQ+GO
lztGCXJLzVPMv4RzN71oIg6DgE9GD4KYlncfKsZBRIPLS3fpYudLamkXaDw735NVzYjDGWfpltkQ
FKlEOCNId1ipcWJsYk3XaC+GAUQ7MKuOC+89P2eH4dFPpZTebT83d1160x2GlGtFe2Dxj+NcufRY
1gmdYmfcPOz0ABjOqdTCzSPJ1846GG5G/YnrTcMv82HU4OKY+rUjwsbIf4xGLaHcTPFgY5WVw+Pg
jEGWjMkc9E0g4Ea8Oc7b0RAT5GrdUdUKMR4fw72z0v6ImM5UYtwDOJxDYGUWyX65Q1+9lGSNtaBX
jmZictKjvlPpRWHcvxciG24IFX8nvgDSTpmUjRCbSxKmxStB4h2jmVcDk/RaERql3yA4r55SzBHt
pasI2wxWYnLbBfc0HoMVC1xp5LLmYvrrHUOwue1B1eIsKvHx3PbidLb9KMFZbS4E9tQOzuEKdTBS
yrOqQg/xHLNVLBm0d2GhqfRAKkQATvN0cBgdRgo2FRRKPfXyCRYqUnN30l9+Go3KiwJp/kvG0u3z
x6U3RmnRyUPNnU9f4JC5YDqcd0mdxLde0anh9NOdwY5rYmqxxhGESkp3NlmTAAlx+3joXUIcsCRE
AQNbzUfxWRQzMhAnFmmXM3/uyBLLs1aNSujVH5/1XE5x7y/IdnNAyowZlNey/6Wva6qJva2+jQoh
nuM0sM1vagL5WzLmLPkLMHVqNg04PJxSV6A/hup+XAGPPuT1C1PTjYWSUp11S7YYPnkRfuMrh+Qm
tT6rG2pZi70D/nwmZyeN12ee7CuPrVf0onblDrl0/3tQla1J8XBwKMC+mWxz1L0Pm3KDW7WONaUn
/LpHLFGJEhC1GGssKmMrIX4lSBy22Nhk+QieWIehvj0Z14jt5jOKGoUEGLLY6EAQc3amtilIyNar
RhJaxLrDd3WJfRaJ6udLU47Iemc8SGpPosXu8gR00pR3i4abtsSJFsaM07Xlr2QgKtTPhrpNv5fF
QjZCnkuIOR4RRMc8oXcRb4KNnnq0PPHysqaJ6i2Eh/7L5928DxFIQl0t0WCdIGiQVJx8/KXyNp7q
h64oE6e5SGfwgl27D5vTAum8//Xx/obcd5UZ+F4WWDQlAAh5NB8A6flNBIgLRb/ViUh4YRxkvUfM
9dVbRJRBw0PO6nciKNJAwfKzb9FGgjVBUoNJCW4lMcNMobjXQgIzzTJ/NFy+XTfU5jBsn0Wdebyl
ZduW0hEz4LYdgMbX0B5y4sVRDZD4/o07wfsT2Gqlh7F3eqEZNd1Nb0pNQepwLb8orGuUA+CLHeoS
4qBUmlpT1A7uEQS2yLfMzXZ2XClo40W00fWMlEvvdNtMwaYmBOTl0Jhidl6EKDTqQLbUkb8KK+dI
zY13QhixrfnGwXwSo/ewA3FtlmJ1IRrgRIl2wYYEx5ECIbM2yWsYxRljENhyJ5LY+1GOueCV+eA1
6BZEkfJmt5CZZ4wBeYfoLzyWiLvtxnekWOA9q/YNFbIeUidpi6D8jiShD8mjRYsPEHYJOOFhHrz2
kbGlPgJs0U8Ps7V3CYNQR/vRHbQUXg1uIlAeCI0McwpP2Uwc1NQFIlcasJUxhJj+pq0EAB4FvBjH
gEWGX9wTVKuKUx9OUy1AIPoMsvRbjerMGPxxGGUxBZ3TK0Z3OmQUEc4PaAoUDRj7LGDCWkp0S1y0
g3OrKPQUFfDA7mSYhgpih+7QQ29KMOKMHR5XtZ1Ms/U8sC2ygr51bNotiqCLp1WGwWDNnqsfgqnX
xCtshyjDp/D8zN3uvMz78runHMaY+p0xKmSu4mNVqYDHGoWZChVp9Eipd+o90Ib+XazDnJ64c9LM
WPH7ZGfwPvtpjSIyLCm/gxrveH/vjmNZfx8k58Q9jam4nNKGSdyV6Vp76OHsfKLurAXoI52Ksbj3
BKSxMggV5VjMHLe27OEF5pdbj91DLtatdZKp8+3QF7wRlW48tap6ZbIfFXE+XTyvV6FUPGFCuAXf
vhMlsrZeNNVop1HyxuMzXx+j15BH95WZHCs6jgH1dTcF4cFFn0mTw/mqTqyE7oHCRS+mJ8T2AOj4
ilo4DYa9z3AUx+nlwOm24oO5Clp6UAvWXuap1fRhJizLS5mAaAY3rtf3cRPHBDa137oA8weaL1oe
DvKJSckw44Ffpv+INRe0MhkLmfB67mv/f6CU6mMQlbctq636EN1C/o+Spfep7J6adCmvoC+kE+t0
C/v6znarGFnLT1ca7jY5TmdZsyw6oZbrS+E+a6LffJfidR6ecQsCjI3HiQ+iMNdRg+AeGAYwkqde
vSY7JbHSRwh8wjzsqQKLikAybY8+wbfJHNUkxBk6TFV0YyxkZS2NjbL5oUfJkTowuzi10vINNPH+
5Y6PAa4rE95c2QY6aokMdQ9cwtGy3M3Y2jgK/HTz41PU61XyQ/8beAjuMr9X88iHIDh45/BKti76
i9EpdtKPbn4UmNbSEKKrcdgMeTqvSrpiJzCdIw0clRKQicp7OqjTGXCiE8jKoSxjheKZYOIClf6T
Nga0rnzzbjmZsF3t4X3Xos6l+HaQHPMSzWBhpV/zKXdpPq2R4yiCfLnK3zu8Rc4T7VWlsK0+esb6
a7aVFmiiF91vlcGZ3d9Kd/l+6C8hHtI1XCepZoMmzdsE3k9yHqCUXDevvHXWEC8avloItw8QvFWK
tMv9JRAa6tLveZJuDwWTDEBtn/HdIBExl66aFGTlge19W1m++YduI0okYrzFQzz9pZQCw8C6BoSx
HtXiO5D4YBB+FVBY1HKPXV3NdGTEzoMX6ItzqUcJDltLdEOwqSnxzRJR+8ZN7z2Fe9wZMjnF6gym
ieA/82fEoYjY6URTl3gRmB335L055FhGinIOMc+l2ehnFHnhShFn1idUkqu1OhIiQCWTe1Hf5xbj
vLMpyqzhusPXGwHc57mEBDxXye/te2Trxxnaw0NFe6zdqhpOgtzIZo0yBjcyIfGnmBqI+NqSD/e/
WIJ600ztPAn627EIekA2xz1btHSeCZ6c3574lZIAQ22RhpBGqb0wQGp7jLXvIqMrp31nDO/crfNd
RqjXdksfIsXGIZC0DxCXFlJY6B+rvcgDxfjHQyKBMuIUCyDtR0gC1jFQldMJ32arT+tBCJI2uI6y
6JjkVralvm3MYzRj+l5qbovsMniWb7ZZCo8ZPEwLVuDTPUR3qCw2gozhVGSn3nQ7EvmQUDcntB/Q
h+fTIrlrq70QSOBSAcQpX3h/9sAB0PzEw2Ed+ASxyZ86TfXuhGc9oyDUMfAAlVRcmZOkqyiBAAbc
Z39NAKi0MzQYgzCcUaIi5IQRGFJzaPAuoAv4v/jmvg9RV5Pky+Fc6VxUI88sCu9ldpbRHvVzHhHk
tjvQiw5Zw0FlUiQb1sg50VW0VelBHqUyZDBSJriU0+yx4x4CE1dclX+dBz1GYscDEtFJluQB0eAU
9GL57tOeuL3ZUwFpUt7FEPqDSq4cd2zd+jVGINY+dtc559sgjDHcdk/tpAbi/h7REVUe5gH6cINA
hc5NbtZ8iG4KUB+MFOw6nwER1fA4k+PsUvnXUZQe95VNDqViabK7QDll82T9JPRVNL1WRwCG3hik
zfDxNxBkdcuKmHQ8s6lRgMktZQs/mywKx+A+yNfDEkWOeOf8kNcHMbXB/P8LQ15d9+eJRc5vDpNt
0eiZoYI8tYYjC2tQuS2mNm4BtD75CGQnFqYujKPYXWijRQJCPzF9uJLpk11GplgNHaYqDd2BvT55
eRH40GQxx7g3TpDlxy/yL5hmIr5xb35+r609HkpJzPCduqC1gJ5hXqa7PBQpsrrT3Wso2x8w20gQ
pXuPWAs+/x5b4BCVMpx9GAbKEzQUKIteryJRewbHn2OGRDIDQazZbhXthfHoJNR9KLIkMG99F/wt
LAjACLtABpbdlvsV9Xs2TwQpK4+ZtIk26wFYjb07f4oXQ75dTa3iZiJ4h+qgN4s6DhsXvDr+nXBt
anDo/aCaaoVAXju18JfUQqKQhW9zWS01k2Sa9ypfLmveCCDoDTBzrEtNh3Qgk0t6VQJwo7AEO6/Y
56TGe8KR9A3dNtxonHt/Uj8jHLHk6dWI7pSp1xbqb1rX1mMQz6HOi7n/o/Fbq9r1emr9KV72aEkE
kCZqU5AoGGpShK9S80fcOBjDsSCTnITpYdnC7I6GI6kwipXGKur1k4o1Gt/+UrjVMAsy8DQutVdF
HvGslbyYzID6y4ThsfmqVhXMJk/BhgVi/2v10oK5oxwzCI3aaAQRFilQ22+N7+xGS21WWKQ0XSRg
vrGQQma/TnJqAz4ByoQWCfhJFLfzVE1Dqik34ORthQYflFu6Z2ymrQWcuj8Ltf7iETPWQR8UiIXh
aaml7qKI7vOPKrf1mtgzQDVLJX2+Yf1n8ltZ//UXRmB7+t/wl/ae2MFAli4y1E+EmtMuGnp7nRt0
SzHuW3ULt79VgWeQWAAltllmSGtpyOCJtI2VuGyFgZ73d3RwxHhFG36qnRDrM0GoPD9rqp4NJxrG
ZtwMCn+9s6YJ2LbNXnEPWJpiL4rVGdSV4wXtlSaBhC/bd+0RU7CJXPyoQH7L0IsWXrqlU/W1pI+R
6f2mUUJ3K//P0Zzoy29KZXbAcrlsZDih0Lq4xAmYAbOlGwo8+8bOrX8YgX8lr4YplcePw6N/yfQT
Rp8dbyzJBHIqQgePeqTqBKNfZF6Dw3WcFihSiW7ZoJ1J2h5p6Hd6WJotLtbH7T4NmEMiP6xrqmhz
Lou6Jk84tMK/j2uyXz6BsxzFZjgZa/UXSYL0CqYmVUCPK7CJWq0rPQKZpVOCu1ujyu3MpM5zPJpr
Nu+pt+bRxcF6eaB26lZjSnYX9J9EOLpurN9Qf3Kcdkw9YmQCV344ntEGP3M2MAAGFH9HZq4qeTGG
rZ3NLmS6sSO5tPSnCr7uSn7aiMsJyVG09iO/RJnNpjdhBc0hvAxiLHbK3CwZ1NAb87o4OG4xzFSJ
1nKNG+HXv+6pEfS5shWqUYfgYSc5bTXF2oAQC8k3s0XMu10LxonCiO0ANXGqkuoQewX8R8lWn84Q
FRRgmtRuNcWDiUlg5n8BSBWjnw4oX3TKTYVojO8EHtoEhR4yTJTtR4060xl3fnkHcrSWoUUrLYum
YHq+LzEwcttmy8uP9HHPqby3iA1X5mgVMBPtH1WXmfXI7kl2uMIO01985+szd54ovapVp7JTfb3K
JOqCOnsRi8fTjKGnZDF4d3sGooVfIKiViap7srhXNqGnSLry9ttsRKL6u1L4Oy7Vz9k44B2kYtml
dTDyOpagYgIXxzUX/RmLihn32AXdvMnVQ8NFqdVh9mosE8EH+kDMmcNyuQuYwjFY3BjzEIM8mBPd
ff2CLmg10Y501w9tChUAF/rBTBkS5dFNcRSEdkhzr31gebi9wRhYeDJDcdtgXFNPimcPaaPGogXl
LqphDGDM9bdc9M/+Er0ZszVuG9CxntN4EXcv3MQ6Jp0YFjuXSjfYzLisIOh5dg0zoS7EXpx8qNvW
yg0+iEZGtiDSzmUH9TdjudAakj0V6m8Vsz0XMn0mJLZuTkENrtAkT3J6g7V0crHwSRb5uy/GRXij
Z4q3F+XZKrY5fM9EDunUn74rh34b+iQO55z+GmQh8caguVfeBPxnwZqXEFGPnVqT5mw/jPS12L3z
cofvH9cyGDSkWasP585dMrNIBYnhXQhA7z/LX27o+aUpJ21d/Rz07tab6eHwYBqdGWfNeAporkK/
7cORcIO1lTXnoKzpV8dbPU0/QlpvsPWQVNVjcrghY8m6E9OHGtkASX/zw4T5AQSEHy8blUfAAR2x
/2HlGV644VqwJfpjwVp6zgY3+Ep+FD65SPt3vq+k3thFXCNcdDzYhJFu5YO/4Ky9hCTuTNOVqaAm
SF3p0ecZbAfuVJF71AhZEvx0kvPt9CluBemmErAGcMmb2nZzQ/uXTHLYsNlTsrIkNYKRM81/gUwB
VMVfezeGAl2e/r+jIZtVZbr6DD15pvRbQnsNKWEwbpzq9L/u3LZqIb2nWyxd3Z6jQEE1OCXH8GaN
QMUctqQ66QVLBrHPpxHK8TAuvUSurpZazXpXa3RYv+5k2H/py3uHSgRIDob4XOOTJIpNxYWYAXK4
pq07Kg5zYeLcduqdDpDqqg/fDui+FWdzzDXlHYJ3rKZ5L9VI72RdYMICtkG5Fj1zW1mErAf4XIzJ
19HeAmzLD+Frty8rHIKdXrBpUq88SmvprXKNyse75VF9erWWCLxf/r1xcjDgcCMgKfA59xgX50aT
LTXLrkt4SX33I5xrEM7ne1O34qaessMILKPObIJ0v4DZU0Sa7WEembDg+8mKv28FacvLyzcUNb0V
bQOVJEwj/iMAu7GUFtrgtSrJKo4MYLqoodUoKoKV7y8OfMMR1DVVaDlzquS8rQ59o6eFRHOz4PVX
qeQ3saoWknsfq+JrpkOgwEM7OPI772vHDMLw00mbJib+WCZtmaRETNcWLzQXNgWnkoUdQKqoS9o0
xO57oIqTJgHFiodewsvjBMd0BQaV5s3arfA6wStulw/m/jOiJd3ndH8UU6IUk9Ldkoa9x8EjkBVY
miFxXzjRTh6ZYUvh+50FLYpNSZhzdOkqhQRK6LZGuCitEjKoWDSq7EIoceKS90omkPaDvPa+w1v4
iVaxWnQUq7hfCPL9JHwVGvZGoycmTkHwfsHKrtx3wRcD1zpmlhPdJT0zBr1cFWqSkjBZUeN9Gam+
gVUm+CJTUpuyP4VVvNI74dS4Yi8IkZ9JlMETeRaNFVsmhjuIvEw0yxPnjiOriAdwwH359E8yDLRS
1JW7Vr/tUfHPqsfObQS1YaReO993o3PF99y9nPg0PBMYRLur1zID/wWKXHpNDj7codgrPXamSSlI
jqh7QMr500e6Ip6bIsXI1E7t3Ssq3uur1zm8LWB/Ubi85Nnspz+76ZYes8FbHIUHQEPfTchAnRDt
NDG/67g5+V1RxFdoF3E92pxGEqcp7EmeiNOY+5+sGuhfZAogcUgSfBEBIxHTRMwT7kvYsqul75dY
d5+yKZbqIhkKkZS/W8lNxoKy0093CzN2bDFX/Fo9fs9bPL9sOmn06FyqI1zPwM3uUWKQ0Ne4Bu/n
DQ9LL5S7bj2eIR5i5f9VymS7QYVk+yQ8OjYlfRgaMCHcVf99VPlgHwYyrC7A7hcNnS8fMcAzm58d
+Hd9+tSa4UefDJW6U46p02+N/fA8pPNarNj8KCDZCKH+USXbbMCiUjbnX/mIKbOzyz9BYgks8Cby
4kUXVieMClvCqC8AAzTvMbDp7Mfk32EYsmD8Lh72aby+7DB5IODz0836kd+jFmmLwbXQXASIgLcp
ni6+iP+SgyD1gh7jSILdSPlX6Q5VAiGzfXBqIFNADkSLp3yntB0B3vlGxVpAjD4/6hP0RB6elXkn
Z5VYoCW58W7FK166ov3/HVlW+kcSgy5VEpIFu6FbDrk9Ja+i4qhB4eQqnrKQ0T4xqTRa+S59epfM
tVLkdPlR84ovXFWVqq67dmB3EMclYOisQViswnTPvT/dWxM9py7eyrv/0aW+XgiPMdv2pRPnI30i
ijpVlbKY88ro6PKmZbFNPPxsvFFJan3Qu/m2FdfW2Ox14xIhQdYjYwpttG90GmQg289F05yVdPZG
ti6TAJAhygqzn8zadZ3UM/uyPGJFV5WK5BV3wuIiLc1ULofqktZzmU2K8wqYzXs0ed+XfYKMNyXa
GIRal4+GHyYTl7BceUSCpj6TTr4ip1vq0Z865PRSGaEZ1FnbZgEgwHox0MKgb6U52/Jaal/1Ad7C
7XaafUhU4YepiHPIODDGdTwUJEJzjrZF8P+tnPeHQIqnk8xtsUb++1/ZsO+6xLWpfCMuMudPM0MQ
nZiTzLkSfrjtgav0kRHRqFaSjFA09vKucjBZmU1VzFSv7UHzsy+/vE6OPL5mn3m1Ley3p34JwGcf
s9fyoUZ/72OGncnXiPlDDrY6xXzBOPiDMISIu76MwO5jpVbl7dnkQeqk2z8PZPr/imlecrHviGOt
gTMPv5fjJwp0wfxxb/HAC2TTa/HDb4EuvMSP1AdauJW4qnC3OkGn8rSf+tMK/Kuu75oXqr1hSGI1
iwwaQadIzxQvuyvKhRjIuhR+7oL9e5Nw2bimXe8Yr0P9Qy3mL/QeQu100J7lZF/sHP+hmxjbp2NZ
6BBGwzvUbo0+RSjfCH3wfpnWJv79DV7KRI5E1ZsXAP33d4BI3puZfDe3PG3n3d/USw9Qz6/mBhKX
PidWh2eI/KQ/6KYqa9WmkdJ4Sx+NyOGlw7zeGfG6hHDnJmwybLBgEXtqF27SulemjEbA0GOVwX7j
ZRYjqtAInqDQBpY7nqvwrA4sasGr9fE3t8C+iVnlBezyvv5irK72XeZhOB4svtNOX4I/nEqr+dox
nG0IQrnZtjYGQuPYjbAb2d/ClAJ6uHBu0tY9PtxOlDZg8G+piCWgLDa44S7s/fGWdtZv7PnWaa+C
CP8NlPFmj8OlH92zfoLPj9v3iKdRXxlSkQiTtkVxRXe0A2BXNejz5v0jPNgkCQ35htjEoi3vnjq0
LgQhZXcuofBP1ZhWfmjTVEJKWJPJnTbk2QaptW07JHh7OdEler47w7aPb+G+V2tEgKMDUaatecIy
2Zj0aHv0py1S3nMuMS+Ct8M/Hyh5EK/ne5naUz8LGnlvjJSFitkd5M0mp1Lc23BFiYWar/NrZlpf
UhaQBbrTSj8YCpleqXd2174VsKWxHAFHcQm/J0YhJgOMn3Gjt2J6eK8kypWgQadME6WMG0vIJSLS
MowuEcw73O67HZVGthe7AcNUq5ty5Myna0aURf/k3iCnCE5Eb/rzUPpoHpSa3cfREBHXkb+3Rtl+
LHNok4P7NAvvNe6rnboRIj94QEuyBL90rxBUmLyfuuygmsy9PNJpYUKQw18j7AlK4y+tc2FTrDbW
Wrsf4GjsfysNa3ZYTF4l3vqWHn0Z7wc7BVL8A8ZMlA2tmkmWjbi708YqL6sHxpZy1EREt8E/E/vw
a/NtGs/+to6HSALJloSo53EVnKbAJmsJQhW+Wg3H/vwNBwcCKA+8KbijevVsX9Kq8ebbRVhVPH2n
wXS0PoDcULeb27aU4BBpTcXYPLc5MdKpGc6MGFSZ2ObuTFaIQW4nKtBzxnpo5tzKoL5oiR2vNeWB
CJ0r72p18F+cA9hpTzD4j+sAWYyABAES2aayP8QhsE1refKQq8lb/KvvJ36w8NqUNWMl8GWw4TOf
z5dNT0FYCFnNZ3NEOmPMZj6NhhMR9qkEV+F6fe7/z1WbadTdWweOKcA/tMHLOhf7pSH+lfAe8OFn
6PsNo28C9HaasaC0+GWbJ6fIipkrC5/8F9Eu9GZjVuf/F29YREU85eYNinK4kRk+66nAjcJWvPSG
r9xGXdQAo7vB7zAxmnJkJhx7Vot72DBTNbOIGXglDZ0AGG340D1F24ukrk4RKXqhMw0MKbX5pkX8
QAF81dMSJnZloqabdE/qKcmIWkY1/gsmz2rn5X/wkjPf2IVxc2gpY6LYfYX81mm07nC/vtXqgxK+
3IbMcZ6OxqzWFcJzSRfhNTm6fQujpj9ZUhZwOv+Fyo8jTtfy9TKxqFL+PmMDqwaallxRG1oGgP2P
zqdeHxJnH+nnLlUHo6YahNlVoi8uyLP9msXc6tft/kahznyF8qMcopSXxGNyj+D/2kHKVUsVPRMf
Ss+QwZRjB68R7gaOp+U7kKKkj5qf5JbMh2xpH7JHCm8JpuSixko2b4QpAUVUCdqOUHJHDOTEjCKS
6ht3ZzOAt4tCR1DM+wO0ZdzuMqTXNaW5g73mJKJZYL53PH3dcLQYm4XpTzPFDlwM2waw5/7V9Lw4
nOKeR9fpucNIZiH0njNyHqoGdHuTMGd4MvtNNIC83n5F83mV8GmeGJz6gOvaoJQJOWMR60mzZrOz
cn0eG7qe4Dffh3nIUnEwM1b0Zxb+BZS2YCaRLnizVmfDyfB4ht6L+eZdXlKWtJYbnHvrflAHR2qn
ifvVWU1CftrR70FPeE5qUw0nq3ydCv9zWGec2G0kqF/swK7bKXZqb4oUy5FwobQT3yjguNFHPDIG
TM3b8dP4ueHfVPqvG7PvRB5wstH37CKiKmwgAmXca3pTUo5S3wNXTdSb7QsdlWol+L41WGImtYiq
t/bZ47iDiHxiV1c3OsMPnMFNySWR0ZVBijBdnAosyH88Zkr0uyO1/e/CacQeuCXeFQlY0yG09in/
/XZ4QeFiljdQ8fYRKOq7ry6rC/uMSSs76VnlXvBfxs3gfQ4caPR2k95bdL3IZnBVlEOiBnMHzcse
3pdW5OG+kMCDTD8Z9CD0BsLhDzfbTlaL1RoM3JnWgZGK4qG5Bo3vvx++yqvReomHQk6FUmZuy35J
ih1+eRF4LF3/PK6rRa9OysL/4xpCGVdF+WzBN8ouijerLoO6LV16FoKE2TLbvveEByzQ6E00EY0Y
ix0msI1AbPbjuum+JaGsoxPBevQcGO49uE3Pxw3jxHRVnqBlAiSyKX03q+cP+0UCy0ykx2cRUQD5
H64tT5J3vP1OisVdZ5PzIrX45y4IUc5X3OG3Y0TVJg+RbVGJCPPBlOaM++XQIZEyqkZPSbjG0Nct
/s5fnfhMnbihE9m45tiSDyE1flXNQ22ST3Vuucfkog3T574J+rjN6cxvT5kimjvKlKxqXSdGR3q8
f5Y2j4RzhPmEB20GKJH48Gxu698skkVbt1ARx+M8SFOxmwbzFgR/QdtZ8q9GVazUkMM9cBqF8G8F
k+ccszYS8/v+veb/oKFMXTnVG2YhpH5+5Y9KMVBpSp/ylPjUHYCBWWzxu+f6HUeLYXhiATcYomiI
kCVPaAvsnlJ9dk5vlQMka0Chu7nA6ZYI+XmAnW7w8TsxXJLutFWivAWgfcekYsLx4ZQRhF2yopJa
O1Om5gp9Yo6nZBUu1xcuSIQsxtkZT5f4lhHUXoVxA7jJR93jZvOMrf/U4GSsAbD7Dmv98lV9u0yY
f8uKJJ8Q8dhMlJnd+8wyAMf1dt+53KQKEmuokZAPHWjUh3riPJzwL0zAwIyQdB9vltv94lDmhNgM
rHcEtf+wEapZY5jibBkm7eXD3/jJeoOFWc0JGqUnOz8KY6BVQk53H9xeF7EIDxvOsqAbikF3ajxJ
4tFCQuOvM2m0st5k8kN73VaA+DQg2surLLaln/Nl3OSBZ476qGAdSXEVngdIpqNY03a0KkDgqDzz
YZ6OHsNjciANoXndyouVKndfrJv1g2OGfPlnb+IUEpZ23Pjsym2WtIXzxe/xaykRV7IY8MwwmrX+
vI63+5Ioquac4Ac/j5zZTbv8XZ6nXwSrEMQj3n4OU1d3Mgr0eqENux3M4E3AX1fKGGjMpL9JjFy2
Hjb9eWJUD0TDfYWC5SRbEgmG5SySPaCCEbMqhjNmSVKLrte2c/ZwrSpEy2RnznFfgCLm+mdH2KqK
KlG8XMLtnooHkJCE3Q/KGoF+Uyjsr8gACFCWvlhFHCgL6kOi5GoAshoFQZNo6AbubJgQfudyySWt
vJ0iN672a/1FWGn9Awf+1e/ygTJfWZrwO/DiXz7wTEii7Q6bXIyj9buY3ms0LtX7WiIRwtOa6ON+
vksSoSGakWuccEoWWBiwJ+V9KHcr3vKD/f8r5Is6wn43/v+GYPSr4V1piLGz/pMvatc9CdA0pozB
VuCtEaZ6Rek/y2H//mb6Kj2jwarx5LSnYBxwamdRpSTT2L8s4uHMdin+iwT0qkb7Xs/4QhEv3orS
2om1x766vpFJnz8daep3fjxl826MdzAJF/dQkN9HJlsniuYO+KdASEXpBNulDW4cVao69+rFHCg/
5zISiGNZjeLvmZtWn4nTn8SeGmt3BO6PZs4F1lJwKCzNvRYsYelaVL2gSNCzPWUSK4HYMxh8wkou
+qEJQZtd0VUN2aRwvjNAgDbn1VWAJ/N6ZtHyS2FcnRNu2GlGPWNhfY/jZdaPfBYWXgTICg0AEIRb
6j2ELonFjURnAGeaL9ONFVB8wm6V8fXHnpzPM/1+CNgupg9YXLh5VjRTgJg5/mL0be4n9r81gKIz
KLXzF+DGYzp3grPnxgfjcEIJjw5zto6LrTdaTq7zFvnCpGbztDxridRpbQQcjjGqopYUkU9T0lD5
FuG+U6lJbUaI+yF8rcaG0RG8i2bSA2sGS7ybeNpMnCz5cJOALGyoOzM5PuCas4DIROR9eC+WzsSw
4zlpoRv9nW4oQLw5gvZINVxvkmwa/BPQtvs37DO96XP21zR4tUVPdBv5FjolxDG2GOQyoNwN3MIk
iGJ0t0jGhkFSFZuktHwyANvTAfoeeMBz3m1IOC+nak9yZGw68R151iZewVFjmKX7iUPpUSuaxFxL
LQhQceFoUNjAs1cjWFq33LX9tPAxnWvXi2O+NY8aBpsSVgWoUNqrvPSCqG1IalcSpjGUNmlAO/5/
KxkJMYjgLrJC0Yn1Thu1uC5jUdkMS6SK1V0pxqZ/25Sg0p4COxhRc1vBaGJLjG4uZ7UYs+p+VlXc
h9v1BZwUS/k5nIOwF8JDU5S/ltL2ahDZxLavzJfEvapUTWdjo4AIoxT0nBWEjwz1Z7cBbIjD8IdA
TwWs2J73pNOuRboHjXqLNzABO82mF++F658vVt606yX5HLqyC5USfPA3dpPG0kKW5VBTjbPLmWHk
YEBfsHQC0++7NjSFw8n5gMNVzzM+6p84HV0eg0AivWZk5yq3+QOPkbVDC6ldAoo9hwtYHoZZ4qvD
tjC5QjSDoVvYL8V7pLF1fdXS9e7ptssUDZObwlevOM6IwjZsInbChNMx8gi6XVFKPS+PDhzXvP6t
ZSH0yzcacrzNh+CPUF845B+7ShViw9auwK8I4xC9NEGBMxWxpmDz2qa7tn2eclObS6OgumNh1vCW
xFPgq5Xww5Sio1E5uVh0t0eVt1sg0y15kBWDb3vNyLInYB5id68baO3wGwLW+qy9EBlyCnl949qy
jgqumeh3Ac9keyPKxodwGZhCwvXSqsDj7Sg2y8KM34ZDVarYKwCxhTrJLqnSgbi9spAQNezeppyX
tYL8sT1cwvjcK4DFpY0aqBdHB6SBMR6US3tyL7d2x6578N15Qwzu48qoAmwqfm8wMKqAJ1Nq5zIf
/k/822mtaSPqW5JFwojseunlXjvY/Tpy6PpXKSVzWGSFm3Gsz6Kzx1KQ5ARoVd2aIl8UB7dvwndd
gvEN3pY5Uw/TEqEoTKQVP3tfxCNoUybkPziO2oqfOuftIhO5QuWcqOTnMBlZ3PQGw/zM68JArrHU
mxbyqnt3mnB4YB6LqHDKl9u0vPiDziM8Xo7294mg7JujCbUc4qRegXK0jCa44aoD935tCef4AKz6
/9ohioPFiuzV751+gK7zufaojcMU6Q9vAF1oPSZFQ41DnlZQPfvpgnCk1EyaKY0r4zPIMrejdnag
jAdREU0ZJUM4US1uYyqmuxCABqRIX+HiIzW1TVd9jSiG+1KO/LlcQ+GIzihbhM5YV0kFu+bEgIqK
qU0dvHV2nvKdtSKmFRcohp6QNwjmrG/4MsTTaozGypUaVL21cLYDhEda9JFscocMWp3NMIaZNHvA
1nSc52JTEZBU4H+tRBOnpInPLgNJbzfGFwl+b85x7xzGw/Xk8rdY/F6gmpzZHcC5nzYtbGFzcxoe
0FaBzmN7SvnKLQX2LKB9/jX58yiuWf286vS5WiCjX1vfvych0kPyswS91/ZEL5h+KxwalKFVSFFv
k2VgCr2Hse/W7btFmuQ9uO67iIyi/frXX3B8QtQveOj6ffWu4I+5KOJwAC+gZhKHEOcACVeArupq
+fjqUjMOMzJqRbWbNOh7piS607E7AFKdx/xW986LFegrgWNAltIpTFYOdWIRe32OhVG51u8mSHfL
jG1k28cgmpI+tRm1U9UfMUI9mWtI+5YtZ71ETFlzwu3bA5NHJJaub7ZOU6nrm42Flh5jp8oIw8LQ
brB9NqUY7DSgkxhALroQZQM7NJwjacmtbI9skBCGuDmUV1HWKTc/W02y1dhlXuPHFRsUbeURr8oX
AH1zcAFpATRNmKhTN0TCC/iC0ipEiqqjQCqdPtd5vL9HrnGtbQxfkokzV4B0dZiZZkLahMlDiDZ9
oWsTu6hzcJED9pBKb3BNNDRsCi+MVfR7lZeFl7gIWXkYVxXGAT7uzOmLg6bcPi5yh1e83xtGZpMx
YtrLVY84aYcopCHJtzcOp+nm+gZFXdw347L3chzAnjplmdz/cBnzkAmplaQCcUB1utFOzSkyN5iX
PMFg14PiT6FalhGijmR7aF4xbvHeVR9m6KWPQBBVTLvNsQ7L+Z2bWX0ZIl1QfwCaaEnQBmiwUgUH
VBcrgOla0T5oG29YaFouN8en+duA5vdBSRJmFL6quXxknZf+x56pxyuQY6AFYGxwfxx6m8/Taeou
YpHJtYqnAeCKdZ3J/gvxQmisp1iN4kxmzB5uHDBnzzH39BbtY9LIxhR7mqMOpcPV2+kO8k3NCbSu
1uZkMwajD2n+p+8BeICrunvvqfeY53NNP4+V4Cep9rfUITr+8AH65lfWvkXuytf2Twz8Xht/KbZb
3yztmmocUJKNv0blAQDMpruMGQOdA9GretYk+Ale0eikbgPM6tEcp1LDJbbPqp+ZW7dVNEuP/jO2
Ew4dtw5T7OvW/1aErUn3Ro594p0L0bZ5f5X++r7GiHJykGsV/TpCOtYLZrUtAb7Dtr20vPYi/hIP
sJUWHSpPdzcKxdD79ye0GSw0J6lrEvfAbLkQ44y8tOTojt4ZgPgGpaFe7jhW5aCZ/3dr/ey1L+VL
X9SCg5Q2gOwVuq3RN7SJH2IP7b5HD0Zqq9NafMWFJayfZxW6+Z5lOg1NFpAc9A1Z5NQN5gtr9sBV
TkubsbfAeK3CixQVM21ElP52Z0AOg6DhTdIGi5+5cexKIgFWxgkAEzv4xhaUyFxgmYRbYQ+Tvvpu
496Klw71KGSIFPCqs2jq5910YkWKh+qzvZKVYOQv1VDfpSt2PnIIa1U6md0KD7IOKXKxsQIUMphn
aMpfYitbf0vApEQMrWBTgfIY+IEZrQR615fpEPuIPWM4doSa8OEwZkgIFwJj/GBE5w/9cgZT8Cjx
8N9GMhAJlSKBnYpC2igw92D12g2YiSHwm6//CYriWUfQgsMLjJBJaUh5LxSN+TrG/kYyBZodGb9n
Bc3Cl8O65CECCp6PqKOtBsNxgxLEhRpjrvca1UEHjkFrLT1cju7jJs5tspxdimQNRtEaKwDmtM0+
83O6qKxux9mer+6oQkFGT3WS4r/T/TdS/0sywdvQM/idbtyama57fjTLW43m7WYM43KkJ0/NlOh5
+86U1Fwfhr1q5JCM2nMqKQcOI/CIGBfKcLfOcTP46Klv84pliCyfuj094bCkXnQJkwAAaOOvOqzT
b3TmIVu4ivFPe+YXzmxeGiaMDQ6juALxOJnpAZ9Sxv7HOgzta7EjMPuqdFWiuqHCt7DE5IrdNTtM
+UgAhy4ejaZqFBwIH2hvLu7PwAsFuUQMWiipb8srR6r9ZZF9LGp/EoJho4J9kue3vinrTFSiD4mb
wOrDT9kuO0GzjVhZu43FfqNaziwn8Ap8vHlZf35rP9ky9NIHLSr/5XXblWNGUTSrPVDdzT8oGJoO
G9jrhHZRa2WQpPxR7BhquprSyjY5/18hmkkiHP9td71itINaAP9LJM0qv46HF4vCRobh8pkQ2oVm
rSs1Zm40ZizQhd25keyYuMNMjVQhWs3t3Y4/JoBEfx9VDcnHgGaOWKVuo2kEWIh68j86B7NUX6sf
Q21hw7YFCersm2JSLN3Jxviq2bU4Di00mHao0ZcaPok00XFu5Q1gQHXADc4BUgWMAIQ1+/iqncF4
yjKmblQbeodoEBQ/An3LepW8r+0DpATTacIIErVpNYsXOKXupCVrMIhpfWQMeybsRcvi89275qT7
Jcpq1+gmN5g+oUF4Xob4K7ZWFRr90966vpPP5DY7dwvn30BbrMNndQlqvEWLEWnKoIUxuNsapwky
j7KPnUbC3vHGOPpOASoA3rVhW395wHaW8NK7RO2gltn2Wz9IqcBSzQVOShW9UU8QH/BKVfFJKluB
cwb7BWr6bCWacYtxdgwA8KSfY4bMZY0Gl0yMrEP77SOX+LYkTlZTLKTZJ0KKkQynCx37w+pphytl
jZ/4fNYejcx35+qLUOjOtWm6gLefsUH+54hKb1JjuDs2o68gvf8puuI1Gw5HwJcB3BVDh5mZbt3Q
NT4xBKfcFV8jX6sHw5PW4CnLXBNoWyYBdzLHWp4eGDUbLWaJdJvWjzWBAKKai3iT+og80yqcnmsg
kW4+ZKwURH50GHUa3GOaRkaj3xFwo0LxpJt/qt+RvNUPHyvct4Qs2sufEfnAJRTge/CcUiuVDhuO
BmHWmVtJRlqM2uiHXkSmjvET37EkKgFl1RhVRCvfGjocWavkKtqaPEmaNqG+edLPU4VPeTLpBhzj
/GrfboWcCXPi0tfxdbr4sVXZgiVP845dYShj8kdBX25yp9RnlndO++8Vw+dWj/KA0TQb7amwOAMS
ZoLWWNy5Ay22nP+AdBeyVZJkw1R1DzQU3gnxofycrU2msNQ3sheXzi1oNNRTS49au+T2fDTiZlWn
0UDchfpZrukPh1sl2l3z6xMh3ymwzPfitk60s5nzcYeZEIJls7h4L6qknVqle+rLn+2VoqId5+Bh
o/zijYtj2d+rAzvI/LR7/2BxUHLK1/gDapQoOhhTlhUXkGZyru+TxWrA+WWwgP9Z286+qaDdFbpB
MHknZyrgn7oJ4ON5Zmkt/WCqPYFEggMysxcEZo6aONdA2exs8f2fYS9pDzRcO0D2C4Z5JBtzcO2L
Nai/Ks8oKi29/Y8IzQw8bS99D0Yo4X4RuJYLRGevnTwjNxTu7ciCoe9+V4CDXSquFBJknhCBAexy
fA1GrXAy/ETk8lE0NKejfjHRYpmm8/ZDzTNTrSet5yxviGNQ2qpbIZAw9HdPSgV+37C51lh8cR2u
ErBzCuhO8iFVKdc7o2q1soKosRWBzerW9+REaJTT3vV9FAf6b/VGi9/ZdcG+Rqq4a2Xl5THVw31h
TgjJbp+A4Sz2GQsyr0gCZJftpN9iTHNneWLNngClvUjvjIs5RTn7TBxOsrLXHV3jRJKNFFUni9uw
Na8eNaJPprD2+KIyZX53ea2rT+QONZAPi+G4GBQaV7YQ/Y0TWa3iqBIBUshLgRT2W6RUvewH2ZyG
wivbgBoW16fRH0uKECD8/etANQOiLl4z03ibrPHU6A9kaOGlfvmIOG6+whbH/vVNH7YZ0yIJSui/
wVJgSacIwL1tUItBaH2HDhuk1Y8FUHCjnxTlcs3vqovQPq+Ldr4Wk7hvD8AQTwz7Dco09TIlH0Bs
IKMahWcLEqHOtokT26rjNonwpvlErfAf6O8aRBlYuHQQUm0XW5fWKHhZ/OigjOUatDmYkslDPkQJ
+PwLvi6IkJYOvgjFp+a1X8/v35o+CWkaRpuyhcfg/hsVE+L6+7EgDketNX0rTSsc9O0tA3+yY5Ln
11gi9tk03SnMgA5VeGbTzWLtBocdFMCiGy7PtaX4HMUv8/wdq2CsHdXX/GaMZNSjHJbelhggmgSW
OyuaV+/it923wuNyM1Km1jlB++Vlw399cmK69QL2ycTaAj3bJAPhFKvC4G0L4EqDdquoXKZ90Hbb
j8r4wLi6JbeMKpaoE08kJAcBO5Sfsn3sQPYPulTqrCTcLQVsd77U8AgHn0dGOat7xKBbHLNUfVcL
fUVxMKJRI+QpimtZZZkTgCnj+7VogEvwvDn2dqnJ30h9Xxvbh3iH0avDqF9REwPKqimhWh7zogrZ
jptElfeKAC0YzSeW8xrIFh0d2I8PU/UlPbjrukqUfkTWQ5UdpSI9hO/2GHxEE+x+Bdg2Ukla+wIL
ZUAKUwrwAaIRQ+AHeZi884In4r1jFqUoDL7OL9J5HpCZcFoX4GJIMagqiD75iz4tlCiKFOR1k2We
bO59eLCTH7y6/Uqeh5Sr+9wZLqfJ3uz+PGllrcFzvKIBot94FkwOb/CuzSc6L72WAF3JnPSUbBvJ
3YKsMLJh/CHDpIJHSiFBIr7z4qAgg5E7bFwgtObCs8OxoJmSZCw3IN2Y3xQEIDbrM1EAkZ+jaCcy
NmWHF3EV2QPFdVBCmC84lVwKdJMTx55mjqCOkxwUMaHyM884kZGI5vObXYUpoVxNp1SaeaG8KGfy
Tet1rmiuxOkotBrjHF1zCvQjiYdsRZmm+9QPvgjcv6vLNnPj00mp8kGoVFtDnO5LtzwSOVhq2/US
coNCKO9SQfSOpG1bAUapQTVbE4bw0xNZVrmCwdQBAMxLkXs5h3sOKtTRih+eD8Ue4lRbN61mkHtv
ja+ZEPScXjGKlQ4GGgE3s7m2Z+URPsebSJw1fiRrimVxSFOj7yQVUJ3Y6jY6NQcb1qGy2phvhViP
lW8M18x0NqADrezPBgF6cKZVflPI2mMvVdDadBBGMLz0jlKJNCzsh3ZUS/FeUVpLhqsJCUr/rUaF
uu/Zi/OVa9m8T1vMUNtI9YL4cy1BrV2VFm11hl+lmjaVJzJN85d+tum/8fI5YuImpgH4KeSdCBKk
AP07dqqOe1nzhtwTen7uujqpJY7BTJNEahRMwf20fJ/X1tmLRy2qecHCoXc4dXzetaXb3rgCix8h
aMOi96K9NEfaLfWiYyGhV/mTQS87CILhiOie+Q1oWIJ/MO6uF31LkpjDL5A0he7lu1R0TuJB6CnK
VqSyQ9HUdGq1yfnZ/tBUx/Ao239qpIkNYC7QSfJPpw6r26ang9x9edvXI/2AaX/SM304CYK8BtpI
p2dYti4BHITLZgCT8Wg2uEykmjR82S6Ae6IS452Bht+d4VJt1ve9Ep30x/HAbpd0SfS0gd0kLbnQ
5S84UBq65OkARPEjLSCakZQ/2/0pRQBciqJihHwvsnx/jZdpulxcxobJ5mOYggYsclxOgyzpXCy1
hQFAg5UXYNryeLmpf/wQ/2CiYyNClN3t6OSzCqyRrNSwweyxLKijYg0BBVJlUN/46srSlNBlvJfW
pdhw7MW7VLJg8G5gG9DqKg9EFPL0S9v9WAeDhUVefzrlqfYjTHMg6pAExtk7Vz34ERf2fnXUpJEw
ZG/NrVC1ufJGPUNkzPGqpfTekpXpFsGLyNId+JRbSouMqoF2scNe9HcLosUr3lP5JJ71X8jXgSx9
KM/a3WrJ2IXUEZsbzApm7nvYPzSu4waV18BllQGknAHbcqaox73od37bj/tjIzM9X/QjoKjhN6ZI
I42rWcZjrBADl+mbcPSBikOXnahSxIoPv2ZhQfNAcPJ0910iYuuuSAIHf/YVq1shpXGYeNh8RgYQ
gySqhe5CVQ2ZU5DrGIshxmqkwi7AY78TmNOZL1qpKinASlvsk/gnSUiUNU8N631Jsb+qzYopH8rC
S2O4HQDsBoNbqwQKvNEQGoQv6gM3yFs03AYecngmbDUKXv1Sbq/DVmy5PJ5ftHOX+fNIlZinPjh/
ZF3ne7vxbNozkJ2VmMKKixuMjsMICNDB6gY/ZZXvNjdr9sx9Tgg8Y44u4mMogk4NRzhFXx7qjCL8
6ft0MlJoTPlrkO5HFlZsu1PoM76wbhvEGsq/FU5yB3fEi7xFmzQxYOLhpDnrilDMphGZxwjxZPrz
re+mXVyjnDsU3nsNPXtRv+mQ3oMv9eX//rAOfiuZ2PEXiSIDf/iwTTwpmjreuGEmzKxL8uukU+Dm
QLBvOTR/Cb4dV7QzoizovvdPBgbRENfzLH4YFHhPvMwrvrdUXZy73tXmOp+ws1r8kgc+5oIVXshY
xDoz5HA7uw5MaMZqcO/tigzOr0lYBEJCaDSfxIClMyAfBmD4x7KoPy7jYEwtVcoEIPP2SYSPtCrV
45fX4NTlV3uFMWQCUSzs86Sr8rcjlNw222VqB5Y9EFAI6aaukhIUBCDZwYRyH7fUnw2W8OI+BZ9d
W3oD3nlO3TWvsFJKnQLaUgx8wjYSyeEdlH3G09VVh+SYtQEWfGbV5Op2NtPA2cA7SE87wvl9kB7r
QX6Q5UMCOeFKAnqrmWRUWWvKNNPRavm7IO3jMCxzLowtp30utAiF4FKUqg0aBSDlI3LwgfHwZlTy
JgFUGi3LP4yfqK6zYhCQ8MJk6ZsgA1nD40WsTejze/6PGE7orJ15l/Gn07CS0cFMshAPFKI0Ennt
gL7d97AsPALjCgWQhyFHTxnyTLTMzqjLVJXKwPn1kjs7uexVoOxwboNAIR5D6bZc8nGtqSY1wgGc
ZwKv5UwSvNliyFir/eeWTc4ANarN8Un6lahFk70GF8g9qMwYfyVSFgPDYOW+PkgIqEOLWq0T3R9w
n5+fEDxuXZB2ajfUq0V3/zZSBvtBjy1svhGQB3enboqUMzwIQ0gu6hMjz+YjwRNlbbfpMfwa7aV+
tr3vHRehVuJrkpDLvUQCRcNMg25GvX2mTrWDQ8U6z2kNgwvo5hQN1xyWHD5nVQbNS3OSMWq2SqV0
SUN7d1T80ogbIKRsY3bfuCzze3XCfeFcUQMorpzuCQExo9VDer7LDAbI3e8+0/e087W9RN9DD1Rk
TIogahv7AMof0FsuwHkZ1XSmZPEqNHdakyWroxF12Vf4ioWi7HN84E+M3M9GRQDGMYgIvmyVBvhj
6uZi7B9EK9RpWAOYvNYBOiePc+4OKfit9SWQs88ekWezdHOLPCBoexRdc2X0XPpug0p9c2XmGMFV
6YSKG/nh/JNJGzLTs4DkrhRwISbM9FPDWfbtTO+UrKQHxxHryd1qlMj2Cx8OULJUmo3/mb8b08mJ
LgCNjOlK3h63uBw6fv5vWDjIUlA0qjWiDyVYBjqU1D67M7I2rescweUKkHbPKaVeMhOwEqA7VY7l
jjNxT2GI3kJ/S+lVduqoo6UJmwB7xGkhVciSVHtIXY4T4DesGE6DlTTusd90O3JYShEhWb8pAtqA
Jlj8Qslsd/gT+me4kDWCOTvaoVA49oNaHA83NwpAoTI8aNv6mV/rygaH4Ahhb0+BsbdG1b4azY4H
82zCPjl/2u5KO78qzV9zmHpausBFSK9tFhfhfU1itq0fCwt41xA9b7gwz+RByN1mKSMBvFO0l09K
F5kEGhUk+uFEFDvxD44h2/QGA1XLp/gKMul76a9OZJCOmZTiIFEe2ajlNIIKCVP1pJHS+nBYaIDF
TFviOHqrQk0hW1HSZT1GPcGDtK5xD0O5wiA94GacQsSrDKx4+vSwBCfM1RPDKSh05JaMWREKJXzP
w/1qtawKJ44K4EMv9C0Ecbq76rXjTJFF0SEMRSmtBK5fyCMYYtJAe/3fZbumVBTAfSywzUZh7sp7
GOcweThcJCHaa99oc9VtbfG3QyiaqqBphBL2eImJ0yn15nZrHhESKewHlueichvOCIMPnvx2nrM0
GwmUlG5/HZwWMPjM9qnK06fiSnONkHMcYPA+kw3DORa0t1aCVCS11LCKvGfGhNauNoNtU+LLTknL
Kh4nGsuHtKKhPFncFNkWX92cIuMEro1K/z11dEMoyYTG86niruXECl7Uqf++DkhGDhvgaa79/bM/
HDVKtwkkh7+YVhBa0LVub8/ZxEPfWPREHRKZQYwup889esyaSYOKe8sBZVG+2tFa+4iya+KKKKpw
NSb6VeSj8miIe43erj9g7XEHW678ce57jgoLNlGCCgK8Q1FIp6+8ZqN+76eZrOvt9qlZMu94IXLJ
eM9E12Lqz6N0QEYDTwPvs2e2zxeM3O+G91T+v4nxD8PGUiO6GeWJw6UnBYjyY69UDE+MNtz00243
xf80WD+oF1yHYbD6AkCAhx2VgofWCBezI4lGxHM2Ig+yWr19iQVnadjB53eFpV+49vxiQM2yev4B
3B3y74uC7dMpYv+VTOfMuxMClHLSQW3u30eSFzgXcaUv7t6jI/IEtYUQNbOxkmlRvNMr1C+u14NQ
AP5O7AuJeeFDp7Y2GXq3gSJbsk1uxNMUsrfJEKYzAr1nPK9TWQErbCWX0B5f1zFZPOYTZSRtDVqH
adTOkC7Ouexzh5udqCBphHe1xovKqcX2Zulj7dlX/5GEtrLznTK34VM/1uGXvX3vxaOify32ZSZQ
et/6ysQwt0Tn/x75JFP4Rq8f15tBXOvq9bRgcPk/TLXUjKWatg8P8WWGMX/pK+6A055rbqasYmBf
SO5gGqTzBm73/qvDs8xaNl+iiLc/r1ZfBPJAQO7sTRPMcSp7/Czkka+4Skfz8+7erKIq+Zii8q+g
KspDltu6trg5rp4arTcCB1yZQrOtOoAOwtlT2lCT5atP6GzDG8GA8yH+89o5taHw+h/h4lw8B4dF
2oFNV2927wuNfn6Z1jwg6vI6sHWymRkz071/ylBft5rerAM9FiXo1CCwlQyDUwq8/d9pO25LsqqO
7htf3DVwzLjUH95ShhPuhGij2XBgJ87RVlJ3dIgvPMYz3eggHhKyZ2pOcMEIu43hBteuOYNG5Vq8
XR4Gg3FVG4FIUVKnX2Iipfi6wMv0jdU7BvLCfRRQs+ukLHyTx/vZEwCrgGqpEQZhqF+JjEPkQDV4
IuLwrT1Zj4mIc1Ciwm+liVMC6QI0IozNzHqKM9UY+cM/FHq+HGsCIrzVi9DWg/OwZ/UbSeahiJ7t
j+oPiWTi7SeCmqcAn8mENvF9KfS75kqwTLXPGyEfDkSfyQiN73R6d46bKci1EPgQWwJJ5IBCkn96
EzkK61kZLuDZQzull9tkJYiS9UIjlktJQqqkzhpJCU00PefQEM/ax/BSsGc56BT3ZIOwqLrVOGK9
ctADjRzIy4CUn4kzqzGuo1/nSRMDpOX4eUbDmkGvFq44OJquJnkRURyheOEEIxE7nlozufUrhQMV
LSyv9oTBt7UYBk08nsUBJq+43Tu+v5Ir8qyvpRmRZK5VsGrl1EOyKXliRcDe/qeg9xQ8HDOb8aes
iTyTwSDCYu76Sy2oGqXPpB2yX/KVgG+2/gJAK9gk8mEaA7M9rlyVj2Qv5/8dwQgNIn4C60rCwpVN
BJSqYf+a+f7PTkEKdZzTZPTVMZgsZDfTirH8f7vywe0rOEAbqdbYuDcmjMVSmKXJd2it3656emlY
FIqon4r7i5QdPjWsbFzCNvNsxYQY0vckkKT8V/tWbuythN+i5gegatRm9zpJTly3kGp4Q/jg8vCp
o9BwSYd1d8t1gspj+lSh6qUaHl6SUXYPKwG5t568KCT0GjK7w5HDWueQWBjqInjn5AcJKxjEup15
MHRfQgUCvO1bqOrntoaCdJvTY4yJDyqXaIp2UeDEMXUhvCAGzM/+6cVHgapF1jLB10vysb1Wd9NC
Ba+xFSfRG1c/Wh9QClEiQ071FAaBok4ldGN2gNbKNnUsJo4A7/wIVXeS6OjFW2FgFylXmWniwSXo
XXRrPLvLeoSvArUr0nchS4S2CvJF1pywfZ8TYJHY1jBLiuqXGvDFcfQWUyAp0dO0b26rVO8H3rED
+eVh63MBxO7YgFnSGiMmlX9sh+I2VGoLSlH1DXDH/5mujOcn2+y37Be0e6dKSw/qnZPechUIE3K/
A7YMKmCIsjSjcMRCMfHX9a62W/3jpkQUjs/IH1tgj6Hs98CJDfBMqyMmhOSt5tK6UDLM7weptnPS
rWlSKWZta6cAxRrWFWLMFODWzTSV8ol79zAVzpllTyNTrhiSLWmalFRbsNW2dUp8m7IzT96AD92K
q4EHJMs4TNx8uJvmUm5lbVfWbrSnTrvjaPEd6RQVHPiZ9cZMbshmnX2NVrtFL9j3+gWPN2yF4S1r
yj+2rifZaVW0Pr7h9V9Q8hLAkDwalBvcAsavmjGRTLSGTcwlUGDBDeJBz1J2PxzkrRuzhNHTcs+b
Uh0w5Sxi2SznImucsp43/zaWnSngm0vMpuZg8OXX5Hn8XakjtQK9R4KWSLZ8xGxCjH3MeTsoYDxv
SYsHg/Pqi+4DHNot42C3/9yvspefiLdEZn/rHbYiRsaSLrGJLY14B87Y2dGYagHK3qiWGz4k4cZ5
iwOqIzAbcepDDXJJl3MpQv9X4JY/kByQiGFx24ZgjgwB7bT7+HKsDR0KQ76dcwrhckhYGED5q8cO
SRfmCuBHqo6+e/eZpW8smphtt0j4uVF9+L4Z/spHhintrg0+PQsJkfy/j5yPCnvJjuPjKSg1R2om
OUcWVJrljh22IIUziCKY+mDkyJH8KnRHIT1oHNSgxHViOOeUTtohN5/vBztLbHNU+pxLzAUaheLy
Fuj48RI8i9msQsa2DpKrUNQHzdA8rVTsGcSrWnxIUhGLfn6Fw9GhfOYVQTWkP5vUAv5kBAo3yc2y
3ZXrRAIc0ixIgYLFDwC7dmcHvHxLbdqJRuX00M5wUH3STahzTMfHGW4KG1QsYvKGc8n6x24TEKcQ
KGaV4jAjiaCTUEzLUlco3HJj0uZ213IPR5+BCYaoXxl74rh3NgUYJ8LfacLEw5yhyQFEmnZiiXHc
r2TsYdry6opIF1QjhXS6xnE+UJLbyEVnoj/IChWnsC7yTiUWpJa76DSo75OuKg0ZTGKSJwI95RC8
9BvqfEffN2KzQx8lgYsHgUaYCDV3a5kjOsFi3GwC0qKPM2rQr/ZT2WxdgliJmj8M9iVzNhyZjf1o
v6RvIGNEw21y6UXRnaFPv3eHY2XTgO0Mlr3mCAF3a3u0eOjBFSw7uglB3quZVdM/mey8fWEUGmHb
OqTvAIZsvbBI+HSyf+Nl+m+6bZ5i7C7j0hGdSMICvDKRswt2rYByayzrhg9hEKO4z7Lk7zIvH91e
aXDue1iK9XRDPNVe/EmX7/IWH4HSRIptpoYzSeESdX0E5ysRxvsrI5ryzfOvSkXWblabauT8ip4P
xr3OxYCbLQ2CSwXYjt7qgkrJCZn7H8G3Q9mSpBy4zW6AWwrjH6E9e3xhhgvcCTzjj5zUCK8QmbYE
AMP0ug0vPW6UaM1h42juU3M6Mw1Z6rPxj4/WvDE3XkoNqPiARpFxdmdqBRaqM0wJJ6A13q/mmITt
NY6DUnrYw0xmL2pEQdToRfWpOHn4VfcPWSkJrWXqfPMexobey7GDngedpQlCH1srj5FHZ3+Y0iNk
aCIcNmxda6zdmah78cVOYosxJWKUJnt4B+274MMuAJC56nJo/7mdBiHvLQgKXGGkKjNfI4rp1D75
10x3zOh2UTPKrY2hd/Ds3ZRHWRNSHeWIdq1VV9OIyiPwM4dwIa72kxeYNZ36DRHGsmdhv1+5yKhw
da3srMbIbDnAHonSmVnfWtzBuVLbVKv9P5QdYmZ3PNbTwNUDFIblgSPF9LlBLZi20r69g4kfai2X
L93rSYnNcyKMZFH71p+nDuJBe43pVhkUtswtfq0Zk5kt/aQplUuDE4zGLBn0Sc3xr9TH8JIWXuAj
NSjdbfVD4yS5edL1u8FSC646gTaIj6eBEuotyyMotg6QqyLXcZlgxAzIWzw7rcyNnjn1yjMs8CbU
Hhry8XLlB6ectU77x30Uys0JHsqSpw68F1BLsHtL2j0OwqZskXAtxWpGCYrpivX2I0gN2rkN9OFl
R6dNymMW2Hm3rlbE4Mdj9k06yljyLzCFYPbUXvX3TqCFXmq2oIPVs9QZ99V6ZUMz5zNWlsPt05Py
UHOaDrYi0kBMKkpewvigGur9/gokOw0y96RkBp2vAyW6CBear+HkQ+vQ2KcYrFokfAuAF3UpEBH1
B8/fvZ+GlA3Y3rwa9JTa7WjGjkwPdtJJs0wylItA3qyXdW6fBc+qLsnycrDcoyWDu4jq5XEdjLG1
F0e3r7DJ1R3f6jZ1Njyk/rC1+OigaeWUPtc6PiYLcyg0lbCzduYV2hsnX/gZADATjfCZxJrbQqBT
Q64TrGcPT+fAlTJENjElUnrXOo9KjCsrtzyPrubq6sD8MFiGlJw8jXYYrgX7qRlS0g6IY9vXRL3+
vZp+4vwI1meIZRPsv0mlRRYyFOlv68Uj/43s9ZF9Za3l0QEh1Ht188PaE/GeAXDIkt/yeRGiLKvM
MGjR8TUmY4bTIylvHpGgGhPlB9e1Qt+D1zbdhqYmKmyU8mEiXEkCBmPHMh239s96f7wwm2G8pEHG
jBOe9lksoU4E38OF1K5d/M2gBFIDE1kiZt3EmiHkiZjzWyMlolFjyquK3x4RTi7avOsrgGeCF79Z
ogWNyUZUscb/bIOkfxXjsPHG1mh0P0V23yDRlBDwcK5Eqqm9PBeSn/cfokGVYR1lhiQkYXSL7TFF
Kb2RidW8WmqnktUF4dWvLUfWt1olMnUnvG7IQwotez+SuIWgWCiu7SyPPyr+zgXxbl4aGe0lK6HA
YohxyXUgajI8VuQmjFH+hUDTKGwby7w19463PUI4et9B2nMEnyMC5TKiw0o0yHNHTCVzayahWFZK
U97mdzLyWZ+kYg3HGpVsiPUGqIiRRjksgKVlTfeYwPs4oh+6qs8bL17gsomHGHlLJS/zH/mtN2Ju
3heio5xdNHyeDnvtFjEhWynF9vclAzcnpbMNkzr37qowY8Y1R/UMXKUy1Aublfjz6fVncMEbAxeT
tGJAt3S+HqC9ZyflTgRRJnV2tBfy38xbMWdvCL+F/o6pBlkMt3oPqoL06ZCM2hhWJiKE1X+ZJLO8
s0N1QynYZN8qYH60vO6SNJ9ntCG/0nC61OrnJ0r02YGMO5FYTMkdz3r3TaoY93ubFSf5HfWhNhuV
LfdDdcYR3cVyh/hivi/5Reyn3SfAiOXOwFF2qORytaRl/3UbVp3Nw2Lm3CHy9tOvP8uSVGFIIIl3
878uEhp7LrcIvg4jCegYWuCMRkQmcrbF3erFNqQ2H1MQJ93M3Q9Y9HNu2NayBwIbGPaagzOCnNwB
vnKsZn4uX0bDKOtqRjphZnYLfLlIEJxkPcKH4yWk3xM4XbPJUK6OTud7azLjYDYWme1WboW+6xbP
qmIxIAG/wMBshsdUOZI0O14Y43QFXZJJaS8eUsc7FaZtTx72IFKa3R52dwk9r9jWn8mrWEApeWWH
x7RubDjXgmRAZWPK9iFPgCyztIW//bqRVZWai9iHjaVapDu6JJH04RJa/9wiX0FsYewWKkly3fEp
BwPPp2NjvVMG5aT7DLm5ZSpG5k5BgPd+SSERS5qsKdEwPTszI3jM5e9Hh0pauLWP1vPe1yjicppr
eai47m5VPB3s8g4HyFueLZZW0F9WeZ0L9yrOGe40jAdphgefZuowbkN87ov5z6q9aaBDn9vmVs9M
RgnwDpzFhUCw2FK88XRtyNPJpbVKqv+4p4JSRE0f4PcG09squOKP19VClj7WUFSkGEcC3zS2FS44
Jv/ywKM/20uvnI85rwzXst7HHZuaW49bSiMWbT+eZTn8HPaKC/r+RHCCCWMUklwFOP0xTbwsqJek
xYawHjOv4jEaWCjob0oPB47G1AcvjfVOGeuWnMrWi0312qX9zx/lwq1hf61NUG/zy1aaS+BGU/hc
TQBA/R4IDSw5vq0yV/fyuSaXgnht96mEsJ42ZZPhSlCT+xTicp73kSC+worVT4x+9fHoV/YDp9La
BC9VRCdRCPHHI20NUmBn+wb+aRA5lhJZkupxbJRlcIvAjjMHgxpuXQ24J/Cg24TrZ9L9AUtqjoet
AeVO4fe2wpbyY9FNss4QNbZdGQ7jaBXnF40C56QyZM1TCC3eovuhkoCZrBwab+asv2Px59GbyRU4
ujmvtG2fEEpBEa2ji3mlUgMhDDew3CXy1aXjkzo3Oo7eZRFQkQVIsWJHz1Y/o1gJkKMqlWlQMzb5
ZXrQ3j2ti8/Cz7LtnayrPCDeoNvLmfr7mnU7gUmbdFp1WGe7Z27hTfWAabvzBwLSFyqW5EN0DSbV
IIsZGPAcK6IeHpIy/8o1savPdKMCLf9N/4k/t63wA5Yk8wlupIfszPf1LrtmwZ0xNviNQKj4PmUV
ulnRgOr2JQTsoA4vCre3XeLymA63pTN+eF7sSL124L4Im9ruYmVm1+7lLA4VKpSw1pAKkRd3tc1A
7k56d3fGs3s1A8sJ0kOxUksh5Nqo+tTNYZeFB17f2Hvmo+xyXrG4GqNabx4ig13LC4NcHgXcTDg6
6YgmOmv7jR/xMJ/rovEAT6brkIvrHScZ3++KFU5DozNW1G4dGI3JLawGDWo8LPxsvCIPmST8mq3M
IMfTfhVSsBK7B1Dm+t+UqIi+jRPWo/ea+KwBhn1mPjoZ1KVjZFGNVmpISsuPKXFORKPba+Elofx9
wT4eiqR+JMH/Bf8E+nSAcp+ERXVklhi7QRplAWhaYtiOTtQA+TlCIaAmwHkUCoCNbDNXw2aefkdQ
z1uwkRZUhmQ2fvUYHTtPAZTs9zvtG7Jf00EOFEZm4pa1DmgW785bbjt6s0eOl6PApyBTRFGzmMyR
0n/4+p7jNIYB0fffHACYVoBxXreLbemNsZGfFl7hc+chf4rf3U2j579izkKcFrWq5eJzuJiB40D7
+ZmrYOBIX9uEI+xxwOj17rIk3ueUf1HWyMuI86XwlWhdfRhy7id8+2/KyXwhlgU7yGhJCeEck9lj
cvBzsBYzTZgaMSuZCfqjg9Saosej2SPaTmRLKI+Bh9UMQ8+NbgpAI1fIrc6Rd3gUpoMTubmRpvY/
5CrV9yDOv8xRaFF8SXt4uLUS/vGFkz47ucgUFibSnwnNrwjCkfe+ajb4FS1bTmvWHiVK4PyZHZ70
cRhELJK6n6trSAoPFpCaD1iWmd9BS/hvuTzmSuaS6+m4asn/7AYK3Pe2zUGTVeGQPfnnoRV2ZslV
pFvmYHkPYgjeD7E5qvDXeTc8NDg57h/RRJ3lr7IS1fCXVBn74yUatQaGqgMX5W5cMuBDaBkjz+B0
UaRprfoMnglaW+hLe+3kvCuLLSQ0Di3pBVXGT2+Yej7ZZtmGK5F8RUUdqQHnXsDIn59rQeIka1Kk
EJo45xAavlirbeiYyrJZpjleckdJ2qqr81M8E0ASKSzNmSnJRu5nYTmswBmCFvz7gpZoH6/ia/Yi
9PLjtqn7kGZXAD9LeP1uHCa2zCH4CwKzNKxARHbpawLjeJYpMhAFGs4dXoe0bl4XydJwuV1aFNyH
3UtoikofkLam5SzDjbvgobCHCdQ2jF3oZouqSBYwhM1sTFcF8w1EK6/ncsVhOUq7NdRaOzePi9KN
+FQ28o2lL1x1MrtV7MdMSLvMwbWnqEf3PUmirAhPWkoK0jjUJRemJf+MEgPmp9zW0bkgtOQV3UkW
TvVUSCZtUd3bxCin71hz99ttzQqSo6dANEc9s2k/MBrNICM4bVgWarF92jfSn4Lierc73FYsRTn1
liQ0Dy5C3u8HkhZiNRb+yZo9jmNvgAeqetuTZUM99TCIJDUrPD1TwVvKFM+8xnLIHsTpk+TOKHJ2
8cTHzG4gujOBFnxiiQoB0gG2ikz6HvDWVz4WewxbGGnEjRL9AK04g6oI6DOo9nrVWRYmCZKKalUC
gL4XIu8l4Nb1DgoMBnD1S1JToYkg7Hn7WCTh7UyQwZC/QAbJSYFUwMfk9sRKWlBqHE3eQnwPVyn2
Rf4jlzE5URwr8xPWSXyujf+ZHex+g1YOpjvEG8n9gDMaq3Mpd+pZaHsrvG0VWdGoOjrWygvwx14T
o++tOzTogR/ocoD7tjOHMD5vWy+BSxAe1cxB6QoLHMYmTsxPSGRgUJ9ALws0SMiClK74Ms2IlyKH
GQXR4jHr7syF9v0z+2RDnQWCbUelkmZVd7D1PMEEYV/o30iAeg483HRPQwQ1Tfp+d4ffQ6sUnJpB
wH4CZnniR6hfmkObCQt3UOoTJlZ+SRhEZZAWq83kdV4anxuGtVhr5I0WpWe6cevFWWkphnc4OfRK
JQaIZUs4ZNHm5OhzlcsnJ+J7uuEUlFfYBSt+PAq6msVC/4TSvZFPKHNN3d6bTxVSZWQ59g2odYYX
ZsktczA3Gmvn4LxYSfRKbxaBg7y1ShtJ8OQHTCo7cMazH6IoZ8jDVXXqcZLDc4d99EV6jB0aEGNl
CVrvnxLoD2PO1Xccd3Tm9c11epSRVss6vxYoBBZNKtJRTY1+9nYbKmypgzBIbFl5uPDFuQW62lZv
WzczrN8zDuaTjWLakTHmTrDEtSXXQIf1lSwkMkN2xfY6umx++8l3dm+yl/TyOXjZr+vwsmmwWmF3
ERS+NbZosK2gOvRApGaBzG0fGfD2d+XMoWt19fFFi3e8Nzm9H7sS8fjPf5UE55kUM7rH2d4AfY2u
UMD4ZZdc7ozr7otyUmwEcmSPEp52N4YRmc0dagWhz6p/U5LX2xaN5tB4C799FtJLmpvBck2uttyz
RJlFIpNq7v3fMLvPAJcA9qA/i6Ve6wHg1WGnsk6G6FAo01900flQi6+iFUZOZTSReFNISE/Yqvz/
sa18Anb2Hd+bOYWUqDrsrMhOu6FNVyCFnN/ns/Xba+Owi0VOWBBYm0l37giSD36rPOxfBmlqTzR2
89MonGmRqMMlLeOHEEe9DO11KSapV2WhiZTp8dHIDwnb0IlA159Wa6aYPFW63CY4TI2doQwxcunb
qA2lXXEy3J57V3hVAEYe70OPJFsjXFxSIGw1YfnUgCWn8lIVv4qy2HCIuqL1Y0wWxOAmy0kqZ6/M
3/gZy0m0aA9Ae5dN0hkrApuWugh2Tp/mOtbR2tdu49DfPCdTwH5qIlC1wbG5Wwlkg/5rU5A1zERx
OhmAeMyb3NQdFxX05qkmIkBk3LhD4jGKHp/HyrMiwV4bJyIC2zzqi0HQUteD8fgAlxDpAvfNwMFy
xdZS9BbPL6nL4GACnnV1VTZw61ZgbMEWKXsPSZkbLaFTbOTHfAjz2wokEHPcxu9Z8wESjVYQWhEo
pfxyJHZKHFzoknpitIy0TTSYy7FnxkmRgddXvFnJkX7rdj/eDfFuE5U8vCbzbUGV4w+ggn/n2drX
q+lEdS4VnrBXigyLHrxFRIvQ1VPJ9KgCK0qauB/iPu8YpEEkRfIq0ACunvoQTBiqFWr/bnDM0MvP
siqDgpORsr3N3ToEi+bnKE0mwULMjOuYhcDMutuzlW5x0gwJQaivleVW6syEK0qOfmIkSB/65s/B
X7jP6bDX7+qck83R5MfnZMDlR1Nd+rpcLK0AUSHiuU7aJhjh3m73QFMGjIl1eHYZgYuc0SBALovj
+jbsrUHzUi257uF0B9A/wP+7P9KDCioXIBNx33n+KOkWvJSnNkWDQ7+ZJP9ktQHdpdAyb+EHGrov
zKsC1EV4O3CnDgXRyTnbiodrBZOxP4eFmA+nM/MPGPQwKPmWBTBefuOcvRdtuidzIkE2mfXF9j75
gwtMvDP1iulnPTWwy9OWEro6AcSLipW59DUcTptxE45f2RE8CPgFyfEMNhB+VBTK91D70Svgo3t8
LUZNWVKQg9c+bzUz29FnqIpPGN9FzD6X894oHxG/ydcd1m9QkfeVnW3bi8HCbNMlSeEUR+X6JXG9
JGqvq6bc9r92lQKf9NVHw/g2R2y5SdqUqYMvj4Wh83gytdScKsHiRaal3YrCgLkFOQXtLHSo42qi
OzcLF/tK7sgvSFurIdX6GdvKLxwEq4ugjVPWDeXx6q0Zx+3AzGb2MF9UDarHajdyDfMWOAzhXseE
WJy39oWVeV6aoPgVdjSpEeAGnig3ZUz2v90KM+SI+nSxK130KKGxM1KD57VMTOZ8MJ5W94J5w4G/
ttTQht0JnibWe8KgHUEGJ11sLHA3ZvLwgWx0OLwbK8Ee/IIG17PUy0LEOaXG+HSErU0kfm8gYWMV
gggfF0398ODqCvURzvuEV25KD93SDmygx/XO7mIR0rr9wBJ0qQdwuFH5Y77uOPkYY+qxPOzdjdNv
yPwWqZhSyolz+0ud3BP12kXsNt7YjFI1D1WKJulHvM4kWZwywvrV5uatt+5RAhgGlqs8EEAiJkDj
OZcbuRkKSpEgS9sfypbd5YaHmeuTegQd5ChiZ9qEtO0uKhFtYwxjWTmckAf4L3cUVY+uEmxLYQe5
TTh20Ovo8906Y/Oa0Ch9vk9sOLkBGAljGtelXrBK6QvmZfVDZA1bK9loTi8OS8INH000EOosx8Be
TQvJhn5wUGXmcHvmidK08jl/3AFb6Fle9Dem76+KQL3MqDiOLL68oZGafq60Ok/nbs+KtjoP574W
icOT/VQTG0f3VuLuLsGS0uRE+GNlWnnn7b1VF7Sy5v3dXNA83tx8AtMgS5U/8EAH1jDVJTPTea+F
uhcKwylAFTi5cJq0lbGorUO7hcarL4PJzSPAaGvED+cU2BTAh2VSQv9ZNv535/pw323YKf2E11ho
0lAS5IPYmW2qUxH25niWK8GDRaEr6eJaycMudB267UOeHBwwQPGzt2H/N02GXxcg2HjLkh+WR7Ea
c+bdrEnjUEu2mbjVzZh0MYd8QyermHAK0TocHjbVWHaRaCadNn0q7TU2bQlNuscX/vtLjkP5HG9S
D37ajMtQmfmpllc8SKriM/96lIBokiaQOyFwpeobzNg+G8/9oPNAhtPedKwWHNlt4dd69r39ZNtk
EgOi4HJv77jGoMhatQPyj33MeVDic7SzlkXiM57FrX8kZuBNJ2aNI/YMY8+pAobJ3COKOmJCjN4p
ETSyO224G/pBBVk3Dqep2mqQ7RZ0qSmhbFOl6DovGg4HApNh31Hh0qXLyS35zpYoC16EAQvB5vXA
2bKGfcp5t6arDh+a/G8ECnNo7yO9lU3DJOuVlqKJ3TmpBFrHX6AnxHRja9q2NVn2p6pEJolK3ae6
BhTm++YjV+JE29HUrUKaL98l4hRUppJHu9Psx4jbchg6zacJjP3cVIjLM7HgHCgrJSGBYZ2efGdI
qZXQaA94t+yvetu7nXhap6OHlgZ/7sH57z7BsINI9uHUKzQ2f1MPLvSeNLLYQJB0dfGQ157HCHHj
MyslmGlQTKbbtzCNfftdTiViVJ+X2PS3+dZH0fyN8UELkstC9kSvf+cafZv5vjk2vE5ZPMFRVWsE
uQ3coQ2SMnIOhuWVePoOw28CQDK7b0PLbjBmwbmh3yAu8gBWhV21UNxV4cmvR7czwcmpreV+tvDn
mU/urXVo9awsq+xltACwKszxuiWIndWAc2SlrOp1xFSwGhgKM0b7yAV6CeNTLQhNUOpMT0Y9tKGI
kUwpVBnpeeqnhCNg6UDvWYp8qzxpct1NwwGxAJdxD9JLiWUuxMIY+qTvek4rZW9tmTei8vEVrstz
ziXdzZMkZesYANVHHkw8TMOjsJ57V5F6cb8HJxnLuCY445qIcRoxjqG3YcWI4jE+f0qB7uAtuAhu
tcnhMEIDUxQxAs4r/Yubkkrqeb+HZAexOeaEBpWzfn0Cek1If+GZ5rfAKKkdq9sL89lr9NHfTiiz
gXEy45lgsYiIxN8z5PZP8/mihTsmQEFA1HrEEk2fg4SLsN8gM1XPsVI3FQvqf63EjKczMpSaDylD
W+iXqPAt1GI0UTUMr0trDnzKRvSE6VAeMuanyk9U+d4rvIadhTKKvGsJgWQLl/f2eEFFqxytx1e3
bU6QqSRQ1aZB+69V+BKJyJbQLRZTF37ZRJOddFfy33AtkCvAG+C70RyuuHjdwukguc1AigqKJbPh
SIzZKGOtwZM5KRC/V0/S9I/cXLWeVnau9AhQ5vyHXZN7CAn+XhGpqdsIcBnlTiDktzmbojHEd/8b
CB5nO4B3bYuF3aLBUE5syD6/+Gj7yhrOxeQU3eP/H6sPIGLOFt8HquIFjzgvQf2RzyiaK0NL7OYU
aYRM+ZJ7cn3ma7VA5LHAvW/Kt7Q2O3RH467MeLTDdFA3F/ZF5lxIAjMQi1/neEoncbDjuJtAerCo
c1YO6Sue+sxgBXdETb+r9/Oj4CTpuqqSYDMPVN3w2GLCei9HL4MumVw2SVvci9Q9vGQQTUr6XwnS
kUpFQ+ZhKVI6CgugMcoxjSGgIf/rVUK9gEkuTQZFX5Dg3V4hYwLTHAIIhUC1M2iIzQfPR1N3ZqnP
HzGx4SrViu0T/R9sGM7sSrZezy3gVPQQXhEQlE2GfUNegWmo0wcqLAKOhKjTG6pfLcE6cbwjgdh5
8pr4dYSyh1IutBP7NXyQy4EU4jEsD1/6hIgmhqEVKeEBZObD98tExSyFwsE9FwMo+0OBXfEB3Npc
Bno/2jYZQtSUk1LAj4NrHVJiayeGfIBx1e30PDxqAFftzTUwpIPWxWo/fHvFf6z9ZG9uL3WlgwT0
jCL2dMXpmckE6RzfkaNiQUv+uBtoxamBagPVhZ+tcpJqZjRjUTPg7NHig+mQXiZLCxMxI7vgcHV7
s0QOqzS98Z993H0SSo+OB25LHcKW/RfGyYCEan+lTlnnwPl+AFJnAX7tgORnBdDCbihqFWIXkGv4
t5YaMsjSJFynjokCjvAk8pFSd349SqDxAfvGBxgE+1vEvyOqYQAPZEQ53PRtUbErMnplF/p/k5yT
sLNDmYCL7HGq4iasEz5Kgd1HMEH9Ok3cyMO9lH/wy5gzi8d2JMkeRn8TmzLurpbKUStF+Kl1vFYN
o+1sbB7XeG0eixCJG8s1rkNG687DzCFHXauxZ3SsqlQ4JtRCxYBUvvyGwboNc2yDhoO315771j4C
yhieMeWM31xw6jCbHZZqyN5Uq7pg7+Bmif0GoBXHZqT4vB38sWYmpe4NZlRd8AoMaOWJ/bBdO9Od
1qZELNB7EVT2sQMM3+1QrE/+3VR5cg/k9AnE8S3KSJR+TwmPPuHp+Gyi6iV6QM4JMGZ5HpOvUJdc
0/6hOP+71x25jBbb+2eZr2NQICkiwN3x+BV9cVoteTSBp0QEIupKjtO6rMEkFvvMmqEmqfnQSsGO
VNJdAweXZTMLjnNfsacRJ/QOsi+YBJ27ZpgVTH1Qa7thwk1aXSUYzcYPB+nV8KNHFBChQkhM6k7R
IZlxQuvfc9ksBQMm1IKKPjssSie5LSTuo/ezE2c+eaXZEbb48sZpK1d3zKXMF24XqeBgplpPkmrQ
zgMsgny9ITozOM8orNDMW2JOeSnP0SCSBrZo8sZRPjBV9U2GIeydN3bnKVt3j+to2baakT8o1j6f
cI7kzj5lOeK/IVPfWNaoNEiWdzuW8cRYuXho32S2V6U8IszgQGgicPfcd/+Xy3jt+2C4pKKI2rSJ
BjHoK16BmiKwEqkJQlEim6ipO/u5FKHqmoFKHiQktTZvzIdfqXu6JMS2qxXdbCCJOvJJTnCeJ32u
H7gVYFfBkNIzSHtS6aUR9ZKYLyf39H3RxPXXpC5SMAG9pW6PhfK5PXe5vdoh+FDT2dX71Fc4+Fb1
XmCfhkaeiEaYMbEbQZn+vUiGr+cWxWaD11mekRSrYSl+IPuMdTimZ5ULlVCDKWFqTLn+1wmo1fqp
RKVo0RfSll8w1zJ4hohu9qhrHsu3b15ol2LWDO4UDjhKa8dImvcUz6B3OPFCA8jQlwliC4Bzwsac
mZWgEoxwA1Fsvt1yktvVG2fvyuVYUrZbAX/TxE85EA5orPRNwfqLRC3qx9HceKInr4pxFOnspkXb
9fUA3nZN1iqCwpCMzZY7TiCwQoZLBIGDWw/f5Nl5nz56MU4dQEMG0u0+4Qbx0n4Qw9JigG8BcUCS
YxYD+dcPvcLzZBPKqnxnEzKYrQ4T6UE238CzNU6pS8r5H8ZBAkXmPZYBxl9JxQgd+Q/5Fcj3n1LU
GLo0KTmqS6hgo3lABNw7JWJe2W1fJ4C+dauWR8FAl1k9SVgeD/gzBamwRpjC8IVza5qnBwFL85Ie
6ILMbE9mQADDJATWTSNHOfpyfr3cacK+b5BXmQQ/C20KwPoYHpnJ0uSdwqb0+ZQQUeOORxj7iGfv
NrDA8OaIVAywg/jvKNvHjiP7Pte9FqvxLEwCs5awoIDUe5xwtZ6LDgpG0ROl/32MWoDS/dmvyX5m
bLn0a80uXkuxGpysTBBw7c44ExjDS6/PkedwdW7HTHucVS7MHL0v/RmUuiRUcj0LdBXJ/zgSp8ug
NawODBxnyAFzCuf1zBozYLAhK+ERTOLM8c4H2uVq8pi1I5whHFYZxly0KdQKZCBsXr6HDrZznnrf
tHMTbpQvU0S8ge0eHn27XtCKYteMjeUkbjm+CmwqhpYYTgvDISuvwV2oAggDATLNwwL+fCAUqMTz
VLdkK7lM6Jsi3n3PTsClebDP4Wsw9fZ+FBkKaV7ZxoyJCRZmA16YLh+7NYVFooIdCM5l8leuTdzG
pQ78rDxC7ONmo49xiAcseTEN3r30k1hZl8tknP2uNe495toFFQNMxJSIQiMO5jD93PD6+x+dSQ/D
xJBpnYkKk+kqYmd8MbxjzloO7ezrY/jsTEmBGXyHzWPOJbywQZvJnPN+Z03Mf//x1KaVprcyvMHO
8PLLPUk/i2puE0b/g70JRzqWu0uWJImWPA8iWCYFb72Z4FPtrSejjgRg5F3QtG30fukNR920qTJ/
JYKxVFbdogNyKPr2q4kcXuq/zxi2cnNKMFMSzVRsJqFaeTwfYa922Dq67LngIQ2Ecvlq9fnk1pvS
jZCCn185t5X8rmB5M8MbAXz8xDRT1ejh2p91l3UjGGeOOmFjm7SBSj7kKliIHzwIibrr/cZtkwg1
b7EUjevLQwLGd5X/pdTuI30NMRF0rSG1WBwNJFrMZMVgzSK/j0TUOnha5D6c0CYY5dvvAsHQExXF
mBhnTjuZVT64+nODCoqZf9m6s/glEK2UtlJCFVvX0ind50J9t+Dg8Fw+hmx+t7fiC9D/90Muscb/
u5TTi7/Ycv4/JpfZ9xfpwWim/s7rkEo0m+8yTwWeku3X44uyt4FYwYkmKmB9KdppfcFDeS1mCbeF
77ycrsgLgz5wjzKp7d6HGusp85xJLfvU1vjd3FyTn7nxEwCGP5qINzlFuktch+gDZZBLHGa40GrK
4bRApRiZHIJWKIIIycrmUSwNfj8H2kcPDtD4ppaBmKy/HPrP0h21oVaKtFlrfNARaHqH/ZWB8ceX
gvjQiZwOZme7bkuNWS0uBewvbLdJG5ADQNc+nO4bpwSR8rOacItnpZO/vpI/nsO/SorFsmRmx983
DUB/FO39D7b7kGNyljiHCCJ8GXlLwqPD9lkvEQgFaaCSHr/JLDN0arsY7v+Qo3+ou76149UmIIh4
uNG35LMkWRf22ivnQF5ayKQn8bzUAT29sB5vFQEI+6/6HeomFkeuR6kKLsJ9Dz/oDU1EEmRqO79o
oM3GPYe8M1WnXl7+J9k3yaUoq3Y7QvPniVNxP4MgK2CKttauZoktmoSdmk0mFWImU+R9hj4DPbfJ
bIRGXRl2GN8vgcTd67Jy2cEdD/L/LUhlWEJZELOf+Jmv3nO0GVaVUKRLGCW7AuhMSm452wDZQi+m
pf2I+9sxdLptd8ZGUR2cRisyQFvWI5BeDCYUFnLAakApQVpmXk7ep9vDx8rWRK+yUrDu1K9cOSPN
Qe5KcOv1b3bBn/Oto77C+6aC3BqjrD4AGs1HpTLW97SA5rUPsJ1t3gpjbpVF1yhAmEcYNYSAyrut
QJO3XmLgJe4eQ+U+eO1b3mWyM8x7Rw2BQ/cuUqW6HDM3JBEPR7mVSE10iV3tPKu/5H1AQG+mJFV6
B1TPvHuaoQVb5sjsA7n6vDxpvhmqlkGqORO6eKjKi3wsPVj0m0Vr0N0iWpIo4LCq/i1OYiWeHKKJ
DfxyYSGYuD3y6/UTZ0yvddnBRS2LVZa4XwYZC1yiNxbwrGrS6s8BWOWxanCHwQPJX4zZdh7NMe7o
oB1EcTveA4EGdd9zuSHQ2UcAkOCbTeJbVOU9FyIzv7/mI/+lF2KRXXmFeVjYEp/sCH01WG9eDfKE
k1GonrF30aAoIPFujnQONuwQ3KPMWjgv7NoNa0mqX5a6eASu3YWnCxUC5aTfkuSfppzNwswWxxJS
kKGk3uslvYw6oZw27s2GwDG1mQkB3yQi9I3lUiIizqIkd/L1EFZBAqPfik+gw/PM5hC+tysJgcag
RyFlJ6w8g1KUBUjrhRVKmPpcXhOsnxBFn9miRF7k4LbSSIkX067TYZTUA+ccpLB8FVOIqmtQi58r
DZxbtbPpwV/yDJRG7ORjqG7DS2glP+TKSL7Xa8ZmPYzC8sfE4EIcwr/frO4jOzn4YV/CfwYB9QPc
+CZhSucT0I3QrzDKYaqo/hgVpzwvVZZRMCIE5QbKgy2RjEc5nbT7/FbF6edvYbpFAU/vRmB3R4fa
mE00wynxju8fET/9UksLiiQTBxcCHqP22ZDUxiXzDXHT/Do0iC7yagVE+rToaFs3DvZXr8nXqG5r
dtEptEu9o8l3DMj3f39J+fY/kjbrc/Q1GYfzzgypWqkYj3rGZElXp17/tEo3HPnQDtwtO1gA5ycd
8tv26B9PMlCvSNjt2IHDUU12hRRlHMYBCYIMCLv0i25Y0VhNvw156TmWbtdHpTB9F+VNLBrwqT7q
5Ih1r4vDFlErUZhvaR/SOF67sFanCeZ0+WfsAXbfM6SBTVvLHMYQqZvtykPxmNnQAidlUeehbzCs
HMtV2WWtA3mZJ+Q0KjsP7eLl2y0n5aH/lqwKM8CJVOYZHznSSy0WRYcZbIuQkdvdKaTvDlg37cUR
oC52Ve/6uf2Z1JML4bXvPdfsE+zsAhSTfbf+zjMXIIDE1ekDO3QtqsA3ZawQLl0tbEXZ86TlKQGP
zLorq/LF8NtsDNWLhl99YCD7/HvZsjkIqFLIIBBtqY7m5HMelRtN9eZ1RVHV4iO7fejIt617CcAM
K6C6cBRbcdVZKgNkLTyjmtUqQ3XfBqKSAQNra1cGLT1MePDcW3Z4Yr1eewsWu/x6yp4MDnvWxiuk
9qLzePvLobb4V9DeeO+eGxktaiQuwrj7FOMu/a1gp3bpvoPOYNuAqSekDvnClE9jWrf7SbcMfdPf
oTDPQJFKjgCNZJWpKFjUYI6WqXSBOgP4XyAa7S4+kz3trcIzVifza27wTt6PxxYehkYbOfWN2uKR
ihWE5jGtTFHDbz5Xg1XrVE984YqzrAPYMBcP3e4/Ige3B+O7c4+aLqoFuq78QjjsXWdI9ugMn9b2
8ikzVBKbOUnqKGMbOLR2Poef8R96jCoQDwfc/cs0Cb+njC+ngrQRnl849Dc4XHc5BWcZhc7F7wEm
KjbXzXtiEkgjsN3T+g/V+yiqU0ircEjvzwV5AKMlyEr4sa4pMeEbzupuIbgGhit2m6Lh8hJSFrCn
X/YC9id3NJoCo6Q5e5am5f+wCjin1jb/awAdh39TManhvE6YtvN4mQ3FDtebDc3pZuE5rvv82e82
S923eyjvhVj8XilYOhClbsX399R+SW3wFkotcabPXEJdi31xRhCTpucnTyAGYrD9RoqqLMGS5yLz
v5+ThphYJHIlaVviD8y6qigzoRiTBP+AwSAghvYy/PO4qerdyjAp8O/ONp/CFyQUoMt7NDeTWm6k
OVRaXZmmuoX/LeLBwQDFEH60Mn+P3xHVND66Hh2OFUorzXUJDzNhkhRBGC4jyCAybZRVYHqqV1sz
R+ePaR8KsgBFBj3KCbE1XkYsorUedl3EVRVAGLqPewblQq1gIkgERv6js/dbB8491dBnJXhh5uQm
L03sKXWyfUsaR23RaMcyf929Wwix9z/20ex3r+Ll2+dNuJUIYW7MiatLpu45Qu6OG7Efah3mNqTw
nFeBobrSEZBa52ThL8SQiQj9ttWeSAxC6+2UywB7Pl2GYBYc+q5jRZJkPzgjUzCthwmrxD8WyQAD
o9ZQt0v26G21/vmA/nFIlZ3+FpYc2aUlAm5phRgcdNZMMacbxOh4O77UuZk8F8jNz/vn8GtcoEhl
ZvUum81JaRZIvC6dXemsRYs1NbcVD20HY7YmG07B3GsB7a+PVkCj8FnCKOxVE0dugzm5R3DOyYyn
s0grpNh7pA1YjYrQj2eq62d7kUjK1zy5BgEP3s4FqVMRSGD5FSN5bVbvSZvAIKFJ/JvJDKuMFVq3
KlxFtfNQeAGpo4UQ5OzNwqDvSxIgM3SSgkkFmeTCS+12N2lA74gvUA+8kTA/2HCwYCVYVc1J8wTn
lijK3/DAz0042TZODPvr2h+q143MsTJCFcD96mdPdTZ94Smh+AC7KhULl9ODIJLc8gZlnMMn8Szz
1uFk4Y14eCbzJPjluJ63JMM8jlS/e9vUqlXfcyYKnzl3lxhhG9db3Ae5Tv4hTu6RNLlsyr/iEOZv
yAq1VJo6VX2/UCiNIXPfz0HPmilHayE5v7dgE1R/IwXZ1CtHHXuNPIApyXtTx2rO2+hdA56UNrpP
5dshmXw1L3wH62cKqO8DHvcF9x8id40s+o6z4QzyEhjCVCGqjieVZlIqPjCc8y22UhQ1h90JWTBP
BrOnv0WNUHImceYM3X4hNJddtl+2YijLr0etcKtqGpwW+bhp2po2My/au0++98RlymfMb+xUsZ2h
WM3TmliF8RKzXQQE7gc0xo5QmIv2cSZbgzmOI5+W14DsYAuNP6NW3mcd8NKVVlU8Xm/uFukcVsWk
aF7qifaE+o3Cx27Txmfk7dB8W3fyGQuRJQ8rm/RwEovXesuy8y8p+vRBW5vdriS/qQ9BQVyJXlAd
yejcheI3wWYwQkEwLbACvL54pMyvETwSp3MS4ux06NllDE6sIby3wHJtTp8BwJaAYZM16K/PVYIc
B+sS8w+C+hK/dm+mJ22MnkZ3Z/80JIJLo8fgWKJyyfwmh2n7v9KPIwNBNYGju4Bp6PEKt97SieWH
7g9A1n5RnEoBiJzm1HB8nBXpU9oTNOCo+Xt8KMWZKSTbeDM1qSlHfYRmuXJx76VlwJUipJSYB2gQ
ZgKNSPkw5Z8JEOzVkz0ILmvMeYTzpEeLfFYeK43wntw+3ylheQhu4rNhmxG39QDAe2WXytO4Kgpb
vr3j+3oWpbYipcQy3YBbC2lGRSZiOFszpl5i9pVOT1UNp9U4oAFejaNsVU1iBYTDRfYRDr9hqHn4
2Xqx3xeDwf0IZkE4jp11zm34uVXL00YEVzn/Wu2hjHmJr45twSt5KfrTDh0FK9ethsGAXuTpr6cY
0pv34gRlVEHrkKoaRbr/QG86nvR1B25Ybo6e7UzxO49EssJsBzLh/K5g/LWZDlHtOGnIupjoG6hC
CIayiC8+UmInB5hOS/uLjM31ImopUVDsOWkWGxk0h32P5gXc81FQ6N9o2p+P6bMIyK/Bdr4aR9KX
8ljvRfJiaVM4uXiG9zp+jb896Y9E+CO0eMtn+c3wVAAG5ijDvmElAX2Qta0zO12/iFcrEgPciq5A
PvoYBq8l/Nexv2pHV1YyyyW2AHVjudA0/kfkvD8biaE+foU80xj+t9hwztFXdCXdXjccQVsiQSZy
3vSjfLwbrH/BWrTLXjRbLE/lNoYEA2O5UnWhZn7i+A7F5D5CAQQtaHTknmvg+RQg0ESpM1RBa4Ma
QvBYULOGqbm/kHd3+Po7f+EG1o9H5qZ2rahY2sK9gb1y/H4WgHBReXezmfOanGW6+Pq5m5aJGZHI
2/LdvELVj+cvmMBP//5btY4cATAOZDxsIEix7eEHvRRQsI2vwG8ktSmFVDhiG30NKsbBTGcuuLPQ
IVhC0gmSotBO1HAlt/t2T9Z3je707JR+vVxE6TgYa28qBPoEAB4vcgXe0tDoyeyW0LIRXg2YMtl8
ers/gYYfrEQyOZlPPm3NGe2AK2uShWhNoW/7EaOzZezIgp5N0VkVyRaGWIv4Nr0ZCBovsvv6eJc4
7mCWJGJdqOj00YxVHr1V+v56psrhbW1OFgcqmnAQ+ALnyUu5tkzWlI9MlQv9FFaoFIsx8GI0aZ3Z
/ZJrbZUFKBTQnH1e7C0JPLYkvoQiJ5TXxE9nYErpoTvC1nNxYiVedyXVhaWkqO5+0SzyA8de3vTM
WJdB8QGZYxwxBS28g0myWh5mjfo3HxjtkVbWdesyjaAgqhpY9kURdlauz1vi/wijxggtnhtrlw52
MxDnMbg+rR55v3P/EJsGQ4+yw5xfj6qDu1tybjHgmw+L1E9ctFAy3cLCHneLXqvaLB3DAOiBImql
IaFYGlZVanld4mmkZ7shEvf7gL96QiLZH2xhX0UzujWnvJPMkDYdLzbgo+2pKt4q7wAM/20N6Bb0
IOrVFyQHr6HJ68Y3ibh+DxkNHf/SmfPF3aBxIw8LWChuQZSJsWW1slC0XNs8Qmdy/2SE6oBDk+S4
zYtGc0TUE2kgEe9UgY1jwf8rdqoczzDb36uwyvHMxhos1dtWHhdl7psbdDn74QPFn9QwJJvs2KOV
f/bvFjFKlq3pn3oszbA5g7XTQrkkkumgukacGePx0e4tMAeqKN5YNoJIo/zmxyGQSxJF5lLIEh6V
F4AsJAqS9WRB/SCil8vT42fXcoIykpzXL3LYIiSjSuIbHINRSRnLds6amo43KRzit7yvmJ3w3Bvy
JUbOCqYil2Ife7YHDwa+DCJTT5pScUb60F+6zfqvAB2gGPy3Yu7JrkT7DrBIyUIqDzuSOVr5fchi
fs8WmIou/Pze9WH/Ho0dBu1kiUgmVOmxnJEfh557o3BAHrozGdg9rT5LPpEL7APFjTICbHOqUroH
ZX6RuRb17ZEJpnVGbNHK4tyYntFquPHhEnSoyppFkl1WHsXq+0V5OZqVUqeUF0oj5oQ8kRZJkdMY
49Gl5r9bZP/w1DFG+F1Py6Dw8UgiNqgsloqJms/izHgW8f8A0e40qjnXpoteY/2oE9xNhP4gwq8D
EZKxSeCWgb0jSSpxoWCXFg3eX2ycAij+wj9WRlYT2R3aAFpbRJRpGVS1MI0UFLdvmn2N2PXJj8Ch
0Z9q82AIkVNvpEwsVSdxNq3vShYM5YpASxUcpFX/T02EWW4OV4Z6Qv7PVFSH9KPwS408EnpCbxVD
o+V+4PXETwmqtueySme1DcullT8giDHGPLnCNmOqmcOc8dA51BAIPD1ryxPmxuIxxG/MQVBa4dG/
pq8peWyJya26z7KY8OxDbxQOUyr3StmM1y4CJkBexTSofyIGgmIljOu0xZNn4hh0GnXEBJaeSruy
3ed4QIqE4676//SpmdGWr/7pzd5p0dFkXxH4ry5ZvvLm5ygIWoqpojwEb4MIEDMH3M/MCTRfKJLf
JO9P/EehL3s6Zdg14p7N0elUGrDdG6FF4sWBG4iyNtyh2+kDUYke8zt+p50mSVwF97nOgrQFXuUe
HLoQgDu2cukfdng/4WHdLrI9gwmMMnpu5/GpqAcuYGu6VzbeYtuUrIj13xgQiaoqjGb78jwjlAz2
upzU6UCZccb+o0MY8wZjE+LsT1gk2HxTp7AmzsY9LekUL+/ZOy78MF0Cls7Bv+HMvyZlZGJdbYWX
2ShOxlX490q6DpUOpdIXBH3SRQOtvxco4hOhA6BKmdO9fZ9EVnPbVesQBeZ34NweVYVhPEm/nGZ9
UC3lgzVk210igUsKJyll8+eVMrCKDL7iqk4uxGn7MA5GHL3pGE8Hi5stLFRUbhD3FzrPFVietBCp
X3rqkNi/1Vwz+wX/SNKhqVXMnorMTHwrbCQKsLiBOD60ZBARcjc5wq09pZZGsoBDff0TVZkn6uTS
FtpXK2tNGYp39tSgzwM+LvRPjtRY/fRAy0svcL8SDJO4wyJTsBXbBROJckc0/yqdkYrPaY1BKS5c
XTd5e6NphvLRL8iEpLGGv6QBAAWtDfr3hbd8d2EroGG084zQ9vAj+pKG1aSiWsprygKA5H2fsUcK
vpHhKMfyCaVZ9B432NNDDpG3qCcP5d34B9zOnwNVPkNGz1qOYbytRMeBRj6kdS1HlL4+YCVEGofg
rICxaMo8K1Zre9fi3bNp/EsG6CHficNVS92nVwf1zZJ4Ji5NC6PCbqB796Y/QlsUqVEV75HpSrtH
coqTNRliLDbuTlXFzcGNfiDZOHZJwe9wM0ivmtxdxTXZaKWDTUNcncQlAYPvlDf0a4O/63/vR5JL
679Q5Mxqt0r2zRUNyuYYGdV7cd77Mitu3QVBN1btBhgsaU2azjl7R03QLxtEdhcyHtbo151qLwqZ
Zkr6YW0AvYnHXnlfBBHR1Zd/HfxC3yXRq7gE7cU89URLTWq316H4er8q0Sn11ungBTzI8yPz7Azp
TxXJVRTcHV62RIJlHyj6OOnJzafBC9/3mBaLWNu8HkAIN5aZJQXoiHX7w3i4t8UEdodrhEAQlab3
TXWGI6w6KcCwvGEZcYbPX0B6r/Gu3KCB4j9vBtibWL6IJx/IAiVqIMBsWIN0Y4oT5o0wx6t06r5V
AMaeTZd2U5/nDPNXgkcDAtRUoEnGYSNsQ/rbWFWLSSJOfgfa6iB3IwOslfdSvqsAczK+Nqv/mKUd
AlHGqhhsbIHZFrITkqCWpUcM7gyv5E/pQpR5A8zDemOqlzj0x5JhcqH+7lLWnLfwtBwQd550DMzU
Q0EVLshGOI4DqgNK/djF/IWrU3ODZz7aWW25Tbc00pJqOSMfV+gp7kEQVArEccOjzPH2V3ag2Mcg
i4fM3dMnLyectsiR4+IcOx86eoyBuGdHNhUyizq5WMwN4y6zcAZCzyo4z7o2YLUNQut5WK9ULiBZ
1DBFGx/IGWZpedJxfgK+LTgPlPNhP2LSiW8Fv/2G61mHXgJVd1c1EKNm28i3XU2qv+dXJ9OzqjU+
NsouSKX7RDtYY5ibzNuf57ZeiCNPVK7fEyvIrBvvChV4NHnXbWcQEEt9Gd4zF5pIenEYJ9LRpaxB
/dIzrfIkEQ/3ZzhWGw4QstN9AqCWOkm68gsFqAw10OOZv3tqjVF0+4oEtdSR3d+ykhINZNjGQHPa
bQKj5XDy5WbKt5k4WUG+A2q3l+SCHBYLLL/2VmWCK8VKnNvC7bIy+qbAgE/GnosjgkpAri5+Ry3K
9cc7Odbh91XkgCcuJoX2AYE9mtm8NG5/6z2GknHl0gczxe4WnvfVxIBCN0h4CLpOc5mNmwPT33x6
O0TtZrSdmqpKA/iNEl1lWB9ez0Ivroj1rWEgFnimany5XKPLemVeSzqCZLnFMoEJfecZXvJo5EgY
dnRN+h3pvYjJ6QYvaSncy2XxoxTLdBiKzxeFI3JBcw9R0uRFmGePpwmJwEi8JP+GOJnvDUDR3NdZ
iVMqiC4vlPEffSIPCiqx3kxrK3cMHawu9M5XfhZHVSyj86bVKUPcKXT7W6DoLrfK01A7ovF8S9pv
/0ExLAo7veHEXin3c648VWF7yfdZbPvOLGW36WKyXmbUrbxmEF0Z72OpHUu7c2ECZSYxwLNzNVFN
VaHVDjtwjsi4etPbHIxMSDmokVhbuvwW0ZVaD+UcR4oLsHHlLKneB+e9fNPqrqOZx1d+tUJ5REW8
GpkMaYuvquAdoobdt18r+Vsp4vAzFwv3ph5XCECdCPR/wfi3gGdzsuV5A2sQHDxwktX4YQJr5CDU
Xg5MK0gY/kuiA0oEcwRqjCizxOi40UX23HkHw+jtKwIcFdwZ2Uot5O8C14ejIRP67jfde5nYErXg
jPQ78FvQytAH8EU/G2OyzMZk2taBGCHMKjzGcL8q2FQT4xrRllfVBCsqKhWF+zU0gYLf/d+IzvFf
CknWqA+8jP2Ht0Vii2lcYHT1VaAG1GHJbz6HrLbrCazESvj+A+6yuzPgMe3oIFm4wXcmxqfgo2jA
9n4NekIktEGq67syLeka886faDmJhM4uTZt1H2QHX2/AMDxkNgJpZHMS42Je2kGDLrKvee6fZkbH
iEXRPg+PoSDgRa9f0vUhQIA4oc3Lqk64slec1pCz2OYli9+esJYi0qlkQDsY7y/KxKdw/gVeWn8Y
5RKyHVi9ykLGUoaA2mOoT0+g/f8dshv2oZsQ4auQp5OsYxqtq8MPvgR5ymKCg2kYCiingyKQig8J
Ss93lzC3hH6V9bPP6y0o94BzncPCq0cxI5wgfg7tGEN42aIxlK1CUtmLupWw1DNuEfsSg4LbaEnH
8enUBaU4iXVjiBY3+xiMVMpK+3sNG4T0to6Y2JzIMurIfe7hYo7Dg5CeNjzmHJPMVg5OJ2KX0T2v
uTB2NPoJBFgsERifHbjkHhUwRQ0gmVQyjidkhzXkKYn4BFgEIbGczNKlOLsn0ktr8DWf8Fc0s/bI
dR5Ph1bZ7xn+M5K9t67ROwA/Koi3Aj6lBldRiUJkA5WN4QiE76kG+5ypeFZk3r/Js9HNB1/739ma
VfyBQ4i9Lcr4jczfZZNOLNwhteQV4lKlNzIMvMplCFCbwtBQJYmSYRHL2yqgCmofzeZNLF5eaCCQ
QRu43sjGeMVp6sC1bn1D1foICbBv2UBwm4DfC9lU8Fb3PPdPjBOy3OVe/qIiI1UAx6lZnsa8WGKl
wM6zEmFn10Sm7zFSOKHjFXcSdSdzpuK4qNkyfaSfOYeES7IHslLDfs+bZAaJQ/XMt8ByxA7MOatw
104sRZJyCC/cCdGAEkOH1NWJFyyJAML9nnTUAo1x78WmO+T5DAatyV4Hwx+giA7aSaEycmTWckBU
HjQYiKKjVsW9ghfBu/nsfnleevyJQ8YYhd41JfO0dWOJfuDDNvdl5nZelF+xIY4JmlvBJX80CoXJ
EBYujrlba7bwNH2bznDVCDeRQczVuAxFr8hbOh1kjX39iLYluXtXdeB3X1Pvh4mbznQO1+CPF2WL
vJtaGgRahymxQZOaaWS+SGjCGk3RrYAGGzmNVYBn7cqRIYLRh0qe/i2RXebkYVa/RreyRBAKDADR
jiqbhiMKFaXAZl3CIvRFFx9IOpj3Kbu4sQ9dKzXI3q4BxXVIDs8AbpInW3JiFHSvx2s6LuWfPpg/
nHXujvp+V6WTEjOCaT7FycZWNaBLHq8h4jndhJDBm6ihaAB8k08He978SdTLYhpJsWZJeHpZ+KGm
NI4+B6C7vrwAyBOYxUMGhee+vA53WWiOHBQ0HyoHC9+O73lu1FcGGuQs72gXW7KXUq1F9fQ6tTfj
cCILvv1VjGtwEKbR8h7CzYxCYlI+/g4G2PPUjppAza1i3sNg2A5YVshKJhGyTc53i8tNb1glJRUq
MBOAp3NU88pQA3uodEIsaoT6TBD+vFY1RKGKW/lNF1JoKiziEMiVnqzBdt6Q0IbodJUDD2apuLsv
rslH62atnYS9yqLgQ8zjMD8PnP7TlBfgGrYQgY7R/cHMQM55wPFBdwfL8ezKWwkO1/rHhfntuBaV
6ycHgNyBgKGF83KDtovWyK6i4lYmb4Vn7difCY6pnAIbRZWhS9VEprvIVjJg4JCoiKFuAwVaW8Tt
djDiskLqXEI55+MHLxHUreR8vBdN5k2lqyOdZDR2xY2Oe0dZF/wov75eTQwJ8pFplHJ33QVd4V3Z
W9dFrHBdEely1cts5E41R2i60Xn3wITXtVmM/GJoMc7aiHa3ZSJJXkm0sND3XmUZBOl8ugy8WtNW
qBXdLGrQH2tn2apRKaq6qndOuWR3lvsKd8mw0pTcA9ziN6urafdXTP9qevtMarx60fv054xog9lB
9q9CMu0F5gTKXrTTf32wZa3BR6aUZ/MlzNcu8CDXBz0mllfAwQLdMd+S6T63rFk2XhaBrzFz8tud
cVvabGcIl1wcSyURI1u7EQhP3qMc/3MN/R121aIEGKMBsH9spGa3I+Re0yLUpilwGIZEbnMMDEDD
4h79n2C6NJkkuLc9x/VCIuHyj7XVlKKMLYsc8IcDu9cU4uYOpO/Qp6yrBilU/hbrZmRpSIsK53xx
BWfyY4y7JWjuxZGLMEki8Y5fdwTZ+GHHBTA5Psz7zaKtkx87AUfA+I6oclUD7FRdcb0EnTz6fgc9
g7PxFiE9TQ/X0i6ms3tK/khZu6htCabcpKdHmvNQEwbq5FVIvTX2PCJbeSaUu0Tr9iiHjSxtl26M
ZH/W6uQ05pLrgNdyL1WnuNaVcXl4i/ftjPGtIlslrIZDrSIugBdoJQ3oEe99yoGSTN1bsTiDvL8/
FuC0yOKurU1ghUc+jiwccq2R3YEodQHKdmf6lYGwPpUisaRWQZuDleIj3sb0RzJ5/sNxZG2T8sih
nyXBcb6hCcQhg3NhbumFq3prMjM3xmXUjnaf7cSL/Z3TzJDHddqppPX+G6maZXNVrhanQpQ6ARyo
Mb7VwmrsTgAU973S0CxZS2zi/Ydm4DpA/ySRLWJMhcG7qw20SmFPs5zKr9V7THU/B9eG7Ql8pkBC
7ZDOa/OZT77RYYWpypNhgzi0coFB2ScdZVW609xY+aXxVrMa3JO1e1zFgl0uzxgoc3TyQFxOlLGW
aIXt+s+02iJoxLXLjkevIz4Z7ITGGDNKJwVRan7CnIcB+sHx2P77vWEz1nEJSNxmkzH/j7qvL6pN
5RvYDwb6YpZyKh4ckEEWGZ1weE0IBFMeTc6RopmrFB5T0YmpsWT3q0ph5LuhErThhidYsVG8RLdS
MGmiIsi95ttpT6A1/RsnHT7OsKdyJpc7pwYbwPZtoWU0aXO8c4BNKvPA5h7HAooA33lGU6B6lPMf
e6CIpT5w+rSYgIaeFUgcXugk+mQzt7xgAI7CtroGXktKx5es9TkztgBoEhumtg6e65wGbZ7pd2Pe
dHxv7AKlgxI+qbNj/CsNm/nVJN+8LtBx/36P+wMp6HskO2rlhc0WxqLrAVxZ+xElmKpy2Cpe54CM
GB/PsPNmv4Fqyvzlf7clE1KL1M5mjSSFgnKO6cs77EZk7l37+c+d0qEVgH2py7R6LvkEF/hpk4FJ
kHmAAbl6IL9IRe4rXYUhp9T5NK3ei2Qe7kUeX0ZGfl0d4B3Y0KYilldOpdWQClkhN2eiZmj8MsuJ
FxY/0dLlfc3dxsr5vL9qOqDmkhV3a3Fetjlp3DoSZP+uWUgEDqykvX1HddzsQXAi/j/ejuB35P0r
z/KebeSBxHPIkTaX+SJEb+oY1o+0DFYWb5hhSU4DcjKKA7hN56pNnB3PBfZEmEwzu4qo83v8dxvp
KNsotd9bfuetm0RmkdZL7mY69uSm1xTt6mheEEXmS05Fbum7seLW5d1aFfEPOigVRhowHMdpYH7E
pgWG9nv+yVaKwdQ0gm9IEb+8HTYgbyrLF/ejQ8zIwyPzJcWTr3pXBtPnqTfwtYs0Y3s7Wx+58IJW
wp6C4kEj1aVIfboq6Bh0voRnDtG2ahp6o3zlTdxl6B426eVHm+bzt1O0QY/r8Wt+lA74e45ItD9y
0uUm5fLPu0GDON7j3hGVlhJ3b37BmzGxGMfzqV/vPHMP42GH5jOXQj4+tRvceNpx6XkeYzWu2yto
D9ey2ucNsiiuCS3en4w11hoZgB73+5Dp8TPB3cMXknT5HcLXJVE6IkRDKHGf53sR+n4q00cXKzXw
Kvrecao4jA2Z8z6ruB/HVocMg1mrZWkvle62Fncf1+c2rsqmplvJZsSRr6apooAOLaCbvjiayow0
L2WM/Evu02wCgM+UMcxui88/G4GgjUMaN1xRHeRMPUntx7vaqgIqcKDb+yccK8aELIZNsBpdwXAE
rtu9RJgwbbI+SS9wCyOyZC0tAKPg2TamOUhvwpzVmMuh0jHZ1N+RBXzrl2fRPpf0C15Jua2uJNkq
765VL7kG91zBFMFUJaSrdYdJPrNHTRI8hQdkIMwOE80UmRLHEm+ciC6/yvm2trWQw99BVSWGXkBr
KEQZ2Tj5c75J0wgc95p0cBPNNk86MJCixunvAyP2HXEwMrkdXZwdTJvSW/dBASIuC2hw2R/XnUzo
/yYMJ4t8oVFRlA4MzW7Pd9/TO6Z8xGbBhmePoEEXnoNjoH+pqcSdDjBqcfnrS+fwchYibtMU4SRX
MrMH7WBE+tigVwEPwl+I9EcGUeNIFn+387/xLkJf1tdH/VCHcH8/2/Crp2Mb45PwpNoK2cZZgI5i
0zDWHknclLkJrlTV9TcxusbHW50mM0FNhZqCKfnoXdkBGdbuwPtcqxkhfkduoqvWEeKMQEm1gPSX
/fMUhl80LFaoLPTtuuMs1zEfMqYpG2JPeg5yaYhPIBP4Y8CaIuuqBFuP1WisEwKfeX8rIFi7Rm26
RzfrDWmR75tvgD6Qwx7aoRGRz6qvbrOzPXf8qar26NyueD1BOlKhP+ihSOWlsvlXvy5SZa76nEQT
ivhPBFv2331NAq4tYSIVRBXNfj2BKQKaajRKIhfBYWVKpbT1VXuV/qI1Bn56qsTa09NXI4yBg/FE
Vra40a6JVGWP0SlrVpobCtOabx2DkdC/z2tGWph8I3DCT+w67r0Hp65ISg5IKPi1bfOrTf+AMZ4m
bis8MnSYSv2B1jcDsCGesoh5ZuzLmI5F6oPW6oabGoFrNoCpYr7qoPF5dMRsVHWC0wujLrQYJw/T
8XoMUzn2A7MeayiiTvjbJ9Hop7IoQ74i1BG624L9XSbY+NO3V3t/i4TOFIbQ/EhYfh8NI9VFBosn
yAneCB2FLDY7FjHMnn+c/BF31wcvq6FIcK40jPcXJQaQxP9VxwOnsZ9ruS/radElCKOcvlObp8W2
IOgakU8ff4t5ZDMOGjGj7/p4hzfjbOiGtbo2CzdJcRVjXWMPb3Py0mvb0pM/umhZ3kc+YAP3tlw6
7QOFHML5SEsKqOWFKdurboH8UMZAIOLxExTpwCcGYzE2SstKaLPNTaA+GKs1IZJj1uFDel0l9m3S
GaBiZxLHZWYGcGbh0wc6UlE+dHo1otN9i2D3kDIDjJW6JmlM/sKbT/bJoe1GzEDpo+9VNFIzh/g+
SNOc0wcjGPkY/K2cGJgp7xAKNn+h1uU5LG0Q8wyGiAA25CNruYxWmvrTjNIXDNmIgA/okfJvdqN+
9+JxAjdp8h8+nucZP/bbqt+dp64K1lxfO890BF/7duwout2qjRkcK3PqmzSudD8A2qiMetCQcvL/
qa60wmK+RKhweWp3bvZ5b1f0GOrg/AMj5CdF5WPrilpWORSdpJvdnF5FinaByVKYe0ofXORKNaiy
0hPUjFLqE5GAOLD4WWInscVYsGEjc3AriXO35I4hJqrC9IqpJjcW1GwjlUBm3m334aPPtOsfYcX0
aCIH9rePqrGPIt697omhWuMRxIv2EUG8vZu78sqD3HmZ7s3fuLcCvHfC/jTTLVb6m0k4J3h6jKBS
u6QlJR6fqDBaZHMU4WiOmHQ1ioZShsK2jMU0pmU0fkqLfAa/gXg7Is6lwLgsrIEYqJ1EJ/uC1Lke
RIhGbvKzNpCynSsGkovEbo9a496HBzTJ9Ib0mJNI1pYT5Epm5HN/Z8BK+NzRVoTePibqtxXw9BeE
dO0RoptNkOFwRL6NdxA7/B6DWTmf1gkjGbcn2OMILXZggqNhw4nX6k23GnW04BWEF6HX/csLSwB1
x8tZ3FggKrKEgESP6M6t58D1axy62fnFC2XjJX5Y0J2x7Lzp02+W4Ouf3hrzQLLaXPacfi+CCyC4
F/PqBT7phe3ZS/XZTjsSRqDsrHchO6ZOfGpZGnKeRSqXRwX6qnG1YfnrdWqgfBQ8pTn8+idoOwQ3
1w0+3fof5xdMFV8eV7lFD/ai12lAlaiOZj07v/hk1n/iwciXHGv419+ARlu9imrhmi+WqOdXdOqy
c3+2BsPpN/9phkM1eTS1Gl4jSi3Wz6GUd1unyanSz7WZH1jte4rvjjPbX1YbxR9d17sG4Mf02/nH
tAup3uZ1bX/lDmWU6QZ2PruJYN6nXcyeX0pnR+mFkhy8+DjTuJp6Q5TRieEn6ygernQpYwa/Z6/0
YomuhY/mYbouDsh9sHV7kDfipo8dKoiVZ5eCymuP5fF/0POikyXmc6bzsg7i3NmqeWoICEx1w6K7
vVRhGXiIfdRc0tVSHPn1hXZifbk9M1Cpp9TOWa4bHd6gs/10wrzOO5mMUoEBLTAjHXoKRgRKh9Iy
slNKKbLtzWK2WPtdjopXhvTOrKezhIANr4Ys6aOqftXiLiKj4EFfxUTEhUxt2UtkyGPnNnB+sa2W
oHfnDTCgR2iMdh+gmKbw47odyg6r0GsodWZhX/Ev5iftygIJc92I+RkKGOFomTU/pRkHzMAKzps7
Phd4utpAmk5RGviTsRYoDj4FNZswSkoFrY/Khzjt0nm2vbzoC0FMtl2SYNa5pL/Z/vVYAFl9NVtT
SBLbQnw4LhjrLLhBm6omTMpFEW4rJm7ZooA2YDBYeBV02MUiUmPaFvcmbwhwNBwG5nN8qm0g6FVO
KUzVcocrQqrT4muhLTw+vQB4E/nezHUMZgqEM9+i5DJ5CvtZMIctqUUOmneCticztqtNOYFFa6W8
WgjUf+MQPfoZGmZOf1grwRQf+Hgh0LRrdCF9UqyHBZnm8E3ITzczqD8q8TMVqOMfdSEHe3V1Ta98
wczQSQOHkt34aBk4UhBXQw0v00/xbBZSoz9/Mfn4/ZXhT1PcmLbrKaLGLSjfJSjh6ZtyDBeJVrjG
mb5a0ifcYrL6xJ98c7PjrZmibKpSYSeWekEYX7qzF91cfA4tSAf5D8NuTBYZdvm/jE/K1v5eXKs3
wdJseoOUNTcBBd1U+56nLB76KPQcR2+ochZ94GHaAcorL0Uh1L65ylWWDpPnkkLNJNgdbRV1Keus
N6wvy9uWUIHMPnGWbNjeILc3kTVhKdtZyg/cSr+Vp3dJw26fmyX+d6DccGGcpbiBg/P8Uvr2lzrz
V95U5E3xegt+wVOtGEZesNdzSRSB2MOk1qwZYq+sgBz+1BgxkmzMULMVyUJ1DK6sST65uXTHzn1s
2uB9YNINH+Lzsz4HQ+sHREA7ViF2fum+Ia7M9u9AbqwrtrkZy/4gIy+4kjXMj3dEs87SuSrhCnw7
1915DO4EasvCAOiu1Ynn7+Ktd/Yzc53/Hc2AVMFylbnEcM1eZdYcL8v1a9rkNGpeqH7rzlRbrWwv
Y3fwqxyzTUborGk1wOe6xDf7nMP/C0Jsd0WXemevK6MyPXINb63Y+5CGQ9T9tVtum7z0pjKovwP5
PdF/kAcOvkhFEr8WPxlM5F5+Gbhc0YSJRVujnKLZ4utUCk5xu7MWJmG4ABHvbgUzK62OJtKouEc1
sy29kVdel3vkbs6Wgse6PWrUfYTMtZsw5i9HMcXPd0AfuDhNrYyWvg3SwBvFpIqapJKrAhqkZVZc
xbgA/Zu2mzNyG+W21SvVnObucZUr9nUlrltu3olnjHGKNqL6rz2bYuBingFn/2e0IzX63/eZIXdQ
7urv1qgdtQW0dxb65hvEESp8RvuX2IDjqVrazH4z8ikGvdizeArnsHDqGS6sF2UUOeRXFimWRurK
CKyevdi1MsY0h01GUXoW504ZNnO84qcCpQ6NR+YXjngEHYvxjlxNiLXKdzoy0iTQMH7PFp8nkNq0
XRwNmPkRtK5iqXG7jC/Ta6BXKXGldzfNMazBcASAHSsjffK/8uQu/5caqBtNQt4jQkKrZWZhL3ML
ycWWMTqM2ThZqN2wRvBdg0AmCLjyvtOheri1DDsCJ/xfmrw5kfLcqDkqc8gcASUtjQ5hYKRerpWn
XQgJueUV7/ym7VYyNCvSMUK8GghDY3cCZ+4ciyqkQ38pZKgwcyPeNCs01FKc9mITlLjHoGnBEX97
QhX+TlpW5U22iBxuo5uSQfjxMqHrDvwrEKTMB5LsJh584EslMHZYXsmSXMi1RELB7vrfXkl7aQ5L
LMvKsLGFu0Ls9i/+O7pw/v7BGeqAKcQuGiPWJC68OvQKkMO66WFcBoVRmEf1dVzq5ElO/NiOJPMs
vZxMJUcP/aL2JZwNtAgdVETmPYoNycppbysZSMisIhGgJVnjnyQYZiU3OMUltUKW8/sn5uqdyUKk
qzXBapqcsry/jU0lrUQiCmCWm/BGfcx30+OxoFwxy8rjK7CgIgVP9S5UfYcL8LxadWEtM6d06t54
z7mjj2LXAt1OtDRbk4A/65rE43iwrJkfnS9FHaTV3Ukzi4EKTbXUml90TpsNx8erknIhHAsVYPqn
D9b6T9E5F/ebNsYIbHh05eVgoFnNI9ddryftzg7+AI/kFTGcyClMT99lA6inGlVkzggpXzjQRxyj
DFt7F/KP6wDAT6WFfS27gfHmQoQHILAUpwfnn+xgRyYbGuByO4Pl5IbjvLDsLTTDQppPBj7SChGR
5PJsjZzT0+Pk89vBgkRBDwK+DrHjpB5hEeRgW121nJ1saVyB6xBZU7TLKbfFyHqREGJIzjUJKCc9
FKc+DXpZJkOAZGzSi9iPXDmI3k5+Iwt1QTp8LhsWFZJ+nN4wRae8uAbEM3J+OQw8QJAqKXr317Lp
qAryZUuivRCtPw0TK4nBlWmJ1RFqlfrOs1aSCA+Keb4yAzKNXT5/S+VZj1VgkPv918qG48asNsr9
S6nydJIyT+Jr9Xm+1obhwpJzSG65EcKaKY/PJv4H5UppZvEV1MMdW3Z0MdKkN394bcEPaJzX5/qC
zRHdTU+L97pxFKcxIfOMr6QoVR9dXOVp20j6ob/xjR/70KbcDk1iqa5yy5qh0K2yzsEd65PT/ku4
ryIIdQGhYztv1RrfzhTZGjTMcm/P7rDf4CR/0uvXQXd1lD/SkskTV3/8UfWexX7Mp8G/EOPsUWfl
R0na7/B1XMqoGH2ikh/aK3DntL/qXCm6mb1iJhsExMcrBfJmOZU99WjDVZLVSr2xh9wEo6oEZXuX
nqimjqHAWPHkLQahgI9ptgrMCft6rqQKiEVAbHjDxAR6Q76RzOVzTxmqQkZR7QNIqoKLR1OCBkQz
SG36uhJbkq5jQw/pmOaQ71YOvZYe+wJIFd4v/yqM6sO/3Zkjm0X678OsqElvBFaz1zBVn4g5UIpa
D0wwM0P3qcM/n0EWvFaejSR0kFcFE3EfV1BhuLoUv23XUkUWGCUWwf1tVnA+Gxwozcvi5uKU6EQ2
oECljCZQcVu7+rX5vPCwhJqJB/aq92vPMreaeyZdMJgWhaXBmFPK/b5447OUnklWUrwIIMJM+QAX
pOV5iLjubPP31ae6WcEaXt7sZtt4mHvxnSVPYxUhD0sZATAuIB/jR3CxVVN6dNVu3oxXQk6bXAE0
8FrxlvHjba0oLie9KChFS/WUph7fEjny4b+wz2rTg7WF3PAONCrV4195Cyej/n7T17W1m42W/trq
xO4RLSugAsJuSxM+d3jDogUJWn0w0w21VIWzQwfNgHgBtLlOEAnn/N7vIUlpRa/zC9gcjdYEBx0v
BQe6/yqYb3gA7qhoxZ+FUrv0zXBTCrT7xal+yj31mCbqr9wqYsRJnZVFGeCj/a4ZY+0jVmz/EN2K
Ih3uTq+1lywp1/yTwDMFRiJPB+KZVVimwhYLuN5DJKkkcRhKXyt9Fd74Nw6WZGvSXavbhlKj4CCH
SG8ANWWv/ttaWkRIqXlduYgSxoiBthha0XhTymkUXzZBwzmrBtwOfSlQsxwUPvMYOiW+b42oqCz/
u9DvWJ6El+SCAlsnBZr1ex+mIqO2lru2jGqQWyM2zmBkwYPGJ+wQgB3wCfQuGfFopPt1SRgZjTsb
GPc+vJnQkjyNNYCr2jcIj3qNrRw6ua5o7sMmwQc+FW7H6EfXpA8Ia22GLgUVuiRk4yVycfR2lGj0
+tyTXIuMptzApdDSloqCxxIhLv9ZVXcCV7FsmEXTdd9QYvwe72fkEWsrbD8S/gq5r/FivgwjGR+f
N1JRjLXeTIk8D2md7hZee+ikEuWYV8uk0bhEbtPN28jPgGDSphWtt3RvLxzDs+XSYVR14brOsSaY
2LGKZix1KGthy0E03cepe7lv5wJqbc87GNKo5M5rKqbsxTxMgliwBFzMSB+DH5sZTauPY6NX7aVt
WEn3qPKYnNtRGHcaQb0fR2T6vq2gklPWOvdGcmCuiKCrLbjLM40VFBWRkUJjMYdzExo4h/3wsJPm
W1L9/KuxhWa0svroYz34MrBbkDTerLr/140JY9NxxHIfeyXFKWcsdsa+qOR/uL0n65JvMBRj9Ayw
fNYJWGeArUylLvg4a2o6hEcKaNiqhJ8NHcMeOfyyWQAykCBjZ7gcrDCCIghvoUnAEA1GCR9eb38m
0rwpyRTNBDGX/Qymiev9Y69jFFt3pb1nave02xNmI80utM4bxD5DccfmLVSciLtGI4LXMbEg/THh
qtWLj+PeGZ8cuMbQzL6r8MoERRbQYJiDE2pJ01Qt0ZxZCwypA1As6Je35M4LASrnGoPG8vf0orBN
ITkGbmBd3hQcvGh+B6hDXOAewEjSu6Z5IV8tGrG1oU8UebtAT/bQMsJgYdZp3LcdD/jpvz7hzndA
DebMUeeV4hAvV6Oq2zIUgcBJf+BS+JAbOTDF12c1R90UJS6mKdLWyRNA+xGKHyU0ZuPYKWAd0sba
25IVTvyxTNmJq4lm6ILfGQpW+xRrR0may0xYq+UQLsaGtVvhurnpRrcCCH1O7Wj4waN8ZdMqkoH2
w6nJaeEDwtIyNlycruDrF6bIDk87SFDw1Yd/Ryitx0qy2MRaqJWEm2E4R9as/qJtVoE+d9X4I+W4
bVrgu2jjCe8KadMxBPlUrNoD7CIVoeShy4kuQTS9rCuDy4zzXC1B/iIjHHBUm7ESedrqUZpP7VMa
iMey2f21GIQ4Mp1OX6pjltBOwYr+arLPsOZkwwSWkcMYpFwAcHSNA8T3l3IKhQMl38quo1K/O36l
jwv+powT8LP5tc9lweopxJXwCFvmzyNR35TSHR9gjm+REdAyPIYfhktoWarhK4uirMK1Hnus4CaD
10XrDI4cnHWq50wQM6FgO+rL2ScmuXOSunrs3GnKBcjKIxuKaeIRQvHoNV+aojZsoRpjRcCRK9rS
y1z+m5Puls7/rlIeMyYUeupviEyA/xCoA9Mmc1rcqTtZ1nlKd4VeufkMuLWGppThZo0iGkWifSB+
d+6qfmTbXlc5Rj0BB313Kuz8ptWDMNlKDRT7SkfkagXqjsFfOGDXvJeK6QluqecaZHZzCRoYRaxU
rTFdNSZM3I6ncLd4EizKQCvMDdavxN9Zj7k/HEdw8Z7DTbBnWdcweFM6y6MIaJp6J/B0RUaGmpAb
4LnmbZm4ujHBZqKQHp4UGac1g/nGlMF6M8hz7gqttAoCkBzYqNVBwa9ekPY46H2mneTHxTayhQQ5
2h5Vtf1rakERv785UC91J1GQrxc+GFFfeveneeTHI9ktPmMuWYU28yBVMXJz9wmSDjRq6al6B4dX
VpOAz77gmbfS4RH2G+PMwig21guBesBBcxLcaul0lF+Fjzwhd4bZAEP7hjqtXFKQ6oGLfC+OQrnz
sJDMNl8oCYUNjGYp2+ZcgfD4bmnEq0ZUGjLQRAEgPVusiQz1+auRY/UTDBuVE//RcJjEztdZCtWm
EzjvBDs3NRi2ft6PAoYA+aaB58H/gWwdALNEdt4CYHFFhHqYIMqs+so8TkheS4jjfV1Mw+YCxjeq
P+mKQ2Rg2Y0wboxqV3uCIfMIJlPm4EG2Oxm/17/Hq9brZl7fWrExcwoCMw6HT1EgzG2GAge3OaCh
KoxYJikHw9fuDgSi/v/vqjh6tqa98LNNyJb0KMOUlOyM8WgGDb+GuXPDCNanGQb3Fndiijmp+Xp4
1/RBj9WwBFT2iwYrjdcu2y7cVza1zm76gqnh3zH+gI/Se6Fz6vo3vVkTds1ZvKRmM30YSAXlB/qL
RtxmIfyCLJ9TCOJpF+VfuIDRHec+nJibtRGh7gVWIjx5EiZHTkHTFh4uqGuFxdyI1Y4l1TS3r8Ls
frWwuqTqzoDCYds4gNOOh18YWymKO3znuAoWUe6hQ7an9Y8vLg1PWu4mYQuyBI/SF/gR5B5KzJlz
3i3Nrm/EGX6yKiGq/cYrPGnb7CHR18PePqiAb8XshN6JFKm55/SfBPSIugbdRmL6cfjBRtM1v7e0
mCdSUcIyB0ZQbnPr63DG64fSUZ5qYAl0ktFI9FUedlPkpusG90fheTmRPkw+IuAhlBu++EZizteY
IVazgT68MY7/KXUvsw/oRu4AmJs/jg7TEOlLvdJoSLQoUvnZlbFHs5olx7Hc8XnbwFPD+/7v2lNB
pyeMRcicosJKUdDhWQwPt03ZNDXYBtwIXw9hJuRqA+RMbmO+Ja1BSK0URsQvrhtt8WNeMNERAT8d
s0ccEV3M5gjjgXFfVNCHvtb0a9KaPZKugOwLpu254q+itfR+BfPF0wEhnq9Z4RLWRYs7BARW4QDx
Q6kTBpdxkQUAxAyOsV/VEWQdzyM3P43aWS+BvT76D6q8q0Dx8cg+DTy5Y5GrX/F+dx62QiN9u7qc
gSNFkBHaap5t0lQCA0J+HunCkgxw2q2FOc2YfFrweYwe2m+ho7G4Ms9Mu6uMQSK5PXKZ2hGu0J0j
wHOCwvugSBvqm1K0CAQuGi7pw9sb3xWAks4aERIhGQ4Hv5LWVGWhuj+vRduaavoIIG4GFcsteP9i
1+i8kT/I/gkAt3yjp2SxGa0umgcFVLser+J4BTvBUbhzAtc2kf4BMS2IHRdZ7sz39hycuFYaG5sA
J+IpKW+84B6Nt7ZVJycylJ1jz5mxqwJ+mAcDgyZkb7PTUuioW3/t3o+6Luui2i1/D+RqrQThJQrz
FyanBMew+Al5KAhg9HHZBMY4XuOAukzV0+g9kbWiibYCoydx9l57BUu8pUb59TUxzxlVvA9/x9yc
Ta7s0QZ3i9Q468+t1XtmS8KiGhJpwV2IvTXbzJIwXrjJVIrt976Htb3q26CbVlZoiyhzpizjiAUg
z7B/awk0rUjpzblFkskGnqQ2DGGR8k3FQNgyIi1xkilBHyReerpA9xK1HIOlrZSuhSiWNinOPpmS
FZ3E13PoUJVykNuAm5cJKqPDWOcrrj4z5wZjZNc5o/wbDVZ0KIu9n2xxr4iVDXb3Zvpqzr8t4Iwf
P/V6FbcgACwT7ukoepexERe9+sEKnHbi0kxqt3SKz6Oco6V4tn69uGFpq7rzspE2c6uSVkoI2otS
anGNrlEky4QbTshObqaz/c+ZapRrqZdUdsmqOYYkQxP052mzNoQBM7zSwK3/rn+oq/2qNSibhyes
zXpXB9xm1zoMLy1IpdpCnuHc5b237NUBSd+W8QM3jr+fJLK5KdFPwRctYrYVHfrFjkfotoB8d5gb
ra1RyYKYjvsFvOeP/QG6SEOqV1/BAE7JLNoXi7jQFoPD9OYi7aoLMVSzjSuViEe6uqyyRIKDEixk
Ynm6THd8Ur7/CIW+VEzgwKs0q6hG8Y097re1y+iDLj9rbcemb8QtEwiR5m1vqgzaUmHJjcPZNozn
nLp5UEWTx53EicZ/lZ9K0MnrzLMPBVSL5OAh6vPgoqUeL4d/kiryBpCG4HVedV7yFRz1BFLj4lK1
6w7sO9wX+RgxBzFHeEfeNtNdo0FvWPPAbsZGPEF5hVkkD4pWgfZDBKpFFiHVAvAcRsCPZoV3t9UW
QjKgguVA0+CUU4DvWAiAMJrw3nUsmyQSy30eIOE12ev+ecdrc0+kNN+eN75AOgGejtVbWKTrFU47
dqBVMRs5sR70qgxwWwjUo3RF57QtrutLlYJgzAidOlcfGcVKoRpnoC5lbgrqr5bK0FCSXbr2Jt49
BxEMCFFj9IDMyk4k6fKhlBCoSzSeelGlLKinVG0wY2gK4tsKhcS0IZyFAVbxlcahd9Qbkum9Z3Ly
K7+nx3AuxVxLW2N5MEHao0/IpsaOobwUmREX/SXvAZkL2r/WU4VygXyO+/o1JFEOT38FAlvq5r5C
rUKl6cs19PL40UDgh26NERaS8+C9104CAag0cfC0h2d846bS5iw1EHdyrwujAXw62LYiRYZhj3Gg
voz5MV+fxTdrb33ihG+JyW/NmjQGlfh+IIsci0yWhXnlPQDZJxXe0mE0v74lR8puAMCDOuT/fEem
23DAB1g4MDm46dsMdfTzFH515yVR9YXIhqpBMHKpKjBsDwSGKqjuBnKboy27mjzKGvYlNvWskb3U
WYgGk4s57FJP3P6QhCCnRIheF32OvY+VgrH2ASr6GhdoGQUB2u8W8asPI5Gpmi0d8orVg2ibLBRa
yeE0i4XIYzq09ALsb3m9FJeC8/KJur5LfnVAYBVCLghWWcFdfIZL+1iBdRXgbaU3XYxyr44L+TX5
OM33ypLLm7CzoOJ7rGhXg27zPLsajdOHupGIcRdlT+8GD9Kf+zJ3LYQyPXsW9Vd3Vuj82Ur58JXG
aU1/e4RiJ+H/Sg0iB8fs1j7gREXumMML96SpvGTZktlUoxZSWER9GjphBxRIdeJEafATfbLXlxVe
r87Bp07Twao1KpFFnGXIODHUzKks0VksIQW6ehCFYBM9cgUhkxwJa8hGGRBoNLtHqlc87QTWhYfT
AQCC2mUfEF7o0XZt9KnPPlVzt8ZHiiLagQdfP2bnmW9lFl1XNajGpkEdYHGPaazMElYGVbvPqquT
BXY9kYQZ8w43xei+0vFl+KTl46OhQeUfROts7GjLfwxuoNEVqK2BMqLsZAeOFsrFslOxpeXsun3S
Tb8o8SDfclVw3Fhomm7y+axyLNbp+IL2/5q1lXxXo/l50Qyg5TYmwzZWnbH7TZw7HlR1NGXkDpa4
msfq2A7aGK9iKnunryZgtAXMItjdPAiVT4mqzAtz3fk8+a0dpYmVrQN/NvwoPDZ1A5WWhHjbWQ0a
m6ZM1KMK3yPAWxrW/cTY9+r7bZEh+biv3tGQ3AK+K27RXkYeMlkMl6OE8QK9Mya3doNpRrNlwjIW
o2SP+RpkCMqKVtEcic4aGn51J0UrFMfJ3+Pso9U+P1Krt2MfyBBvuri4QlGx7dmuYUrs5lfcxhyX
aM8phvTRPyb0xPWYoU1RynixXjnE+THsE3bGG0u62Hdvj7cMsA2XH36NIvyL6vgOhWaue4sXo1nH
hlV5MMcVnVSVUVOD/8CiGuRDwr7rAd8bbOfvuzBRomaU9SJOIkCMIPMi5+W5KOF81GsQDvoESicS
zIpbfd2gl9YM+JopPONydvGqKs80CQ3qETXmPP8f5x/aKd8DRw/TDEQIUF/FRBu+cmorTigOfn9B
4UP5s83KWsHYctQdnSsWEQzeUlbwSiY2fq5Q0owy7niKPgSnxtaN7dDYMLhDYBIqLMfQGzPd7zwe
x0lOFN9YlAwH66pZod/YofvfU2UYFO5z6KXDOQ7s3NtLg5pHKT09AZSifoLnZh52QXZxTWmL2+Ot
H15wo0r0Jb+Xi2E+XJ/tMlQSWuRrX5rQRnuMKIRRoA3q5vUkOCA3g1mjj2EFhwRK8rCsFdf01a60
4aB6CgNPrC+aMzmbOVlguDM/dA+aqSAn3ibEMo5rD3B1Fenj8Ae3hHr60vXDLbyTHQH/mG2csHnp
qViEteBwECy9EIrLWrgFbMcv/igtCMPu72i7DPi7+SfNtVCMBL9zYl05TPYUpYGQiMBoaZZVPWNO
vM5lH9PvC73Vt3E6SNawD5o+E+diuqLMWi19FT0OLL6/iF1zZ0vJWbl8uvryLvygchzEm6Inid5k
bfvM0WTrBOzQ6dLzz8yvTrippIK8hM1K3WUEvwo1cMQLAl12wgP64mOYTGd/5nqRZPtBJHttA8qW
uM3ENclzAIraN6PrjyrNT4BcpNDg8dxYES17n+aiGd5lhYwb/PczY6FQffwlLzLh2yVbl0PAVqaa
VaTCJtVpPvn4V2iLGvmcuPC3t1BaCGfBYDqaZ3C/ePRjB5ac2EYd1+UgSQlFyZvw7X4WCR9bEVKz
ia7M+ku60MXrSJvURB0N6bm1oYfO68ugrZsOzuNEG1KezG0FZxc2hMqCMnCo/a2LU84pYUDM9U/M
wk4TBbL8/j3NPVa6hoiNuhxqX3zwaUWFJFSbE9WfBkS3w0UsbZFQQBvETpk09OZuLiR7BpkSx3B+
jv4OgbA7DO8oCHSpJyX3aXYK3BmEHMzLvqaXSTCjzhHW2SDpTEQxf3lVlgJvLln4z0HQ18Al5OTJ
iujk1Gbp8fQihBltN6Qcc23uyKtP8X4wUx/gWLFId8WWHYDNDkRKqut310ThPmL6vmvKDlQqVGXW
iv4MxNaLrw+zRcNWtcPIam89fss3gHEJJ7nNI9zmm6wTIhQZ2mZGWfiKWEr8xu41hOvfvbSqgMHb
eAo3FdHxcY6HieK1ATJW8RksMOU0LbZGDwSqnexb5o5LjYXgjBUZJsoF/G/r7OeJCqdaBCeGE0gZ
T/h4G3OU3UNIxGbya5NLUJxnQ+3ZrA8pL16MrwfOeW5L6bnvoXpm/MeRaBVuMW8U7NlE0cwQVcQ7
wBs1oQMTG+Xzs275p/ul0v83FH/tvd3wlPzKp0ItJYleLI97Jl1B8rXbmgUgZHGCaWGoKyk6pS1D
d6b+eDGMqbxcZGD4J6N1WlP5RVpbDsI0oN+AdMMOpvhJ8VSsljnEuoYdBQyVaT7yowDxCYRZQ0Kg
SVf2U3uWM44LcjXVCrQ3iJEj3nqwkg9Ddr0go/05IdgDUGVZvaiECzz6Ksi7zxQ1WhlbuE2zn2d4
W+a+gVof6UtLoBXl/gQ4evTZGjIovspmgK9SRe7drrWLZQwPCZgC4TjFXgX93jCBKSNzrB1iOv3k
VA9HkDL3qCYUDltQf/Xgstco1AmuwFbHt/PeT+kiiyehfjx2WkikU2tNSQ2aTipyiX0eYE2JL7l0
BHYm8bxVi4Tbtbd3edqqXHyFm+mXV1HLcU0J00ltJtsWf0o0SgJIyiZS8trH5k/g70sJe4Z5WReX
vNr9AV/lY0v7T1xzRInqUWLeySPQ/yx8HTHtDPXClVplnnZxc6k/xB2kd7HJtNsfs+lhy4slqqFZ
WpPbP4ORXB/jGZFVF3w2DgKDmwFRe+uL3KUzEeSxiANIe+mU5QQglWuDFsp9+Jla4pg6sKguYJLt
b8vb7+iqY3YCnHFLu8jw/oAHnzHIPb2IkfvlExQ/RP0sFnJnHnE3lsmvfV1PQOuXHbeqO/35wGeX
07Rb2cM3QEc53oPXzCyCudedxxo8V1c3PK+NPGPlgO6O8snpedhca/pYGEpyPEC6ebrYi7Ktcq0Q
CDsPiJkr5kB9ozpPw7YFNl3tOTSkZPJoFP5Rx+Em2p/kTvq1bDOrUZXcL1x4ABl+Oza/BTAlmrLj
qcy5bx31G/mMSZ5pEPnbiaPddRH70Bu0Xhc+vom5yadRM5pjsPzsRfGN8odcDQwp9kzBWnYXCT8V
tidCucxGx/veCmBbRM2PNk7U+DxBwVospJJq3fz/05peTm5hLX9lmbgpdLAVkfFdsJfanVnhR3h7
y/TgYYTARJVgaFmr6qvVJBWefuzagYOV+ePqhgFz8OhjhOlgjv8MFpNjtLjvzwRvOrXRgfKaO/rF
Xbbkms5jIf16dN6rYI9Eqo5xXdSSk5neBWu5SAdiLqx5QCxdJkK6AvxogHvn5Li6LKDnWFR1gmK8
BV4yGyzMUtRNuoVAB6u5DU8EO+SXrQHOrpdWQOCe22oyhk1Qsilabflbu1sU9p3GfdkcNtSpNvH0
8wcJXiY5eS4XqxXaYiwQjR912El66Y30SI3s/gNTviYqxioa4gsJiwj3RY6+gAYL9k9A1ERv8K0z
qfwcmp5bSJCvjlPC81Zezlx6rfyPcl8VFd647RyTQvWOJiLZqzvcBOS3VM7MDiE4mphA8cFIDa9f
SP/cGlV99rY0YAY+RYV6UIiKT0ggyrr3oPvlqZ8bTinzjYUulYbW+js9rgJKFyL/OUBN7J++K4iG
vgZaH2m70fsUc5jby7VCqq51oafIE1ugz7Dbjrf9j5XnsLa2H894smxQeNpfvTo58g7/BMM3/jqG
RV6dMor7vTjth3s4SbYBPLbkkTiYRr5pk+Mb9MHFu7uPYBhysfuJcECxujhlbycARekS5lnfHiXH
5helt5Y3kc7fdhblDrCYFbsMLFqlgFOUwrRieLJhCzkYmWP9QIXsw74zQWlT0vNhyQ5f5Xxaz5Tf
7Hun/sgcPzhkd3d+KRtzmoIvnrG6vl0erLVRtta4puTan4o6+HIXuY/+sO1v9dlGmp5ubU4jwJUY
tJipky8VkI7EZ+KJR8k/fO96iM09RvaBz3vKXxx8RazChYiKCVICc8QxDkpEIz34kpzaH0tl3ifX
UVdlPGAxieXdYd1fzVLjwCIGOW3CnBYvVX6buAYL84LMrOS8XG5RIKTeOPlZycKjE9gXnqjRARqw
AJmAp9NyYdE4qL/KBvymuC6LbzK3esDQesR7ZTTdtUHArMP9BdyzJrV2ntGapvhKAD04ogINtMVP
F4QF0h9JcMMp1oVjVIp9be5CSePUNYo2YKCOAHwbBkW2NYHxmvil7PCZFDFUisRIStXbU7Gnesj/
TthOy873j5qe8Nvodgs5HaCwAv12kPyhL2g9pg3ZmCl7sZT4YgpVJ0m6tGDw3fTTiTq4p2NfEEQb
GVg5Qrh2eNVscaZOSvkpbNe0TdcgK0uJ/eKawkXTMeBh3ueNrhp7fZUwRkz2sZarvnkpj86PeNo+
hothaDVDsj+WKq9xZE+12WlnVZZdG8sAiNy6dEV8MhTB59YzdOOBA1YPZm8f+1nt1MV19NzyOGJH
nTfyR6ZlP/nqP7M9ysjcxKhmc3YQ/jukBrB9ZwJBEKmB6UtV34w88NX7qZlv7cDm280Yd7n7BCxn
w9wxjrAMnHM94+Yxic9hlfNvErWUAJQDn3R8M3QcJxyCyzwUeBgfRdK+4V8IcWOyCo3PcWIUAiQI
c6G9e+evhpkA9+i8QWRZqAZRtjgUaCzrONT9XVxZIjZWE+wBDZx+yidZGk0pWkrIMA9uvq64UNaS
ShmHbFymFKrER7x1SrCoIz2iDf1YDQWnVT9vYA/F8qkYBdg8ApplNE6fJkSHmikDJRJiUZde0OsP
E4/JdzqeWrcGsDtksHQYYlOhZefIwJmqijh766+ONoMVVHTXrHCZ2o00UIMfBcuk8TXhpJtC/jGe
r3Ixk61h8vGUax5QGIb08e1lNV5j9l0ehMTLW8XoYVkhz9WZFIMGK4cdBkdMfU+NcTG5P41uzCkY
xLLbu7Lvt+DQEgH+doAc/u+62MYj4tTYAu0gJFWEAwbbNLiWg9GVAUtlJ+qsqI5wE/48Fy51fhhP
haEOKJb5SwlXJhankiAxPVTUt7HMZT/24H7wZItqep4b7o9Ybr+K631QW7GrFCZ8EQ0UqYymtDjk
p7fLbjsPuVokMvutCS7Wjb2qXrvH5SajZmc4bEfHKc+teaiEfI3LWULQNtPG4SIWyMosDaLnlzzF
cwEpOtOp7I+XG1Q/EvhCfZnXv2FF21J4gK3g8wbVvt0tC9xzEGEwc2HEprpPghxk88+nS+FSMBxE
ti418U2m7t09CVIy+LcAnfWM8dCOYmqxpw8MpNIrwBLUq5vr3xqT/9hdb68Zx2yRz3hVKjmNEvSk
0C95duQptR1IJkdcUsZX/Xe6yBFTc1itIyKcFYx/jkUsi9RDT3xwO4r/ouzrfmNSAV4aw8apjTok
ii4Aee7BG4iSmwZY1ucn6Oiv+ZCWRBSK/9AsSUWX3dXaYgwJnOG1x3ieK1Lff1XCLfX7qKESzvHu
WIfjJNuRDTLD2+rv6foiAIXwze7MVu3mMs35jrh5blQJ7liEB71sRntm2/ZVsAgxWGoWvKQUV+EM
p31Hqr8j2F14npmpT+8i1DDXFMF3NG+YDEF7Q++rA5UgUb5sVDEMbEDvdyjZYzwQM2re335CO1Mp
c5g9RrW+R6VQD2KpKKhucuIoDU7/az4Yfg2GV4wppomTNYzs0rd+5UhYxdzG7sWDL7W8PkTTULFE
wC22/zBjpkSbUjFXHm4EvhKQiupCRkrh1C4R0XuKvWanmrX6HcqsCoWwZRI4BbzLsARQcUbGkZf/
2b06biL3PrzheHw2CmJd52yulxEAqWWvU7bzTlteFmaCjhXDg2LTajWTV5PL3OzD3e7h3N9WbEcD
FgafSL1kx+r5M6CeSSL2LOwTwcrtm0BBf7x1b8Mwd6aC9iQ9bfNO09pvnmqLpVDumQ8BBMecXFrX
GcsC60kDowPrD7I84UMQyuansWoIoj7mZI16qEBiJcxhBDZn2JbSJce21SKLF1GTCoSaMzO4fbsU
MxhMLAYQrzSF7XWu4doClei8A3HaspxCzHy8xRUBEQ95HSp62lqLcieFhvNtq0a2YoQ7usE9YClP
B9DaTgfbm/byCopKtWTAiN7Hv5kfaj7zvNx4Gr6ZvQ9FuxHCzHVVY+I/tx2KrpAlxl+TaNQb4A1v
scu/OfV+fwcIKcSQ9AqBpREE6Id8o0Pdlk3t+pLeNNxLYNmcnteCFclTiTdvJy/s7Riuu8anQtvg
Q6DMHzUqLaWj9RIC5XxCFM97QGyX4V0m+doq5P5lPG33ld4Qm0QCSHinyaqLdgEN/NjrY9Ush3J8
FxSynJpR9DfIKpe9VHzT9BSMRGBLlttvIgsXs4ORNU6UgGbd1cTe11M0LlvRagiM8veh3RukRgnM
K5p3lYe96iNS+UvfrLP88TfxAIOTyS+Clodrbykxj5YfE3nnIz+sCgxN99O7ttyYKy2W0pxkpNLM
wAHbt1eBzE8+40K+Wy8SNEeSJm7/wokSIE0aaInJGlsEvPkcN94/PAgAtl4bWfzQc+AYfmLXNMFh
w3Q4bG4efkqFw/wvSVFhLs0XNTfKdMNiIdi4D3CPCd51QqM+FL4GDM88kdHumzVYX4KxcyS9BmaP
pwh3nhdbkzCvVK4cxmiqf/rkUrgbbgP0ulhSuyrDAs/x8cniClMARhj8okMjWHyd6EPfRTx4U3NO
XD9Ylr7exAlw7pmCYCGxFRdLtzATgfXn7H3qnmKKL6Zn1T/IFAvsOzuaIovFOgZPj7KgowW0+ak1
4bvO7LC4cYznxDbeLIB4vK91AdpENlnEt6tvy/DmLlFACni3TYCPiYHQVpSLjsJGoDpMeh1R3Wmy
jIbQwWi9/ZhTWZSAWHbBs1RYPTuONE0cBUquYuzIIstDzKpV711YdpuGV3KwoBCuQ7z+a0mmi1xD
9XMdL9r6Nq5aq4uCkPdlQw4FQ1fIJs/O4NMPPP6wSwVP6+vQiFbUDB0yMBfgf3cS95pswmMvIp6K
FLBB+VKSHr5TpNbi0Gl/NSHxsnwzE3/TL2J6yaERi51pOQ5CaV2pnSWkiOj3jSjftvYF1HAEW51m
7aOwj0OBUSywDKb0g+/Tsg/H43G4aSbbKSgyDd34OWOBHzwOTsUjxOpWKeC7WEdHyTci/SktLGiI
0Fx8Wyb7NRr+w7Tmgr1H0Gq3UzdYipQ0NZY16KQ51qPky4LwPmNTQAYjFjkb+pUHxcfJQ7ki15Fw
laKsTQ66t89x/yotkcFXTGV/Jn30GCCWSgxntXPCp+5p9JtCYQ3wEDyr9nCiQSzrwzychtdB5UoV
LGADFMkC6i7qgWYoJgCxvI4OFwb/tjULROZPluF3ac0DJJ9/qWl/H8lg16J1Y7VoFdjcpANlcc37
D5jMPzuVqz6fvXld0Pnov8Y43gjoYephXHDHvtck1dcnT8oSt/V4wQ/NYcF/MY9x1+Nwb5hGQDRG
Jlw6mo01hxkhWnJFHVDJGFK0co1bJSy22br2L43WFYE3hmCx5DMK4cBcLst3l+kzJ4mWKWbfcnHf
xjZmfMlNXetEhL1LDvqVCbE6KiFH6PRkkjB5y+iwxNlhmTm5kj96l1hwDSGKMd1dj/nyOI95kBab
fOOpPz3SKmjEI3P2pxKvQ65QZ72n6a/nyCBy29tHc592ovhydhduAlI2uP7MmhLwOa002H8Eo3UG
2Du2cGmbuQ6oiHgAZcS8YCZzZGAzOtUab/6/hIbokGaccwRhHAYODvW5gje4AhmKcG+2Bg9zHv2J
po56BgjpdEpt43FWCf1RT0ChE9soWpkpBEMTEHwBwjeieupsU7GhRK2BrbG3yvB2rRUORSESa+PM
kLeox3dRvdU3dPdpC42hM2gI7U248igpozI7oWjqcQz7o4SeuDuxn0oBxINCL1RNo7sRHOA0f0in
p0afeG6m9YGaoW/yIM5InSaKbVtNmk/bqZboajrcexBjvo3ZfNoIJoMwtnU/r9JZqMNV0Phc4gGl
NqTEOaKPfloQUg3ZfvCkhVNb3cFcdjAWvj6QaM5zq3JT+UkfnfS+B4l9HbMOJmYsMAp2QxGr1jh8
MF/e+LffxoC/Qt3Nk+8ghAXhHhMgR+y9GxjeK7X2zW519nsAgUEUVlx9GJSy6Mk62l3mMTP5yaoV
5K0uxtiUhPZnfNXxLP3vGA1k1grHJm3RUcnsMhnf9Vz74xGo2/mcliie92qMwTQAhpmSU+9Hu4cL
ooTpkY+xUASF6WI2dd5Mm+vk+7S9ca8TMuKEgEk9mAqu9DhZvPi62aDm0vYJrfR8ixIo6iHDx4vs
U2OITsPwApo/m/cxWeDs02R579FnsJMpT1EMrBArDrcWqBzJ3kZpVhzun04ddwDcIQUTBlR40NpO
katerd+TDERfiDegVki5ZGE4wCePLOvMClYbKUnvVMcbfMPmZfqHLWDsduVSye20Wi/NgQBLqkNr
ITam+ujiAVm5BCXthrexmVtC16if3K3BjrG9/cSB1ZWuFs4ovzwmh1AoMjfdD2Rp8iAkksPCKdpT
k5NrREI2pVnIhsAJl0FP3VUt3+ir45+j6nmUz84TGZYZSSyFyHh5HxrWOwDvrisRLESR3LtRif0J
dngbgtm2Ob9h1moa//7RDox96zwooW53pxcAJjiNewxy3qngxvXaufkS1BBbcZwT916jBhOTLAYE
mglerzvn5jIeuXe9rKWkWhHrmt2mj6tHo0UP9urDknXvfKWvCAPladN+VMgkH+VIFGVAnzGeCal3
Kb5BwYOGWTAEi1y0PakPSq0QbbdMEOtzhi8k56S64GsPJNh3rG3fgGvYnvD5hjBwBTnyqQFRny49
KQn4dEDbtA/MLkEpBeSlQBsgZJZ2T/FSz364SvhpSxxMDIlVIdu+3Y4KS+SbOgKp8qztYRJrFRsM
o1tbBqWvJsVlncIFlDKmvjvMLWEV1gagztbT7BqoPdJvHcBpJt2DaJssR3lwKsFCgeNCq0s8HWIH
F5F8zB82sXG5CIAol70Zg8Xrm2wExHe7IQ9oiErHmLR9KhvB9zdQnCInGVZlTvqINPCIS+imeUHM
RaUsmsZBi1FbRBZePsYEdXlqZ1OIV6/kXCZKvytXGiYLouNR3zsnwujLuuO6ySS5yJaudzksoH7q
7CAl8b/G/74JIKVXGCCBYUjvWgBPZN9p2ZaA+JR4hlxvnOBriaNSKQ+QIqFgknCQ5vP44QHS8rXl
VEbF2crKtVpZnjsTmkskGLkKBR0F0pJ53SKQLGOE50QqThvgkjQOIRpPJH8qKfaMycb6vsnTth74
2jpHI4IvbqvojY59af5gKN0DlqLIX2Ar0Jw00GB5uoCnIygzB/6msOMd2CNHvqb1kL4txXK3K0PH
e7sl2XIQ16KutrPUl9hMV0JjEbkzoRkZisSAgg8/f0p/zy32qC8sPpPeevrOqsnAqsqllO0FjBzL
vLado+VSMyjD2wDUp33IgGWeb7RbA0pzdYgmRgL5lNG/ozMBx6qiwHBO34ciQqSFoJPkcM2S4/sA
I4e+X9IPoCe+MevgziidxIidWuRZN1XBotlVvHdfIl0nscW/1TCkkuQb/YWl2igijV7kH4eM7Ls8
1/dwTgKFJmqWTM0CUF4Cl4i3EJwdVlbsQ549yr9BWlqHOvsGsUkeUYZ3TzemZeFKg16CUjBrw0LC
w7F5EyjCChTScZ8fA6G4SbZ6gj8iUrnCC91zTri+jtCXVo4GBAPtBn+qP8/JhMEtN48kiT8QumZv
9TkoFWO+l/4pom5vyKi39O3iGW/5unggLKWUonvyD1TfN7PM2fb6Wuk/Pom4BkKyND96vskJ7aU8
9VtLjeUeJnwG9mF+XiaVI6SIQFGyHYDSWmSsyrisy6izu3k4hc0hnjMX2vrEb3SgEq/rnb9HTa6p
4pB4VqdMYnqyfodYgXvLhUHuhHuQOPfA734+abGllWpGEba7xktq9jC3A4MCvbm+K5g+WKrd3U5O
bNjgjGABI0s62kKHkF7hqdfxJHN6BielWrRQSYiumFX5omojA5daxnKfgZC0XpvGk82UJbtflVyQ
4wqahgwpqF0oApCsF+2jUbIX+gfTyXXVVa7OSXfea0I5uVKluOpvsm8ybhjvR/fa7Ly3VU6i/WgZ
neGkAYsrKwBTljwDmQzbfZf4CmOtKgAtCPl+4IuNFq+IVa/fDVL1H/zVicOcaHZz9tMK753uK+uM
gyOlNTJo4L4e6eku0zTfdfAgaylUmSAcP08e4xi6vwr6XeWVHmDXKuiu5QccbsYRQwyPQ+MRQXII
m73wRY+TpxdCqneUljKiq1uEZ4sD8lykhr+V4QYwFz9f5gprIkhloT7JxT0YfLhpG6SwGK+OCOdC
Fa6MNL/4bVt11OZlcRIGfBA/vM7c59lbOfBAk8gTPtv4mJFE+1V7mIPFRxhj4cdkGWMh4SFA/pKe
au4pROptc5uizExg/lPzoE0eDqXn4t/ReU2BzO/0/8oQ+khUL/1NdnMotaNyUaSo/WJmvpHVHhQ6
68e0oYsEXhsoWYc1aYQa7l4tu50UKdWwJHFctNq3L5qUMdpwFjb50jXYk1pF4T9jOxgafbliqfUb
6hSEL3LvOK977oYpehPO8/IV3HKlKgDNd1KWlnjhDlKWfymIjq/NLC4oZjre+PVyAkeg5sATNB9e
AHo17hYDCp6Exgx7/NVGZpuCOEeLq+knwT9M027D8MBZfwDr1D+xp/V0XRHFucGnV8Mgh54ASKgC
piitD8vGQmuE1mH58Tclw1bMgTEnDnZ0CVT9Qc24pZpkzwnoGbJLrEfyyVTozgPHty/XxF6Bva1Y
oPHBMZSZU+nfniGk6AtfWF7XQh/Sq7Ue9zFq2qzPkxO7s+t2990bshp1yzJWRO6AjwlqXyGN2FXb
LOXJyPuN5qj7jDv+RcJrqWn2E0cpEd7IuBR/BG3Pk7xugrpklJ/Kj8T8ga5+MI1DUaWKKNvAb+DD
NN1lHXE6it/L051ElgrBpcZuxfSgV7ruBMtBU8oAuhTWEMnFHsoymwsnc3sxQ11bsCOaHfJABuvQ
5T2J3N/wpe5jW7ei8hwvDB1yQFGlZkHX2jddcGqcu0LSDErb9/I+1RuSgkJvYJTyD3Kr1bQbG4Zh
KuMM+kAWme9T0VAUoBzEKfhX0p+sv1umcU8r/YFEO9EiYec0RFRRJDTuDlX1LOfCR3y96HitptGg
RXtgvKZFLoTmRJ9DAW47yu4sLIMhjaPGzskXszeClfhWF/y7tKuNR92sHzMnEhve5Cn8aBXANso5
0xwR/Zr/npa4UtTcp4BgJGnqUT4dZa2w/GVhrcRxaDhfd2jpy1Q3fdOiVBDAuV4ga5Err5i5ClJC
JNb4ibXxiQZH+fo21ZEif3prNX4a6q3HwO5AOywgE68UxBrVMpYSdcL+QA85c+XvpMGivqk2PzTh
orIop8zod0n9vdL8EuKAK5rXbmPAUvVcZFCPcisiCwSeuYDqqnM10XallBEtQ6AH+I49blKXhl0N
GRKudqKcdngWOUOEYWawprr/33C/ZVy8CBo4Dqlxrv+zQZYQwvzLYsv8YeNBjIKXElArn0PLOIJC
3JCbxcEJAO1GW5JCc7amx42keGRt2OgD1fkNiZ1niW9oqAqptKsWJOwk0hsl3IwyLEo7Q6woKU+D
CHWvSSKn6bXDYO4N4ntPFnqJbrC29quhavReo2xvBNUBmFe/z0XRfollj9vuXtHyRKSYYUETzVqX
3GOTFd4uS0PusBtl4HN6Ea65YP8+U738/Smg0hefa4S8LmseYpBhYuFi3O+HIxWqBbChLyycBj59
sDMqsRnAc6kX6t010NyqPiOIvdBiyiRSgeFKhSb58cl0GV4Lry+UfNxaacrV24DawsDTHB+E+B3Q
zOCW+ZmKYm5ZDraJCqyEEOKAwkXP2xlFWIOJrpEEN1fxaGBtbk1ntX9KVx610m3Q92Gi/SQQJq8k
k7ytBC1ceyvlEOSsIpDcX++3PK6j4yhlLTeublfl9EglfvRleYRaK3GrhQ6MLFokh43zXCNQXF8U
kVPQeG618A9EtvAwQoj0aNCIZS4lNfDkQGboX0JBshJIgWb4Q6PUgnShuAAteQp6+CgTf1LCNpZv
PWHamdjvSH5z6eqCJab2pVayY2J6PbT61NAktLgLfmT0kItUp0vvAnCvQFieW1fzb2b0eZuFv/eA
k8G7sibGDkzfjwH2rAsHeUhD7vBIsmxYDJ4PS1v78Ivie7iRY0Ffs9MottICh9s79y67FxpzASrU
D6ht9BwzTcIekUIQ0Rs33VCJiz7ceQrrcYzVoTSXvWi58y8RNLP+FsVeztCehQAGhqa4QTfGSv2X
cc253IseDvs6R2oD706fRyf2Rp1y4AhBIf9NCwpp+0QPbbzPqlFxilsnwsZPkNJq5L6jtnM6eEz7
SPYvdSXafn8ATCN401FmGovNWmykGTMmeUMyqPwYsesM35X6bxVHA7N1IdXAz579D4xt+2Y9tC+b
6ln5iqEeg8/1BAL6kj7m8a73k2cIIe/dacs/4o47jSdCtLY2N1M+883S/zK1OUm10AmtzrRTn69x
WtxC8heZw9vkztZJHZzKWAeVp2FEnlkmRLnicXGuIOZhd3jWqTuPNHqw3qm3bNAvEp0PY5xaj8po
D3N8/mzGwyv0KGZcOJwJmjLTnWo9ZrtHsCLjN8a5tPpvLba2ilmjEuHpY6UDhRK0vOAihnnMwzg/
z5EFUiW0CMpkivaI7HXIVJCJYvD4vMui2lqda1JhfRhBaOxuwV9xbddhFp0hv0+KEHxAHjmUqZRO
aSBnQHn4bF2IlwDHY9Yo9dJYoP1e3CGrnfpSfnkqfalhjBkzZN0D+zRusK+0UIlEMhVyXliLOREr
K9Q8mEY4I/gYpvIgvONtSqZlrgKry5ycZlrQE+ZUkssX0xAUam2155S5gpgaSK1d1EgcxZ/8Dgy4
tubFFBMG68w1j7VKAvFE/1SzswjE6dDWlyCT3pE+tBDkPYZhdUmY4YEJjYxPuDTOKAT1+f6xXB10
eaV8eyw2KfiFmk6o17AacZQxCfHONx8FXOT5BkV3KdzH57hfCtgKERTb0mntmsjzXDidOInTR56B
go7GTecUJEXsUsUFCn5ZomMLBahwgiXGDWYyN+nYONOtZaNjtgas//pm3QbxMHSTZIMNYV9vXPGv
inWHVCo4IdZzg+ObJjMnBarUPCHv+ob1cF5J45EmvsSp1yT69Io4SR68jqyNTpsWrLhFQ3hvbmhe
ldxzV0acJzGoffmU9lkbDKoO2SnFKzKcd9IbYZoKTaiFQCp5gn6UYRm5Uu7Q0Jc/hxprM79G9wBQ
eLA27LxzcyIQKTKPMY5/gXHEJLqysOeiiLEEVYuU5+f5NAmq4X/llFOEm5agHt1FW3nxh/SMrNV0
YRo6kNwwpJ1Rob3BDB5F33OPTQO42nmvosi2bHs1ZhlRHOX96qqnoCENztr2OrxFo+izT+LKW7J2
SlMwf/p+FpV2Drfl/Dr2Lc0mwcvROkn2YzSIbbxBe3K/DEkUymtHSukQh6LVv0WAxS7wlUM6v+YA
sc7PLlFg8Ewu8HOX7/2MIdbqO3q4izy11Ds6xjnIW0HRbsXoJ/Yyhaj86zF85t/iUSZFrZmQkxps
D5zqpwTkQ52F1Hvgzbx1nTkgb3uuf0MbPdLEhlivL166m+sogbWh/PLkys0ye+2rPhBwfHAVF5fI
dnsSUI1y+tbAdtV0s9xBAfs7+NlSS/+hQXPeVrLXGpplp9HVQ6mNag35YLHK7yL8G5eQlBruVFRh
fplzqx9GTZStNRLytJNcit2+3SgTbLQm2WoYkDENnTgouhrY695fzCj3iir/CxlONYNH8Zszq4zJ
wt+xc9FzmSjNLfTN5I2z/CRaokzoCyvuYlMJ6FI/YJ5dLk4Iw/9M6klvP6bZpwXdSA4FTiPYel8P
F3ywFYOs6aTOWUTIPGkatGQxoFdYegxqkIBLE2vXom9AOAGvkiyvx+n6pscV/7PqVLCAmjp/tYy+
7fuK1PGXPGu7r2W7QhPaCrDiwCnz6S+e7ue4I691y6QuiLm01x1L2Ck0xRUpzT1nBSsh4THNLOX6
Ev8HADKmAEtesOKQICUmGobJtkchOBqDPVeWrescb6h2sVIuePGr61UChkB0buZKxetvlzrgZgmL
/3GgviZLWRcY5vQVMRmYhFXRnnR3g7O8ckA9KVSkWVXq9tUZ6d6Wlk9cf0L//9ZRl9N7i0yt4Y1G
c6u1ENxtH9KrJpJOLzLmTj1HMqk1GSx+cgBHocxSu+PZfMpLwN9bexEN8XpwSf9+GFqSyLlS4XoF
9G1UCsM8TzfuxpQcIcN3mi00jN14cUe+fnsQiitISn/VmtBa4UolpKHAncBXXoAVGjSb7o0UG4Xf
IXB0GEkj18SsXUMp1NvH63Mo6PhyTxCM1rmR9ieqWigoJCOcj1N8ikoL3RMTkxnaqlf4ZKC+FYYC
DYDSxiRhUcmoQ7A1yQwk50b+P5HKzFh5+rgy9DwjC+L4EhhWW0DN8fbzDKj5atEKTd2aR/zUWDrz
yZVtTYk88yZEbKmrwh/cbir0KNuzmegsjsbi/EDfhk8jgmtdojUcRTztCSYaZyje/e1R7rqv1Y9U
g50oWJbBFninMs+7wRrLrPs/FU9TJxv8g7b2zJX7o4NjT85aeLDhHbMSY6BOaaZLZ4iJNxWvrwA2
PLzjzbWNVgATJhJ4dLq2VqyKxPsZp3PO2C6CigI7LLGSqEGWYz6bvpiA0MmCEzYhg7kZ7xz1A9e9
UgGzJ45hrz8oEtTcRkauDjHjGKf0LgM2XHLU9x6wkzwjSPi+qY+7ka+Tn0Rd2BmUrAH2hwWNy3a1
jUITwjU1bYkqr9Vv5XdY6CfVxPj67gzbSEjB5JwBNGCVhrRbyO2ZKXCkwCrH1CJmzpzubjiP9A8S
nAS8Zr9pqpXvy+o30pUfAFwkkzwXYyTQqHQeTg8shjUkD77wld8zfFId+tqzYGpn9br8ZaQjW2Wq
u3ZUOKiD+23p5hcqX/G0Igs2e5PVpUBcfY/6bmaFYWxUm3cn2HPd1eQV0e/gpPriCz/5EItdj2x0
FToRvqrZkoWqRaw61Iy+jam3ljtn7FFYbCIn/5VMzUnJ8RxHljazmYuwsjheBxx9MA3Yllm9FPZI
EqY+X74xNPJdZvbimPO5PpwMx8AsjzmflZbIwVoBEaDGbgMBVvlRSBAed5S5wngil9ClbQZWsqcM
C85OR4nzaglIZwPQq88wshDWlqL+d7ih0af6qifRsxmZ6Y0esKmgSL3UlXlhYDMbwYsKNhViw2cA
HaM9RYxk6h9kOgiPzAh8ZvQ3MrIYam+uGriCFCR9uh/DP6jxquCt3JeuybIumDtLkpIG+EZUj/bH
gL4HjvsJyZVInN7gp1iOKNzTR24LKL0LSFObxRBvYElHg5dsSAowyxANxdJOu/bDTb4fZ8DQoerT
yzvYMGEHP3EbW2ASMbS8kbcN07P/8Ct/2u+1z26uEBymMTf4OvCjZI5kVimLCBogyiatNiLcmegE
6j/p26N0L+2eFRs12uYFvJEm7/MsYRZM7LRctd20Csy1ic8gfZ/SMYU9qaisAqf9gyO5twJJpbgA
6omrcLtF5oCVslwDM0iPAVexLqfY62RlZVhVOScT/2a7cVyTliuYzTtUu7qB3QQqrHceWnyfmk2G
cGD0eXHmXRn8pt/2Rkr31F5RVRtRGQPI2nH2iPD9YXue7IBbeNphOQsUdporGBG7fhCKPJVTGVOu
06uWxvQHCqIoGfvtfW0qWzMXP+zPsuIzWGEEBsWgM80qqM6/bgvFrVlQkfXbr/RQkb6V+It83xyO
kF6V0q05jAJS1itr9eHlsRli8Zf3NouU31G6i4jsjJB0wtKQmmWcovzqSH9Jmje6xAx787iI89D5
Qht656enAGLdPfGmQE0w3seRXmgQW7Sqwc6bCj5IHxOhIWa6T/x8twd7hKYl5g5vzEZyDFqSmsuV
ak5mZgxohXxijEMDsHM8aa6eRNHwm8Fc0hJbAQ1/hhIbFhBnAtNBEbL+1Eztl03nDIY/VSqWRBfY
hlJrboHXebWL1Lgm/YCdsBKetyQNuyRt7gX8XJ9DPOgnjs+aF8FRtYLunQciqHEYfCuM0N6452y2
PdUMVLg4QfYgyBFmxgJfMoZ5PKTTdxaW+J5+atmpGxE1dtf/4LT3B4iaiHmkySOXnE9gCG8MIekc
KLvvhhO+rhOnP6KAT0rKGx/IOI0p8vjRW4zaFv447ac0sVGVKs2zy6lzlJMz9mz5U2oe7mlU8wgx
SbqWukuxt70IjlrnU2ouWZa0+R++g9fI3ZmeWUh1Z5wbbuBrOrTABBvA/10+u0tQEHnjzpTHTwXE
ReTR8BAdwvVW6etZfvDnp+zVbWJiZw676LZegQgspoDiFOmSHWvDZrRddA9Sw/EeBFDNuc5el7Zl
gQOyPtgT0XhgwGreniJDuZdUkHcrd8Sl5zCBlZUrL8qcJhDVPhijAEevYqqX0S47rf8s2H9aP85f
j1QGHSZk3Oglpdevzw79yczDT90VnnM9dnPnnsVKQWK7qSS6FggUe6TxH9aZB+8ofOSPoa7Xh7vg
ihRGAJmtkxSuHihhB1VIhXoEvfOlWDFi1WQLoEB65Bx+HCQmbP0VzS+Wey1MNLhCKXWmkJ05Cyiu
zeHZbT8v18feGU9lF2zT3DFOv960ZW2a7LZxHWl+ORS/wDd6lYkc+MrhvuCsZbEJfYZxI7/h3ZYA
3u0d2vM0wzdTc3Xnz+XzjyG0w7TaYJ8lZzvKxmrBJc0/+Y/hlMsoXfIKzj+N99nLYIE+Tin4VCLA
Pas7diLL2RaRrLzBCsp46oRe30sj0pEw5DGEJYxuozFgxO4Fx1oT9vrVvDhgTaHKd8r7vS1kN964
R97ZMDMwgUe41ISktqXWonRUt74M9Qe4RTNl5n04iEhsugSVpUpvQ7pSicXuEVbA0aGk/4xapnOw
X0OWYdDZR95hRaeKh1ofwmGnM5FpKNLDj8o9kR5fGujK3QWvdfJuxThoqIQUnBibOQY7o9e0gvya
q0gqstDZLHjU9He8CHvcVVaJfjLHpREiTDAKcoJSkfRhA9bzzCYFPgyqvRvVW7H3MTeDGB7CqUdn
u9U1ZUi2lTzDidivpHrGVg+WDIrF1JwU3TB0oFY/AZDhg+ERBW/GgYSXAQ4SWblAOCSYYfkuI3QA
e4yK6OwLoEGOBqLX7gMIzh+jXxwKO2gtflb4a+tQsiJLHFKKf67GQqawp1xsmWLbNzCAB7SMxBgr
4UW94/CkoKX/3wLQfOzsBgTl0YCzN0c4GatLekbAk6Rtddy/QEr7oV18M9VmZNQY9cUpvzhUgwiX
C37cAztYbeEPlbRD5LbsEBP9/2k/ZAn/AKkXI8Dw5X4F/Uzw4YicQiaYxnmoTmXTrvGp+nzZhmZe
b08YvZ/xXUdWAcHDG8ywkYMuzXYN1FZXg3O3wzWh23Eocnei1W0NqmTQyVk0sHSYx6mzr06zqgt8
+qgQLikX/F/mLt4K81m7mOfbO9wWAKzzD7B4TCAg2hAdG0d0nudRHNh6s3pRR9ESHcLIgT3xUfus
yhki3iNIaWY+NY3ChctP2BHsveD8xPX1j0YhBiA3ryokHZn2H5khrb4kcrlXZ4R/HObaIbAVcSy3
SbQ/ITYnbphETUGGfWvr8AZ/0rLZkz+EJjKehyk7zJgsFPmQq7wQQBAsMKHuI//3joQFMdIqo9V8
Hd5xxiXtaqsD7OiKfYpG70RnoT+rAaA5IgZqhHZN71aQSGj1Zkg/UQw46x/AeJdrswo7Jir7owQK
DIJjmRdbQSUO4r33QKB+AQmuv/FOB39FaC9xiIb9bF2qob4rb2GKRqcT451+YUYtq3PoVfC6rA1a
H0RIt30hC0ftaDJ7IBfayF4RGTPwxlq0EcSXP4PeywMUtAqtLSJxVG/IzM/iFNFzbjUpxxpTqOH/
3S+teqproyUJ5/v54TPFS7Ch/B1YXRdMNuJSwBZQgQDbSdMKg/K5NDeL3m1I9tyJT3F9qMl6YUve
mZYOnXhgfLQEHSRerHAPr/U4m4gmmUBAsUO/Fru4WY18NyopWM8BvR47pZ1PqgMesAWWWMhacqmU
y4P3y4QQcJjV/9O5AJTWVCaJRW6gPhCfURZkWSKoEFmRtI9+D1RExBoU/+a+F4hVAELNxgPFWEMb
nIBUCRk7mM50UnLJ9YUkza7yVsn+v9x8ujgATTE82+A+8EdpQnDxrD/SR/9ZXRKlafXNp8MAAdjz
irYBrFGZ1aggJ04hWXoXrJcaJVZaM6AFqPn2Rw1MgdQIvHc6DiW0PA1FV1UDNl7jmtHrR+GfFCQf
VFp/0qmmIrO0t2eMI/rg5sT/8dhwA9DcVkwj7GgfCn3OacWDS4PSalF6h39CSV9R8Th3MB6CHK6I
2+4fIbabsDWd1ngw7m4jEcQsNLpesXk9lfRp9O7P8sEHrPfn4h1Cibfsxk8bMdqlZA0BlpWQTVug
0XPrzxCz6rrBov1BVLLliEN8rnoWxZrhlGJg7OHT6/KWKIaJjuT7+2+vZU5b+A23Hpyn6NYfEGVH
vjR0McvxeNLJfBdzroTjOIJNl/VjXXQUHW2c3ZaDVwO/6YDwhB/f4Kc9LveQ243UogAeN31henux
b+XYUFuACEGho/820K3eGd4FzsX3EtT17o/9Btr4wss8a5RzTG4sBihOoD4d1AnpC6P6GraBNqop
c2zNWJPcI57sciUdR4pKbDK1tAy8LrtMzQNpZJt6rt/d3mdyr3txVpmFyAtxDD6w5PazpWZkloLf
D+Eg7V1gV7v4VjeG+oezabso9eKBtw+MZQ/cwDTfGOGIKwh6VIkvLuIC7n/m9naxEEFieujU6qng
tZf0ATEoChlrGuKs78gvFeaTtuBTcOl/xR0M/0wuybCdy7Rqs4YY7WNvelYAH75MxRUc3S+blw8g
nUmJtodMvCclvrDdZZ/zioJOWHOfq1Dt7BsU3Z9VkilBEPzdQrNu4aEyBez7cHdMUhalg68qFloS
GGA/RDa1uXRktDtTxX37lVnMwORsZQmMKziohry9vujORSR/4TE1ZjL5kJu/DINgATITQTX2sTfL
Ba/qrzbcOdtR6ewezQTv0meRZLCKv+7eOKuoT0i8GuRBic3bd2aCoezSOAoM5yjMDnMMuIPuF17R
aPsUlsAAZWguMKqplISjFwHqLxmokLp5JiVxYRBe3qPls4ZTNuvFQRUdD7kzA5FGjrvKb7k0IZd8
EIFmV15SwTNUAd0S97qq7Goz8Ab7d2aEmpcRqEKEV5lBokeFZsZQMrOeoyhNg76UQT+vDY5BT2MU
z80OLJ0ryyRQbdZ081Zr4KNMhaMrmlbOspgZEakiKRV6Pwzn5fgVW0fNesB9UkL/L20WhY7phud7
sXa25pa80nyEPDDnyDXT5J3tQwcC9Ytzn3gCyM99odhDrXCMDHhonMdypm8cVjYMun2EsbkXr3CE
HRBHcgtBFwvssSiLo7yEGNAZP8gJl6ZdwAOhl6F/6hC+oJZSu9Nqi0EaKsjQ+lsBGVhcZLNPyQqc
78t7WT5BYT8FvBabSHVm+SZwYCbaNZ4BwqE43Or+vPm4M2VElU8Rc/e1x5hWOrXP8eeyrWg4Puwy
DSEa6byrsASkCU0mE6LuESxzi9zCnd9AnNAQ2SeAwQ559Ty4CMksqJSoePHg3UiorI9t6qf5zgc8
H2UNkiajQugV0+9oQuPzv26cPBNmhQ5UAzb9wSMEvAajN2cxqdQ2Fc8BW9kKN+sj7vFWQLVFkbjP
tKmoZkZ6d8CujkQyunhZ63gT5nY3IDAdqh7WZHrkidFx7QkI/7yMeiUvel1ska4J1H0UunHPzhGB
hNMElEQ4JhCiuP6L9N+bWLyFsgEGsKz2ZJmyj+MnxTj0r4icYZwcBrV5z0/8wFVnIzrY7JGlUWMV
E7ttZ31mlWoUnG5GM702/9cbosQjugDNXRvr+9jaCHf6EiSfLOCPV6o4Y1+PTUic4B4wM/zwURwk
TNoy4+mSn7UM6spNxA5MDwHU+YTVyPK7nxu5lfgjS3+tpnREUe/RFpgfnMZb0DCR6lZUmlKGuwOU
54XpcZOQtSYylqIMUZD198rC5OHN868oRz+VvvvfsS7dBN4LxIrr5EY7DPOZuk0GNpZq9SB80nTr
LAf85D3R8ktXBHJxzn4J8ZbZGScrGvprC+OTyFDyjYR2I57SzDCl1GRBb6AC8CgusgX8nCMyQZRw
I5V3QvU43g3rH2iZbUN/jcc6nLk2M50dfJ9dk5zPE/aEEaF/d7eNGbwVxNV+m+ZpFRYqyohe8AR3
hvYrVu+V6lmLBm7Ojciz4UGX8KXD+M0zKx60aq8yJZT/60+Trxp8vTOqUQua7iHgiJ2/Pig0/rRd
Dc91JRL6FLJLXIX0otisWdZjEr2PGNYBdRvWROPdltE67swspzRieiaJ0mYL19cTjbQ816F4Tpxu
F9eOD21+FDHvlxcDRSFwt4DQeMzBEN30SyevzgHnrFPOLD1CTHw/mRf3C449xo1AuUI2Ex08WQGQ
4lKmqFUBO27Qmnglb1wFzUnbjOoU8ez6hawF06VSKNxTPLK2bZpJReOyLRmUQLXylSADjE6ReLcY
fSduyMuY0MNTtkEiX14ITao32RbvxNK94PZzaI101i+WQdRZJVNUY7eG6BOW2132nBCD63wy2/nh
JCZJK2a/fl74VqplxZM7ZEbD/EDIXtIiw2SnVd143xElKZmYgGCSf+RZD3fk/puDl6WsDtHZRt0/
GJna0M9bljQznnUCP0VZfDMEUNxL2FRdyHgUZA8nD2/MeY6dfakJUQwXAC35mCFBmPs8KI5Y5x+I
Kw529qhmkHJRv/yPyfRjEqba6G8k/9Wp9uPTkjwKOv2nKFnTY0lZClV9dMl9q9TJTsCDoPx4KjjS
zTSObK5ghsPSweFTPvWBs8SQImFzfVNIj3TJbO3XT5KFk2rbbRxyPG9R8gzF86+owLVbQtnDwBSp
Bv3dITrxLV7A6YnGmdHafWgEjE0UnYVaz4eGFJOv7/+TZein1Xeh+g53S2B2WnSW1vv4SLJhK43S
NHpeJPWW3EPA8w2eAmBnBK0PpIiyFGf6DiplLuenh7Yf1X80sQROcC/oPJ2KPY5g4+eZqfA10NUb
wDDC67pKqFn4nkMXTKMeQ3+cKliS6v0AMhkuehFA2YME7hs1aJp3YiHDmwH/y+AjI1PUgPHxlmTZ
h10IqVRz4REttneb+VTvNa5o4GqFk0T3MD8Uh0rriwUTELvuA59WGW1FLBHn+n91Gxf/m9Xyl+GP
NW6Io9kPGehS9Uo27F9kTIUjSc/sXthL8z/tzIKYtEKEPsX1M8UCGqpFvzS5kh9RPM4NxL+aQcph
N4vCsg9caJFxVJevcxLKMc/GPgTxFzssqMWwbu5TrNLrqKBT6o4vdYiXrwyCSeZzRPUxQ5uJ/x4B
miUj6FZKYefP2PBrP1ScE3JiFQs6D4hfduVQIEAPmthzIpjFVemVLCn6PQ3v7mDSQM3+xi42Z+/F
n+cF5c9N47LYeBixzwVSBk4Q/Rc3gC8tiGJ+5T/pDzAYXLed+clwBeBeV5oO4MAPWBIJch71Leii
0u1koe3y1zDBEIuVTmO1Nn/qDnvkNjslu/vPONeHYxlj5hlg3cSsjpWr+YLTG3/YuBQZwIb9voWN
qbCiQEKtj6Dh63eKJ/TtM/nMwhrlZmayq9cuFvZB7jlRytf5DaXJQGpEGOfXgR6jrzHwAeiOloC6
a0E+6q7DYnttRuhzT9cnagjNaAE8p9ISEJsdN1v7n2spPPKYjeQP/ZmQZo0ewxoVzj9OFk/OzCYJ
RsuNqtvi9lR9cOxoZMv0rXnMwqFYEaujpQia0vsFb84BFjp3pzC+s9CajwiSjHNj5aHNIzT+goOK
fp8g8IR9DFhpHSSts+5QPOjA+XnIv4wzzgpFz4Jx2cORHOVCEgj/HUwUZTsYj3EgGXl3yVnGTm5v
lMfkBXdwOkLPNfjguXNeA1htdaEsJfAhan7QDiZ+1YrafG56/E3cZt2mjyd1Yly04Riqt2GWbbdH
q3hZo//uBHvUsljeNtDecki9BGD5fH6oCXexZYeqZ29NdYB03Ii2SCDAYYdSEK9pfBLpSgyt89CJ
g8ZPf/T6xA23mnED057JaYdyd1eoMSTu5tuu2X26gU0iK+Za4ia6if6GLDCJ3zGMbQT34Rjh8B1f
NGweZSX7sosLmp1acujGoNgVW6MfqX55IsbiGM+iQ+3SC0Fcq9oZ90D8HuBlk7X7A++MacNjywoA
8Rn6kRvdjpwOSueDBQ064WJQSAGfNQzWgvG1z9qzlAOmNW9dzzX6Gqsg/qi9mMR7r2+OZUHZU2ZH
FOu3l5ApldE1h12ATo/Y3SmPD0HtX+FcYizYRq4nI12r0v0TUJx6kUZD2NRRB/JeF4NYCzUiPWLJ
0ntFaziRg+vly4NMSkNFuO1+tMGy+N0Ht0NsS3WPlCebDC/nPZamMGLrwSpETudQF6u5/YsUUyyr
yBox82xEXXIG/ZQZ1tZ96JovN5TUVXU26fyM4ltNInhhjnndys+6masEl/6JC7Sb4ls29Q6z3P/y
5DlLF0LV4z2R0oSG74VLoMwe5cKoOucwV7+XUOARszmZdynv3pE1AXE96GUaUoy43KS2cXG2NHoq
T/N5RdLBoNmjvNssXPPHTD2BOoMttzlXCdGX6mBCGeGnMbrYIaOabf2u+ZhCwjAKgM4Kt3P4PdLJ
Zu4eiIWxaw55XufStwz+7x2Isi9YwwedSLljZBbqjmL9zZ52PkQ5Wzr9d5c1X+dgmrIm9xkVK3Gh
5Xvm+yQ0CJTa58ffWlKISQW0sBSguMU4DsblqVoGmWUER2jPKGTEDab2oA2nhLfPgyZHOJ8+8SKO
lpzVsv6k1BdSvUGMFY+v2vTgB/liH/k5cavphV/GUtUtTUqAa9TDr4Sy5IzLTPpO+a7Komxp5oKt
kwovwpSK9LhrvkaS2m8/8RZ1bIjsUEa4UrnZsK2oMtP/HsBAleU7aNnKLgrhjdhnTovQtefDx2it
+735A75ZpAh5xPewy6bQDTDbvmXoaaB9C39OVOfiAXeEKmXmrWSolkjceEqdgT6SuC8bqN3LV8NG
KcyvhE9Jm+i8E2jsL5qqRwv1zNY8qjrz2377c0TWUvO/H0qCsAMxQR00aLVGVT0FmOB7uh4rw7KB
/5f1XEAl5VgcOZhtbJGobYukO1vXr78S/92eqQzUeIUVh2Z9OgGyrInOwu7grXjF89aeqnmajOI5
Qrsy2obmailiB11luc7zPw1WcjXalIhoG3AwxjTx7iDnrZEKmrPTQfbKRovvoEdVd01JZ9NHvD1+
n2JALSYNDmygOrXVzeQSvS3MInAJxxsGFnMx5BpY5DVp5IIoNG9e6TSwekAME3cpkgRTJKwCEPAu
bdqkAIg0X3W+Gmh9c7KeKamKN5334WjuolQdFPLoaZhE7Di02JcEJh0vQNRp5iwRBp8CtcEsjXQO
EsWJQDvKRTccU8puBL7aDEuenwk/jjfnIGFsX0FPmaWUUg9F6gNB67RcNrdpp1Fes2qpimcC+/nR
ObUBWcHJKWYe31/ETP6alyhhZ89DLUH+44VzrReSMG2GaNZTm+utIEncHIuUtZx0lQwnjv/SJ02Q
aGcwVnd5cF7JFSsDOPYwYk6NsKU/XC7BWhhcQ6JvNcclh4IDEMkiucTD0BFK9HEeO8rFKyQ5lse/
+BAVzNXQFcsBev+Z92Rz6n1h9Lb/yGn9gMPvdMf/0bsMxVm8+joBslF3B4GxnG/XAK4pBjlB59gG
wIZ0e0YvHpvqgnOeDs4lsvBgeH+juKREWlep0wL/3I6PSDFMkGk88hYGUO7SYMpXjr4QWvESYcwz
+UsGBV32R67404oRgUqK1w6GbfZd9pCfYb9OmiLLh2u1cO0uhQ9iU0+vljxjWx0QtlYkkbJ5XOeL
fSiMBZ/EYII2argDXmQPxIcR46FI7NOTYoLMaqinHU9SjS5KtRO/XJmJPoDQ1bjBNUewOTL1I0Eg
9Tv0fD+MnjxJsj3l/9djnCYZr78C9pfW32XZdWKvs/HkPcbQ1xDJRHTfVbd0Lc9f2qiFveFyWL74
AZ73daBvtb72uLeemK0sy7EJtZeXzjoHhd+wrCVxXEBDm96S5fjPXye6bMAzrmKSjtqJbyq+MzxC
Zv2f2Zc0by/Ivwe4pEdiy+sq2ChHtjhphPOSncTZ5fiuZHtgc/n642Ir2svHgtR8D86sj5hvlwHE
5i/q09G9qNj8lG5TrgK/BH10JQcSzX/b/laGeA6fyCdmzI6Iy7/kWFvTSec6XFuxosfchj5UOVIw
MxQNpLhtAbGPWnVf9SCPV1HK+zDDQFMm8UhH8P1kEi1UQZngyfKhqJfyBHMGcevEWa4T0E89Zsrg
njbx24dGVeFJdkBY6jjDy6Sd9R5MuhIcT2qn39pELGmYh7o4WjXHiKraJKGDXdSCPWCmyMD/9Zfx
QNrcSo/3UXEw0F1AVhQvXC57jvzsYW/uhqp0GE06yqXOXkGK0EMauNtz215uVNWHHlRFtSY3V83k
aWlDS4WimlH9BxpVxMMwxQOZs5YB7bCyIil78YwRKsrvU7J6UlftoDHhvILFXeCNOMHQzTT9Zl5Y
iva23qXiNbbsVxXVVTd/dAKiPW/6Vw47v5SYbngRlVbg/4I43iBm4X388JVe4WYhJ+AgTqCKNXm6
nI6aa8jJg/iNCHnGrpmsleN4qiUcOdq/qJDEsMU2huOsShLCc8CyZmnnUlNrZvoMP1XkxjVJ49wq
AF/YYIsCOOyniG8BxzI4mzXnpVe1t7ca0isuwmjC2NzfVbCM/v/x6ehJ4ia7EnjVmbuQjIfJJIJj
Jm7onPzVKMh9NuzZOSIzofjFEZ1dnRwP9E/OCJL1sqVlJDKG/wMibj3P5hDG9aLGG+D71G4sHLI0
u87sGuVm8S0DaNjoIGzJdoVnnMVjDJi6VAgS0r4r6WuR9p5x/ju789PKXKRoJsNhYK1MQKCkKWC2
zz+HI87D7C0/iqiow1OgLSokZBLFdg7A2HBEI4K1V0Vpds/LCtWB9IF6j8RhhdyWys+BRMvGfntx
vd5WMXR9RjSB660scWZGCsjJNRaYf5J/NI2lDFt4WIQJZMJaRtaOsmLsO8clDlexgsVPQ5MxU+Nt
ahUnWZSrAkxXzZajBZ/wFUdL0HnhUDs1sHdYPj0I3jBxZqTD7cgLU8+/k92ab46ZybH3pFpafGUO
qnBfwJfM/XYElUXZ1fBJCeFuisyEce3u+NWgkUBtN535hmf8Ny4kWNKknLnaBGJISXgngDT/qdFV
gAHN5uuuX54VKPetQ7NyZDybxdVZSyLBhwnwQ+coViKWPMw2L8kxHj7OcIa7x+A/0Dq8PWT8DS47
/RSzyZQLjwiM5m4NqCbknuj2SP8d0SCvPAdVSsP6lzIKI8jfyzjiNrJV7U8spxp/Q40JFTw/1eIl
/dgGaMUs4ZqyM18GKjfSMGad6ZTESZmODx/nFqdq12aS9xowhD4luW3zF5Q75+PZAbLyxKz4kD5V
PE4dfNoB208CuH3uBu043zL9qFn7C96XJVDg+qCidLkQvgfptvXQ51Ya3sBueOCDT19UolaV3Um5
4zECLaWEEp8WJ92ee/GCj1gFlK7YGVSq1SISooUKTLvnJ/BkA22J4HeGFVyoMlb02Zt8Rl+7X7H0
D/9NeyvIuIKLwTW9CnwNu7VnwVKrZIcZ+pzuzkS7fx8oVCuPagL31whmGxNJ2s3DYsoXnkIE57Qc
2AjaO1tQ4ediPZsbTb4FaGdj4JxvaJYDxyQ3JPoIj0q5Il+4ykdRKZnHBIQ0e2onNJ1NufKqXRXK
zjfOikGYZWaPQ2eNr/S6d4zaNsTo2Y/cMxrN/FwQxg2Y62RkVRzm4q6WgRZFafWHM24O6GzcSIkn
qeJasjM0D6h2SELeXorNC4VboI5w212goiToyfcnNFSycilOMjVeA6oqgxuqjcG6RhxqQzIW8TUB
qtqn2LoO1VsgbTpvIJPcenUCtKnTNO5ikfp0TeW2XGonHQin/W3amZthRmwTC5C3OMm0yZPlj/Zj
qyoOuYq4rB4NdIwdxDGw6IicRI5RPHVlS0M9oUdTs7zK0QRTa3i4V/hrZnKalCNCrpZWr8bCIzMg
qZawl8tj6ZfGRI8bR//TZsXABpUCyAheiAX73G6Zr8sFDEtQG6HEO2oM87SwSJ23e8oCCZ4UiJY/
usJfAViVYG9Vwbq2BZfFUp8mm3sKi8gqtI6JqJa+ZLIA92x6ht7UIlnp55fyIysN6vvSKuojAADU
pGB8nQuT+Aq6gLLqcWNLpcr+6hqzdR+8SXeIw0s2Y46/2zi7FMow/M8wVBcjho9eoSdMlvi/uYVa
Ty2e0dOyoHLaQUnUljEmaWvkcssOf7Wp7/iyNXtz4UHVIbWjw7gzWK9PpS0smudRTp1kRzMY/OQr
zriQD5Quu9rLGI492FU0sYykyN93/wQ067wzCWjVBSoGR+WQRsH6ooipUxMJaqjHAyXbsZvbTZbq
aV2kNZGyppAw2+GmnyA5svPaKqj1MOJjacccw14vKf/BCTWeCZYx4YPthRFHxD+1TFrqZopr5oAt
vjKZe7ecywb817vYjWFm5Bgk4KkWqMs8kx+Ya+jygzT2nu5MGYdp+jtfCgeulQd5tyD8eHxxHCj9
RrKNI5u4Wge5HdXuNZWoxV6ovyD3xSR8x4jKS61H06HDWaUDQnPgdJBBb2d0omuuGuHbQSzHwIB+
3+8Go1ats5UIICFuw/1rX6FRUEhyk1wVG9ANUcORZbKxGA+kekdygGuDmJJcAwHVUIKBvQNWj07I
zuHT/6YcjuG7WODqW4/chrGH8jpWB9Qd7KNqg98DsdlZjQ8tazwjUzzkd6ekbG75OPGhSgTIWqLx
E7jQqtDPp/wDOSQ3mCZqje07WPFBzXLTtJR9/ucgFjcP/cqhydTL96g97Bm8IrxLFZcxpq7YYJ/x
HwdP59DqFV3lkvdEHSCcA2ZKm2X1BMw96kJsBzEyEpviA68ySueg86P7pCUJ9arkI+H80MX66Ehc
ZdC4cQXv+22zEhiOczVpOH9jdIhQBOzGCEa8Ha9edT+lsjpVGFNr6kFkEhGqxPb9WzKXuK1h8Brv
mVBPy9e1pg4/rv3Yd6pO4GuAacH9hRDK8X78Fhe0vXk8OBNM3Hq/utLYwM/ezbOO/597cQuJH3e+
g2Fl5IlGlJV/FBTqlnwU8p/cwBWK2uR+vft/tWj+LaL/3B2MK47W175LJ3jzFkd1aHkIeUc5olO9
p8xKd1pw95jbRGQ9Mo7LWpm5UPUBu/xB8anJ4UftqShc9Dt24smkS11Qzp7Sg45U6MGRP3xdgc29
SeLB5iy74ZLqFAvaJAkYlG/eLH3EqJlaKH+91PYCRv6pn2D2BqU+bw+f12Y6IFmmCTmgJnXBzUNC
6ADik0ybRstkwNmx28UedX/baYq5D6HdctUqs0MtVboe/JC+2CvZ3afj7ewD6zbGou3d5BORJeC3
rhLpCVNu1/vRJyPBEETWlaBqvC3cdp96uqgrZB515E4J/X8FaBQye1+I891WJnGfQ2gjvQaY59bp
WeVwJn5SPhePHbAfSwjgvbWbWXDL50aTfWl0bt7hit2GPnM215KkfRzoL0Wl64QlDc8tTvErFdsC
Jl2BwIIvVjv37hMDpidQ9Sc5jfpWYbep5da0PChWz1qqw/SwCnU+jyUfZqYugpkgSeVCkEgPIPGv
vXgKG9AWsFnvYxP3ZC1/66T67AvO39pXJXAEvEhcnTNUMNKUdb5fc5fQoA1wpA8yldl8nemDDd3V
wuxgWVOKlGuTkIVKoJHJBEGfThObVaEh+v0i8QVpJ4/AwnSgx9sUF6fme3iPsPyJ2CssouWvmIJc
rXfnBqABBFjDwsE77HLU6tmyR8gDKngwGNxIZaDycUooaA16e2dGuwcn9dpmXk68rDSSuudVfOiP
mg9wQbxHxHBbuJPIjEVKrTCzIBAwNLhDFvISsfocz8oNgtnt6ySmMJet/dreSSuua91iQQHbSc7k
ILshDhwyGhnh4F8wlKzw0+cjxj+C+/8UD+U+Wvf8L0Hijhv1ftswyb4QlE7Dyt6zlAR8qXNURZqF
exfVcbebW4paKEZjMZRkp+5m3vsmPW3LnIDDhzSOTWbfPRQPzz7dDLP0lpNIUAL52TbDAZKVwQby
w1r68fMfVw9woHrz3wl8ymjR+x7zRWHbeJQHUfAPaVurbgPe7hhAQ4crCFtn1NnBNz2tFa0Oc23z
dBrPjzEaNKt1UhBUgPJgtPLw+JbsiIvDKKJlXEO8KGtsynL98C2w/JaGmgTZ5C9wD28+j2ZN9M+U
vndENMLC/mX0Np+VHNAFB2X0xiqK3WhenIkxFJd1JmetMpyAeUFJBseq8V9lUeEzeXJRDirrtJiw
upCGJW99vy6OhatU0TNCAOVkFhY+nH+GJkejFNBkhvAwj1n0UmjuxbSwdloiH8BGcWYtABdxCAMx
oR0WrilLSvMkJ01zGGXzpe1i9L3EIUKVLIzg1tQBpVgMw6CPLNQnbfalF9HFIV/Rb+HDE3yrmoh1
BQ5hHRddEBBK/TLUU4vcB4mkmlz8ghF1G7c/4Lz7Ww/PJXTEWOHgGoSk7q4RpuTaMgSOIXa3EZsM
qiKJ2p9EFED8UZvSv0DF8hBO6GekLB4DkRyxuQ0f2BlvWj8CuBGN5do+0/oMubJ2/m9lK3nU22Us
DCpr+6FBIdnTdcFpidrID8BvAqGPAJI/4O6t79rwarpbGipsfG7yjS1LIpRauQVomZsebptJzp70
n5qSAsP4ZavvvV5hYI89EQ2zU03+fPiBvrmJcv9/4dzrCEJotpYNlNE0sB9GVDZX35NU5CCiw1Ff
A0RivBhBeyTURc+NHMaZvwRWnLZhtTZ64GYlUzFEx2RI49hJayJgx5A8FIxYX3o6mJQuDdfmjxE5
xm190iMUyvEsI6DrRTvJE4T7IhNzFZ63oXSjPuMgAFyIVrDtN7gxI6uYaz5fbQlxklKbF0hUbn/5
UaoAjnnR39XFRDs5sVGsXlHmOXYohkYmRo2+956MGzILyNVksGXGkqtScnsit4IXwFObnjubpiy1
Uhd3eeVivsqcPKPru23g/Y2VKCcdoLLMWmi5FxU2fmEQXbhuFPDDRtBk4WUyiXoUNKzsglyp/iAm
JZuvXCSowAf/qXdMY+QPvlrLPB6To8A/8ux319rGsxPybiR5DJ5Yqa1Z/zAAFJDrpsXGZZ82Oe8r
Wpwb+KE1/2mg2RtYp6s+K5Y02LtUblc+HDUEgiQ9QykcdzJ8C5GiVUSqh8z2eL1+H+HUSpWeDcS0
os2LszdMpftfx0pGB3SUrH5bzwG1ZgZtymPtUAMFdXQY/ORfgAnlgSv7OD18Y7knV+I+Hl653d4j
ZemMvJtrGYwmAAzrDG+W+GEDg5hss8+JqnnFQIFMaBuli8S13COHpBvguHZYhnPgJP33lTi0brHi
ouoMYeMp4zrRLYPc/LvR1Kxez0NdHaFS62+klQEdK/EtQEwYRd8kMWqmY/3UbjKS3tUyDYMuXsj5
BfwzjAP+JA1sQdgKX3Dq/i3H6t7P/cxjXrUhJYtx33pI0XaVjff/X3kRsCePPNT+9VbCs8CJEQGC
JtJZbpiVIhUotts90H1AAhM5HI8hND9MziiLgGktnzNUcEVFXcxKwncReE7iSc3ivUVeQM+g1pwl
kuMaKxE2l5Ea5wWpfP6cZ99gkG5uv3+WHHF5F5XPwX0TnvsdtI0elOBGvm93xOsu7LU8oeCJQXFW
Jacm6dduMuPaWo5hM6UBdWp6wj+Y8vUQRTa+2w9hc1iX+RUa4mn9layjUfxx4qouI1mui9Yh8L38
K8PRXqW5g2qFzDWkRKT8xbNnJ3vJ58SBj4fl1BwtbDxZwtvvC47uJvGmhqAtnSOVU/W33AWsN2ik
rLoMURhQDCRWxPQ2onCtyA9nPzHAd6pvVd9Y9b1Jad4ykKxthJQuna0/NSvtTfqSOOpuKi6ldtCS
tICnKXKPWHJ2prQf/jRO/vEax9ahRlZ4wtuHAFYcRFzt1jhbqsps6PbI7vuMoIjpSHaKF0+Pti66
kKAYiC9JpNY4wmzymZunIQCXi0ZmxbmbzhV3ynnjvEyUA14tG4EXNixm5PbdB3wE4oKVict8kIAv
qFIwdsCZJVTJOFgAOVv1OZgArRR5IvFyhZRaiceQDeuzTqysQ2GRpeqlkMB0/gd1ABRZfApduORk
WKLD0Z9o9TO54zBi58Jo03DQDHfA7319mHg1MqWB9JgxlXzBKBu3fEE+iveC7YE6XVOerDEnR3Oc
V+ccJxEP1tDjsVL5AWbfhhpv8syhDdGo49Smsl+AdURk8BUjyKMD4Gp7Np+5l6ScmD754JJOIwrc
//jZakq5iB3wpVI6hAWBob4sP7lEOpLmspGB+lTEmvUyKzWbRSF4DmR9PwUOwEHUixyWCpGlIjyR
xc6w+a8ARy0K6SEJG0byXm3WtLQI5KCkLi2AUPTIbA9sN4ZiSHucsc4elXwzgmv8mLgeKMh8N/51
jQiOrXbj1oumNHQybRSPtjFmdxKiFIGkDEbJcw8Goiw8Xg68YYw04t/EB2iTy6J04cE5izAVLnAC
pn3ekXHSk3ZqhFbVpR1cTK7Khx1W4HHVA8LR7UYURKF1FG3Yr4HGWMedMKViyaK/As8WZ6eRaj2j
jwyPv3he/dIMcDyZdmDa9tklnWCghmr3jcBxuTFn+QOOvjy70QC8t6ngG80e+XUoEX/ydktkqdAG
GhEFEs4S8VaPc9N4hPYMkA4odpe0paoLyvunngBGSWTgZ7M8WytlG4a1v/v91iQMT6EZG1fR9vjd
PHa9KMxXmzHe/982xu8/aM1mHwTDN6SPWbee4may7Eg34wHUEwQkW9nxH8JcVhXSgls1PeaSQLmV
4J8Fwnop9OtRIWsNphNKv4j6cKFvsLkR6EpJecGt1eFJi9P3Iiispnf7hGzE8UlbHaahJBsSqszq
ZEVN4lZACDukTEl4ID9J7DOizlOit68hl9w/DCPt3v4K8jNgdziitCN9u19OFCztaYS+YfmJO6Ya
S/xjNIliuYSsGPQSToTIEEJAqEI8iTUSF8L2g7AOwxChgWtI0OUezoFEj2f/Dwm1uismL+LkObAA
KiohfcfPuFPBoyg5y88rGDHVy6ZUsH9K2+58daPKtejnmOAlTQAGO/BA7Dd514qUyz2igFsC4upf
q0zzivHJQ3JrLW6UjdyHISb5Dwp0eHBD8GDtYsZtiaPKhLECY0t4TCOno1z8wiqYAF6P14xh90FC
EFB7Lx8kh+jIKmq/VpKOHNETqZZbyZo3TvHQOFu8bfiNY1MJ1A5xNRbA0DMxThPKN6dE3Tkvsq3N
GUFvouoKeEigw3axQdEHc/PbAu4PWQdl3W6bcz7Cm3Td/1RJn/yQfx1hNjH2C6xKkj3pR6xJVdPF
lTs9VVJLjXFm6epV0CRy013oVPE3dzo5v0kk2liy+3NeArD4QjyU3celGuOWRv3+b6g8y0pjBCRs
FichI2fo51wwzOhQ4vzzusNuB/bpJNC/UQxpjQfjYzJTUK6O+RRZB3uurXUABIGPndJDLz1M23B7
o0sCr6ATaZJTL1ht0DOjpsI1DjiQFWHnwmBeRj4hr5FDHyfC+gvJU0INjb0UjoNDsAVbGYzDfpyk
mUvToLJffwc/3FyA9Nu3bstcUqGLAfO6e8WC5SDP7S8UMFJ3ptc5Ip0UbUqQDjJHU62FOKK7iiV7
HaVhycOmE7KDQSkgyYwyAKOCJjge168Yr9cMpkoD1zh1E9VIxBqwy7pB8luWjp1L/5twHsrgiG6E
7hjYSvp+7fgjvVTtBjtcplK8G9i15HkXebL23fGaZqMYWLfF2aREWB3bcaAqdOuO8+V0Kl6YJtHJ
J6oCZZvJOUFDVWD6MI3Wi7RJi+ShCsRO35NGcQ4ulnX6eG+rctIDjJ/CzSB4CVadZ5ZnslFj9PJw
8jaHM0v/COks4aA6e3Ny9b8qllerMIj06BK0AAbG3tUH+0nDSkJ47UTkIQ2+xvxw3A9y+ZJ/pEgN
mai+nZX+ujUrQAbj4mph7HIAyH9+gP4BPlo44iwAvprwLRgrwPkQW+UoFPUIHiaYRh3wc3l+l8oB
51pclYl66TxWOluUfXrSoTV5HFdnYp1G6Cc5eW1mtnK1MpfuwY2OQHR8Jf7DvbzCOiVHRER/AljM
Bd2sQ2M4xmB/xAuc1ODSmlg1ofWaIylsDAxct8haB1BhgV5gm4LSCwpUIi7f+WlDZzAuSFhGt3PC
wB/3YroeaXgQh119eG44iazwWv8mDzrvHsbyMTjejrLd9EhxOJGaz7zB7mezRHAeJdzk4czg263S
+j5+R/gb+YWEyuz+1lzz1lQWUmBJHj5zEm1oYJCoUPszumfQHqhdchFuC3FYdoTZroH93JDNCKSx
j/eTjZJz1C5NbetnWjCNai+Jm4LrJtgj+qUkDhJyJdVvcagTgwEC7dMcRcWBLovbqZZu9mGThx4Q
qvKqro4656Dmj4Y2VgkpvF9zc8TVp7JPsLltRigaukTegcMmnOdPQrAOGLBOWvtpHQ5YQJN95Xv1
+5dBzEoaMdyo39wIQVM/zBE+MRYvcPXjNOh6nFOD7N7sClFXj2D54wnjzyKHCwPb0KMaS5Kmz3ZB
UmODM+prpg/9hG0f6h72zGLwRAZaHMaBdk/pwQ8J3e/ZX35qFymWIXaimuKqq9Kbg2EWrXlxG6T+
QlYcoNZ/wd9QjBo7jzISZl363nJz3u5r4MBjE/TiO7UGCSs0snGdfISE5COSL3L9Ml9EksGGaxMK
zsjeE6nuHyahBGvyp+F0hcMenYEFS3kuYz5TN0FjKFtg6AvJEvCtRTFlZ3hh/YD8S9H8VeGGK2Oy
Tmfi24tvYx82+yOVtdlY5wNMK8hFPk/pLv3WX/lznfB4AeQ9N/dc8RzTqotSqrzMGbgJCbH4O81f
OLkQ5C1oBwsgMm3fodDDLOEX0fNtlPHcEquNNJLb4kBALJvR1MOVpUniyTa2u0Gbdp4hIEiQa+0k
6v586S3F3FaaAOQFCTUmXh1ZL6CK68NEsSJDGy5/zyjfwuuZZw5DWuhAzeJiqjbnz3dGpuVzMHOL
UbQb2S3ejBkme8Cpue25mVXc0U5N+jq2qxYtavbwchI0Xuae4D18wpn+xPwOfd1DStJKlTAjvVQt
swtUzwXcIOHQ5s2S33W0rP0nAZHJBxSgitUoXcyaJsbFbMgaropU/IRpNeXTuMvB7LzqKtV8pBCi
wKwsID1bpqVreYJU6tAl7FPiYQRlzlIKysiito1LjuKhqx1nNamQc39QpCZLpsMoBLcLu+qGp5aM
E22Ec/28uovnsNZf9CVyen6Ry5GkxsSbl3Yvs+TL4nazdUzYvjq4y+KBBIC3+ju6gAGUH0sFEFs2
SVCUwyEWQ/fQzY6sb/A+1upKnpehg2s+D33pWOgS0g1V27GZJ09adgtP9jJDInKHUJJ3nZ1zgT9T
nojVyPItpB92PcW91T+0oEr3e/uJwowaWUol+b/zeQ19kMmZIt6/h4HgYgl/ZuW/YVhGQidW+mwE
ldh3HQ/eICNND+p7k8UNp5ExZhpnHpMA5TOvBbzNti0VERxxFiTka+yFegNxORN4tGAVVyVRecGh
qNZMoQJ0zaMYRBZH8BEgJCOdEXakiW2lPv5G4CInPsjubA9MKKXw6GZjF+WLHrXQVpH1oXJoUYd4
NOhO/TmmF1fp7qvj33AzYPh59DvfZHfoLZVlPx4nbfeiaLoBDJm8bpW81GROxNh27E5kPRZWS35A
uuiRr4UMC/vmuf6Cwt38qNPtMkia+HaYC822/W783H6EgA7Cg9w5Pdj/oj3e42kHTrdLZfUkwyBT
wvsRwAg1wgtf7tUp/FpSTH1dg4L9OoivmnbzFWOrhZaRTRx7dHxGdIftZFtXDW2/K5JGh0nmwlaf
HveANtCE51h/uJT3AzrasC5EsNwSilzn0eknvUuYx0hWmJRmR2aFBS/8RDGbHwMvY5dxDz8Mcp++
KF+663BNd9h/gc1bz896Vk1pdnzDeHtfL4muxBIGsMBIPcVTqHO3KACV2Qvz70KRjR2T1bl/vIS+
OG/cTQYT1P9GAfFMeNwSIUEBvLIVocrXdtTN+Ehh+aaC0nIA1PF1ogMV0JF11exEgcUtdXYgH2kf
/Im1dVvjtZmZzBZvZuuQ9LDDbS+e72ZJolYPObp7/ANTF9/uU1xIpUpquxYANtDWqAIaddBCV3eQ
l9N3RPpxaM5wnR9kO7RJha8GS5A8O6Y6ZmJSUVnbquYpCilskFoowzjrpS7q5qTF+H7MKLiYlJsk
9lrF3oQ3bxlgGDfefL0lAYQMV1EvgZUeUZcnYw2PnZbGUqL5CM/pAQQzTOhhXjY/i/Ms6H3aygR9
YXROYIAl+UsbdSuToFubVz+piw6t4Daf9h+joHEd5cKiGTEl41lDKSsxftwW7XvivTFVKk3Z7v6K
0ZVoXsl8xdIc1HCWQNxvxjLvS5TvaOLupqX//0jlMcniV8/tDvqsCxjNkStdMOM1+/c5z2+4BWt6
vzxMcnkS4IP+QqfbhK6Fdi+Okcvf00ibj6vDLYsqeoTr1C5l1cMvZsAD+c5Av11rIAENeAk/d1P5
CEg4IC6yP0wpmKIfmwHPozhHdGayBbfvl8obKPldgyczN9jHtte97cHKxWoi1/fEk81OSOzs52ec
qojGcj87A6o7ZvTj9QGQ+6ETqr61wgVnPUqVJntFW3qw9vafQAy7pmbuVS6rrRYNWVjzaeKw9vd9
1LGIphMDPMj/rx5YoqXUQgH1zLPd/IyP1MJjsaYqwa33pwKYejNnEDpASN+qoMmLVkZwNggQyOLq
0VfiznIJXUnJ+3op+ZttJw20if5tOzm5sqyYx0bGR7LBkVd9OhOTh+bcaZ/2fVrYOtNZFlmC8ROn
bAudRbJYI8/2E/4ZBzh39ZgrfFtSocnYuQ2VQ71fNqd0d/AQHZ8lL7pvuEHXVZKGyDqz2Q4QcvzN
U2iIKBbjYf4beStAF9V0yov0GsGlTR0wKkUEziXyhKJMuqksHU8xjOCUtE2T15MFycXVLLjpxhP6
xb9ms0QMF0xGQI3tdmdi4nCFphiStIVe/HJS877hprkMB+gPpk/WyMv8H3Zhlpl7t+Uyt9QVMneC
bxLLI3ISg1O2oM1k4n6B3CHRnqiCaiW5qvlNMktJpP7xGz5w9hEB1qN7rqlQhDXuiLqFCjmhlD0g
aWz53t79WCblaT/cOtyDcw2D2Q2NtpEvhGSL2nIt+oMdBHWVUUMR6mNRsdJBKBfkzNqn9zz0fIUh
o94c5t4qS7FhU3us4Od28JW1Uj5DRnICsb33KQjSyrF2Tre+uiF6ouZ1rE3AKPzmnqtQ3SBSvA5o
sYX5KTQ0G8f2AxcGY+I5kcuH4yRuW6pLCLo4TKewdwIB494tCvZ774uLwec4h6h63VTXRBXREU3v
ySIqFpHTvmv+qNWOrSXHSuIxFkeHGIJ3fR574cSMeq1X5kApHyCsgokXSLWrVePPiHz9ViloA2N8
LREgt4ZhNNulM2fSQJiTG6dRYuBJD9jaTtYbJqKHBUELHQ2l0dvJxP5tkz6BX5cFRCXGjdb3qXbL
P42U+FgDfuQAlvMFB6ahi0gSTOFlbvEHcBCjUQMPrwAHhRdL0aBey2QMC7J0Hd66nYfl+dZ58Mwa
i95GL7MsFvrl/sToIdMk95+vBSYGc/tKfy9UYSA1aMXvYCdcmdWmYBt7dPmEM6weDZhLLzA+iZNX
7i0ggZ5mvHZHHwLz4ecOOIDFa927vyQy2MEEHlp+hnGAb3kBwd3iH+Y52O8ELQe498TSmBn9AqSg
qjjqmgApwgUx/0Xa9CjUdXnbcChWay0+xTX0vlScSYEosTLRuUa12w7tEolllDElpXCsd5N1h74c
ormsm5P0oCma44zCJ2K6h19tRS0t7ZKhMT6c//2+iOm+z/0pg6Mys7YumYtVhZ5O0bIo567kZ1mC
J5CuIVh+jqjRr+OQc7tYgxVpxHLOBCAB7Q/Kr/RHKsq0EbrAkVis7Qs/n4L5Wa77hZzG5pZjtCnE
5jiYg3GN9IBDZxHtLT03mjVYqy1PUtpb1s6H5jij5XAMOqGMtDXwyxZsA563ZGCEXszlQ128gxeO
FcEfpSDQO2/uBucF5MDVQm+NcZ8k8fRKghwNGI/lvCezlh0ignpGcvAQV5JAzlItk6USntIt07Lw
F1yzpPEsgnSaiNq8j+hMWhzna7QwJ4569V4D6Efe7imvCsb0L6eWwW4w8Ht9umlPVYtho+BHJu2t
/js8bPtXAyDMQ5pXO2EHLQFw/uXNDtzt5HB5vQJNEqBoaAPEl3njEu7Fc/KpOcQ6nOA6/ga3rn6l
6glHvoBsctH4cUfRzsYIG8q/Q7lZD/SfMr+L00kZ8g13CqlGjnlWAhWIAK4HxoZOpBuhkQKayTeg
uaBjXOIjI8PIfXplGTqnqkDPAwmFGLSZDh1Ut1+IJb+ZylONkcRv9fyYOwHiFGUDK0PALzkA8VqB
NuXV3oCsLU4g7pdQFcmIHuFwcu5QXQgzwjSl2k5Ov/+SGTqLtv6VuYKEAH4ZUjvf1e2TMSpl5Ofg
YICk4wVfIEcCp2eizOV1VsIcLDIklkNksNigCf270xw24Suud+mfRbPKaBbHvp7Zslh6j6BXtS19
TeD+hi35qno5JRDnrfFNLcqp3RJWlaXQsx8T/JaCpNbyrlIDueL2sYNBRd6riLvoN7zsukUS0cfn
UNvkPcLuMe072ClTszVGWE4O35ukpdBgHoNl7l0NqRTyDz5PhtP4NEuEZStX0fXRSDqAj7gHK/3t
NjhplR8ADFxkiUjN9tCVnTxgYS/xc/aQB5YQVgS5L8lhKC1zy8Q4ba9Co7XM+a4gUpeqp5OojpVg
snLhW2El4kl+zr3z6UjLLvY6Z7If9C7g0oxXLD8al7cRI5JEIqvnWCCojUJnC0UYgz3EwKMAmNxz
dnjZjM9vC4mDdX8UZYH9V3wXJJAyNNe1mZa57xcTQubUrOZH4ZZHx+S4t0RvJaw4E5aTBapcRNvd
34iGW1vy4zlykASn9GIEA3reC7nEUD53du43h6h4sNPXnVV4h+EGYSMo5lR2piK5IVFE2DjZETtw
tuKzP5BN4jfdxTA4sU5Xe7+OT5CrlFXmz0MbiYQ4dzn3xL/hV4WWd98PqMor99LFe/+bCNym1Url
GfbH+tuw+ouZi97TAVtOyScHMqWOyGrb4tzIZYv+8h/gbTtcjRFzgHtxISzExEfbqxGn9iJfXY3F
GfQgflVyay1Z3QqLciGVRvFvdfQuK/Y8uI6h/lozM1z5cR6Zvp6RfAznEYKIpq4diEmz8RsWO4GV
rSKtKeW5m9AO1t97zn+XcSRtC2kBExVJQkTafwpcxHPKpfwqqEsLEYdzVsNc+BA3T6vZe9DsYI5S
ys/j28AWQs3FThSJrKMEUlemwQr05pgDwSx7fI5HevFyuoxax15gEvL2rSXWrXQ1F3JxZLpbPxlT
NkR12taXSYwJ+oghCkl20bhGbtYU/fZydh8ocJRHFm9C7t4XAg9q67t6KNhTXbwsoQ4qn55njtN7
FDuvbw0ZXotyViHrKQsxeTNPuwCBF22Tk8PFarCXMHws1f3pWMi7TO2Z2G2bPaEV8VJ0vUxmVoKR
dSkm4PPHMo0/i7dRW8p/KKzsL8VQ45NijDbGUPdB1yOchmpx1V2odrLrM4Pen+BzZM4BZvGRrFWl
gILSzMh+Vwy6bHgNWv+ejwRKbrCxEDgEr1gmH6+OrqSBiOcaCQsE6d6GZIjNOMbskxzSPP/+DIya
f0J/gla95bCQwBnwgPFcsrKmHnzLO60rqZ4a66TeBNZFuRT1oAg3osMzXGJxsubBY+e7F46o+smm
aVoQ3Fq1uTcRivDfnFChIaHgCi9N5Pv3pgKCP5AisRaJIxscTkUEmMEPCmft/755+YDIH7m85QyR
1T0K83BYQ5OwPAZd37buG2RTS/Rvg2FW+HkeDqmIX4piuaglmiIB5N0sY2KZX4ycgQzks/tDFb11
+zcNBF+lWHt3QHiKjpuu31YX1syJl6q8GEiee6cNl5BFlXVMzorrPNeNXwu0jQZMGFUPV2OZXm0S
hOe6EmOuGBgAoJDu7P9sHtkpJdxFDV1GZgy+EZiUDpZ7GQhjwPHa2I7+y80aaJq9eeqHUmEAzJMP
Z3wL0QhfdwWG1cknIJSP0VoD16coh6ZuPI2xICR2UC5gGG196Fv4Kvu+sCRDmXFYXCIRf/04n0Yd
D/3S73rb64fye4/JlN1SJcGFFgeE7mmVvZ+qxu1WXn8kSJCft17PjjgCmUs93uiGvENTOmWQIWuW
ROqupuhDalp9MbFx4sFtk7+7jWK+wBpbFJ73ZSHSf6e1+Vc/Yv6NnHTiK/JfRel2HnaCdZ+eJwOV
1GxXPRPj/Ik/EQ582tFs7mVem5DdtiJ35md2yzlDG6J41w8V0ugD+Vz1/TKfXxp8fVXnCIDJZrD7
tDLS3qicRehWlkguzl9aqz4r+AwEy9i8VjJfGYD/8MwjgOU+EJYPDmXZuarub3tg5UdEY2NlMn6X
kBQfsrpf/FwKmNVlb7fSoy6Ve0D3dPALS7JWIF5BnHygAFDi8eiY3Idp3/ry1naqeNdZIpceMoHf
DrzpTljN4VFBrmSXcEvbqE60IpJ1KK5pQNGFe80RBRvjLbzQhVvd4TlDDXpmRmhOgM4z34ndnwF/
jftR4phWdtyiAuy30h7Wtl5CejlOaMha+5EyXAOvvNhA92P5P/zeBdniqVFmTdQn4I0THHQcvqzD
UDJ32TwE4j4RbR7xLFpLLy7iyReMm08LS5bGspgksQ36LMw6q2eGfsL0/u8zaTdcgFmopgPdQgVb
yRnUC9Z118YZYXuexmDY7xQEiaf8u2DQVQ45OR19xGZ+0jun16WAQa1+bBQeU4OrHT2t9oLWKrkb
Edy1Jdjn4mOIeiAjJAieMZJ9zdpZtNzWNfVSgibCrEbpYybgmrwvm0VQSflfmRaGtthKpynId6mA
in361R53yoIiFjS680IhbUbTgfDiiwCm9BTIB+d7CuE5IxRPT8WVMcX6qWRDqvmjjIWQmPirbjSg
TWx0EGlKCnEUiaDlso4D0v/r108Oh6OD77PJtY5mJIFCq2SgKtt3BOOX/Do4a0aQfORN8Nq9APR1
CbwuzR4bA6edI0Rknffyxmazlkp3WmNfTvpvwn9/IfuMjzcHIdpQ8A0ZNjII6eDH1gTPhahbkxkl
onj+3xqvq+PPCwhFORRQVCTZ3gUwMarJvmvCyVT5QFp5IPRmcIoHxtZBUpSW3r8yDqJyMEDTyhWx
f526fvr8v4hEolYeyItFkaWymCfF6hpvrXbRKRvmkiTBcQPQ4mlABDpeYGY1Wt3kOyVT+7wCvzRJ
TY+MW0ynqh9Yp92690LBClr9WfNYqdMyuFgiF+qtv9ZoaJat6cIDMccXbkGxp0hlNpI30M2Oq7mi
MY5AnONEfuvV8sn2HZxdUJ0dPtMS/SMJvcQIZ79mTto/cSy7iz4KYHfvKkmdKzYwJUJ8TYYOHwbu
wSJIK27tdh0KKZpdxYvjEQPoUlk0n/rC+Xb5OVJviCnT5RfqND4bVwMBMsk8pRaH34XXQRU8pjrK
m5pgYEC8Iz1V3kLCZ9iU4/mB9oF9/fZpR0TDW6zMbo7e1rYAkWKQS3VUfqosT7bLEccD6Ep4NOJL
azmEkYMHdL8hu+2kqd72+4GkCQOQHy9FSjRf3aerhHoYoIH5jl1J96cSpDWnj2kdLH2FALUvbx63
CBFP9VL5qZBbR9yCtvRzHaSw0yJWQS1/7Uge8bePl7/mziYlePyNO8zc37DEop1u1OIN1wY5WGZJ
nVAeekGD8Dczf7HeFW+ZH/WrHyvIRzkj9Mdpf9+OmEXbb7TcwUKsEzgCJ3DXX05zglFCS2Ot40/V
3f91NF8BX9gPk2emUnCEsyWUwLm9W8H0D2P0tuvL9jIjX2gOrF1+DYMKx6j1LZFJmvNTKG7VMeYJ
lCqYfb7ITUMmKqxKqVMsdlI+2mIdx8x3VOyl0MyPke49xxRNeziMqWbalaIups9qL1zYrAZam/0z
DMr9y/9lDZL9UeEqPixrh/aLH8e8QJBL1K4gdotVuW7XPFTBAieOwAJ4tLWUNIjZ+svDHK/ylIFi
9sZqhqbhAuF7rJSLZbdyUwfBBRt9qCrpENc17dZV3+HVp2rR1o2RaCeIJs+mIZR8K+XDt+HnIZJY
lhQ7kmIHXKmFNmidautn9JSsjxm+/LSK8xr6T1YABD2uiEmefiOCQRVjyxApq4rgjNFrh6hsL08O
jbayxTuI9+fJtKg2OHOv/uh86vTZgXBzzkYKzFvwrrYNGfHSYBUSIme8Dw6gRPAqXkkFz9wOZO5k
P5nkkBE6+gH2Sc2ER0hTIxfM36dHFlu1xyKTW/t5LQYP/7TQONWjcX9LjO083ZB4Kopp9hLr4Ux2
x03kznPImfhg/1onD6wG3Votxpwu8yi22CFqyPSdUpsHVivcUeVt6e4zg5PNrKGbYmVcMN2HUtJu
HLJrT8SCFrcK4v+P/0K3lIfeLA9+NgWDW6T8N6fdQxGeaM2xh3TPN1glXE5g0rrba8jIsrWiwDPM
a3Nt0v1C8YC7Ir0+BF9Ri5mOXQmCvPP7+/2CvLaD5RIdmuLcV8afGHpfKc95nQ7TrwXtOT546fW5
1KJkUqUdCVaG+j4QX8kLe26c6+nG+0hsR32i6jwHX6DMITXEPnxQALU//EiI9buPMZPZ7win05p5
ERmlbKHyfBLdzxyvnax/eWaZacnz2QhLm0KTL0TdgGkfbVmyPKU2mS1O6UAVKLYPwQtF9254v3fb
LNXaQEV5oMOT5o1vkwqDKJh7f2dXeiG1KgnfKvrszq/Ean3+8/bYH5pYHZPgC3iGJyV2fNrzLE5n
GWM2xEQuIJHTzwF+1qrhq4ohGDJKDWL9kRm35K+J5BUSqKGMqIvOH8nKhl9j/fLmebUK1UzJeE/l
lCjmWKayZ6O+8GyrKyk1CmCoEfIJFHw7CcId4yc7AHzKWzRGiM7RPGOgCD+qj3PIkovhKa4FpoQ1
PABql0SMALHfOGkD9iYXtrIJyrKdt13uev+hO9o4LorVI+y5W8k2tiP6AtmZfzPGZC0qzQZr/Gm5
jQg4XVIIhboZJ/yqp2iL1l6A2O44QoEgG6ESqwLy1vd9UbVxNr+JGthzls1JiiI3BdY+Kq1AFxQQ
2vTgWHGkSZq2+br93RxB0SzTiEoEw+AAVS9u/EL4G6/YgcAIPmXlWiiIwcHkX27vjynJvwFUji8k
x2FzPoaAW+TuYWubwRho/2m3GYmAP/9sT65I7W04YcLk1S2Rs3MzenbQMdRlu7PpKy1YRPhw5M2L
H77FDD9YRIrh376uPegBFtw8YfVpRAiMih3WhnSxcckB7o1KmfUstoHcEewe+zDqxKvO0obz72om
irqGG2sDyAZXFig89LYufBfbRfdDwgm9kiffvOlo1AZtivYarTdF6YvPeqVeG8i9c2A8a39ld2vK
yfUgZNWQYs47RqwEKju/+LpfvKfl8OVDHVlwZdIyosTq+22+RqUS1DvuWK/katol/qBbFMk31LNZ
mo1Ds47EEC24Uy19fujihWVxaFQSSMugfwdNYpns/VL83nnY1GfjU3jrWhBkWkWXQanxvAOgkyIs
d4BdCQ5d9KuI61WA4edCKAc7cHL1SOFebU6S2w64zVh6n6qsiD+L2f+bkUWjX/0BVpgQA6Rx1woP
bkNBiJOzBnw/INOjZFagNZIYiXB1YpO06yQYzWSdH6SLpqb1g74MilcQwnP/eEqq/PDlYSSdT2DR
20bs1IyE0pjua0R930J7RcBp8Xco3SSSXSL+4XEqDkVoztR/ZnpYgebXiLexxqBwTnU/1uGBCiCK
/GQlKAXke51JQiVEvFYw8UjpO885JpbhnZ//UEIqxDWQ3tDJX+/T92YS8qn9PtjvSzvsu9jfrt7h
mLrnbeU5rSgTO270x4cuWjth2wjuKs3ItZ5EEEO8INKpYHSIDek6C/ClXrbpgGzoZltZaIHJEi2n
QlgTp9TpsHQKTidrTVie9v0lXxQRtmcRvkdkH8xgDwgsnjzombQkteA+LFnXzoxTBlpxStqBaRef
fzD9VonWIXtH5AZE1IF8am1h8Vj2HR2eDQg75S6TKlVYu4oGHIFYvh+bZoE4oXVSaXz6XlZRhKad
vyD50SdpfOlSdIz73hKJNheMX014pvZtLJB0+Zm3ApIojgcLMYeALT/BFa4XHM5f9UDAqlAdMdRI
G0giBOS+kuWlzbZJ/76JkE755t9lbA5pAWAGW6vrOAi+UnmzGpSZbszGc5ivsfP3L7HvEjT7pHzb
pDfbPKQdRePc8jnPQKhCFkJv6yzjjvynAvfZxdFUfIdl+bnX49tLmexEqFlxAmMbi0sG0O9wIhk3
e2mo40jQ0w7G8LIrknu/0u6mwbFD5fxWqIy3vFfpbursiDFnHOm2DbsSWfQ0VUodQnESSDwZRozz
qkGLEffwjc9c2kMCxn5XjyzaReMCPam8jLtEarBTktqwbJ7v5pXzIjK2ofMJ+x1vqkVVPA+SpExz
0JphOGPlQuTvEdBhW/Py8GLqinWxZFPEgV8l88jJ7wMFledvgS7dwGwgFLcVjTO3Qay2sFzlx4vy
0xUrLC7m63tH8uEbl7TQrW9YEq857xgmxjyd829osZJmKsskD5dW0rkDjoTfFqz6nD5Z4F3xCuUi
9ZNDFgAfSLK8K5MavX1GLaOTbdstnJe0LdNI2oNpIZg5Vt7quRDcuaLerVLZiS7q8uEri6Gmdg7f
8EzCt5VFC4H5+vaUyEZ9x2UnImDBcQOAPX0nZUpPYfxQfB8FP/+PvTYHX9vG3YMWo+RvwKRIato8
KSt0GpY8RdT3rEik5UOzfDWC8UMkmTUtT7octSfEpIloL+7LBa3WoZxA31XLfdOvNRXkE59Nd7Cj
/+X060AMH+jZ5/cZsigUVnuLiWUTZeBUc5YROOwqVTP70MT7uyHbJZK7GvvzllRdqEQbxT5H6lCm
6Q/fhBSJskDcqg6NCfumJq2HuRA0W7WnRyhStbWcS33AKSVWZ7aIY99RYYmlibDXzRhsH7B5YxWE
jSKCh3QWLMFhUZZMIP5fEVDvbb+KYcTCtB/lEvblPp8GWP7JnJKeeUCgRGNeMs87p+B+fBLKpJiR
+1kaEUrYqBZFARxN+SuWfjHVAxBNOvEoNdS1IutCOPz7XfvI/yuoTBdIyYyA8L5SjN8vKJPA5JkL
5Kz8rWWL3PxzHLfgRqp0nZ/1i1EY+tSvQMu9HjdY6M/s2PF133FlNnapPe+s0uDHIz8+G2O+HYtf
9N+mBBOIf4mgOrz3LvMpdgs+mxN25vD3nmM0ynYlHodENopFq8iijChrg/w5U22Pt1TxCzTk9nHk
3P2ghvaQGkKPwJhPe26XoYUdsxdX23G8HMW+DeLuMuo29Azf9DNGnQAL7588RrjrKnD8uyOlOkNA
mRLgZJpXfsztTqos/FIiHmzFcOZJe/qDA71js2kbShddLMB2MvqRJVhpqeTfOEMpUIDLnHk0oq3U
YPrYDqsJPKzEYdnp3j+yaaQA73UWsE5w0sIyay09uLR7RuSH8BKlE78IfR0/fRLmUtBAZlGoFEC3
x9RKVebyPwY7jlHN3xojOL6KZ6WpRVKLRkYUiwXZN+AFj676+bfdzAIqtTqk7G9FIgbn9pr4+/c3
hKYNox/h8qg84J/Yw+/OuM99qulZkvANxIkbTVZ/Ic9hPLQfBdfEQRikmt0+P9fAUf8kddvkPC4r
qoLHSIk7K6KFYNulnz8uiERalY4wsMZEna5e/ephkCpypCFyzUwCHeSBQib75t6E4CjBdcoDU2Ez
U6tZBIn9nLq+qec8HtvAzE4oD1x97f6LieaQ8yIG7KD+dmQ5EHVca+R7VikHzSQwC6QV6/HHOki5
E4KGnv1uXIxKgPs3X2KOp0X6gy+qGWd7zWZjtssXeWHNRGMjJhlIIg7AvP55mIdjhbWnRpdNyCE4
ch2Vc5GunX/Lqk0hagkC/R57j7qSV5DTj5fV/jVrn7ajc7Z5tnc+dQyB5UjnVIlFC8wjqNg2I/5l
1NAU0MuQQ1m//YUGU8iY8652GafGmCJN42cHXwojVLgfUhPuqZez/Q2+Yg2njyXeAzFnBbiG4zCM
Gj3/yoCnnwJe0cqmmIrQR3QTXSMKU2GwSyYHppCIE+9gXvQhjz2cU935NckY8PkOgn0+rDt2xDQV
sMqOP6c0ozTx9LT8Lq7ZRKiaHjSkgCbbI7y55cbq2yDYaQoRSKmftYJ8yzjdo4/2/zN4uoe9QmzF
hh+FXm99IAmvAp86E3Anh+1qW1q2uYCc23cqFk8ILr+tD+9XS9MGrXYRGwS0O6YO/eINkPSsnKP7
4GTimo40OGCRulWNMeqEamH0kkglx4H262SCXtvqVJ54QsvfYlgQMobw4FOnDHatUOGr+H5foqqD
StyE8CvpqO22ho65yHiF2c5OvaJzEjW5ur3TyaEZCz4sX5MQ2c3fS4BaoSIwoymqQut305m6FTit
NRqhr+MG/O7YLcKciW8OpdSUX0w20M5ylBN8T1ZKH7O4WK+B8Y21/1VR6BxgNJCy30XUU0MqYYZI
6W4SNzyVetoXbcS700VSXnNU1DXna+6IV/bU2IT6CLN3EdztPY/pJqev1qbWPrBI2Xx5QB2Ugspq
GkEfFQ22Wk45yAyqkyVeUEknsayvVhIS5n5/Nr08cQroJPMFgqeFQ7NppX4sl+ZsMOeu28yqk5ot
/8PRhPLuHaaGfrzkFWwCeZecrZ2dBobigSZb+bNIq/EaEsLJFFZlHScpO3iZNE3TCT/lS1JqkXWH
5yOpswS0IB+gAgsOadRnRhHLo5mNBl9DFIfaZUJMs6fUlsjQhSpB7HjhJScB1eCbhMPAVXUvVgm8
sRFZy7+M/DU1Voqp9LPyvap0yswt2zhrelYJZmh5BXGTEs5HU/rLgbXK4qpDcOMk2FIw79P95GLd
kbtLhXvi10lZxdyL4NkmLzaoz60CkGdQXIn438kB6+NwqiZc3IXFqa8UtaUneoEasjydlV+u9bt7
SRNfC06FfEgSTKvLkxCSb3rlPELwWgUb+60BoERLDuyY4UHRzfl3Z07tlGuifJQGk3yIpyepJZvK
V39DDpqS8WZyjAtrF62i5G2vv8OY30XICQHu9DxSGh2/GO+3muMLPVUQXqbbimctFMjrMgc0eNf/
idaJzPEtHixGRXzh2lkeMVLTYiUfAXmSPfIv08vzx7tCzokz+XJf33jzLE5EgfmHtFGO8kGKAmbq
uJZz4I8ne0Pw/dCRr7UhZVyvy/DiJYW093KZexzNjXPihTFbQLhKIDWEswzlMoClFk/IoZWAWahq
QzRWLB//2wxjbHeB8iaH2oCUmWgHkij/OPirqskUH062S07lE+osq2HBCc0xoOZii4nM06bb1eFv
qve5V64Vygt3zhqcRdCQkCoAjhDr8U3pwhCo/EoIWOhYDeYtm92o2Zw7GyPS/wptzEsar4brtA42
mZpdyfPsxuIoANUAbm5KXNNRQ4iKsmhQli9AVOLDxY15w+rO9v8BCYZpLuPY5PGAJ6eyxnwZuqR4
/KW64T7XnVRRjI/BVl2Pp4DuNZdeTmXAi3Bm9edIDiILZwWBXtShYAHFtOO2QSWLf+dP2Mhf9R79
LXo3hDLsatzO2o89lMpcCE+b5JawcwqttqZNp7GgC7bJy/XWCOSoCo6PhN6jwDZE0MK7p91SKBs+
T6PtJNXVHwV4am9kriFLpYRVwiBB4UOFd7Gw79cbL6eoszgM2erXUJ+tkqdgtPu+ibqs2zlZkbBj
F6qn6nvrT+b2v5XASj5bazF0sy8q6yQ96vrXL5kzGiSkCPXZEbpCf5pVxHk2sF8a0QVE83Mt/ggJ
2jGrEJCErSsnfaq7GjqB37t+ZQR4wiKt5J5ZhY8jHjrhw0wGrIwNm1KYTq+6F4VmlRPA7vylVH9j
bi/wdPK7YNu+jwUtVwWUqCPu8tgaQWicWCEJElOKf5fZURfSazpXBk1jRSPgGjRvQPFKdeJBgPgE
fGm4vGwMw65Wm+sGI5/fsBdX4KVOT82fbg6UmHlY9olzdqkhricf25xTsQDyCLItc18MK18y1k2C
Qkz0TV9tv2CcaPcJA2gmS2opsIciZj76iJF4V+KNwMKUVdhZN1rXOMcd8V9YccQDPvDl+57qK1dv
KaP5560g6cltlWS6VYglJV7m8638Dfz4zdZOnsS+tZz5Xsyf9ya8zgHeGmYEuDS/vwhnVDjpKQ/6
ZGzN65ShGKQVOrEyEsr4UD0YEKhuQtZZyDWRnBU+6i2TANM8ax+4IkIjMpLeXuk5+7sxp28HZ+M0
2BibrHAmbAl9GImRHpTzHyu7Jket340iMein47X7S58sV8AvPDMU092z4VneYuQGukZKjXWFsFmZ
nN6xeH9sf4dfMhNkjV8L43t3crUuOQ+IoPI9K2xrJcZhzJrbsZktA0jY68WKePdzO6OstdGWVmqj
6OdhU4LcUvO5hAHDb3F0kG2SzDP8YXjWg3QLwwWaz/o8wR0WOrd1Y3TAqq/hczp+UYVzDXNJRB0e
iIKPuZkXnDDTIwAJvqHfMRXuA83LxSt5EV1wPDc3lhnIaGBylcijoXeCGURQu93iNIweuWNWRhbs
Miil9qPT5ZTzup01O8xkh4Vu6oK7tYPm2YRvCL2s1S/S7Se/WOx0HXWGhVLQVKisbrqFy9aWL4ro
p0vvQ05+GfCSetLtp05KyjFxVUeVY71DM3nWfQOZzIetHu50HfP7FAPj994yZmQ5PQ9BmECgVox3
BhNoMrLY65u9MJJ90SlMgd+BjSgR/EpxHchYZpGcDBHVGpZVmiQ/exJgli4s7h5xJJDZuixCltiq
pLGyXkOjaJN/08HqztNREmcgACs91sNuLnbN/o8hEA4to8P/d4vrudo/Pw9OmuttLTc5lReU4n4N
e/abylKvK5oVL6Vqeq70Kp8aUgS7jFXF7kxoQIuBVpzNsyMgYuf37QC1cgMeWbRyAcddXO7cJxSd
oGWt8PNDwBuaMXlO/3FRZ+hCHdy2PEjh/l7aRcS8JYVQJWVmaXVRZEcvwFflTG4JJWrJXwdPY3se
YOffTx3UROgOrdtPZ9X3BQ8EnDmNbWzCakN7cIhRAsESiZO/RYnbhIbb+ECmrC94redYnqTsKGEF
A/3Yyn91VaTV03VixfJu6uF9ETx+jp5SlsT3RgKO6QIzsCXE1TIW6yTbYbWygWgcyCBtfdNYAo0p
gd3aOKaAjwL37HqagQrcS2JzgTu4N7f8YBlR3lspFNGRFCMo7HJ2fj859+qLmOQy/RBzo5J29M+1
BSABcEbkuUG7uACRaLNvnozTgbD12KTbC2A3olrOKnVxyOO0bBfNelU0TnRMvepZMmdRJV9taRzN
Ex9EEMpNYgDDrLom8IXhfRZ78G9wjAaoSAgxIucSCd7n6Gd4Rfm7lMEsTpnti41+43Kpy5upyNfS
fnQIRxGZqTa/dK67G3extgAbD1XLneiZUHQnEUyUlh35UQTZAGwPSxxo1nrx3/dpwmgZgS6oiigI
Nkz945KxDHk5unTVEH1lyrMMjIz91MshIwTCV38zMGivyY+2TZ9A6pXb9YvOfGV/T/Qh2ji78hJ1
uKL9oRkXZuUkw+MHOkTQWw0eprI/EEABQ+ymsjkBC9ovEIW7xEBhy0CHGYzyqgMMntmi4apnfAXl
9TbbZM+Lv49c2uTvQwfdag/Zk+2fOY0Hx4PpXS8idXeLhl3X/wP8RB511wHSp5eRicjZGoJhbXG4
93K0pQ5jVfRVbSDYP1tPqjHCSbqlVXyKLyHPLjRx6GcX97QrVyAFbUi7lVm7wLBP77Tgh2dpNt5i
v5AqCgqNFSdbhrOPhyQFDtFDETyATsZQPhfImwXtPyjEB1PrwT+Bd69eY9agbmxe2P+wBLpkTxOY
xfl1swE2Gyd+sQtCHah6c+QtSNjGRoMrOP+joMGhrWdc7Zmpw64rOXxe+5kGbvhUv8BfIQCjdY34
yLsZVOo1u6r3wb4q1U/XJRyGMporpyL/uUuB72apFCkctRQR9/9DL0YjdMjMUDwASZx6aoWqSD+I
EOoRnWtwyGfJ53Ij74ZJXDPtPsnkB+knXQSXJLLO3VpWivZ27wUabWBtuxo9kCY3tyjBnABmxe6v
qE/c6cVjj+71wSc0dd0bRnsjacmNJtmYNDLZSBhPK17P2qRFHs+dDZpKr6WX67NV3o9uBFUeMH2Y
UdjNf/3hw1uCZfLtk+gyVfZ5/aoSFB0hcVFCL4YTdFC0s4hbXtU2VTb/EXNtJjY78TnypjiCUrlw
FxVlIPXSvjH9E0EQ97IOgcfWtLEet2h4pramvwtTc1ElA21Q2t5aQ6z8nw0DHKe/YhPwn/iEm8OV
q9n5Wxywis15z75AzxR9Daj16WaFySgl4ZJ+VTdsUV6PyN/ElrYvIun5zOzB4bZIQuHoY1K8446w
nIqnF7UJTlN7cnjhDjDB6VH9UCgf6TlsD4CEHKadHm23lRhh0vWZCgny3xNVK5DEBtoaCc9cgoD5
p9qR3H/GeMPRVzqPp1X00LRBOa+nQQFjmp05aZ7V8j0R4629rG6lCZZgXbd3it8oSGNDyrq6P3UD
7Qu9MAV3sxS23pHqJSwUoCqrud93OOzg1DedTWyXC2KEB2Ktp/jEYscq3GmU+mPkWoxxnHP22CXV
jg5ngF5s5PohiNLrSbI7g8d2wjNZG1Y50YWbkTPyUXNaqVUDEjsSW7RHpm3Hu1K0IbkLQGihHTol
5KogfpefmQYYkhLWEe6fYcgism8pRzbmgMLkvvwn3OnIJKQXfJ8xBMHlZZ81OFf8xXgCKIkf+/x/
EljOejqdsCR+gFG6WwuuAcyLeQ/VcMea3cFO+md3l31X4W0LjJkEgb6i1GFalNWnpvxREMo7TLGh
giEhCCXeBF4Q0R48BzIdDD0G0g7bBji28Jmq5onpDje7NOYrg096YdYrmfdRVyHcN6YAX+qROLuL
D+25PIZccIx9X8WYJCppoJasssSUy1EwpixMq95NPXxUr3Qn/en1XAC5J1Bgbb1NNWfJ4CE3STBa
sGmrKT+TwWGe4ibyxy24DYgUMGrA9+i1YvxT87p6nzi+8rYAw7ucfF/Q9aqqLPBaDfyLRGYgXj06
tt8baDWq7IfKbXaTr6X/83NVh7A76HaDIPnrMDzkJLSYZ9TGWyAScgRj5uBKQfyOarusEY9DxTR+
8ZFBgDSVVK1wtxO56HxdSLnls+qWqd6FL9e5Z63+hNykMokjMuHaj1PBf2A55q3nEhfaAjiS4eql
UC9wzxTbMDATnm9ky1UCSpprVEMCCvEtZP1qInDq973YTXw7w33/PJbgY7X9jheRshIlIPtPXbeI
kaZio2pEd7PkHRxRlZH0P2bNAPsaH6G3h8tAN5P9ilhuJkSeL9zxdDgirC/rgji59fVW9I6xWEWh
tX5nNDMGCmMQloUTc1ZaYCISvkGreMppy0XL/3wjEWuNCN6hsMxVfodfvmYooWXuz2irXsv22yQE
zz2fvqYinI2acLS2rKPmQmUSs1fky7pxb+xcRCE+IFx/zrRidqdcLqUAiPCNDRxUonM0xdTtgcs5
+pnDqPYkMDCcpobUtgpJ/TkFvvXYn5yHYqbeTu2xgvGfEjx7gkgCLQmBHBJxLxl7Y0BCIf4k6PPy
xOhUMaCn9ULTe1XGo8N0gnjFmWO5zzDe4VBjmdBWDPzlTTXTur3Cn6zpdBbPxaP+b7CJeC/8ZEd0
5OlIWpwGZ8eJ4nEmgqf9DooZ/e2FSpYJM+pz5RW60YWdSwNs3GW7PMQ7G30HjDH1J/XB3qc6EoRr
7btW9urahlQXgpHh1SX7qjfzxBc6mE2xFSEK9EvA2yCCqXXnwXtkUKxuVhLDGjo1qjFr35FfMapC
+vE+7Q2uel1vQ16IVPe6aYTz23M8CFfpCi6wv9iBMSp6MIzH/1NvfZIXatpmtHKYJWFH+zJ6AJY9
TSXY0PA5jcT2/XSt51PeLqjtdC9tICsnMXdd7Gdqg1qakjOPIB4DJygiXhj90TWT5UQTwpweVHKJ
F4eKXIeElxUmZr/dvpYRxnBaeycLn6N64nW0iSf45quKqtp3K9skM8c0s1v+jDUn1h+y/vrvyFVo
TYXp4xtTVK/7TkD+z3/eMzw8rSr3viMRFgBPngQYuxzlcM0XS+jFVymIm/IGNYx4HLDOihTsFjQs
b3YP5UUFdab+Vnv4THD9vTRtoT6woXdlvL0L75EGY8QNhjwMskL2xQBHEkl5KYC0Qo9RdbVx8prR
PiUgs4mk8U2pmZOGlIWCmt9Sv85ue3Iem7jkRoxuvezK1VKO6gNz7wtjRfJKNOgB9Y1TO5hNHXle
Ep+c04hBNmFiRaNQMxRF5+AQGzXd/hHuvnI/aLznP5InnbxuoIJpGhzgdwVpVI/0BZnkQ52NxqNL
KTTpptqB3rn/b7yNx0FwnBjuZi9LNX2EGGeoUpaZUtCklK2sd5vFErkn7bOaqnokjRQUzkxLGCpe
NMdzakYxYrNFD32T9haI79zLxX9PBDRSttd0BTww3kgDh5unBZ4rgi9SRd1K3kPn2Kk15cXz9cHD
zDE+rrPyzxlHG+iImtx9PKdO4daCEtOfg5/6r2YULvNoJ61s3JFO4ZbW0lEDUneDjlfyrcmIm45c
Y8ho8Usrxd4bZW+40e3Q5WaF8v+xQhbQ6bQ3lFEovksGaBWQAy2YjEb3cRDoOryZFCziGsC6mv1W
KUXMMCndjMMPdCDO2BNE18Y+RWxTOXBfDs919rARy9rlsEnh9ERZ3Se8WFQSdbSGki6yUH8J0qH6
Jj3j6qNwje772CZqXNAnDW/Z1tJ5SBe7cpIeHeJYjcfVQ65CmQSnhXuuj8mlTF3gEzI7ykXvPWbJ
ckEnWDl860+K1AX1SE+b10S0gGWz7FFTC67nbTbhhqzxSjUhV9EbzlaiUF9vxs1y+p9vla9f2uiS
fzaoB88E5hs8111GvffgNkwSpLwA+wFp2cXpvJGdFvnRdzknGM4ijXZ6ylp3AzzMNMYhPlXegQdV
A0UJM8QFATU6z3Y5HfR9+eM3X5AOYCExdWXwdkrf0jEaDnTBJ1YrNbF04T+p+yTHGEfENmiIvFZE
0Fn4RC9KnbcNbaob3rXUn4byBUWVkLN18FCYoMPdzJuc2fsWFlFHnQsUMP/wEgfyaOKgpBIr8vva
rteiUORX5+YXY6kwbo0s15RxzCxXJQ7INiWmSWbzPLLzRziZQi311r6vL4vYvtosoKAtjh1+gGKh
frH814KsYNT/bz08t7vWmE/AqaxBQMNCYQ9Tz3b93kljoq+Ei5QUbwiYVsY4IvBIkXyAXEkfoYIA
Foe5YEVY+DQGHthKoTVwsupyj110VxHChnQs2YwTxtZKiGTbWA1hHevMl+/DItIZp6CEhi2IEne4
UjV9y6vnqBNPMq2Nc7St1MGU5R61x1wuqZwIMUdxhydE3cEqrV9NzDEzUx8iG3Gbw2wVLnJ3ag4L
ryL8rCGy4OUKpi2kEkED1yqS8wyYvlhuCLPnFNAB7YbCQe3KHmm6Tn7CoaBFLICbgRsrSWoYVpqQ
CTAah2CuI/pj3V0ch17sY0IxvPmXvnQM1Bj3b/cvrNXqnJ8oUwR6k32uFN6hsDFfZsiXSUlga/K2
MoruPWBuU5lJtsZhbY2/5r6N7LCRJ2h9/gkyd6wtUlA8MY0Dye1uZR3oSMlReso4qJA9QMi/8ziJ
kzSuo9nieaOk5cHwubqApMPUHxlzN16ntzJAopt9IznohLPMoKKVEZACMw5GHPtA3xNsg/tEcslx
cr6rwnZ95NWvZ2r3AAdKzbt4Obn/DCETFpmpi2QgGTm0vsyPisSsjkuNLTy6GREtt8PeIM3znDaS
mvW5RfDsggzbQw8pFTwhm66pA4xWDDnJMdmU/LzoPvgEomv7KQxS3CmgaelyeHzfEwg/WE1Xt+or
vXyoGIjMR7fo9UGycMs08QIlNzfTyP/uU7Hn3kJyZN/UdWpycCEkEfPLVXZnSpLwEKZqWAxcQZOn
DaFArcJdIyvM326mgwMAs/o9YrZ+d/OvHi+Erzic3D8oIQdsgQvnsyrJ5klHSkB4GdpjMSOg37rz
I93EPrZdzb34Zl19UvqbYWU4IIMr+NEXOc0IN7ThlmR81RPSHhMaySXVWJp0DakVWOTTMi8vuC0Q
Cd4GIYJ5rkdgpTm7kP7LQvrveD83qnSehLMPthVHBncBzRUv00YMu6E6Qx+GvmTmamCOSYeZgHuy
TvSExItTJiNiLRhc0Myuod44gzrNE0NcGw9sDnJ46lBjl23zxPxqCjRQe+NL1WB86dPRNwEM4nIr
hZmbWTcziMHjd+iJKNs+ShGZmeWiYTTfh+cmPzHyFW2lBZAemWcxn3qWWiyDIU46FBdBTga8yQt4
lKIv0gLuvaXpatP2goUPxEhciK1gkT+XjNrp3DfQVS/PxrPKcJtaGK6PXkyX8swmQeVxJ9Lm5N+2
MD4h1U87B+0mmytyaO+oq7QPpa26H7syqDljbwynIhR8AVkQaR7m0Rj9y2w2OfYlnR39wjn6vMZi
T4Vf7nXZ8THwrL8t6Bw6NE/2lBQIImAUfl7O0IF1AQk8FJ05wxbHdMybcXXEHc3Y79WMEMD5YIOF
ZuwukpGaWA2HnJi7wTq5KoK96buVe4CRyMYBnSMhlJfGUvgDdNmFxiXT75JAVdYtjlzT+EUOxjoP
3do8O46hUfvsK1LpV5sGbd4ijjFc6IVPWKPdRQmSPD4s5e/q4RNoYPMuMxyTKH2WGZ4tSRZyJJiJ
Y1SZycfEctQ+P6BLkcLkub+5RaU0WK9GaeL741ztco0vHglVSoWOUnI+g2b9xWnUYPD6/Qxzaxx9
l/6xFsSC6JWSuxPu9LR644rtaEztcdWGeoxVE9xY326eHH82e7oUNIZxYnvvBYdaYQGTp5/7MkdJ
udt5vuxMnMheYmL4F/vWrW4V19skUXAIPJiTzjD8DdeLBvquUGhhw5ePkpeY1lD4lIkI4wifnTjh
jBn61Q8BZ7jyVUeLjTBfsUF6IofzZ1EE/JMhwknwfwwehhNtdkhLfsS1GbeCP5SBdwL36SicOnRm
v3fclc4VOcSpue5KvoOAd+J7t/r5nH165E807P+qw8guf10M4Dmfl1V86SvYHCB+7yDRxPspr4yi
oipnduaKijn4eG2/m6wNiy+39f9ffTvnXoZoq2DIqLQEX9/fJvjYTfHNGcUorBOES8SeKf4Hbx+Q
s7r0yMD5Ls8kiZjs1ml/yOo0ow2HhCkwTTYHm/wtKn4TqtSjDIekalsLjM6S9h9fNNBdVYGjd2wq
CG66Nx7yCruFMPSkm7dGiVxS5rIEyJ1qGESNs8Uc6NfCUDqrtFdar9w/vPW6/8ouMdmuZAmBFRgo
H3zm+ssloLmRxFmbgByypXBn00XKW6pMHDgVdZVr21EpUlrDXNBd/cGAz5zfY74bb+vkTMAjmOb7
BuHLGK3ZK0RI9qUfT6fDZsMDHZYXWFCeTO/WKg5C60/BzRbKbS/bViB3fxVCOcsKpOBwV1d8fKem
a25yrZBbRHirkwpW883Zv32JprljhRJDKk+rq/9/LcaZ8hoYWYdZNFxqk4EU8y4zDgrLfGPcaHcV
ys/ohX6OekD62qndnfJONeyVARpVhmFG6EdRwikke/pZJXsfT52qredYbzS1qhUQdN1d+w/CwJnS
4r17pZQvogiA5xgRUqeuIMyYgqY9LqvIl697bri7jiJziE4ecXAjAsqcLcF1GjMU+LdBFrzkmgiS
LUqBzXK98dsR6ToeJyR9FrYI+cBQpDPOvQSUGRE6Or/ZHxObfV7I535kxp7ur5nqSi6d8VCUozH6
CjQXZJPXypoVJM6fwrT87e99xS8mkM1LLo+Jb7PwBylKaWg4Ac+SjjXq6/teTDN5GgiE5gjkuvAh
m8Cwa5ajPZQYN6cu4x8eBm1dfDNFYu/V3RnaNhjufPbMAWHtvYjapgCLH5JNpDcCjdzeQn8o/gtp
vPKvOK2TlnTz1QKEMjyZgGYazEjQ33jAPawhC0rdJc0mJRIAGA+1T28SSrDU0Uz/YhGFythE9gpD
LewNR6YEdwIut703bR062XJq3MpLCYUh4NrcbmeLCGBPb6v0r/uznL1ZUCfDH1yMgfDWIkpNOP3D
PKamP2AtMM0gacWoMFS5bZWGJC1iElMqmVw8MQQI7VTw1j0r8fmlIETmzRdjI8T3YkpcyrTOG4eB
rf0tcN3Y3fsjwvZLNk3AweKfV0bTGNecT/pVlzh/q0rGSCbKZuLGgvSdhpgKEjFDYBfyBSU5ONbT
3cgQXaUPa/PK9YGUKZ3M7OskwSQS3QTaq1ghSDhIeOS3pGX0EX8VDhtgJRRblH1ONGF02mkch/xX
KOt4r3LA8t5sT3/AaJbz9e37LmAN3xNLb1X1PdLY1qvjEGtA46X54RL6ZmuPICY35X6yZvCdnNQo
m8DhZBRIJYzaHNXQyDfp1cvk8AZjL3bcfwmjRjA/C+k6Xvr7nFghnYNQRYFXvl10c+vzy56ZZZsi
n8SjKCczs7OQ9MkQE0s152UktN95fiqRQrkeVeeFZ2gXCG5CDM36MY41qJ0ELaFCUL8N1nWSa8Yj
ta47XPXFI6WYBUUvkjM+jCyXinTnIbetdW/Grh2Z06d9V+JVxx302OXgxAg7yH0KNLHmuKSGc+pR
FCVXlaM2wSOupM+aWJjimkZo6BfOm2xT5/UjonZCayvzDI93ipUowRbHF+h0/LN4lmsCTMayYcWG
DfxNAB0SMEtVByqQcocgC5JrTkMjUjRgNNzgFpcQT2mFhqd9oO976zcLJ5Rgr2IbQW+r8xtrqBRM
79/ChQiuy30SC/s86wkm84hYsArLCDlMBR8wgalbtEkYQVlqn+shLY5rUepjI8itWqJ2ZtNQE0DS
fy4B17PikEZvJ24Ss+GQBeLkfQNDx09T+YZqc4jLdCVR3uI1ExgNe9Z4RPCndQw7Yql9Tsj4/yus
mLz17bHgvxBfGJjgaVU3MA0NzHgVmXy7c1W8dHrIeCJvU1jYJaxZlR9ysPZZdnNjJjJMsQCd4Gxx
vAhZFLI6G/oTMkGLf7XgDGwF2EsQBrQDAm8L+ozHj65VgkNbL1eqBRQl483niksrtdY0uxXFmZ2z
GRGZKaBiqRNeU1ySKKRSu6DcaSBCqlRcwueBoZbNwIb61fc0lVPbxxNV1gJuQajvVYKylX29Huan
gh8R1y1e9GrhwnVS+f3SKgG5iEpZMprA3lQ0ek95AYGcYew8aaZrCcEt+VwqiK5mbLZu6MqSaYYb
8vL3ko/GGbZ+f4aGXOLhl1gNpLPG09l7S5bFwR8mPxSFrglPEz774xPLew5uQ53dfYR0xRElVYvn
GQyynX+t0Wa1Cw0+Malu0VpLrSTBoY8HiHExfRVsTgDnTc8peQTIB7iyB7zk5h96tkcBW5bR3jjR
RScicuXgvIhh3nLVWkESPycLhxV3ZOj6OJLnqC6t+SgDa3O1TYZpe7zuZba5vcl3ZgQytR2f57wX
OSfFEs3TR99LovGM2IhpOjk73r1cc08cIoOe7PgB7TJWlmVmYwQ98SmhrXaEtUUuo9cuMT8peYId
ur7F0eWDpXQPhTg5VFTiPdCK2boYQQsyi24fdkZauKwpoaFlnCBhn+8HXfggBmj4dhsHkVJPlibq
4K+KcWpknhnJwVkPvB1PjEHKIfgwBJW7IutaEwYPioOIr35oAEN3479wjAlXl+w4/oRY6kxHbQ8B
1h2/cFJJOpafgWUploEnUsbQZpokp/ruYjAt/9Yv3YwPkff3xG3TTKilloXl5kf2LtH9uXZ8fIkH
SYl0nP8xAqLeTkSt5M5ngbP/i3ZniWEPWEtVXCOw1F9jJJ+dHG0c8C5Q46uA3medaPJHyLDUJwNu
oyfbVmLA/I8Rdh/J8sVAAY7ddDwP5UwzijzGeo8bZoGd4PA2ZEwrVnclH/lPp1B/7O/8npHIs9n1
kIoQlVCz2suHj4nyGbdQXbRPHzjg7QswCbevFW7eHnhqxcN2b0IXslk76nSzVSolxh2uQdcTvQQw
e2+U9eNqL2igVVOkQQqy+c2MzSN3YwbG0ChAVgyKiXop4G6GLggvjBgtl7TVVCmrbH+r85HYworS
/dRtdYN9mLoxrquZeiztQTkYjMn1HLhYUzE4sWuQzCyBx2Z1/LIzUvwvM1U8ZBo/qdtf52Nx7pZ3
En9rVfKn09QXyAxe3tXVaPzFVVwwOosjsXTfTG8GjX5VV+nsd5OJ+pk+ujMtuj4K9fola8Jn+nyW
F86lj2QKwbsIidH2t5eb+1du16QUirPTkhFMXdfk89orIqAfr3n7EMwwmzCj67VPuHCqiA+r/5rp
R0NSq3OzYySe4Z4y1mijRZQddjwTXrQCnKn9nCTem683ua/B8NBV084hkZeNU2WXCPZip7w8B3Tq
OiqT61Dmaoayby8W61vTMyjIkZJzrpadBrKYpPmcMHvNEZqCnWwy3T7Zp2kw6rCXNfPrMjLzm6ay
o40GsODD2MkrNK8w66NvhLa+zlgZlijitTFSUE2e4V9DtLdp0nVvHNV6ARuKM6L9k95nVb95xUR/
rifxkVLDuTN3OhWTdE4N7iFIYazP+7wuf/1a5i69wENeTzmkWEv+T1+TxatvXCkBwwUuyHkQWXvL
6r1KYXx8YzckLdAB5RnR5qdV/cNT9dLQAPr2KxL5JXaEkA45uwW5yUNz2xspm2MSFqqcvzdcn40o
cLyrdcYcKQ8F8V5JyyzLirQSz+Hm1mldkeZuPje8hmZ4IfGHqf/uhKLf9BHk6zK9vTIozx6OPl/G
FgjA44ZwH8et64a6nNsaXPQR/l0Qa2CxLb6IM1sUSttoPlds0IbQ8iAVpXbLrY8dU2ZHZjtKh48C
YFUkEXP9G0Eaxv4JNQceJnvzZ2HNZnnQI8yhuz1SxZMYPrnPUPr+hgv7+aKXDtRDMzOTn57E40Km
e2MwO17guphRHpHJeEKkGcHTU0X6+IqbMZZc+bpTzbUK2KAHwfnCHFYjwbZPGq1WDnhb614J9Eql
RhmiutK0CKk1Qz5mLDJDcnRgL072UoIvD+Piv5QxecT21+Tl1Dbn7Pq+U0btGmQi9K6BRPPfbzXm
HqK3PdAK24jvKbJz1Yc/RAn2X+ZDG6xPACohscqZKga/+zspcVx/fyJFrqvS4qDdE4v8xVnjF7M2
fgAZ+S0D4/eYHVCQkmHanNlFJsewUFiF8Zeu5bllf8z9w9QXAy6zKUVz19bSOzmX5FdoUHE/4sBT
Fhj+eliUEPxeTvCGFIRrYMRM6VrDL+eVzPYly6mNqQRHB8jQjPQhkDbDt7iHSbCMhzCwMx+IauYD
xW0El06/la2tC2jW0sNegisI0uS6Y9Ixy2ZGqwNQK8ur2RCj1/sugvP3O9LDLQ02jox7K9+B38eG
PaBpkx5r3fYbb1jfKhuqpgajitGVlp6ruT1Uu5qPEwPT6vMk0BbET+v0CHVO/cTMo46lbkUN47uL
L8wI3c5kU2GG9gJFxozpwxgclnBo0xlZZtzRHKs9jWxg5g1oilUOfwR3VmdOOBA4Eg94dfWfJTa/
gxUMXAmv9taLEhTbI8toJFhWE512JYS1ZTnY8H2m+ofpnpU8uki+opEz6LiOk6BTBp7jk7n9zE8B
8d/KxYMOFy1pgh7/2M8tvNmpghH57t+X6TS4hD9MXEcch9rtphNMkL89TbzkbuOZcevrKX2BREgQ
/XO70XMR2PBWeym12cIZ3GDPl795Ozp+dfpl60Ji6PaAZakYnSRBgPMYWNL+OISnOenerPV147pz
OoqRn94ABmOFX8tYT3PLuaGY3g+Gptuj4XJBt+uSUeHDsPj+HEV6zNSu0YT6MvTwVsf9iZC8wDuR
YlKfjGi2pUULbHpdVS9gMMIpKCYshdocYTWtEUJZy2ObBh4TfuT0w5QzK2halFyWdMPRiQ2l6oNE
fCHZl3fFlfxIEvsvM0kOraeuj4l+7T9JB+610o0lAlut2x+DC54AoVWtjBfTbC5vkSi6SK+jpQ1e
Yu7nVUDcwhjVQ80bimzqUGUGaO5cyCHk+vrLu2iU2QP+JyPxRma6jSC4b9QknxGf5mcKmbi83hKR
Fh1+4o021v5yGNuBqMzQWgnRt+RuEKrPr3fetHG1eF/hpcVYCmFFImnkxnkebTnekB6g/DTGVNmP
Si5fMOAQqP2jzkmP8yjJ01fPt73C8oUVkd87jpLBh1Fsn3vGV/TvgXWDc4rB6ISQFosfsfl12hLm
TlAbaq0Jnx/aqAipy35rWfFEWmMN3XrGIYlBVXf4lYpsffxAfYQIqYFYesFgOt94yC0o/zN7kvol
BW7N6ahGk2suQroNBQuihVlwPsVfhdPRlLhQ73X4hVfbk9NX2qdOZOHDbT//BEKJNRsto7xgHW5P
fZ3l11kLhuJmD46HUJCOxlz63gunBiTBQFE5udiFUNwdJgycsOBXek5Y/H2Kow2AiqS6LsgZwMb1
HoSOAL5rqdv4JIkSFqq7hTT/co2IrG1SSuEiTqw5SACnsVSkEgdNnnNfLcH2cyaHRLxqfb7rM7cu
uoBhkm61cDsrS0AGlj5jaJPcLgZWplmvEWStJvDVnOr0jpOkH1qIIJ5C6EubfsxllW7T8jROSLM6
TMEOz8ChaX/wqr06Kn1RxgXtFkedRltrSq4XzODaZGR+V5rLe5Uj8r3p4h/LxoohNSnQL8TbL62y
2DxB8ZvpMyk4rH+O4TjrQxSvfwO0JWkNSEWl1prhafHytTJ9hB9FOH8WTcKBPtQJJqVW0kMhLIIw
FoOiJg60MoRfuyOhd36utm8DcgMYH04yDfCCy5wFa82d4CNIJ5H85XO2ILVLR0QZ9NjTVsCfXWxo
M5cJdQnv1cXnY+JbbObodM5f3N2ct/px6pq1iGeREa/osotPoPnmpG+SYOZ9O/4kFlWmgLW/tYae
+sRsXPz3LjtpvLRDVNnfpdgoWCOu5TaXCOjzElzHbr/SwCv3Za3DV2AQETlYoVKs6XJsdGr8uXj6
7C7KfoVIvMmjPQb66y5k1XwrIM8xPtIiNqp/1B66cRdaUTZR/Hb0A6fXanYY26C0eITHJXqTgC2S
zHkpz75urnrgW/et1y8aVAurzeflng0mXR1/7x8Z4VdhwSpGJd6bHpqHYx5pmkOhU8NmePESY1xM
jPcT4sNcoOX1sGFFgVvxXgozHiLclw61NoZoasvUkPbLvGgr3uwuok0Osg6jv71FxO6RjFMSxlIA
EBM0rrRvTrJ9RK3P9E3L9FG774Mx7+c/Ae+Ri7LmRlzeKuoOCIftnPq18TpPTVayidMLw9APUISC
UJ7eyEkEmMw3yV3HAe1icJ6f8EzDvAPJCPaGPKpE4MvkGmbkYILPHtx+kHQfnUEcKsK20+B+f1dG
1xaJpZAYYZw513qS7NXbCKmiIi2wNpsnKApwidbT4K2hrLKhbnNghXUsS9oDlRXx3zstghC2FNTg
J/vC0Tm0Uga+ugH0+igRmLUsUykQrUVsFV9Xp920Q4KZ0i7bAhnrKxERfls2F9cJ33LMU78pTuh3
1+60r1qTzl00VLlNfU+KzXoO3shfupGQJHtGTeapc+YONNqwRdC7+AKTz4JsyESBGH/+KpSnAw3U
BTX4KRcqLjTRIPfL9ftOwN/FHmCfzUWfQVzBpz+nV0OfKbOejOCaV6p8OCQDFXgD++s94Fh12JUn
ZRt8aZ8vfN+OztGO/hpApL04Vh9ZdX/1d/wZ5b+r/uPaIXDCstbsumtNMcMyqXsHjkLh2fCHsp9e
zO20vxMvyC76OSGtMpfIJz7TPxfT+LV5McAugN+IwlYGqursvwRrEKO/dNLLoJp0e0nKI0n4bUCi
Z4cvoP7W28yJTTehr37SEnjsu85ytLhrvpOTrXw4jUjAwdEZSyhWnVmjMMPlnbAYs8p/JvOC6KS+
4813SNXKtDosJ4pv5F4ghIEyURXgny98op6yIUUfjDQwrTZLwDMnrV5uZ8U+IfnRC4XkzhBzG50F
SUoJvY3hLf33+5+Y94/tsgGj3YrsL9+OIiCam3fG9kUxvwWMkrXcdp+GcbHjALwXjrpYn16rFgiD
YFzwuiwFm3jKuBGMkI/4iBiXxv4i2F0dOsO54zVDvSyMRXtgFZtJawiq5e66wyKsOr+7R/ZlYz7z
ryXgOmS/8nWItUL2eq0C2eeuJfFtOwoepTdZvg0u8cfSoCO5f+jd5oJ8px7ii3vTrcTK2raHPhBS
TNg03MRUgZoxr4j7qlRFp4L8FKVEbVu7cwIcgruE1B2K/64G8SzVn3P2p59/PUN/rdx44nfTel9x
P68O9lodwFcbtOK5I3RFFS9ABUR3SQe05UWOLaAq4C+I/zzdUpgXxGpNr15Pbn6XAP816p5vMMkQ
FUXJIXJyZ8kNtRqos7EITDhj/tJxPtIRPl9MhUnsljzUAIB7WsxhzEkjNMN4zfFtTxKdDdfWP5jw
JkLlZLm+2d0GuN6PE8A+H0550sJX3/YL2vJvGxYRCflMecMSIW0eRb3bu08ymIwCjTVxUs2F8kkC
ZxDEb53DLITJH5Amxj4f9lXu38pSoVbTindCub8lJLqn/ZBJve64fZjlfyG2r9kfV161h7K98VoH
xLFgebRayKhESgkVhUpEzQvHnXNgXUOTO+a7HrTCci8YxcpAowugVPNfXpbhoJjcScKIJXeqWZMW
dEXIXSK2NWdWwHKsOBM6QETDHrXWrpFoi+8sStYu4GzE40LaHUwaQwYMvGSMJDYWvVhpa+3keAob
x3HhIjvEMABeC41zqckJqtPaf1y1XxNJDygfEk3ZmKkDuDI5xbfDqu+qy/ZipJ1VHqzP4ciYX+Fa
N8Dwx++SHM6hfdnllP6Moggy628KnQBhZPMKuMi4SvfiN66SIDXxMFCcjt4JrlPOIwHHOprprZKh
zeiT6PSKvZIYgs5MUNizod37Mmgp7ghuhYLSN86rxxeL2Ty9F16o4+la2UvSonU8svC+geF4ec33
PyVbworMm98XjYFCpkbXDPlQKYLjI+nQ9YO0bzBHfxFyr8kJfPDFK8vtx3YAbWuIDi9k4uZ96K27
VJqhPZ1u+FQmJ6Z0z6NSt320brCsMKFYLI2nDsKGvjH07YPpmsWsEJC5623gX+7nCV6OYmzGLyVK
iav6RR1xbLjRPNtQvDlrMV90ojDY8MIOTFCXe24mXsmf1LeYt9Fw8ASUR03gBEL4bA4HXfbdtBCH
vSxpPuCg9G3lUUeovNWQg/rr7bIXHcCcqEfX4aP5zORdlp5QsoOCOFtK8q7aB0RhdepGq9w0Mwer
wDHJgi57TFqhE8Mnuq6zQHUSwsJuSanLC94GOVWHAso6C0UO1nhxyI+7EHmNbbcJhxTcTrf+u9A3
KZYPfkBo/lGmKOaaReYQnZujP+z2PymDz5IXVb+Tc2m2ooMx0n0IE0GoEHSq27/0p3xs4MZ/P5D5
zQnzl7ElhGdqMjkoXRH5vJLLi4b031TN/kbupivc+pZt24nrT76IO5z8X+u1nBFKsC31M2Nqgx+1
Wzant9uvBcF+to2FAyxHUlkGTXcZYM5l/hnGGCnj0fR13ZHx4CzMsTav5Y21BxtIVgBQv1o2FSGG
n8ZUl1x8BtRkY3GEVwzWPF5daJ54x9yti2rhPw4SArObHyreb8qDkaA1xjj5OpDCh1iu1vJ0CKK8
qn0SrTDKXggSw90ALYGGhiIiKkgKCyPXmLDgSkEhZayK2zSdwpLPhnF6t/GTTagA07xAJO0oESj5
mXSdGQ3gYiD5VoFzoyiXPHpXbc+wqO/WwIF5j7OOBKybLO9rPr6aRNdm7xbbZPrTPmYkZaToAnqa
iNb+iG4BhPDUtyyDdrpWiMlPNFpqoNa7C6hNIn60lw2JFpVWcmoAigLsci0ZtG+etQKaXK9ja8YA
iXbDDESH7gZ0TGdaIAF4HITT2w7vQYwyQH+Qu1zRXTVN4CkWq7j+v/gVggOFnFBpIK5cktBs+AkL
6rX/NUErZXyOA0KzWKdlUV/2Q//6ffNqRwWnEETU175/y49W98RYBp8r4BhBsTDwsWTpDzXjF9KO
Oxj8zDi2vSRPjvVHieN0sH0wUpPfeOhg4tLFY4/4KeXYvyjN4gx4W69NfnW0NbDd8FaCVLR9Yn4o
SSMn5H76NiF/qCxTCvGtCZ1AHVSY46Wu2XZ/6qdfPawd0RFh3l6g0KjIUIMQWRQLUAbvE5fRdbDL
ET0vD/627n4ZR1FLMXe3gnsyf6y+RypN71rJJQ7YwTXVKDbERlsL6u8vSYrEPe6E2BbfYTrbnYC8
HLNGxDDXbByTP7poOSWlyhW4nuDrHTiybkd6vxiKXKZUQnRvuPb+fNf0ZfKBsX6I38lyLT24KIEZ
77rvk49I32R4SttHHfQmgO9sKBjOdnkrkzATneOQaZd4Xs3zcNg52F7IIgpa0oWibOjwrkk+xt70
8m2p63i/9fA6emJLaGTdkAno3LlGLSKTYMM/wsU2YOk6tbouNDT+/bfger2bSzZnZP/yrGa9xzA4
H/2GytRBjMtRgXr5qI7CyBDqX+JnyrqIbMNLmE8UmzhuZQU/WYMZhGFNL0nAbkiJtyA6OslYYrKm
ajnsmq4QT84E1AnWTzkxDp/HMK/fPpKsGytMqmGUD66k0KazVGOiaHKXu2ykql5agYrPme7O3Y3F
nuqRCQNUftbFP03JEGfZQIXl4z5fGMI+o2lYgWckFxWy/qzKMQyU/NXI66rTVXgpAnbsHoumsopx
vxHzj+2KP5yGyrMkH6tGAw7XVsnEOdGPa//Y02D0KhDfTQUwXs6EEUUNTw+R1HigkkfaaqZRTzyT
OcbUIPJfeIZ+wMRVcHgvnGdPaHgkRwC8SO9IuyfDGGFoMmW8WuNkrtX/CsQR4TJYrzE0OK3wKeky
3+9NWQsYa2NzkYisPhkvxTmihfwRgqMd0JUCgMJHZ12BVFPX1ATyLelZvd1g66NUdtnQAvBilzu4
M8F2cmgW49acbzxYbsMLPVtMuRPKrZdX3i0g1oeN7/lqkHW8aZfGRW7gGft9hAR4Hkeq9iggQCYx
avD4GQHkHiCRcxRiACkJr0kqMQS4BJ0hiNEP0fCbOPwSyiylGnbhIOH2bzRgcPIedxJOD121vGNO
FTeeBhknkh87SySKkqSotHCzze+2Z9ccD7TidcG/LZAXm+Ty5Z/WVgz8mAVJQx1iCyxghPxjdRUr
CB7HW+KZWJQoSvuAcacI1qLeDeXmPrxXiKi2v0orOkGrUm1qm8OVwoUGlWKn2ozFOoVzXFmJ/XxP
wEaWSpZZWF7HjcX0IU3yMTrzge1szGWfUKKEfBU8ENj1PJT/+vearr36mwJSta5dCbver/Sde9LD
zIV3MLTSaUu5iesWFuBHZ6grQVtc48QwfToNnR7aaNc67Gpho20iUuI98NDTkSxdE5DFt1dbPZfs
k5QEvaL6BvICyYQ38Fp+V16f63p/v5xGfBaFIalflriDJ7v9pZqwy7bAX3H3sORRHKOVJ3TpBT4z
RSctXUEQsVbR+N057L1EfPfWAZFED3qwhPUA3srt3qNYEVxWybtAbv3mlcp5vRtwfkWpqtdVnpAh
peJshE0pODc/M+HstsJ9Bvu3fnKCWuxIIANxElLiek9+7zWdnWnwnW/y3UX2If1M5G5lBesmq7eM
Q2jli0Dtk6nWcus7GXvl4ko1+n3GdrWmeouRI8ZhLf/xnVRsg9hQgjB2UOh7o1/aG0zr+JmAUHUw
gj/iO5mzPFDVp1DErG2PP4ITqRl4mCZ7bxSqn71idenu7SLh0GigTYkkY0iC/0EAQdgvcVvkQRTg
Xnvf0vSKKfh1XoUh1ORQkoz+kAYwxacF/OZ/cO6I3Je+McdU91fk8lG5ymM3czNEzTgeSPQ0olrF
QLGHTr/Ob4imAW3NheL9/WAlcQAxX2avr+lrp/2JUEhVMXFmwSXmaDFfqU4gk6x9RbMYifa+yQkY
e0CNlNFl+NAYHHZs0p+vK1FqowZj/xJ7K86VdbOSMHSYeNRxZD1XJf13gagMJrtxjQrspySBG4Pu
TnuDwF1OTMo48SmxpfudWRUwApNDGETxjKPlN+LbaNrBSCnn9MKqckN24N0GLXUG/7WuT+UWB+dS
QNNrk3zI+cU4039JGX4w97xoQCCBqR0887PSDPjjgRO+4hLs053pzl0bDwIBNMGzFSM+JvZI/zj1
1N3NxafEpaMLCl/KTqHTtM5EHLI0CgIAAUiqHzveQm+nc8uFQYHCS9jFZWe+f3mO3e6xvu2j90nI
zFmYQD8w5L+H4a0HkFzXBBl8qZw9j4IILQYgxLTerSFMwIPtLercWk6HnDqTK76s77nb4GTmTz78
tSkiRg2ZDRsj3IIM9Hk3I44JsKYowOpQVdrEeHRZdnNYCcWVbi81czd9SkZxw53HJrPwyB26Co01
W6wLQ1lOmHgwEt2rIQW1VmarIEKASQuRD/vlH1rMulELgYrkVGCmLhRkQp9jrwG31QBoiMX6vxZK
9MiCz+oSTEiUNPuHaidfuTF6oSPxQgSV2XXzVjGdRij0hZ86iBDMpY+5iS5rEnQGxtfd/oe77AC3
IuV/GQHUVlFTyYr2lGjcZLljaQfHlaNNhhSHghO3R018pH1VpFHCWfQJyL07jdBy4vhKyZ6zIdqj
X/h+qqjA1ZDVLIplUdrG2aU+ijSXR6z0jc4IsNS3Tdm4EnwTdp9r89gc7Qs6Jspo5EH9XKnk16DW
OaKlAinbYEGZ+iXeoU4fySJ8kcHZm4nmxkpr+j06UjNbWL4VFI5tYU0GM9RVhorI5yl01lfFWTkE
AO/Luv6n/YFGjt6Sbe6CavnAFIRit/nONCzo77WXViYIrcSm5A/qaqDezwPdrUXOroLZF/m9y99r
fOfl/hfT3nwpdX5d90soGcplMzyWm2WIhoz0DJfoj7SIZoUU9bWY+SlKkRJhktTMvs5wynPhcWHp
iKzymbIvAmH6xIkvz6FZOPzCOfeGQ5ptFJRzCO7tiM46NwaHuuw8DU/Y7ZyosInWamIlL++vAOLw
reiAZ6crjXfoUYjebWV6Z5x064ghLAedc+nbNA012oWcE9drTN+uTxOrRtOrov5eHNg72xVReXzD
YCd9kSroyRURBIiNhUlaVjMy2/Weyr/hsBNMu4gLbnCIcVkQcSU2Vi/di/jYIkAbFZvBUMrxbFNS
JvWQ3tF0/HEHb4akYMdpUMYKc1dyFJNJBKEXpUP188lHVY68PDdoBSsqLPGr6SzzH8vbjxZJQqyf
69WiOwI2RWTetb8rMkLXZ3dcIgOsvbjiyT4XP/CPMjUY5Tg8/eDXon+efNfNdj1AtkvdsYCcJe4R
YUECTrbaTsJzE3uyUirkzQ41Apb08IYBgFzSmD2iDKGUNeJbIr8Fi902dSZB2GBxyGKxME1vVU0N
v8lvIBcWET9fdA4EF183bFN7sKMmxv36ogLh5PUf7BVZ+DwCuzqS8CGt5PtQwSCKFPhYUTfBZhS8
36BxQAl8UUd/KgLxCsJvUoAVMhZm7SKKDl/AT3+jFaQfWaa6W7pGpC+8Fh8svzadiuv8Jk+0FwEU
diUV+KuIislk7xTBdrw2KtjIqOhJdrpSpwDwU2j6v03LeLXNu9V6lYXTiCKf2c84BV4M6CDC+ZYn
mr+ey1Hu85Cmt6QSQkU/7iJGu5BG5xItcxUc26rol6yEazWYBYKbfQkGg4CGq/WbJ3l4zWJkxYrk
DHRW4RvLJRptK6fGKKHuTUAFiJR5AK52GPRBZ+6MleAt3xwfzmlIhOHG8odvWPtbavK9obaaIJ+L
Qnsb7UB+DmyWFKYlf8gM6L5LSsJAde4+azLHYpqRxIfdmcdwGis5a/DiH410vWIGCHYUzn6A+T6a
9jbePPjfTbNY1BnGyxhVPHUbPqtXT6K7zexlJbfw+BPTH4Z7Qbp1cTgdiYcSf/zshHs7hEoGv7Nf
OGjRiEmnBH4HdFulEvC8Cl2SHBF7Qzr4OECO8ktMOEUAB73K4xw5CehQ2xEeb+NU9yXx/SJEwLUS
p7GmRWlFxUyI3HhmKkpxaIUhSMV7geF86nQUa13NjqLleBDWj7RZOIdEpGVPsohlOCazlLaa5Xaw
54YBeVy7pb6TyDL8slDXS53s56lexCohMUwo3Ry/Bz9I/g1HIDpau8X1q04PoeeNpUd9JVfv1/NE
vmfYisl0cPvYtWToRD8/4D1offpy0yfmqoKZHWvmnFbBwgsJXnKyL+7RB4939OqDR69YGSZbZWa3
U4Q5hlhJiiQ15Ph7ltbN7umATvNwrVQABK5WUtkmtAqQITbrmZoibgFPoQtNvI4c/UgcSOiajBvf
MmpTwWQlO2a68bLewY/o6Pt4KH4FQdNwNkPkSVOtFIor7RpSzOtQ3VHTkRx+0AfsiiyS6sPVwtq3
gYUBceSlc3I1UzM4ER7FISEX1wSeYhxrmPnScEBArUGNbRvY1Q3vKxXT8/UI3BNWoBO3n5Jd+TX+
VyYRA6z/tVFZKtxnXC5kvYzE7Chwk0iLu40r9z70hsoLzAo2m7BfbMjInPWeQ/ALApnZdVz3HJg6
L+CWK1/hcWP/h62c9Q4qUFT103hceuh+ydlo+QnbhVSmvId5k51WmAJXxPkS95FRT2XT+CMDYyts
yxrHUMksdwSnEuG34qgop609SFxZaz/DoU6MxLTc6VobXewjkzKLEWymHSZNKY7BwoKC3SiDXZkX
xFPxpTI2yqM83FZJ8XoeP2cSNTfTCRyZOCj1ReKQ2iK9lP0BRHn77uose7rThHSpn8rH6fne4sNb
InGxHOvZx++DbZ8IDN7Ge5+1b6HVu3PGAeVJG3RgOT1n5ZZ9C4oDgI68CAh/HZ092Dr4SUn+B3m/
/zVDerVkYET1LqnJhEXwf2rnrfJmmScUwUsE469PECAb7wy8H0+5A31IeD9uW0hmFxZvN3wY724n
zeNxbjY3BgQ5TYs88SK39XQDx5O6nrvVZNKnvdGO5ScmIPKM+DnPE9bcN5IyVyJjxEuE2okAakPV
6QohE8wPa7ddWPp0iaOdBsYG2SfegAScKTY1YsQ2BaIb6c1Hb4SW+/NmxM8ii2BSgv3Mt/BMYpKX
xvFJFEfRBSt8ge8jqbzCM3ViqIPMMoFi3+ySApy6CClWZ6OUGQr9PCJlFel/P1AdcQVGA3ZehiEH
MdOfoMsGHycdiAG+dQADzfvauZ7KcumY4qb8C2PRE43FcwPbRZkkoxR9cdlafLa1QcR9K55Z1nPA
f/+ET/O1FgGEiipHOhRjqGvihmtt4OLYnvo+Ed9swa/eVqVMPAt1r1dpk3QBnDXNBocbNfhJatXF
Wd2AnE1nZNX1dfk7Wr0U37t9CqopWGvKF34CYd2XwWmmBNyTgA5SSv+1CcB+cM9wmt9aDysUq7SM
AyZ6CiW0H/cKyEA4tko8ZxH7AvF4of+CVd8cRy5m7gAUiu3n76HG6ghsRXim00LLCQQcoHp59SFk
t+nLbeUMbroHVlOV60+nK6YucEhyVDIez0gv7IDODeIzRYFfsYUihyPnVioeOITeYyV3AFad9Twm
ujL1zG1XhSzDCReJZmixPUMIhHdp5jAZUBixRklCNwucZ/EEKZgADjmglmjRtMsH1InB3yZWSJMO
W+9xfklMB80vMjelcUR49JWjyfH3I8LDrSH4gT2C+e8IjR/bpGnkC5WE+AjXw1HSq4dyUzbzYYtu
/6R3i9A3yPqUIoHE6qMyoEVXYEp6WLKTPbGs2+KABlDVgy9culHtT/YnTRzFBJKKHKkF6pokziP8
TLzh+g9MrwYZB1VxsXQXvnSJ9MaopSDSmvSq3ZgxoHYd0MSJSbYaTCeafnPqisssTt26r8bNM6AL
kPbmg5/7iQU9Zjrb2JlWRcB/OFFozr8gO03PMd5qhyvMXq8geCw7VyLXr2fWeajYWKD23jlxJHR1
mHusAfaFHP8tEBaKnh0chYkPBFcbDSGGJWtlaVS7uQEd0f/hvzmn5o23V26v3OfBZ1dGCNcSBFnq
YXDe5nYYw9U5opwZ6TvmN3tyQfFmMArg88zaAJxY6V1LvvZGjlH8zqknUtTS9PY5kYp1VpZZsYfz
L7r7ejtqoMw6V5+ib9GOni/OERXKx67F/YI0gKsqOVJY1uCKwjP3ggEaMAokGs944f0TMDMyhAa8
VAA6aZ/LaM7MvlTCc5jYjushKLwiCSmbzQJPmvXgfTGWl5mcY3LEd0PK2u3LTKIdUbAcyQrRkhZ4
IqY1eq0GYgHMiVyv3eybC8+4eor34lxgOK+fyY6juo4JYN3rSosFkkN/NFEhGNe5gKmQgWbDQNoT
eJYxBtKcBjkoCO1cUlzgINHf1RD/gZOfuYbBTQ3qh1Kd7Lj6cHZXHCSl3bKB07GiYszUePY1jfpu
0hKczLg4C8EVx40G/v3z2jSS1Vgpi4M5la+SM+4GK9ULntUd3fmU1pJGUZibyKCScMrSF6mDcRsV
6uZgoGv/ZPfQMdg3KjXIK9nHiV6socZYBS1c1WX/EhKUv37KAvmLKf7RE2+H5eUZ544CyMmzs1sX
SVVZPI+wCL8EHUxriU94VjxX8tawfGP1Y5Kf2QB+XLmiLKfnL7PC56MWHR87W+rUWv70DKNVVBLp
mmwCuealftKQV4E4OWim/IEYhmG6VeWSIVvX6Q9U/9GHbbtpPlqe/0Q8Lrf92TS9KhKNdADfcWM2
6/ZOdCOJkG603nkYpaZGOV/pO8msSkkA0QdLK9xYRzOhRT92+12hCGFiDS0BNbmqaurEdTs5GojD
4ew7jEfLWeiBALR+US5wv5Ocl18sgtRXsYis0XjBwpUGDR6pmG13p8HpjLyRgZwzsGVGGbUmFMrs
IKy+ICH6kpcaRcq8D2jMEHzylLXsObhQ293psP0go0e/KXhhzD5gc0r/3HW8JyFjJwVDhwLKivUN
wYB4SbqAW80LMJFdOUKGC8vvENaRJ8NS5Zlibcy+oMmN9MPIWtk4g5l4MGSpmkUd0rYTPWNNvUM3
woaZ8+Xm9imfSOj6YgIXbbS+pyfZ+Y+ozb9epplfzcqkWZRbfSdKObhPMHSjqFnVhNEAZZOg6Izc
TShDR7F06ir2FHTfahZOhwwKsMJKUR21PSYEaqcfxTI/83kE9pmJisGejG57Kkh3qD5OAwAB1xe9
d1ACNQbHMFXzebACPhUIVsfDiii/m6JRBUG8UMUAfPFPAf1Pd/F2quceZH8EPjtNsI4okzKHU0Nc
lpqEW5j0CNUvwTAko6YlpwIEeVUVZB6w157YXYLY6Ulyee/uoxTFA+M79rIY1tObwLeWlpOVwJq7
hy302tc+bg36SzrbOYVr24KOOcXKh5kb2rYpF82k4YAmu0dljIfKkdbDaH0VfoEfEwkR32gFekNS
zJtAAYTcDX8BsO6Wf2x7Cn7tMfSGCPhaQ5brEmNFo/85AF8UcWbPzf/6Dh83rfOurDTXkx2FG0Bt
qDXuSo3sI2qPgku8EfWSk4TdUBMWcdg7mG4MomSItmpe8H/WpjKeDKXmwlah3QEmqID9eX8QYcFB
Gbtrl4yWj6scDU4kIRTDk7cCr6zvKdvYacD3Iv5iqenXHg6diauT1lHsfFZwb5UU0FnR71N8Pcn7
TFHtWt6W7rvpdgE6oOB8trIuYuUrpPbxSpDn/WGm3+RIsQoKIhYjVlurcf/LAm9O0ilcvGnJKPxr
nOhnOwbz9+vJBxXAnARQXRHHDvPtQ81u8FHghajvnVE7lYD8R09s8JwNdLLmcD90oxZgGLEO8PPF
Eu3k4vA2PZYURDCbIAhojYBpt4OvqpdKa7ztGov/OUDYVhhlheGsaLN+jgAMcA/D5xfvjVkzgE25
KwyfkKJ2DnUBNVQKo+W+RVjTvU8XjjiZ0PSt2ywyIcVBB1bACuhYUCojN0Amf9MkAUlYjkx/VWYi
fVLuCWQRfLg/jtBIJa1x2vAuA0sTe4BHbNwev924xicfKcZ0fOpKRxiVCoN3kceQ/7V0Eboq5ZCa
PD0l9cSHGNNvRU5A/2nrchthmsUofl5yG/GaAoEHtNcPoaPz//1lJJ5lHK2nvJCApn8CWNYGajHb
vjseGLGL6wPH/us6ACc7hqxhxKwDy4alzH/jYwdvC2rd4t5eSkw273CMgtU95OsLT/TziJFfLFl6
0TZJbVazCHH0zr2O8VwEo8IFrrJ24mhMnssstND+HYzj8hsuJCVI52oOk+yEvVtxJunrv3JPMQDd
f7Nqg5XHLKhpGU95rRrS1GtTvl6/oo9ies0I+NAtW8vD7hAkmiRkl/1yPhx8WsgleKcnj3/69W7Q
jHMe5ggD8Uyfri6CnQ4ywgDM0JTlz3H47QEJ6UM76fLnb7m6Wz0TQIEcEDN+GyL42AfnH5A4DnxM
r/619DCqGmCIrywENHC/0Z69WjIoRjYGOwAklKM6LTcEZ3s5BDkbsHanDf8wuxC07U4CwMgyqxze
zWmA4bwbLyfnhSByHdapuoTs+vImwUTrjjoeCo1YsIS3NWouuaFA9TCRpWRhc7xph6EI/NBJ9F0h
ARI/NSrixvfAb2Wv/IjsDbInXZEkIBDtStSn04QZ6y9jFceY45CBLQfOrYF2VtfTEKBRMRdAscgv
4q0OXGTM6hGOm3aWQe6j6D/tlExmw+KZsQgPCk6FVytufwAhz7maAav4I9CJyb2imF6r+Qi8rIPy
BjXAsUG64T16C/l+sVffAOf01HX0tPDkKRTUebUtwGLDJvF0y9cJRxez6/Bptw1J7K76/xgPj38z
X7/c6IG6MoSu8nxaKNsyLoZyKDQv0O/HFGum6ykzMYoYXieyQvtlBDnyG2aYVK3Ddnuhq+pqrHAC
ePGr9mp3eyynKCmDo8543cemZOuBZa2sEc6xlZagn9Gkdr6mvtZ3yD/9Qh0nZiT75T1wBQKcxwM5
twahRX+ugBBYU8EjMx6uRzV3w+QkSb86THq2602SQvYA4tDl2aA8crWMjkIhjUh0cloJxXtJMEbm
Yc3F4ePnDX4i2Q1o/3Zic7GP0QvuFC/sXw5VCtlmvGt6znAvYQHVTNtVyilUGcwGmWsVqYsNjlus
Re6Nb/Y5B5DlkL9K+3fd2yuInZgCjee3H+I0ehvJwnUUSyMFbHr3+4SEFR3yWV9e5rIRVW1rBmya
Qq/j0S8Zwkw5pNMzu0bZ2+wiS/GahkLDVySykYHAhGpCjcEYM+YYoejmcrgsYowJk6onQbfOk0su
/qsdt8Mo1xC+wbGokpKgFWYfh4Lanw/DXJ6utHDJ7X2mDiZkzO3lNEP6waZ01SmNmPbEmobb8xdj
E9tfxqJ0rIG1C4juFRkzwLf+6UDUtScAWZt5O15TayQvdqFN9sgcgh/Sg9ebfhggzvhyOQrOi7C4
3z+wus4sgd0PPBZKRmdGVI9O6EX2HRcr46/JSCdq6m/kOjg67c35/Q6pnKi5Z80qrFOikGR1eWoy
Kx+qKzjnPGq2IwgQ8py1lYxc0h+t/jaeCdhYvDmw8MlzriGncwDAFByAgkLvjPJSpOJdiRzagnOq
aVC+a2RHAMJQMQtJ1w7pJHy3xx+UKSvPI0mBgcY8/GNhR2i8G5DYGASmwcZ7wB75PiNrQKX5SWlk
CuIrhl7UBEd3sgiZfUWPl59AfVMHXljVxXVfp1JFKSLkSaJ86DLh0PBprgiayFB3qlMU2I3xCbiR
J8ZmS6xrmrz1joSJt8NtGKJrFSbv7rIpIAoYLSe5yq268sDzygqp3+U2OKiwkJMFESZ6zF2shCOV
KCUUpH90JLmRrHOLuT8JSG+GfQt4ou8+HxJcryjX5tXaa+Zk0zv5CM/yarZiVOO1dc+bNLF/3bEu
S+/DHx36a9ss0p8B1/a/zapwVxyXE1SetzjlpC/01SWM7zS6V7E6kXeroK0w5r0EXWWRZoFw4iJ/
8xsB7e6v/SVWdPCdg2TdIKnQTbkFuE0gKp7dy621SDfjVO65mVEXD7GzEPI3fDsSHLOoq1PpBX04
v+u41jda8vD3YRyeigbT6U4UjsDdyN16YxQFrSV1DcxOxdsFquiuV7GVVJi/ZRhoD5EFciHDFnTz
V5Q60Bzw08f7U4tQjHOXxeWXuOyd2kCeryjdoc1Gk3HSAJtziwd0CszhGrxIAJz7WcUgJqkrK/31
xqHxKwDH6UFfUaOzuOemg6bAYG7RTn4ZmzK7Zds4GqKgF+QeRAvJXaK0Lm8vy4tgLMVIUCK8NmPJ
LzNrCWyqGxd6PsNWmwRm1b30qVdUzcXxH96iNoJrbhcOghpMw5xWGyaYKLf+7mt7/a6AO6Q6xVTU
+ze1jY3ex77HgxXiX4fAsUKGxoEppV9HfXX7cWKBGiCmzmufvh6llo9HPPctxfCyQqCn1bZIi9Ju
/j59+Oow38qo6n9OL40PgWxbrKs+dRMGEfIMV/HkFLV0qsulcKjH7w7m37gL/8uyxuRCPpfAQodg
iYWv9L7WvEzHPRRiQRXi6Svn4jfLBjAC+jxQEIZDL7a/+jCqynElv4uNF/rTQHE1o7cS9UfjvAw+
Cjj7+VLHEVPBI2BV3oe17ZFJitvh8FmDGfcleH5y2HjgbdYv7N2a53I+sWAulvWP3Y4TJViVCA8g
UUufClDz3nLUzI1Gafpwv96abqyQ/nvCJeQTl26IGg14blHYdFa6riZtAkPE420RLd1a6/pZB8dp
XMSdPwSZvbDooo4SBw3MnFWzoeb6ZAbIlnMKhpXQeca8HwQGhwRIUnbHd3WCb7PIDW9IjFq0a43e
nDYafM1HQEQfKiCStjMWqX8JqUK9sCelZdu39NX5fZ+Nuq0eYQtOSimiNJVepfirm9bTxXg2GRM3
3zlc2aPgpUiRpg8VxoX6RQNnIsximFKTFeNWyXtEIAHiGznT0/MwGC2VNdHDQJ7eYLQ4DTcBgc1Q
WH4hPtq3y34emcKKNn+GV1ZwahK2kctSasFS1PKJcrziIRDHzTOkF9zFGs47P9vAwYCdQ4o8XgbR
np4iMMLCxoaQHCSo0eFIJMTAR4Ig4DkE0whrkd0ZemaAkl3ZzRf7TDrqEj7NFZ9MwJjCD/v1af3u
IwIlEXz3NmMErzARS8l80+YwnJUCNBZ3eLzU7oxerz0B6KlGv91kAzCWDyMNn35+YF4+Fb8d69BX
cLvIhJODwPP091F85KndjhIj9j4d7n0M0/7bJSJRfSoQ4EEIfbSDVBWQvgPhgmPT2oHLXD+LvayU
bFBVdPJ8HWNW8E/WwI2Ua8ZOOiqcP8AraXmmNwV1isWZqdPw27sdCXJBcyw8L+T9n5MowLsinKu/
XfPKx+RsKlotuqG/A1GqquYQ+cXZGw3iaXQ4IhJVoBRTbbe5Nv2ttpg2EunZZ7s8yAg3FJScjjLR
JoZSCsN8Z//YenHqTkMxokv/4oH0oQ0MTveU7z4Jd8uRdomRXz7O1WY9S5BBtc96KA7ICLfBxB5H
5wiN9flj7G5Fxle+CtxQwYyO6UiS/783HF4+sE/gpiGxPkqDqTuJarRUR/4apf1Vg/P2vAJmRqyF
9OOfjkIXqyIW58E8QoiYmMUDVzTzrj1FIeecqCvpl1uCyJbd6Vr9MH8v2W51Mjh6bkQlu8brjLnw
6EXc6A6sxXzlIzkv7uLkSAydspxZmelFOKmP2XJWyOhGqNpNVPRcy+NtAS/W3gxcY75RsSd8FBHg
FsJljBMEVxFCSSROw7CXhQnNlL656SB3wKZHnBXy5kpky23B6uRUsjWXcDdlzPjxOF5wjn7Y/FEd
EPkjnpXxNs2h06fcooJCBDqZSAItz4jzGpHgYJR8Jb2S1BFH+zXZ6QfFtCmCZ+6lZoTOljouqPQU
Zm/HEzgl0Ihif+S2v+FG0PdRPc+EhEXQHeUXyGUWOJYq92S7Um3J4r6tiT8mc3iYygvWAeWet7TZ
Qn0J6Yzc6rGL1OVGGbX/gK5ksJtTYfAavAOB81a6RFKQDm6joG1A13O6FLvBH+26401vE0E/8nO0
RNqW1nnDuGcJOM69UPOAZa36Zd4CVsZx3BmTYAqptDY/A9VX/bcya5oiiZ73FzFZBx8Co0dGFNiy
DpsOmqdhzVgDDe3a4STWvDicImoJ3V8Q9mO/29ds0mIsC1InSh9pzj4Ct1WmSC5wFmNra/DbkuN/
n4mdtYdrtN/xc0TzmSWDcUQi9V3eR2OEJNkst8My6tZCBNFty5UtvU4/3iWjEvtn/9LOOyYmQzcx
wlNT5MiivqR7el6aF44aSKDLXccVWu78eGKFNh3o53uD4AvphQos8zm2Vrj+BuI0JgGiSbr26yxJ
kxUOqQXaRnDexZgzibbwLav/0aV6H4y/HTsH2UN5T42zyAp6XqE7mAm+pxuEkVJqtCwlGTZt9c/O
kaDsKOBaIiojjOY93TsMhB7AzvaBXlXec2OU+X+1BylMXME6aB7r6bjPglNvTxWupq3O8amwRzqg
7/rGl7M4jXi+P/Gs5WfE2RsiYvtU6aPVIVfMfVW7f9KoGZ1b6QY1ZeoC5OYPhR5IOC6bgRPwkrCm
8uEiv3/owwb8nO7HI3Sr6vAPkwwyj+xlxxgIDrJqimAikvym+hTzzDuJIWtBpwfJvETeuPbsYapP
xhagpu4a9pmLaZfETL48Fhfq5fAxlo94k6HXXjPZ+DOoUglI6RmhTCeTCBRJgAEpDCzX30lggVGj
gVbdUMh5Ebw73w/bhzYRqyo81tRKJFSnIDbYu9TF0unSS4Yz63ZpERlZndcwZERy/Ox7gdE8GGmz
xdh7rheYt2B4T0280pG7aN0Cwly5UuDhkBzZgMqYR9HRSQd1+R9kDxuGas1y1sUeAr61YHaMWG5j
AvP3+Nm5YZzoXY2ydV05VJEcNSztTRfuXoBpIRxQOq53d/qcsTAEcBt64da9aGZ5BioslOLFCDU0
pcHWmYAjiFClDIjl8cXMDJ66RMRl+VwBRu4YsnBnRd/YVPBDgP5VFqGK0OiJFjrfT0gjoufn3M0k
Gx8j44cIt5OWBpyvoKGN5+tGuf4YpoFD0pyrzypzw8deDoqPxB0vibBeWDan7upHDwaoAfjuLh4j
itfrNv5Lpy8DQR+Wmi2FX2BhxlIyttgRBsSrjQAuZ3NKrDAk1gbQ8BNALC+AfCdenw5K+E1Bi1mS
Kphzq76crA8lfiCvpzTzHdxw0ga/KPKZRgkNlzTgB8ybayhZnhSYMwUFWLv4LMG8DQjWYTG74JIC
2nGXl8S4tRI+P+RzGYYQbEV5cYOf9YXksdgWa3bbSFbpZ8VXocT+zHmz65Ne3dqjq+zHtbS3Qx5I
HPp9FP96rX8sT0Z1kCQrHBmeIMG4B/W5cYZwYnA41yEthSH6NWlMBrEsda9x4AMRHxcqne9UdQtB
lmE3//aTC0G9vM2aG21yB94zep7ThO+9mjYYTPT0fuglWjvb5VZr/j6jMp1cMfyOW/nSzgjniSCJ
yAn8SDT3yw2bLnfMo+TpyEr9ivXhbkBQfaMhirQkk9CxZur82QlOj7Y0X1ct+EBNw+eK9pvEbfDn
botrgwdfAyYcG6FgUbO53FIe5lkx+IXkbdp6o7rFJhN3ue6W1z0Vj8M6whSmXGegqRFsFnTtPG9c
g3pgE9mNS92mBlo+EMGa5/t7yVRuINyowcpUwxCcKnZxTtT7wBT4XoJJcY5iq5WF7ieWxNVWgMSl
1ggnoKLPA/zeQvh5J2zzXkwXJBhM5bn2NTSAB/76n+vRJESTxcy9eKxGuv7VvPjOchnB/LlKo4LE
n1PmZ/YLTjvcIWng82EZ78LPAF4ePNkdQTS9faqiChCNgQ6spP/gv0zoMDJ9AaQdLlXe7gT0G6Uc
8RaCAwSD1NcZmZgkIWwHsPUSR15Aonq6ec+plyc+lxvtcMXJBOMXH3kvzd38ggngVT5H3Zy8VBLV
1uZCO6aBiQfuKzKMfyOtY1eU/QsBQrBB9keqKHORCAS3Lk1Tzw4LNDqjYp6wM0X2MWoTONQ+BC8w
oP3BSeOJMrbdroqzafAJCPwgIAMafCVdpX/dT1UPF4s2VgzjY50+Q4fT43H5osfA7tir1QuMMgal
4sqx3/8n9XPEhuX0HIXl+EYT2L4xuV6xvmYily5NgubLsQVcscmB9DeHD/HcB7tzOHjao71cgGaT
uGiOv4VKWplPm/RrxEs/N3o70F86hZ3Lv1O8tEh0oK+3KAtljeMr7650I/W0Xzu3l5iaV6bopUur
1hQPuToePyvO2/4Fn7YHEEMKDnatoz8GWh5oxxmouq9Gg4QoA8EsKwmatlVdmYDMu0ePYqNwj9XF
Hwgbtava2ZZ0t3R3AG5HlaX20TMJnfCYNazOlubohWe8fWw1P8YMq0L/oD/r/P49FSV/PClSVYc/
F7idAlg2F+k4wPRFfUjR9VdAJOWXu0oo5BZBGh8ndmvT/pSHD4pPnFGFhHMF+t4jtqxL77y8wqym
Yta1t8TkU2G7XjKrQdj3W3Q9JDDA5zS5lzpKmi/ZipkxFxTh7YlEml4bSEF0oA++2MjjHggbwa+K
FUGYyyTOStBF+I7EnleI8W/X2QcUFj14ZHfA5BKTPLOOYPoVI+abD/ynmL1YSXc8PdVI3I6wNXo+
OOzycvaAt2Yoa9U58Oeqxnbo1NAIqclQwW8P18yOJ0VteakgJufG8/n0VoQa0seMpVuwpdjxMgVK
oHabl268ZyzgVooT89FrWdcbG3dIRtwPXy9ceWusd+39axSmR6JxLXlVfGj3SMwR2CGjCYLExPXz
eJoZuQeQa2ibNUUz5W+o48xaECaf9PuNkCB9jtkYrImrsdmt07povJOvSQfDhseoBXxiLwhxOjrZ
SiaZjhwx0cajuiJOlXpiUcQVhJ1t+2sY1wDQ/yF4AO/d7lqfha5xTiO9riHRmsLcoishYmotcrim
MPOzblGKr9II+EeHkm1j8pyH9L7lZIWybIszg5VHqdtFuy2lctp2/Z0lcSZ5FDUSRaAWY5qzSKgT
AKg7lqRYsHUdSXUfET2vFNK1aQVBWdHNO32trL0wdE7Sr71A9v2fuw0zgbuM7btH1E9AZ8S8k51S
npIzrfPpu+b1LgetNhlutCa0Rn+YzLmIrSZHs81Q2TfyLj/7lrrBsmUKi91d2j1qLcSSrBdhPUnO
xpZvu4MWMQdygVh7DWtJcJtT7Ga0FjiWGfW7nZxNqHrbubz6N4kF8UBd/QtnlTfH5iPkhgV8bAHs
ZV+Zz+k8TJJwgHI3iSRkL+Eo6QZsBY6F8IjmAq8Hi6+p8lpT+03cLvMLa4e3lb/9LyMBc3afinL6
gMXCiWhQ41UCwJnv/uKpZC8ZoS0Di3DT2a3QT5uhBmFN6XNR0leoRQRda5qVJuUQFewbt5G+DbD9
txD105Cb/Iix0E2bUWbor59LL/mQaLJjod2m8Sm3wbTHSJMjsO/MoOsOr8t/NbC/peNNFxYnYzz2
ZBIgzzRBGgCHANDZ1q56XU23mWo4coJc5VcQRMJ0AzaupJ8tzZM5n6JsCg880xA4+nHuSEiWtyCF
/J3zViH6RxMiNId+17aJSjt5I5fjhcBkZUlMdVXe15O2uCHYwzgDbCsQilKjObJFuUHShHq5jM9T
tIEpTFzcqdmP0Wgvm0WYi5BpZc6xX7THKR0m5jknH7stiXyzTocOhrDamQuil0BUbremJVDrpyv5
WdZltJ5oZzr8U6lV3cqkLrv6P8ex9osu+u0IhpkN2JBb5olafcR8RJWil4u0Kcd5ZIBky8pWYLLU
82MijoHOhzapbQwOmcRbO2UowHGgq30w3xVmadGwi7rYwrKA4L26hMYzXCehkmWD8eH+HxGJDrh/
FCt1v4nNKaS8dLI9tdpXXVjtExtdB9cbrF/1yNKgBFy6S4u9lC1UurWnldYIwNTw4ZlbWvPwW7Bo
8SGBvPtnJWsoISpG1dIYsd52LkeJ47dGGqaTpMMNHii6HyuAdYENs+ToBgyQ7SUEyjZDBGaPhD0O
yqLguU9aNeFeIyE/Zh7eMd0UVeSsevNMIzFZhhO2LfgCCuupbqdCDvOlUXTqVYLCEogz8rpqZSj6
Utt4/TTecCOP6n9BadPd2pF739kZJXkJOj7XCFtQyRJJOWij5nxdMyWogjUXtBlO8hdMkcm2hVxL
JeuO9CJEaIKOxAMiXw5C+ZDdlD/sfgeMk/tdTrkpr/T3SHhfeanTk17q7LYgRXEQChd07yvBusDF
QkwlbnFzf1SGjTTx2J09KlXss/sgOyFRACSXVBAGqTUJlIqxkqkK2wwSWWtWCDrGTLIsqQVx9/I6
nFnQOXhT44O62xEtHoshJD8VdUG5LR5dM0adUEBmL6wzoJoQSpplk1MARe+M/15qdvJ/T55AkVlP
oVRgnmkKdiIr4ck1sXiDrMP5NCg2aCy3EIf7fOxEAMN2j5Fzm16nJL4rOK4BETCEU9pF4mBF6j7y
zDgfWmbMCND6+ovAh/cu/xHgUso3QdKioz2oh7iIRwkInu82jSeR12RVolCHnondHFqesXPp9BDk
S6EYrvtI5sfb5lGV9GZX4F5Zc3f9G8CDJUrwI5kCQTv1quEzmpJ/BpHl4oEm3hoSiwLGeVuEf0gL
GkAa5pZF/oIQft1TGuxMvdiapWhIWmTjxGFCSnOdVGKpplri7Cgatc1166Ibyk7W7kmkWNmHGC5F
wiHGg8U6NR3bhbVwpmq5cmE9SN/Ddx8n9Gj+27nXmu94ZonNY6X6/d9UcbrvaQVDysUDd+5wrdnv
i5JsnX2bwexb+TgHWP9xmViySVW26NG5ye17MmZDkFTCcCnawM3gCjYiSLN5QcRs91gFOFcCQEn1
QnQzHXYxcA0QtfCrtibFVr+uLdFK4mFXHI0tZ+t9uWmfTW6ItEiNPBr1I58Ae+xwFZts2p/ZKaX7
G3LKU/MtxIaNzJSsmiLb+CACiP0V99afM8/YCRbT2PbA8BP2Ta7rVHOsjCqW40Rdx3kQ1oUQNiz/
dDIz0Z9wzKSD3cr1j3CavMQtMGLd/ZMVFCxqOnGwlXMPL6ZvtFceK2qiB2NdQRT5ZnrVCQEkmONB
FFDwFkaL/MPbrRngbsbv50rjGD6Ew1pQCkGDR4/7X0AAwKXxJQjTNUlKQ8Tqp50qj54i2nshO+s0
8fZ7LLbJiAuXq66S0lvhdpad9uTp428Zfq5URKZyZTjUMLCIwwvwMdhvJg8GrRwQPrJGSn1WBJvK
1OkDiI4wwJKp9eRhbgAUo4tQbFqdR+taNRLKH2JafVRScsVCIeb8roDc5LRPjkgYahEm3LV46r1X
fxy3XkOoBOiZfjBiEwbc3H187+Ec4u6vEL9eOizEL6wEr7TgR3oeJelKiPikM+/yUT4pZpUsUIqk
nwbtAsMUOtjhRyy7y9uuIOzl9JgaCu2vKQfn5PyA2mu6+5T1270R7PJTIcvyQ6YWEPk/75areym9
YmYBb/kxvHw5jky8zSRCg6PBYL4iLka6jn70j8DC9wWBaT07eYqHntburOM0fAWSBQp/cglKSXA2
qH7ZM/O9zzWx0EUmdANhmrPChK8Gaf85Dp+aMIV9kN5/xEZ7rXc9wTK3iC+W4Ap717Qg9O7uEgOZ
UBqLhj2R/HF0fh5Igbgzzkv+gf0S0Im7Zt8/b8KMI7pD2feS3gyVpajE9O/rUEgzOJnhuheqFsNk
FAGVJ6lbZKSfIKXqxuHJMtqZ6pxRQskcnSbvcGcMBhww3RD+EjemXykrGNN6nwd6XGe3AmT4IXMk
mmSGERI+brXphHvHEeiQoqElWM9vL4ih4A/Gm+JTIGU4AIw8GdrsXVlJEdS8nC5QOHtzWj2m8hsr
1LRqe2p+9j8IKam/sldrBWX+I5SvMB1alJrn76YMg7NkszBfcu0gujSnWp+04tpNECLxsDDPhiZI
NQjVpGnxxSly2kZDKvOHM8CPV5xuhYYca3OO60Ou4zyXzkSDebE7feQEoZWkpfGXBgoeqSSCWst4
Z19OXJb0oNW03GZ/hvhJO8GpBxKYa3ZS2D6mdDu82pH0zCpB6rYxzG1y2rg9iMtghz6+RwzGms9L
YbCD09Oh7TxaxZjd1Z/iQ8Su2mFYhA2VdexQ8q8fG20adbMoErqgkJS9/tjjILCSpLCkZcZ5OOji
C1saSac9xENVQckTvu7Pgyl021XAUHe8tvLFGl+6CXJsX11R/Y1xn2M7vFoMnjZFboWajBTV8KFw
C9ItuXkMfosO5CJqJCM1JTZr8WBrE0pOkdlo94dIn0M1Oun1qk3j/Abx9oCwF6zmovg+ti2jRzae
Dg4CZAjswEsufActKy1wKhoQGI0uSgoHhHZ9W62ZerWtcl23qVdGHnM7L7wQzEydR83eYwOs22Xr
rkKIQNT5Ksw55lPZ1V6DQHC5T5VZGu+tAyETR80KtYXtiU3VdvsiKaOI8IlWefRgW3nRFTGOuO/3
Rc4vRaBOJ9wfNPD7q7u/isszdWuwTd88PE3lgHt439STAu4XeAdCFHfz6WjcJth+3HhO8qF9gAmk
sy0Q862Ap6WkdsfhdBC6zit7MKTBbv1oKwC/zRlGupp7dpvOMispAlK35zXKs1tUexaBcrM7ie9G
YwEWgJTwXk6FQSgpZKFXQSZGORgNeWRYPvkByxryLYYppDGq1IJZFx1YM5DY6SHfrqAbFcaYWyW4
bbmB3fUXRiMqzd2L3w2v1z/K8xh32uiRRYNWlGizwHXn5iAjI8ch9YMD9VSmZPEfVfiYBNIrxJ8f
tbT3wSy40G8jizG5Ha6sHAxbiSNHvbAvQ9xAiyJGhSqpMvldlTbQrUpmpiOcUkncLIMBofoKehNF
Y9FJ1lmki5ZYLbPLe06Vka28s1PRaJJC80iNBm6gokdUKqf96ss0AvhTTnly5HWGidZ2JoNJxUOW
zhdWI0Zgw9bNIo8u+ZDLl6YPKqIoXL5Z5g0gqhrDhtv85k59uL0mpTPVWpDyjgC+rWY7OUTFT7hx
edD1JBhkbmEC4kkQBLqFcJBJn803rw/NbuuLrmbPGmHA4rOP0lnrN3UuP885CvkRixXcYfWBV6/z
GtckIfUqBVv9EIXqeszuKDU7S5Gzd1DDnCdsHIpColYQislEKdaMjJS7hvVoJc5zwD7KpsD1IPt+
/CppN8clWLWUIof8UAbwb8G8FETu/1hXJY7qf6toAIBIeKCoSHdVazWcWa9jHeKIpfXyDhtSsmzl
W1Sr3ZQF/bESyTdF2UcL61ap5Oy36/MbTrnLPfisEmn7pWaJDmynEAHOjnQSJVFtQ52PXz8QWUgU
8V/bHo5StiTcn5xgc+mfVARNbkJ8eyij0gYsoaKyBLV4Vc09Q19eJNGD5SaHXWBnnJaQ3ZSD72gv
4DQxrYAECZXwHu5j8IFdEWj7psrIVSbkl7XUCLVStk8GZBF1BCvHZ9uHVBTdrwV2vpIcal1U7Btw
lDIIefdovKJnDkQUbV65+geV72uzgxEJ2iCFYJlA5WaWrTGkfx8lQwG+zlC+kLmvFMZYF2FrFqCv
qCS02Uh8rzr8ZATV6mw/3Z8L9jepCVG9mnhAsTz/88oszB4oLQAZ4xJlSzV0rJkG+HE9uOWcf1hJ
5uLkbgaydN18BUSHqZU0QOA92WS+4Lmc+rnc4ZIhtBLuLXXYnEyNE/C/+v6l21UvsIqOLntAEZyr
cVLlx1XFuqAFcHQlFxrUVHdWx1srgQ7m0Z+ofIYAE9rFKtvqRJXDbcrPRzztt5U3i4biJzR9P3gi
znPiV/qX7W7g0CJ0g9mus2oN6KrkS+iV+AQ0KvguqEXWpIMFCXz7bWhOGfceJSqFfl4paZa9wbl4
gcoDX2Z5oTJZrH0gpvJrqiz419Jv7vEPxO2S+rv8uXHB8bK8sW9hcxJxFH2a3lhCQK/mfGAaRwLc
6gPBbff1OCW3Yg/cLcK3ghC1zDCcEU0QnC3NASa4yPG7nxTH02Iib90x/iJKkdSljV0gMPqqDHo2
vp3waYotGVgJ35FYuBWaJeqX9DGluEmLKd+PJ8kaD++WVYyfRZ10wMS5NSFINb2nh8vl6iZnWy46
ehzYJRRgDJzT06QOWn1RoDeHcbZsq0vIJ4jrCs3jzLbcSyg8F6uJjDoOypzRgydssNuSa3TV9Yqb
Xyot7yuTXlxu0blExRokKMXAvWq2xf2iJ7WaIcgELfExQ4BAl7J8rKB5/r1i+i5g+7itnQtD21pf
ImBUEEhixNgkxrqp2GAidf6OQbsZi2QRlC2BwFMyEmRFYi1KlgPYwNB4IfFEAU2c6fr+D0RMnhGz
ngIvyIPBnQFigW4t3vg7Uua6Q8tHR6axxOyP4UrwGEtXWrrPovl8BOEc7tbQpy1fmI/5ZLk9pcaI
9bNKDPPO4UkEydBMVGd80dC3N0LYtPFiwAK6jc9+eVJPxwOsmjgNYWPAxPhldiz15G2l8O94fUqU
YrMclHFVywiio+v22Go6qW3bU8yVNQ1XFV3uzD5X7jqkXx/wiAlNR4eJsVQ9yHpl2ezFwLm/BNSo
3Vj8LI+dVgTZtuUXvw0GDmiq5/tgrWxc9GuP0AClK3zpFpYMFVliVT9geGO6nOeakTqdNDywT0yA
GAQW25OL0/ighaQ0MJPbN4c6OwWVMnhac1y2DX+C2d9u7D4E3q/a6M24OVg9VD/UqnTbFl0lFy+N
pgtscL2i6w5jH3X9Ax7LcLcbEgNWrUNGqwPbFj0UO9xD2+M7Mx2Q2s8ZwznWx4meu9mZAl0tvum7
dzvxYhpI0OXqbdMvzYUmFQM/UF7IMb9k8ZnLrlLMplZ2n/r9KufH2ecPLSbdWBPAge7dkrAiToHC
FtuYuqTguO+jtenR8/YPIlA+Zifdp/MJBoQS8VqVNzDcNJbv2zYYxpZQChE8MDEGbN70EXaSCVRj
5+0VsvcOm5M3kBhUL2qenaDnbC0G/5sjdOClisYpjy23Y4maCPYKf+oIuxeWieveGxJ0lq4iq9Ag
IxYQTMshqSB0DQJZOKGr6+pmuOYL2d4dYCKR9ImpAVx760y/IW9yLBL6QxJGqkGEPtyAoqfvS7Uw
xDdiysrUeDAHZfNnaQiEkyrBDUfp8KityjoAOcPitcLBxVnazw3k263uLMacqmkkM0Mmq72H61fc
awE+tu1zBofqYw+2QE63Jja3fQ3zhe+aFxntdSKsNmP4WYmvGllD059UFMq/zoxKESpbtPMC0JFl
tff3NPh4WebM3HdC0ykz0Xl3ZuQbsgbN76mFgC1dsyvwiLi05En8t4XFe7oXczqZW+rtesptSaQK
opCqAuOLIh6tPtqTpCHr4cB/y44rUJpuTYn8mju1PDBDl9Ht1VeG4CEPQapzMUsU4iqn80N01mNk
D2QJujzV3e2CbF0oe0FX3E1C0a4wY5f7kycw6zzx25shpva/UKCCIFL4ecx1u4dRqoOOTZ8quu6F
wCu3K9z8xrLeiCwuJDeenNNNCw7sGFHBGWYsWw29GDim5SXPvHi4/03gFACG8vFKwD+Sm+MtmPAR
v1+U6w68OFS8pJ2ObvLPh3O4nf4yWCxRtlZnfaE6lQfFOaazCn1ftUPyiyVlBXjdwQj1ajzZC+dZ
ilvcsMJo2gm0viSrp1ieKKLnJFLp+nTm3HoIO1zElveOv/iwNkMOr15ybYo66JbxnkWYDl55oLba
b5TYJUaLY8n/2eqsDuylovf5WTVsbAJ5ByrQ5/RulB2D7yhIkvReIpP879p4hOn9tChiP56WS2q8
i+wfyEwceXtKy5YFbNxeMJEtkjCq+qvNm0hMRdBdkXE5BHyYR11uESX8lFfOa/2qU2i87Qv6c+ij
iYbcEzEGIzUQNl6reU8tuH3hbpBLp9fSKsx9tIpkx3WY+UXj/j9SLkNq3mokKNFQjb4TNR+0WYSj
Ho+ePL2cW83uKZWdSfi/4Uzk2bCZGdrqGrWwUvQjKtvTbV7qW9k3BElZNOa8qdTJcxLhCbBYeCMi
PRLjFY7G9NZNpDS8jNqGFe2M5c9Z5KGB26yA2H2ye7xcOewxAzWnj8A5TwkafhsN3FzKdVZRHM1M
cPwk+m4nQw8qq3etP8+6lbDg+UkXNWWECRYrvaG/sJjm7/8O3Su37JuNUpZsiSW8nY36g7JizMpB
LR7DwLFVntZ3MgUkpt/O8jh/mWeyPO3Nc/v9K1XAbvrwc1kz6uVCEz76QyleYKcktoaTE9Ynz0AN
m0kaNSjMQrreRKHayWBldy6gQnAPHScbaMwk6Kja/i3MYG8AT2uo/dlhzWyaqpr/563kqrf8KD1S
WZqQU9orP9ABWw+eux97faXxIpqJOXaT8x+PYrPvo4/jnlZCxTxyw7pgiId7aEoelsPz5ATRtOZn
IIwIlZaVadQPT+0Yshw9kkrWlrUfpoa/CI1ay1ndA6JvY1LPFlKYU+kZfXt/yJQ8yeDn25fVbLtu
S+uvNLb77Yy5rCCr09wOWVOn3nWJEwmVUC90AW04JIlnzuTux0miYyxcKHvQ0VBhG9L9nzu//x9A
PanE46NaQlxyOtksH2vtVTLielHHE/3tftD2IdXy6RfXL0o6u3ZstV9J8kE8opABtezs6OTyLKdO
HFq9PKlA6oBuTfLeDpDAxoXRBpQzyrrAi8wOQH5QttL/klFZboT6+SvZI6kB4K1f7JxvuCcrVhfy
Pdai7amGmQIOfWtuLvg6LOeC+HYEg5ioQaj+UiLDmIVnqPyq1g4O321aMrClkZESKGi8Qt9vPLsi
vlBKCV175qQYh2/xFu9niu7wqH2cEaPHiMbM1Q7/Daa/RdM+mM99q2l1mHdJGRpRmaRl2rB10/n4
1S95oxGm7j+o5yA5ev+CSafpXy/XHRFlauucGx613JHgy0a6XdoqG3c1c5vHwwt45af2ZivAuQi9
JBtiMMsG+GGWCvrDPe6bma3Gzet0WVHUZZzz6LKlLnEXHa6BawRi3kZ8S4fUcEECkuzOBuCdk1z1
9XsOtQBcC+MA8/68KuzdOYg4O3EoKpLgrSnA30gUQbbU6ESPMpbLk8y8NOMvrRmrlwaQDix4bhNw
FVMi28nk7CUwJABDXpP6MYke7izwulhsovt4RBWBLCVSbEaoI1gsEWmjdfj49W3xJJDOMG2MP0bF
MM1vyGitqPJma5TYM77sXFNrOo7wPxrqg/t8vSNYYXOsz2Q6OjsxR3Kkdi7nzmnACbjvOMmIVf+d
QGfHqKydUGwk0GQLifkt0kgLJnbvh7FEO7zh6mKANNHjcfUQ2PUGcGeYe5kGuVdHIQIMOiHEdUoh
6Cfq+0dDDJbRUB2EYbbMhzXC2S5xTajAHKCSDKf5Cbxe38ss2F4qJpJQMjiFHxba3H9hm0gCkPCC
ccj6zeALSRncJOEhWU7ChAGw0fyo7LazutM5u4HWniBmjLNCysZ+YMMH4x4MF7Dp/1Df3Oby3b7e
+JkK/mhEdweBtAZZTk32/zwYTLAlHEUkryJWgal8R7hrPdQBAp4Q4HG0LYj1+z/7UXvmO2y/3vn/
menbnKVLlTakI7sTn9YpGW501iizISBK6t8rI0BPukvwfQ/+ctZ8W6mi2XZLWUkYn22fV5ZSJrd5
DZ2WbOtI6ScH8e2k8NOKSvxcmPeiFYx4L2JyI9qeKaIDmYouRyLlpNkv0jQSJ503iku3ct7I24dC
2KK8zw/Hh3Rp/fsLWlzv9SeIgqxszmjSGNPJtxVi7umHRNwPFiF/7ZMcwjUIp6zV2plaaP5xwyN/
8mqlnv8scFypgeOerzYR1bo9o4n89yBEp8cb8O9jx6YG4bSNGd49z41Rhk+sjCyB2AO9bUSWNCU3
XZC5c9Pny9w97sRNl/c4Xj41ivLUdebGZpdOCBMdXm/6OFkmNJj6/knRiKew1Be9qnBKIcufBdhV
iloTwo3zqge4+yy5myUezTueehUe4lU0ZFJp3pdFbSMU1JfBoD20rz9ZDEMU84e9k6AfSjiM8ZB6
ilWd/bdgtmyfB2VJjlth1MVzwMS0DSR3bXUoSnr/N/8IyoQt3rQzSEp7sGN/MPAC4GtStktyVnMo
SgXMEw6uagu2XKgxB34vx7YrmG47/SuE9zpAbqmp+r/GAqNgmC0Ek5p2FToJd/PCWHFPhiDXtt0B
YIPwuu+8uTxwoYMJfgB+LmsYnQh+/ZZmSHBq7HzMgQUEwVdXdut154NHVjFA0HIe6nInVZlLNxrp
wzSIEUSV8ZXuSeKl/SHLjR9RNivegaHFZhA+yF/10pCwagSmC36hQ5//BpK2NeAE5EO7N+HZNhK0
L2tyEctx7gviiL/cbosI+xXz5XmZDCdBwdItE7Z8H/0bjlH/NMbZf8pH7cvqHRMMiku6nUlwbSyq
KlYRn2K9NMqrUOGOzEpPlT5J0YeynVIkoSyjGlAjtJDyS0a3YMIojUz1hwpYnB5RWCjGMIEcz7/R
PBERm/YB8Y/0zrgb1UcDW1XYoltWgAtpmWgSet3iyHHvaZAevqxNmjkFyDIfOMbuGHN7wyW4+dzP
GmSA0De/pf/T5axTcZdj/f7hMq7AaVpRoJkSBQNG52k1xpXThULCVXwSEGz2/cRIqKjY/SpVx6rn
Fe79yiJw73CDmNGc5ZptRG/97N0VYc2Dua8ruFdi66pAbj9PZCQPo7oQO11IJdN88C7zNtEe7Gub
9f0g1WuvNJHD+hcY6zjGvT6R2+CAjU+ulbqr7bXPYCNxONzWLBIb+BeMviZjoGpNSI2bvdSleOi+
BhbeafdziFyIEPcmSWYVwcknFg6ENjnw09XVAn+Df7e2Ruz+fkmllOnQTuc5QAk5elp2RP8Ft8lM
/SKWqhL3NAjs9xdqhbqGIn1Ue56uUElElINAyvEmi1FZl6mihEzSh1ZCcSd0JC5tLN39VHTAH/+d
YDtd99mA72H/RoV+gLnbYRgC1EO56Trlm2spK3ajEC8IDYlFnjEdT9addi9iOZinTQUAYnVQw7Yb
JtjwJ3BXKeagyVnbd4+OCXMR2TvrOTw1ieFHToEMcRqhRs7WUqevi67b+gX9BAvbi4ydEPmaUgm9
R6LeHuW6pTj+pRv7/MRssd/s9JzuUwpaGVt4y+fQXbYEg6C7Pxl5NLHn22o5StVqtAPYNb9Nsl9e
cw49MhGZHBnW4Bt9IsAitqBtMbnHYcCYK97ifEAN0wzNumn+FbQHNwuMSIbm5INNrtkSjYY7V8xJ
+yFS16sfPLnN2JyY+cE4NamXid7P4BCPgLlNfnCXKrv6ws5o1+nvLcpsMKF9NZrMCIghMAb93TJQ
IAo6vsumiXGCKnnNqrLA3QLRe08DwrWGFfXAVr7Gc3VYiBbBdxRrmtv0xYLV1tcI+m8h5pwP6oOH
tu23NmGRjEcEQedFnO1Rv3Aszz0VwT3L2myKt9xhZck24ugckhw+6UPCA+l61U+UaHyGG8EKum8h
GU0RzoNXwyLUafuehqz7IbJDF4CiSor6TjTlRC9Gc5g1j+hSLQVOMvPR3fo+OvU9nO74p0YiNFA7
17vru325urYleJ8Zb3vBc546BUHnrNtQ0YYYgK1K7HPfp5Z8AlthEdv7kC8nQDLL2X0IInBpBOty
hpKHtX/X1z3fNbo2pCm4CkkGjXmZYzS47IJbtbFRtJF5tMgL6kNqtUxjM3sBwLxhFBaYjn0TVvny
tbanNsONVCqUrfzRAFhRD/9+PI2G4uFd4V9UgdCscYjlb+vxCBhRDKe+el1Z/Ph5qJzGWRY7pe37
mBkuMTTESBn3Q5ODgLkYYWY/dgvUD+rHDjU42jhaPBH5Uvm9RtoEZUftM8qezu8kKxss8QzvQPng
AJTR8yug6j5m+nEty9y+VQ0fjdSv8aVwTp6UpTxX0mDTvW/qni++gh7Etz6fWsGLezptCnILZ99A
WOLvJIDH3SLkfuW/Ex1JmXHJh7stEqskouDw4t9mICR6IhWY+i1Bi1CAjyWj2C8vAy0aOnbm+Gw/
5NHAINXK0RPcNo9qoK0KLnVcNNuoMMRt4FNDuVHr0zpc5vmHaG+4wUnH3Sys+c/3cpc56DOXvh6t
XTdZxIMTzTO3g+5RBM0eazvnAHybqhI2feHyF21t8v0qliWmI/Uv4BdsGFuO5uzbw/Q1RsR2ixA4
/U5MU8WVhDeIn5zp8q4t7ftwbn9az1kZw6vQMuZDnBzEwTQSF191vHmpxiY5Qa6RaN5ghnLHMInZ
xaoFaK9WOCmDQWKcrwqvJF81e/LLsHCUaU8xh4Qvqlkk0yVympupNX5S3FXGo5vajbNmN/SebTIy
S7YYmgtQ05MJTZMP/opk1ilG607LMOpATD5G/tj0Sl/9TSm4EGx0M4VGhGpgp7iy5o9r+GDVAv+S
QOjhIvMIJ6DPNHInstwtlAly/2S/uJAM3MctKdp/3PQZgxMu/axto98leVhFZmcAoLbM0Zb6NBJz
GRVxfdumbfJ0KzrqZT8nlUYZ5HwuQKGr6FJA0kyBjon/kNZhdjwjG+cbLaEfcgF9D4MGEIaDOpof
R3/bhfe8S/waezsN2JpgpxNMS+AXKogTCFkWQnMEP8oW/kg9oSOowOA1GTM5/iffne/IY1B97l1+
47pRk85iHFsBk7ebSdPrIJV2Z/gExKDSklWwKU7YlN1uGUbdXWFAWQ+Ps9iXTiQTQvMS2H6ZXYjh
CTUpfFVzrvxYbhRusvRKPlbsuMYFuM0MBNFtb4peLDleVnmpjLh6HDUkR6iaMTJGAPrGB7WksgLc
lOiiNAGt0NtvoGLMIuY19ivvXGxkkUQSma0LY3EA9G1Yrmp8QkoOYxlRvVXp2E+CbjxtQSvbXCW0
nRmUOGIijDSDnI7XN3mIWFTE2GfknTBxwlJWvfGB5oD+yeVNnn9jNKn9aMe+fgpkzt8v29hVjKmg
HMMnEdtOy92opf7LNgtBXH8H99M+/vuwHt+Zu+ABNRNEF/SdK7v/uoDfZtUgvrmxSYCu2NpA9W1G
VtsU1MG7G4GF39UjeXPcc0fJawUC5B6iveQ4Pfmt39fLD//86DPMb04sdVfGOPlk9xigo0xt5060
S7o1+FMz7EChKrDJw9huwO2NNcLUC+DOOZAdGduiSbgEjBk2r80PRoBb6fx4ffKN+WBeJ9Da6B4g
rU6znqBI/QmZEMm4S5uPcp91Qs8R/c9G2EKt7oZdzIdG3jL4ScPZJPivhPBJPMW6U2hUj/Vo2xF3
j8In01pGkimqc1TnQ+jrhVR6TFRH/aZ+aE0KAOfKjDP1J+HX0Bryh8ELjztoMAdjk3NMBzahIfMx
RejL9XHWsFCiAYKo3Zf9saxRC+sgcJcAg1VrBY9jG6FW9vz0fv21hH/136fK2iIXulrtmV0Lxm9R
GTwRHgl116qCyesZl+bXM4MxDueZSC8HB1CnerZH5CiAIS8Pei25FJMVvex1QSC24RitI2xT8ABX
dUQUdPow9y7Yi3KQs/02ouSNpLVXu6HeZFD61M1+QwXIFAFbHVEpEgqDyvGcuW+uAThTquyGs3LA
gjG81aCfFUSH/tCGzqAGKtZGPNFBpm1qXIoWssbUCfCArUmt/UM0lEYolqFNDcLeKgiVBrb/6Ms4
9qbOoTBP7qIifqv2IKApn/OUHTaKYu4rdEtLXy8Uk8yX+omz3bjFRMCWkIi2nWnJG3LKrRLylZUU
jN30Hy3tviRSLQVPkgfrfINq/vl99wIGjgxyOxDDerotswt4KpxDTVsfiqHhCO1AOt7Nb4Sbvsj3
HLEQr1w+2XvOHWeiWjMjv/SgQM47Qw2oxywL7RsC0PaOlB7uFjeBOhG9iWd5SEXEff3DvvCwgJjz
8iUauzeDslFYKcBVeiyReKAf+5+inzN48IMqZnDbpT87A77tKgbP8vEMUtmjHMUCSUYT14wD/DPI
xvWnmOV7jcZCFNixuB4fnWZaKkbDShxHFDHsYBc+0q/3FzPKIHBWGRG2xHQfPVLmDa24H+YF5WCq
XSTvrOymlmo6WBUVupa7fhc7pUmPiPxTw7XFA1NtJQYDFLToC/lXaRANNye3KmqHDLM1fc34KSVf
eKW1QJUYmGZBmbMUYE2o1lvP8oqAkZpYfqv+N1T/otybperIMoXQDfWor/U8JRrQLhp8SGdPKf9J
FDUvj5/LevYM48oA8kkXWRbd2k9Bszchs61qowhqRrqhiT/YRou4OL5lpexMEyxRhdTPapqg0QWD
Hov9uI06Re6iEXaVlTyIzug2u5WtXpXd1d6bPAv7kmTp9m8ipCoUX0LCr/6i3S10FG8I1D/9yqHe
684c7HyUW/dRYEKDqTRXz/tHRN/DKJH9SRIMRDIzBsszJYQB/6KqAl4C5cvzhiVaJrEcNrqZ+cnw
qZVz2cFaeM7f5AoaOHZ3pUKLHTMgoZiTZjbxcuW/zzZwUGcqgKk7C34ajE/Z8CHjAqbRZwXt9crq
4kLmjrhOQL3+EhxdnGRptM+UWbq1+Zoet26mjcjJEPCUP8AXn+J0EhCSfwYjHBXBWdwnOwfzOk8K
U+FnuaJKoVCwJ2NhQYYAaEOkSl1saCJQepD6vm7aD3mdP9heS1RF7yEmqRDyIjQvi3EfZVD6QOax
uo98I0TNfRdTzhvvMnElhZtNcWlCpEduHkRMhf8yV4I0v3B4WCPT0tG2JUgGyOCe7K86nwxQYWR7
szyCKv/rE6Pfp5RQT6kpyvgWckXe59NwEHzyguC6RduU8avTMwK72968A4erG5+aQETStmmtklIT
6EErrpMoRgyH+4irP8g9YAHm63AgXMS3pi80rriKUvETo5Z9tGRYHN65QoC7j2dszey9FNR9YKhh
163Nf76EAy8z4qxToRy05L5UBFAXDTcMRB7v7pJivBHQWnjwsp56U2ubBMOnMJBFhEa81MBPscDK
L0PF9dGQcCseo1VwHKwZvxS1JYWg6Dtxd2FtRxuCrjL4rqrSey3EWpBWVBmUbcx6i8Z/4/QcKXQY
pyVa9foHWkkBlQa5h0ZFBZGFNc/KqrBhdLW1ripmCQpab1sxsoVv9WaprtfzvJcqgmfRhtp6Rude
5Gw5t4H2m0QDQB81Axepm1HVvkPi8AFI4CLDo5nUWa7SVZKZpHFBh8P4hj2o5eWyOjL1ARb2U6TA
blbmmEZA9Z2niR0TDfHdk77LGEQJLPH34wF9YoHstB6ADEdTh/z4vcINP8WdghiMuZyWa7SlX+cz
9v91TyKVYca9hLv/YfkXwtOsCYVgIz5pNVkT+IFNwNxb+TNedBbG+wdMDaCjFFe0tuEM/i7xHybw
0y/++RVZLva66DBHCgbV8Oeul4e6nAxKvlNWR97W4arfhSzsPjDp4hxeYznGxrEnetKskZ/aDg+I
TrQdppJT48EuaRcDT4ES9fnpmfW0KI3lVwd/D5jAp9TJhQC3V0n5hEhkuhrj3zkMk5NIuE6mXA4k
GNwYAcwkI+o5bVFRHfs6N6ijNd3vFV927AJScUU3b0SJjRQHzfZrzIezfpYZDlNiPmfez1ciFMQj
feINuFICpX7imH8xDb5MTteBz/0U8+YCXynIZTvvePUNnNTzYf7fNuKBibRd5waCqgL8eKocvvjh
o8WLFd+m3cmw3SkpJL5Poi2kq3coVQz5fAvPHGVbBPrwzpbYTtLo3OnkqmHdGnFRSII1HPfuWGHS
P5Reqh9xzDBzlUcSSiJ+D9aQdIM+pnaT3h0ueELMlm6oSMJeWcaLVlSw2lBjy8hvfPDcr+5a+3My
taEdth7hILCXQEDq3lehiopLwL9lZgBF3138Dp0i4JhyymH+BSXg2KYam/qcg79OtUXvMzSfocp5
JDKV9IF0INZnk5ybHld4L242thkQt65rOSBt5u1EF6ew4Jx6V7nho/LTxWg0bysCDmbn+bSAT8EE
BQE539mYEsTpKL7yYvKebp+sIUJbySV1atR8MrbjINUIXFuez+l1QVJrQBJjA62CAHEDi784HqlV
rfDKNV3gdcyFAYnhD6AEo2Xq87Y2ZiaaAWGmdl9/xp0L2TIr3eFIXnJ/X0Ub5TZdiWLEQOaEEdqp
BAxc8sJAeQsnVf8+f1YOOy15GuwShYxSsm9lDbQ/4M21TpiJctkJC/PsMF54MY1Dz/utzXMMX+YR
pU+Cf3HSXEfOL71PBBv18oJXEIRaLkyv6tBs+lpy1LXM/1/zovJwZk2SQixaIAGcm21Fgr4pL+fk
/iXvpq6lq1dT1eLWi+pCKlmv1s440m3Nxe05iD6FkBbY4F67BaMagxCEE2INEBUe2YqHsQM6FILo
J5R/wE9x/ZVc9tyD9H3dmpVtkStSGlN+Pi9R4TxQM9/S/ENRtp/io4lxqT0ETTF29Lyp1Nsyd9CL
N3nmRYm2R61DZhUs8MwBqtDbzQKYHgSWsnCqllK0MVeUgibLJRfT/B8KUXPU/VZH/UKIXYiLO6G7
RbQUwlpxXh4HS0dPIKKosKggH7uHVup5UGpPOlpe/s34kbr9ULLzleRzmLza/qRmWjfRnbe7zCRs
T++Pn6xwhPWx6kDdhDfq3Sp27WI6hYwzKrRh3uoHi5RKr3WCh1wyc2TVPNrA5My1snyKczFCBsxi
cx3iRCNhkwu2XlmD2ucYPh6on/+YkKxyP0DuEE2EG+UucLuhBt5BCa9J3g9bhjsOaXj7fhnNMYqD
cKeWWy7ovGLVJFuWLAXF9ik5L16dIqazX6W4dx98DXcDjxhI1FU6UbTKVdPRVhn5pwLiowb8ZTGG
E1lBUvaX8OzVEGg1RnOKy4tbD8cljWg2agyyzqs41fdPy+S757bpSB3G0R62LHD83uKygjdrWs28
z9mvWO6bBAw0aecWr1GJsZ7THQTEUEmLsSI0f5X/ALSAjCffY10R2OQP0k3JrORQ/bbaVI2bkFqj
TQ1Sc/xBXe7avrCBNSafSb247zB7VJoI4sQYokU2fiEidDnWYzQaQc0QzYEAczvAaHpilox9PheV
b7+CZw4jFvnoqJ1Q7buT9w40EBamre40UUBsqSx0tXh4Zv3ZU2HcIWfEkGXQVFREFgwbGjdsnGk1
7oBC3mv4kO4NKXg6cz0IiASkD8nmg1nezT/eA6pizDf5rUbO5ZQwkDAde5OsD2Q4Ov5dsg+Cy4oe
UaXzPYXGAQpJOUWfKrR51E4Uj0R32RCAbR8wYQdcONUS5x05SO+w0kXA4BCEY5W6T9+CeVJn3mag
SG0FLbuHe6V3WFY9o+o+kiI0FWfloeaofDzdE1F8C21P7A+afHm58UaihYkxeTkOUqDMN4TOA3d7
uxnhRbH7Ibc2HZmpjlIBvWwhFmbe5yfCgeIu453nLzWLAPppScI1au8LvMi57g99MK6zym/jHIgS
62TBX9uLtCbO7VyndWxP+y0dPIFv1DUJaLEGtgs0pa0ifEYmBPhQ3iOWMFv+LWTRjSt4x/9b+0T4
tQx2a5mXdAG5Xku/Wn1MZ60DIlxXscnD9MtXf87ATVdCIVkz3ZbpVK4sbc7Iq04fJ0cvIRODyV77
Ta9zuYheKqGa9HplV7LLCQI1e1mIIu7wHJHiA1jHy1tHRP1LMdCh8EdsUBrdVGfRLsw425ylE72G
LrGr30oqatu70aVERF/wpYX8ydlNaysVRNMA3PsW3h9YjGzJJgaAlKjKIydBWehk8qwefWkc5FQS
yZr1L3YFX7+2OUukRw+j6eykH8/pPp+xnC3NTYuBssK/fJPwmJOfn+Sgxndp7xOaujV7qOpEG20t
mz53urpmKpzJH+C+xzJVnLN7i//SxzH5oDxiyEq2d54XyQu3WVnD5XGIFWCjZK4+zmjiVdnOqlf7
9bN9SY1nt8iSF28OF8FpH1TVZYwN+kCr9mVgOfksv3VwbucegHE6t3VT9W4Kv3xzXr63BkbOMphu
1aB1vsjpRtget2BZx7K+m4/RMnUORy+SwhEuDvqfA645F0dJ1eiIDNCfU1/GTgLYkWRa6WLGH/b8
FkeYySYUi+nK3GKwNeZPQdEazx3BybEJLpyC5r7/U2cSScM0F0vQlEBUjGoUzROpZS3Wd1UXsvRG
gscZc/ZXECj8MX62v8LGWHlNtPTppBN0quna7qGyWfRormyVBNQgs6BOTWwUY2xxErixeKS3hfPl
nYmbnMtRGtz5V8y+FLN6IGBkvmn7CUKbN/mECGpn5cqEZoGtS6F6A4XVZaWbQT6TS/vVAkaJVowa
f11H/F5KwXbN7GvOVynRpRybX2FQpMGJPSH6wpf9cDCNJWGxFG23976/BzoqhFCNXU/Qyw4rRe0d
7EwG7Zqju5Zn8YC/yS/4+jbgkTnuBP0k5C4cR8a76AAEZq0tdGbCfzhn+p1kLYs5W3Z0qMJ609tv
rqo5GcKtZTLuqXD3UhHJ7Baw8a54F+tAwEfU1fCQCGPJNFxxSVVxyrQU9zgw/76yf1DUeNTUKWKw
GtawLKl8U3XeLH+yhGgvID14MVZgStGPk4UZnvjJ8H0cj0Ulz4uKxR8z1A/FHkHYY0SukQAl1m1Y
wJnOuR18TTWBdrdQ384HzxM9YcXh5wsSe+b/j1SPOkXrMTHD/ldJe6r7RWoO//HRn7vm2ME7mXt9
xowlX2pVCLIlatAXJjDXW928/Y59xtUGcyjRW621Wbjy27Raa3NkUVDZFZ7AV+VC8M8egnVeSJ4E
S+/8fJ0aFsynuX+8aFNlU043LWrt3RsLtKXie1pjhpFCKfbmc6B/yuFUIRFccRmBxBTDGQ1Gzw+J
9m9zqcTfpLQFb3iHWZavvXe12dr1BMYGyX2hqeVJ1UAzfm9XRNPtU+cj6EAiiRwGY4TOQ3wfkrS1
nwctNgGfxy2Msiw6pvpSK19UOA14Zc0hgD3IOG+zkUfWYKoWE/K4PeZZNtLGsZ9A/ekBFz3wPupV
Zn5KlxzQX+jSSyHiMKZHPrD5D6zYoCBWAOkH4tLFpJpRU3n3RM+czf7++JB/IB9LgAip0mpTkcwg
6DpTkZat61jLEUcs/QqJ73m3Vvlvevy9+5BFqr1EQbMMKeJLp0bppyPQ4lKOCk7SzYQ8DVPbmf/z
oOFskGyiKUX6hYAhuxvY8/K7HrbflCr4kT/ja+lfXVFzoSj//jrc2Ky2KI0bO6j8V2mZbGaPpQQl
SicQ9FUqUDhJCWyHdtyP/HNQZMRxlnbijz1N5vGZBbTSQBZsg8vC5dtFpDDmfbJCWhNKckOP20Fe
129vLmisK1AsIIRWWOBbjqsDH/DfugH1a0cAajR5NEfis89gENQJapoStjDOAk62fZvUELc0+xg2
SOOJsSDw/zoEti73qfTxC1KxFyeLAceDM0Zh9jySPiFDXo4Abkrw5MuMaRViu7bmGNS+nEWcYlXU
/W+2vmKaSO+fULF0Y4ggzXYaeO+3FfRRLNA/i05OgUw6MusUL/P9bhb2cyVHEZ9fFBqTFPf2JA5M
wUbqfJzphNDbERDksxJlmKfP6XuNlXvCoFiiQwbI9HKSzA8Zc/wCs11FHKNuEo+Fosx9wQXCyPlg
tuMs+ygy8UXsP2xSOH7msXoJaXLnPItdHM6aiBJ6WwJcMfjAoQS1E/0JrtbSdrS45FU3yauqfdXL
jNl2J80O8YnP35/j1F0/u1uQPm+SvxsQvVhZX3Ct7dwEP+LgKfNaWb2EojMrtxj/TqdU2eWNZXGP
3P4ae9HLbHPjNUqTxIONzWc6BNqNjzFWntvpbPbLh6xf53NaK3p2gfFuJykY2aPsv3GFYVLQaEfd
R9w0Kxv4y5zQtF/tT89cYroz65NLIUG7jE8TUp4/J2uFjDdXaX5Vg7Sq2Mlzt3Uh8t72XIkFwiUr
2quNu9Qtm2QP4HxwXOhVsNj0LqFvkJIsKMO2yVF4uVz5zQPpgxFBQKiYbyHBJTHOwlM5KWI7FXui
uriz/sPyimeUQMkXUDLp81Tm05cbdBn6rTETtQTJGBANUACWjySHlx+nCVwsVyWLyISBhS9lCZds
+axdD4UtMQpFni/lseqy+qyisWwIL3purWzW3zuiQmRejOZkw0bTC5XKS0TSeYXNOl0MUB3wMRFY
PcEYC4/P1+6nk1QnXiVCN625Y9bNrvViUe7x67K2UOdXEnwwTapqP9+JWWP4N5bS4l85i7Cpawds
/1uI/2zPK40kCOo40Y4AV8fxQspdNmi84eqSdYsUFFnJFqjdGQd5Ck6KfEZ7Bsx9FJNgLGup2GQQ
k2VXuOV3d7odtUlKvD9MX5vzn0Eg0krUoNlpPb10eg6DfDbxgmXoyACRT4J5VJqQfCZmJtKilq7I
DX9RBcOELo2MUxzEKl07ZVeZ4Z0XjdT9k2ISB96/VaQXIzYs8zhBNyK2t9isitu5E33eX6T5hA9A
jAcIMG1qMFxsTJTjiqD8vqLiUU9ai9T9yqnG5CmOuL3BVoOhVHMdmkssxnCdfV0tNPqDThJ/h2zs
le3QayHJPjj4EY4IAJSG2nW+rA/TgvKwanvcfGG/tcdbjuPODiLrwXHVUzP0o4RlLp0qEOHuKqdz
rjIwoQ6zonnbuVDnbWyv0DS6QDwS09KExp3XwUrNJIMEE0DBLlk41jhG6EQCr7FaUl1+0giOcI5I
Y0kiCeKJpf+Hee3qe2Q7xUpsMkvkdXS3xXByuEc7OsDjZG8Ip60d121GDGwqSCgJy6avr2+4f6jW
JalGWcETRmFbm8D7e5MDhr7EYlmiJPC4aGbfvBvzxZsEgh2zLh+L//JxwGRvOJYbCmvS54WneZhT
nGxffxzbfl8Me/DmqoL8r7Wy0pXwTAbs8LvOcQKvfqNVIh2nS+P1lCxtGFIoOnFzYyXKp/Bd4rCZ
y3rRtLp8SF60fAGZmLuh0HMYUQzqNJ0PBg+r0K0bsB4HpD5dHZkhGml2qTSzYSmC5DQaupPK/xNm
p5oCRQxIHnGc4w9lipILrHDoSCMmThjnVayu2yXxY8+6oNiyNkfRiqIKixQ9MZYBlxcIXEP33IB6
LlFeKf8ua+ydHPheQ5V0gBYfbYkqXUeSz6qK/T5m+hrckcukqAgxvkmM+DuNm8a5FTFjFav5ygnR
7W8wLMS4I5vu+HKwoF3gzYRlM0O58lQyo2LPE4QYicS+GJGpR01Rd4xDETjqJzCy51QqPohYfz/2
9GiZLOK3PE/2LZ+xmGMRETq5BV9hYd3L6mvT2zlnpB2yZBC+yVC3/960S4PD9IjAhHO6kw2hwUSf
5XUt2PGF1PWnvWfF84dWrhn5LcEXd52aNtpa7VDxNvVXVc6r5f4bghg1BOdOOi63LqapJ77PCKpW
2Z/2rPg5xUbgS9IrfrzpczSSAsOGXs/UXBuCdbUnffr6U7eUsAubZl6k4SciZXRC+rckjP9LAUkl
tdEdpKduDMYM1/IgQG4SaD8x3+JxAGKZHwKuwf138qk6mSYhhcsCrT5scQfTp89WVrXveYzMvnzi
kdhxTr4ci0m/O7peAXJ71IZLfnneKbtYFG1AnM3qNkiX4FQ9mmy3tqgEEq1fr7OKu2X9bWSvIR1h
I/GwDyn+BeagphBgqUc17brKTfdCLGfdDDflT8OUuCnv2VYCoXNMiSpOAJsvy1rGZ+r4qF3wz8rV
jLxEOyVOInCJ2/5/2KRGcbeuZCdsJH6fhhh+qSwePat7XQQNf3Xhechikl1lWmM6i+Ns/kEf7/WW
N/OsLRJP98SexjDA7D+rVyZH+l3pKpT11YrTd+j+raOQQ6A8tel3dDPm9u18VHYw5/dWkvkXbgzh
UnlSRSARvuDb72k1954coG5p+Dafa/M7TYvdRm1fl7p8UlP63VEFccmTHrbeyXRq57Zg+THf9PEc
w6E9i5lprZt0oxy79I2l/jY184nYQKS/v7Zok9j+dHHayHv2rsxlEOyjAiuNL+UYSW509GCok814
ZWe8RojnXqSvm7oH3xk/PE9wZn+fgrTRXWe2AaicLAA441p9thYS7Y++H+Fb2mV1nMCVz6a+gE22
nVwtq4XCUU9FoBZXEd3cuFsAulEtBTj/pf/Nmi6RVKRa+8PZs0tXkJrzFHStMDFsr0dceaoqbhHy
IOvHzxRR9MTNb7xiwjyuZeQSwYxsvIcYlbhXYOuAiolMfiybBUbzg7YdhTxAlV4+9kbQ5iMlSAhD
TVG4yxHUcLH9dqgZgVTH6WvQ845fGanM4Gp3sB9yqCyKCdQoYE2sldLWUuhhDBHB/QrD9SkIDgh7
1uNOS3Sg1LIrkGyddN+2txOd84MpD9JkNLBaKVRa67X5hgelq+9FdSXXgjJDXz1ujlnFgsuU30ku
r42Mpx/pTN3HU34AS09XW33KBM7RqUM+PgSstr63e0HdG9l5aKCIQnLpERhXf3LHAGLVdVON85tA
h8zHgtd3/jh+WSb36WZHB38k0BmXGmPAANdJCYMAfGZt9tBnOd+eH5f5r2SlWqFwhjjazUpNjkdb
5CB4RvoP32IJidufp3gIoZ3alQjKCOWmwVeGFUSw/RmmXiEgzjBFhh7W/IeF3M8gzAIoYV9IqEdN
rTAU22ZHfJJMql8luGSG5C5j9nfckd4qBCZ+oAXO11oOUordArbiWc3DHzOxLLd3ClAgX+AP9XTY
vQtQWVq/IegYNQxSfsQuj3sK1OVbgMbjOyEbVoa9XEIRqiIFXnSxZeVxh3RnzxiFaxg08vhLo3pc
GJHShKCx5IJgklxt0yNBe7TxkE1Av/C+bv6pfvtvtpBhfTJAkz1QG8NKzZHx7ST7GeL9yO7KgNZU
qTE4jc79KsfHYEuS/ghVp2u7bZvOR1fW8t+els4zj+/mZRePJFdivTzUWakyvWCV05+U3NLPDbCQ
AMhyWS4+YqXjh04elXNvbP2cc/HsKMFkbPL5q0M1WXlLnN385Lnb9eQ064xO2sE/X0hyzIg/PTqv
2dweiqfVzDSbjM77AfW71EqW8QONyCfFEvjwuaMaLB4dzwC1s8IW63jc45wIo4KGOxwZNsVfGiPG
ASVY9UUVU2FtIXUMywGU5yPZYj+fisdi8GwUs9Onh2mTaTk1izVwlF6tXcdOA4iVqswZ0L8V5z2E
uOhuOsMGKxHhY/7pML3FYfwSAyOFnZWCohYkI0iuh53se+3z7GTUCzBUyqWrRQoryeP1/veG8hYo
+Ngd55o+jjBq0xW4XB++kpJW2aU/17dDWW5edgwU1riTAkQYupZy3EnmKsIcOMOXdj584vnbftrm
eYHmW3mMbz12qZoAwSTRHbhJ/RAkvuwAdnQdrpmpfZbfSHQnK0WqLUiWhxCgxFy+O4m8XqmW6AqE
1GFa2+jeEB4caLhRyqEf8zQno9x13iOIcewqrdzi3NQfnk7oS1eMup06k9FtC1IFwikqQ2TAnSix
+sG0Zg6fYmBRjQzuN+ntkV9iWnh6+5ayQ9zrkOR7q8nu9xVL2tS7/hmuHk4zFtSeAoRKpduAgZkj
fXln1AHluyyUmkvy54HrkdN9St5XXc3REmvSQQPwsAOgx08YPi3OT/o6PrzYpgflPEFPR8uGRrZ2
eQ+7lQ237v1nv3Ql9YbOJYx/jT32KYFKbV4rvyoscikklPdBQEoHdFNAcUvsdIduLFa7EAq0vAte
4OkP1uAL8s8ikhgbxoHfYXd4IBpqQZscDyriLfacYD5rRr4DvEnjpB2vp3HovMsIltwg86l8Y3ET
Pdl4eIfUR4rp+sntOJIajJQfNwIDk7kEm4bmrhthO8MaXEq9BLHyBrhOA+/DOJzhJE+STQipv3om
dtAc4skvLDMx9L99cVQ9CfRk1aS0r3egJX5OXxcHbTCBlLCko45+s0111dCTnG4LeMtJxP1KsmeC
8GBhC59QeMiuBI7pWdh5VgufJTuuwb5g1uk55a4ihU+jXzCOby4sTDkQog5bSqxSJMplNp6ZBPtv
A930A4mGc7QP4hNBOLd+byvEiRYFNxbWkQtzpDhuNut/f7LWsxWpyLlxxNVAUTNH4MBQfx2HSS+x
iG0wNunWb4n73OrSjC1yz33BLDP5eDO2/8nq/GcBUjUFiXbBx6I2MTYdLkq526Q6Xhm75NbBCeC3
ooOgd+wJO7CwLIYOQiFJnAiJeJqQl6RlibwQWWsBItezV09qIMVZ4ZL0FOG0jER/PpGxjfeigeMe
oUS6HnGSPF7boFKYi1Q+KAv72x2KS6IGDLTvDP5IlzD/tmb+yJhlnobfvW9JFHUpiA2JA20i1qNr
Eia9ImnJjsFQampxnBI1tmqXE68xP/qyouFWqOmoOsT2Gls4ZmTCxIJdODbeP5fiHGbLapaRRRrd
6NJAaPWgu6EuJ3L0CAGgp9uXsPOHLBZjK8+Ev7Wb8Se/jZpkDRAKs5TXExZNjsGLOr4ZTZK3Ep49
ySwc/ayAYNQNJFpVvw8iNk3em3ZARlDDzEWv5BRij0VTiVOtuTyMFN69bpGBcwpW5+zvh29ULXOb
fB4zuw4YyLARrpb+IaWW5S7bFXIscacZJ1dyLlUOTRuk7f0iU6PpMMwBjvESMSs6JX1ydyY11JOz
CwlmXwLrKYfHDFutg+R5HY/i6s6eqByCLDXnX1E/WtNDAWUJsmd3MCtMOS986DaOetXyrq+WTvmw
co9etzPCqT9C3fdcE/H21RJMjjTNnrgdsskTufvWC56R/+V6o+Zz7AHLjIB8mP2pTCU8t3MCXF9p
GUIKMFhPCqMQ6q/p9nwDlTNqs9Wz+qBTfHtgJRE+nR9jkNmVTER4cj4+WtA1fA1saWaZbj0QnbN4
sJY9Md2tBOXArJr+a7/17LBq1rsnkR4djx03rkS5LL3Oi1LvaJrc76iKuVwgrQBqcCDUxW96i4p2
HLX2T8NRlN8knW04pHA6ghQV5jdYBiqswKq59eBr6qP8DvVjzZ0Fatn6qfT1BneBTeFuK6BFEhWk
mmC4PAWhtLbkugjwsl7wlyAC+adFqt1m8xERPs6J6CLgmMur0EqunhmKgvMeSodiOgs8VufYvCWC
3UBwIXvJYqq7im1xep+aPCMIXAYL5cepY9pzKsKsy4jbMyPNhb9FKQt5LNqZH5TdrgT3wShqKEwo
MmAy7wnphPwcEkbAURKI8fAYmpXDgI2Te5hpRiOFcrdoks1lL6H+Q/fEPtWFqGFl96c4fxfTbyGv
8VaWzPVccJnImL/RGfgl+y2ZOnYQBqNiIcy7WJMgL8yPTvDyeZwVZZ8xuNqOHY42t5/cK1Xz2mC1
gByRR/2EqmkPqamYptHUYfBvR9Ria1j9OIO7eOL16jzclTHjb9t+4AOt3rj9PT6z9y2taeMISONg
KIMaxQMHySFsQzCAyZHpXYa8T5ITODo1TK9uI6xwIFAFM5TsMdBWHJAm3+khBcc1O0KL4GRhElsk
F1CsuK9IlB/xxDGPcfMY5O2DSFhPsXX8aLs7PHYMJHLjkEzhCfMAjzTeIfynghSBuVCaIFz+tR2d
GNkNbJ0E1kk2mxC2BLXS8NE7Q30/+toPDENwhz0+NcIdWNX6+hAqga74D0lSxhGEcSHYOFu00ONN
32oa1DkjhynWIui4QAAuLdGjL48O9FcGTbAEwBP1DklOB0W3MANLNvz5mWKORDFz+WPA9R2b0qoF
kAgvGgIlIP5XpnA8ZYqvfoNz+kUZIe92YwLa8UU4VwOMGk2G8nafhQfQH5sArMCuYUBDDoQ9BqgS
blhFVpjZxr0BCXC26soHbKuBDqTHl7nLjOrVu/1e3K8BPEKUxSipqsAm6RCG7JKodtGJOsHCVJcI
EAuCmWJaZHuZEmjnOqU91JSnZjtfx5h3RR8YuuevGeG5+ANDQB+XdHKXjNxY1WK00ZXFBL1fi7Na
jf0acBDItjeaNbI6m6G0JSiAe56K8hC56xuQCTh+p0S62EE79Xve840dr72FDuSahdrpSJEtomhk
GvjEFHpTxVMsrvbsdLnabSz60RQKvIAelFAMFvtUQkowRs0ckbivvxyrcZgLGOvzQvPX5fsmxaUD
yvCWTSoblgtZSZ2Ouis8sHOgqeAXuLjlRKqmmZJKMmmdcqOPZp+oGKWdKqCeIEMNwczaFIAHmRZk
HCRgDl/z4Gpe/5g4ezPATsw+CN4WBy9uEJvtDiNHfAuJTfm2CQEi3gtN6R+aakLPj/87EfC7bhVs
PXObGZEEt4PVxYVkulECWjWect0RBlI5LpFTZCLmddCHZ/DT5236yPBVzop4oZy3DFCAiQaS/4ob
vrz1xKC4uvFg96An9ZBtahl3UbEnnNER7HkutEVKMpJ5LJ6NUSM3SFKR9LJM1rcXguG7F28jN21q
3mQxI6px7F3oTF8xF2Z8W74o6HwDCM6ZaEpPVsFNfpfih1/5Wvd7nsHJNHScFDm3PIES9Nx9FfF5
MHp/UbHoW7+IOT+2EcUN9twEP5VlaMdHWl22yIjG+5m6i/sQe8ezEuUKoe8A0OOVHo9tx5SXxfo4
3iOYcJaIlJQdDMcAOYMa+UwWje528hWcLCRCQNUjCiWXTAEVcn+9uJ7OgrapCvW099ol9obG+Lfa
W+VHkNHIJxOFPPI8JD53V2w8ADgkbNCTzzRjtRJB1K2Il5gisLGC7PX6c2WA7ULsb2VyeEqlYrOq
Zup+r2ejCohFHS1ZDmJrFKDwday7brVUqpAvCp7x0XUj0v5AHoDDrIIWI4yo7Ixv+Gy4cU4xc4Z3
YCh9thwA2d4Qctq+chcwqbZmrFoGsxcM10j7fLaChyWvqmlyyhDb0P/7dXi0846gUNE1q8toiGG1
E5VYECSLTNAbLgZJDXmcE/sFUlsj6KO/b4i2CKsmyJzRgTEg+4TR/lbwY0O3NkJAetbZUScwL+6G
qjKYJm/FOIbtH8DN/TWKKvlf2BU6k/dgmkF2X4/Qyl6I72Gc6Pj6xpqrm6BYIuKLY2maeyB02cgw
FeUND/DjsBiAOw+9j1N9/ODn1Zc+p001Bn02RG5ZtfVql0YYqjHwogYj1Ateep2defhTLs1/jlHQ
Nk/1DnU9j9QrCVa3X/hd7yyS3+TDS9VBufzrlRHfAlLP1jXPOIHTHM9jmBRXyL2J1w7HQGxovpQL
2HRXotT3ZRKRAPmPeoabxKkDh1Bh4XBdXfuKEA+N7hhQHSrWfycpkYK0Wz1dz4TQ5IMrOJ2PSAeu
zcqkDhUG0P9bn9MlX57D5noT3iHOFdANNYdWJyakQvBL1IwpPxOeJqA7goHs1LpBadmQ7hecysyA
jz6nADq8dYG8k26anAyjw7mtsmlBXdSaQmK55IVXL8LKYdxfZCF6hRZaqYbqRNCilA2t1Fi3LQTJ
Gn6RS/5BbHxBb6Bbow2n+agCXKG+9Q0Er/6+xZlKQAtqoeV1IretHr/71lBypxIvgzfAaI/RqkA2
gw2v3OufD4fwx1LMWJnP6REwA247dApQsDIAiBLyHplF/aO7JWgeya+mHotYa3zEjFWaohK1DaeG
dB7C3Pix9859zru7rv/NoFgv3DY5k0nYYahykzJSTxG1AVV0iH9dyyWKExDp2TMFQJybmul26jva
Vx40MP3p8G1MzRBtcvxwaTdGF0H3HKT0dfXYPBiCQKIRWcgA2WHHGK3onVcUbo1d6/mo7MGWu6OA
SNk0vnEtE2eLf9puTzDyOhXIhv0bDpqhbNUSQ3Da/mfTOSuH11be4M0dU1HkbLykn5a/Fe1goDFi
MQJkH8Q12tAiL4f7pa5nnrNVLOyHztVDhT4knQFKgkfT9xZQvQTUO2LqdXR6tT9NQszdTgaMe4VD
Pzea60CPI0SR5dKPYcdCPAHZsiTToOXW15VRX1BxkDydohLVEDfN+Y2ul85RC8vfznS/9B8LkE4x
M76HKnM0hqkBoN1IMrjGJ4BJuL9mGs+YxzJqZ70xLfMpO7bzr2Q6WRp2XL0zZALyeLL8hWYUZkA2
uow3heHpeEkFMu465EyukNbkiILvIq1j44rezr/JwOtf8pS3P4ci76Nbeo/vX449gpnKABnJughE
crzJ7AtDF2pYw7LyuOcVnSTvzBHFpr0+RLK2k2/f9o2RTe1vVferZ6bMEWyVcPzfjZpHugSDLrni
LJXtssA7sAeKt5c4Wuf4Hbg52uXGVNqMKF2IHUf32PetThAOezxCyePHkRRu6T21pFBd5QErOT+Q
VxSU2Y8vF1+iGatKwyhdL3InB+w2hriGs5wUu+TnVRLTRDEa0K3rmMDFTlZtZiyI1sd28XT+A6Uk
kP6apnAZXE1vAQth8XGI5zRZfQ12Qlc2L4p910Pz9hbME5IbDhFgEu41NrEOmhWuVRpqd1F3nQ31
1bgVYjOqdyN1E2YsicW8Vbo4B5LvK1mSSnqRPmwpUS7ImnLNXsyE+RulhcEeuGGXshzNyEgPjz6H
EP0530Y70p+By/WxSmymo/m6AkIu6itYVlVQl/p6EVEHJ9dG9x99drazhhKnYpgJmlbAAfz/sn96
ONlAflgVcXVqczUt7eAVcv/VNuClO/MyXD5dfMf3+qYOEw1kVVfFYnx7jL271t/yYKZK2KgQpgK+
q0Ui+VpsfWZcL6tfLvR0WjaCoAX414N1ELfgvhqN1dqVJwoM2H/6AMcl89e3Sh4/yzxX+BK5igR6
1gJwnePjbA7qtGwJS9xvp3+GkLyQi5dpET7T+3QGyeJFwRArazBSvBW4u+uEKtx5PBMW8ovsBGid
3j/DVHekZEcl9mIuLnf4QvOisTOot/2W3WFCNlQr8Oe2xkBNQ9v7OpIaDdt+bh6tLTc8HBu8GcoY
UMi/oF+U19LCAMoHXl5vTZIa8egQcXsV+cTmy0pwJVJePFLrM9XkTA1Uhd5FTco6BEIfOTnVVK93
hyPQetz/EZ0TdZmc2l6C3gXMbkivcT1vAalHGWiNkOss7rsuSUDvYz5+6ziEbBrPI3mLkQN/zNHi
z7OSHQpMvOZ4fZ1FSDvnizxFXtdKSKThY/Qnoys5VGNhYQr3b6vpB6aQGdsKY4g5vApIOGYAWicl
uWiLHv5vUP7tK+NZ6HqXcbF2BsJOlGKd4chgHztOpk1E0U/JeFGjC8iknRc6RC33eHvsvJcQWT2h
EgswZuzJPZZYjmJa0aRdYAlWj2ysAs3uKrRR+RhHynTdSkkfkp1F0LtNLemKS2bFtyaDt0wXuihJ
ItufaAKC29Y8DXsmaDnXmN5XAbRMDCMn2ecm/DM+Q7HSqnInUxGvfxXxtX0VStcO3j64Mf7sha4i
MNg+ck9XYF5FfeAJJxdDwqtjkq8NyIx7osVE5fasXFGv6zsdAEr8QK84x+i17J5SbVRbfu/2/NkZ
fTUgSRybmJDTDOMnb/sTI3556/DIT/FfKZOA1sEXgdAdbDXaHGfvCGwoNJ5skddEQGbUa5/1Wmgz
I2L6EDeWK2/CmbicbaEqr+SMVPj6TbYfRmWeDnFZXdCkAxEi7YVmt34iNZlGW/5azclLU9AwG9tL
VQo230pdBihp2wr9W1eQoEBnrn3E/VEvyGYHFt569UK5HsGLr9pTsS180yW+sCirxHN/88129fsn
gKPQsZhB8dMoDHuRDii+ljNr6I3/aVp0mWghWCkN36h47K3ZBaRJjVhCW8qbL/R4Aoketkb3YQca
+ciK7le7W5y3LlE0TFHvFgH8NIIWl9ys1gKtnp/tcMrqFdVC8Z8GGXBilh9tVuthxETUr0AWc0nd
Knkp+Ml5uggXPXXsqjhzxzad3bgh8azDWpc7UuVIqIAsfhbECJo+fQm5fivSv9/qcAiWg+7I3/78
eTwz+lxK2iyEHAK7cKJpkbJ5zSvh34839DUw5zvD7oG49ZjynnK49wRUy/teGv6Fn3rKWQURI7Hd
NODcc/jS+a1DeUoXeCMIAEbqWEsFWUf3ee6m4M2m7g5maRatGGTcSPLaQFqDzk32HEdQRhEZtprJ
z5EO9RwjABBSF9LpaCNy4J2X5yTegz3Rp1KgFT4AJaj3CWYMA8O88URHoPUK2RgfGUlkGGPOT+P9
tIsSybau+x/4WSJXN4subnG3gIq1PHN3eCZ7LjvPhc7fXBA67laIUl3uzNOclpZOGZE9/wiBrbz4
2CTjpNzS0rddp/DpkVt81aaJDGAoj102dtUgZ58sp/RCCDPrUWm2maGSsCCHndSshn+AmQ5dReY3
omS7Azkw3BYWKMh6Z3YkhTBFXovcm0Rh/tElAfKr5p10dBg0vgkjSHfmvnPX9xumpnDrhLLgYTLC
7unOiBCkfeFeTRARk0RotWsaiGe+LvlhL129g10ORTaPgrgYaqPOnDJJr5n4D5LESQ4pmMeqcuoi
2AF94InobJ91Gyuhy1dgXZj+PuRAZvVfN7WbdoqZ1ugdTAnVuPDLPOe3Wo3Rv/W4bP/Ao0hyWAnM
ypBMpn54T/DuMwnu5oaXMFkY6DuCLxD2Eh64bejZiM8pKO3Kn2tBpUIPDH/lhdvs49yYP0X5v/nH
5OKQlwIoiSPOvGMHoOsnxyBYqx7NVuQQgHdxfb4TsQsMh55IIlN1DSw77+LjwALdhZQ+0Yoxn7pT
jmMJTUEpoTSvJVZEp8MCzJQm8HYrhF439E8GPlJXjOdVfPJMGCE/FZJXTc/Ib16wXDgIjUAAVBIp
kGzl+APGuljpVf/9IT1JkaNg+SnY7UN9WIqKknqYZBk0TVJB1uH2wM2iDhvNwRzjclI8p+fj1OmR
qGru9SZHs15pke8fTH5Mg8khJn64/1ICb5yR3AJyVGFqKQxY7vBlMlumqzE5KKW+zOsH4mNZt4cL
4Lm95lmAsAzrvBCtEv49RHMeHUHBqfJ9Uj2SsNos71QJwgfRzIPfT1T43/ZXybJkHR1pXZ7WcSbr
yPJjwrmH4vhxCM2SqeNLOhqJs4/xyHXhXvUDs3w2g6b1iuc19lcrilT/jyrG5d28V/phDO1sBtSs
IjZ9gFk6HxlB4dGOkOansFop9EYdjIxPNmdRnUce96bFhkXOKsT+9pyWxr7FAGkw9vkaiLEBBbcx
It+9Kfp+DD0KR0nUKB4UYE8daIhsginxal++hcsokSxNNx+Pgn9NGmGlC/EPOr/KVKyTDZEoq4QL
VDuCxThMm25f6mVjzrqyMA4Cfl0urJM266N3MgTECVmVQ41Nm9CbZI+HZk5FGZDey6TZwsR5PHQj
VttBAqfI0aW6/2MOKUbKxuG5faubfSGZ/NPdGfpoti0ILGXvAvygoSWSL/TqX81E38qAtdEpJIxW
kC3qIKgt/DgIvmzRhTxMqx4yC/qBWSyeoJaTU4Pphbu1UfzICHlvHoIoI7of3wTggpNlqJVZQnGT
BNJX3JxG5dmeQv+m9eHn70sVDQ8RCjQpOnR5UROsR2THCjNZK4Pel+jMxRLD4xf7SrpFLIGtq+z5
Jv/wVQcs/SQVx92lJ1Ad+yXfNgxFgEDtAOPG1fqAoi4xTUtvh/PbTJTo/+WQ8IxOU2sK8dtKXV2U
1HV+lavWPjJHpjW/IlNmGNOSZxd4EFOLV4p8Jmz+kJuHyNYK7LF1hFm0h9o6MKDhf+W1K8vqiEls
ambuGBBGUfmtwq+7L7I4hbSKZnKygos1uLeSwgNB1ArF305aWlC6NOvk60DTUNRiJD4UHKGnKLzV
bixWgU79GKPpvQWDfDtVzFB+FW9NELOvvi8iIThxf2EQ1yH7XF8EMqA4ht7y7vcfwbTYTxfFMJ3s
8HXltAs+nyFKEqLuQNE4PxpJQlXG8CFQbhbMFzPi+WepbjJ87ajnB+pvPxkiW3CJiO7v6qt2Jpmz
fCGrxsQgFTOzM9mvBBAYCVGmC274T/d8P/m3tJIDvD9Q5G9CpUXLOIIgHsP7fJJ5fQKoPwJYFr6S
acTecT2pXfBtA2DHC8BfTMfEnTzXQVqXkEET1w/WTINqZ8npVcH1gTjtaWCr5391bTlN9ATtHfgd
0DPymp/zcFp8Dktt9qrg08kJhYmlhnuPQo9IG8LT/G1fefQXLywL31sL0QlUqnEhG3nlIcg+aFB7
omkh2YUzAN14me7u6A7fZY+Wg3qIppbVqOpCVIEIYKLdyW+yFI1LokUWmoEbVqMG/3tDMLPwu28k
NcMnYo9Rcq6OWQFrKkVF0QdMO/T5yH9yUpX0qFdeqTxXvGg1ZQtlwVVPyXpIAS5tsldcLp/CGSgR
iaAO48Pc0IPwQ9WTPzyTewzAMAgBcXGPl6lOr5iBXTBGkofJV5c29IGfUZTZfpTLJs1F8jlM5Rfa
VasEyEyKlDf26eYjUd8GgB0knh9hB6c/YWjjfDvUQVl37SeFPFKvFHkBPDKcEnR0nN376vwSzctj
mGXsZj5sqNBI+wAdACX8HojwkigHiwvC9cJ+6ig3IoBW7wIZqs8hZNJeXRT+voyfSE40byf6p2VY
/CNZZRiZDOasAM0oLJxd0xihxc5YkiRb8ge8Z3dqDH566NHqdeKfWnAeH8UU041BTRjPa/Y2de2h
eoLSOKjEiNqTV8/KI2UVfoc89PtGfkuVuP4QibuPmG4PvenC2DJmvXxOrp3+2IRb9q8y6aLBy43E
kAjtZv158tIXyE4DCmBNXLfV+bCX0YvldhIDlXG+j6xFsWbwqWW3N4F6/FmY7oUMaCaNoTJeXFAg
yzkkxxV9hxmq6PYuqMUtDt1/sqsj531VEYDzRTtz0x/Zyi3+7QUw2IthX16AA2tZhf7+g45davAB
OWYW8uPqW/UAZi3eNK7esir5IgAKG9N7Hb8N/Lk3ZPVpvyrTi1kNmp2ho8RhOiE7WVnru9roGMxL
pIIbEO7EaoaghhIzm6DZCl4t3UlQ7HTpWEjFzn5+cjYDP6RcS0YoDg/VRK47DkYDdKNTYCthX2o9
UwROWBJVYoZuqXx49Is7ps8SDXOw1wHREldW8SNy7N6G2yfT0KhXnY/PH7Vqg3oRkPAwXKLS4SC+
ooYiNVfkx8idt0PsrBjCK1zL3Qy1kFj1VNqMHovg1XwRF6OAzfREVYnYNKq+vg0kqvaRCRF2jpxW
AHlv5VOQxgzL+rECewBcbQOHNRt41IYJNd8HG9Su9sS6p4xZ3+O5lWFOvH2WWeIkD+1T3NLQKLBi
w3wLEnyQe6Jzox/g84N/Kqp8A6FiAYaV4GrvRWpGUpqS+UEtOhOrDh41lhWycVK4b9eyyRW6GmOg
yHyoUGhOdGguMMpg0ULSsRtLnz91xS4Vm2I1rtS32+fsWQ70Zv/qV7ob0lRR8B3l8DlK+/f4mm7S
UCK48nY8NxaHvi30Hmj7Skd4Edm3VCmLRL4Li1ikeNOaVw8DBCYPIv5s+s9QRy/uRWIcd2ZMd4UX
wUPTRIVLThuv3Msk4C3yQZn/n1UzqY7kJ9bfuxaIEZjyugiT5y25L3YrlRoY+gsJDmDFWo5lIN5y
bb4MJd0TRJNPJr0uspD7jad2R/hukUJ4WE/rWuDDKd9IrHqkqZSoghlfybxvcnsuXmuaEydck5BW
r8i0WaKrPaPa9KB0NIxks/mLb2waTYym8wLIh/2oaVxSO6oA+GGMlGRu+vS7QU7xZ2Tae0IhcsrW
FqegYblIAyZUMw8HN0LiUPCE2oPPnEMcbe9zDSmKHgky7zG8O6z0ADAh9s4JTmCSaje7LqmR1AOM
M+1fyV1uArrjnZ/OUBqvscKSZJ0/Nh5kCKNNGk27HbYj9CQ6pUmUrDf950Aihx4Mpaw5GPPD6ZuA
asCFiKc03tTASfKIWvAvRem5LIm6Rzj0CJgEvmYBMVqRHshMI9v6+afeZ4ayGkNveK8X62GNV0/l
RAgo3CJAHp3jO+wFtJ3grEnZeoj++PLH8KGzf29EvXC5TyWltf9Jw4cmVnaYAvhQadXspC67OZiI
pVk+n78o7AsSClOLOkS7j3jQgWW3TYvgj6M9BQGE+ikyRM6mHLWpAW5l2OqtfvgsK+fYNyn1fYuL
RXUYsu2K8Rwf+0fo1vvg6WVeGRo8ojiPNyXul8/ho4kfo1sOHTUS4CH+JFovc+1Fkgw1BmyWsWMS
ExBfRySpCnr4umsey45ytk0CNBDBBXPmhB5OzBFcpfqyUn5RAR/qed4H0OZ532rpfe8D3GmdC3IN
HUyE58gb5RUOCXYgzmS5UeZubYkFbREjubTWUQtu55FZYjUk99q1mPAupOrf6acs6KPSIcN2GOhw
rMRXE4MA7g8LnobiVXC0r2fS58jE8Zu+F366aRJ1kGPl4YXJNAbliKAiFU/woW6Ab9vyNjBt4uxE
dBXyqoBI47vDYVOFHyT936iFYsOtDJ6P1cmkDtlYYNyAzc6rhoMGlo0E5N7FosBXrIF/wNwKTAl+
rlcz/ZwRmiCnwpW8/kwNfU7PXxIBfPy3ful7WatQzbGsvZeOljE1nWdRsCYT+t2qi3L9A4NSQ6Mt
OXlF0t5syL1UpBfkFRK4Imh8sGi/2nDiyAZyRJSSbiZm6heBmDrXnW27f/MVhixifOtAHn6Un4F3
SzqOwBWS9gth03fNMQ+vrBprkxus98UIeE0Q8KboyXvEGktT/qMccqQgSCb3vbeZVLRE1nOXpWBr
40cTtMnLaDBxcaSAVUqhNYmbxR5O9sCH1eUJCW+Tmi4fQpkbnDcM+EYu5h/s6j/2g2iFs9Av4lP7
qSZHw3Suz7SydfkpTSt5Qe7cgW3KfzRIWrLUVx7F5LRCATRPt6ug5jLXagpbE+mP6BP/HmB6zHEa
NwlUlvIg3i4nZDq2dwpsqO+7Td680NIeMkpfI5/Ha14vJAzOVYqmUPKyYsQavgVwH8drypfU/UDZ
19AWuCO7JDtTgZ/gnxZh60FwSgNrRrSTxl/Oz/B05Kb2VaqHb6j8szu6QptYvy0RtkUo8if6uKV1
7gF3tmGXrLsThBQhBff7tMdQf//lyPV7ICVfDu19Oi9e2PLYGRSv0+G0UD+V5OCMPv7BhRpL2fhF
IDVfD3cV3E6n4pZa5CxvUDdQmT/ij8KDfM3zAf+QTyIo8RjxOIkG3rZGSFUSuEg9qrOnYGX1wdq2
o1G/2yWEq3XQYNIfzA3xKmrrokJ7Om6WpPgU4u1ETYhlZQ44kpQNmIighEO7DcW8Q0afbRmf5l8I
72CcfZFmvSThFkghgqlul4WCLRNvoQOWWQIBNbxOclxLJLpmalEOlUx2s0+uPU4S2wBzpTfAN++d
BWVfMaPv2hOlscq8XqVpLGNjHJKNDdfld7FvLZxuSPEg3+Q8v1boXpEhMjz72ZpEyRI0tkY+kmMh
0fL9x/uTlGIPOxz3iXDzO7plZwENRLqpAkhdjdKpmfnrOJ8o6boATotww1W5VPCuWQyULLbAKsXm
dd72qXYGhegP0rmyTcoixRKZAScCEpIISZt5yWmH476Z8+BC8ilWWz8fJphch9nzfKNpBxBzvirU
FQSyn4KK72ykQdp/XBbWpXwWB1ltkLcnj/cCi2djFSUPgepKTEL2ox3GlaskuAEXHtcbjmbFifSc
Az+YaoBELBcCAzssnx0tE1yv14BDOCILLImkAHWw583RG1A7q6YI3LP/KJAisD9xfTdATmA/ZG+v
pimGiPdzmzWhnKZS3EUT664yUs+KiTxmWOnagdgh5kr4Dyzt5g8Te1AxEMgQOc6WhTBvuvaTW9J2
A75LlmGQVpQ9H6ySukvld419i6KdzMws3Xw+VVNh/M8c1NulGluiWxDSmuiRw7PcaakyfdO9hEW9
m9tReVxoroAK8QjMUXtSieXqJoYky4Hg5pL5b9m7UdFoO/TYtjT+f5nKXGzyfG6yryVtXYvyKFZo
La0iFJFsjICEv3LmZHIbWxPkB9BKoQm3gqiZGREe1xrohAsLfajqQxO5UwInsJYh1MuJjAimR7VK
dWM1hOGc6Y5rFj87RTdmwjJwwGPdpH/HprecDDdYBFBOIiu3yvZJad9WL5TYdhjLnN4zApBqHCLB
RBhbWGCq/D7fethjnXYIX2d1nA6BtE4duRxkeCZXwHIXIia2JU5Z3rg5lXc/6s919Ivc9sbYJthg
NIbCU8CiAly/8wyv2ewuz4dxqvtzZv7DO2AIWq7xhZv3+0tC1nRDKf2CBVuFCB2QT+ng050uKYVR
T7lYmULPREhpfcqH8RWWUz9EWu+4oxv6iRedQ7hrNwIqLD74+tp6TRD0mHR4UqbFRS3JDor8J5EC
MGQ1EO+aIHKmezYaMPF7nkGgKQDWqxXCfeiF0BcGZ5DPpYbMKP9qhf1KMRWriwwRbxT4EpxIq8+m
3KHnaOBYM86RQYa0DTg3a1J2d5M0GhCAMXfD75gZu7rhpWZQu73/I1LDuY5sydtIcJ8ksbXNl497
WUNB6BAlKkJdYSN3SORjydxPvbV4PeuQYp6YZWpBFqD8QETbHNRVTB2YUs/HKscJR4znNl3Xtu3n
j1WHzr6QVxaDYdjq/dxDydTVKNixSAuNDp2iuiX1Won08oGGQ8IhuyCq1maU1aMx8MKjCi96C3Bv
hBkndc6VV+/X+YzhvHBbS7s4QPSCA0XD5n9veIbFb9jav77OnarLDElkH2Fy+mOCZC6MhZR3cTaH
DlKHZrHH5429zhEa6I+3+KBmEHY57EK2VTEUtDIGXUBwE5XrTgpaR3Sb812TqONAVQHf+NQDPs7g
TRPb6nztHJCh3ovy86q8fKzcRCp9WlRJ6wrS25jBw+9wfKzXuK0+T22mDg3qWDPC69gsU+lgSgcv
zJWJYiRnB7iWcfhcXILIuj/mQBVnDeiKYHHh4d/24bsfBeYdSL5Bsb6OMOHo+EfI7vP8ILuvmvpW
yrZYPyfC5sbev9IsVaFcl7fVzkaPGorL3DgpbRtSzEuXwrUbPGs66Ilyxf922xYPVnSy6ILsURuX
7BjTw3WXzTh5UHMjBQUwr/HmwEn9cDTeKsyInYX4Oo/9tSJcEM7/0LMyLkAOW29pm7zwNS0QbpPm
wFWhNeel3I+kiPK39UO2rsBv2XxHTmf6b4OjiQSExxA3uR7Z6mVZ1Asc/HL2DSEZpmBuyjigVUxx
yqW3Vc4B+nKXWlGSh8o/52a873UaBomrWbHOxi3lbr12dV+y5G6NExZg5HeWV8WQBmCIc0JBZUil
YILnqQ5GMUsg69K7OiQX5E8ehvJJDTPyWbEDVysqusGq/n4ZfMsTV4C+Ha8v5ZhekFePrQhOe59V
cx2LBs/Yx4yxv8O6QVwJwG4vR2QWaqVJOPIIixbwtRoDiADXXz1VxQpfPlegZByLrcjSwkTwP+8U
M5akUhHqHF8U4KFBZ15doBjFsN2Lf8mwoinKRHerD53TEsaDZDPjp7VB9n9SMqgKdQVsv5jZDRaJ
ZYdtggyWCMikIVQDAzWsHDcWjWZ83o7ccfIT0zsnCdZFz+yyLnvt1M8AI7YX+/OELL1hMYkpfoRh
CMPljqHtNqHx1zdCUvhy5xGOCyABVTw2SabL45CfZ2DUpdtOZP6k2OOub/zvaoGa3jRG2ArL1KaX
7UxJpQQzotfFihroZ2+X70A0LURcxlq+Qen6l9uhuX9YXe8C6U3m9NoiZb10gCC1boPnbxkqZFRI
RiyVnsg7Y3zN3uBE9Pz3Mwz7zEVhGD4jzXuu7gcefwh4mBd5wI0X88sP9sriR3Ypc0csOxVmML1z
KeMXhMWjvIP8zHgbxiqLm9m+s7Sk/EOkrJyY1AXijmDB+mCHwT8TGBG9IGfC3pc8/RHIuo1lF2Y+
1wsDLXZMLraqLETmEhs6A3LeDisba6Pwd+3Z1wCbCMRMXhMHYWgRmRtE3ySXbKpWh5iLtlZGmN6u
oYLrVlplti+OiCtt/pgoLRVkjqGxrakAffGxdzKCaiNKFHjwxCls+BYnF3UBUyb82rRK38GeleAQ
8nD0fhZNbw2R1ojNVnufpmtEG1Pstz0/7qHO0N4eb4+lNwbJLKY7+/muJwOvV5WMn0oWvJt2MkEd
dMYfYAvMfCo3G91BzljR2U4JwLvfOXld8xvjlZJZC8Xm2ZabiLEZo08b0sPOs9+E60oOFROPEKHF
vFhiVSTKuFj/98Gtykx5PgDkLJJ0n7pgk/47oT3TISfn5AVEoW6lCjZij9TkjcyRJNcXIZ/umHGh
RIVKfQhf7UdgWrj8ZkuIDcMOqoFAZy+xPYHYAc0kn7UAeNcrIF6H7/43G0P8YEHAheVDWy0Ubg/N
wLPQiaHLGQxdeZoBEju5cnoXyeTp0Et4zuZdT+5ATlqfAl/09NGPn1qZhsShsi3ukMrf2oMgQmy5
RyzukE7ZrnoxXHA8pnbJdQjF97Gcu4nPZ38ubZH3/iWCknNfgCcyiKwmg2cAZRA9l/Ssn7h1owNZ
oU5IOOzxeAbfv5jeOnOn54tbKIXMccjqoiG65mja4uRv/yEqGhwe/Kx9Q6EGsiQqkTai9NrF9haP
YDAtpok3ICa5xIuMeF8cJRhJDM2ku2VhIEvxujdvQhmBGSVF9NdX67QP1P5C6uODjC8P4z3R2irU
E82z3yXVMUo0c96BCPprxjUMEnx8esUMBmb0MwjylIupjSguAqh0XDuBFVxj3OThCoQ9vO1HeorY
OeVUnnae7OQP/U5D2AspdhicHj9gOlC6oe094JlomktTtiViAKV6wE2UBxQe0oY+qvd4anC/IWqO
puXJf3/GUfNsOufwVEG8D0YGqjjMaXqRYHLPE6a2Ba6o+Nz+31e/WX4VYKcQhaxEDfDWWwNf3FK6
CJIryp4vTVZfqfQL930CkSxMTN4uxPlwN2OuLUohSEEP+xy4MyGtF8KgD72J0BVl+vtUopY/caw3
kH43M+LsA/Y/JXqvgYICJ3huEzfQvzZrW2dUAEMbVMfpIyuxOU62t9yHF3AsbSjCWyCXdblVWJtd
1FT4+3ckBRHFcgbWlvmP4TTJdtBrW0cQjOR/zU2O2kPIMts8r4v26LTdfi4pgmqLyfrTCuyD23gQ
Y047kCBw/I6E2FXIH621oSodgXeA4LIL3agV3xFuRZW/CUpLWoATcuysj6ZNXoo8A0RPBpgjb2fK
7Y+O8WqWlsuZgpEv8DR8D4he5czRziS2KJpA1N58IKhXapkJwLXPSnB5E9Y9MXVfPnPx58vo53eS
AwNDsjdv3iYPRbDvccNBX3yPG6O+qhNdN2qeoyTzlkC7mOLljIXFR+T1V5ovVex/+KA11ZHMt6Nt
rRHWRNhaQa/ivsqJz5LrsXWqf0CWgxOURPminSytUQnvtUgkmAUvfrSYdxOdMDVu3EPk7KqnZkkX
DsLRKm1FcoM8flUDDULZFY2+kZONiLkDCVewDTZIBlbmPGFWQNwP7aiYfClFW6sT632kfSn9Mqhj
nXgc/KJwHY5ulA6pQXRDlkHUw57SvXZxiwbB1NPgJG5rc86KL4kJRz0U+EYJHhPE7FMSiLfJdyQa
SfHlHdEVik0FD0YxAyfUQ+dZ4lSPlN/xlRwZHqTflhINImCdd/8BPdEjYSHH2GIzgepB8+IO5/ZW
ZIXahG6imjMv1i34WCZ5QGxnTPM2ioJ4V9qZnUuAPkCIX2F3x16Te8zQ51VipqEjBZ8+Wd8A1Nw2
oi9tF9WL6CR1zrkkQpKvlqLgg28D/uj3YBjt6UiPfKevd2/7Z+aubSMxE6RWh0VObmxo0TElx1cT
57TtLLybIkDBLs9WUflpOBgjqidNMem9qB1/ATbTcUTaeT/AmEq+9w51OXwL6vFxTX5SnpXXHOX5
mRKBvq6MKtTjoR4Klrx/KG4rM1XzA9nJIrezEsVYmdORQBytVc6LevQBhL+OU7q0rNjfFC6TbMxJ
8OYxZPSKmGzwtvw0Gh2yblSYFKoKtAJMO/sqwfPjdxCQ6rrhPqaajjvvffIhqdEY/gicIHn4PX3I
SDQIe/zDU8GsqYLIPvBOvm2XzFcnHv04N83DMCApu4nkNsv6QHu9cAuySQLqaohF1mKDk2GHPx+f
xaulfVR2Gbn6YJgqA+REV87hAqoBLdKwg6xeVFGiSugXMByyxpT70a4j+ZmZxyAh3GTHShtQL0ai
7JceYcOA8yMpa4spOyWk2Afi7EpV3EdQraaIbo58ek/VkyrwaXkPvta243lRmjq2UbMs2DOCzd2S
u8zMv4i0B94qmEo+Hg0+s4daqCWye1SLIv4scTGisE4Z0seKeOcHbpBQXgu7plTaRfzux1ffVTj/
VGNNoJKCbhsoFVtT9fqtZUTXPSgvV9dEMBocOAWnF4qICe2pgL/kckAHPv4S2iivq2uEW0hLE2W7
ole365TXAnK71cdYp9Qj1FKMA04NMjuqBwrIq4cdK1iiSHg4B8qYuHedSdR/UC/ek4k2tU06ZFR3
QW4LFhEAIYFP/8rVeOWut6JX7R9rnz89OsCnC80PScOS43mRTZyxNKKpBzxHNG/fQrwibhU7yMm/
ZznMt1dT9Lrdcz85sbi6mo9rGGnZaFGM9tkZHNxU/Ot6K/AA3r4q27sTh4R73IuIR/aiwzksjKid
S6AllhW5QPugTr/+p7vNv+P2K/qgvcGX0V1VJCFAQYVtm+3Zxj1hIOKzM2qUzRTknAbfQvqoQgaA
FF2vPmX3KnHXRbFZ/IemwNprqz6ujbiiYTPTACR168YDRnGODF8UP6Qyqd+PQWaOx5YPS3f7Cc/X
n7Cfxmikd4APqQfuYI2MRfqz8RIE8V16WBJu/5dllv6JLYyXBfybBnxjmd2h7GGv31oCJT/QBdke
xBJEcK8t9wgxhhqUBcZgH3cMgpSALnaRBVlO5/KJtqqMmHHQq7d85/Lx0e8o6vLxObe3H4lCvtcd
SWwhZHT+LVeUa1hOaQXve7dcLHdkilhI/mrqZCdEyRTtTpnm2g9JNNTeC6qTM7E1LkzcagUxCHwL
bAgur/h8821jLgkVfFHuQ2shd/BTEjS7MqeuvMakFBJh9bDATPiwVVRLCvgQMP0+qw/beP+UlTFh
FgAGHZK8bCt5mgKzz0yNmjhbPYriqrMEN+/71lJQ8XtIFHeITAjDDe6N6oQllXvFjNfhWqdgEl33
mHTTCzwT4dwZiW4KjkAbdSGJJNty2cLgWreJsbvmbS6n/AZwxRjHyNplxA+/ZBOykmRFKMmFMv9g
dqOBTjzW+iQPRmW1Ib/rwpyZkhadxOzXY/V2hriPFwphyScMmk2g6JhT7TPREcjyRK+RhCkxN8Vc
+lpsQ6s9zZFdLg0qn86DhSCnpckIjRcr5mY8X68DO6l65PyL8EbO9tFMQ7u1u26QFpm66FKgAfxB
L3HViuded/8SLkHlJB4qHb2SXBmWRbu9kLtomIDgfIqDTTS+C6ccwrRP2Lram90eUSYP8jwX004o
Ko8HzqqLoiikrOlb5rTlAqwnrTOEHoBhzhDOg2p57CbQcQKeY6iXWbtmWWLpr5//1vU59Z1uHv5m
lvXA53/T849E9GTwYWIQbYyS6XW9+FIQlhSTSXdKIvO07ly01f4uhVCq3kaUYHe08dpjDiyoL2g5
xD4l4qSjDsxfWRX4xtZObcrT9b0TFloO1B/UkI9NkPZXt++jQmCHz6n3dJF9aRz3oXCtdYPtRdPC
uPaSq9EQnjBFlzcAUajbYm5zgMawvqbB7cCsceFGYln5iKe7cYExCsamGgKhWKV78ODf8VDwK2cC
bIzVduVOHLxO/SoxP0vW/ibIBSfp+ptVOJj8AnvLknNbUiLbUa82nB1N6yAhXwqfkEpX8dBtbZtA
OEbybct/NgU0kAQHYiLv1qrphBSzvSTEtZ+qq88Gc1yJzHj5AEWMB5nzfogAsqlvRM7Fs4Syfj6g
vl3nmJrrFZw7yop6CDiaE0C57r8I7epx4aaLbL559euUwE3iNANAiA/iRkB46rPN7VTcl2a007Rp
tDsqXAMn1Fvmpr6QxgI0rtQJCOjSKPJkEbZEn5c9KxAeNK8OZaaRvqUbwoyLOyWVeY3a9Npx6WHA
gEnklDoHVo1ewFFUGxjvYUaaHi5Xslm2q3K7R8ov31dBYrsqELbmYR+hJNlyLwT8PFLMKw1abSJE
V/ppegMtsQXaTOvYTFAwzYbmk/305B+CnnO33KkCnxRpNV7LS58pOnEXug/z1cVMhHrIO4J7aS1G
nJAhqbhxQHa3uxmJjBpIgHFnXKUH7dELyLhwYGnmLDY6rNsxCMUSECh3QzAzcH3CcAHx1lBv7pgm
362DYo45uJ46Kh7Mojhb5sfcwqe9Bi/zeLZV1+ZkPPOZu2AToOhyb5uucm81NQnOTsaD3WyqM+DQ
S6IOv6MEQS2ttMccrPmWfBYkO6ZuMEYFhWF+4u5K1LxjbMy0c+SAIdrG7KcbbSTEsqbCigmtg+Ha
0rCUzzR+FBWa0Va5HfDGAH+pFaS2mXXVv/LYqg98bGIgr8Nl7JEGlDXiEahjLWFwKxcIBgc1VrvL
V5SG5v+nr6Zoa1WXjNpBGbzITsWSTSU1M4P/7H8fG/3118Rs16ilPFrTWa6XRfBat7ktkA5a0tBD
QNtctaovtMyTUSAo1ITkjF5haGIAKUp6Z6iQv8KsWnOINU0m2pBjaKR8iPcunE9zoyPwTMzVH7+S
F31iJ4Krzgg98OQRVk5T4sHCvsb52x55Sqbl64ijPXy3tVo9KQqG8VuFLmz42wkbpgBxuiUv1GbF
NIJmvwlZZiiPncq6yPmE5zbWxRkaDo2Na6AR8wOcnTV0gifYFhJ4lC1J9U2X5Ef9PTdNwIVDw+jz
BMDO06vRC0c3Qjn/rPI5JHgQ1pKiuuTvY6Yud7gRXGP5a8iDEiNTWPflWpj0vhXopZRHTyNddLq5
ZRt5nms2lw09q8LVNzFLkPjULGN9WwyOekkF3XnqRH0f4T62LA7hsWpQgyzjDqJBc9xO//oldXwW
tpGx88cYD4a3ELD/o4bmJ4iA8dvGRBYbWs1EdSXbZ1O4KNk0buQ4rvNIR6CAZLYGVzuP16CVhNZS
gdJSHo8WdOy90NOHTUO3niaeGecxssUnuLc1VyuNu6o5PY3zg9j7mCTMxSb0P3k15AGQ5V1H8vEJ
HnUcXQHQCnoMrKFdzfiXoyg0JWJvYCav8b68BMzJHRo5Xvb2Yy5O+4jxsCesymgQNcMnsi+FMBRH
Jo9dCvTugq20zwM8H3ys2JyZe2Fe/EtWKyp6lHXuXdg3zPU7nyXA70/fFJV+HpHDmPtbJGsBUJJh
41br8K8vXJAOLDbH+klGhXk1iIXvhZalTa6nl7+IwR4tNyREDu6vnAOd3HIccfBw/Jr5jUKeqNdZ
Puj2/LjlFqXpo5cD+YydTDdCxZDSXNPLjoGlY+QFKKTRtfL/5C1Gz0DIxEfRpCJ9wD1RAyPmvP9q
y1/Ip8/2iLbRjfpx1A0HJmNIDXKTutFtovYzqKOeH8YCiTPtU0GaXCMQpFyzGREC8YUumzOFkr0m
caJcpcArqyCtOyFSRoPGhyDglh/s5jdiq1L75tyJshWvHg+CvD5QG/SqLr7j3+8HdAao63U6ixo3
k959132x7vSpcrJ/UVbz3ava4IeKQBCZzC3jGcXXUa3sFpbCdefRWFsPa6lBnOiysrEcgT1t5q+E
Ksdy1CZv37wUMNATSmZFnWEnWJJrw+C8jaqP38PL/68Dd5qv2UzR02b+ufj5MEhbB96QAvZR1DUL
Psoh0X/py9a0FNadcQpqF2VV1NN7MZgP08KUIieXjq9Z8waP1ph/pZAhP6op5ybgCdAA6T0sMmaA
mPHiX7Oemv3QzWqQcP+FIJ1X7y3Z7YE68xaLqNGluWOw4fuiZvjpr8bvfREjzGXiFyVXOy9iicNm
SsHmEnP22K1dtAWWmL0PFhcPBYITMzMeHwhbI+ClfKJBAcatGgDwC21fbqFWFeJ4qSohR/VL5LB9
M0lZru37CZoczehfj0f23sOQ9MsJ13UbgSPhLqzncNGyyvZXd5Oh/3d3nokzIjoMB7lnNye2Jkd5
ZRTINoVSFPjBv00AXogrP9bVGEx0pJVwBSP2igWClO+ZZp1w0ds8+HmnATsbpTRyRVBBx+Ube1m/
Nqi5H1qClL7raGHH5h5iFGo5Q+7Ki6Y/rk+2AFFNlPB8QMhcIfKtBFqC/mcXJaXJoiF8j1OeSKhC
pr60Kq1P2R5Km2/GWwa9tt8mEIxMgf01vckPuhOrz8K2egi+avunRkzPlfToAL+3smgZHM03auPu
t8u/Rw2joHV/sma+wcdLudaC9jkilbLxpzbi+LvFt5fJi2BPC8m4yMwdoh57UMe07ueGpcdRN277
k13ZKfmAT9qaKHAuP5fTwpp8Eq3ltGd2MKOl/wG/FtSFcPvOF/dK3OF8VXOQgqQgJGa7SGYXAdMP
oqY8tD1yizaYgnaK4cfAJQZfJgIaQQnGbPVaMatvm+0H6PgQmwRCNoK0qtaCIK/OZcYVzqIO3ZRY
Y/NVznP49KP2qbYyrru5wSh0lEeiJ5lnCM8CPvY81DWzzVAyBPMfiznB7GgEJ2FtVxS08wWtQwXI
k4ZwK0iZyWmsVAia8KCRvsa/6EIv5MqBXLejChNQDQZZhoWsOhU+KfSZeY3N4C5pWXdLr3biAzuk
SH2otn9ed6QwktqU1VQcco0yFSCBUIQIhjAYr2SlraRTldo0rgV3/OfuQZ+MALawMmURkbW06CX1
r+XOFnRZLX2js0TPXj3JgrBTFip81DOgVwvyybjr1tgtaGaYnyTTGggOmI7vRdkON4K2ZMNOypWd
iGNU6t5Yw2/7bfH7fIfI6jrrjqdmkCmOWVyg+YwOcyoNJGG4+vaPDNJnZNnSb7Iqnjmkcetohjkh
bNzoauFYng4jmHFEyKVuVcd9EqVIpAOiB50f1xBrfJHDbZH4lp2dc/+gMYmaCT+Oh6qNdrRWe2+8
mJfLFCWwCtoxxZDq7euDi7z8TLGzUZJl15k0kJn8A4hHCpmN1zyE5QrnxP1LPcGDIPZ4rDEPN0wQ
kohqc+HkssBS0f8t22T8Bjj7yBcFxxJr8CA176lDCgKSdP7RZOBHVRr4NxvB52Yjcm/TYJf4ftLT
2ISVZf0mTNTnxMfiRsu3rB6kDo5M4+6DKxA8Rr/6R1Ax8RTtmipqqNfvgn5FxcacRzX8d3Qw+BRX
g1DyXzfSuyMUtu4v+HTrUjWwIHygo1bEqDApwiMS8LMHqorxMO+ag330dHbZTqEtAXEn6lz7VOpH
TAMZX/xZMMP3IJpBTF1v2t3lmx10FVj7d4Fa4GdM5MgVhCgVLEY4+CI/l0ykuOkJl5E4ADsC/Emy
pXIgRCZ+Szsn6JscQvX2NYMq3tfjkY04cMxZhqaiHpSOMXDeGKbLNGHtBDdWmXluuAVf8XyduZ9b
I+QNA8wmlHNExqJGObW/lo582W2N8zslG6C5OS5t5pCSZFm9AUofjQIi/gjhJb9AWxZAxrMzL/as
Hy2WMf2WefDERF0uVL+I9FbtZuD7/2gLVrY9i49OlsylXu2rAMQ/N4uB/ZxL3zYQlCf4CcVbhUUI
/qXBoG8Z8Ejl+txQ8m2OJlhEjn0iklZTYRtuE/L1YEe7x9PlIKmZ/bPjimCEZUGPqsHdZy6qeN2R
4s98unewf2f1x5fwri4UhK6L26iOd6Caulek6ldd/OKpk1dPhcA8v779qo5aqoMR7nSnL26pqhUA
DL3NqkWPBWvkSI+3BSJ0kZkCWfxdRisZUCuPqwxFtWd3/ijnZziLt9LYV6d0Q0yuBKeJjp/Bfs/b
HVqUgroljlT25M8xeLFHS1p7EcJwU/5PgWbq2ozaPVKasDWJPVEElz5b+myGZnCp3KPvBkARh13f
H8SMPkJ2Uea/B3nqaeof7E7Zh05TKvotSVL0VVnU0DdJ61JME7Rvna3p3ekHRXCvOmZNLWVYHa0I
VyWKNzwVcPbLGp+nriTouTGaE+rgWQ0YeWSo+cs1lc/RPujDnB4vB7jEJ88pYMK8TyJC83trrSpr
4Wm9FtqW86y8X2oDjMpC0o23VTHNpP/40ri/9HrulfzIymjKdLNKi/KcLL/HKEil3DwchTEqASw/
nhyfR0CIJFkpgupX3ExGED/CmLRzApwnHozrBB81qxKiD9Q5uT+6yd+2KfZBCiT82s0Q9xvbdgU+
cgtnOi9Haxo/GsTfQiDWIn84qlhHiI0epClPLNedih+szYotbJRB3063/Oxuh82smDB1iTTD/bMz
b0Ed/eSuNy9H9eAb+JI6obGb3j1o/sYd463DWqwRSuKwoCv+8jPVJOS2QP4cAc61Ne9KidtT1MvL
Ym5lsCuf2qkyE8ytGzBku+0hORiiKirE/l0NmlKQgv3pDBn4CykvAoeS0FFoP/3wVY6uwSlh0zog
H710GpeccMDIgdJeS1yAlo4fwWGPlaOUQoQGRuqoZfIN7YjDV6pNzFnDXbQoZIbSoMokP/NDhAv9
pJGmgEsTSWmsU/GuHOppyy28xDk268k00gdB49cG+sxa9JVOgaoTOuHo2+k1eP5bQjkqX+bcwJ4x
mt4BZ+5+zQP2XkS5HwBD0o5bO05hk/S9OqmIX0ss7p9sLXORLhtNQEDzYoBxyzV0JFuoNBg6B2Bn
yCZacdlih/PYhmMh9VwIPPGEDbVgY5cBYigX//FiuxbTsWBfcJXdacU/QnzO9tszf5d+28VvFU6y
QGpYPZkMauBzed0bCdrqQ/ECFcpOf2WP96pi+UBVQTE/S7qIKZsW4Md6t8kczM9cQlPQn6LiKs0k
Dlny75gUUqizYby9pqsY/6BhrgaiT1gYAYYZto8puj08ytV+OLCtXCx4zuKQZN+1rvVCE8xXNXnI
y1Ci5sRBwVGxpaRJXp3ZDZUcrL/IYb7+e2stbVzwAr/gvyt6mOv/llfRsOyFmN2qOzHPYc5FFZsp
EhTDcPh1p+UUYiQc2Qi5bklwbANFDORCTd7jT7aoWtzAAlVkOUNw4xGiaUVNuOyY7DDiuyEBz30A
7h56tizJCW/ZVWIhmgKLacIKf7o9aSF+u0eMeKIWdJ/uJBKkrslVA/cwc3MVr3fSI24Dwi+RuxYI
38pYoMoeRRsfBY0zoqrMjm+XhMbXXjZdyp630K2NpWJ20efAyxbnLb1Xuao6iPOfOzjR9FncLutD
EC5aRHJFfLs704q3hVhbn/N10xnZrVkhBs5KsHDOEt7jpuvh7UGj+Mv6AbiWe88Ydog1dZCNsjio
UY3opt38zEfBS5KaoTQeBW9uOILKiVZ9kQEIfTjVKHHaNK7ntiBlAzqbIzJ5p+nBFvb331w/ZhLj
IMFEE6vatsWJwj7OqRMX6mirbVCl2FTfUOTCPTxeQ+xf+6iUhqhbPnEcLdaDYWgezzSQO8KyhgE8
5S+aNg2zJSZ38g6qCuJqAEgffIr6EyGX0mm2dc3SlIURIxWezIeQBAv8PbCfWlno8rm6p0rGvnxn
lhytbjkSwD1HBktNm/7oOLzzDxAo5tQ0vP8P9tbYzcmB5LCWBoDYJoybNdSou6I2bGai0YlabSvS
tElWltJIx1/SBaEMqG+VI4kpg+BfEEUGocWhHSgGRhUl4bIkPKFWJqUWbhxLTGb89/re6xyzEq/S
6RmRZtkvAsWNsPZSd9CfA4u1OCvvXhxM0RQBOMP7lRlad1eGuBiIvyWszUMc5ZnIvK3sQv6RZAvR
K9NJQNkHOEGTuvQGbmu9A6O1No6OIV5EY0F55ljyL2FV8QHaE2dE/c1a+7TT5eswuGYc/0r40uNt
ZBlDqkZ+O7lVUxmnC6W/cm9ZYCScSuZVNstHBC0QHCQZjVU/M6uu4T7WS5ZrTkx+OOfXpWfpwt2s
2/6cXZFaEs5+kXKSOYxX5eAviNMJbegBh46DpFc5du3y7tZzsbMFXRkx0jVBlX8OI+p2IxZrzByo
RTZxobSLSPmMDV/Yp/qpLmf7bdumT9AAmaJr6BRFtJBnYf3kb1Avm/XMHFTOxjGBbgGI4eZtQFP0
09vVg8Rp5ooHjKuEJ7/zyPVowQXzcWcCwt5hlR1cSFtgpkVhnym9LpegpFQfwKScQGwVt0vB0yi2
nzBHEyIkzeoP4VlUNkGvLHSM44JRW0PdBN/Zm2kRYCN5U8JsbfeEeOjvJH1O/2DDuNCRTtza6CyI
uwEPmtBnli/qIHIdv8dRId8H5Hi9qE5vukALgFHNAP+w2AZjm8b7XeBewTYsMLKw3Xrmgp/INDlH
46nRFJwAEoUwRmHWv73RTSu9ly3y8EVoXhJyEiooxfuotuTHVdmyuZkmeJgpoQJnoh5hYq6YiJll
CyQ2uDLcon4ETr33Oyt4Lw2dkts2pwfT+I/LVNa/EHZE4RyZy+Vpdx89bxULAP8kxbhzqwoJfK4D
VHEVweFMHFErGgVDE4J+CMGbS/dRuAtGNtuzff+cOQPK+Bl8T5ZNtBBjC9vE7K8qs/4FvWMo5JfU
37xqGZZ1sHfSBbBEVlH4HOOlEvAheeGCtuhoyCJVk7iTQj/FxKWLXFvmq3nJPOf8taXRzeoMjevd
KB3pyzFBMCmmktlvX0jWyvO0EjyODE1ptrfg1cB1OBvj8Qut6aJ5pg6M0E536cIVgjNHvZHokb8H
ALgM3o1Mxoqia7uPkJ3KCfcjL1HbfW1DmYYuTC4RHODRGGvus1APoLnxTrhwxLDNGBfSt3oU6TIG
QSKcG5r9r7iAwSBwUgePgWaPdl1vDASjnjs0wYMPCa3nMZoTuTeIVrTSlDTCvfzkqhtplLwN+GSN
C6fvNV0Y+nHPVqW6gg4ztrwj6LJv1WeuNXuwmp8k1vmpO/ua6aawyire2kdD1tCX1JlAo6RjvXjY
viJXYA+bIyi0lpZUwgWjx7GGrDVRC8bFOfulXs+Z7cwn8uRoSPFDYkFclyViBXKONWGl5LCY9MWw
X47+uEYYRh0YmcBKqAKbSxNGp3b9pjtiKN8I1eD2JOqrwK/6A63jrHhzF9KtU1ZMIRc29mx7D5tZ
8vX758nPLnv9ZSa+UFdnIO9+BTkVvab2znymQ5Kykv2Zzs56DuGDab/jHXzawnXod63DuDmPBVzg
PTx6rWsuiF1C+XZUBq/wdH7AXz8IWSnP9RgqiNn26l2HJ+J+wLM708DQU4cPXhp0CCfaLnL2QfCN
cLzuw+PdSocjVb7jAe+BHJHfqTB0lCf0sP0yp8WzWx4tVCiNRL8/emT4Gn6CLKr3pz384UZdnSJu
gItTYZiH3t6+YPw5usyODyO4Ap8ZVgYuSLkPpchwwJ7J0m1Dbh5GPMNl8flSkP33QAoZKD2FlN4z
62AWLzjU5ni1rJTuQxIbwjdfjV1aaFMAhAkeYUNYv8E+VIuKB8Zq35p4Irpx0IrayX/g0AsUWN35
V7YIbHv8SMpdpl+vK8Nz8EGhip5MkPrDAG4LBX0Xsygq57JB8gWRMlcnWD8gCh6ar3rEYqXOr9nb
aoDg24TFt55hK80YJtLOij4jqrdrUi+0uAMELVk4ehCdi9mzcv7Ek+SLANVdYIu7Nxs7+Wd7p5yz
tttWnkS0xsAWwEZYq2qwSm8ezCA3cuLNCSbC0rAMGrFGm0VbRkWRP38aH5dSsqAgm8YauI4xXohG
Wi7Zfm7ZDiVzp+Tp5A/gwNnFUhgbCBGzTBegPmP0VM69rCh8H8oDPkR1nrgoQ9b8N/fHgD70AVe8
nNNMGUquDj3YPTJodNK22u/jY00cKckLlplAI+LUZ4eG9BWfP67UudChVOkiYa3RqOTiMAEaQBhb
T+Nbfq2wGnLalwmZ5X73nXPbhA9j9vCyJTyOYULV1evFj66/FHD/QUSt6nz4PQYZ8Za69YbXzzht
DkIBltLkgLnQ6DKXcLcXASM/JzLJ6rln1cWrPaH+AyquShhCHTa+tsWJSFO/G8kD7f3mGuFmP7Nv
dfZnW2/ZZOB/SmwRyDa9JRGQSbPA4tEROmD5B2oJ0DDFhyfsBVWz/uDJgKlYGDE5r58vkIO8SLwi
5CXUk7y92ctGRdm+8no5m+YoBI9yADHe7oaauqbCTSZtzC4vMn7X7ENwtSHlW2hi2myFQ0UOoBlm
FU50pUraRY+PQpk63W1YvbKbSPFWLuLKl6yTzC4AVPutUvHbB933V7F6MuzF2aQP9fUbdrU08tBd
VGpigyzoRLyVZJUvzkyi+I+kliYwbdx+1lonx7L04dS1w0xwpEkm7vdTrN7pnZsMmE0D7rZSYw+X
7XSFJt2hZ+6j1YznX1ci5+WrG7EmuksC+9bPW8lkLozxg9FUyU4PXy83Pcq4kHr9bFdd8WUQJ+gf
LZSc8vpLJ4R/6ypKUEj1cDIxWBKOb2i4K6FAhWb/Vya+jaTA9wWo8RgZM1mCaAYLSvB13XVnK1xo
a5/ih9C8LNk2DgZkD+SquPuRzGJR2uxuSA4ACI01MU+I5CatTU+Z3zbE7U/Ea1rYedTXJMVTxgyV
4TcNsBSwqbhk+s3fytswzexL5VlA7gT+tkVE329cJWlU6t9eX6WhU7UyhXLc8i3QLrp0h+D+kuZJ
hR5tIVZrtWs0MtyEPLiPnxUZq5bR2optF/0JRAkvpqSDd42kqsKwekEPqkDpDuUDX7e0smwjwGul
4uDZ+jcYG2+RSTOpSl+WLrlw7s3NtnqyWuojsIbP9bPgYXbfYLtqJUKIbzmcB4+I0fU9kmRvdY2I
+zTEalwlk/rKH+HnakSYbPic/5H9MUDJozw/21OrCPA2CwZxy5dAbOR4tW6VYu0EwCCJwlPO0yap
HgrG93uyliTMpaoea5XfmlCdqHDrd/BxaKghzbEUMLu5cBpwa8dgMDUfV909G5X23OHFUlU2TBfZ
h2d9e5+2FLxlEPmYaYnW6bhFG8Ty7IH3pGXASeWkB7ai+y91JpRakR+O8cckoBCViN8P3eBNLViO
9lrQ+PfXq5v2mI4YSkYEEU+hTFr9p6+aZ/XK12VuOL2sAEFD8DMbHU/Gf4Y78SHrEcVPPVjmEqK9
3JZwGgVoVQiFZ/dU47i4dCmgdNZZ52LJShGwp/z4BDHMEqKRz3Xr7Eif7Ig3kAPspNLLd0eA88h5
5sBw6zMXRd2tAIZx7t/sKeIpdup+lxWfe7nMf0d8NjqVSRuT7/xUExj3DMJYaYybYSDHy7+ARIbY
MHPyxOMfJU+c1VrShR8sbvr/K0oYy/CyboVnT5AuVCbmDr8gOYyTWxvpZMEXw6triesyF/7ZdG8B
Vj0b0UbiYN5F4LubqAu9shFFpYglewh+e3Fv+bUJi1v5XuINMWlCNkdQ4DiVUS/kbdnIn3Kens4e
4CtAr90Yp8zTUdYIAZDvm9I8DTw2Afh8ao3SXo0vf3jBD/Nh7U8iL0TDVZDvH1Ul1s8vGxuZ6EY2
3QmAA+zRSawVtBYEcI2FJCjp75hh0I7PqnZYvQXGhXQEtZGVpbrKDl/ukoSn6YeGCtD6o7FwheVd
67JsqxkK7OAfWW21i2fsGQGgCxh0gfmmz08rXcOL1FuDbdJfzGg7HOsEzF6MoKu1ahUTt3roxxCI
65CXMTvh0cXdmpP0B0SWKKtQE0R8YHlYu6DFseaOvjO1jvWuuqjw+hfDfxFYddMZxci+WBz7RocY
xO9CgtRB38CQ7iS6OkNuat+T3pJoWv8J3DmIgsUcfsqqEJu98aLI4SJflLYsb7zbVYAJMaD7ta/W
Ax2feHX394kWOJfeGmHTXNSZDcU82SrS2lhs5gl+HEjuOPXMqYsnDZA/VMK4sO1OXZYDa35+T3kx
oXukCI9TC+u0AXBUxoSERGxpiIPgmwiGw2wCv71yuL8+tghVr08X5G/XokPLlHkuzPPWM57gCJMW
z7Nok/aiOzxsGTYdyrRb+oY7Qt/PmtXFkKvw+EIV/L/THXVVuJY7EZsbYiZ+Npq6KWsabJCAtmBx
25PTM6pXmIJyFPCjaLTqnRz1zfvg2viP8R/Fsag/6RBRpdt/IM5tb+4Yp6sxyg3zUfmC/Nsz2Idg
9FkIulnQD4+fsvfx8x+yRMG1XGNPdk1WLtjf0B0dXOajOy6sQftLGKtaawU+Ww4+0JH/x9y/wikB
5XR7yNr7aqiObNabLWni46ewe8fTbAaSp4hubCZG3zW8AptQAtzrfK2h7/iK4e+GgYw3lHnFb0Iu
FXxo7wdwjf/J5CfhqCJFFFl0aKxZdzWER0LG3LpCHfJBk0WCTRrkDcoF/wAVX91WSCyzGIVdlUXH
37gj2boEIsiJbkcGUDdDelNbsV0Y8tAs1ji8z/Soze4/W3HpNk+FtuyPDb7XcBCgJ1JAYr7QYwNB
aXJeSouGiz+4uuJ3eed7ClHrSPCEgtqXoNg9wEaFjxpRQdJ/F84NPBz1aLXcI6kZqm4yYE/OQ6O2
uhWtX2K2oy8/sTHMbSRveVfWP3Rk/6aie/JK1fKNWfq0/MhgEcnEjh1IPfHAJPrOp1ys9PbawE1T
NRWqdFwdU8mZB9RneTqPaiaReWDjcrzjRvZl0o4JzCgoTWdRmeaJMztLpdmORq4E0ng5E+Hcqz8E
K7Ow+L+8E+uD+/qFA4YEuSsu2Js7tAPla5VMk8+0cd/JyaupqarEHyn5nh/xypPCP4UfXEwl63sk
VUX7zFfvnnRZgTOgzgDJKcwigoU0xLYv4NbeDNhkNySMptjPLvjLHywFDQkk/tvZRX4j9alQ/BAV
Z3WHpKiPYj2cSMQC54DoghwplsC1lGKTzAcn5lhRB8D0XJOUVUActAJFSSY6SLoJZRMmSJgIKIon
BOy82usJiZNb+ntl0vTLkUyoBtiMfJ7gkSQmcznpYzSloMlplJECfFX61qiAfMjGXhR8U0XOM2Q4
5wy/ZrDY9e9g8Cd1SAstiaiPld7YHOh2JMRx5jCaqWrcep0OrzUSlhfbemI+3/7iY9ckvtQuUTAw
8aRhf9zXF40RFykuvuXW7fyZt0BYJ+99WkI0akJyf7qLTJmp3vsGXqzUs1ZsdIQTGcL7EeivwqJK
PuGrjDvbUPcwVgYX23UnNM4lkNak97yxeGl23MqvBQ4BqDVSbhK72zHa/MOo5IJRs5FRJYt3nwWA
9uMFePAdH5N6TbbM0GQiVBmKsHKaPxNKyhIdtP9dNUUNDGHEwcoqCMOMlbRIEtRNFxPqW0tXeMAC
knVBh4UTx2/BaXU2z7maljfwJZ4wY/1MhKpqt2dXU8Z1cUgcPYBgM4SZdCTEIAlj7sBLrtycxCiU
6XzremF1lMSzaZhtX3qg4E6EWRzeLsnLikE+3nhCjXYjWo1NYjkwsNn5jUJMJOLrg5CbD4+0IMKK
YdiSLj+NSbR9Ow65bp15awjBKFBbd9MaM0yA4JldqgexMNqJ/pStS0hYr6FIuTgOEcgZIs6bmr/N
MdRxsa5gKmmBxUht7Wk5C/OXlwgAGYR33FhxiPuw/pKp6sVXckFwP787r17F6gtuLlpkNoGqiVTJ
XgOJJRQyu8c2fNiU78ij+yeoeqyXQ/x44IzEUEB3Cdy3+b4PrCDOzlzxl+O26/qfJWI4lGDIxvbZ
fbMPToudpI8tQYlIYYJvQW9ddKtnL2aHc/YIMMrH1gFTWWqpZ5STWyX9W5fJ6/3CCXxllujRT7wb
Me5wO44VDAXMVtFfYWakx3d8RyfnXxL6nRTnVq5WGTPEBWTZbq1BbvLhQ5AFdeFTMnscMrEmndLn
o8vxEqUFeKpv1jsfwyTxEIq4eN6KbymeESzOVpLOop1cCiO+ppWMlQgQ0vA3bD1P5uuGp6pZOfGi
bx+J0M7TCfpumDBnSXutk0TjiHDla/2101+CCx9/FT5stiU29v2UnB+1ZKNpoEh5hDDdVO3nyRAX
nMOzrBYLV5j+v0z6PD4roRStmj/6KnZd4NDaqiH52odxOEr9OWnnKXnTeUutb55LQuYAb3uBUwvK
OPUPf+TkrCe9sIMXEYcCdY+HdGsWHhCXXSlsCqqY75502K+AacC+2ky4UQ8N3KINnBK6K/wFhH9S
vqT+fIysqAim+b0iVFS3FYByi4EAZliew04qL/Yy7Z8e4EKPS+FUNB70+xdXDhfkGZNHoroQvrn3
uOR92MbHVSCgeav5MVoHM0nEBZuoiGH9uaaq+lpPG8qff9Ps4MRtNSZs4+7wfxENqwS970MxMkA5
uBeDY0aYGAUXeuyYwgIW3HpU53HR+crpfZ6GNHQi2Z35fXhUJkM8TUA2Yq4EarBNFpFtHoyGhUeB
m0uHEWHKmlHKb7hWNMg8e+KQlKq/zMwo64c6ykk2tX+oJWHfzsHHCR0o9jLYVaWTvyBtTo0qxGFS
CW0EjUm/SjPhFdSQE9zth3QtvwqgYX9Pb8ZHZ2MJqlSW3p1+2Ku7bE8e9C2DO9h86p+c7S6adfaC
nbIcHMnwEOJdvdW7MU8c1E2j0ee7xHXwET1hsljPNVZcdG+VTkuohZjLsBXeMD3xZWM1nglMXaBL
lXszyBGFqYEy2x6Q7+mlwHE+yu3aetarB2/QB0VDZz1yx+4NxMjj/V0lNtEBhfNnuFCs3x8CmUPS
g98oseGiNesyEpxF2MI1Xo2UgC4roeJmlWpcgzIQvGg+ZCYj2AWJEuDNhRLLUulZh6S4w0CELQB/
lGIXTaT0wIF7lzMODAbSkZhu2sGVDYSB91D+S5M0N7SzSdR7KWitUZz+Clg8TCSf9L4qDMsHu+Ri
QBAoSeGowZ5bEzvGW+ubmEryk+k6IuIi2c8Fto2Ecmm2fzfYxs3jS0R41VQF6ej5OleDgjf9FV0P
lJkETAihWV6V0z0rXSoZeb6uzAmhBB5+iIboJ64XsgEKy0dJuM9xGq+u7aEl4k9TRYaz1j5S/ZhO
Mjxp72UoiKMPk43a6Oa3G9eao04mfuXDydC110CNF6pGCuDy99nUF4LwL2QSBLydnXqdAhUJFSXD
yQXx9XM0tHnd3fJb4W/WWfQwxjF6WZ5xDJeRadMwl3XLADc6ac6GR7ekMbS2HsaPZYoJ35F1RFSU
EVFx2XRWxG6h2iDZ35eZGQktqNBzy8CbYhSADrURN+eqM2q7uy+2U0OLhwiqQIA0g18R6lWi6j1U
2WhhqzKd9mI1HBL3rMddbD7HxJEN6YIbiNqgvCZy626oXDgSTCNl7S0/kE3NZk/VRbJUJJu0S4TT
r9HO3MIZnkjtH652Yr7gQN82Jm8M/QcVqTIjm/MAyNRjV92Lb/GJ28BJpGxInbBNk3ZfTsRpzeYC
AeuaTSTCqOcV8v/k194T86wwM5dzsCpBVhr6WLl1KTPkQhLwD2rAL6chxVp5gVfV4FIghT/+9ciE
ayPnNcZLT800AdCBe7qJu0JNnKHg7sb38wJxoGBICWMpUvWzhMLCStk2M188bqhSD91GAjrhSK9v
mzmgqTDrwggs71OorJPtn2gCTESiHvpiXRWY+vuGSMDftRh2UrXAs81nk5CydR69s6HjNZHOm6PK
FRJEvKSDJcaHa4WvKC9pUENzu9OXKNcy+PB3BAseMYI43XUZMejd3ER+evJBCYqBIYeFHkTmNVW3
vdF71abieUWk7Vk4i0w9L/f9uWjg956qRnQyH8FV8mwJtL2LmN2lkkffSvO05rL1NfAQUFheq8fc
amNU6mY8Nd6JvitkCOykBJ/G+3ijLga76/V0w3qC8Dj7fFBbLz+ZoXHUyQI6xuZZrH4OfvgDaRsl
ijvC1ZMG1+ajuYSCXcnxAVjdQ5sXpyR6NOgEdIo1BLSy1EQcWQBmDdKW+9LD41iUvZzr+q/0FMt9
2gBXTifG24hh8aI/L1IrnlPoLoKuCNmuQ3z+uEpGmI7W7eChxO6LwuBzLCUZqkJKBsI6XDHkwdAq
A/Btte9zkXiop9eR2oRi8G9vMba3Cuv/FHW75PPNX3Oj8wb1b/kFJhqoUbOI4KkhhvdNW2E8LWWX
NuhfRVyBJt8kyYXuOh1/Jc0Vm1Ny6OTeU3giacTDxBpeuQszOTG8r+xsEvcrQsy6+zK1yVSV9r9T
kkW3MsFSBoV+TuyBZ/vbyn5QETn0GQfZpgV+lJI5kwXqIoozYDWvrt6fB+tVAS21Dwf6VoDOD06O
iRcaUWFusvWXahmSWNp83eDcBo1vt0/AoxbXMpanjSULIHUTUUvCIkqFYFD2cQkzHI6WGvznVQQg
GFdDQW8hyzJNE24Epy0gW3W6QkFyrngge5KdV55XsCclBLdQ2hUXNnBUuOJT/rDYEwU8eu6Pp/gy
LyIJIZ72HdehRdXIWyLkExsHO2D5zuLpbkqUijVCTZ0uD/CgTLvGAUuob+0oVKRWHUnB8t/J5xQ4
yDEO2ffJYouFwvKMYNpUqRUj6nuDWLnJj9rxYeyx9siUZxlq5u63x6ZLw4H+DJiiie0RVB/icINV
dpTQe3E/fqHUVJpF/+jqwhYBUjQCVBElzznB+iTRKnivyEzRJkmMFE7PLTcIaPUT0ujI47Aj6KiY
RmI3BweS3I6rOUfmQqPzQWSUByzVJjsTErHA1L8HETRGicLry0jnesajv/VTCYyZ/z62wkFPYluO
3BpVyPs8CA6DL97fboXsplFnvs37yfMSOZbDJ17iJuqHUjQivYK/IU7T/kAtttY6qV3fr8et010w
9ANJLsIIc2vIKQA6yUU5fJxw59CDd6lGvDTRAwgLaQwWJ8sL7X/+NoQuBRyZrMUviXxgr0hASKp2
slFGZeUUZh4qngzRUwZ+vDEVjI2wkmhUlUomAJ1lnq2CHK1Apa/2Y7jbUZdL4kGOhmtvZnT7cVRt
w02oJdznDCByZAa11I7+6y/yP29sTghdGJKY8ApTOkw4xqruEMQU8K8wAbi++Z4iZ8KEjTmBeczP
S50Iwjf1t8MIsdkZr5Qg+jPnSO8/87g0rcIx1mr0SHUBOptb5IdItYPlbncLdUvRI31Su7iAuJER
Q338+YfTheZL5F7zwfrXPHcJwVTFnwayvEEoRzWDbZYF/jLTigcTV5zmlp3HiRKAPSeh/vT5gQoJ
gBss6Lvy24Lm32eAjUntLW2Jvf1V+47QWy3oC/dt/H2DuBrVPt2Y3u4a7GdVdcjH5Fw9i+a4dFsu
nztFAdnt0J4n88lU1X8wwf7Y8jLOWtGjHry6xokZtkNn72CU2CJDAwr4O4FajSBXlwIwO7Wm+en/
FP+80lYTsFskPmNCmhj/clbHSbzQhWEItJqEt53NBKxDfiURpJpb/GfCXTJZbmcHH9SsDCoU6b7Y
4STNXta5bxgO1/QsLaZ+cuyG+UbMMwgkn3odaFyhp9Of5aKKsMVA7qiayKPDeZV57M7I2db8WW6O
6CKSNa9oYp5/kRwRyqQu5HDJLHTzdCnmf9D1nPVtMJvRbYeVoz2A11k7PBSe3OyxsYoebD6NbZeb
PeriUhqqxRK0Wyy/PzzRUjsk06JTCTFX22eDaX/QU/Zr4mAIfOrqBawOFoMmHJLuEpagcHGGHQRD
meyKsBj2KIGIriZ4ZzU8zHgPFw1M7AIGlYPsB7wlXKpQOa1v9GWXh2Oz9fCEspz1ufMahu033pSQ
Se5eT0HO1fo//a+fkjBgr05CFMkEBi7L7Feb3ERQqGiWEPnkVWH0hRK8aryaPY0ElytXVAT3SYmB
KFePAfdkH2WWiA5s2PrNu2lMSS2R3UCO5h5yRsjdORTFCz6NWVoYyemXTJl64XHzCFNA98zJzWjM
RbY3OX9fSB/zWSkEHv6GtkZZDnwB5cMmj38vvzNxWDSTWzybvj/DSUoVE/pGOHMA9kZ6iYubZ11i
dJ3oOAB4619A6Ykbt2x6nNYUWiTyHrjU9/tE4rjIviKdtFBM9DnIE2dJpohf8Ae0Om2OciPbMMhH
/BtP7JbPoiiz+shddIJ9OCFzWYvZEKQX/HdqrYFvSiyYRlO8lVy+NgAspbfAggOBA8pa4VOjY5sj
m4PWtOtWqtqOJtT+N/iJxy2AaMBD7E7KY7aXBbxgbPonh1kUs+4HAbDSAsUTOQS6MtTTuiTR7U6f
m8OFxq+oarxSBzgPlYL/cOqwJu5qIdyS5LfIgpbRhw89N4t8vAtQmqDkitl/mNnqUMyoT8gPczaG
RbgE1Cb+t2PTh+E1iN4Q8+4/iFMqL5qvm3j7TCkZMVH//g8MkIq7933SUa5yb6oXDO5GVkJgPJoJ
zLOxPH1Ed6UyzABf31j7tMC9Z+tXH28XRNZnW27USd/mdITLAxeIY+tKmWXaY9ET2tc/2IHBl8Y0
QiKl4ASYro+Lk4cn2UJPEF04JwLcL6Xjmn7A+bIUZZPV/3NDUbLfShxmJ5r7+y/t2sfJiSL09laC
3K+YzJ9dibJhZEAtyd970AkcNRsULWxwSc1S51CNIeV7TUblwsI9WJTqdUoqfcTIlmvNvQWy2gVi
hFSoPpbxJyQ70+LiBY/C8wdzNAVr9ssP75rCIba5zn4LpFxziDBm7m5fLw2i6/93Y2nM2BM3Vfyl
k3PYAcu1gxqpZDptwMuU0aOy3MKC538QGZobM30EtFFF9uuCFX6cxcinkjEtS97EoflYBpUtR5Ww
DqDH9nvekB9KReY7mZAwZ3qCTTtBYcjAJeCVIbR83geIgMID+Kwypo8s5ILeXv/Gz59pHljcF9me
fSbhPUAeRxyGQNt96vR9lwcDx166/ccDZGlq58VhoDz8Er5MxO+06TL2HgF02dIjwjM9Ch9H+nPC
K19HStNUAtCb1G8FoMj/f9lD0Tnfb3H5W9/X7+JhvUd0fNVOR9qrpMcylDXWGqXjJN64TBM58srJ
qxkuGUAbyACM8h0yDZK1TjDIQPaGDPkGTOvYeB0SvcP3DctWn0OKJTMDEe+qeXXpfwvnRsWhUdG/
JRW9UhWUxATHH9bZTZty77bM5CkXW0DsyekopNVUp1Gm2OA4e8PbC65AiQqj4zvnnFEP0tKyg/IH
97G9jDoqqtwjMs97OKNBsV56FocYGvJcaYW5ysi1P9ZlsWaLAo7cjJ+/k4rLHNHIXJ4KK5P/oiDA
Z2g+AuraFXRKmQmqC2LjpReFpvbKQs93ZiE5c8sDlJI8rgYJYnRPErRY0Ln2zgKCOF4AVHE7CkeF
UVzjCA4OOknj5ApSO6zzsTRLKTyR3e+HJ6J8mP3EGvUUVcvnqgtucWkdQbDeoT82hdgRFqkfEclB
47Kfd0rqAripAPSBqEDvLjdJBKYh+uobMvas5s88y1mYfKIxlcK1wOyE0frFifhsb37oXevRu2t5
yawU5P9KtenP3yYFQVAkNhjUe9xr8Kcy8ru5mNkkKROItzWOtQMlfQleh/EpisR7XUfJUgmupc8q
DAJTz9cEVObCExiVNt7FwD/jZyCbhf/jKuHzLpblG8aWuCKDr1k8gPoXaVdCPx8juXhA5S9WkOo/
zWnNCv9r15Yn/tQD31Gw26OceUJi7CVMDfwqdNG3DZh6xi1BcKLJpt9qE1nh+L79CDqoIds/rytk
K8EY2EHlFxlkfAWVbXBSu/tPNkU49Lu4ZAz7LyfIkQayPRGSELCgdAkePYPH5wQpGE1Kk0LxOex1
cGtxcqdvu1dK8dc7SPHsX8kW+Fscpv17w9TrpwcWgNvameGNyrs+vz0LG8upt38jMIKDawe27W3A
S+otk1Mkps/La3u9aX9pqEd/xR4uHR9XUmUZQojvM9BG76FvVW+ijePisG8zY9cnWxmddYpU/e4t
+IeD/oG58HaG8LZ4z/CBkOPySWFtiMlXIFpQOWwcNpya3s/MI0biHtvWjvA1blYy+XOUWHkw0F42
pycm4RgcWt5jfAkXGvnVsZ4nFQhA/3eMJBXGIWtxjoe5NBGLHAxYTa4TIJeDPspSBBuxm0Gy3OZU
rBKSYSq3GMjeobRQInvkBX3NvAZcoWRXZKXcIyike9zBonM9EQD9JIKVNXXpsuMcL1JS7ivSHDvp
WxQ5hh/iMpsIluuyNxlVeG3Q3zTyFwSlwOT/MYRhP7ZwIEQ3ehOzVl5pbRMnfV3Z++3/GOFGwDZz
boWU4igM+NHqab7NhVg9N3WU8opmMtwEKHfcYWtIYy5D0sIb2Mihqw0j7uA4eaJlkcSUC4wG79WZ
4wZJ+C4Ry7ILHt5qKUZX1olqyhRI3PLLM/ex4L7YGGviIG5+WeVr4s5GpkkEQDNjfy+fwOC4obSd
KkR8EiPkNpyRfUUYzN+ezWZwjdaq2DwQnP7hYNtILX/ibZ9nJmebX+1rT9VDyasiyHO0/qdrHldF
d8JJk2rntNwFTj99vg70yquebaLgFYETEr3q3O2N8nuFWCliObS9NJHdwyLv3zLphZnwUzgTzeYj
KQ0gG91oRn52Zta3/4rVEiX374WvfsHcTNpH1pFOZdesLoloQsM+ULXsr11cG3j9jCmIq4SegElD
IFG+ePAyJ3BIMnAQ7LjBDYTDujy0rKOoJuNslXp2QeKJcDVHHGGc0ZnspRkQtOjy/aDZAUjz6NUV
6NfL84AinPLlZaH225uFhXy7yWjuSYpsz+tmqQF1ee4hMYtysb4TFn23/KAWluO5Z1FQf4Fk3TrE
F2NzOhBAPD4banlNqmFtqQfNeInql6muEWHNcAruGnoeF8eFV8i1RyatSf9TeoW4fTDU41+b/0m6
ELFuRSJYTHsL2FxJx1EvsZb1YP0agKQiTgaBwpa/d8ABerf0Hz3ojGdUaJBkm8hzo+V5I5Dp+IRL
9oel2nz4lQWp8qtdBOzyQ4eDagFiVu06GPFvy/N8i7S9oBDhc3KP8Uk3ZSIuClr7WvZXMRLXniOQ
H1GDmq1AKIhnJpOioIhdVhX3XniqAqDl7zs7Sn50Fak6pyYu/LuVgW579CSnuI63b/zQhASR2xFs
pSVL9MyVkHjdhGbSJa74UUz4YKg3t9sNvoXIXY/M35UXMS4ut37v0hOSOPrd76eGHAIbL/e/fL/k
vmEq3YpEk521AD/7YXO09UGuGS78ASK4kTNsgYXOfQ3htxqrlK6O377Js4wvdeiJGo3Am99QW11j
vesL1ufmgAPHvngHMUINKXy3EYgsTjcXzb0I2WbEgoB4bZYZfb6bUXaZi5Z2WJDVhAM1TkHiSTYk
b8vAqUdzKtxAwzIV5usmRZZ7qYwRym3uA2idrTPBpUXuzWyvbCrn1zPP3pZIFayhP2JCav98N8+z
jGdhBIKjiT5gzbx8dA5FHXUjnf+4nBY7pJ/v/kgUW7BFmRD5K/wy7NgRA4kLipSIoZJSr2jzxOo/
sD1g5oyaG1VuuMbkRifC0Q2a/IAmJSv+OMnRxfzs75JZoN7R89fzHf2cDlU7F2HAOiOjvEyuT1Yd
RllUFhQDE9RiVsAUgxl+ZFC0XjZJck6OHns4Ex1xb6gLEln0VOY9blOXPakZ9WQ0aRqnTY3wTJLk
utuOvI7aVNcD19vmUAXlWBk/gDqq3O96UJmHtlJbbcuKR2AQbdSyMJAqUepTC2iOL7G8wyBbm/jA
296plPP6+liPMYdx9VbgLCXZGlb03tJlst6h54hSLTqt1TpiVUVzDWHGsYnM++TQPk8Xw6i7C2KQ
n46XmflW3qi68XKtx1jOBM2zkBFCKfR5IedrfmTG8ishd9LjL+6IvLaVqm8PyOVaT7EX+bdyDFQX
kMuyXc+hiZ3mmEY6YTM4/85Sgqmyc9xF5aKd4+f/g3u0nLyuRjfyLCsnl71qgZMBBAZqWFN79UJ8
GrsEjkoxdvmMHtQXKTZrH1oou2ul4Yiu6a4Gdj3t5UsijCkmfVDR2aSO26/EaCGx4MQqdYN3D1vh
vcjUPy6PPGM3/mG8+cq5/BQBKqnjRk00d78twL3/gF1SkJh/N51E5YNl9/nXd0G2I9WC421KRSd+
4Bm+LgaaFRzCimVZxJfvSafElSWmKZta26MUt9qVxeU1bVqTkQH1PMgY4W8IuxvDJlThEEwqoCt+
+iGkpXWp/2UaoBhUIGXSUEPyFaSuSLJTbXCag4HW6gK29bJ9DrTeQ8wBIzqznD6Y2ZetaQHwx8TX
lmAuRxHTjDUbu1NZvqextpLOTeaCN0ZQcAVmzFaAtBxF9r0n1oJS2Udh8dSajsQLLBOJItzVHGWD
+hVpVDxeHIhnDzEf0L21p8egXeLL65GrzMX9ZCvf0ATtece5IQ55gyajTZr5HtgNVFUrETyIvfJ5
JVr3JUccvNbHaKSbc/uMrOduw74Y2Jad5mF0Ff1OuwAeUXsKeOnsMaejJsUA6OFfCnC+x3AFzhLf
7t88oUpoTlrWr7Py+cXKWNfy6sJdvr1ouln6LA1279pcX83Ss35pZv3Ilual+4XU52+3QZUISqTD
RC7I4BTXQOQP1Sdt/sc4B38x4n2qi97N+bG5Ig9e5ea10G/znd9obKgfjM7clclI30ALMNjcxhgp
5rM4H80lKGLWokqLclgF3b6nqG+tSQ/38Gv0lbD/Ixx2vAnQPZyDgmQlRR2UdPgB/pM41J/YRZP3
wrMfRnu0vbdFcvjZdR7GP5yIDurb3xBhq+LevsZsT7G0AvgqulbRSwm7PWRM15Z9NUOXEgtNPI7o
HW9ZkAPsQkx79COkRpc/W+sd3LTXtghX7hI0kw9C1vGUZ449sAQS+uE6Kef42BUCP7r4lx+Ctz3y
04JRZtezqGlkBWYQkrTlaO68MJ0Wn/7n+Qv6lm689LEMraMNcbraMX0N0T1FQPllmhUnxsJHSDbW
/GUo6ICUKoSOcIvKB7OOs50WIFPT3uW6FbZNh7A2HG1qy5o3YlYLE6NXK7b1a1MNgLTU5SfzLSAd
FWVjhk3DNcWwh57r+m9t+f/zOMFu73/Uw7lX8IGJa5MxFHhbLPNtGs3wAMMPNYCoApXceScP0JQ3
KMggH4rWQq4Rk2U1q7zf6BuDMFdmEBT49JxVvIa3NCYcXz2znKFqYCFGbHxkt71ZEfeCLWPpScqx
ixlQ8UENL3O0/0LoTT0RruDr7tf/wegCfSCsCqp93AacQIz5a2YwZpUhcL/WQd6NFotfwojEa1mq
ON6OGDvGyGqX1YRp44bvjZJ8dtCEcvOFoQB1t8hRIy0EYZicyhfM7/FDgl0eDPJJuqwpGSPIBlbk
p0fTms0l/yWPSTYurWtqze2O7MdTU7eO6cqt/GVW7a09Rq6hVjWdRPzm9+woXoVJB4RhVnCvC8zS
8nHJBUV6Pf0DN+zQW3Haes50ZvKWaYodF4uujX+7gbwVuVkCTgYF6vfZRjA/xDIKkNuzrAw5J1zc
JD6n/Kh1y3yc4q2WuD2Vue62h8WAr7OwnYuf8o1crr0mlUDcEe5E8P96ORKeN9fFaFyZQnosAm7e
rRyK7o6XkcVa97JfBMCNaiT+LMZaLbN1lGJvx70whzPPIABWTfG/rMLI8Va6SPWQYn2AT+sZwRDO
AM19OnWd0qQjWF7ssMoW2OXcKBn4FDH0bqfLBDmGw9Yp7R2ZMbQMSl5rK1uyu+rj+hBunZ0Dvuk9
yVwIkJ1hEfKD1UVy51EV/yDz91UzLJ3D8InDatwfKyO1C7jxOMbdRIFShJjGQutgfl4EcYVjs2em
pKuXoo4bmCeTFeNRqQxYXZQxtXD3NXYyg5ojytmZzm1SSXRxXKFMNGIaVL4Hh0ej7qHK8ZcVJXbu
tnThm/thHbLQIta8W7CI3VBUPEvT4iG/u8AKrDCaunEndllgVxjOSrYvQT3hy5mF3Ya+kxUDlyQW
Jr3/WOxENAix78oDjOV57E8eGgUl/B+xTEIj4ZxJSLbA/MpdpesiRsR5VL44f2xSrcFvJDLLvIhb
1FEo/vz/w5EXnPESPFB1FE4aMfulEgp2nTVYPg6RDWTJi2DvAzFJnvhWFr6iVyjkHFxJk2nN2zTN
+jLmC2SJvth+8c816VazKu1iLHnvo9OW4uDp3XRvGyvF12EYBJr15FMt1xHZz40HI5gBEvDpatPv
7Il0ELJ7QTHRN+gLgLPliyqetxyUugSrxU6rUo4A7wrLgptO/vJRWJqsdZAI20I5VAA6b/RWWDo+
Bdu0BM0NvVjx7wpKNFk6FJYIwD/eVwOCH5icftFzXHLbbmq0wRZvZYydkcDQ0x900hm1RqtdgEnz
I8lV9pD6fyYC1MLv/xHc5eTMGsSyC/n9BI03MSZbq9z3y6EmgAwzOlAaF/dt1VnJm0trsD9Sz5vS
LteSj0xmLHYsNGZ6F1j1gurzANmqSuftCVKQMsB6kKxPSkdbQqQI/rghdJS+I9MSXejdx4+xJ3z6
lnLQeCHvBGV87zCBTdw5vYZWmQlOFa0fui6QVT1JzLpRRIr0bJo5y9LtTQbkHQ3XkoLEhmbMCjBX
2iS4SGUErS7OgrtxRQ+c52E0NbrvLGiz1iSLtNIdyvg8qz/R3YjfYZY1m26Xk+aDVRUEIIx6Irry
F/DrBo2DJf/PVuhO1hTaJycgzkBUxpUYSZIsxqMIgsIWxLq3IsTLkYp7d8NK3xv52K+vdf4nzkVU
wwrP1l4xz5kRf40W9MYXAZK/ay+CAQoskkgrs9sVOy9QlCxMSJeV5tIvI98LslOZFejY9IlqvSjK
PmX2JjrBcAwrGoJ59kcaIh38SRKhziUGbJqOBAtXxS8YYlje8Q3WQze2yuQleJBJ/2KLIsXEllyY
Tb01zjr2HdCyD0onmII/aO+sdx1UNmKhIUU3971rXluvgKoSiJmxCY9+HupjLn5g1cf0l6zHk90X
rlpnU2LwIWHqc+ZEnWvdu1r78MruvHtumdXix2CM1wdP+HBbTmiNXjArYlQtZIAGJNB/su6/hBLb
5n4ylGLOKmcOUbWhgLCI5klVF0A1X5n4bQStZk2jmQvicC9auw4ptdRrjmYpRlOpthxsMpugaoUL
ZxBJGuu8Hf9vY1pnI+w+vamKIf3UyR8LHxgjqSiDIvvsSP43tJfhqxG1TEyjkBwC29MDFan5vTwn
ERFhHwhHO+r62+1moKA07ZDf9ImocmNqLWZGHg+QKZrJXjkIMCUsY75rJH+ecV+pzIOadb3+v0gC
J1WGygvgXHCcgFNpPXm1VUdPA4Ug52gQ6g8khRizxGff7HUcHbXD/U7V2t6Wn6oIBMdA9VbKxXNx
3YhswnsTyo+qt6pCA/AfRYrMIT0Q1K75XuaNmekCJDJzpqGuxSvHmuf28qfgO/mVXsRdIYBbA3lI
v79yF1364SKfIVdeW7uN69Orc+H7msiLS0PJpLlwdhoWCnPTFTtHT1h2O+NARHs+PZst/OqzSjUc
QkmsSkItPzQNVdewrgMLRvViYSis5nm3UDqATHfjB6cH1oWUaB0ja3MVy1qjJ/SMB8XiPyyaJKMN
sEVoXu/xgxjR4/pvkEcITq7qx7xk+4fELFBfDWvSIZucCtSCDQoA+rkBfGeF7Y96hpOqX7Rg3c6z
fsSffigNFGtqyTL52GpDJek5AVzBLfQKSygBwtCkMHnG4sD57toevr7PBAyIW0l8GRF9mO714I9e
9yO67mkQUduQU4E9z6Q2LfKtSd7WgvfI6Bank6fn3lQ5YYuCgfhhK4a+cJfgPsKfniY7DsFhKPT0
fPlO9cGykvf6HMYuFKRtt7YbQqoa1TFxIdFD4ewbJX457JA7UFPC1vrMM6jEfZWV6mm4FjPahzoA
sICHIkr/L0k4hvL2v7dXSkXWbgtb3rdgbXzHc3OVC8Te+fsaDSe5a94LKDlVmWZQDmlb6jDtQk1U
mx/bS/hNQvfeZD2hEUfp4kLWiggyjeSnnY3mApb/JX7PtRMwGp7nFVl5/xcb/zBIrs1DUdPFBpI3
aysjyJ8oPirjmXZ1ozOVTU7ro0YOApqZE2C4iSucbrg+8EdQgwaFBlgufk/SDGKwuj3VVjXfIxxG
GZQKlyLJR67zH3jaMD8U2EbLIKf9WHh27eu6uhOWXUpHp+U+8lO9qglxh7Yftx40I04zKZvpeilL
8aamGMKE+09olU7pfN36eM6K1mBP/mUuzytNDeWpEsaYHEt0BKy6l2ScxgApuxbqzWR4JpIfogTS
0iY/8GDVfdabqAvcghikxt4NuTB2T3EV7o+yTy0NCS6yTD37L0Av8KcEXILD8aLZ4zpaLA2AVExk
rWmiNwTi8cdFuf+ek7t4QTfC4BYeN2mvgkKHA+sUcC7IhNCuHgRQu/aKzzbPmK84+3mzgVcvB93d
JVS9y7X2PC9QyVhaZRhirwpFjPNZmA3Xubs2vdJeLwjkrKTUrk9a59BdmVG/OMxDVTyKLVF6QAK5
rj64pTSVMIhbq6BEQWNCvVQHuNtXMlHgKAHQ2AFQN2QI7CpR0dmmLBkdxx0RgdkAA8n7m652Tsuk
3Z4LkuG10JRA+XwZMyBezV00q9WuIaenYcrBGzWK78ZgYRTe4N+IvCGwDUrO1SMHAVpjDH2r2Wcj
/fASXNPrt5IGRmseCDbacqn8YDtlBjtRCU0vwfBUVuDEKZhjq5tdopWUeE0Sj8gfrxzjHNcbZce0
6dopvVLjMVXteCI/hWTgUxWL6sijzr144WDcsQNHXAI6vakmEhVTNZgbW7oFmZX3pJXhVJPZuYYx
r4/0JBLTUndVoHUOTZ24OAGSHgxmJEFEOVTZ5OeY3sOE1trHIyvuq35Nzff0lpN+H3a9n1exJSTb
TMp/R0iTw6q2SILcVgK3ZXOqzg/tIASWY9ixUVaSZL5gwdZ+p4n5SSwEcenLiS9XTzNbukkoNsKQ
1nqVVP+kWwRxQ0mkdMcK1Bj2s9zdTBV51S+MeMVHdEJm8t+ne280NVYYsfF+HOn/teLQmgAPgWXf
G1PXs/dzq+oFnLZctdOMBIYgP2FOXkIegMQjmAhS7IysdvFVITykJErmf0Wy9fYYsVal42y1Yj+4
YT4EiyDiFBO2yu1ak5D6L3x4oXmEbxWj3VUQjxIYyg3ahRUYJa4uB8CegfCgX6bc+YyrmpEL998M
lFYOQ4QmfThaR3ADvyQflEwpEjXJaQZN8CSzvdBXephqF3RkTS18+eaUy2tmPRd/KrnUA+wcVi6V
yCWCHdLvO7YuYTX0Isp+fevDdQywZYtWHwcRarOTK+fYDhyMbG0ZS+ctdwPqUFcywlSjYD+boJ3/
T0fdcVvFmemdBCewcDoIeUYwcMaHWhHgXQ2AKd8BmwtQlkPqbg8Ui4kYCbpS1o2sZHQFXR7SBRgr
dPYFGKmDbwclV43FCBwvZd++FkOv28blznfzTS+1yOAZedeNJdOuYH3ajHXPaEar6x3GdkR+burn
3co+aBRoTiveZrmlV+1rW413w/BREq11CsDj75rfnXPEz1IjrpWUCmZkN73BatJvMUjyqkLPTpzi
KuY+hOhLp26jKWNocALX6kqpD/x/C6vSVZHHLiWBQ8WrUtW+RjKCGevyDA0e/Qx9hviNCZOs3e86
tQzVEmYcJYtCs3gk56lBnzz0K02TDQ0mICrmD8Z19+Os4Op0HHQu+nwlRvLqokyt35F2QIMbH3uu
G/kFlf75x+bfHqTbqieFpQJaSuPsEKTVmjHU5QiJyZX+nTPVheqWVs4YBCglaBKUdBLzdaDhJ67Y
ybqfuAQTyOEZQe6slByRdRD62Qse6GlmTWfc43DGv4rxBh+GzrPkIRMmllGNeJWsQvCzc+3UHX5I
G0SGC/dtpYahei+RfvNweq+yQcldQkkIvc9sjED5ePkuBebQYT5BAIg6fL7+saAoQH8QtbBhKI6B
jfKoyQPWrDcFpXQGiCj3z+KQ9Wb+gbW3htQuUedhxFOskbtkX+74yoKelV5xXZ9NAV3bX3rO9p18
yOCR+6ACixAkD3hQKRP6kPK9jskFhMapnzRHxhtSoPZPHmRbgoto44bmjhO7WM6dn8uEarxebYHk
aqXRqdkYiUxJzOsMu6Mnd3rYtFmjAv3u4LZLVrni++Du4bnr1WWPHY5CteVJV6Yr0Zsvr0mWGBa8
0DZN63xd2r6XXv66Ti3su0UOHCy7f14eqFX/jYQt3x/wle8jjThxQqjLbUEwap/dtCCKhJj7DvYA
hyqZmFKFhzxP0SCDCjUAHkWomCfh04G3UHsf/L7J91ERqDhxfOOEDqbo/tvSXlAZ38n41nPasrL0
C5iM7Fcz05mcaZQDK/ABFbXcNwLCIo3v7ywxplTqXHy8vAV4BAZ2oLrTZhgI6LecILOaAy7Q2wtp
LfPYW8JIqPL6TBIoXfYHJdiaxvRuz4ThfRA6BYn1TW/aRrWtuzr0HoNbZiVDm3eJXaa4fZjgO7wO
MaA1mCwl0wNup6w5QkyVVPW842Hupz8E/rU/V8aQmTLGWCl8tdkGRwITLz/SuFx+mbonTWyqsleP
tswZJdyK1en+CXteg8xM8mv2s0oJmMJUmNjLf+6e9y4c7GuJBV2NHgLi06edD3+VP7SRS7PIhco1
nbaMXhbD4T0LMAi6NNuK8Ojf+j5jLXFBk4/MZfDmRuZIM9JSnAU21d3dThnOUGY1fisMBplouQY6
yL6Bl3/OjLhqDHFrDNKalBwz3rkG9z0wlQ0VZTe6lmNJdA3/WxCmmbANH9tF4WAbZ22C4T/Zc245
hrYIN+RfjMJUNGXK/SrH7yeXYEfnSJeApYNo40gvLGFbPvg5/xAAcXsk32+FF93U1ORTF9m0pDaP
wowtKUlDIjiUgyY+zQrl18aH2kHqRIhBhQzGbUdmbx3UrUiWTlxBGF6bauF7q1/5NaiPmwgyFcnn
6jSFvJfm09UWb9gKvOCB60ZS85RblFY41yOaeN5M6nnaE2wBD1Tayvn7Kfcj8Clrwod33weRwsDF
ErlQTNHtvhxRdnLUmwLCkpvn/1JT5hpsV5SYRehOq4QP94obLNR8L9F20y9Pl2FW53+Wlwq31oE1
MJ4RxJBOhAt0bG6Mr0ssAMOSCNH8T51n6oDmudUuiAGty3SSjGNtoCly/xJEFvmMMhWljSC0ZDaY
WPdaQUAj6a9pRAW5ygIfUrCBO/+ab6ljM7VlwhOpBxzu0Eb9YX5P/enGMCDJtWYm28LfcN9boR5l
pMPwiO3PKFb+zbbb8IT6M+CwtfgpgFeJogxp6suF7pG2+1qzxgs2WbU2BigeLge4J6UsBRYJwCDJ
rFKOrexzv00buuq7DrUsbuNyJSOJEWxjjeqDpyObbXDKG37YgdHA2gTMQ3wg2D1Uo0TA9lycEYB3
I9xOOMaoZ46yy/s2OAm5/nLtYkrH45Vh4QT/hy7ZO70DxpP83KnnP7WQDaSG7GOupj5Iht24Mtq/
DLGn6aPvr4LWLX1UTzFaJSsHD8+5s5Mt63PTy9I8hQKh4N9Q+FdjewiTzLk/OWzkvm/GGltvfuqq
upL69YtE41P5ob3YyfEk7ey5gez+HFPOr/TfPTDDqHuY/65Tj+3cDzU3Wk2Q5MoFWaeyoJ6JLcf7
+sfgpsYrvW3sq8RQAxTCuoX19iqqiPPS6s0Tlq8NCCEFXMpXsnosOWaFqNpH57brzSgywTSgjbqt
p1FW8MOc9MaqN9+ro3jaUmKBMcB3yvKF2ddVR4mx9ImDvHPjRVplGySGRYiXP8LtXjdpiheAKeAz
l+E2ZvVMr5bEUpFOnBw5zKVRlHJ53IU437b0rMx7J6A0BXyafnjZyZP7KcpxXjH42qxE2byouQej
3EH33fePNbdDAX77l8yYs9zmLtzcvlE5TwbfES3NPpSq7DEEfDmLzYxtr0WYvCD26cxpC5LINCKn
ObARHQyFVRZccMnftwPJ4TmjhziT8xfelt/7iIvanr55m26AHKmSXjkeekpVIZSZ77dE6BBEEgFg
L36eVY+o8GC/1sH0xXT3R37Pn9Pknax8gdlY6Xpi3KqCKRgb59GmzVhp9vTZqv1uH7xz6mptAJ7l
j2Vk+/WnJowVANgxOumsTV9/ThNH+DO4Wso1Lu2zPU0z7d+tgJakzg17j2kyaEF8EPXuBJ7LqIJA
6Xq6CPi5GbR6lr0c/SWhmj1ELme2xHxAFmQypWmby9Nfrbdpjz57Kvdosytt1zBD3R1uPUNoriLk
Q7O11Vvs5gHk1eMUf+jwtMTFJEwnr8yjDo8tKh3i005/HifVP6fXbx6Klk4c82JQv9KFZmG8820v
bOr6OmWgWkPzG/xW9FxCZ/3kOVmrSs0NESA7yS3GtjvfX8LrWkPuKGcs3QZIRIIfXdVn2NE9mdAk
Pf4PDdvABNv3vVXX2BJkK24NqzeWJNmmV7IhZ5d7VWVqgwPJtuMzPl3aYnY1sVuePEX2ZXSgUfGY
2fdv1rumLpBjkSz9hOzOp/z4w1yuUb1wGidOE9W6IFQksw/NX09j73zSXmDhFgyjy2jGQOPRitLs
vnsuxtt3X4CIlkkH3d+C2desbxnNtoX979kbdKPnTx4Iyvj5q00Q8OwZtIpIlNT/3TdsXosTsHQq
DOyPUlByy9OyA+4GEzdLb9BR8sZg9HdSD+VXvnz4KUfc3MKiQdyxOh5k3WfNMt0gLYYZCzZQ3TVo
TCGAZqDj7MoYOzH5cRqbhpF8dUQSmgpUJZt3DQJM2w4wydTZ+MKhRmDhXtn5pi3CaeIKcbTBNMzK
zVeicbDP/ZAQGwCk0d8gCqywQYM8PgOe2a/UAg5rt1iiMAb+5tX3LYucRxsUzUNzNdZf583AeuUQ
Io+c5RCwegXAurTP8LhO9yluSXYjP++sawkBiCh1ksG2TFc5WOBWX/EO7rD8UnZevLzMRsznm39K
dy5bbZCD2Xr3CYlM08kEQZ2WLS09XTx4ze2tBArBkokR8WowHY63gn8qTkFPdrzN5aPMh2usoY03
66MeG1fMdosfK/zm8IwWlHu+azgjh9SPBDzgpshvOq6ZOAqN1hCCRt76EMoXWL4ws+pnNYIWuFCj
bCr5b8sFs3uxWeSpVAb9TKMSNADe7fpBEYNj6+8a+U5VzeSVVs5fuXhF8ABfQVuajsAXahqcAf31
qFt6VzJ5fmCb1wX9MRkm8gQt/BDmBCykfdaC9Yxpl/JcH9LSWBjkt96M6EXbB1HtqSNxR1CgnBxg
dON9yy0QZMmHVhkZZ6zY+8YvWJzf18RYHB8isz3hYTg58lfYdtvceuX6T/4+C3/wUL0ZIEw/6gRy
D4XfqQlGsOi/EXNa2+nPXQrPJd0rrxCWzCkMa5MiJHLhTYfhDwGXxYDpqeQvdYFvOGkm1SdwT4Qm
aQz+1aeDfXtquE3vQeGGNWwmEZaiWdlIjtWBZLfZCIxpdHaTc66JnM77ita4lEXQ2ILanGtaTgGh
ygOSXIwfYfYw+yZUDHrjGfvyqA2w+j994TUg7EcNvGHfi7lHjw4Hx+yhWlCpw6r8du8/bZuvUM6n
jwKRqA5jMfj7vm0bRn2a0mq20Wd0IOwqu+1JnCCk7EjyT+GnefReuG7bvDpupdNOytBA/TUcBfsc
3dETgoLsH8U+soDn2GY14A38PSqMWXP5Et/gU9UNDucIm/5fbhqjQd/YAjKkMxay9Sh5Z++vLLdq
U19RYu3WT5GNPyi2S+b9JG2lHA6k8aMim89Ra3/r6Fe26PICY1vGU595q07T8cguGXi5sIvr2XLV
8NwUbSM46gwaBdm+UknBrSEcJej3sgVvngoWlV01uMLkp8vsU1eDj71Z1zhn5xmJT5AnhBtE6NFh
JpEwXnSX+IMJFuqq3NC3ftR4m0hRWv4s4KtW2JVl3eDxkQUPTmPGAt7bDkzYM3yS6gKqdWj23TJy
1jkJ5dbD/GyOguY6KaLBN5YwSDj/5Z4kZXPB9itR3PeNhm1acTezKTwzgnpLLUrgCHdEVhi6kY3u
//rS0uvh9FypdniLOArWLxHAoyrTFk7WQ0tXs2yURsU2Mc77+dkyefR12vzkluMcN7WLR2fDw4f+
Rp2gK5ZdRUa8Mucg0EfMNwLcgZRBkX8C4sSEJMEaG3S+U3Q7I4uGTyqc6A90ghXorpzZ78dWuxTo
EmJd5lxWcXQEjoAzl/2JMLyAP5aj14OVO8eXL3Gd5NjdYCPXDLR5yWIFObYrk6wLwjW/5+LOVlTM
YOYCPjvBql5Yen7e/TjBXNW2Eu4KdM1GW9ynvCXeVCHqa2se5d+ABknzSATOqOwPkCt5OUAtISeG
54RST1rLEkYfaWEw4Rhh+1LeHNnjldeClSVNDXRejhP466g3sc/fQ8Jia4WZOQgEXvGDr9l2SBjd
VqObXX0/2pO1Uu0U15pKyJF6H1iqCm9co6N0fWzzuEq7MWeIoEgUoYavNmhE34eKO7SPWMtj7DlE
DwUPvsWdhTKEcID7YJATTgrDGIujFsN03+p26NPnJwCQTfTMTm+cyksNrlO17FqJjb/6LuvBuNnk
25aSTrqgy09aEjf3/TPlLbIhP4OjjO+/PcA/vDxAKKgfFxRyjsfB6aZBu775dSTV5Vm2cFUTEv9C
HIQPxocEDgMPgbpXnfviM2rWBVpEdCptTN9wTQ7cPW4+yuv01uvcMsvlE+LAY8I3X9aL2VOMDCCY
RggUb9PYtBp+nWuyEBr4G2LWN9ZCzDPdh6AK4ev5TcznrjWODpw2M548RFt1SIz5Y5ymWxUlRysA
iEk5OkDDeqFCFRD9w2sj31aVFv8C4aI2tSZiTri7kh0MHW5XG26jbWeoEZNHmInJZlGcTxQFuUcO
g84VYChRkWXqdbwZioBb7A2L2UQPZDQZ0ZXif1v9q9TCXXgErMR9b92Fr4QzxvolkVed7jJ4tN8E
eDWmx24XBVJBdJW4Wcva4w7TXpelJkdIWdWnKFPZhTRJankSe/Cc3kcmoLGKx00/xqVIsmE6Y8vK
ffIc65CrnTWL4XLuoiytKjQSZQynbw63qBMNpG4o36zAXHFkJ03z5+8uMaMcwoTnT98XslMkWahT
jgg2eWRpQEpCAGAVlz5Ybik05iBVBnkGzgDpq/jOLE73PQ9MgZsjX861VUtijCJ/ehL6PFSB4WVP
WyGU21UQLpUTQzcEfbGpJmLdG3ajYTsUbDN6O2uW8wlEDo2bHgwfsxQk25t5oQ5qeXrvmYDbEgvK
emdxzKxdVPFttfFJ8uHrJrfx8aPMUHhm9IYTwfPdcgVoMD+7nFbwplCoNr3uLqyXYsGCSee875qE
txSXvCw5o0J6Ue4wVRBeypfRqQb39Q6K7mlb7P8YmG1QcMduCkPBty4ipjsm9BjxiqeqnTLLLIlV
liNdY27KX2PXWBNmIH4fMDxzsin4LXM43kERqB025h043qO5bHVe8uJN6o+C9lKR+2WGSpklO9aa
L05z84dJpH5aJbxK9D22prfS1URi12d+KMDz110waZnmKoIJVp4CoZ3QpM7JCPD8aIr+cC+N99Bg
iWnDLA7XiJGc1ncXE8WnSwFUASW48PrQEohGKTCqbGnkYOJCumNGX3i6JRB/x9G1Ox/tZuxd8/75
2qAmY9JlgeUQjna+e51ggE3MZpXlovek8M8DUjwTZ5Zzr19s5X8o6WI2NzLBq5rSqn2oCLQedM8v
Mc47STmkP8sbZNAVOnVT3AyHsTCdO9ujMmrmrhsJfUxZcY2GdmwTB07y7uGWd3oKecLQ19+itr0y
edxyyDzEo8a7K1y4INM7+IItC0uVL06n8Xe3+1s+QxwqKWpYG/r3DKi++t4niDsWtdUdaIdwAEk6
k9Bi9uO5L70/BnTvFquksncbN6krTRPZTJYvu96pCNFPlyNuOcE51AGcN20t7yiXp93nAYXs5Le4
+Ql37+/nmNtrlWfKNKsCzuuVinDrLbLoGPqtEYyt+DJYLJ92eQ+vBF9KofJenF3hZiKMEY8DXdmh
CQbBasryr2pDZ/j9z6zShodYhDRlor0m0YVZ8Bo4JFTo9MFYPtsLDzudaVZeDnG4A+r9DG1ze8Ka
YKvadbt+W1l0n9oYbpSCRXh3J+n7S39NTa7Rd+BgdQ8S57RJIbwWPlS4dDjv7y3YXpbpOEVLBD4L
rDa2B7rqMUIKxWcGCU1cvOJ1a/8i7xuhsEppuTXf8otVmNrCg65al9HRDMeJoamZvOorN4Tn01Gt
bKnkuw7FhYjtUXZMm8XDFsAEGIK1YU8WHCDDhf5z1sYGUcCvVTTXVQ3ULBiNPgxxybCaW6XbUrUe
RPnK7BcxCYPgmyl4zd3Gkg4GqY/RB08qcMmNiJEDaV0Zwwm/lif8d2Oj4WMRXlMcX33O6mw5amzu
EmZjOYwjnrIZd8NXdu7Nq0QaeBOGK91iz3niJL9U4Yu0bdHdZHc5ejQvUnhhbZZv8LGPgZGGdbEb
oHRjCTMB0ZWKhDgpxxALsdkkT/IAOhnwTuHzBCLFHaLfINRy48aSmYCnbrMCd3VHPr3zNsRCK/PZ
IspTeYvdWmSV+RF36DHda7BOTW92UVk4/35gT6eW8BPwRWNE9jRg40iT53KTB4F5Ssy9FQDCQ9qf
wrbYzVHd+jsUr76A/YYTA1vU0UK6eF9D/blgvY323vZQzbRqnqQb1TAFEaXokPPxkF7Fuj4LaSs8
3iX6gmMc8pWhT4xi0XCPVDasYKBew2b0HEgPgV96MwMQMsBdID7txDVeoJyrkuu65KSbsAsK5fLT
+ReXgLdiag+EAOS24BDxC890VPQrMtJ3Muvd2AhKUF7X7zAYncMg+U97r4uIHYwazY1Wclu8WyvB
QwkNcjOcE3mxKtYruwqqBv+U3F5YZ5LSCpqc+/O+2hcy/CiWVSzFTsf9LJBe5netadPx5SgB6aJt
kcx+qSDWE15raoB6Jyh7ryuVta8roU1QYQ6/VAoeyVl+tSamw3EK/aVS4Jr6YYRsPyTQ1qJyAY+e
4XQK2NPT31arU7huaz5HJCUr1ikZkAv+nifCTEZwa3SVk5bWLN6/NvIrL5XZtPPC4O/M63JL9XHu
/pOOO63CD047TVa5nl7yjLZzmarPTZQJs+v6JjAsemYmmD13rUmACLyqC5n0RsHq96rRG/pka9sh
LsVaedulPMQ4lYMIImaFgduA+/5wM3+ZuCctL2TcAoq4Syaw+jDacHG3HV/s4r0ZPoFoB4e2Jsno
YkXo4DY9weYOCnWlEEb8uOL55JuWk48B23W758jsazBMUlaK3BLLdS3z03PR9IH1g11wfZFrNdXR
3/xcQxV3KwubjNnUGgytv7+DBbcOcqJ7d5s+N+ADNltA/RTv2vxCQwO84rtIjjeIccSVtd+TMOWN
EyAXaZOTGUCZ0Q33Sb5xZCdkTGDdXGygEy08BSderB5FZA7d+SxsS2JJWpA9zFBBAEwajNxc3Toa
HeqiS1XeXx1LsW2tjHl55sB/5cNJjpvcZ4lIukReOUyuLuEQKQ8d3J6hDPE9nOghCwzp0JkhrUfH
WYF+5YTi6XS36yUD7mNP4AJh49BvER2lwhIPMLatdDAymXrhTyAZnvd1faLNmuvket3jfX7BYGx3
VtGW18CXgGsUtq3822y6lUy4yNmbRR0T+fWFMlAB2uU3daN4kwK5FffvdAw1+qy82WvuN1BCdl7f
e7esSJRHCxQKM7TgUyIGuugU70z9W2QWk24DQaQHNR8p8LusA59/9Sul/uXfQU/uP1AApMND/Wbp
FY+7w0UGbNsG1sD4aqrnwXSl+hTwkKEqg/zTLHNWSOE1JAbpVXRMmJsHyQtUL/J/+cvd1GXZwLem
xOY19Y9Xyk7VHBoBWuQhRNdohkeirORsgogz2CTG0epE5zTS2V2ScEzQuXa4hg7Ug/GJyCmsLZJA
gPZ/d64MqraRodMTVgAqG/Id8EiDhA9MqzCbGsmnK854f/IBY8UGxNpSg/U8lIMrSpS6PW1kQmUw
8sOMFdrsUwjoSO43uJBbsKbZQuJFRHjBRvZfUGfnNzEkYQO2DiylXkeECMbffY4FLW8veUxNXgK1
kJ3XvIHD5Q9dDQmReXEibdgE94kG4/5X29ib6bpvfWgLFR47i9YyH41i9PMIv5JyaZX+DOIAFKJ4
XV3oqGVWTE30brtZsVGug2UEeEWgzngxK8hkBn0D/5jffZ/uvpmPkvbp0S73VrywyO14a7UVIrZJ
3zWlyE7tDFRaEGbq8FWWzmzdpvlnrQjQGxLmH6fpPmjJNoUT9oKhGxsYFqaxgA9EdsvwJSZcKvvn
LfZIXH7qR8W1S1hYksggdhjcNO2x3AdH6NEkNVOtan1ZLMarwAVK9VnAWqKVQY3I9K6fmenMKq8V
4vV0K8dyVsNdCD5S5atPhJEfDt4ZhYh8QR7+hawZ+zAhCiAXkWwnY1ovT3Dn4UPA1itrlb+K1e4A
zL+w/eicxuYMqPLd8VkM1xpcXxu+Vs8vmJuiS4YPKLuY/bNwEMW0K2YqUo+Amx1fPkjiPdwMrVzP
Ouo98gnjkTZWmZcM7wPixK1jZNfoR6IJtsM2Slzf1/saieXSFWkN5tCbhK6CmOteMEfjEte998CV
63QI53EarMG5uLLcgeCwdUtPx+d+WL6XgYhDRYVcwFZFii0Y0KBxFTRVCZSvsRhR07zKnaBQ+zFK
gCZ5cGT518C1Con1P+dWqbz6zJxlXRCA22AMPPYtQjoifz4+l3ccbHGKx/lZG6koeHwMNGuS5F0b
hmDT/tKuXUpgew9lN4sG1xiINiCAOOQAcZm2V42jQaso9rXXqYLEtdkRMBNN+8xZqwip2vJ+BKRs
aZq2L5WxWjhKZ/5zD2atzvliXfMX93sKk4T5s7ib/hjeUwvtPz0d0ydIGOPRH0zsgH/jNzuB1Ivf
PEeZhAHCk8fm8DiT/ghD+Kp2P2kzJdazr8SbB9LJjW1ghLfv58nXd7rQ9EzeQAkMaL1+BKIqhA7h
2iMA7rfhhTUgCAOH/mkKKchYiVoHr5xGvAylYO+Zc+N+cDe/8HLu2raBLeI4lTrnMf5ZP5PPxf5w
kG4oNZFTFHYRyf5mBHbPHhOop/uKgSYi3GoTglWv9vsmuVQiiy3C6oFV0Jm5ZPx8mJrIn3hyW8aG
d5nDUteau9qTXFpSC/x8cDEf7xzGs0f3nybpb8LTBKASaiy3VAn/vzsdBKuONwKfRwoEWu2RJyBY
b17djPGJOEpSMAEjY0vRct/Im9J2Qhk3nYq81tGBsVkvUAK/z/Ryh5Bb0dGzd7NZk1Cd0SGxTsHX
W1PHn0hrZTCX8DKEYHnVzVtexfELZT9RxKS1kurrYbfCOw5DMIY4qbTHu3hRY9EvjhCwzxVXXFaU
nGd3lHJ+jpFv6xGlYxR2F+fqqNtC7/JTVFt3631Qp+FJ8TKdz1fHd6/OfgYgZDDw3uYuGh5yMvCL
RA1hahVw0thk2+ROD6B8I+0EdYl8A4+myPnNV0s1LZRuOwR6KIJF4amFvsMYo1ZKQtEVbCs6SR2B
doz+Cdt/rY1Z9Koxh1ZyxDqwtfcVDLZlsNTBHk00ifWGmc66YTF/q8ZOfZF/QoRgvIT+x167Eybt
R65juifQHx0XGcA64rOJz1ZkSUWWwkV8+tF0HdpwvHr858FtP/Geg/YeEPd81AKKY8pdvz3DZ+LM
7O/RUYNmhYKwgtQSWVKTXjgHqsQ3FA50oGHgpH9ZHtczfBO6KzPulJHvKv0sHH37RDeWAzY3v2cb
Gg/AQx2i7N7IAqU3Drm4zUlzHWSQiNdQuWS7vx1K1hpAViYTveAqS+tbXG4D5w6ixkjEPx3Ur4xP
d1nVI5Q9k1/mu2OusK8Y6x99hzy0lmsOnjSlMVRDP0/rxUR4ZFPUgTPUDw8Ya4KRFuydqhQ7StZP
pbUlzk1URQkH/LoX+kDc04+UgxI6CEx2zSiX2bUvLs9nE6l60rjLINzgHhkeLUohKDpWEqT30Sz3
EOubONiRXH4QaTY66GuzSpW7U29uXWtihCeduXuamzKYGubUoEiAvMbcSEJu8NJ4ANDi8Aq188t/
H6EFhRvdZS5/fqaq3QBJztfTTeN5JgbZUqwmDsL4hDHL7dKPXpYwjfDAIEt7JhKdVCUqjJ1K7yGT
+Yy0u3yI85ENFvV+5CtP6g1W66G1KqEm/I0+gZF1NNpKMpcm5RJqAsSoZaf96Egmqm6q3nPc2pNt
bDKg0o3dKY3p8xPvKCc2Avygee1dXpGSxqyUbICHLjMq3Xs5GaRhxvNrBUSR5silmZoEz1k/zY8v
v+5c+NFPeiZ7UOQnxa2H5bLKeBCUenwRVzOWJvda4yUZQHDj4UhuqztDLkPvv6caQ1XJlTA9qTsD
awH0L7TS3GlJ6q6fw9ThqFWOzFgMHrrbucHZjJvTh+C2Z6YVH1j5RR8s8ZOWD3d6BXjACFTGJqXw
mPi/UgymYXm20FzGIb3pHS9stbcRgfOH+4YEXmN5QtvnSIAFZBj++6vrxOHn0ml4KWy74whsUmWQ
C/E8tn3FTHGqJ/V+ULwIjCLrkDeGyfJMcWQpF3/09WoRXFhVx5WlAFPVY+uIkt8F+sxhf6eaIl/h
9hqqhkna2ZlI+0XvayNCtOn3+ZYgPRtDfEYcQIkC7VCBsPLAIYF8XsTOwR7zOP15zFcv1Pryk9jy
DMu6OQTohUi3rysi06H8Do3yAGq1SBhDjSqRyEASxA8CarqVLNW5c627x+bnk3PT11XaJJEBwe+8
Sd+2wshz1iKKMOZwgcBCrbktQy9dtF0cJJzId7QLbdEz9JTUCdF/IZNfHO8jp0SVivQisH1o1oZw
o2dQeDwwxXHgcoVo3D8QurKK4n6wQPiW/0jODMYR83hDLRYjcZolZBdLnBRxTmpC8+EDdXmZ+bxW
NvravS8O8LGFUOJeDydTkCTHCcuEtHnTTOS4UpfDl2Vk2OdC/WudI2iyf9onncqYYdbN01yotNY7
A1pBCe32AVO84vIoBGJDeJi8ZMjqSzqlxrm4spZiigz81ehoUwsdjbaMLqO8Tu05n5cA9Z758EX4
AGY5QNwbIVGMvWtdm2UudmW3TUhcPoe4FNOY8WoS5LWvyZiCaYYT5WRZZfg3v/1pF5gK9TJrzn/i
2e2jhHmLLI0mhrX8lW2uPE1dBGpnKW8vJ+7nIXgSOaJu8gaazpbx4alfcN/3l1m873LMhRe0ZviO
NvFIn9vo1c5MGVq1Ev7AUUmnr5kYdJqHIrlK4aBzctImiQ//7YSHdSTvzOXkSZveI8D8UHRNKfFv
srukFj38U+qgdhFmnpipmvrbLXV8C0AstRkcG687aOrhCgnFaLYakOvQrxCekTUdiXAudvZXWcmS
vMBipQYW8Dxaz+i3Q/iKaxAcAln9H6xq5saGW18dqMEN/1r14rE8lY3kCh78E8wgqyELxXiRCL0Q
GSJPOS7aBBJLjiHQnoXpy+AbyotX0Z5tG/uhZG0c6QeLLL+SLgs7u6MJHPvQdjspbQkXlESKF+WD
JiA1MvPNyMWjNGIHxF93dk2nP/fao00Rh567eCPm2TBCsSvq/ny6yxe80WATaId+SqXkotL4fdi9
4GvnnowUPytNB1scwBYiD1zZna3f4jRmW3hKlVpW0lMSIUdEIZUuS3XtqAPCkghx05rxKMd0TS/I
4YKD2eqfD3OxaxZcWLlRP0sGR0hCkR9NFKE99jnlENVuWm5NthbnOoQkNJypwP4UMI/YgFBWYcE8
nKMf3IQsDCpL0O0WweDgKE8lBYre4I4LBIJFSSSX51bcdEEVvgm82YtWgsdXIVIXIIq2K4PfDIl0
u/ff9H0uUOa9k+sZbHMuNuE8Oxv01mIFKd13D58h3FM1txNe5zCyzBYd3HWyGUL1XdQNrT4fndlb
WgCPw/CwAT2wRDG2HoHmz0GI6zXCHrTWRDSBg5dii0bUjQnjIp3WRcL/SrZEsDnQCqEpLQCWTQhL
QgL8XrvaUjF9OMBNWH0jemNUhI51lGXhVSHQ/K8JMP++h6u61cfi0OrJrGjmp/qxvegFVdjl8W6f
eMzYprTt2KPsN5Gqm3UKhOD7s/FMjLRgGE806OWuK77fWCTCry8iGXHexIkbTjvRbjsKD/Z57MYt
vArDbd2SAVsXS/1RDZ6zhPxagzI24EI7LJSMZ27lVAYMl/2z57ktjNg3eP90QP+Sgg/TyUOoSdq9
Q3DoCKmPvfHHkoZGYsuJ9KPRKGY+Cc6/GpCpxcMsDeHV+Bpdd9qJUQ1NeSbQm6qewICe6F9ub+zm
B8nrsiwK/NdFBOXOThVaM7Q99KTetfIINu6AATzoeT7z2mqYZ1XimpNpC/+D0zr8EoMr8bnxAE5V
BVJ/2FpUhk5CYKMDuOwPtWzoOfk31EnKe3VrLky6XFskgILSEQBLzwB0Ul4pjPE5IRGpyWVvA+XM
tgtWX10+A+8wbqE5FTrUAMw8P6VF9FFsELGWrJ/Wkrx8zaCCyKGHRXRCMROQj+O/AOp5hljvfXRR
qjJPRDqhDgQ0iZ7j/axBPl/yoe8NhLc+KhHL9GXUYcdqt4fVUQgkHwvgoEkOzX47xTH7j8RbZMJs
fzY6kgK3Pi8bpc0u3JORHu/dIkxRghcpEWWHAk2q4wcz7R5vAR5TddBw2wEQYhm4jU40PBmWINFa
pdjN1o80hQlksIfCsrS83WPvj7sCmJ/G2kqRhrgx4/N7HuCRE0bFfY/+pSRxMWcgNYd+6+afl8gW
tf9cHrTjC6lPzC//chwyVxMKLbfW+LXjK1WATVP4FzOVVdCyse5B2RHgw1x30vhv/nKen4YqFRnU
7dWgtAhWwJakMZPodSlS3QUEE4MI7nKHXb9vt+h4UnwA3JqK0WnplcTp7g5BzNUHPGtkr5SMfhBG
7MjlD1ylP0RG7+GKQsf5XLzWWG7jGhd6dn+0cpWB8px9DQG/Y8N2VWqI4TYwjHh2orpkfX9H4m1E
U+RFg3EzJZAB1PnJfJX9jPYebOmYBxruBJHgDv/seFW/MbAT+btDtIHQgryruzgTxspZy+hMXzKC
KRXkC+POjK47NHJlLL3mJymQD3wu9pgYPP0OUIHm1gP+fmldZvP8XgkfW76qABBbiOOs7m04nqrn
EQUWfVkh0PgfwYbkDTbfU1seUcdTq7IkfoZKWl5/oJ11+V4Ma0n7K1v73cnm339F+TwjFMho/SdX
xMQViLHQR5mM7zrON3U/6WqSel/dqsn0dRFs3DXJ+ZFFLzJB8fRnVzPRdBOX2F06irfRlVbnRSaf
ct1UHbfBRTiYLBgEs+3Yiw5MgR4FVAv43xWJgNosdOpk0c/mWK3e1BgF7NDDQavQYv/1fSo2lrAN
YIf+1YVworlMPx5imuWuKRDNQOCTShQbqUeTYlMp2acVny8a1DKQFZchVOm/y79u1TgzForhy02Q
1NY38mcrZav9SPcub3Q7HqOUGjCtdXYYAKQnvH22EKy8ioI4Z0UXT2oqe6nR0munS6EcTQ706Mji
CqoaazGXLHT8vddBsZRoZIEuHqDsTfvYj/ualXO6Hidiok1GLywOz98CRlVMPTAbEVr0ALioshQR
OKF3eXqHqw7bk11SSjklVZs/jYoxCjY4lDkHei2FIDudNnMRzt2iB29OkmFi5pegXzDFEskV25yX
Hg9PPTyM41CmWmX+9QOJVeGYXU4f0THBS4BcQt8hgOQ2OcaFMcz1EqzVr8FHorL1iNRmFkhEOJGN
OcvHSL3xEYCWspqW+r67CbZ+gjVHV0m9Pah67ea6REPbskvAFB7NSvJSMMPq/S/vNR55vlBwdfra
eB1l4IGM5mg5L8judZhcdb2wfHW8aIuvXL4YW9KlwoYhXoE4YIY/+6QsYCi+Dc8rCl608LCM0ss/
9SD5bNYtmGkeWc0Y11prarMQ1lRmiNDJroShlqp7hhaVAJUO0Lp+S1kbqKgEztkdl9nwGCnt+Arl
hvfymc0MuDw5Xk0dBOYfVm4Su4aaPp7r4r9m1UoJrbD6o+bB0DZiwnoiTY5XvjZHXXmdwysq5sBG
08W+TTwhYsT1RMDh+rxm9jiMSPavo+zokqfH/dls+jA8QwXDeblgUHklosLbEWVQuhROeBAmaFRj
hkCSCwvwdJFyTwJ9cDLcQa+1GK7O1cE4XTe/iXQcTuP3ijR2UoTKD09cPCaxJfYNzuxBjlRa+SlZ
DlClUk7TJ0u1/gJ8Z0KuoCDa5/7RRs1a5C3a+DngtNigYXnB9KlBUBe2PTHoFIpWoVIZBN3GkaFG
3+hcBnZRvH4GtT1dpPUCtPts4BSMI+k3i3cOYZ7jp0psiKdhHpb0ZWwdeJ3n64wTSYfwfAadpk43
6HzA8VuBXNRrfFkg2nnS3HCewn41tYmMrcl1HF6oDEHqxjJFUGwANr1Ncht5MPOmXL8rZ5LhW2AD
nPsinkK+w6R3ZHJ2Ji9kFXxjfGHEFU2+ElhcW1ZRxGKOm90qePFj4E+h7sL4Ej0z5W4KNpKjJ1NX
COZgfWgVWN+YT/CICgV2nVH40wnLZvTemTo1rLipgbgTFpuNb+wFQW94v8SX/EDnSFbJqHrR5Diu
CMUD7Ra+KZmqD0Ukdj4EpkI4wWoKDG5rzBJYPNw4t3/ZYMbq/1T8VDa4tw02foY2pcW5tMxaYrNK
Cc/qYg94c/lCcYZL7hkhw/T3xb5b02AUAGEGtuYVCTpY5h5WLjrKUelhgf4rApZKWM6SpI/3qRNP
Y6ZnttZss4RV19P7o+xrKXp30Wtq35YGzkuwPy2hPw74YTR/RrSK65KAeZasdut9F/o9h0jrafTp
Ko7Q4jnTXJ7ka0yytoqc4rEDYJDw9E9YZOlm2n23dKYypNI3+acz6pL8atNy4ZYWLY7TaN9/QYG5
S5IbyWpShDUisSHNf+zXMRBgzkY5kWJWFaARduy4ehA6R4LlFLgN4nZ+Mr4LgtZh/TUFe/4dGMxG
1cJ2K1b7LqQPUGNnB+AnxN79ZMMZrpJNDUOq15mJiA7L5jp/mWZJ9eBFJkOi4hlJBqXQuPJMiZW4
Z21UEL4j7pWPd7TIiL1p59sIAflBrUS5SQnj70xaEJNPcY5m5ybK4VQUmu/5IOWddd4gMOyD30tm
kUZExX3LGUfcC3F36+43R59ICbFvZPFW9Hvys+LB9XSb0jp+eOAZUFhhu4HVJ1QbH8/e4aqmquLv
FBGZABuVbIznlN+4Cvcbr7yuMM1NyinRCwMwEulLGYiF3y8o3KmKcxfP9zHI6LCyK1COPM0sTi06
krRuoxFBxb1L5/vhWIndbktOSvghHYoa6usagtrRLiVdf2Qtyg5CS741oSpaD6vD53SJ89KBj3lL
Zq5GJGv5fAo2swKDbQZw9v720FWmNrmvU+1rQ9fZoTIEEN+q8ImTUok0ANUuh55rEuTFIyzIgmBY
bshwNApd9dHhnIKUGsQ0Ew8VbdTKOqPAzSm7Q5AJH/iUcTZAki0eyg18TuhOCkB46Icl6V/uVvS2
YhY3kxm8fbbjFwYTVdypqMwEg8FtAy2zUDqrocE/mlZk1bh2XmvfYRSQpBfVxgNanj1wAwAOBH0q
KLb6duhjrNoTNrkG/vY7yYXKvxbbd9L7dYOurIlBxZIunP+t/m9CQsTqflNs6qZWtK/bnrDLoJuX
QN77iZiQ0z7iui18lgwDVeU5TNMMG10XKXxEW2+0h7WZn5ZXJRdtlsHyGwB5yQA6NjsPStw9X9wX
KPFV7J9EMkKhCXXVMYApfjrpbyq1n4vnyAXdvJrY+btzgWC41CxcVUnedAzyUk+qUWwvFZplII9z
zr9nQhxoqKzeDbhpW0GYpogLLNQwi6sTJ9D+uiFp/lc1AOqXOxTRxbf2VWCcTnUThjDGQSjwmjOu
OaYRTaMB9zqt5iAKQSkmHmr+xhFoTjy6hQXOmFTNyqI9ndZ4h30ZRym8ecyD4X9oS245AWZvBM+Q
vi8Oo9Avn1HfIqwAV50QUe8C0C5BRdqjCkKwllqp+ey4FSaPHTZlwLEMQSkPIFbqrcwdbqm47fze
7vodU9/D6b7z5R3cXtC2AcdzQiK2o6v1nS7MKdsOMD0/WNjjc6WK/umB8fb5+7QOl+4L5FZiQ5qO
dNref7kd05oCsWra6h0X6xT/cLgZJe+1xksOaXCcnj+0bdS7ZNMhD/Ews1pfarhDfzwzWjbBlqWM
w2GA7o30nVF/uymxK1hQbPlymdAKMaofbSPtaUduLkT9O24k3C7FyPatT/ItBts/vDDfGXXasNvt
hiDab6JSAMVVT+f1ESvgLqPGzd4Lw+lCuhrWfDqtZ31RBJ7P1/OkL0wa4HeGKa3xnwfQFSQVI0ZN
ItHIaCMeoEgPCl31WaoZJ/hE1c80xrlOL+lBnIyg6d+cVcL/0oB+2R+8QxHqPkVm5k5YvFivhT4C
wtW9XwOYi5NLYBZ2v10FdpATvn9al4JK3aC9sDnUENyqIHDSZbcaHrph0O2EgS3iAa16z7V2RGvP
bP70sCsK7NIRxUUkGANM+jF80oxdmYt9P1TSgVmEFux8jxN0BAPsYFgj9Kh4fEAWZTtPQfqm/xR9
Q/Jskb2ZZyvHKyu/kx6Ou0we3cmnQlwExtMd2N+9WKWtSG08iCAMaMaGVByMGwcOz9C/Imk/sECV
EFNuwTPc5O5kK1BTaxuQi9Z/pvA3BtKEu9KjYFjhHIXZXwIrKxo7gT/UUqdtoxM0/1KsTbkcuzRh
bmgnoKyCXY+zdjjYh1oBCDLOZu9UQZNfwKYm4/a6F3C/ZjZoZ79UpFCfbZ/p5jEIjNXsRblV0Rdx
2v6gF93mZFs3APr2ay/w9mLp6L5Sv/xtn/QRgj/6KnE5ODkJ5EKfhezb/5nTUUp8Ni4NBB9Jc/cW
yLZdiFtWYaYVO+LqN6oEVC2hN6V2YkRVPKVmrnOznI62g74VFV2j6yTpL7pQTzwJkrQtEtN9sO/7
H4yfqZvTe26qSOyOzvqtwUrJqPpzfDEcRuFjcWJ7l7KpR56FOymheMExnpRZrocBGDfKnoSb5+Be
9MX6Cnm296+evZ5N3KA9QUiEtq45xi6VwXHgtwhhFzQgRu2rE6p2lWgNcW9IOBQREm7RyXZA6xHL
paoqcTPQtbQCtimsPRaJ/d536h1bxgFYg9jK6VYddBtG40RfnFj/Q2ay0sw3DvFHKBmf88Df09qM
/OMEkc+z4MqIyXGZy2O+RdDOy+TWGWNmX3XZLYHqrhr32b8K+U0+OJN7/7ttB3EhBmprDQCdxdPs
Tmo/MJtbtCGzomxy1k8s1bJu/s2pFKshnhtCZhVlae95Ys7oEr5eomgH6KRmoAfejOe4XqWadnh4
3eTAg85s80Q7xX9mgcBKkldXaYawPLbMQ87hshAm5hvfEWwwsw7JsZH0AV5Hwefy/HihZcOWc9Ur
BJw8f+2Th4CWnYqFvJwKq8ILIu+jbyP8T5mhe//xo2ob02JE/ZndLgeazjEGAtBoFuR98DIf3W3N
loXGQUZb92VV015I/Gfj7pQcekP+sW4Za5sFY4jxLv5eRNlBI5wcsON4PbolV2rNyiU/bHwIy21m
dz7ft7Rf42cdRcmH492/NJ3lStqscxCJEZNAHcaA35tEeGQL1TczneBi1qzdhlnB1EYXt68JUzqP
Tvi1RVGoLY686/O+cwO8xj59K+jKto+DqgnOSuX2zusNQ5Sj8LT2GgAsC2HbKRPavuDoChpbGzET
uWZ3jq08pj/W8t8TWcry3eNbOyWhiWY52GXiD8KeOTqtwF8LpB5db4k22wT1aM/aj21UNmAGcBEP
BRgxOi2udk1ZcDOAx5oVEvEks43XUKpCU1Nht2A3BrJ/h5E/f3b/FVcJ22BerVGxjpdooC5Dtn0+
Y40jci0YMLvK0okXJByIVpxP/lEDGWdBb4rttq3WCAD1BTmzybYLAfu5tFfDOXeSAVcLxKUMykzp
eBiaUe5hMRA6EsqRfd9qlJmXWKj7yiwXAa2phdHbeGf0CJ8f0KSp5EMVlEG8CBZ8TOA+gpxxCoIa
7qvbrUWCEx50hx/TXEl/shr6ChrykG87eL/nOKN7LOpjt5SOFAk3DXy4FDlzU5oJ++HuQAXdYbgb
FIX11Od41HWkC9O89bpKKDF5gG9Bk8Mtnoi+DeqQFgeKdwFxeNr6CaGnqNW0Se21PUiK3i12t7/o
ux96CycMk1NcuhpPJd2lsHldNSWfmmAMpZLXDP1HwAD2Jl+QzZxbM8PyTMr/PxtWy1Ni9IRLWvns
3S0wGfpj87+Bl/WHeoxroxO79A54yLAYIM6cM55oaNLcfxxBPXNfEP1PTWQBxJymmudUk9/kg6aX
MJsK4h7voKIhziWkrVe+AmgddIRXWXKUXWOEui70yWTv5oWHbtPxyVu5sk3OhHA1XJ4Db/LlF0+b
8zY1Hrj1cL7+xR/NsfMPHbPGGzLiHgFD7xs57o8rtVhmXJA9A9eV5Y0zJpOA1m5UetCKtRKOxeGw
C0m3HvuMihu9el6TwVruheYgcuvHmABsZTRgpQsVgxLxjc1wF1c5fh3S90xxENxOfaQkNjy0G60Z
qMEOUsE3fjkkfHDOZc23uYZzSYesn8PK7da+5ehvAwgy7/fUyyhEX1bjUlW6QxvXe9DKvG49pQmn
1Qp+JjbEGhNvU5L0AegwKJnenQqJtsTgzs/CVxEKAyy3e/o9L+HxO/4j74hF+xA+ibg10XFdKN9l
4PCdgv035j4v/YBLCKaWjkg6gEkvuO4vf2ZIbJV+4GYPOOGBkRDqEIkemwBGtDDGAHQwVHiaz+qz
aXKTJi5hrLbPV+O+BP1KlqYNa4NXsTAHMZUvXvu9vs7ZgmvY/PsOKp800akGxcbG3bhLSzNauicv
WnQqpHz8WpDqRsdrqKT7g5I8v1NurLGBeMcuXWsHmQeC3dDR3XGdIdrREyO5o0mThU9WJODd9HXs
70UT0T3EaBcx6Zb+Yfro/gwS/eysAK983qWE22EtXx8Mhhek0D7c3HHGVEAZ2SYh5pu9DGBaV8gQ
JzQvaaIxb7Cp4XKkPGWGYEweWg7h54r9XZIqhdz/e0ju9mz0P1aukwnpCkXdRrRgTQVzWgx5mLYZ
f41NRAG7lGY59PanSd+k7znbQt0cNZeOb7F71n3eq/77swAjN0173dQp020ECb8no8gC6BogDw2i
XNeh9oyUIAUrk6P9t9OQ1hqiNeITD9tp9hkgQKWa/OCpyV5KClPOxabtaunwHeGZbLJ92u/1ZDRb
MYeZOnE2p1BLQOnPMwG3yUTikie6P07I1AWiWUSAfT+nxqqKUwt1cnx9koWFdE9hrUEw79rvAZEI
QhN8ZBjIBgoMfR+bROG1TUKIDZDLySBLsTkdqOUMTYLnFiU3FMbh28q9rYbu30+4a8nUCqloh6Bs
t3rAfKIDBiD1+3gqakqhLS0ZSaT7+XHNq5SHVWLmFtkxl8a0Cd/diddWg5yWTxqPhBhl1is/71E0
zjL3WF2RN3cNrrvJj9g4O5h1dXVOCGysSR84T84Dn/uPIdIb5t4BpQcntx94YBrsvt7qiuP7e47f
4aoHuVn9bfrCzym8f3wIF4TmLbS29/aJwQUWwzsd/l77UidXr5T5u/gsGjttxOj7NOX5CvQym7Ge
mKlqTARQJ0S8HJ1PdzfYM31ZutYqOzLuHjKZXL0Ml5rj9egnUeybL2LgEvmB8jgE6+v5V0vYfVz6
Jq/0bxLoY6UCbAliSkVuIB48NEzsCuxRmubzPH7o7XOTCK5ivTEvSWRAamk2mw1wXyDPa0iMah1/
Ui+8qW183HK2xK3YfOmCckdHkMgQLmUIvGvR5hHgP5m/uxdzR+55sWA4sOFBS9nJu9DZJwBmTAtE
QYouA6ZepJi5W2in+PYrPBk+gACmHjk4E4CBDdxPoO7+CV84HXfNZR70ymDZBieRnhj4M3CVyCRj
WirGAJFTWvdX9KdaaJeK3ltTcUE6cKWiXNMYHQVvzsgS2KwMhk7jwnWkpa6BSgba4Po05r2pNyv1
4akOKPXadPyVdzplvxMVT60wy452Ib+7yuXYUM/F1ZRcanzK2eRUueu/CPpjERW6p2wvHzHkt8CY
HZh0n2DoW8tkPPwJR1hJxfYxi4yJmW+hCJRCkiL/0WQNka7x69V6TrHPyZyadku6G+sOzSjyGSEv
NAfcckuVSN+RMpADLb70TsWl0xUIzHLRtgRPvqIaY/YLW2A7Rs2+qXPtgnvvw/dWfJAPxyldJkiM
cjbyFyLcqNBluK2oFKcgzGA2TkigEs8OjR4JF7TxphBaEd/y5LMCQHnGPICG5g2/Lm6DpINRbZlq
huToru2G/1FSTirNfOiwGiEQqD0fsMuwvmiPrJc5F+v1fRpkhFj5NZBzabbwPxyisljbe/xUIb2N
oRXiEnHenPBsve4998/tK34CeE+zHCpSQqRnyUdrGI4bZuVA6QpWujBUBi6KB71fh2pBsQ5d0j57
t65ul8N+QAM8eSRUySuY/Q+JuECsFRWSI04NdWhnl0Bu8HDgTm1uy88oNzVfUtLQDl9tHjQcza1s
YPJ+oo/YX4ZV3LQI9N7j5Cb7fLaZ1nz35xgUWPUmuJTq+/QlHiaE9YfNqM0JmiRvZMqFjsJxg0SV
n0lBOoNvvySvGOXUph5aFclE0/6VpjXEtYEEtKAq0i56Orlea4zYmiXWqt/nMFxXjYoyqnRYmXjw
emyrBpMArCiFQtHkGukhcz/KhyOi1dk8INJTxM2ULywbe31BeQ5VcH8A2irc5y7PTEpD9iaadnaI
q0XE2kU3FDfYyLx3pGJgcbc2Bj34mOkhZg7VjXJv4HoHffudafxQ2HtUIjSlej4p4535XBaNHl4c
EItg6aLDAJg8AoKLj3g0XZAm8d+PmXQhE331DE6w8LjjJ+fllO5va4LXlc4aiT/XIZq0Aj/UEcVe
4TcAkQFfm/TUxNIkD68B5LYZrGpxcJMwZVjUinS+ul3p9SdmFp4Cfj+ZFPUb/nU+FhNEXxHclzQ9
VFRDRszGNQOFx+tm+9JswY3Ddtt2XH9KkFjXR870PTAfGiEUXqB4XmX6jetcuQuOkMQJpTCR1m2n
pl8yMl8L4J23+lJTIzBBNm9tqxXkjaK9BruKqKinmuWGlgR+XuP0BpCFCT6UdEnNJ4Fhbz8Wizyo
vKAmxfenrkoWjRzS+IWU/23TG1L3fL0mm7KOKKvMydUBIrOfCSjuMJzqm1WRaVa61oaN7xbJ+WXe
Wy6+GRL+01I1JpYKAk34PbdHuP3tBu42R9qXDibpfkFxv6gKaEQUUJirYTr4zR56dAItDoPRuKVo
Els/HIoyqRnFaNdfJf6Fci7egjS3L3bGleZC67VDpmLPWNgEsy67p4QrVTd61JeCvCosCv8YEjk3
RTdqcT4FGnfbgZIaKGL9noo4w0SHLIMY9hkH9+2NNSVhml8eUtMnAilcWHvLyi/aL/FmOFn0R0md
ul6ofRw4LnxysMSW2c21VwaAA2Yr+MFhqpQEPtvei9raGSd1j0RoeGghhBT7nav0NsV1ONoXO0jJ
n38tO5tfm4Gti3/Xeg6AHEhYgBopM1HM3i2xtzIt34X0KWAGkwkX5u5xJNdt3WHs8Cv21U27rLmB
DFfJLCLIjDVCT1e6LhmasMhXZRQ6Cjnu52E6fFHQo7l5+XiT87+XrZz8OZ/n/O/thETdW90U9TLP
hSz2dSDv7GWhvVARo546EZ6JFqD9Z1q6PrSPs4la1R36Ae5qonTELDjRiEnHdgbqh+X5CzuHTIhp
Ahcz5lJUUIeSZVSUlO5TY0XkrhtgeAX5C5tNQN4AUaB2jiVksizm0psFF3W5zkdxPHjC42OBnJIu
kraIgj56SAQCtnlactakofFn1UGss3BX1LeYV9HxImUpcORn2xhYVTPxBp+iusCdSODQL2+/Zjav
CreTj89kDdM+x9FpF62kL8ZoCVLqgSBcFtQcnLovcTnyKJDO/JBHAW24t026YpAxj0+1Y8uuwIZP
QOfdhYqJjdj/9lrs6uw2KxVm03aWypNfsllHmTV1PaUZs8BZblma3Q54DhARkf4t5P2pmgFJiDmN
bPsqRvIBKcE6h1Vib7gaef7/D0SmVHx953T79Be7Dx2p3PGWcMCeamcLn91aoFtz/scPaqSFII6s
mu09/quaOoLD14oAOo2Iue4x+feTcDTUbJe5TbOOwBMtxuB+jAWSwnqxPJDnehHDIYToXCWin8Ku
xv/bIQeTwAU6UP8OJzvfK0+S9xMQxexw0tFwOo0D8J4hnuNolZRCb/1v7HogbbSmv5ExcdJt5/Hk
CKgwT+JwUdu4j6YtRD/pV1uv0poi4o/b0EPBDo8FCcktAMIY+11IAK6d29+lPGkTIEV9bNB1Sdlv
Fx1EO44Kx5Czbq+q0DFNP9zKBCnOFuesXCjOK6pIdpADr5juNIUF9FlhjIzP2G5Zai9WtPA8aQnn
64VdMQJHchK8690oH/ILqnq33OPC759xP4rxUJwQhsGaufD+ap3ENO+ZvClcuhxx8e/OGp7/ut/N
WJzSJdQIN0lhrb/gKhl8ziIotZiHCF59+UfdDfaChUD7GFwH8JweUsd76zoNI2IEBFjBhaBiTNgI
ZA9V5ijl7ULNJG3vwI277RLQe8Z8lpwDMfUqaNzUu3/iQKO35yAeedDucZfUT1ePQvrP0s4V+l/0
HF2hI2vdNZswvREoIx4exwbchsByAk7oqITdVcnRIrc93gR6mFjvrZc/68U+FTibhChLAs0xS8tr
1WDFN1RnbRQ7ply/xQcHotX3LtzqOL8TtoheJZcSf6pMfKZZq4ycuNV7ItL0o9X24AJiQLZ8/h5B
l80RojUFa+K4gyGQ3dcGrxTtliW6PXmmqIN+OddZ/08GuI/fZiPXSZ6KDnwTd8iC4B62nKxFLhYL
uS8mdK6AMTSeU/H7/8IN6W+/M69nCmeRWp5aL7c3dT++OMs0k1gospHKZAKk0xGs8UXEbgR2yDBL
cDeOZXv7s2/zmHdC1B/5EFJhXzAtyNhUYliQLxjMFO5/01SU+SLYHL9NfKzirqFGoV+vovHe3QoC
s/FBtW6o8MVOlzamXaf2BOMLuNWbqztlXDQtTqds82bsTVB4hVVh0ppPs97A9MP2FoOS8Lw9yGnM
FZ4edZQkU71GoxihayPQNPGdnI/3Mj/8CPAGJTRx4d4+Ay6Vc8o0E/8alIPvVC+jzNWtxA2L0VDa
AgJBZljtkgM59YvGao7w/N9PsCc0YT8GSR1vh5ulPGE8kN/AH5lA9lHuk9tdaY0tXhr3yBiZyuco
4cWvir1CBezBkamskKJ+1v7vvcKQ8ndeFfGdrIeAjfPzl8EDmM9+CSjT0eu3QexLQQl1Jo268Ehv
RycMDiWQ+2GW519NiUeoW0kiyrbbkUKpp9aadfmAXX0mHcmoxYfeL2ETYA8NKZiSZz/AoCekzdIl
iTkqlQT4DS7+gDhjuqJclA+pfv9NGcWMPCmkJ8iaa3uw18LjhXUuMoEbhpEtGeOTZ7RkpM67D8SN
0vBS62N5RZONpTjRoYoxRXNy7o/DzK93wYlnwsqY0hRw/iMf9ZjXnF3sGBNi/SJYfavkkUQ8IErJ
7/Q30ICPtktXMyxCMm/tH5XX76oGv/m8h2aW7+RcD8hgi5jzJaNLZxKmZFqq18oebXqpoqcX5T/e
x18qGGVy4y+W6fYEHA4Cl1v7rylraybfdhLCd0N8TugemfK70sVGzmHw6Md9iAbDdb4+Lr3BSuMu
bBRob1WTbeqYDQy2XBkTY+vRRmxGHVGi/4Yy+rZaawNWUEn88ttOOdM/WuN13sn6QivqotPbw7A1
FnsSxeknkxSpu/vUCWvIvC5xQgeHl6sTKrV/QLFETPYEK/SLHiSfXyaTZyQx+/bPJsQoYLG8Vs26
egYvtdNqELFxu1+IPdchBsXDSd29JKhq5wXws0iubBPQvktNT6y/cU20B8BzC3yumE11mjb4iqm6
do4bJAxMWRg/VpqVzcH1LgxZbWA7jVMrgjh4nM7pRh54mtmnnnKVON0ZDl5kG3PYbZuYEeKK7iuv
xwfxXI6H/MZBIjb7Z+QDClcvvbQGx6Xv/UHNngcpWaUgOqK6oeLNxp4IqIhGceKiATHAPM8Sytw9
dfJcI9mRX0ppdv/Stol7D5RZfmo1dquIP4VpmncjS5mp/53/4ikUngoKXpCtBbe+J34ZMQihepOF
LntH08sAaaNVyLMRba6HNiYSRetkCB0go+YZ8kdlYaEEMWwJm+qGrapc8uNlpOUEHMBRU2x5soO/
WKoj1KWk6TVD2VTgUpAVbQMFVn0KVL1e823KgIag0FCpKihooa55uqsXd3k38HiblBZgzaWdVHhh
dLy9kZ6SPLNeuujWQZWr9kCHSzBdBCWi591lQoWTjcYZHOQWhYIEAVDSLzGIFR75a9bIr1L9EpoV
cFYdeYhtYLCWuSNDKwhB7wCPbNTMcLI+7slcImLsvl3v4A71ZBr+kZwxZK2FbGoU9P5XixJAkGG9
g4CWjc94sZijw+DDYH5tYJkrsjb0v1uPlct707HEAMht47Y1wMVrwN0cd//Q7eb0IFH2XHeebHeX
PA5HRKD5Ly96cUZ49TxYzIMVplcS7kaT0kpzU3fwzmvLmuoRRvocPMIb2gzXZsZW1u2BikVlSrIh
Jh4DQHf1YtbH1WbPomRL+jvoB3DgWTDVcuz/1Fffs4n9Nmfs1Lb+aKi3288q/+DPOYdAwtWw+/Nu
Yl8VTXrJCPlhCbht6lg7m1GFonuDXKhKyQ1nC0LrVsak5tZnULozYpKq9hBQv0wX/n46Qs1BWT7E
R/AMwtfq9NwjSr1j04uzzcs0phlFOERjO8bd6dbBm5586KYuAt44IhQyWW5fNUEr3RdMIwdWYeJp
N10ScNnhTeL25J7X82pehLcrDn1tbrnkf/ufWnnoqrm9WBk0DoquYb5Ou8McF2bBSyEHlVxoyiQ/
dCByQrxmrU7KRX2bfpSIehbvoViPn0y3B3qiRNYgB1Wlhk/O5BQinYGBg9hbKLODZqQNUUwxA5N3
PWKfTbGJRJbsQE0D//iIeo8uQlK1+baqfP9CkcL6R60C45rkva/6rYRCxxrw/Ct7oLV9AZxsuDj6
oMiz2szkMdqkN1z9mx8rLLXUozxzBTaR24OezO6hOF5znYiu/cpAcg72I3UOzJqzZS4/cLdSUeLC
DY70VlBicedaUvzLZ72pIqEnqDg0lHwMNzmGmky5/TNt4Y2gPuj+CJPEOYTNz/IL1PJuoLQVEx52
Mcm4XRiflCFvTV+TCRlgCzIOo8ZIrgLZqPkvlGLSZyDHvyPKFnGkqHcgDKmZkfByCphSyy0Ijj+T
cWMgB4Loum1zt1Anoa4t26LuDNBo8wQIsM1+2e8mHj+kHdCYNKGkn6O2sAj2k2ZFdpHW/Ks/Tpzf
q5e/JodUY8eaZosAb8elIEs2DWSxaXFj1Hv09js+HZR9/YjVPJ+kEnEQ2Vhv5/Yh7gqGj89JFliV
z3xFIxx4vC1r/sbyv0l6Da8uxby7AUqzkTFA+OC7AfqOVI3HGj2kj5Bp1T2YKKgxfBV5CNP3KH+Z
NL8eM0JbyqXUs/jaB9ADKLtC0KKj05nFiOlpkfBI9ZSULFW9X16/j5INcq6VhUW2Tr7MYSzJ8rls
b+26nJUveat7gliKzXSqZaGJn0ZcAmz4VZ44ErQv6uikG5Xl6hBgojCHVBJ+bRq/dXMd7mfr0Bab
uC0GMhXwuNMt30Lgv5QPqxQOOt0bJNjn4ppkQ2HKOhx/CMYrH5ZtyFuuq1fd1FRchaJmPoFyf62l
+MuGc3GBhUqKd98WgyPMXoAtUp27coexf3/hTJk/vNsVzQrhGknGP/qdU3XzFf104I4CQ59VS309
g4Po8L55l5y/QK1r/q/0s3QFIQZQB7M2Xu4eaftxTRxTWSGOFrA9txDWT6fxu9e4G5QRgbEGX41w
XefgIkXSJlQ131RKGIE341pPNRGWK84n9/IX+YNSfNoQ+8zgbydM7sGZNO78VhVXmsF9PT1JVtAW
F7ij7h1qwJkzJj7ISOuEcj/op3kEBkTV5Z4F6O561wANaC59quwb9SVGKQeDzybZHAupKa+EuSNn
q44KL5jRJICX6hFmQPQ/cGv1JoxtX8oUaibjF2WNaZBlzYVvAyd1Y0Rd6YZdZK8eG9FLTumIVodt
v1id2fCmFpHXyE99/B+9XYIWJJuJnI+ogqj6YlqQVQeSLD4apcvoxfZW0+YoWdvkzTlUpKG6zzs5
GIkWrkTrPOQI/6nYSaF+tNCyh+klnzWj39oRzFDdrkMmWdkryZD4Jv5SKtXdPsujepG4SwPZ29Eh
1DET7xSSEcyvA/qDzmmumweJ0tDtJVdq1nfyua5u26zl+6PrxUqUeFgHSUIL+ZJkM1hcS6FM4C9h
Isau95LIcApgTm8K0NNGhYzW+Nn8zenVoLFspxZsvu8mrVLkECrRg+fjj7cdeViMKVMFunem+K1s
Wm5UbMA3VRiditmhlZR09iVdWvl3BNXvbHqEIfFvQddzJo7G9HrFCn3baHYYsW3DvORQ8xduMH3v
EBF13WxIUK4z9KXZ9i6WyjUHekCjXQu8QyrRpFvCeGBmHDqbUVI5k/fSO4Lm7TBH2U46T+dnws8f
q//K/glyF/0n4pSQKRlF7TMzHO/6InKPzM2CyrueD316OF1uLzeg5kaOffmFCsNJ8lRZ1EExNu8o
jfzYoi//whcryF02D7seASksmdyzqf7jGsDd1tJCIJ8HvC2CPc77Vk5ysfHQuOTlsyZ9R9hRYq7/
k77EcvK84tsmYN3NnGorCu2JjaFRh13y68ZTuiHs1EQHIBB/2Zu0U16YRwT5fDI+xBP+9OBdr3yC
bzgKygItFB2xsJB6n1aXVu0LTkrh0PrnOkwSrX5l6xYOEXASeZrBufepOqgH4pMAJAq7Wm3MjDQk
lsepEjx5hBg/XfWU06vcDc2nuX4DJPvljlbKTZzCT7rH3s9ddZbl8RgRn68dqRllW4fyrqOs0g81
kn6Ws63V0IYc30VvSRN0Eu7C2i+HtlJe2GZayIF/OGdchRQAFFEUrblHMtnr9zBdEtdYsv8aaAEu
d/8cjVvbfV8mNNzab+eJ4EMquFSlyBraqNIHMbDiFyqi954hAAymXveGGYcLZ7TpeAsJCQd9+sgy
PbXP4mUySzGSBdOAmyO+gyBrFQIGgYHbXJ1q6emMRGyixExrtE7aMiaWF+z6YNwRajVIe52a0ZeX
VrjJWSyrXL6lBr9Q4InsRw56mYJesCW1kMUf4hx2PLPGBwtNu5TT/w0RPZbBzjF0twrdk6DDivHp
n8Te97OqR9tQ2UErJQLZe8HhS7z8eb6HlZQV+qRwRMfn5NhJ8cbUgDXlZ3tAgZqIDQ4pgxblZw1g
m/LG/pc9FxDef/aNoHFJ9k3vtHM01WjYsA97lSGjuJU1gJFVKW9j9zX2waaL+5zwxLgPFJidlR84
D/njBiDpHtt1ASwKX/1g4jM7pFRkW6Im+cEtUO/5Hk0r84xcUUBS/OuKWqHtNUhMO3pW9ji2w1vL
7ktXrzX4wOgoenJ7GkKpY0oKQIqsQqNQh7fPVL+K+u0KK6wuIrMqPqkp8w3PUBekrUXCvE+sOqCw
i5CFfGF2k1cujp7ViBnEqTM0WXQySPnbt31G7BHKV+sP5MxWd0Xo/BLB9PXMqmVIqYoNRxxrDdLj
468R2GP27AeFcaPDgIRq1hYaurIGJeTR9bxQz+3VOsE5B5jYz3M7SH08cj/qFCQoxPjNVej3ALvH
aqlMWzTr2fgkWCdUmTJFQ+JO2XawarjwT536JMz9wytj+hxlduWKErnQy2vTx+OCUNxrrY4fa7ep
40ZdszcgIWhCkD4AHEidWfl05F95YuA7ia8ZAWV2KZh7tDzLqFeBnzfXLa/TydPLEwTIf9h7O0tF
3liAWuIlPBqdxA/smP1ZqsgNGVK5QXqp+Ule5AEctRxGFY+VFZ268RU2LaZcfwMM7XsLNikTF1AZ
GNR/5T/hgewHGRkEooaW48dJ9UR/LL2sJfGE8G/bnPxtCkLQDKHlT3e10+SO81xwdaQpEKAOP5Ri
Q8z7BU+GeqVb35puLR+9UWUzmcJOjXHFfSsqlT7WuQCygqSU7AVZuu2bE801LrONhkgwtl7KK7Gu
GaY4NrwXPhJb5EvkDBAyJeSSlkN3t4paJyF0ZVpLk72NR2mIWEbZ0zKXB2RySMOJkO8D+QQKS+g5
r7nFVnQhPsiWTphW14VCI3Z7kGLUbYUPoXt4jXujOsjUkZYSV5wxyCmO/Y3Zvb0KtAq9e49y/UVg
+boVX1+mfbvr/terrk3EO/Tr7nf4wPoaDN/OULD8pt3bRxG3HjoucErvtJ5OJi1xuQIlRk81OdpH
SyYQFFzlNczqTjbB9WUozkyATDZ59Ly/mAjywiCmE3ZgBnz1NmicmnNK8eYQ58I7hXjUKpakoyqE
CVeB4KVuH3fgUYb9kd5ZAVnsAKibMTgOh0d6qujariLCL1a1Mmm0HBWCVIDuNOPc1FBEdPiCS/9o
30/bVdzo6HugxrfguyhhZmQt9TXKBGtB4u9L3YmyYDRD/ruI0SSmIo9bX2LHe7uFDthZFsP/RKq4
etXumA1M1MCzv43tUI2UlChZX4EpIRp3UTF39VctKykwHzqO9ldu6k04TDU8UeatMyhQiSZ8bc2G
mmBwtzbxsAGhrUZ35+xfgZIwvJNCiyVU/2snhoQHr53MCgSHhEXFfHkQ29LzF8EFpoypRbU/F4qL
1DwUr3OptZJAwE+eHbn14LB8eK9VgIi3mi8t0mfSaKoILuXqxD4PsgI0LbJupP5vH2SmFdCfh0gt
wAVf/yNfVtizd4p2K+ICD3KM8a+JL83dB20l6zraBbBImrCNLZp0kFjXmDiWJjASBPFEu2I1129z
zKlcdsp7nVPyFPpNB1xWjrU2eMQqbSXbxIco7pBcq92BKiTwjpy0za2c9/Pvv9JYtIDaPpkfnDko
DKAW8HQp8MQgxjB56KLiVKU2RVqEkf4dGjt0Q0R8KKZyk3IPHhOkSgEmFlOjuBgTXi/FXXZJC+zd
67vt+wQLU1J6Fkx9U5CkUuY8NTTJOVNjXzkvwWrE8A+Yi3x6t4d8UCmlTzrhkYlVBlRVuKSLhDr+
X6vdueh0bL6QRaoSR2vcE/yaPV20xIS5nLGdxqRpnO9+5emsye5ohgzLyXgjGvM/vNZkRO1OssF/
jurRoI0nTqgAHbP+47IjjdYxUsp29Elk2ZEATS1fmG4cXwvRKxbvh4KxIfpui9Sd/uU7QkQkE0fI
amLV9SPCX/dIYETfrieJDaQ2CihulByePiFMHn5eWCbBbzq835qi+Fjy65RyNIkTo6E0+1HLT2xY
ptdRo1b0gRWWHAW8NJ8vHyZ2IM1MFL7dYiI/JSbC6r47uG6Jddh08Peb8EGbLL+sJQoOQ2CsYfVs
KvZMJQrzD3DVy/rx1N5jjopk7VxOvj+PmpqubyELZ+KBouyc433BhHflq52V78+x9KnyPRnQ0B/S
zghtDadrb0ZRNxBZl0wRWApzIMWfOgB7iQRNPD1IsHq/Ah7mLR7xe3lc7RkqA2U86IfxtQpEGJax
YU5d12Oyy+WVIHdv/LJ5yN1JJr5MTlHvwmOb+mmyvfV9a766ASDYL6CepYcpSEDJur5A2gkGlKWC
dBEukVg4pJaDcGZUEOr87nmwIIVx+/DGyozWZhgQYTepAa88Q2ebmwp4Ng0jAnAaRTmi4aruMh46
At4ac9MC/ASNGnoKP9zinTe8nlBPOlcF9hHvq2Gh4mN8uYKGWV6I2HDQMfygwb42Jnph/ICLj0rg
wEPRPM3pRjVfgQkjKJky2CBuS2kKZcG4JYwjzEIBkZXzBy5v3tl0Mwzhf/mQ9RVrlrwGXvn3SzCC
PDZzSln1PixBWpF8hYiVI5YJyhSzx4+KWXB+nKAa75LPJPIpfw+YcNxRxxJ26svTaGQb5qANVdHP
q9/TSkVKKmzrOcIm3IX3nGxpLmp5Cz32KmcPfVn7jW9PDBM7GAiNbYh65pcR/87TvvmXpUCOCAhj
243yvYRU/K9ueiPJRG5op6f4yOOEpH5dyXWHPGWSXVIVFiKL1+Zw2XqBkFNKARfeW/iFPdYj2NCu
mf1PYF+84AW8d9PZQyQv7/qk3S3b30Ly6YrHoEFKA6KIBInzTsPiaxWBrJNYI7WhydTpU+WvdTSP
fRnGlFQo5gyiFxDQvCIfRDw6cK94Tf/3ASis1reI1sh0fyP0srK3t0LotHM9emFcQzHiB9weoI0F
xnEREgyhBKkLjrGYhNy3Q8ki4dfhlf5GcKO+NlDLm8ELhJ9fDj22LjJdFf6p5a/LRgwyvkLgH4mu
WXjthJPWN/BqyYi8OPnybbKIYfNSHHwHfCp1jsusY0M8ei1lENBK9h27pA6MNxDampIRgTH+Uccq
5HvDqWWPHzUqWDxX1lC7x99ezNpllcnza9HL7KR8vE9/ChrPEQPLkQcgDoiCoqdfv6Yid4Jun5uh
nNj2hwS2ztrcuhiyqHYgBOxxuidMWpVJtVIMQ223v169sbLL2yZgg9ESDNJwGpb3B9l/OJeunEU9
RxMOTRHptP2kiiRFmVtsHOcFxwzVRFV786uRhC6h+UCEa3HH2SHU2e6rtH7kgSGvz3EpvzLmDiBw
UFoLlBZczv2peHt7kOf+leD0EQvMpja+vYGLH4CrF2f4oHE1iyoINzTwMmuaRwEXNDOdf1ThgfrZ
ni0Ckrjwzt+vEB1Wn2O4nmChdx9Uo4vifzDvxc9TL+zA/fY0+Owo7PuBiWE5vYKFcjk4SKpxqH0X
iJQl+Wo5xjHoN/s/1H9aGL/O3txJBFYdvk3QSnD6mFMP9C6QbsCoz0VE3r607Qp/XrwPoJangjdd
k9N47cONoIK3+MXEzXE0t+57DMhTSi1v6We3qKAkfr/aKYHEQKmFS3xlIi9gdJaGfL0QvmLwqqY0
S/1ZKXFLsMldU3sB0jumg/gE6IEu8OwQLGACeylZF0EWV8aM4NSwwu0gEI3ll9fpz3bqwGCyuWOC
aLbQ8yZ5eziO0cJF4Momg4+R+YXXHgYh6gjK/VVRd2WnwzBWqg5cazk2DyN+65QHMXCehKmUkQ7+
/yyERgCEVRETzYL9GLQeHBaC8M0Wvtiy92o7gX7GtNEzux1X0mTQnRiaM73QzWc547AOMslk2WMw
uWz2Gw8g8XHVAECbVm9vCHO7ejOGL6rLW5CNm/jt7MzZt/x5FH33q49PVlKaITGX80iFUmJRVpVj
Rc81pqEOtbOMssz9Tqs5krbjUxgLXxMzLwurbTzGdjILVFZ71CGsBv9v1gN7c7F1vzMzQQxY7eE7
QRoKlExJz/Wl1FXReRzeufjRfFyfJRb77on+mJ0Zp5wrwMmrxPy1NjW1xjNvtldIYHVzEA0+ISnt
Z5b9our1tKDsigToIcfK7jYczZ9IhSb5t2uMUvwfxk5EjHVWHg3XhYeA7yCTKm4379s7mbhaY5NS
c8oS70Wp+fWompQDVZqjcsHU0p+Gvc8bUp1+JELhZVuCBiio5s0li6uo2pbiernpFNQNFO+L5SAQ
vfUw1ETASBzp2NTSn+9v4OY7+gcr+y/XHxD3knYLJsWiAjzhFtz5hkuBXEIuPEIJGGD8Twc3V0wD
JdxyykMDMIYgePmV94BnzVvXUlhJ4otEdsjz5EnglXhIepkRx/NYzrNnYUHqlR/KP38gw2Z1wSTF
qlH78XIckQig4arTep2JcygduIW7kZVLMoP734+N8fP2udIMyjexW1y+VIBe/+GLbJzr9phJDVLc
LDbQuhWQ0kpS9MfKnv5pJGN64TMeD/6zU7g4LEUAvugYmWTRB94i616TY+SUggR8EYYfxjk/iadw
IwZO5MYYP0AynlrhJtd47ZM5yE2OySpJbsTT6Px6sxPqFy+YoRslUczlQ9Yl81GUgwk47BGAUO6e
VXOjnZYIYRUgbUizv/xnk2OuZfgA2QECwcKpIdMeRczJfTeBMD8Wo9TIkilc/R0qTJjNeP0F4giw
8IsCnYaKVk1pNEgW1CHDN/6S+nAkWOffgUbkNrQFbLSJkpLdPrn6hmXuIySKZ8VuYpkuo+4V7GaB
A/YCzQiqo5W0ERQj4AWfdSPEpMOvxEZ0v4lbdxll4HMWmP1vJ+Vs2jfaoWrP3qV+o3YnPE4/fiWa
APZMOV046QQGXAI85RsTZCB2dNtFlZCNDSqFaH63vgT5O0Pl6qjMf+vVnk0eTLQd6HSD8VvwHrr1
jPAdQutS4AXGoC67hRw5YZQHvjl3WzWd8itNYTfGnrh9pi6puyAvhWPEjtiEz6PWDZhSX+iiVT6E
YtGVWU1F/yF1N3x2JdcLAWbvhduf4pITHcbFctzsSZ1i7wFdThzaF/Wm7cEWHmukd9koQDrbw7I6
M1cbsrd6uAS8Gvm2WoStqaEILdn+kRJMUy33X5o7zGgkgi51Gv8pcS3LWC/eOSW/XDoRBJFs63Hi
FBBlwXYeeMh8BZLgh+QRHIeCG2b3upF/BO2tVBImQQy0Tg4h8/VunRznof9sD5okkVTuxI3NdpsK
1pin/o9fP+L/zvjaJCrekLfxrc05tmiILRbpuB3QIkTHQEQ1vG5a6b8eO4a6iTu9slGq2S7HrbnT
48hCw6y/qA2d/rx3ApYjTlD9YmZ4tQm9KO4+4o+4+BqycISAVF0UKlJ5GEKa9P+tMiQRHkbjw/BI
f76hx9M9Iehz1VoU0NdNnNKBUj/1pNSOYDQhV6g6SYaljC+69lrs7qGsdqeyX1r4kUws4i2zCLzU
GDGI7y9heV/gPaFYX0JJUwy52t8WSAlx9u6kcuUAqIGeyoNq8aFhZ2aWFy5beadKLn9RbjwfNuI/
GJn6mNMBStjLDsf62rtywqd9MF3w646ycOJMMUJtJWNunBjH8Z/yGFvpWSJLAS+jHjS3g3on1nfd
c6ZtaZOdGTRGovcnc+T53Vo5aeT1S7ATpEwtOX0ZebI+/PM9e0K4FtnodF6IqPYA3ja8IsoeHDph
tbNnBAkGsYchit09jj0gQFFB3fLpmqppqKZ9doKPdge6lmXtfprn+yKdlaxOkzlXj/cI26tlkoYS
S29NAxI0YBuU4kuMFGUXq7rGvYJqxvO9f3mCBuHGdC53/QQAhqAf90Gblsoz5/wmjiAsoU+L2HfL
WzCBQy0lusmoeo8I4O9yecfkPbgkyZArN11VoH1EMR+dCpz1Z9kkX4n0wV/+WRPt9qoRuMtcNUqc
BjH71eUpgbBXOvvGNRJEIGXAWe7cDx+tV7hzIiQC4AuWO736PHx7xa97VhZ27D4yWqnv66LEHiiv
lWaDa59xR3RBclXSgzLWDRVZqFjL9m8J9DQdDfHUbUs1AKYZeS2fzvfMxV1iQtaHzCaWQJsEVJwM
mYDbjL3hDp/3+Y3NgDfIC4r5SpNxeKki49m7iFN3kJCXHzSoxMxvnotjCTkQU/nX1Bm6e9AQvivy
deDCTVGfCI6iWZi54OKXgFAKYF4UXgHYWKO2r9ZP9mcp0wJk/F046yhZAxkHsOXkPd0PyHhl18z4
wEIDu6fYFZIamehrrvuO6tK15VgXe4HYuHHZ/13ahSRQEQ/0SF3zfhYQYI7Oc1U7ML5lbIkgG31m
DFXjGH78yVjVFRkV9L7nlO6q4UJgeJrkdpFknF4MYYHNiLz3c9dIwnaaGWfJw1jMxhanr7F7nFNf
c/mCyAEF8Y4YVU3foe3jiSx41wzL8CcwqJeRcVBXB2mH3ycqjEXVOW7TH8TLPfKb5w1l9hhoL7e7
SF6NNSL/TSnSWEPQe8hBCQ1Rud42DvMr+W7eng4arCJoq9UlqmT6oNYTO9eutrP8qz59N1GQBnKd
BxPO7v8MveQUjh/voLnNpmbJVX5jsWoJ3zgfg82lVI+AkD4QAoKLTa6b82TIvpSyu+PQ7guexi6r
uMGcWt8t3CuSPH2czR5RrzXun3Cyvaig85O6ypedsNB39v9v2oixJSw6udKZvdZh4T+4H0F9tGKh
uazvOcT+8SpsVoc9Gs7+jx04qpOMEmGbWZTzLZ2mC2ef+jenOWisw0BZiigU4+Kx8WHBmun0zC/2
Wx6C3nWjT117eCaXyT50HUQQIdG9HHmHpJ6qepfj0jpwFqaVYe4LWZdB8YEbJftzCT1ihGonqjci
tFyrTBrGNk2j+qiaF0duCZjiT9NAM5anv8MRomhmgJYFjTUcdRKvDGFTSsyly40h7qw5XzyXSdiO
GEDIwXtxqqIJ9D6ImAZqPIrM8kxx+I2I6OzUwQH7zyAYA7tCD4kRswowrRn0S2fe3D1kFqhMGyLg
/1tsnCIwW30IXUsWthwBWUnLnQy2zJVPQRIEhbQiSPpJYWJbQ3MiUNrEAkw7VITkOMuGvJ3JuGKC
9dcPth5mLezCASXVHnSo5ogifmSRunUU+2qa2fMt/s5927x0DGKpEl+75qVZZl4n66GBj29Aw1Q6
hq6k+f9jhoJeE0xFYgTw/OTClozZmgkMwG1ZqQM33yAEcvQZKwmvPpCYxgvhzaylDOTUG2H1xSyD
ekhoF3wmVZJ9Sht/0/8UQQWcqAmPyuwh2ZnWyR4vHjBDuFQBh05zJGvH7aq4APmAV9JP+Bss4TMD
4wfG5AyMrhw2bQhVv51yNEcg3BfENzmBLqvG5S+498knwbvK0oPdZxtqnEFj1D2yBZQtLhfGqI+o
+TDTZWHtjZ6Bo/Eow14++Q5yR3qGjinBtEGKBb4WK5ak3HFn9xSqagWwZGu6rrX1gq6EkqxfiqXy
pMamXW1mZn5mNRZjI6b8gB0074afW4ad5+B5/TqM8nYcRnRNwFMyJDVQk28OyLXDduLBAosAmYdv
qPVH0NgjUMpgTE0C2hG76KziYdFp2RAsFUhVQ/GClO0lU2ga1m0QRc1IJeky6TrDuHixAZoBW6b5
Y3/p31n7kFTZkYnNL+9W/WYgjueVVjr+jr1dSF+mxqGuIsTaYjcXOCocQiMfSJ1V16ECtpOmIMWE
WrYzuhHz5NdxxlmTOSWq7QDE6ezAKb8ydLyHo+vHnoJaOpK0YTS73et5hLpLkYhsOprmXwYATvBu
1wbFToQ1SktgHmcUwGOZzHRt4akyHTFa6dwOcUY3iWlpafcaWHoW2j7WEV6ma2uqUAJgxtxL1iBq
VqV0P4RgMWx9gvspnQSbXr7pOHZWN/Wi0KHEOMG4pW7TbeOr9DrGj5bHyk6yH611bcSe8Paqmh4h
w3NEwfoVSj3Gb9pn9HN78YTvFDhyewEqEmdQrUsnrj1mKm8XqXLorsI9aRyNTV5PAQ7E9QhY4HQj
UYsWV0e0mSNd/C09NWCbtFXhDN4u8B8pu3Q5AxIdimorYjjx0g+dodvRREPK5be3zB8baUYgrC4x
WtDz4Qy4uHKBtcWf/l68pSHu0oUFKo2z7ngHZLzG6IcwzQrcR4O6NEltgcSv6M0FVHVMi/izQPRw
qjmdtYbhRnKmsHs4Io5gloOzouEDaWgodY5K3tgzfgGKSvtdnTyLJPGWPF1mo9SImmeyNZcT6LLg
EbEiXLTEF/OIvr7NP841aQYYOYLBnV7qfEiP7EBgR5d6NwS4taK4xmJTANDEJyYwqw6XWlYkxAOd
ctmttxj/8CyCOLtURMvGAZIv9xYhp3NskkbXl8Epn/9G7x+YjvM9c1zOhEhonQWLYxbCDGvw2Hkw
9gfOHZIpxbiw0M7ck5Hjbmlp1tP3gvO/rrmCzCv1uvrP5lVyWTWzC2ywJTXxSSOOk/KCfVD6rQR1
AvSuVlDJX0PMIBSfa/LSlDkhXTQmWzX69BM6FX2+YS30wbpvVPRwbnfSCTs0bMofw89oIJBvfkIR
F4kK5VmfyvLfWvTM/TPBddGmvR9HthKAzz3u8shHFgY0BzfeExWrJLKJp1cytVhkVCveVH1gqZJV
HsZa1kQJWkAKUsPdm9FPk4A+DEzEApP1uanbK3a/1YZyTPpqeW1zgJE1pEj2ayo7WbgCb9ZhNcAF
18XXfsrXqYBjo6RIJstg3Xhj2T+9yYyiExmmHpR5ZimPcR1yNjqQNDFzp4zLHfeLNOaYlVqJJ+la
8s38uN/FaPWCHiTVlXw/F/CFdPxWdKmhFLFdEdhhA0ykAkAvtdfJ7wSO6+0K+VeCreY9BacmoLMI
V0JwwkIx1LzZ7b/6vCEHjVooBSmMM+d1Yk3/R7Xn9/BpI/DeCmlmOB/ysehCZduNimnvG/rlPxqZ
up8d5PQV1av/EyWFLpN6Mhl6gczLv2+LK7lm0M6skzkWDXuqErKz3KxWstqr9E6HQImVrz/KLFh6
2qCijdlyJpjvLl5kJQuec6ZBpxfDoraPm4ec+fhE9lMKklxDZO2iD8t3iogVyHN+TyH0Vbaa5Kb7
yrauXr1h/8VezcrqsQjIbKdc9mMG/unbOOzkl23Axnm6Si5O+GqFUreI+jP07cZSYG4kUNI7GIv/
RQJDRxAml7r9cT1KgpSmgr1Q2rnrNhAk8L6HWJCIR4jGFg4h6O4OkMJr+qoXwA1cLumf7oun6N+R
AgzPV8tXyhgbawa1X8VOhZancy+5eTQrAdqYdp6hhwf/FSFEcKEfwcK6xjbBA/ZwbedvmMnrhwTg
+OXwLNazeNQXugKfCYOuK7BbuhGLd6RjOKhmwePMeQAcZwXvJBmgyOi4dFo2vDqGmlJcwALwohFA
SxYLJfimNmEQOIWs+lOLEvixqfcGyfQKfyoKZgEfSMM47103WAdX/YW/szYptuG5AjUen35gyRrA
9zvVyskBdlgetsU6ZWfpDsvJUw24E5myxOfAP66wMA+L/rO3xWiIVa0p2BLSpLYocla1dmctlFoz
9mmwT4I7rFz7Ha/y8VDGQJVjS1W5bXWXmUYWonOHczbrN3y8qem7T/IYMfgwkhM9aCWlYirGJCZE
mA7xlqMX8HPoiWoJLr9mTcGpFOmegu2MTBvHrUe41q0g5mI5Vnn0ItyPuFr/kbjaZPw5lYGSYrCk
qdggxk2SnnEEeWIg5PzIUnnRSAW48Fa9KrXuTRcq2/dnkwDCg7wDT1v2cZ7HYYnR8siVGoRJSZh7
HB9ZuFz3Y8V5KfuC13Rr7//TX++x+jzmopBfBzEPEDOd22PD5ciBGuRIMUFUF/fpX8iq6N+kVSnb
2uydd6f1QaZabbPuMya0E6wH6NQ+dNoz+aGkUUScQWcs5aEbZornHSgMlzgPSp5VI6+efPsssuDu
ZuyOPCunps97+EsYQVuRIAuLlQO0eOe4Fo+0FqT7o6ir7iUfOJC812qfxvCS/kM+3GKFrYv7OUfC
kAFpZPxmGtOjieM1LZxB1DRYiLhEhUYgKuNVs12RCl6O06K6CWLj5cIaU1AjgYoE3uIK2MS/K+9q
V1q8gMk8BAXh54ZfIVIBd4W41OBZfNKRqBM5VYfyv4FQ7yVqYJzYCIjr5fwYiX/Yxy01ijA7eqs0
+Qo+h36Ojt2wGjlGInvw6JB8JhzACwspplwZzqPostltfZQOIuZEqoMCwkZc21b6jPtH6jDcf1EI
f3EC1A5I+ym3OAR7OUspdDEVH083SJLF2P3cqKu3u+07gHbBV9ZGSiPJx5sTBpa2nhmgmbMp+Tit
7Y6E0y8K8+5NefgcGnn6tKad/HX+nV+fzHAlV0uMBpRDxa0MM6blv/cf5+3UHmOIdHhtge31FyEa
mXMNVpKTR/jJlEfUJDlI31pqYwnunpjnYEK74yeyAXcdE2YxCVuyWypMtZ3auZZFM3xw4RlIUBmH
Zlezu5hhGxcGaG75HEdxsoMIGldtM3jAqTfVN8QvTJ9srcFhe+hyPse6LivuoUxXUdsYLSMoOwvR
FGq+qzOgj8xICHUTnK1Zt19uYxzmePbRPl/gPEI+148FVy2MArEnbgamCyRRZkFOuBl+QSiBD3gZ
4nteccHsgwknLp3K45Sc0Kqj75rZNmfUK/YkbqateBcTqdvSO7hSuawSuIjm5wJ5y5S50tl4RA3S
IsiMY4yat3V1kbf73IzuXGU4NKtRnHXH6d3fzczOCy6ZMdJFMFsz8my/DKvrECua+p9wd/lD9aG1
KxhIv4T+TXO6LilIR/fOgAsvKomL7HwQ/7c7krOrTH4J/HkKVT8pzZCOrt6Vqe1kbOwrxO8YKrGQ
DZS+akjEBN5peiZjodu/pyQmf8TVhWPVdlaQWSempi9UUi/XvHb5Sv7fbLKQK1yrTCtxIIPNm9It
ZpArtw42nPfEv87N75rpz/4TSVBQCwoHICMQuYMHgzv8QmyDr6LitNOkEh7YmfuqR0P9igri7HN9
kli+IIcAKVOF64a1rCGSubjH4bzlXwfziWmw7N1ULU4xTi2WpXtqJdkFfdgJvZSCIVV2nO7Q5iZJ
tdyDjb85W+LoDO0vtX6DP7AXOcMGRoOWFFErPZ8Iwv07oan6RecDI5pAWAAAAwgLtiWcZT4VeI82
L7+BhJPJcYPB1fxcZ/zCrx3V/pFrGXHhqf41/GHzBAWzk/7RvBSr820ke+IzXcStHf8p6EHmJP8C
tKPQg5lKEggV++dYqApOitRmg3EMTrgeTSre9l+Qy+jC9OUukS7M1t3NbB+6T78vTwCYN+LXR2Sv
52hP6WRVmwIDwdEOkVAi294nhpK16IfjliteJYkFYqgBKve/LrtGiGkfQEX9c19arfUehADsOeh+
fJTC1PTlgWhf2fLosysFI+7FkYLPRpqTA+RQ26C+8YNsoC1QtwAWMGlRHYB7bTzM1BBshvOxYK7q
AorJbvzE3jAxlRrIMBR7rtDSoqrCN3US1CztDkxDxRUkkeeuMHWUPX14N7p/MaCeiag435nbAv8e
vnIUz5ZV0otu8csmIvItFheI8RhruncRLnPPbKRDQd2kEIoaDQyO5f/aZuM1dOOpC7EvqQ5Foou5
cnapy3qnYllqQIV/44VqxAeD8BVU32+VEjZq3KE80OQSrMEwdkwb5Ivu3A47ABrNQ3Wxhns3w4Hv
u/bbocJZ8UKdTaP9ALWL2mJ9y8Ml7Ml3AkghJT/m19NbcS9DjD2PeEMPJgKJb9YIs70xKKQSA6N2
FfTgtUQZ6HZqtw/5XSwi7ot8Epf/OvEfRFh8C5EcrhU4bgpoHPnQqt/EI9vC+BMaYXHLTU1I7o3+
k2MLG3QgMBjhv0IswZgKkjyBZae3naNi3Oq7DoonkL3C9UHIPl1IFyEjAUTpBluF+fLvuom9a0Ds
GCxMd8aPGG3QFJPm9Q9+CnP7NSet0mdQ7D5IB+jKa32kUI3e/CwP0SQiY1y7bi0YoeIIP69Kr49V
RKSnvlMO2gSald5T3b66rllodrGSFbbKr/eMuQiPVZFYbxgmJsnhx8mSVzU2g1/qVC3reCOZYruI
L5S7WCTgSRPKtVZIcHoX0Tt7BCG4FvqJB4GNZCpxAkAMfD8sawkAob5HYQ7KLpB7CTHKGcQy45jc
otNjFdgTG0euoPxzz6zAqd1CnD9yd3kLCE5wQFF8uONKXdj/s7d1oa6VbHDa2Jks+TG2VOVBD201
9iy5fOARxuNX5fdyZC+jJ3WtcPpM+5VJpiiD2WoL04XyR5CDgvJqwmLjWzZi4+JfM/uVBD4XIQ31
XGDU+OmystJWMm3UDlTYf5AgMcTP7zAqdIbdLtod6kUAf9WJSGhEIqANS+XpAHuB6do+k6OoF49f
jqn2/fAvi+rlryLXWTJkDxNumRlJgKT5PtvGB6EVKHt3lWlZczZddRJxQZCjvureA+/yzVcJGZZK
CgxPnri95AVlMdH/nTnzf7MknlByFESbqsjhib0ahRHqMKbomXVgaSZ33KvKzSFWDjwDtXWKP7al
QAAfyZVoj7IYbL/+XFiGK60h+oMSNKU8sc6bc+6OBInmUHsp2n7F94hcQ7p14qMiMXuIz1aMy5j0
ONIY+rQYEEVGj8IKQYikJ57YFHswZ+XGTsVO/ClABHvj2K8rwsJrYS3tH3ghbSO9Wu6qa6EOVm19
5Mj/zm4/oEsy1ZUZq7+YjplGFtGfs3j/T6zGWMWw9NkJMyG2AMWHi1c04tBZNmk9qp6rDjdUGeA0
1ozj0OaSP5IM/dR2H6goNr3lx3ON3BYAtIFgdP+K9xtaLnGEPRmHdPhymHc8zz+9vBvlfnvrJ9jz
VEi75yfW4QTOMS9DcSspHDoC3Aq4ieOMl5oVLV2C9mVOEhd6cJRUuZnACEwp+DhELRJc/tiI706W
5Bo6YOc9Pri7JRi+ahTwyERQPt5oQoigmVTDV0i7MG1g45pi8E0w1Des3XxYajQt0dpRL/pYQSjB
3uDFGRryHTHr4+A8W5G28RDuI+WzOenTs24hBq33s1vpmxIbLe1Cilm6IuGpVzI6NIcpqTHnsDW8
xSkAczONxKcY6Y9yq0JmYlWo5GAykYq3xo8cxzUs59IlzCFH+L8GMUZOKQeMpOzLH2PyImnfCXek
RanTQYgLTS+i3g1klBefxthQK2iO9q2sukkP9cXWi/uN02inturIOuyZZ2FrFwVRfRHx4K2VLMx5
60C6MrxFsDy6jJlLbiyEHwJKlCcoml4khdQRH7Tp9696d9MzO27RM84MB6yBEUUnFheEdxnYEIKB
4ZNR3CADJTHiUonNnPMuGNhll90UhuFXe+hmIoc0yjrQzCZ/wpyzpsoUchje7UMRg2GBmqC6NKUe
3g/DngfehkgJfS6vAVTj3XrJj8z3MsSJgvB94Rlcy01+RqqmOLhKUJi9k7BqDjEGwn66yziwIeSM
lxoP7zQAIYJTLYh2gy3rZd1NU155vYI+IteU+h9OArWpn4iLVPWvUgNNPu02ozAojcBZNjQYwoPU
XDD7tn+BhHVwrIBD5l7XENp4v1guQ3l9jKJeWwh8BokFWfAyg1TivPq7gJ1BVEGpZ7RNxEkrQU3k
cfGyl3w/WTqtT625An0z0zD2YI/zt4wRHKkZrUtvLqFJC7Jrms4uIwHi66nmIhHfVc751ZeM5zm0
n64Jg/K+l4tPvokdpf+gQu3v5f9eQQcqq4Ld4wvQ2n3nsKlvzKLS3zH7VLNBO8wgkXgIi++UxZs+
QWKIqJY+9kvpE2rC+SvXx1YCAKYUOMTu2vBXZUiYKVkrvBPDOQNXComYUpCWUs7r8M+/4WkQqqLj
pjKHczmbx/O4/+epvYAif4JvuYYL9YtlIh7U+rjqtJFcAs4XDymyVh/VIXD+fPjaiWFKNMMs1+Qk
R8hAncQzlP3SQXNAhGXWq71ewKRLqqt9z6zhqRMgQbyWOJZOQ1JEULdUrCvipXgBTiOwsMaK188Q
F8INApQos2LEgXDO/FNtJPXUYRHKM+qO2Io4P5aDQO1L5qqJYqNCvtPSCr/VEzqkXSHhh/MARogZ
R/kEour33u7cXDzI8tMJfLuBJQDyQd7XJJuirkFBxMH08H0o5zw841ZsraWT+oa36a/nLbi7vZ7a
P0WGTum1oeyf1UvXyRC/VhAHLpS0wtT/ryz6Kc6uerGWtU5QRdpEoQvCT6kbuTMiIrCPoPd1/SxQ
/ekHoDDFY2Dnxvy3SjHZu/4xRku8RKhXgQHn3GuRMHUbAYXhR7V4MjHVAYL2UI4c6eiXbGcij3qG
1+lmP0kH1Lvk//UdangpShIGFgwp7yyyc5/MtfX49iVvF0mrSoNlNiaRmBb8ooR+oMQatH7d0e02
4j1MK6jeVfvRZXDxhGHkJgBlHRX9JbOb7zzbMqDergOhxZAKA4PWG1cOYaIFrsuDvTUPNKkbtss3
9zPcmkayrsl1XPj0nICwmOItuhU243ch+OgpzCe58FOR/WAFJ67MrXNaTYEfhGfYQWQu22qsaiwI
aHDo2sm2JLKmVAIho88M8aqur0AMVIjCekTw+es9cbTe591KvdzL0YehcdarY8kWoDeV8VYIfQUp
ymjzI5E3eukJrXc6NBuhQ7TMDENm+5Gy5EA2xNfyghxcoxRaqxO0pfU9FtfRSLWAAobZILCwvKrb
Vq8f+4ukqfC31SaaGlQuSvMvdfccHPqv8eN9QhtWSY21L20HdLzARv1OKvg5SbQADQaNMXpNxgvN
++f/SydM0yjhF4c2MgnE2voWE95q2CV4YctH0Lx+13hNGG/JCeK5GHC6TSeaFm5fbyej6z6isf9B
sL+hc6z/CIu+MKcmnUCLJIyeg6RW6iThdoSA25F9mbEbWVEDhTUOt6LmHExRTmxaLm7sBLi9oIVY
8SKNht2LpjLsYgi5g9jTK603qRu7JPhjMN83KW/UtKeRnVKTMSbd6CXAaQEWkFDsetQ8FBXvHmSM
CTsSeD8hTTz0qDtirFj3dvICawYi6Gv6SnE5o0Ia5z/aM/N4MrD0shN8lcyNZPVRuSbDj8jv/Ioe
v2Y0Ik4XWnHIxZrQCjEwUita3tz9UwyJ12Dz4O6rJHggMcVm2c1zL6BqZNd+uI6ud6CzfhbzLKOS
DXbC2or514vjTG6Up9WQSJAkuRf3kUQt0IL76v7ii4BeqZ3V0F7PCnfKoEsczMbwW7mm6u8wqCjX
y63MVvhDamvEmqR1cZ3ZwhHK1VKtrYx1mvAyZ1nqXJnH9pGV+l2dNk58a+Q7Bj37qipVgFnS7Jud
LgLFH+d4BF7PsXnowRND21k1ivcruYoJklDG+dBFwBryfbsGnvrW02uXvx9bn9HHBAqF4UGm3nrT
2mCLvhoVMX/lHWOup/g5cL7tM4Bc07rcaBh623N8tp2ddE1TKa8Qte3OHnXgEH5U9nGCURcUijSt
mHKzhTk39Scn8J+zj0+NfVzpeRHVtR1BKXhR3pTlMsDAxZlH9ti/o6Wz9GgQ+vBBEH56kveEqFq+
F3CtzekIUHbpPzgg4/cxAw4t0P9plj7T0xK4QGuUahQyKbPX3qgezN62JYYY2DgKdxLbMR9QxYqT
c5oK4bfnyRVUHCGMmK7RhGv9KJBdiTXwuVyi952c9sJhodUWu99ka05vv68bwPWE/+DKzN3BWIm4
vPwrQ+0CeouEmyx+8lhAgqH/rGbjymRgax03PWGWoyqvE/BSM4dCa6p+DjQIOaurNAlQDUV5ftP7
EG4PHvJNWnHoZpjRzDla1vUz3fnk4hKUFkrbnML+jEbzqCBjeQF23zRKPd79gDFzw5MKOngf8ima
AgkHM0z5XAL0BhIi8q9fQlaA+dKLv0Y5d3PTU6SFn1Kr7coH5ixeanJS1hmrSw7nEs+9EDiDpOjc
E5kQEVjS96a4j25ZYkM6fYR6Q+m1L3t13dvt3Z2Uq2OYEGS5cZwCHKprFe4V0RyClVhveEBncsJp
J/CT5PdBNQ9llt4WjthqnjtiUAXH96faxa0iWuU+Ul25gqrEBiEb6w24BSd7eM+/Aqgx5VTN97ZJ
oecRbMfXguTYPqiLd6VBu5hppsgMGVMvft81nudoXth554RHZB6SK4kMAFx5ivYh3SosEMjECbP6
9vIYtq47tuibrTEaMFvpynjeG4N8PeN+c3HxzaiGXvO0btYGRqlgkQPKyhpRNPUinV2epJXKWCiU
tHnbPkGSCh/Tn05RkOqHteqLWPax7RorlcpQXKtGwGTh88HkY0GZiuppFnBE333l2AzZyR0+MjEO
IUOC0q9DQbYO6vtDKCoD75V6z4YvJNrLyChgtdh48114JAMQdSnyh8bkpw3uCQ9ogP5Rnl54x+jt
xHCXxl2GeUOmN925cmAW/0c2ZOmDQ+j9jLsEw7OhLORXd94m0MGQgHYJA6WXuhYNETz5cUX6Dg+x
9YFyafnTZ3H0DaP0P7bw1dZyMCC+hmQfkuXkWV6HQhy6GySGawN0BQs0/Qqr+FvtiDbulemL+sPJ
WfauGFnN3PWXq8OVqHJVb4WUdmb+na8NW7B3NJPWUFA/JWjQvWX7VpWjl9y1MaE2Hn+P44H7weD2
cwknQlPn8mtwPzC20BPpYusIuK1UJCXGCDzqMxexyq/Yh3hNIXlLOkIjjIYv9E2T4CIavGK+4chA
O4FuYynPRYwd5ro8qL50Z/NdFJo6f0e5DkzpssiA+irt7oURvGBJrY3UHz3AvzteF1bzGXFQxdUG
CK2hdWd/8qJVjuKRBWAlUJv2wkUZpidnYbK8DjMXJa2X3l/XAvZYYomBJ4+sLAyF4XzDnRgJy2yP
vfswCoej5NdntqzhgIs1GTFeATVSN1rqzJZYAYNsRhYZt+e10xd+6kWKfE8k7NgQ5Glb/WKbjZO2
K5E9/9QGQ0pFBVrwliRkRYBV2j4307LpR30VVjY/2WOai3nQIVwgALTgq0L9cia1rYUEz5QO5mn6
TuRiMJY5CrwmF48/o7spx0k00sUBLpwUZ9IWvXDJ8XKTCOqELJx7yMVIVbZQV8aZoaTQVqzrrPce
2NV8uYxlkRiQ3tv4wzXIuxXqY65QNLDQlxzwP0giqdDWdDWrJOmsPGoNBEv9Gk4bTFr5llW0y0RH
yvMbV7VqsKYGbkfMxY1d9tnhtP3kuhuhyj4OBZYZYAtr/xxaB1bwIRKn4AUAZeG5vBtlUvxjA7Z9
PaA81KNvyh3XJb6q8/9JZ0/1GTySBMfMBC2IDk/OT3KNDk8Ej5GjBoFoRMNLDowwHfh81xbQSSBQ
b/RA2kPZ7KAFJfvm9MT7NgFvdFPQR8HmzqXB7oB+h5nxgRsLg6CyAZYpWxrkIoVdOS6FA/YhtnlD
LH5SfOU/qDg6cL1xWUCD+Mp4EasAZX82jtzDBfuYzrKiDtTeShOK7sFABh+5LMQ1paIZYyIcA5S8
1bkiBwDHnG7EQ4JpGSS4wCUcwzPI9sgPdK5FgG7CRmasai/JFKM9Sh8+xraNxyhFSXgOi0htYXPr
P2P7JJP/PH6NF7TP1wpyZ+DHoHQuG2LYQ11TUH8+AB1vA6nk79s4O3BSoAqt/YpfTT+5BoTC2mD8
sLtILDr5jEnWKmV5p35bpFNuMyVTZF2x8GMl+mTfM4xip35OH0+k70ZS8xx5R6Ks9lyyRrUR3FIB
Z7h7hFEY9YDLTB+tuEEtzo/ryIRen2/jvDi66VKVYag/P8W1nWBCHXLDQIxmGJbcIYvnXkZCY4m0
DCOMFx73/Wb7sGZwfu2UAcsPIVfRxqXVzbv0HAKzNdHiRNGTDSXxfXG9hb8ECTIXjhFsAEKRJ1BW
q3ACUKRyhxdVT4DcDrJqe6psOvkCnpFiDtruWZgeruKGoEJ+XksZirEkFE0lZVgM1GyuVGgaO06g
4RD4In6D7jap5/mcc6Z1MzIZJWE9MmtbIOVuIo3qOz68d7Tt5DAI6RE34sFrrZKFtcsG06/4vK+7
TItsOytaQxxFLEPrbjJVHLVHLLLWV7WmaT2edRFqbVSPNc2p6JjHQUNOsCcpCEPtwRw3kDF6bFtq
nfNQiE50GZyXFYTunTWUS/AfyvOT59fh/n4zPrq6PQ1Quqvpk6rJwgvsEmwM+gUd8NtYleX4YZrz
nyj1v7MZFsjqSb6vid+5Ci2aLNMxtJUymC9aMG5Zyo9P+K+oppoXiget/ZjZQ7dKN4cwbVtPXN+T
WL73CCtwuRf1NlFx+kGMMamI4Um2sCkHvU9QsizwKiIPpLlPwcMw1MIJHRxmYh5tCJD9L7IbgI+W
uihRJy/CJT4l2lAhP8mUsYkjEpwWzBco3n2ClJXIBSSP7352kEI8JO2yVgPMq3d+r1a11LZFRUMs
3pLWVafZoOby+PpjOyeYEpcVSlI+eUfNvpKfCdk0c3es6HS27SiQYmpwTbOpVpuW0AQDSAYUCsto
jUbKxvuTuWbYuKzLwUKdOXhMIp4Q+JHxtk0g6ZrSRugLXPmaG3raQYcNs9Ztq5QsZmcBdseePxNF
zCXXnChT6S/44yFz8KZwAH4HHBU4XfAa7FTCZUMQsVdHqD0tKxf2XuciiPUXFNRvb7rq79kW/rc9
AyoyPZcR8tr8+h3G3l1I7C2+mH05EdvHM67LyNbUFWKFNDE+efXKV79RwfSEmUHQOzJmqm6QQImO
tsb/n9SK2PBxPVA0eW2tir9IjzVR+QoiwJX0KSVLD/VOdgUm5FJKqr6ewX3xEC2xpxxg4T8SMEBc
MUBqpuKoMAe/jwvOYno/IZRiep2vNsk2+ryH4XtOhu3ISvkzVxTYI0gWyaf1awS6mzv4kolgvukd
reRVyOsoT3ghlfONps/z5Q5Sf5Pztq5W+COlb0L2agheRlzRZkGI94+fMaFpgDIJXPH4tTTwjOj/
by8wfKVZgUV7eZWHEbpmmZDrTQI3I9Mg6XP2zaYsrWFrUOp3c0pJfD50/aYfpjZn+b+z8O+bUAuX
65R3pD41Ed0BZS+w9ybvr4ctac3sExFMzl4JpqsDCsp4jbcdXlLBhTjMLkzalOhZ2Fewk/vPElfU
E/92tCfvG/y1agCIIO2y9RRaZSbQ80ymicPM17HtTzjd9fP6gwxT4E3YpKsriwB+8mQGBPDGh5+0
fu4TwqS0kDbADIWbcaGeK1Vgl3n57Ilh7/6+Of3iMZyz0TUDupo07b83wqBLzhcYfKxtH7IDlPPt
0fjY8ws642B1R3zCqMp6wSee8hanFEjXMESwnWkBMO6F2VTi+tm3s467OJMKOmu0MGFg6QcYUqIW
ldOq48FXhG9TOIWonktB3h0efWvVzq24PzQj1brMwbN3IVgD9p7I1z+b+jNF3659BHdWtRL0Gewl
kzgc3SzyDGMKlRXWjoTK9MUfbsJ1cDzst+iv72RD8t+xqy7L+gVwr9vzlj5YLcy6GHkjUs/rB8T5
h0ltbfXV1LIBXaB7x9EFejUpXm9P/FAklJDfzVyeO/J0JADUSSPOkkIt44wnevuuJrEg9V67jQId
sRN+2XXYAoNWxbZWFgV2IQUnez+ntL5oBa5vmRb/NekZvrQaLyeOgmHMrg0E78NXBiOBQx5qgQr6
AM/PTleAAmaiFbmNtAfEvfru+cvzt4H50h8ETrueG1t3I3O+ljk4UHsCRMaKo1EA+0dODIfNkfpS
RxsVK9jydqD4B5zeCCWdwPwvyYfnyy7h0yMbfdIwZeHkNXivJpwkeFPeE/nnK6jLhiDZFtX4jDO/
L3CRwR6SaMfDAgJtNvzdmUOFWIoET/Uh/HH3afRXpPRhLB/QZQv+SWO3z5vFBhaOH5aHvi4KvwOP
QlbVETSg1/Ojl4H8qvj00LIJx2i3bYavRyG9hs3kIbpMzIr+cRcm7OR1nClYAqU3XW5CtTAqRJp7
LYNnmJ4Ih0zFvfA+hITrreLI3+ahXh5cBKdRYbt/UFaAoZUOJPBcyJhHDOdr+pJsAGqogvhtEeUs
gmjeyW6ra2xXZRZAHhseviSEYm9zrq4HyaFFvDR/B7iA+z4LIwQld+HhlQ3i8S8980dJa7BGQNe8
Iwya/RT5SrlwuR782ddGJ5cIGqG8lf+zNMDH3MulFblSHKmVVeo9V4miDbBQfnBdR7b/JQhjBSu/
SCQiCvaeAGwEJ43P3knehSnq1jDy/N/sNf/w8jq/M53JRithaA8wIWX4lINuViX7C1+/CVtZpAtG
98u0fvTKxIfBehfn+XdGgzLZTzGZorBsvKZBBqgWoBdVAKM0/cFK3S9a7QuZlxujbEKnvEORCu2n
ePVg6mhmOqScNQn4prbDDDGQmklfJZmWVrKyY0beannYLrGjA1c56o8tAuOnsLgkOfRrViGTnFnW
lmFe0g7wjsvk1ej4+Eg9kaQxBYfu8LpkdSiWlZWTjiNI3oGIF9ybuy8C5NhpVijB1IFm6LYFTOZ9
xFUorBmtOQTK758nO2PoiNTJXNjZQDUHZ5pKwoMyFj9Ko3uowbSDWj6f2MRpHzbZGMYEdYtV2P2N
Ixejp4eAuI7Qvq54FF4AhupReuDMWbCBxPIv1B0GpmG+4dP3JMLggvkcF9QPAuK+/TBz66YxbZGW
du+rha89X/RZXh2jvBEcxqAW1tIKxdGxiG0uRELiqypwmcQiEtmbNlHKqzpG3rgYEQflfeydYFEE
JhZqekMpOnoaPWr9u/J5waXHHkT5ljySLO1kOLRyrSQuQz+S8bbBq36WY3FpS86LoGDG7qBmEugh
rKpm/M3EVsdx/orMbezVAC78T+KSMSWk4Owuyeor5CQM/XFf5XSGaX/h5MKhT4YQcXBwoukbCzcR
aGgE4SzpAK29bSxBxcj2WlTEO9QrpKmOF+m1h8IDI6s1l2wqwZiwIlVep72lDbPnXLxyk+lea5ZY
q/cZErlVg9GEguTJxG4HdXVTWvBnhX/KmcT1qtz51CVq/FMIi7xjLyAJ1k5n1Jx0w+9HRu1sZt1H
PXr48p2PUr16U5uYahp64BqVdlIxJ3lojOC+hc5kCJWp0QnqOdeXDHd/+Wg7ctPBNUy+v2MCurtM
jbEFOXZ49aCr2289j3UPSW5Uqsf5/KqV9QE51W3bJul4jKF4NgztqELkbncdMTAot1k9QV33ynkA
iIb/hzNwl8SEwKh1Dc2peu6j3ZBCP1GEpxHNq1xvfQrgUqjfsQTjZuufh/PfygwUBiRHNVhZpoaW
FVMLdSS5uBEB8nxFO3rLERAevGF+FwlZbfwDtgivKm2Uasfdb/5NLFpfW+cFXLKtrj1Hx9qm0oOv
dWF+M1y/c1S2UQ9ciWbPM0d9oimyZEyp1BtNT6YIG/odzuSqBSyg02D8qB8z5r7s02Jb+AB4gRzx
Z5iT2mSVUGFlAhP9gruNiSicBYzTV/xsDWIoVS0N+Col8Rpqj+ZtRxXWDHOQyTp8A+QchtT5tPKm
TovOWzhn7tugFRImQlR9aG0jyTBeb0cCrLc/FIknZ7tIt1IvkotTev9M3ze/Y/VsKAGHf9PvmZxB
SrenKrHIuNuWk4pSS/raLcCk616tu1ifb+/cZmXK/zbTvKALP9cMzbJI1blibwHJkuPEYrWuvhTZ
8x3Fq03ruhvOD7C72VqayILtfS3Oi3gI2J1k1kufJqG1i15TjU9/iIw2hZ48ys54aiR5PnrtwzJ9
U9fRSBphdwhqG2C1UttPG6tGpABeBZU0yqbsDIHWt8yRQL/BkDuZ/yTmdaRKjD1itZAEe1vJXhLk
1s6ZkF7JZuSII32ZaU7BUzQGxcvglU+ObKpY+BYK4xejssXGjTr71vEPZEhS6TaGPUDXIbs2wduN
aU0OM8cZ0J+tgyTcir2bfbKu3o4nY0qLR8RnSVawxnLzefwVn1isT4c1iTuOW6rt0Q6J95kSj4mP
61Oo6dQeAEMwiy6PU6LJ7Po3ror1hjxJGFZyUkqsdrV0L5BANV9N8w7d1SXLMtUY+KLtPhips4CR
14rRguP0HTdwkcsGeDmHdRPL7c3H3Nqko3sdDhLbf2sQwnrBOfeKFNR7YQlV18yfFrex3bj8EI3R
fwA+PyB2mm9cCsKBQjBIRLE4T9p6NpSwPI0MzlY7Ne5vmVOGg/LGA9V0x+LUMtgt+Ca904cMlw/3
c8+RPqpUrK7ZOnq4BUQJD2H/fb8r+lc54GN6BvJGIkCefmmfaivlj+F/Jezqnx8jnX0F82A/uRq+
2knKES08FIEsBP8UPgLQBf3qrFd8PMNHlzb776byjbKjSc+6U/ELaeZUwn84L2tQGa5XhF7xq+Tk
ZfsBlha1B6xnSwlRXCyFuoUYDFwa6mQ7mtaVkpmP/aAIOYQ4OCOPpy9qQ/pFyiCRsoBtVZRC8E/b
wnRANsPf/unnbMzuSN5ch0cdAeSqsqgBDW0DYRDM2JwSr+fbAnOALlF6zUwYEe1hUxGbpk/IwHLt
LOXbIfKWPFBkiWYeHEFS1oENxrVSuNq7EtQN/ZCa5XsH1KLUrUOgAjuMne7Cyxum53BgjHy538j2
dD/1IPamotaVBDKrz6RanV8XFgKMHBf8sQRlwVoGyXRzgm0A9um1Ok+79MAJJaSsEQhruTlVmmnh
GIpsH7KEr6m5aveq877hyW7cPUpCjR9K4KvEBsFpgD47xpfNaanodxIWRQik+1jyWCSGSw/ZDpiT
6g+O45qC5g0IHj/mZIG2UquY+WpMRyD0YPjCL01J+n31Ll0A/2dWc9ChqW6WNdLIKDtKaosjpHV3
z2b2xrG1xy1XIRDp3qGN0H+t0OW9BYFMHfZqqIWudGWIiRCPKAIvhrGpZx616GBksFhZIGEG61nm
jH0y6cMUMVTv3MuUDyAZmhfaerFJEBeNoQWMjCRXaPJKB/0zCr7UbAuzzByjD7YlYeUy2jjV681M
xx7yXfXht0vSZ5EHCiiek/BvfcmbR0uxrEw41W7OPHiHYYqxzidWUQBWqplbc8SYhiMn0k1/cyPD
ZQ4KYsW/hpo4cZilU9CXT8pm8xYGLo+TrRz+jpUQcj28L9fJ7GdlYREKELX8l+fHs5GynTGZBZEX
1n04kISWAFRbnLmhgjYheTlPw2dy2GnDXaS/Y1H9pgKdMvTJTEwIQ6bf4usKxuluVuc6kU2KPoFk
pbwcdIJJ7gqCrJoSN9GjtCe+mqlJMLeEjBgXXENR4RmU5pdOmuKAz+oCp5arprzT12Fnr0tMqxTd
XpIrJeiCADwn6SKj/gG2Ucxk1I/ANHI/VNuAfiLedRJ5/UabKkSUlOXpVx4MZ4ZowWpXTDKhgH3H
qQDELWgM1EOuubNOMaX3I0q1EFMWhB5ojIDdFWrQLLq8vCck1Yz9O75t3+kZL5p2dG3qiv78DsTi
zaWWLkoQIzyYy6Z7Of7ZbMSBIzjSF1BrEU3W4ck3WePX6h6KTSv1y5uD7yeJotxj6PLID7PsQsZx
Ed2ZqrPC668xRNKEgIOIy3VnJAxsjc9r9J27Zx9SwIp8x5XMgmzNHaTrDpwNZ1ynxwAvq41F2gwe
gcEGjj0vdu8z1ZR86F0MItWCl/hT13d7DbOPDB66nkSJZjGNTSw4nrr9edkRVcdwhGUqrVXMxPxp
oHpCa1ZniXo0btOJJkz80SU1Pb9z6dezgzUi3fsVksPX6uIH7VzFDMjR4ose0izWpESbhaiFzzf2
7ckTphQWIQdMSLoOVZamuJE4vEfrupfuBDWP2DLcblVTPHrQKjqQSb6PBqP891/qYyzpNy2Fc+I/
CuceZXiSBCv6xP/kixj70BgKynhzCeimvYpLMO3mwH7GVupSBSErImtDp0CaWaCgBzgdqr4bZK0h
EhSsbNrTIBKl33uUC6nwhfx7t0oc/R6Bvw9piHMJDkoDFs8y6ZhFidhhyEf9X+MJejSwyWqrdiHL
vhx3Oizx04qm+uF6UIXXtg5czbWw8E5ZZf71hvkjumsHVv8SPyjNFea++8oQvUch6mWJYR7L7jJn
vSJQYEfdctN0ttYrBKjb9Ub9ORueETcBv5eR4ITcjYXMRimpGXBddHMFNl9Iyyilu0xzVc4lmrjb
2RTR6a6jj/cproDsUTEI3w6+A95nJmyodsjWELfsQCRlQ6n8zAJ2T/bl4I4R65iaJ5oT7xLNv0T9
oos81Bt1U7LAebSQxgub6lOC/9j4Jdldyk4CMUzCAz+e3l2gioSSyfmEivAr50Opqvvz20ou6Nlp
F1Wzo4E0a554uUUMmBgpJSyq82iI5dEyl0GR7KgoxVpG6sHjBrwgtjhDS1bNYzAceNYeWPHLNpH5
kum3/Kh1Ew1lgeOfEEmasBm4XwyxYDlshN0g7zEOBdT5xeIzQClo4ffR8hI7Y5e4nPGsdDQS29Dm
y8DC2ln45w2pk+lb+fyjIuQTEK92eJms5Oq9JcazYm69/Z2FTt23JekO1auOhDfVVruJCS/cvEXP
EihrgFyEgq1wuuyrxHHZfNQq/bH+xhbI8NhET9wXGr4g4F/TPXFFHwwauKqnmO9/I1zAj2VGiQmV
GVwq1Rc7wytyNBrHyuFbKwqNrFTmwvTQ7m7vssLSmJDvCnRLambQNiVqTtIWQneZov8FAiUJMUEv
bBKMtYUuJQgmBBJU6R95NZmuKJAVS69vj2WjNrzVDZr5xItso6n7fp8IKZNZenCUvUt+xhIGY52M
bnoecV0nid24/h8uVERNvEUZ62iqM0T6ObInvXuR8iGNe+zfwt//tZ4BmKcradL2ZhKYVWjdroAO
SnOufJ+iwMs7L1BYwitLuOENyR8XEYAi75OXlYayfLrGWB8L/hlMayLftDQDFwgi0GLizkpb/Sxu
0TnL8sIWZrfRb5kk8n0HboHn0ynizXZC027E7aP4pVpk4egrcz2j4+/xHt1K5CrsC8eBsp69nJxp
YVojy/+qZzh2uwSdXzd/SvhEr6VgjlpDjfACnG7FlAxHX1AQVGTf0F7+LNnJr1H4M2Gm+dam5qVX
prU6vIzIKBAHcKP+8/wrZoq54JfH4lrGZys9IHBpbjoGnZFeNsyP+/MraNgzBOIQ4Hfv2pLt0BvL
T/dUIO1wa675qhBkjm5m0pisnLJEHi8TEvnj8nB2DHMARVSRzEt2F3KvIf2bqWBYzA+5jnDzdFPs
I9JDnzhj55PdEv0k0I/4z/otOGq2NtOkqNtcZ/TD7sYd/3/69PohZSFRk5RWA2TNz+nwFZITyYwl
uGRcqcdnHsf6LWwN3Z7tnhwvhINd1pnvtKRhUdGNglIFzm6LvjFYbkGLMTnNU0emCu+kcXAbmueJ
qugl9OQPPvqqDetWpOHrWNEFpI2GQPXfJOkmqMTaRl1SWyMAW6hiYxiMfVJWMkVEoZsckXzg2RbF
z7OqOkGFDNhIBMb5VbxZodiymSguMwLiTm+mZLSUSJRVusooh0e+pAW4Jl4dUgZYMUQGb8vdRzgd
SB8ifE7cBrX2cTug61lX8WxuRZluRKESqISi8Ksq1Hl9lMQk6n+xLmtkUT8oUTpa3RejpoGYZXzn
+oNDn4Wy1J+UFh155bzcxEub33te9X0ooHvRLy8f6AYHQw05pfvIulnixEwbNfx/2lXTADFXFUw/
JBF7RBwA3yArTi9HUFjCCWxn8kqKIKzgimBf/WWylSgOmLlq2SteOkUXMAcPiW5CaJzdlWAFMgzp
huuQ+RGYeffeljgR+qRZ+jtAtROXOkYTWeFN8Fl0csvC5jnzXLqS45NqM6uH63EhJilm4wHgGjKJ
b5mAIVKtxCg8BOUM2mtANkY6FH/mfAk6nejxmmokCVAjyYpEOfGIT2yRrpjOF/vbCd95cD30LJn9
unbJd0lFmCQFgadsCOQ9TjBU8m+AJDLllhSFzNcPDf4QMmYTSFtMUPlh7yIIgh5q+ChYgf4eiwEt
dp/2WULavgyDKGYqeLPo8IQW3Ma+6Xan8SDd2OmW5XxOuOouyeatsgpVOErQof5XkaF96lLQoQxj
eqynR/TzCX9pFTpiKPr91Ex8eUABnM2ElTcBFiQl775D9CK6ZgzyNHsGwOVKV1W/WbZOZCJ3FcEl
nzjfpjqTcXeoaFwplaXHRUomQP/2ljR0GYaGo8WPD+m3fVAbkeL2UIAgsokbLIleiHQ6m2faCe7J
5eDNiUP/6OkodXC0k1bXFhzPMmtUCkW+eaEUXwDE0ZnLloqZ2eDdBI3etK17j/2GpVvXj22TCXJM
qVS69Gw473NV/z4xnk4kB+ZBxAFXpy0co/qRchkvryk+OCt3I7qDnvd6TRcjgGwCiBPt0LYnyyQy
goeyvuxAEzm3BBHYx28MCL14MiweX2C3fYMPvr1BMwhPv3uAsbTQYpAGujHbMfjsC4vRgs6vJ0EY
G0NjqSfR4IiYOAaLIwtduBGZFurf3QrBeTEW1aK/MqouCvyDSLIfhIqrrRjiTHTjrQCKSlshH5A+
3FYMwUYRuNZ9MQ5AuVK5dJzM5Jgy85ay3h7J6FKSMGfGeTutu80upVmwU+n0BOZGtPfypctT+Kbs
cLxXA8uo1oV0+ai6jiIpn64rXzNaVjrOOw4rVAqScofTd9JV1p8Txp8ThOQhA7qJRsjxaa6zwSxR
5acUUuh72rzdd4mn6wE8etWD5jMiAdT3tHU89ifRVTtMHFzV/8q3Zhz4x7bMlwXwjFhFgyCnnTuf
ztWfJv24Uu1IgY66VRLzgagMwlHiPWWF52JUCIZhEUHk8WnAsqlpU2fmJH+W2u5PZFtp4wGnOAx7
OLwsltlSWni7CY0awkiFoNYc8HSTxZv6ZOwmdDX4XEfo0Y7Kt8dodffz199CtW8x9CT5a+xVdnaB
o9SGUPrE1jf7Tw1AZD8ZKqh2Z4fgbH1XQSU5sLMTyU9gUyfxicWLlVE4sLSuvwIP4TL6jBNEJJ07
OQ6+2jHn+pbBJNU4A+w1Ul6g9fRSoi8/zNEqEPm4Dy8hhAXCKXgHYMSV/mfsFMoojlY2Mi63b4h9
8RDLAmNS965LqQ1AEAk6vazk36GCL+DtzX0XKh2TQzOMEt4A2g3L37IDAwle1Tq1/Vq/UpElY+eh
PyKhBTYEQGgNE5HcJsYeRCEkyXPm9lUVUFJtfnPgIi6iQPAoFPoMARQ9nFhRLcw4COu27jeqiTt1
oU+RyHFy67TSKAChTnHbq2sG5N/ONQPdjWt+rQwc7kYT2VrdY7hLtTdqot/samK2EBJL1ld+5fht
XxdFF4PLGCIZMBn12hZuHk2ftBsPlyf9PyeDvyDGXqwcE+9NSMrYgD3szha5YGCD0Qmales+oxfz
Pu5kcQ8rIbDw4RGUA6O89K5RatUZRtoN/l9UsavY+Uh34faKmC0RhdF3HXWvAVuEqcoaC1ArgQKI
GHubwiNprydRfyor8tW3mQDU6dItRnl10dkKp/CxxoMfAZQrxMmZqhpAg50fDnCDXU21cEr0bSbu
eGAzmTifmV89ssAYrsBHZWnn7thqoKNc037Scs8MAv0+5q88vPBBqyg07xY4RCLWtOU1A4mWaMrT
Zeai/ZcKv1pw9DFRMeptb6Oqi43f7wZjjPqJdSAmjDAGmyqgCUDgLj9QQdc9LQi1l1YaMsdE8FoL
7Xki1IOeTjiRJJpD6XSezCfYC1hhpx8eAVEuPVsJD8eYrpHXofrbsa2Zdp0ze9/Xu4WsBkoCYxAF
LZmj7LYPOGhCvnKwfbFu7foQOy7MFh5YgFFsN5w4yG+RDSJk6dOZz/j/WMFDlmGtvwlJbIqhErps
o3mNtT1K115KJFVO4/IZYpM4e2wD5KY1KVOSrJWejAKnn4CW/YzKEzVkN7tL6T1tZHssdFGooJzb
gJY6KkyYazRNcIufm73dSaSR14YN7kW0KCmtTuhMuU3XUp9ovQLsZwoZYJdXxh3QERGbp2Vap9J0
aJBu2chXjT7zwD0/aEkEzezmRgoJQ32fQ5Kxqa1Zpzog/zVyBIzq593K9Jmb4hmh3udLrxiZBNI9
S4hZiTw9cRAo1meZ1sukY1GesGLKX14D0RTMfafyHXKzdxvtB7iyQpHSul8zjl8LeqA/O3YoHAU6
yIM6nNM8/H/vYBPAwt9Rk1AjZhG3nZLu7yRH7jUVn94aV38bM1Cc8I3OcNFo0207/bSoKU8MoqeC
mrUlHgYLbFwNPv/zqRkofjEltOo45dMH3ZWfiSUbvh3BQo5/sAkSw11TIUvAqKQCWnN7UiXV01PF
mY0Z/F/vw5W7sx7uOCb9xV1kneUtTq5nluILz0u8LenWoo+ba3+cyYt+chJ9Fwqo3MiLQyh5rx78
aP3M3qNowLXBdlFLgi/USkuF4JbirGgdrH1eEjqAPutran+6RXssmyP6vOE5Vy0InetNoSmQYMHv
FItZcxODUS/Ss4wNKDIzl6Bjt1XtJLrowGb0r1zqa6OWl68Tg/P6kPehyi5p1xpumG35GRJgTyLv
ea+A9uexqZzYGoqV4Qy/tjw296VGkBeVGV7LwmLR7BvV1vofCDTD8/we0SGtF1y9M+v3weL90B5b
Ezl/uza9SsOzNTfEkPS3QfK0z27SP+VJqTFKKSNnanuhs31pcq6wY2q45aNdbpXKHwUCbQm1YyCq
IIKwipQcmVedIMuMcellwF1fHgmYZhqmncykRr8PRsCyBf9Mqk6rxZmGFEFPk/xp1YRapLlJFkbe
1UJBITg/YzKkDes2xkdPLPq1CLNukkCD9kIg+aRUciL6VKeHzaKhHzfeeuPb45Lf+bSy41XzqdRk
bBCUqtxZJjmfxDAybfvD5f7w8PXWaV/8XvbbPg7VvmiPaXdjPt9IyD6bZUQIRVfwR3RLbv6x2Ah8
thBohccPXUgY3lrR/W1MeDPPkE1nIkBpcEkrQhUXTV6I/IrGRrngzD9iMSWzZAtZDlmBk8bGGADZ
qI2nDTdVLP/GfDQXwfwJBrsz4kwOMxD1Odq73/yDggla000pAuCI+YouPfclpmsqWYQ4fRyQrm8Q
0RRGD5v7qqABQJqwA67hKn2lvt9zf1R/RJXAGT4jtGTHB8d2sPCAwcfhcTiBjoIZWZmi+ZFs1ozd
U0XmF3h68pZw8Rp+ZyzcEKGdyTTSJabB+cktAoX0y0JWPH22BoGCTEHEHg6HtuFVk7SL00c99nPs
5cs2LMBBWVJnN40X6JO2QgkTxAx4UHaiZ/lXCoaBzkcRukdNQ4IIByEjO7oBslNBD3ZnpIHOUIhe
j4CBAQ3hyNTFmhX8oiPt4Ne6VQl+Xo6kXle8U+W4bKDqGZpTll8BZbsTk4u373eoayWtwFCA5RVK
8L07VZ6OZRoBmPEKtOg8bSsB9fA+nxBxJfsCN1lXRmtyRbRK5jki4J8YuRHuXJ9G2Ip7NDAbMPJf
s7j9Lt00msb6R2rsXOuQx0vJOQGtcLcPvEeg0q/R/cVwFGmZrEUEsdC68WdOFsjHOVcrYUsn/LbF
CUMOSiNVzIiJAO76akcGzCorKatEkd5NC3wH4STCNDYu3Rb7ikyBxCoXkYakM1EDoBRM5yWDa3nx
l7QScXc9ZvrVHQfGKvIIWFB5iU2Naci4AqQyNzB+rCX2omNsYl1wjZ5FA93JGTATwmnR5/Dzs9LR
eIW+S+LzgNAeRdbsd+QTC1Qu3oFX9MEtAFau7J0aOc9gM2L9Y+PLBcpv9z9FDJdTQVj61pf1dd3p
fT4QLWUVyBYdLMWr7TO7O6AIC+L5Dp/Ezgcvsay8huE34YcJRMXCUEbjUyJU9zwWY7XiUQjij8jh
olXTLFjrU2DyWYsenZR3zQZJ0PLaQfQ5Pkr0JFApozKRflquxtcGbDPB7oF6rAvV+BklJhToc8yK
MBO8+SNrohJjM6raoYN89GYzBrJTr7S2JdqwQhdHQM+u9NmH+Foox7mCuhQHBoCDL81OKxCleox7
cYWR9Uey1sCliCw5V4pwyT2r+aQjLRdDxh4XtFy++wif6znStsfpsdiuT2WArwfdgn2V78bOQ0oW
YuVV6Nb1K8p/6cSsnUNHGaNl9x2j7WOcdhzIXT1AFw4FtkElACQVK0ztWn24dx5DrLBOsP+cHsOk
2q81cAzauquVcGNXlqVFAHaa8NJCrG6mJO66t4uQDJSNDH1Z8CWH5laXEtvOn0JSQo4/EhSLGlJj
WKcBUN21yzKiq9bOpLYJ0gonCOC/8oco0wDAAxofLC25E51HWWdvpFzxVOdCCeq8xCp4F0DLah82
6ZOI1uHBoj6ez8Z4uEJ1LgswhagwUvMAfP+VRzc4uxg50G8IVTSZ1W5ujQeLTfSF6DUyxdV5rKal
qXWWb9SyfVLzwq2dQsLA6hYbjQNmtnBZ5BtqzN5HzdHGe+Rtq3Zhgmo92AXwYnhsF6IvYQrn7U3U
wL59fajfGQ7rBL3dhRde5rZYTW5zCaN2DU/tw80NeR+6W7G1F4L0AQjYttIIDBNAO9QbGq8TCj+o
u0tJw2DqtVwo8kNDRE+pAt9/jgUtYr+ZDMkjG/bob2XyfgiiLx4YAmlWVQ9rM20TGoLtalXvJ5/z
V2EDKTzwq+h47sqN9qbqiiYkbxUIZPlpOH4vkH7LuFb6/7d3KKxKZh7//2/uLix14GWRI9ZQg+9i
MT/U0yRMxg01wlr70TWKFchwqHm6eesoylIq58XqiwOuO5TE5VaSGzZeMu6mqB9DDz9zEgjpikiE
AUARlT9U0ZbqcNze8goOLB4iOdZy4jUn32NYu7caCoTriemf9kAsyfzhtR+6SVkJYB2lKqwTEzj4
jPZG/d3IW3vvnMUcEqzzDn5QLyKR/eTWatNWFRcdsRyVV2L0817U2FuIQFk9rZ0kHczzZvktd7ar
94cxkG1A8saUk6sL7yRT0xth/SZakNNN0iVrA92kCPFP29cY8O1CIQdCXRrWdEcl2QfKPGQZwwaK
c3fSts4DDEKyyGDgEFrNIN/8ZlukrH+y/OmrED9t6czEHhU2N2WLMEkXabdEa4XGg6HqUiE0lvMd
7An5hw3pkCLhFii9jkUbV+zL3gOa7z10ZzzidS7aQ32LskV9Q3UZXe1GBmCxsfudF8w9V5Tu/g3w
ShToICcVKbkDpCChGn3a2pZ4vHeSGyDXlLlKMn5qTzBT3NV44+YoID9Orebv6vg8B6mp8WxWe4wZ
v4IxVUafDKk+v7ib88eq9CWH6jLsDNZpYpsVGmSlXg1n3tZ+eFOkjGUXEIUcEAWfsdyrrMMdP0/I
CBQg+AKbqOvqCEl09Yk1qse6itMacV3t9TrT/LVEd+1AWuQHtRvmefziUyzNAYo54VoVe1zZCReY
ME4FaO3Jzpkoh6y1Kf1Fkioevq6PwYKu6XEh5zIuBVOu3FXSIYpnoBdpgFu3EMyUqvn8ItGZtv9k
aWV6MIDXql6U+Xtz+UdQWE5V+fzIEZvz7UaVapbQXgPJwWNIuT6Pa/Ql6XBGKQqT98Ln6rZnDJi2
aLtYG9NiRXv2W+ap7pQ5P63Zy7cLxBEKVdYjyS03iWoLa2LEnhc9bgn95EfbQhcxY+xny/bAprBK
xEnXEkcA43ZxMNmUHTsvDzoGkzRofUwJGor7kNukcDnuRze3j7k+Cdh35EaQa8I/cfMe5jHP11tW
fUPrzo9Sm1tHrSt2WBt0Jqzz0FIK8yEW5Fjvd5+zA1oj2r/KqCe9QYATyk/X7+T0EETrqjbKwAhp
aac9LUpAdREdjsYZCpA8x2uS1XgsniAkAniEBw8ccFuZpe3OHLtau4M/rNgUrfHUeYIILkljMnQ6
aDyHVcIS2reMg2AoVJRYo4BB43z6lR4qdrBqH8BSaO7bUx2kwYbd5Pp4/Rq9+LL+o9+lyzLwJR8v
vReacOfi2shjiRdfcCoeGMu9DKhEJfpePD/QrLR3FRsL0dLjqlTEFOp+h4UgQcIVcQWV1noUhPlJ
3opqa1Od6oVsvN4gYHCMVQOV0pkUlWVkw7K/XTxYqVWK+nj3fxT1/WXfe3JOUwmrEz5DgGzqAAGJ
30dVazEJeuy1Dd8mNml1H5QqT3tO+JYJBdxWnf0S3D1S5P0vhYKWo7qILP52VaHlQ6AWwo0EuNnL
94V/oF/M55TZR2K/Of+aXSPskmgUUBgxugwlJtFunhMdQ/fvb3Y95M5TJ99JPpfqRpLFzsE8zhvW
a9EWh+OLfNQS9faskvG2BRuBe+jbEOAP6OtcZHIiteq4xV4UYkiUjaejO2xr/4tg5lcGunsLnk4r
eewVCzvHQZpcYWmRET1cuvnQO/jAeiGiKHnlm1bJrp9vGVQb6XA7cT+QynT79OeZGQ+wEtycjQr5
YJXQjkgP7GuEi1sUyJF+hCQ4hHDRpYbAp5S1jotKr2HZeBHAgjaajVyOEJ7Wl2mCaZ5QbKEcpBJ6
C53r+vjo7cVfs1L09mHLVsL5r15qSiipe0Mf70S7oFOGDpnQlA0iGlge7z84UXS2Qojjot9TF2/Z
g8EYQDYNpkRbL6JQkRtYwXGsaOPQxKiz/wLwiT38TN4WmMH+EmBL4CRHcUvtPJ73mPOJW/pPvw5t
qKOKY5GV8PBEtqoApn/5h5aUDmTdPLiIvkHDSBnPr/n5WSPELI1vYtDeb8B9nWKsxBDFzsyaUzqW
wnoXBrVUm45v/o78MjzlQjQ6rqoPFQ98DUJytmACnQgTbgS0Gv5AMpJ8kPeMwiJnXu39z/UUSY61
w4ArvkJVDGjCgjoEheQdq9erh54XGshfOvIWvmjU2JE2v/xleWsIll9LXt4u3MByqCbm6HCCh7dK
AUT0pB8VxL8Vq92up6QTLTLUX9TlM/4JI5wsLJS7yHWpgj4/Xc7q90sVkH/yMCW7wO08C6Px4G8o
AOojwXImiXd/WuCN8iPu3+VrYKEKZndfWzhTv/nDFSrlTbBFwLOX63txrMqEZdB6ppJ1UVYZ2pHA
QCmI/WjTmMfj/JKkcjVd2cs4TL1nniUSnvDkVkh6vEnDCP8G/3a3kPP2frc/NqMJfI/eWkUIlkdL
Nt2Frz5Zq4Rx807FTRoOe/NPCv06RUE/k9JZZN99pf/4sV+3zqxwydBrHw2/DrgRvppQXqrbh6L4
uK0GlxjMh8ELissWX68vcuR8KgnWyu7d8oKzcWOpGvVXIGQXu6IE+wjNz0qv6qt480IVNcxc5xma
71eRYRGLZ98bUXByHZGsjD81u2N1Yf/KY6p7sjhnVpdIcw1MXPQYlqe+OyfT9OOxee3i3U6zPytn
dDdT3Do23soqeCzr5voRv/RQyk4QGUJk+t/NM5e3m6b3iFuLXiLj+XGle3SEwv3ovgz0BYZosUpw
is+clZbp19r6nPtpTOtSdzilGAxsPDr2S85A10uf3P7MDsBPYlVxtsqD8eEe4o214pDnb4ApPzcP
Th8zW4AAOIF8t/VSuyobkRLVjscIn7QlEJhQ1s3p+etLVUiLPYI3Xe9/YBU6kzn43xqMKAsTFwGC
d98nvZQN8dsH/c9t1RU7USCZRagZFbz4+pyaUHXzk2mGixbDKvNtd8oJc4IqJ7cSqmnXL3qPrVVA
1W2TUbS1xqqZxDg4sVlVpi2jSwLQb/NmNpY6xudwQRrOlvtSopmBCiLfoHkDtU3s6KJXf57uV58I
ni1DW/2U26hKHYqlLcT4noFMcn/jRS00iKZvLbs5TZssDhxhL3/HNCgNsesgfN2kJ+3ygr+AMi59
nbDGXjy4RP1hnTSBb7RBIHMg/J4gN134Yy2ud+vdG/RwUIticpRIBe4pHGAnc4xZEd8umCTmMprT
1QMcFDK1TmoTEtj0CpydUuj8DKCvQmuseGUNmy2WJZs7kV0Gaisf+4PN7Av4qLiSP5ECpKH50mxp
ce33/sgKihGdptYePpYYQKqCgHw1xoXnGbOEphLFG7w7piJJ20dANTeRLRaga7AT7QczwPyQFoJn
7N3xhMYv+ayvnVWRwcGW0N99Zkd8iBI3JIMix6cRw0gOEXybQILyPT56NapNTIJOdzCoUX33tF1e
1ZhsPRddPAdIUsTpn/JHpSRJN+R6RZaJwBhO9QXfzWDDjbzOwlyaKdrG/C+4PXxDBAIQBav4CA2A
LSQAM74OtxDbYLITQTjhzJJi0MqL3mc/0JSSIO2Rk7bEqVajCGx0RWwkBQzFnMyCkoLVyq6jS7y6
NDK2B9dqFr348Y8Z3nL8zdFo5Ymy524oKhdfA80/eiIRjPRwJEzuwQA8AflBMrt07qMmLyQHOHp8
vd8AuYNGGHKjzYGuGV1hL9FxEIUerT+1OjN139+QmkJ5o3gngHqcljYnPqqIpxc3qGWTFAvDVZjd
DuerJ6VkabHivJ8iT1jl3ynguoLeMpyTawkdehllqs3159BmbFeqvMz1MvY5JK5gQXeXBDUbuUnd
rcsgK0dWjFo9h9SGujS7nXppuOaW1SxD6a+QY2ed4WcVah5lquVCkHUQy5H0Emwkfw6P4JXXiYIf
P3HXvmksS948alU+kRGWtN9tg/mtdb/xTItDqpIbGGJT+o/vUbiryg5yRaoCaE9uPZuYC8Xbf8gN
SdUKVZ6dX0mpFCxZc+9/8Rkkq35lGKwcbdOhl3e+sW7Q9sCsvA5FHrKyLT4tZ2IbmU+7F60z+g85
6+RwUpCQjyPy626zhQPMfd9N2xTb28nVXZn1+28KHgEe+g8XKfCWT+lfCYQc9MGzMj5TcpEYz5f2
cIS9v50iYsbeq0v34LbVWT1zsHrVWBHGf1v0mQIAKpbTb3kvYcJK5bWnJkz65narylj9uopZnVR2
fNH7k0PV9OJWTMYLIwTyqtfm8vrp+gKWceHuMecYZKIESUALotzHU6w6K6THg87+wCTOLO0INoxr
XLNmpQZ7iQI72okBKOQkEsSTC9Aafh6i2RF6SRJV+1Wtb5Gzx8BHoGnAUWDFzCRbtCfm9B5MOcnY
LQFWXM0YVytKZWs92DIXwPYBcWRyn9Ynje6dqjB14T+RoZpTdQ8Ac2Z4uOVtIO3HajiSJg8yuKcQ
Uws8MX1oPGz+hPVcG6TZI79qo8+h8+zUqVayfLI493KaMelQACd96UONVfm0AwL/YWyi2MbQ2Ihb
JAhTr9D1CHwFaaY7IVyEJz5/vCpOcv6b0Hvv7P4njfOgrtkjYJTuUpnXZjKg+NUiS319gsoOgf6E
b6KpPEaMfw78OoOvLnFfSQ1dNJj/F/bGNMEeD7IoRXD6RUpcoPlIXs3un3PGisDYwFHMbC9e65BV
yueOBW4Rpha2u2rb+v7U0zZnjul0U/JQnPOu6Fr6Eb3X8T86Foddoxh6CFVeYJUoXPFX4jKxvtk4
Wt8nNBfsZyxee2bHDcbA0HEtWn4QRF66HcDYFKWsyOOmNFDypKEIwlGOcAzonXl3bdHgpQdA8bES
SmeoH0cSDuaFMhdJNX9pHxPpUwT9IZ5zssZBnEuOpCtYv7Iwbq4z3KzIXo9V2pl+hDeZRez9euJS
KnvQClvcp5s0tLCl+zxPGacAN1we4Ett1zDiWJebJXTL3TqSCYbqdExERWwUCzcBoNP7piU6dGM0
YlEqJLN0s3ePuHr1o1n0AlSB391YacjbYnWz0EQtGIuTFyAlprSq7693gsjf3xhuZmq3R0+txGX5
1oedyEomewjJPZbyoJcqz6ZaABbqxyKpx/2hypb8d0goYVheBQoyKn2G7Zv/j/HhJquFlowIJKgs
BNRZwfZ3bYAPOFLQAMWfUO7apvxeg6iwRutJrMiTx/anTUSXCL5bIox3e4cnXCu5Y8HSwlF3cKnW
eVIxmeIoEz8Jw1es0dZpGB4Ab1HjBvmapnSVyRtk3n6L8jSBpCkuEj6QQ/GZNZhcuYISZMg5KAAd
86ldY3V1D5p6h4XnNjL16r+fPbLGpozYwwkPvbHdQxDoQ+5hKg3WwzngBnCRC2CtSKGC4DpiODiJ
IkObVovfwy70NW8bn48OTJ4Ecx7JInKt4DXN5SwA/2cQF3fEM8pKkX4WKBNhOq5cWenjmJNLOzTT
P6h+14csw/GGWMUtpUjM8bZERkxcGvTdl2alpHaMQ2lRaRMJpnfYiuJTg+o7qpckVw5U+RjlXQAo
yn2ZzZ2EO/0HyqUwfhEqkwh4uWQCtAqSRAyYZhstaKvEZf+jXcGqk1VYXVpkR/F6BoMWRU0lvD0s
RtE0Tv7KmBdodiy0Nq51sw08JfvZ3XzcSJDDb0iKn2xT2LGHvDOQyEER3q75BVyLO6mXJDD8aQfC
DJ7FOL9mieN3Gr8oM1qCNU8sT3mypGVAkKwiUvjX0orrWG2CCKtrLeRZ09uYvcre+Fxeu5sCLC/U
wIUFvTAQI7KpOh92h9R2ROAhGXLr7iVYdvdk0wnF5QAI1UFA03abZuvQDOyabC4CkGGtsS75uAZh
WSTWFfndkIusMKLorSxoFaU6UYu+3R8xvThdt53dcw/CyqXkBLpTSL3RJ0qRZI1IuUu4vv5wdUNO
0L3NTgU4hIKPB5EHVZWDdUqKelrPXFcdUZiEMTaCPdB6rJOZY05FexKY8BZluVpaeEW5cvTkT4L3
UvlI/sC8p2gbMnMTn3gJlRdjXSQtPiC2R7nt1txDFouMR/vTY1EnB5lUnKHB21gn3S2bBYlcY37w
4SCnrXHeuqCHOBkq2ErJi1LOL9IMqFhN3nPS5T2fZUIrHlxQsFQW9I66JABdxtoqW/dOllHcdbbX
vAc3E9JKf/B6YBVtQDew9/X20ovZQPoWBSUU7meMgjIro3h8vx542T5Mb44K4AuOrxBD7nRAQOG+
I+mp0snrAXUp2LKnDdicf9uU7whDMRPpTzK4EE8PYnUrmiGVvUkfh9nhiCw0ifMHyEKqNJbo+vD7
7cwADNJovGXlOpUYW1WmiBLpdiQbDwuhwQdpZPNRJQDTLHs7sTjOEvW1OFcRbiSMdbw+SzqzPbLp
8Ch13GDnyUT7mj9hfDVLnqrpur+uxfsYBK9zmQqK3MJW8dwSoYjzFdbR0LmDX1s+XiNWHlRcJ3jK
cBFjQhawilD2CbOPcSOcD1+H9JyZtL/uOL08eaQvTXa/29aFEFkugxSv3oPMgdzfMLhnr98F/YYS
dEEDn7LYIaxOTQgxqjBjjsqjt23cnt5gGM8XV6UFQfJpuFUMkyFBvI6NUEqDv6ZgKZqRmjf1zeZV
A4y+O4hWFuKAgR6HGkmMzMqFy3az/4snadja+CQZijKqJeLBG2nXGXNGTtdvPjVvGBnb0wz3tP3L
rIT1pcQzeBx4b7HyLDVoF0MNQ8vS610LX7tvT1fTQTZ53UR295sVDo0PqbQQHCTkQQBAxzgYAesF
7+aKQU88B1uGygZhKbU0BUbaGmUmgvxgT+0c2OTCbP0iPrGyVu9irhCoe6NEWquhDBqgb07G28FH
kiGJYqyvNBUWeUQCVQGCxtuORON4kJ/0gKoU7rZqDkAey8R4oLGBq64EoPbWT8NGkZPOuVNWL9Zy
NC06bmEODgKJy2azJoF95JkVleQ1kPPuBaBR5j9o4da/n6t2h2R7XJKFklTaUJlHR6Qj6J/Jeel8
NbyIFd8gOydDeIcKsBHPgdWGdT6hjKahkcVIHP63I3OB39ELadPf7W7SDgu2LJvFDwCM0LJgiAcv
qmUiUaFyF88dJfNy1D9Q1lAlReSU4Z3g/8LaW7FYJ25cYXZBiW32t21bS9Jro7n1WsoiJpQHqReB
OluSGUg3xBoFa8T7PdwfCcv/t1nRsvTOe9nexiLmdQ/MGHn2SCI8aSGpNQuSPniOqTnhcHP7uvPW
b77eWpC6bUMeBt2xzw6MH5bldt3ygBv7YGgZ6f3xbCBJsk89U0wmebd93viEdyvGIF8PEGquuFKf
BkTgVjRWJ9SCbEfLQPVQ4gsobK8wxVJoxGJe9B32p/DdL11r6Vv+kCojGEj6CPTVz5ZhZPH96gkI
KfzBCcVbpp2zUDc/iZZrwy4oSpu11w4Ye280GqNzvesHU+N+M3kBEbL4tAehBBBIlGl8jFsLFGBg
AMQkU5yzWdXFhyk/Cp/VICTAPeZW5VssjovvNmjDL10R09J1RpBsTSXI6s2cYGjoNzuhYRWWQQQn
8LsnunGxdy/mbXO2QMnN+ybslK+l+QNdLcvKFRgZdGtYDSi1tI1PiKlCIET0k2H09wDN1tsjklhe
dUrrMOf1yJ561Xgl4dfi7wMe4aoGOLTUhyWc/XM2aNhmcw9evttappA8edlGCaQeLWONiTBjQN6f
aqmUpZcv1ANaCTp4V814vyROD3zF/1r/bAYxxuDvhItTUaVV8aAvgLzLLltzbVLeXsaL2/ayEJtB
w0x9tX0ecgPPa6bLN/uoMsW0D29UpdS0UdW+vbfbDNgUZLGg+ZF1x8GWQcdG0Y3GvBY8kpWa6lSn
ZYCjY9Xq6Ca4OgyQqV1o/wronBDWCV9fVqr4myEyIyluHCyx8CZt3578B7rI2WPO5fANbE0kiR6x
rfKokfvSlxpsLR7KGCPQGOquz4KlrHoeRnECeg69BQiGnyEnEB2ED6OAbbc447LggQlDiH+4vBf1
YIrUs2n8F1xWfWBBtzcOGG3gaM6uifiBVERdfuO8kJOiry/7Y+tcQW2+94ryVJ74oxdC6e/3yFC7
SMMcgz5tO9PeyACzXkDQX22NT9zG+A03LAVHOQPbSMgF70eGXzHvTAmBLctRPRkDHGs5NDKg8lmA
LCB2gO5dhkZnZybeTmsK5Aj/BxsPGuGmGN9ZL7EX0mtsKbnTl+aaIRaBpFVZabQY6DALxSJK1z58
tf7NwWTgKOUhLTq7M5uq/oVkpAUumJc1YjtUKSPHy1arnNuWW+42tLqk+WaZlbqqObHI9VuDpl8q
Acic7s4o78JU1AyFWDCQkemlbLxt9EF89gOc8XxdSKfR94y85T0K0Z6+lEH9OkWfezYamZq7f+ks
SU33LQ3spq/+b7cO5YyOCHCHx6LmzdvZGxmzHXLF9jPF9UD8YR6/OqVDJ3mbZp6awDsD6iSPFKc/
prAtsziFV+aUr/Wo0MXzZrxh9SAkDNLyQ/kpWi2PoKIdcKF7RR5eZfWolyOZjHQuR0+pVeFaaB/h
kZ292MamsReiTt7b1m0UPMkLCrC4QoPjNhViIOjH797OKXQdSMC8birDaUwBfW7SabNIcZ+NelWO
/+RneK9mSodjvvDgX6F4upXfgKj2VPUdoPIbT0hIoojYLvx6HqpzENKxEimDcEpH0ve07rWuIMo1
JNOpd4IHTwLt75pM++l8WhuBqGeCyPma98m7cdsRFB3H43p/7NspzOZOnTkMx7XqwX3ojCurDOUM
fqnm1+Qf1fnlwDcGJL8b3hiKvxSyVnMVXT9+UeMB8poVfM8nTT4Em0BP/FMi/b1wj/JbVfx34GAu
Hdwhb29KxxQuE8PhnXPv05Kv+/epcUjD4mPM9W1KO2819lVatPMH0uLBiipoZUUkP29t4P1+aS68
9bRgi+vENpoytOcRGOThsSsFpKdZJvgWjfgJR0rGnosDf/mrgI+yKPeqkUi9YHxSJUImZXu72yT0
p6FEQhwBrmnaMvRyFHyIYLWDa6Q/mT7/HQcbL0Sogk5t9McTMqKszUq5061CttCzIWCscdpxqCCw
SJ9D/sUB/hQ/HmjS531H2SODJzU5fmQ9sRtIzKfQUYtq9YHW3ZWsAro4asufivaCkepIaqWeVLNW
btuheC3DN6xXiDTaKYewp4OnFakayMrUf8IXrRfgq+B5Jgpj4bj6MpxU8xqgWhfihT+wFdwdLgfk
V6bcrjEGf6Pq6WjmHrhfqMAp+76uIGauuWPfkxA8PoAytIZbLlDg/BsifsNKdPo3hOgY4eiK1Zpp
uwWdUCDayXk/IHNQjqzdRBIAjVY55lVmZKSqus3+kRcRueZiK8lcStWsEYTSAG1gyubkzpP5rdyL
RzhEIfdUPMlp/oLoBUFOjsZHyARqp4e0H9XWthlFnDidYKzbERMC7hHzUjOAp1Nnyfs8MFxH2IGy
GjyXyMemVcWudWY15DdWChyKsDbagd2PU+U57vAytrDg5EFk9YSHaZRn7qx1T+8C4QeDK8/FyRnJ
G91zak24JuiADHDsxFB6ZNgRMEhSAs4hI9YGmLoqRtlpXCh/oMpTAlCUGHrhNe2YzgqQGOE663/2
2YpelBBjIeOeDEbFk/WaydMlQ01pu/e1M1N+0b0emDpxGlmycSoZljBHA/UoHi/gRWunweQOOn12
eiuj43n62AKcdR4LbRJlVznBvQ5x2vV8jKk5gA7Z1LSkelUHRCSo7LpGS+MTJmVow0CGrq3q/Uh7
92g2lk1/XDoEGBCsFB/0sjod8/hQqdqr/PclFR8oc7bNleE/aSoxlKkRljG2BmFqM8CLa1ejS2qH
tA7v2BxEvg39Wy9q9El5fSq4feBPW3cixuCDTJ9rWbOiCz8XpR8AzwOJyF7xuAj9iTG4Dau5/bKo
hcxEknpzME/fBxLsSR034ZVSQ9izpPMTZXpA5zdBzJi4ApQm3qYQtoCGiJCVLF6C1cs4Q6j+xXB5
b3x+7idnMvusNix4H9PnJBX9s9W7T4U3D6uObAQ75PjYcRNfPEvyJ5QjhMoRMtEnHHpFJ5dpSP/1
PoE9Jfy4xoZWG4HzCMw9hBLudps72VGqnVjea+LRml1bcwvZZrSJV7rUzitI/SA9+5UIRaemhhdt
KbXJ06s32ztgc2ZfexcbzT/WB0CHPM4RPr8t4YzVAY3IROhfvwp6zr/vnB+lHofW5YXOQa+LAkOq
X+3/BLIs2z1uzou8xMdFMHo1FNIPQoQgPEnJiLRGyMxbTK2Hy3tZw+7+NQNW+b9q07U78VvQeyQy
xvHfZHHZsp7aBFRu3Hu1g2G/794Gc+hOwyP/9COtvPLC2DWpuHOrCquCmOdeOYyJWKPnBnLUV7v8
v/lV338pQQpAWZ0YQUn/3uGu19omXGdyUe/4/PhbHK3cWVz6hccc8jApL8lXC04H1BKV05c8vB4Q
X3GvvOWSGL8DOk5vmbBoVnOsP7RUtrkESeNYMbYBKLn6PenhYUjNZhEhLSJANArqSUJVSApnv4Wh
gpazJRpG4eMVQOOvhQkaxIbFfcpS1cCMP6KzaLfvih+MNgNuumUJoxKTZ9NQHFtA69rFGAx+DPoJ
7BZTSnXYrc0MVhjXi7qlP1/Zmbwl3G57oh7t86eYp7Au7JC3eUn855wbOARYCnYqu6Yzls50iIgN
QDmtQBjERRoRbbOll03g7gUIRlnTDzeEdEvRSvc5oM+3tyEluZT75jHzyHjtAPyR7UhrCRZ+lF/S
fwulCiZs4ZIvtkWIbmbKNImrbEPjuVUFj4JdmeeOjgJAOQbiUJNSbf+FbkIW3UpHg5STnHYR6U/o
FuSf3D9QnSoPee9h1PBaVvUxKgBioJyJY8f0AcLSceBoNR9mPxFArQtWSbsakRgm97hWDIzBmqqe
b2GX2J76bquIh3Wr4WhnVBoJfQbTRFpThuCcaLfhymViZzwGqiFkPy2n7vwptAWTZTLqR40DHuGn
sbnt/3hMiuGVwdTfGnFmQ1vbR4FFSqoVWTsJFeFHkyu2FYGbUymRxQEk6afd1Ml0wpXUTkNuczRd
GaKIwo0TocGVE23/gvqR79rUHhzvCIuvUf/DzkPM7Y9q5XgYAy5htD55R5+qA0aNlDVzkYdJFf1D
HISwup8ts48cNOBABUj9KMuq2leNTn3JHTbaf/af/N546n7fHHovdlIVd4TMhDU94cE4Lxq78SyP
PruAQoKXsYg/BuzXhMfZePUU1lsRI7vEyXp5NHN/v4P4oQYCLTtFG7HZlLbYBb89KQVAalSCxSby
Vwmi2qg/oPzRPhk74Tr5ydTXlLjQK0apAnhKCYvi00LHJ/Hc6BLe0hxQBALn4HevfnrKt++KG1jr
yN3x+fdAMLuAtreG0G/Foy2aEXVhTXLE4ELeyoSNTd/9Lnv/HOow5dSe815tTBBk70/y4KemzUyd
4Nclk7LUPJq/pkNjma6C/zjVqbyfgu1RnM0aoGcKAJof5u5fOb4xUM9IXDmKl9uN3PrPYzWu4m5l
gXeR4mJPITgv4iOA84mKrzpOmzzxkO2+bKEa2v4JnBlvduT3yv6SmyTGLT/rgnGMAWyxmMCl3KS2
VI9HTWa2cHhcYn1M/D2UFXPlLJI0xXVyXjzGxV4YoYXRI5ae5d0f25W+uy8+Cfooow5Zau0j4voz
/+6vtVKn8q9RrQGuIe4Rp7Ts+84wr0Hvuj7TbqCF4iYiybUsOsVhfm/tD2LY+vpPXklZK6sHeqVN
HiUaXJbRqFymPd/4BvyHzHlPol6mJJTiTC+95XLRARD8E7JGdfddRgstphNixlRNUi9tOYH1t0LZ
tF3P/3R3VSYLXl35b4KWmFvSWvkwxtrD8HzAAw75GzVxv2s+gJzzFCEporoHLHUZhrMmUT05yw+x
LPch+jtcd6HEYPazFpNj72Wz57WqKih5rBAcgzMDKp2iEo5CNH+9uyNMhcPUt+Ff+FtVIDRULmFS
N5qvghGIeZuI48r53/ixWTf7m20CrQ/e1F4C+WgvhkytnPnpL2HDHq8tyaHc63pU/S1rPKtCdBRI
YooyAx5+buomlKQvSC/qzhGxIShXAK1Dce0FM2j3qD7PZMjTPNwQb55W7xQi3QdVNWbbPkuS0qhB
2TkgwWG3sL22zL8SYCFJdSFlKrxYXXf15nB3Af9CmhyXT+/QrGteeXhqi2TXVF0P/I/A3hRxLOOJ
TU5B88JS9dZtYC0hmLwGKmmlWA7gDcK0zK43OP4E9/fJ8aWdgy2vsV5n/0H3Elr+g0rL50nFXQLv
guBPPaHLQH39KWbeUtYgGY69pYfjvhecpSs4shjJPtAnXk3xFzGAi/e6Q6wk4kjWVNctvPvt9Crq
MUdfEVy63JYYCFJatBMriUCdBQ/o5FYAqRBLGIUxm9rpB0ns2V6U8pk1x43WDigDfV/jJ8aTOuTh
bs+qSicYqLZd8Ie91hQXLAb44qsF2MZ6e0MwrVG+cGe4tkOJraGq2tj0TH7c7wlsQ1TxtJ3IhmmS
0TrcbMwQGCnnz9KpqnzgwzZ85b9GUNGpQPNt5pz1hxii5zQMZjVJ6YQHOU/9vIbfwYHz5CRSRend
+tlv9ZnJgx9SS0W5ol8qHwRRSLN69X+Gzc9jWCNFLb8mYJ9BNeF8ZuzrWfNQnIV0z6gtU0KKUuCy
DuA7t8syM9BPw2P5tY+GbtI6s7m2eo3efJ+dH1/ZBmGVNA/03dE1x/9oh3aij+IHs8I4iYObvbIq
8FrHeQ1viPNjQAwg4ZR6enyqKrIYBGCeblzL3MO5xR3sWx+ATX5Fk6Zc20KPXRFwI+nY0U4Z4/MK
I7ERaeZk7HUsJztK4zaecNai8lY3stCZRKdT12yJ8Z9z2EtGNOj1yiAHw3Y0du/U5LiG7jjCYqTX
tDh1f26rIJZO5pGfeYyL09q1LwCIhArAxRmUCd17GRVpjZ6nQYZLIpCd0N5KdWjD6g1RzzB567lH
ACMsLxmYJtxM4qbf7t/QuCNTCvGvfVzlkHPSiltJda7EplKgiLK+YCsUurPQJHJ6aQIckQn+LKIj
oOGtfyH8JefJ9qOg/hrwNcUPllsznCKzxotg18RwOAOWeM1YfpcIavCyomxF/LOcmPKwqO11TpMJ
BoC3zwFeatHHtbFPKrpbBxIZrhDlpnhyQUylzgETWQNGLelaNLwxskCus6lfrAehTVg/hzmI0R5x
l3MTf4Wqb/lzxh70v9735YGZ8lEPdPJRDwZ35k506/EOB0ChkMN68sN5NVz7pqP+ms7NWd86377C
XUzJZL887o8xL6sf3smcUUCzbYmPyPFlUKUSGLtGi6GjKaD/LF22UrUat3VrFKkpUx+M25jC4aYo
gZdvawsPw+kwwIcz1jyKLbKsHp3RaC889CGa3WhH0mMtrkTivqntrlHdnUOaKcrHt45bZiQ9YDum
OxIUQlzqnqWuLFcv+DNgQ1LE2YCcgihzP5YtcgL2iSamRCBifmHqUiSQc1Lc+WbuCiByqm5BnkuA
7aNPvh//bfZWk5VteXfjrIAdE/5qvH4HNTv02oTYc9rsQ6gY6K9N3V/O9DAK7SM/6qzxIVicEV0h
OdbxXmkbovP366dLrnaQeALbTcUDOjUhYfygs6LeU2qlUYldTsGKBaT59lWCSpLm7lDp2ROKmVMp
cxHy9K1HRQW1tziqoxI1FrVAkw09qoi9mcXXgtCdbIK+/w442VMMv2rU7SNek6TyNXRZlVGxcUbV
+cYeOIHAp2Vckmmke3/GM1u1r2YPfVCLLkISNETCkIVDRjbL/bswZ7aPUxwnLcsW/mzDhdZXp6ey
HRw/4mElbvD4WQ0n+XXnHEOJrchnxrvEBawdx9NtSys/HIXLOlwpndn0dUKjSnUCVPHayuw4gBEq
QQ21QoAH5WOIRNAQgG9E1E5AEVvLnej0cV73cRWFLTVkgoECBwu3PfsVL/lJtZMIxyEW6xqMDW6c
QSPec7lhKVRkcQHzU9zEoUlPRrMo7WDm6syLN09ljvSHAraSHwyqQ310TII61tSqTZCqaEEswFvJ
xUPCV5nPuRe8NpY0icM3QiyjJONPBN4I/nuqGqzhVg1kX7LUihoVbP3OJPhcxqVPoRKmdrvkZYRy
RfvTXFap6+oc5eV9jadigI7TCjtDzu5ziCuMQMQo4hBUYl2PGUKGmch/GOLVjgPArnshQmQhKnIQ
BHmgVLk4rPJ7bEkyUKlBOCzUysl6tmhJGI7ZC1NI3ZBfAeLZ54a3cOBW9/hB069pD5ohSwXN/H6x
bLo6s5CuzeY3vc0PfvKLMDXZdh7qK0Ci46Ju8uea/DM8/z5QALn40JL8uu2joI83xu3rEF2wck5E
QRoIHTptOCOutpzYbTQtTKZDII3J//2pGLZUzlbxx1y+IIMyEdMZJMrS2qVghHcF4qb791/7GNIl
UnxRNg6JnzCSLRM0V7lgSuhuLPboXnH3GrJNqjA5Khq+BvocLMT27Bo5XmyvoLVLK9jlMr/gORtr
uSiEBJ/Xndtc/JXsUlk8fBoGRmkZ88Aq0oJo1rxUipJWqwVaI/4u5H7F2l1v76psXRRMYG6h6pDH
DBLLucpQnKa7IVv4EfT5taPjEuMFn7kEV0KtunOzY+XHYWzc0yEp5+Bwzd1QyxfVFIQnb6nJFyWq
/eD+YoSdKbgHIFf+tFeq5cCrASBHMls0VJ5E4HMYwsN5Xxpl1++z51Cy3oeMdEbFzBeIsSjKMnB1
qAk+WyaDDPfRXAopmpc3ri4To+2dzLTt/LRao2yeJDPU09scT1m6sZjlVO4RV9I9yOVdFyeKIVjd
ZbkF27sMATJ06QS5aqhkLWZSZ0DLcZDBgN9zxxPxVamjsT7z4M+JDb89ha7lxsmTfAEzbJpftzlB
WjaBDDMyKCQihf6VFqRaj/JjqQesjyY/wh+EEF9ITjK8yHwaZOI8K6h1tx2wzts0TG8zA+V1sJeH
SBchEkhO7+cweRXhGut1DT925davDEyosItLURBwb2QPKEbHcI9qhjb8YzDkzi3K3BCI5R2ZXcub
ygk6PN8ESYHrXAr0hBGLB1D8z/r2RQWqYp4UocSQ64oOWcUDY0co9ErHYLvAxg06VxjZsrfFLh1k
RUivaKxKJZhmCM9VT5ms/cLRZkgeH0Hg67aMz84Va+kMeoANX/CHOoiuzib5jxdj++S39NzsW8B3
taqrRubH6gWHCQtLaLALICgEO82OYtQ/HOOQz0uudYKuytVIdehae+5oSgCzSXmUn4Td7eKspOj1
wSTHx17xGgscEBU9KFgRW2LaDsNsY8CwH0VKrgahCRUtPs6xPcaYahGDJtA1fP6yBavthBzSFSiM
+IoT/sLA4Zp8Hj1EiWJgAB1gzTzw33seeNiyDozIJJNic9fqD4vGvlr1oxa+wtBfJ/khHs3Hiinh
d6Lrt39l5+tJH2IOzRkvc5bTu50CYTMmW83514G/K6BvmxhCkka6Cxrr9y9duwpX+ENZRGLLd1Zc
fP6+UyEWBTjFRUHKLYBuCQ6iyA4D1NPZCU9kaLdocL2Q5EUSvehLLyzfBIBp/vj6ACp0ns1lqw32
4PJ2J6a0yCu6HdrVAyxaE/TN+gPBQpNww834+26ZAwEsgLOAxh5lTDg0KzYX4Ek8DDdr5WKyIgH9
mRRwzaSGRoetGHDN6yFvs82YLorfEBoGr6nq26nq1zGh/S9FXAfbtp1rI38sF//RcGfVbTi3HZYD
byiuT9hYr1fieF1YZVpyLCvkVwvwzRVkFV3qYDS1Gsm9sI+Xw26t5zCQoFV+DbhPkMtUulAe0yVG
pu1334yZG0SC2U/DVTGR2DdOo24SHBJkdImXi03Wa4KQOn+6+eKF+RjSea8wBwOHQuRgtTB11BEq
Ogtw+BdsTJN9v/Q5lSCPKmm3Q91BWH5kWcoeykdBOc+INEbf4MNhsASIerJEfWBEQKvyPy1VUfVp
8loNTneu/zgWSediC9C1i64WDpnZ8WCByaOqjYEeEJkQXnaTWndbyXazrtyAwcPY9xu823GUZILd
XiwXY0J5BWRy4GIUXfozMUoX6j/hl00KgsM+7zJFBlE5qu/cGaKO5FNlLy8fz0FptyZXUE5I7T61
dgeWmoGMytrqeRy1tI2tWGscPs4wEVAtlJVUKTP9shx/Ps3a48xRwlNhrm+KIHGOGSzd/vRDexpD
ksRQ9WyPeELiXs0Zt4+x2aUDx+5SxLMPIUm2+d7wXE4iy/c3junIwNyL21hanYtgMry1W5xh0BjV
l9GV+1G+1Nnp7Ti0f1sVg2j+RHFQYuvOcpWbPuglNwPDWCWw9a1JZJWRIgNJKA89iE+Wn5Qn3nVA
l0dn7UmGubmnhsq4ePR0N9fvfwS83cwcVJhD3M70y1PJqtPFf6Kfd/Upiw39xMaW2hD3Q8whIeGh
Tr8RpgLm4eVaAj/HnkDSZkL4LS/IWqmY4YYO4gz95X1/LZfnPkrR2xJKFOV77pyevN6BJAbS5+R5
S2M6qiNUp5Y2q5OFNukm4AeUE/WpwG+2s1KenntP2ZC+ENpxRMaHn0EKDpyIE3gbaCxz+lk/CW44
LFX7nDe9xNpQwaXYvgfywCM6cBcCilrRoRNCBOBG3j9Eo0ZoZ1e642pgnQuW1+U+BsYRoxWwBz0K
Wth0XUC6RVmqoX2A8FMbvO7TD/PbB/lcxQSIQMDuJO/v3W12V5pmqLKzsjoWYCT5L6XRgZJi9YLU
+aY8BoMWq5JooKKWDO/kUiULzFd+mBzXG1OhsiLwFssZKsAAArHXQQ4whvPd+UbeTuV/86zh4CpI
jYTiGJCdbq55ncIXPf6AzmbXvmf47mYmHb+oGq7jRVEUKNPnAMAky6uGdc7mfASPDLnU5dMP3i+n
lnk5/fijh32hNShOg0p4DR4SEY58q5W6TG5KcvkuYg94qX7vGrwm0x3KL7JO2xBQY0sq5lZlf1G1
MKvwXYL9nB3nHUqbrOI/BheJeYmG344tZG1wzX7rU0VyZ5FGMyWFmNQT+z94PKGVn1qat8HlMct3
lgax1EAwzU1UkqKsxmjVUGQR6qjyxewTo5nWsvkaqnZKCA76OofJWBJXs/me+bigOFLxo+v/E2Cs
C0+ukOqdsawXGywIfhVgD+a6F+V7MVCJZOCGfsSXtEEYaxqzZ4nx5+Xb96CvEH9nH9LSUxHiVjKU
K3mjK02IxECNggKRnyx/6ZHl3OlPXVWUYzGpxAe1xpMrr1Vbc7OJtSWCl7r73lYo/k/qT2HNM9kl
Y2L/8iTWtcWatt57gCFeCj/XtRl51Y5EOTbe8VG7hYSRygzZ7A8d0hTSXScGNMqd0cbi+wPL4lIy
qHxKmnCl08iFl/cEAJ85RSaEfUbrW3Q9jJ86/mHz6zGJm3nGtXm+yh5fxhj24WsS31oAq/iwCCah
+qk1RqBk4kp4hewZ0iDU25sQVphgf+W1bOTZJXiHGBSFXk1NDn5n78fy1qQktjIb+aBVl9WGmY4W
cSTeD83JWj5JNdAPdylS/+PW9OVSH3SwsgnipI4WdAMyqJAdChWtBHghiqmRKGuOCw2QO+T/TiiV
O9cTMGvCdJMYI/3J+ns1xSdiLVAfCGJalkI5fmJKwren3H0IgENlF9MKa6YArtrYtwNjLCxq7IWF
RXahxUkOANdq1EUKFMV1RGToBvwDikokWxFA1+6N+zbtbqdbh9tAjpkwNlHLP7WDIe1AcWttWgvh
lJItdvDsuuLBjvT1eeMwJ2HfUuEyGz3A3RkxeYU60NRE2MX55DgxgN+mAhjxxT+3av/nGVduguER
EhzHDQrAquwW76aqOxcXV+zxWW0zNz3eV2Ops7bb5M5C/CGVHPNimZaPQgZO/+EZq8Y+5fT9LMTL
fg//ioUaBM/d6qveU0LcXey+V1mLDLs+6cNAXuEuYu6wX3QZvcVqKanDVRgr56iKuvIXQMvFY3cP
x7NceYuXl/gaX5jwbiZe65egEX4ty3S2PeqwKpEfqb51aeS3FSjXP/CPa3350zqNJUTVZTRe7a+9
PL0fgAgUbK2tNsfGpZrk0qZPY7kj6DS1JXtY94GKyarEo4u+M0nVEKjCo0Kjk6QnwAQQ9t0J9V/5
+inyoc9tjvu6G/3V/BWrq/hsBGIgQYSHeNKhWM6N9Hf5wcD4ehSUSyu9HliSMJoWvQl1Tq/vUqV+
NHIUbsXzftpYri0Tk//Ct8aE9N7kA3epD31+yi8j2y3M1oPuWzn0FIgTEr0IDpDfwEm4COrDdhs3
J5t3gtv3ozXAkxTXqvD0ynNELX+90MT//BMNIYylB93nsYP5WgIJ2ZG5ok20t9B/XjcQO2Hx6wYV
mx/P7ZrxBsCUx/sG00e+GemY/Pb9Rtmeoq7rSGKojo8wAeOdN9YcbsVl4hxTatDNR8E5yDVsz6L2
3MUHzbyD0E6DblGfEtfT6/Cri6Eiy0Pef0VnHJKgYiNSYCdRsKCbvsGAcHYd6w92xEJPcJHbMqEc
F1acQD8dVDqBRB8hD2zTumOoiIWBwgMhRz+S9O3KHqBkQl0mLkZGJOTJfvmIyS6Hn8QEILRxgJDu
P3nsxEX6brSQHDzdDg1vA5Bnni/EsubMoV9XlydLjdWCE2ORIFUCIM3k674zZXe5n1xPrAlVTO52
R9BxYULAG13w0bOjfF6KcWOTxzaum6ikSoSjuEVVAXp/POqoWuUHlu7b76HgGGYQVSJnx9wD5rT+
Niuwj8frYZaUSqe3SClGp5WugUBhe/lAdYS39xC/HaMJfvvX4N5jq9/VZbDuk6ctCp1pHCZia/3q
xf9qYbTWfffQPFXofTABBSaYstSF5D843GGEWBcPGTBA7AolAnZZrjUQAmq8Ze1MyvOsvsEGy68s
TzyH3EpuUTW67od5HtlDlvSnwG+5QPTU9HLZQbVcqPIpbrm5jzczSNA7eKZ+qdWTvr9/B5sddoKa
M+2wTcnk2bUeHKpxngj/NN3TauMg6SpUUFrEqi0l9uQtkG5FiBd337aWwVZOiGUoXjWZkkpyZ2Pm
6HDv2Dn/GqKmBvMwODu2FSvHP82JNhcZ+qpwpcgTFjEpAMg6ALzoKFeMaY348+y8xu+Xrky4rzZ3
7riyYAWBDeWerCmclO4pK7R2QmxvRDe7WdhIXrVRZtxA4PHgLTPPN4NEAWlnvy8MBZp0kQA5mGPb
A+ea+uTMgkbPEAA1shQWHgSFFW8E2SjGQMfjQvB4SPeuZ3DNvTwA273Xzr+j5j5inQ6akuO6cuQ8
WGe1pFHkHmK3S72mE3uRxycm0e5Lh8CX5hJUM4yTXQSM/AemgJwyFXH4jteL5OiLvLq9+Qr6mNaG
h/6gYWUaNbqoQbYBMenvqQLj7M5dMJhzvtOX5DqdU9RhS4WRwf/Adz+brQANdfK6ip+JkbDFTiNb
I6AOrIaIhpePUAenApODwlyXlnzS6HPt1sHvR+CwfhOxSPXf8ZU7sI3YtK9XtvRLIUI9kHXyxKkZ
3tErkHjPqwA1ykl9z/5AILGkCQ4YXegXrOjmOQEFzj6nzHiMPXjzYBqTo2VJYPoZCPzlG05M5rD2
CWrZa0CWUGXnIJEUhoWQWlROFK5lPUi6jMwwyyF88B+CDoLhCc6Tx+wu47CI+4lRe4Ku9fqB1jo4
j7X/aqNaXwVsJW4EsY90l+yzgokDnZt65xSI48RL6TC1LQldPXAjrikQf9wuP5lLrA6s4vs+88VD
/jDc+zRmAmHH2PWyPFC22l7EgKodiRIBaI9EFOFTqQu4FPJn+zAf2AcBe08zYJxRU0FJxWHGtXB/
fhOXnPPt02r0+R5F+LZ7zz/DFC7C/yLkE788VoEilIv16yXTt/oFn45P3ZtjAr8Noh0gmyw5zag3
lyzXY6NkDQQ+BiTWZ1tBoa0IQYfvWlwCV/cESKAOVP9TWE1NrqVfP5MK95Ex1qMMjbsRVEK21uTz
3iOyxu15thm2iQK+zCmiPyJLJisgq7mFRcQkxHCTkNsRNGzhzW7qMgA0VMHu/Fe8VBuNLs2SDKPy
1UttJBtPR60oGFM+sNp9VANEhop67MMhYsvgi40UZyGMLoxVZUCVMzJl1vVLR3x/Ptr/q/ZlT7MF
uxtLJ1h/o5sniJiqGGvFAIIln2SaS9PLpuu7LYeZwbJlnVNox96FqqdgE/PmVhj85sX0JtFVJ4wz
pYG4XJCrnu9ensjHGb2K9sbI7T6DjGn7agM6o9AKTCBS+diy9DswEoFHD+6EDke/czIGmWDRCX1j
rF6aZlfDaAyL4TZRb0KBMgJWsVsC5Jm9k2Y9PTpPUw2sKeQWRAE6KxRFHrkuB9rQ39eTPGeaGo3E
PNUfqn6dW+YE9EUu4bivhw3AqOWRT54+sBn2yKfd5KVYAmLtGydKFoOC6qKltcuytI+q3ytPt0Td
JfKKG1oq1Ehnph2obNEtgOLb8B8rJnfWsJrX6jOonESLQ5UGG07/uhVNI8nG5Ib2Zzi2tiMSLZgb
A0L2cZC5BJO3jHVknqVL3bZmfiba/DPiEVjq0ReQU/VB14bkXho8wsYiKH9LUtQ/mKlihiZgleKe
/u5MMzaMrZAWGqYU8eT/2+GNI4nCKBNaAA7uCrBSUgf5GedtL09EMvCFzp7XHM2apC+ghVUgs9UB
VNj1m+j8F4ddphXQz88z8LsqacHvGQL0RKltsIX7/fiwVPAL3G62R2qHj9tthbNWjol2UdOhPmm9
ys+WlY69xpt0k7BKThJ/j1203EHhlOGNDzDfCWBeHGc41SV72Plj8B9KkWsB50BT1aQdeWQgYQj9
NMkwV5zm7Hq/uk7PRx0Yrdwvam947RCeo+6XVs6J+LnFCU8LBA7kWWwCkk9RpMjzDbr7XaewtNhu
L3wRF3td5tPTtQs+Sm7mQ+JocIMzKumphTf/w+AUwDx0+egd3UoWNTOXhviuq8hC/sm3p0SzJkHb
7XloRLAk5mR0nJ/6DnPBeWslqLoxxGTfspfnSi68FgscTK9ZfIFFyeibz+54cYyqmYAvVbZlFfj5
PJyzU3bhVeFiYbbZb+96Ma4mnAGE3esIKgMIML6hQ3VuRte7IqZj7TmY4Dnl0Nz1WFw7QzabjlyU
G1mPG6ddgFW1A6WQsS0ZrSzbemsdU2AMrbalYq3MvMcAZWO86xxW2MkfF4rKj6THlSfqYRsK6whG
WCNqpWPP3g9DVidoaeZkPCiUAPTSg7QGQY2tEb8PcKw5ZzlMxePUglLVdj4DJrIPbHHRRE7G0oYz
s5+uRlGrwOqTp5RETz5y6tniUHpoxAXcKLK+1TVaQrWAJulZA6TdNgoyuWvkF4+8tNL1x03mTkEC
7H5958BwsfZcjZpiHcvWJx95snyhsanfIXnjmeU81c/H0YeKAeHBB6tYXRojNgryWSaRbikEV3vv
RDVOVNp03cAl+kPfHCLMmRVqRcwS2KHA8Lmb1jEezszX9gilZ3UgC1+MqtTWFTPjXe0iqP7prGz2
SQrcrhgnmVLm2xmNKpJq8ZvZN4nWZyKWDIPslBQM+S4M1YfVofDbd2YNa1g9hvJR9QcjCWs86XCs
W4TVRCTM0FD95V7z2z8IcwXbg/cRaDdZPWi+IvXmG0AJAIBwFrC+TnufU3dt2B2S/MnMlO3rVosP
6rJ1n1KbxPS5T4XPfBhxWCchAqyrgQnyVROBKBJIR2KyYNlql99lyA1yrgttdA//700eVhp+Qvg4
73lPkI+Xj/95rqt7YaAJ1sn2HFmHA/G/7RTh2pPOEX+ysw08WopzVZ204wbGrvN0k7WOrBELzHD5
aHvpGJLDTog2i5/dhF5v3ieiCUC3cwB0/GwEmKa8Hgj92EYE+ULLVYqKxQ1h6ViMvKdbAcEv2zz1
5lAiB7EDRXG1GdYHCPBivh1vi+GAHabEEk0URxNT2PyrZOwjws84Dvpc2L1fcbfNl37N2t79njMW
gk9WqORtYB5AjVaIFiBU+e5Is8IKAqVArbnKgibggitxD5XYP1QkaRMUw/uXjJxdy6JVN0w0DYqf
iUKNF7e8KnTbzAjjUo7WzMFZ9jBiWwQm6Bl/+P25nzStpvVU8ow5I443wywuHikI2FBBk6aojEXI
L1WHfKhAh6ngeZ3paHleZIHxxmXozQsd2iK0L2imj6P7rjhXswnezsNN1nGHxUeHao9isDK8oYqk
ifkYXH5HuLSlVfLBeXO/q8R914DxOeaApbsAfZOxPR9YrH3w2yAJ9++JD0asUbsbJlyolULKHkFS
vMc+XZMXReh2DZ79FV8J9D4oVmHNHXPM2ji7wi8lAmHJlSKGqVPUkuylakPI7e2h43ihL4cJXuPp
pCSZZ65p+dRStM/hionP/lfqU9V5Lq6Tl0uHgAPwRrQjd3mCx+PC98b72CNZtYYMJP7lEZCeqlxa
iKRFvGCvDN2i9/PsRDgu9aX2cVvGQTt72a/Kju2qcaskrzrE39b4CNdlBj0ocL7T/rwFBnICn1pH
+r+3fEJDK2COHHjd9WuNrMcIop/9Pj45mpCkWAwSOcj1yPr3cwVtudoT+J/3J+kmXWjThEVNTYx1
uChoYuBP9DM+TJx3LtTUwd90q3OHo8EeMsWuhM+GVpiJGEyxKXVqCtSnZRscUnQtr9Hr1d/Np8eq
6mzVv5e/jRhVsnioKmqQnGwyU7eYJbweQMom/OjsnobkDRNR2nrXAvJXOcoxF+H2WP5LgA7j1WhI
cSIjhg0dr107NERy4RgivRBu2HOEtQ5MJ6TXlwDgLgLm/mEAJGbhnHlLDrSHUbAMsnvG3RXkSS/e
pONG/6nPfBKkSuYtHgGcZI9I5tSprykC3ZTPEcC8LkJhTPLVGAWL52SFk2mVprggvOXw+JfgQelk
ysz2anVRw7b/h1iEG/5ZtZpSOEs7Fbqo8k7iDrdikkG8qV5whiCduUuR+u/VLVS+zX5wsY6RuFrX
N0ygH+DX8jjz1BDB+knVd9COpF3nP7TKXYPr+11R85rcXpemns/EChXWL897PZkPf4aAg3zYc+Mx
85GVdkhtQR9HJTL32YTvzvI1oiRdqL3EQzR3r+L7dZRjCw58lO0AoOnHtCatLj55h1lgCfKBdTmf
8IHJoCZlLPnHEJ3BPnrLo64ypJbSe7UtSq3DViqUa+2RSef5/idJ9ED3ty/gBulXwMCGtnWkz4x2
nxuaJyNhgnXsCEeSi+A55w53Th2kgi+qVHWiaPKyV9oDWAzt1azRbNrQCWJ7nAUMPmac0gQvDZvm
Q9yqiIciz4HuptImxo6i2aOULBiCBKY1gt9owW8hIZFD1F9gQJr5+M9Vufj4Vn9R2Ci3tcglktd8
OGm/iiJdJefc5DhP0v6Zy48LCo5c6jpMcqrYxMPRCegdOSKNTvK2iRp/c+EC2Qurt0DejCz6QSXr
79WLW0zNmqF9G/ZTpNiYbLxs5lCpWB5cBXr8nm738+7A6VGJrEfNrRNOvOIAozy8ZThpqh33CgKh
vTEDKGp7H4m3adRQk88a2pjciaEhszYuP5NkTXgG/9VNaWD57SL4ooKjpxcPDOvELm+Lqh/fU1qJ
kN3boIxARO26uKMOKq+Jnfv0qNjG+R3PfF8RFAXKL5hQYn+HICYxlJuI7OM2aFMCb4d9iAa9AhAO
Yh8p7mkQ8O0rjrARysvSz2l/Mj3aSIpyrjdR+Sn3rsA+jyEk5/sYbROvKPD6O7nT9UoJMI7sneU7
Us1+/4/m7avXIeVsz2jwQFWtS916AWUg2oYphbhu66oeoDj52/VOtsfiez9BiY5Q8wUsDB239InK
u5Tmq2znYmInLJCC2gFm6sx3/tff3rV79KltevPI0IY53U3IXS5OdWffiX3zk1JgkquOdYoQl9An
WBD1wtgF/NE40vxurynf0VKV0efg737Awyc77Pj5682A0rXRjCSoQtZx4mFR9vCN4nAmRXLsK5qe
4254JSc5t6ZWyRAp23PhMHMOiqpeQG9Ly8U94fi5sL+j7BLyqlVofW6+53uxAJhgVRRXCmHMeO/b
M7QmrbCU3woNvkA1kwbGkyhjudRbKaUQvQlFJGnbW2dg6Nst3oLbfOvodsbZTZo0CcGbtT4omsqO
EXzdQagS1FD1JXwKr2SVJratTMqIHNbHAhFkjaT+OeavQm7NuWGD9Ht4O5qZnkQ9oxdcsTDySpHv
HfacJqDUwXB/2lZPq33qqE/ar5N5yjpn55psWnwmNMgyAcz1l5KZQihARLTAzyKpa09V4X5N/PsA
IibjuHF3TqhoR6tp2dJH6XCqtN6bYMWMiZ3a9GhfZjMhyK5in3ajXdrD7/tiPjfniYr0YyOJpAow
P4c3dAWnip0Z/l1fi7wrH8hrWAi60rHgUpPR6aUXn4J0GkTVCsU6Ig9cDGVRxC+GIk7NvB3pGSTa
KbnTzb2bhpboP3T2UwzNU578ujzqZBXPrFmMpe6LdtFUYdPs/Sp6RzfXagrVndn5lC0fYjW3OymX
1Un6Uq7L+7iBfMpR99AJpC+ry/YTDsBEXSI5r1ReAOmbqAjq8j3XlR8DswIIyWEh9B68ednFDXiJ
ZZpFTYuXzCjeXxnl1EDuwjUxdq1ICHr6tuuyoOzhjePfVg4/NKwTyoIjHy6nbQ9dwkcwHp6Fonno
vtsbxCNpLZraA1u4FPdhrvcM6Kx8e9a4cNmj0yeivED/fRB4LE81SjfqmVl5h2gHH2tOEotStzK6
+urciZAFMBH6bwBEh0WLbZ2f15lyxfQByILrSr+7aznLYc8S6T0G5l71UGXoddX0xSiTcbPeDBC3
PN6tzLwZKOElGmqGznLJ62XbYj3hhly8xlu7YnJB3OfVtG8LvCg32n0gB8oGearSRVxnMG+woZ1w
N27NhIjPpPdwwYCn4Pb+qGuuzukydV+Z3vcwc0FieYuEVth8nbbr3QP5W4kEL0GakcMSOPRt1MrO
/K5B4ogTfp4SJiQMrlVCvml5kuMCvhQbHUX3fjWKMa/BgwR73kaC4ZRrszQOSY38Q+WwFikbru3D
zJX9aBa6lj/WqUK80jzZYzbk8YOoyonk095J8V8VHRsC8fiQRkCGLUWb357LBn3Vn3fdVBAU7iIZ
o8wAkQhMjaShGY2t0yrs3PfONYjXT541EKTD9E9H7YTkzlyCYjgoEqmA78x5eOC8MTIdGGms61oH
B/JGd9aXm1yKZHPskvT50whpqBnZPj3q1KEYyfeeKlsimMiz/eZpBoK6pTffdcZYF5HkiHdxONJ8
iFQMj/Ep3hPF/Tlt5KnR6/6hC334/i08xqk0lWIJBOP3R10lS4HFjw+HGqvnt22m1A4suqy3cpIC
10k7/dFhUhavAsexCutR5IDdUet588mwv2RuDrofIyW/9J1tf7HpJPBqnKtxFprDa3qGbPl/6dTe
9Tb3izgFt7t/TdW549b7K0nU8bbCRqAjC7Nx0u7RxojypOI8yqiD+c1phy8Jnxlg8+WJajb7nBkq
vIzJP6Dap985o0qCe4z81zjGnEAhsWCeaZK1KzPBC8Wc4c1pu70Dzpk5vxAK6y24uPDK8XxMesPr
S8+/5pihchShdvi02BOnkAvxnrT7uDhj1x5E8qCBR5zNIYQVVjGdS4K0SROzgspytlitR5joDiP8
s2JPewwynosPPiNrmA9/bHm7HXfqs1d0KNJn1ZJXVjZAjrSxXiWAB4GsL5nNZu9qSoAvuqCH9JTT
2QX1sLOLqw5DIqhqL04G8/eCkPLkJmrRoj4KEAwg2UC3ShcwVlw4+EFvzYcG6NVEzw1Cw/xNeQ5G
PpTGojTJpzwvO3D1WLfVPg3RKqhp04J6kOubw3O3gDUZXqb00Gu4p9IdPO/GtqfJZOzkr9UPFneh
T7ZFKjALKWoEX39c5+go/i4KovdJ0qFTM0f69uARVK7zfxUaQFnHXkr7G87mRQ7vpKMeCY7i2Kgk
UszzMVyb+q2+VYhaDNbnIXFcGAMFXko4kSJvvV4x1BPxXGJGYS6nhLwA+tezywT8+H4GP8MoRfgv
XZ5NYRu2Jy6VahAtSf/t3mnZuxnbuZ1bktN8mzI8cycir7xDpMJ7xeOmUeyzCvmoG2ZZcey+CgK7
7G4WkpQcmqRfcJz5enwFEbX+NeGvjZ0r0sXaXX6sOrFx9TS+/PT401xpXgD2XXjKEC28dM0+yWWT
jV7roFIFymAqUXjo/U8keKBCMzfdVYECadJl7FFgowvJzh4kPOKT5YVcyZgWfO1UOyJljSmBz9t8
8l3oWMow47re6yUiAKaxbryTcbjeYU9Cy5qvRoqqgtW2cbRYLifjzAr3kw3tvqOI0FmypzoXbWdy
tVRhlXISuvTfj+/bGGAbEtJbAJbg0C7koouqVJYw7Yh8kHSxCT50YU6ppJ2ortMHNohWvL5f7+kq
ANwmy6V1AvyTvSapf0yNG5qGEedXEvLeQt9tUGTlesVOfNaQoTd5/HQGdMTyGDnbfx2gj/Tl4D2t
eqoz+JXqU2YKnd+N8GacB9CyNCyPqfk/woSsLW1tDRijtmTiRrypmAGkm/mb/5GawOp4v+oNA6IH
j15ZikNeWz+GRqOAEwBI4p+0rbmfcFMoePoCtddcLFbRZiDhWOJtPHY5Bwl8CEQVBz2bfJuVieyz
yd1mTd8+vim/FEKxbywQxnfaktM1pjwQvn42NVz3n1HTSUcn5qYT268N8+BXXaIH9hBdFnHa8VcJ
J8NpteHCSJn0ocGc/DHzq+1GBRYY0o1VNkZ9W0+0lS/wyjiELM1GQYuPohzQ+VO9qKVbdtvLyiSS
u0KJH9JFmUVZaoC/Jz2kVF9iH1ZOHCB1XJJZRHG6r9Lu//lOJNkk1LF98WkRjBqXrJHbw3TL8lV6
ZGoAEngIoCdqmMBudclXNZF6mJa4OppK1B/UU+Lg6FdMEiVx2fd81kFOH7mmHzZHkvGpWkDM5bN7
ThTsNXJSBjfgZRj+sZNAEBun8rDVqKKQ9vv0xQ56SjxKb2hhKb9RzJ4q3locXXDDwnSsoW44V5no
vEd36hZHA6LEUXfXPoqr2jdsiUdfgkVBNCBLP3cZTvX7sQ1VLX2mDGKZk/B7F3gvvOzvlWu8ctTN
Rw1LJuu8PgyxouAJW7AkYRB786GuaW25OucmmGd6HacOUhmxeOOkFg6kzsJawGyitLlcMkT/AOK4
Yu6aXpDdWa/4olFILGPr5iO9sJ4AawKeyo0yMl1B/X4cPNPcpe4wBT0B4i81/e8fAf3cdSKeweRZ
HqOh1iJF14XsjCZbS8W7FhJ084cFg1tU5Z9Atdp4GlJiHPdawOFdSs5xgvtJauKeULNXtzvLt2wS
T+ZMtHrLYj6xWtWkKYdnb3IH6vIqcwWgqrqB0guwXE2jPvLeqOwNxOlNWfPDlBCsqYv5GFt459R+
G3QrFA3f2pYAwzUj4YIvXvdvSvaQv8b+We/Loz7PGbX1ksV00u2fNay2kZyn3B2vH+uI8jmSF3pz
vNWLQZWzVRSIjWk6549L6hKeYZbvV5AVsUb3O09/W0WS6/f80pfMC9fQyouZ8sBSw1QFd0Y3doxr
tof0OjzOCHx1wBjb/0H4AsWIEmCRKR0DTBZrMYS4YQfjgzTzNDqwEoY7LVfnEy00hi8zhPz3Zw0E
bIB1zG96/BitR0VE9+n3dBnVl9n5Gzrz7OXTJ4ZFkyZOp7lHGLCLWUTO6vKTILeZ6U6sI4y9rBIA
mZgZdE0Xl3Ome4czlAZdywxMQ0klZ1G1TtIj/SRgG9JoN9g5TBM72x5C+lUPqSs4sP7JC5uk665p
IsKqr4OM6A69qjXFMW/6FJ92TOoBOTWWAaJdISuMWObROqgyM/PohCG3yAqP1ZQ4dS/aVkjYzOL8
Ce10GTg+jbFf1WWS4jJnonm0vr82YBqyoEdftepn/RtInOzQFexpQxJlOiKqFcsuILlJJbSeewAv
IE4uWMTTOXLDL+eOqYoqyPhNXbNNcHBleaEl8sRQpPPFoAo3jp1Te6i+RaoUpsiM+ruymKX75I4c
MpWc2stMSrf12fnjNS9o1pA4BE3+1ESuLGG67bHSWprRL0oV5cCVPEpfKzrF4eVDh3kRWh//nriz
JPrsysqJIdgO2lHqS8MNj1lBk9NqcjvpYi1gy3zf//av3yKId/CLoR+JXJnqBCDS8Z3+EVHlVSdA
umMWCS0KbEOzQ4tsQt7UwF35l3UMp4Ipuz5biTPJ0dqdg523HM3Cd9ZGcDsTz4Smul/O3HwiYjt1
XWhSq0mNUkGdP2xGiN6zGdgTeSKmgw0JPpPbza0I2aKu6fpMrgm7Solk0zf8gA2/4BD58atLfUuL
IsUVwJrlf08RU+xyQ//IQe4l2vgYiY4ZXeDD4iCKPnFDhV2zBkTr76rJofBpNgqjqpAnx6St/KzU
DZjunBOMcdocSB8YlWypjXyPB0SQUNePdk8Xl5gQu+zvx1TqNSAcw3GFu5PScQBBhw/mUyfKBQ8t
6hj4oUUlBFEV8UUXtYUaiwZRr1XRPATW/rWUZbbTsivXpGGNxDW2y30SJCyflnTFa94Lu5IHIlIv
3GGTJroQRHn8Ef+1Ykh/WuilY0IwT1s9GH7yPTZRuGmahzNOluGuYZKMs/keBcxAHMCOd4kvKp+M
GRrFxAYMTBOoshFB5y43h+qa+4lZDn2SamAMPXQdyO68uX047ZSj0dZkwJu+Zj2HpE15IbbG1AVH
GyIQtwqeb6whPrY53F4gOoldkX4XRpvBOePDHguTsUQxLu1tmzanH/+jEMge68GjD83hBgBgHlxl
eWNs8HCs9qcQ23Y6AAn2CyPhdw3SAk8lljnb03D+PekFCr7F+0OaJZuHdoauh7x3diQD3AHxEL6S
JPnQR5dY5T4q0JAUZVUci2aqSGjwFS73hvu1BVaj2q3QU/UV6Oj+HDwDx+RqCXgP65riZ9pj5lS1
vc/94RCpHkLI3zcfu5DLE6PgHzs1Ht+dj0LdrF3RBAES9mjpjr8ulX5G/xZmLq6+qmE/Comxvp7R
sj5u3I7Ll0lLOeaZGXh8pJ1Q7J2LqosW5koC2+3rqQxJ49tGwFD1L1tKZD9ja16PSVtJShYWkaCB
LSuGchlGSP+zoXzoAX520ZNag5gqV3NJKoq4Ij1TUQJTv1DAeSLiT1exwtEKNah/8zvIiHsHSTQm
zqgoFn+beL7LhbymlqUW5C8OHw0MxVnrDlEz3lRnikbL7ZHeZ/q9rgXiuQ3Ig7NOV2B3QELm70wW
tNgpIeCa907euctd4TeDOQqsFfGRn0lDMsQCkAVanh9DP+cCsTKv6/HPdGIgnarBy3kqbuPLSMsK
ghdz4Hj3kgV7E/4S6+fbmQrMdOJua7l9ehaMerKWUwZT0iqUbXjY0KfM878PLCCtv5IMnu6q0p0d
PzcdhMMHxqkI54O9cBFiqIkq4aPz86DSzwDQtMdkcoZjhru0PK2Nnmo0llJtwI9Y7rDVnU2piL8b
81P957MG+R46xp8ugt/mX5Gq3LWiydVeHT4ntlLv2pfd/xzkKpSGKXj4Micit4ktr/JA7bpOsHeB
ViNr46iv3PE2fm4NvTWDYwa/RTIVxTMxIQ8Q2anTrr4YbOliLLois0nYacuazMd13MLSU38ib2VI
RADOqXUiJTFsiykcuWQi6TxoGe6OHOwQkvEImOOn1JIElFpHMJNHJc5wO9Lll2mnXiNzl2R3Y/2z
EMJGpZjWp92WDJijBt+Opk1sk4cyQl9Xm5e4lxR1jQ/nin/VpdwC6jaDVwsVZe8wNr2nYespf9tX
/YGEbiO71RUqItWdYH0bazzSCMUk7lzp/XfT99MWDpn/PcSZoMzs4s5PgK4Av5kDqjwTh2SL4abu
MTsqcb1xuaYPEgXpUOKa9/q3olRO28IrVlZDDWf3UVDprmA5SDKoOP9EMqyqg9Ii/2HB4iK9vPVt
xtkHpcK5D4A+kW2dAXV35qhjAZ2bp0sL2UvWOI2VMjA997G3ojRK8GNa4B26SR+BmpXadaLKfqJj
k/R75pruHCdcKpMyKQ5m94vJuw0AW0KoM4HpZfWTR0x3Q1ECJVvUBHndsQnMlHOxWauzUNFhPqYD
yQdmHckvY3JkRNzUUnyty3Is9GqyLOLbG4Ns4GFxUsA1l+8jqvDHQwCTiWqKZ/gULtR5lHaN6XcT
vDPYY/7v3r/C/BfomzOmE8i5WGWrObabR+W3EUvBULkL5aJ7Kv3CHgXhIjxdP/7NEmR+pxys71xd
MWwTrIJT8bVxjGQo+PnmlVsiydWTlwE+BXhY0p/rngQ+flGB1IRLAml8Qj0Vty1/6Er+fg6cIW/V
Se6yHrbqAS2KW/MDLqgzH0pF0iIbrua8oxW2Aw7I4t2SwfW8i6yCDT/tRSoAl2H+qrRyNCJYx8wL
eBl4B7jD6UKMSXr6qnx6yW0xd4og6DjJvuEgnHES+VGu/lbrxGeJAkni4/iTUmPuA41Pt3nlvgd8
+asWcJveGyoe7X4McNgNrDdDK+MvNY7XDbq8sNevZlMcxk/M+0K2N4dyA1dCKlnv/LhcCiB3bPJc
tbJ6tP9aoETK36LI8HHjLPvSG7P40Y2P0c5oHX6fDafQjRiMhjO+9TZDx7Nf8goAUffe8F1dHgFa
A5c/jDSEYnxDKP3mzFk+rXaS/0T1h4nNwDbH2Czybc7xhFz4ievjVtySQyowam2hS0py+Ff4qRIf
POtdLn686ZVsSxN8nl/bfWg4HTlOYgXnmTWZ1FqAGgzW/DYhNO+i18gzO8D34fX/39k0nbwih3A+
KogH4UC1PFf8RSEL2zblip35gZXtdTkDmiMAjUutKYC/tjktPNM/T4Nw6xaasKERZFQ0zZiYEKfV
NQZeN5EpUA1dxb9kvpXVBoj/3zyDryqr7GnHvtB5+bpsfOkYc/8SOIXS1Rph6F5cezXRGBfNv8GG
ha58ZXlI1KPMm9LWNa+gZ73Nv9iCIYYpf3wXaMF2sMQfRSx9rEPTfZb6dz+HUWG/34F9YDqt9HYh
Ht4Z4NUOENY/scsSS67o3eTT7Q8uI6Hd8WX4wbm0pgDVsL/lJ4BL2EtnyNiDUZlx7f+d2nQnpck7
XtF7fLdTxxhQXtflHChqSQYJO/XOwG3Or3o9MEv4vhDCT631DRXdsJcU2vAimOd2xNXN9ZvwNetJ
0uXMlPk/dPTwvY6rAY9koaZ9H170q6xmBKtG6WtZM+jPGYF64/y2eztOSBNm/Qb1F5mBjMP7EQS7
GTHJKpQZ8j1MbH2UCOHz8GRE3vpGlYXqxt6EZ6BaRYi1K9JRe6erER/uMNe4klT+gpnqNZ0IqtJN
Q+sVupzRhFXY7CCzivmf3SdZ+REtKbpqS5w1CEl+nJuILcHRhulKNDYrqX+8wBkd4IXbvhWTdkPX
op/m+eMkzR+9xUeCBFjyNDr+2aBjj8O7j2hYk9qmyPRmNLLq3MSF8Rh98e/lRHzz9KRodXywhHxj
zM62z1IMmq3NQnyklb9G1CCSliJIbx7373VGwxbaWk3pqi1r0ido63cp0WyMaS8a+cW6LqTkQqOg
2U+CynGmmp+XbpSPBIJIlcJ/JZna4jC2ue4OPH3IZ6JDem3CmwXcu8iju6GsKNexkYZfs/j+b12Z
YycWra/7UArpvFBVf3TYN5KXmRoEwv+2y+ozmmqbdMG+FjybnN4h3ikKhbOZA3PFK6F0gGz+/53D
28sZcbwRnujuehWc5ckbavrvl3TRd8TA65AgDTGvq9IKgL7hAfB7eRBmLa0rhGeRld6EO/1iiEE8
N/lf+7DL9XT8Zo3ZUNzPt8dpiYez7Iw6fwUhudd1ZcIf+tDSTUx3y+9K1Ieq6nKrRjE2a9BZB2Yj
P6NbzhwLw4uxDVtg8luNgwjTh/aJJ6LaHoLecE63zemMb7pOMH12upmMCydJUQ1Y+CFTsYJEK3n4
lyan5PyiH6K7wuyL5wIkhzuqh/ymPAF3GHaWOz2rX5mnqoU3im8N4QGJFdSZTp85mdxleieaNJiF
qxKjN3YrZumcyF1FOetkjZSoH9sz5nKjbcn6VkEQIEpf1qEVUq6aUTf/1dH6wPe/ZPWDD3+f72L2
Qyon/03BhIyA03Shyf/AtYWOqt34mBIDdycqIMrsrj10fcbFaJvGYfxPIkt57FaKwq7r7sgsHIp1
v2LB6qjJ4e1I6gSDElIu1kkhKUEmObDk0TNmwdLkvSiFW5tu6AdUjSKj6FZamQaqKR/GagpXiYLR
tUab+uZxVDClKcY1z8z5GEFTsV5tfp7sS5FlB71I7mK952IZjU3PzQNYa7U3nmqnDsjYIpTHeAP3
N9ZCcFI89AHqJGXfvFGcUOYFwn2wpLxng3CfaLK+1OFMYD6NLO0GrErpRFYqZzXuvkZWak9WSGfX
lveZyhz3KDiR8Er5nL/cAcNutRGuxu4Bx4zVLeuGf7vC4SRZf0QQwiYifOR7ARxanWVQEtcecUPN
F1q0oXdUTLwCvlo+UVfA2yOnIYdX2hjwgjmNsQa8ZhCUZ+1bjeKy7zo32rNZfdM37qmUL+e+bsue
TkUehMUCj7VFfGEJwFiRz7xkLj8hh6IP6ZqKL4IDZLlXfORUqac2lBIerpUW1PXyYp3R4p5Tolrf
7x7m+BfdCXz04wYH8Gy1qp4Ipjh5DmD2O9lUC0ZSD3DfJm8YisNFk1YLWbGje4ZrW6P9O53TeLiq
T04izBlwKRPISYxUOF7aBuN9EOuunaCFXa5Qf+gQnL3J+0tLRCxu0GudMIXGpTGR0eeGyq0x750S
SEQPhT2y45cX0kEKoT8IP90mNu/Xo0Q9ojOya9Ck5OpW3oaG9jW0DOQhzZ8WPfBObx2c3MqttMEF
7Oi6JZ/VNXQxqz4wLRSJ3bUu0Z6F7wfwBdOnm26b8PO9OeButcxnk20u0ELVDZ+cjxIDBr++FLQg
xpRJusL1HtreG+fzDlzsUNPLk4FxfLXtDQdfkSGi3Enqm52QGCSACnR0l8inKs2RJyub4J77mUFL
FxzJKa2XXvGvJk5ptzfPTPJXFmvi207g/VGPe6s84iQi88/V+zGExaWpJ5QxqwrBhnlCHD3ejRmY
TcrEzh15ALmLP3/7DjUfQXGvh7ssn5/UZElw88dJ17ihY/mXzVtI0PW4J9e2krR0V+z++YunwQ/o
JxsQwFyr2orzXr754cN8ROPDOzASJHS2m5G+GabgoLogYvL4XmltrEYjUJjRd7ytTTAjDKd43YFf
GQnUOFgMK1Ej/qCyYm5e1Is2roCwIUlGgw1EZqTP+JHPbNlIrZ4jPogMiag1B2j0gWALOQijtcMN
Hrcg7xwFKT653N+eYYMnwkazNv99xHu1ojZj0aimDSW5n8tTWrmmWX94+R15iL7z0HcBe23POqSq
EXmMrGg+zk+FH2zUH+bVrffLL/JKEc9yYRFQarg759X3dPZmFyOrmuxL/VYTw5Kre77EdEIo4l/m
ZwvLO5z/BY3RNao37iIyLi8dGXAe5FwWo5hEenQbVCvppgFa5G7H2eggev49Ls1NbLQWj0rigY8d
wURHnoMIlYIW1hEQiwHinboBKrkZXsq9bm2IcuD35wI9r+6ZH8p1Vp7iAKZNLs7Ev+Jhl00BcnZl
09GhceADWncIpVR91e2GESdFER7JU/eSz0h53FSMzjlgAXyBxGpS6/EHLxRDFLCNWMDLl5myKWj0
MNFMAmTkeD51kcieIcMzGvdwskVF+Ta5EONQ7ETakZtjKjLoWMKrddnHuyvJaCFqunLudGjDUKuu
MEAVFXFzRUHendn7DZFgO1Oj6HvFp/+9wBAJ+ObNQhhEDDEDPNz0GVdlJHFlBWRsdNVSViKxzQbn
Kb6fiDyETO8HkPwtrI8aMzoLPpF1NHPRKOtAihW/P1uhwrubupt5fS2diiRoS8jG7tVa4getUIJh
cKJ4m+X4eCUqMJDwV+2pqLy1/UHBpSsO1fID1eQqYRqLu4UZQmXIyOjMUfBYJ0TOViu0yLVAQq+r
MQjckO7W3UxJXN+mXeE5QvrBkm45NvKTn1SCYJngwPmHk1vfmLeLhV6j/cyT5WOjBsMuBHfVplm/
x3Lx2aiYHfSJaD8LZvPgZZBHxVPFX9pM+eNgn/LrK6fJDcFZICU6WI/0VdV33JPrgQW74BooHyPj
supL41p/ZaAgzEgq0BYO8AOZB/5NkQiOEidJZ/e775oGZigaF4pGeCBYecGH0RCIdLpDZv0LPkyh
g0MJ9vnnM05YQJxKr8hd5ytIMt5LBA7AHUR0lOMWCktUAIpKQuIOL1DZxf488CQGjLyXPju8jCNq
jOuUCFBs48auk3D7PKJ08hguMI+Gja9wxXG65w2U6sKpiiHeArsUDp9mUpZ21T4qZNV+U+tX3Ix2
AJwEyY8VwDO21HqieKEH9fDkTnpRgPqCX0EF9VXnRBE2qXISJX6oh+UKy93H1wLL9qcDET07uGXV
CCxjFm+He0fSrRhpwUKT33Ypp9Bj5JT88th27uKrpJASgNvmh8/MWSPSZUosTPZ309FUwhYMci60
hvzeB8dHLLq2AwXsZgShW2dpxPteQKqnWn/7TxuXvol8bC4t4iY8JFl4ZKFDIIf9IlnmGhReEy9P
ZVnu/uKhceqvM/AUJTfWOCPJHvOEPonqU3i8X60aS5A+RpZM9zyoxhQBbiVTLFYZrCnD3UUAKmQ3
zoHgCVTl58YosYq8WdBmc7r8sVIJ2wmIMA678+3mnee8SULr4680b1tqMr0xv4s9ivgbyLwMBVoY
yl2d4vCGP5hrbVsrKXccgot/dVDKuy64On3jlu3bkFiQR4MRQE69A0bosweWM6WwVqOTV4kDTMRt
9xKCEbzOBKsUK6zOHbGKhLE5attKRzwq5uaCt3Uga/1hF4aQ2FGTlAV8ug1Gf2YoX7RC+HR5Zw9T
ugBdPoRLT08Owm6pAsiXb2m/VINJJV8hAusosh0uesIn/BYO+cd71lP2oULkuyn23KtHS92PZCDG
zeKf3xJ1BDym+swwhckqJwO4rMIDi3LCftdH+8ZO14d6eQ6Ozg8Vz/a1jLauIeRbvVDu7fFiI/sa
zpiToEb4wrnboegxnhH/ZX85ABg4dwjZKRxk2ULPGD6n7GdGp+We69/9fHs5Q0KzZuFAvDG6ke3g
CVvoN/M1kWYJBE0bfR2BlwDzH+4mOWHhBg3b6CbxcaKnx42Fb+aJTJm8QiY8DpjqQ0LuihMdn/9Z
WJxCmdYNMoIv5cs9ETcs1/lS5hTHcflGW43NsZL08qbklO9VnUNuVANBjM/EsGruyHgZnUdvOZkR
1NVotCnQsDfJBzBeAPLYDqUBjsRFwNfacGtUYGYN5L+O49x8WnXSWaFmBObktYZK8b+Dlgq+1Oc3
WhvSJol7fLpiH3LXDE+UiYSNMQFt1J93GHlB3ycbOemvlic82WG69Lki1Min42EAOUu6iKtbc0mL
N5bdkBj7NnnFipw9w582p8O22PJg9sv9rIkE7zaqI3+UnPas5CfIy2bKYTXQ7t+6W8TQttrv8xcu
obfbnw/8nJU0TtHMxSykKp8fe9ekw2W/vy+24Uq/MRMl+0pQSiHW/CpZmTAinw0ABOeJm9Tgy4+L
m/7vUrPfN7076mCc2/OoOHja/Z4jimNEpCr6c8oWMCc/rgvzlxLKP3AirThVzqW+Wksol2m1sXKp
mqsOVuAIfwJ2Z273E1x1T9+crFjcYgZRbi7C92/lVWbQ6aanB4FKSct2NuzqVSWYUe//RdeCvQC8
5N4UdfbLBmoJ8z/GznNPhMiyXeItV+rtRiXe6bMxAtqLxN0DpLwAW0Y3brcgumlB4hu+JNga0/W7
28DxOTehndrDK3ClKWv6IfceyyfzNtnOnE7h+hv1b/mZUk/nw0FwaRfyVtTGwTcInWfplwvAhprL
PUX1N7uEyEkDRCfrFKBPS0k8J+sgmjOjNH6BY3KOEqjRTvNCGo6nUcOWkxBtuHIVPPleNLoLg2CJ
vGfz/Mtt3Gt5ZrY/aGuhbFOWnwJoguG6uKlEr1b0GlBot9Yr3In55pUaqemcoCO3TPAit8INC2/c
nTKjCxByCzHnygXEYqWQLLRqWBxoiGvJ7ex97tTlQtYtTL+QJXLlZUVfqIaNbBzXs22ZjdAbgT5u
w6uRdbLcSikc40H4xdCSNyASSKYxOu+wD9eo8ACFWpAGfjTACC/0ffE3EUt1Hbd4SJsg8g/RFnnT
VAfod5xhMvbtql6vmp8uFsVtvUg6Z4yrJEsuvSa4P7liU0dKTaN+tW4yrCNdr8iJMq4DSt6GRpyo
d0RGYhS1nX3GeDQ1SLQNVQSp68AfnjLKq9V308yF+YKUxHBk1BNs4IWfG27gp6lor0kmzMTDRrS6
xtFbg2G6cVqLKTsb6EonET7cNRTeUKO0wwj1zrofRX9XTXW/wZ4kwIBYY3x/2KzGl0pVBbd13Pie
o9YETz4NdrRghUD6iIVLGY5fvkDuPDxBXxm/O/b/5Wh+6oEZQwfbM8IN1npzEQXB7yd5Pdoe57eK
XJP2XmvVJUElXn9tOnNcMX84kUs3mxQ7+pOpXd9/Pkltycacx2XoGcENFcGZLe0q1EaIi8NQy/9G
Flk9CLxkBC5xVuGEceCz0i0e/t1V3Au+yDsgPUH1wkWBG/I78Z389+XoFyclgk/New3fKNkCkNEE
T+kLhkZ2D9JpAZsevydx3szlEs4nrMYHqAoPhwECSwad+Z/OpV+x37oZcLdyJhXOSQGLMSXFesI2
ZIYTIP9+fKkOFlqvrpuVQoz/D0B1fZejxEh24GB3xTucTOdSOfXFPe6GMLIad2tkBxDrU0hJXmHT
cAhmCKj10de8LPJkXo/gu+A5U9UP4EirUppiCxv9TPaSTg8cAT6PMOWzpLP2uT2QMZScxmX3Fe2+
sOeHc4KNhJGKhYAdn0NmsziKbDgI6DGLQKYGoMvh0hs4ysWsZV0/LIFxyt1d6vsjeNHX/Yp1ElhD
zXM2+M78Wsg55mStVjQzfSxRmri+9xM0gOERpStlw3AFRHNjuW+s+gl6bjo52KVf3J2i7WatW9PA
N/CQeh+UZDqT4QFl36B2VzSuoG/kYTNNyAx4T4o8BgHLZ6fkVC+DaAruOEkNgqgpYYqMSwg0yM4Z
ldu0p8f3ewPzh7XMk13yE6cUyUkCDbimM6gY3OIth3UBIYrb1lsh7ZQHutIZgWc5JOT+vLfW/CbR
4kusYQfbfCrEAtKMqC5gFiqvfIflMVC5eQZrLnpPvmUmX4OEx3GqBynkwc+0ToHuWkokAvZudDE5
qZcoEHRuw2wziYMhWAlgX+MfxSx/qqRy9ItgG4QpqL9xC7zpyj3O6UjWcEZ7FrtmRvGjWrS3ywoG
+Z8vrNrndBBJslzcuPRVQfYkrDctpIjyDQ9pRM1cBqfX16m6cpTj92XRbxpQOkEeCyMsdOfMewLh
uZwzm4hTpULhp4B3JnkR10Ut8qwld3+CXV2nIz1eSb4X3YEiUZnvnB6N0bcMPUA2Q8Abp6e9P5f6
v5toGo4tEPE9jAX+lWdQkq732udbv//NipbgBDpp+4r67iHGKmwpLX/cbydjwjOe/RC8W66+Wgk4
KnLqyjEAy+ytAOpdGB2HRwUwyRRWsucNH9Z/qtzow1QYkUGNGGfykfzsc29QriclYpSxV/3izUy8
tJEGaX/125Qnm33zy40QcHuRIL656wUP370v/iQTpXX63W7gAnzG3jMqoMDgoeZOejQhvvkhBRpw
iF4SC1u2fKoNdyf0RHa0EfTAaauEljGBNQnn2qva4k8ehF2yJOZJAp4HNp9NqaDOHgzObNrEC6bW
Z9BKvG9Mzxs+ml/4CYz9XlgSAU8QVGerXw1ldabGGll/+3aZsmmhypOzrYLNrltet6VRwvU0SuTz
tgKJ8BLQQlPU0PSueNJTgLFz0qLQw98wMuIFY1l+4R4dpl85xevMWEaNJ3kCOhHF/fLl5HOdqxBX
z5k8FpY1qJqRGSAR67Qs6Cf8YTp7yrG36vkMagmaC3SBf4UrCrb1Lg3AA2O0MGv6TjVSSEyDccHK
eB7I2RhoNcoy8M+I2z9PrxT482m2BwAXE+WVkWjQSo5Z2i4w4FRhndIhs0BmtlkC3Qal31J1r+aW
sqIFfJdjRr735jKtmBDXEhiZret/+anSZH6x3GBDy1ul1QaQNbX2VazbYnOpweJ4hGoYQ1QtcKze
2QeEACkW7n1hGEhp2w50/6V1hn0zQ6aBVsUNSuMlqmgoBz2A6DD8T7FUUckKCAkFukdkkXPNEtMh
DCWu2zP3yUlSABAGd2AWTXFhVKKOi2981ZgLkSg5KMqLXUCwBFwoC3fzdy5DZ/ouiok73ipYTdsW
NtIAxuUNQwbNf8k4LP0uiimYLs/pshMitDHeye708DPBKPM3RKNUN6Rk23VTC5CZTK3DpevbVohF
RmaSJMpxUQlmY0Bx/CE65ZxjQ4K8b3opIM8VExUUM50Y4WnzZpJSyuNILkGSLMX2tu9bMfjfKzoe
/XiE1iW4TxOW/wNdSDCKgl/xCSzA9fMF7lt2y97H7I/Mtl99iz+6w62W62fcSlIbR9iwnM4vKJQd
MJjtSDgmGIShI8aAANkQY9euDJUFOrIMImQR58Fh+ppYgF7AsjyIu+kWDRArVIZt1wZOKfJGI/r4
XtSl6W+Y4cMqqJjJPfH5X54FG2HtWpz3gcDYRtLPh4IruDzfiM76ZGutG+jvvrWeHyOHFQEeUogE
oBygrTuLBLz2/aPzNqmEStIWD9ARuSkRHca+EC1+jPy8rkscb+Y5xa3Zk/nywI6/ogtV3Loruetf
br7PTGSVuR4/iKcvL0idpAHDY8FWIP9FAW4WbvRdUgWX+cxjMI98tpvWpaxzslW9Z+u3X8BUoUPQ
r1BRbkZHLiLbMh84USk1aLnD/qaprR+g0q2nSjbTFrD7QGo8sh0pmQ9jkNoJ72vW6JIToKSVew7j
9P2Un8UWO4F7uzu9z1hoU+bvjFKSPd4J0Kl7+zyCRBWLtaEJYwZMTXJsXoEkqm5U/kCXoEsf7Ybz
+RyQhjbQZ6bBto+4K8z8UsRFzcXPat012nyQo4PpCFI6u8EBTuVwtdofL2lekMSndVxZItnKa9mq
HwV4zkGz50wDicXho/ICdGcNW6TzolZIBki9jLMv+ABFbNZiUyPWIJ1eDzAD9IeBBwaViwQoEO9P
qXOT/D6i9TwLi4/fYjecqUXOT16OGsX5jKtwsUgmRR5nx7TPK9R3mpFJ3HRgddceeQUtknfEgyp6
f4Y0lLZBoncnAyGL7uLW3KQvgqtqnaY1ZHoUb49BR/nDP5my+iyL2QKp4Ofiuu/dHoF0iDXFN9M9
0N/8RJv3R3V8OeF6XG5JiQQTxFAyucN2QaBwW5FSuz/kNq0DgCuP4d+AYZdqR1ov1zvjk1sin7pU
73cD0TSxdOzXUFnb4rV+yyMMmwGROtoAzEGSC5noOJ5nJ11fab3M1JrHNucRauP+7aeEaMslMDZL
VRmyl7v1/GKmKIYpCpAN0ladDiQGDclYTWrP1NjzaGm3Xy1jH1rkeRoS0Bc37rmxMI3u/FDrskeC
kfw60Hz0IVcxhmJwcEIFRtSmRFAfU6l5CR15hbU5Aq6V4Yx2ORlvUH9IwiVkAzEog0W9NAE0Kt7S
U39OlERtgJDowkBtZLW51GGhX+bEB4qrZMqCoWWKPkHALjiTzCH5yXWA3tNUGKUmcXSrU1LaQgGJ
teWmV/mX6lUrtIZo1xyy/TRg1gRtWfm8IuzSW3GKTVLMYwacpMhmGSnx2uSZFrFYoG2t9hv/mL4x
a7iOyVQ/sb7TgspPTI0hCkibiJuIq1IfhayYsGjLu0QMW6qikAlgkz5S5mjZSibCXkzGVEWtfjEk
GpZlONQH76JLdkgnJgsbgQ1akqSRoh11vzAJrLiDSnHAi9q1mGvFZr8WqgkmCplZ2tCQz73ZNZel
OTuiuGfAd1R4ixTwLLfRoazgEB3OUEEkXAqWJ9sMnzmAN8Hrbn1qtQs9KKgUZmo5Y5kWwik/I7FU
kDW7LmCT27NCgwarKS20T9JgFEOl94b7RMP1lhRseDh/134M/u4di0HDhrhlWpbqTWYYtbtYXICa
eTGaVLfL4a4KQjOB9XkILpfiZJwmjLG/G+PN9lzjNH3qCMiQUNW8qhnwHbYaNQo9Aajq7OM31f9G
e1hNvUt4AtlQMG1WNNFl86J6eTB66MrkC7e8WYySuCFygokk/wUl6tSpYJMrWpMoMvElJx8q3yl0
yKLR/GG8BZMT7VibtwsusOajLxupcmCUVBViKiJh1+jOgzym0JhtCa9/JpUvDOcZ2LcjHhzr+Ho5
GPM2AFc0BfkGrwlPEaL9950uSDzoexE/uZb4VUSJoUvqWaY7q3AvpgivTeBrideYet5CqQ6CrV2r
HA15XVuefQ9LaBnosGIVFlBkSoWx4PKgEMkqu833gIEFgsPt9lKlCYdEzNy9cnDHEQe1FyC4Cv4U
lT4BoP6nxm+rbaN80cvqGlm068mMS9dPW2BWfwBDJ03JY7alhTdGT+wfujMDlrOSqCLrBOQ4tABF
JxHzr5gyw1gfHvsac8ZtyI3z2UKm70GIHspVkZXfFq4ATOzNUHjBRU074gBzPw5kaBKXt433V30Z
v807ZczZyo10xPUoT53byQDBlnfPY6ErTw7tRiZBHZjU4RLtIW/vc0qSDWLY4QeCLRqItFZwOQmF
fllSQaoZQSA5txVKDz1Fy2azBFzTfJCuM2k25WFJ6n0tXl+M6RJh/UxtnTCGROikk6L4s1oEi91b
KSuBZHzFwmBdsQ61I6AJWAwJmNnQgekcmIb63sXNXP8COzBbKOnppbz6mZ9ctTIPgV+CptHvEj0W
SeJQudPflmUZt5na2cap/RHyChUZe4uveLX++7GsVk/2Gvr1xhkARblp5ziaUFCDyfjhgr8RucHR
EPM0bbOTe9u0urAewL6kovBu7tT9Qlxsh3vJ2XsXwhOmCTade4ytr+bax0ZPtoQqR2ym5p1bjF5U
Fe3G0qKvM79hauRDC0dP8j1tCgJW5bQxOIYsZg1TbGTzrpHh8la7+zyEkTT3YMRD0OOsLr6/ltjH
Ya9J+xyUXw2z11SxGcwG2PqMqBZhUQBByLad3lO5v9fYfHnJ2pWtJztUmwIme+U3b91/+twfVftG
KnL3JzyAF7t7yYRCd/aJawIbAfsWe3zwxPMqITeUPqY6C1pCf9wi9xGkqhV/98+JlwBJnmZpU1RF
+AHxBorUfpUNHr17DDCo+s1io/Gj+Omouu7zdvSaQzlt8hb6WyZk3mIqxzqhH6w8Uy6Ib2kffSGG
0TvpWpql+XbXD6fnTz2DfsdbV6ik49hqDxFCZ6pj/E6EIU9X0ITeJ7H/b9QKls6+1vkBNxF2p2Zk
eeEIPEqDbZ0lHM0njYvohDNNAjdUsHcgKp7S8id9BeX0s3buDAGy0Zs2ipGbTeudID43i4NiPAaI
pGO1j1sKBUL47x1cveCGlWgsmIhz8sG8tq947q+UauEQcqH4XV4flLRIve59+TzZVY8zEPnGa7+l
P7X0gj0zI3IvXKfGDqIYkgKcUoZCZI62VtCydmV0OBR/XFAUKQzZNADPgf1ZuyLEQSHvUy5HTKJz
VxoCbIG00smoe/Dl+LrZ5Fib/AT+BvyrGga8B3I95xM5MDWx8xVTGYDsRuCcIegsKNsQaOBiL+Tl
A+fz2eHDKAe8YqgCu/kKeEYP/O98eKuwpFGFVi2rV+94gmLPEi9u1b7OhjqKjj5H6mBlAOdJlQpi
lpM4iph9OWyps+HN3MvO9PTnSVE8Gj0322ATRkT1T+lwXgw/R5XRKOidqAlOi5PaED2jBYou7A6H
blVnUcrDUHJJ250zN2okSJjqNYUxHz7RlAANpjusEgShW0O3XkbRSMEpwGFGiNz51LKWSKbE597n
gvwUsc22eJLcscxMTa5wTjrRtpn8NULoq3ikQOEOtwzxLLAYSaA6NgHV3bA4IAOFUYkxVu+dtAY2
d6o/vvYYBJxnkZoC6B9l2nYF9sIdxZDneA6705h3VpRbUfKPLk8grh9VUHUYncnpNXqwqBTDVxmJ
wBty5DvlORPqbQOpO5GsM6x4WhGXN76tXOXrIq6yEh3yISktFBbGOiMQ4s7yDMqfoHf6B1p/am8M
SEqyuzBYhvvvCsId5QvixXBKND/Yt+eyoYX3Cuz4GQcC+XU0RUHIL3DCHvt6N6PdqKiKo8/dCXyI
39HHHmi8uCnv+ks0rbUKciTCBus/qX11o9bbCCzA1eUNig5BjJBR+QhHPP58/c04L3lmIrMjoEiX
zaMgXcZL0BM+9bZbwrkSb21H4F3okXW70lZmE0U4ZEF+2gSQITOU6x9ySyvpPnL7HnCE/TKzm0Yo
6YRpGbHuMb23b0cY4DSRrRaGxspuZOtgO4UFjWJPHEzfdkVb70o6qmixyzXxu4XH3ZS6OsUezZEI
USunZayfkeJVi5QGSdg7uBn2Q4A26YZRrWkYnIKiKvYMS8H3QN0CRoEdoeBoeFuubMzWqD0vakeQ
9t3IIor/V0zhqXapbfIDOWNsToQWStoJiwdNjqLHmGnRDFmbYoG5YZ4JVA7IwBkgIcSGLf/8K2Tw
MY+2IgY88DWlUl3ef7yQX1oUhpHMRDbmvKvzzOEu0+CyxJdAh80K45cr69tNj7FAvtbsKDi1gNog
P7dbJhwtUD0ZWWDF+aZ+uw2sEYGI1QR5EtlagKys/H5k+srdKWI3x3bdUVYeP7SPfT7inwKaY3X0
NY7aikBcAmvB3BCtRjV8AVIf6AE3mfutAdww79jCuEfUG9tYpIPO+SbvtV2wRjbQHg8QZsavH+5G
1qk9ymumBeBVurnkZ4ywYfDHK47MzJR7YHYQzIGe3VyyU4WZ4zf/wqI+ddpe+AgEp01lXLRUjT+3
b+JTagllzLZox15ePdZKmFr/stC2aOy6s8Q2hei4KTzZiCH8X1w/EqmgQEcSTd7Pecn9GYIIGmN3
3Ir/C/Izay5NuG5haKy1khZQPeH5WJwxolJQxuobhQ5Ff4rValagPuQ5HLYA8WKO60oR4NyN/x7B
xoNHX5Ff/uuFYM39Q/yRUxM/OUvFTi7tgW9Zj5L+1F+YU48XVvCzIbZI37zTh78KNetXH66tnwu9
b30bRRxkDl6PZN/HFLl8Qt7YyUbNKVsLkRE6aFFj5vJ7XBS6xRBIOE28xx1zPOeL7Sxbvq4bIWAt
xb47VuI3ce4XNgSV6xHijIdb9saXs4u7jk213vwFFYLRi+0hhL+9gdW4BGFH5e0bKn5t1xIY34vv
gmpjOKtiuPwa23URQBhic4HAkmWlun5/Q27aX0Nk0zJqyjhKL3b8jr/o8UB2c4LGJ39iozM5a5uD
lickMJVuW+sFpVaQTA6ptBR/QEqf6JBgoMsMEGgZ479iZ/Ppe5M2y90D/+eHFh2//rBI4uCdgrqe
uFXz3mni0gW+5TIvCQP//UD+nfW+UzlW0XhxzBo0D5wkzFOjLqKREb020x1EDN42EgkSHhnoua5M
P/DoUsr52EU2aa7xDKwuRZbQgy0JbnDGQXAe10j6PkFHzI/N6cMTvsp7JxvkSO/jpNLYWC2giEux
BRpiSJf/gblWxpMiT0fdagUZ+RQ2O9qKDoZbtTuDxLDOmaXpfnnELyNYNnnqBrC8ZBvSDGTsbTuH
VqJewBQo75/seWHsvlvH9jhsRJYuBHCrHryqhoO6nagvbMrVVnBfuL6KpC3BPUY60CxPwgvIjkjT
baCKcV1KJTMLejPpq7tIbnbbxJ4+nXhq96D8LGE+Sij4IM22e8NsIthkf0evQYm/PIKwDxlLiWAQ
X760ja6EoW49iwVd2NldOKHqydotEluTKW+gETj3zOMB41CMW3V6nlL9Ru/PEGIxrunDwWgSsu46
DfPPmTfZWDQJnpp5NWbaAQJCa2CeXoE8w/ofoAexmN3qGSLtwQkQAQ/LyrEkZMiRlRKH2Z/A6Gi3
xZNE01RY5U9xqvYAXdKgou1zHJcUiD1QnkJtn6N/BZKXN5jZabnCAHupMlTczRSyBFOMkkFlKikW
wbWgT/TtobyiU5Z61IyINB2BHWGd64OAE8DSC/i1489pnW8shrbbllSPJ1wwODaSs49ajaVvbtSd
s1cUZEjfdEUs981/KL4W3ffipHand2iJEs48xfu7cJd7MdLD8LpxNozFtHz0vfoPNQfQ2OCIRWNp
oc8DOBOBTMfHMjyuZ0trUUdPINopF/aMSib95v1J1QphUZtdoHagx4yBZTO7OqNTqxKk+r0uJFvU
jiLMGItR8f+C+Kcc6qzO4XKl79mQSelBZH+5F5T3seXYc1h+HkTTDPibj09sWwQ5bhKY+PZuDbKk
Jmh4LQadpAtXLOlCVilo5Zkc41AwCoRBdCfljJw538Vt8fSwlFnZU1CMFHSw7VC3wkT1Q9nnS+Gs
uE4SDe8mqW60QBzu/tGxJFTzwz7cMvCjDoh/9goKjiH8jDvWfCBv8wlOKc1/H6g/70tk0PNEfreH
uO5mImKylFNX6OXHZlE7Dv5oS0apYcQYcNNrABzYfju4Dj41qieNN7Sk1fk0I0FiHXAMgqnjeK6r
Ac+V7nronDOsKPjsjlhf2kgDb4mRigWmokvCtndgeQ+waPkC2+gPXwyQtA/iRqgzSZDgHdC6tZG/
hFRWOFRyBAYKjre1jv2oW9yubBMOviQVaLmxDsw3F+wvR5psx+4mLhqZ0uIFgYoC0RhD53omzDKT
d/he6mgeAG1JCBdyAnOExpyKArqdd3miOoGkVs18d+N92+oP7yC1hct3nUjWrX81EfMOVa8ssQ3a
9EErI4smIEAlfDGzyRRloIcv/zeXZiMphD9unsj3SD4+L7tfyI+FyPLrBgbRObwgkkCYXf/pZTrZ
m11eAx/Cz3SZ11lr0GyH8D2tLKPPbvJUtg9UHzm5wVuhNp+NrBYbNRYdLp2Ey+jNDlPesHqYeofo
vOuk4/KNbPT8POPcgIphBZLZQJ+kVHVGOgfLxOB1ZH+v39Q5TunNXYRLnQSSsw5jvXNPBLHSb8Ax
k/fyEXGHBT6lQYgFK+Ns1VAVDpaazxhOaQVYBWnGcu/WZ1eXPUrV2vi6kjfuOASGYkto942/wImy
vFcb6pCrPw1HWDCzYshDfOikjz7QFMKmgU3Bch80vBMp2omr8EhUCkgBoNUvq6o5zRjwbnqHz7tf
G8dhwo/zXdy89ZA51H04uPHBfoLLK72ouPU2nIl6luS0z2ci+fhfdGLVq+uJp9CniFM9JxI460lF
aWuucH2JNzuWzMntSrVkCMOcSTM7TFV8Qkhjf/PPa8Hgj1pmFjkhyFPoNyqzsd7gzp2Ch426faWm
lamq/qPXhmILoxYJuhxD5JHIfJE5V9X8CrP3vYiRF1PsMyepGcO46wjKcJSEeT0NtEE7Bzfi1vwI
ieEcUoe7zCQEG6sD2fYRnhsw3GbDzsCWXjYY9Guhb0wY3z3jKjOsCBUlBEWZ7uxvL5g+C+iA+esz
thkvXYWyAYQvEPwtPNAvttrRsdu4Pdzjd7YrqDuAtuN7w4iske4V+wmIHECrIxIPuVL5IhkSrbbL
YWo4yrK4bb23x1bZdfJNhBGvLKpwZVwqAZGtySYEl9PKgmeDDB6K/Iil9l4UpyozEJk6NfDhlVvz
ae4IkRgY/GOqlhWiLNAVO8O9SZ//q1hzA8irunQAJzjGz61mcUmm/tUCAgS13kpK1IKHN6unuefr
qgGSjqc6m8I3gjFAW638wb9ZrETmFKycQn+36Z3/WJpZceJqbRZf/vqKvSoll2aLpfU+k/XSIEK1
QxTqnUd55nFvwSwHEjro7yJrdr2hFwM+9BttyC+rOxf5tayXtiWiHadGhIW7qVZnn5bRer2W1pBQ
DCK284GhfSNoFezNAJpdcTGRZk/6DoJ7JQrT/4u1ktZW0bxDN8I7kQ+f+Q+7yBhlcPvLczuhuPV7
FqiH6t7C/30sZz+d80q6gw1+kmQDP/TpKFUG3exjf8fQuzheGcnd7qak0rNVhbRSKzmDfIAvVy4I
1N2nRQ/G9D01mPHRNPr/JgeOVdpWCNhNiobar8Q9AuDTHSak8ZikJIRdARyxi0XAyvtl09AJtAtL
Ak3VyXqcIvPDptB+MujxXxR3HLtGn2MiTjSEm+M7qF6PVuR6Qbd/1SeV10sFsUaroCZKY8+Yi1ry
kthAhWJkdb6VY/27ZAEUfG9V1A4tPJ/WmkizndbhUw8wW43F10kHj1HMbAAeOElYebXD+xs6Dowb
Nau2l5XnrmJHp/4qOw1vvhFce353j2NTpfQ9Bf7H/clWwFg67lloDQSv6hvJQru352L4Np/IDSKQ
XBaUQC3sdPfvHsI3WS2iys+a+/mDQaJZy8n6EIa7IRtPSh+r2z/S7vAoJfn29P4oRcum9trXMfKx
Gm2RIZHZFJvUyfgUHokkHwX2B+aSF42hnY24yh7a1vJcHsWcXK/EBbmCxUgCBozj8Ldb569gMaHU
ErL+v6hQTU/uRQFq/ojtZR9fExv2OZDPXw3tokUvKbbNiyFJ/uN71iyTqAosWagFmigOXeGoXKTR
s2JW066w26BZ/Ifd8cryFqJ7g3+i2cRJNAWOR06CxXDUNokxBJyUn7pql9XVoF9eW3w2aTB+S1DA
Vqb8OZxcrj3jbBbkHEjNzv9GYloMhtT2B7gCmCK0UEDe/OhIj7sz7xRr0khzZ2sZDX/FNC+BM4GD
dRBDfJD0wEAyK7togJzCw1LX93DRVWXlIu8hT98AfbdXtZpg9ry74Sk6bnkF6rgkNfWS2Jsk7vcH
Ru5FBPlXvKcjpKuyxBJIGsbxAvd+Mkqt2o4uZwcKQ6UoG6cPnGwRoBa3i4jpbktdyjgLvzXip/XN
ioRJwo3EGnVc9QWHRBNu7XvymwgepoPh6+kEt/USrKuewXS6jgO0Zlq8zZG4y+pa8Hx9UfvIo1uX
7X09KzWEdGOSRM9hD+4478Ih7KAsUneEU8MeHbUIsM3cGCnyqv8mjNH/7DfiirSx4L9OKcqMB5Wo
MOR9jMyDwjOPNJmEmkOcZzyGij1TDEj6KSCpkPDTIq2vJRCp5690ktysg7T93P3KS9kGret4Ps6z
WgdoE2nR1CfI788/u039OfiQyVyH96apSe3PPUqvWAybzY+ghL/l5JaRTfEZG/rRvVX8XQS0y6Am
0Mx6WB616M65QMNcpkALOKf68tZWcrDpk1jCkzlLx/57IhCL2xOIDRBBqTFr9kKWgsJjmmQvUmLJ
8L5G/p+552EhDIQYr1CFNVaV8sfxeMhBGUK0nA9maSBeHhdJy/XjHi5cSijggT1VzDovmBxj29NN
bcMzsloVBYzA9f+1O7YrrscpswYmMcUQMguP8enpX+8kOxU45r5dOzy58iAFC8bm+jCITVUzel1+
HICc6ozShJFiHopg5rCgdwHFKidJ9pQ+CVP5/dNMeNE8BUXCSNt8aHSR2ejM1pTQoWpH8ZNy9t9g
ls6avAUu73otixeGWFHf/gEyXMW0U3kCz1Gf8rFPiFgOLpUvZixV+sF5RrZBcq+d+soS1FMRMC0q
E5fCNl9rr5VInunGD1ptZv82bYtnX39QBm/MHWnpRsHie8RATUeLHZN330PF8D0DM/ucRObv0ORV
VTWNy4IHMx77cfCdGZ251llMZJa8s+Jj4gDJIZpSxT4VPIE/pUidi6hr9UiMpG35/lPJf8y3Mj4C
LQ3ChaKKAxz2ub05sUAHPi7iYJNkdFgK32Q7cTbt25EeYowXJsA449f0TNjCfm5lR/P84FJ1fy/j
nBW88UX33+EwJP5HQF49KCB29wPt9EMbTkow8b8Wx1TJMVrWvotaaGYiHNECzujA8c5r5O47/MqV
XFJRCC6mbrCc8itkZPUUFV0NS5p6rQX6Q8rCGUt6C0SB+0abZuMh8ixMa2rY0TzX+byKrg8kZ8Ow
TRaPilO379V/qET2b/WoKcT913+uiCA3lB4veGl9LcHVDv1qdxVSBSZek/gEtc4FrfQp9HxRXsXH
hHBNqY2uwt13cIDKlQL7d+BxZXyFrPPvqmI1pWPCQbsuyhrcMf+CyLHo0fVfhk/hjDlTDNrvyGKp
717YlxA6RWx0Rnf7IOhku0O14H/j9p2CJMB0x6I3BZswweaEi4cH3bpAce4C/5KHXQ0r1FRE5/1Z
7OSewMK/8QxMiV+6ZehgP/2qBX5q7QNtRybzdkH6Qq6NmJiy37HdnMOJy6gsZfIS7rpPpMqTFeL5
TzTt+CbG/bv6iF+4YSWiAP43p1g/503fP/q3VBO2B0+GOiyRoU67X8i3ZTJx4PEANgL+FQ1pm8Ua
HIb34BLLmIW9lEOBZHIKpANMicNLPurDgLqC9rIEsxenhEZ9nVW9qdE91MS0F4sgesV5pV7CLih9
G6DMZRnVWWojM7KU7bEaWwXYEl9KZ34wf0ywAYPMCUC2u1G0YZ16C1LmJYWcZNCrrxXxIQb9+OHb
EOOQfJi/DresWTQv3NGWZjqOgyFFdwfJowo4teS7zXCx6ItiERZ9Zs5HieR66PpgbMoEXp//GbvS
Jzs5BmxhUGSI+nZVNeOPm58hyKZjtPyyI/UVqsEqvHfKFlulNmInJ6bGHO42opw3DLWpDuuuINzw
eFsJGsCAiBAEtRa3B+DebVLyeVOPBTxwj8jLGLY4fPUih9TCpHCzQtCr8El3O3Wa5Pn9XbhWJc2z
zJqHpltFiRwym23qyCPoRRR4ORfeG/UuXFQ/v3+x8+BExgjnrHlEJMAHxaOgy1LRICDZ4e90FdJX
U1/ojjBdUzKK5Od6gQktW7ni26PVGm/t+Alw+JHuM0OnAnJEhA5LB3DVOKHCOlfSpxIAoE4g45+g
7t1Q/ouIHKxsXLPX4YrMuLLSoKat++DR6QUJ2w6QYFojLqZ7dcLiHXmCZ8y8XDnrX0BdEK6qd7Ji
z8yoHjQ+YgB+vqS4uyF+fkwe0WMS+M8H/NK+gT2tDGffxxrEDJXme0dxeJXwwxDft5UxjeZlCzIL
M9e+ZyisvF3I9YTn3SaCWnij5BOKIcHUl4KPJB2Xw2s7vRKiKORfb5DaAa2my6K2G7cjj8Xe0mSF
22QSwKYbKDt3XVLHC+WH2ybbjAuR2jwpBjjA9RQcdFfEwLGqgvlxAurDrxSvHn7/Jp8ESEuo2U2R
6q0aDHSywyPo7yeU4H0bRvNqqC6m2SoWHh2k25EhuXcZ9bTuWpcEPGiI27PFDnNwk2w9OBcX2gxl
rtoDG5srA5wqdQLVJy7q984GbcdQYaYLw9p40eVPzZz0G7eC71YSwClPbKUyFvXdpTSvAj8W1I61
Aasu9QKZRzKeknKPPTe/VCGmzZ67jGcOhUDFKRco1089LucmtyOJUTwLMWthKGZSZXxjCXBtuZoW
EBwSVI+jI+lhgBoZl2XifR6h3YQ8FHKcwP0I7otZ/UW+4vixgA9K0SMbga39BNHaMR+JNL/A2RW3
vGrygHA9q6eGRvAz6TcL1nHIkGbgPHJfCH+L+p6fD9bLZS8Wsmwuy5pvS88l/Kgf9t2VeR9P3+Gu
Ji+Ow4NcW2wuOMCYVvuSB+ffWtStwFlJx5xAhcIr7Y9DOyzjH0dRNs5prcLSKjPXF9x2zWCUmLzz
nj+WNgvQbFzN831+cC/qRSeOQGS6MTEmbRTGtBr7fah9XQfWiRxXpPIbJnqMK4KebJl5xf70jDGF
/nCMC/j7gHue7EmR2wOxTIvTGRXY+IHTIYIv9zgNkyZfoqBZFpA5CmALiQTT4LfYz/8ci41tM6uH
SlqUH8Ib/Zw7cvgepiPZu4cWBrEq61wPRkEiKVbLaQcH6sHpXz+PnEXpdWLD98veK7mXYkfCD03Z
2pDD3c/JG4TLNvLJ0d8DF+AEsJ0pm6yp5nAqPV7qYJS+rQ9kYdxBAuW996VsLKnemS5kwyIjimzZ
qCRz24mSP6Yhda4eGi+EBqohOnYSJBJAFNFEogQRpHuYXeFEh4/nssIusGMEpub2fzksffieBdi8
UPmeFMM/iK6jDsrO57EysQ7fGVYX2EWRHEbmcODJwvd85OfYkwGREq4f/eqav9rLhZ7Yuf4dvvpl
6VJwJjyuOzTJj8knrcbVAjkiVOHvRLpNcsKGQ/O4fyR81ZKAuyjs4uSGY10Ca2e0fq64vhlO99fR
OjAVKAlmhKbThxhBUrdeExch8LLp5v+bae3UsRadOJo58Zngy9hVcEhSFUZGMJPY4wgAgVg4pEvL
g/t2Bp+uGwrJOPPD0THkKfRMStayTdHInZlHFjGOpedm2himO5csfJlhxoUhVAa1mmBVn9sbDHc8
Bc6xY/ir/TqgHdKmkB50+jGHPY6rdJpyUwrDdHBLbfTo1rn878+hToESRIXIyfsK12Yvzc0oQN30
fc5WvhtwlfPkBqC1NtDkCWtnl1JtWY4CMaXgZZQMTjFt9PDtL0bVLRuel9uXX7okTPouBRR8di45
CC/h/gRKTX5WbTPZtGxbiQrWMXzxHz93Cw3hvLPi0BX0/YceWnBbWjczoToqmmXe3u2vb/ZOClCI
LOUfVf8nOb0PwU2B/3Mr9+VwKwZCI1OHK2PzQcH4iNLGtEci6rpEfR6U0drSuKLK4ObR0iR+VO52
wUKuzP5mT6o3B9Fv3TJoc20DUMkVUxhjHcW9H3Ca9mgh4wHhE7V9oa2//4WHucXKnXBNla3FnxT2
fMXFaIm/kTOgIiRvUqmUccPYmVSXdZGol/kRvyeeHZM6xx+zAKlDiBrBF0kuunYLh7zA3bZdd5Zv
HmeVZmk0shwUYAr7hppPiFRQ19moUnIS2jSHM0b0kQ6Uvfua/qlwW0SFhTqvaaogoNDzTbNxfF+o
e2S0SbumgFGIWhHUYF5OTf+DjMhbag0WcZ2CrKE4b7r6Wb5YwwmP0nwgV7cryEgwYGtgVjRcF2Vx
rlo+/0ChrJ/iORK0ud63k8NLoDYU9ZwRQIQ5Gaax0iK/7xxaHx2vc0m9COX90IkHBbw5DmM94OMG
yYEhxw5i5L2HJtvQhIj1K1r+bxwblmQIQkjBRK3BLriHMGk0aUiE6vxQtu2WBJvMfu3VhFdZ1X7Y
ig+Xh1KEdCjSKZ2CCLY3CpiAsZmt3QYAQyFkKz/9PNooILG+t70TL+9gWhuvWOk+naARSjvpzNMF
1LwWax3R06isq4RMiT9IXITR17XkNRs8r7DTiB3t0tY5CvVrMx7om5SFcjfhu7n+smWWwW0k0wMi
CxsdAEXX+2zRse+bPZ53hnNEu03aCJN1t+hSdwUeuCs3mMd89uP1DS1KWNwQCUIstYcQ6rCo2fI/
R/U4xqW8TdWHAIlFWExkwtOuAe/HfheKvon85Xc3uZ3Y+gcDglru8b7ZwvZo2KAheyPzSk1vtNFv
Kx+HGG4EqHkdZGZVg4EHK9Q3DJ/yg+CGVtKFdLueWsxtBVB+GKry08JmkcygmxGLsE/1BrfjxVPd
wx+aBuoa0QkvNpNUJwB3RSnDpYkQ+Q4dYiOTS7JfHCA5WhIgF5FujK4n/vVHdRa32EJ7sOjC1XZ/
N24HUJa/Rs1C5Wwx8ZuVmnwu5yJsVLqldN3fz6aeUGGcmP70tH7Dr0k0f48aWXHr9hoXWk93oWXd
wsoCKDJbj/M44ODQCpQsDQIHAwJdbhd7IcDMPR51LxvZWqbd48S3Zr7E7ado2CoIJxlLMOduMUmC
30GY3tRiVM8GO98+CGyIkyjBKANcnsM9/9JmQFIc5vKamE5REOjBcBuDdQM1JPS3RjiYuR+A9blt
pupX0vw3U+ahw/GUyUwIVAYSURmJUbcSMFDi1Sg1KgACnaesNLqcftLf3+usXhTIsFEYY3kpMlZ2
aPLLP5wJ5iqKTzgBlzU6/6gfzs/3nrWDnpUmOYHb9bqob9XMcrGHasDOJ6V7EaVaMT2rTIn6MVgX
iJOMna9pCjr3DOYIfmpk6kiH9cf6HlGmvqygIGDIXu84GavFGjB2P4+TX1uOoFpzrkk5RQ/JpPRC
rgy9nkYwbachDXtWxD6R4YRengCJioQ5aaRRTZ9CKKzW1Oi/bP93qCBUIZgNYc49pw6wqxnmAD47
MHEGt7yIbxZ7Ln0csuPDpm6B6jYiBR7yKWU8IqKO4/2h3ALoJmAnR71qlXStw6GwLERCXeGyFhs0
318iKjMFSjJzlFPESGQqUKjxO8HELFVWkcSmLSSE5L3KzA4EUecGAfpohZpwFDscBRMVRYXgfDFJ
A3HaklOItV9IuuWdvXfKwQS/KDQ28K+N59I0yDg4yL2QIs5qHnoj1t8FDjqN/EXyjW+zIZjC+nF0
wSJujpLxoCfRgNCismOASDU1l6kduQTJ60R2o8f885uF+o8Rcj8pAXUBxyaY1Qg7QPNl+KeR1lzI
4iE6teI+vGlnLkP0P1pXat2pFwLUD7bt4zoTUBInrau6qWXNZ6cBM5Y1ulFkHr9yAF//191nP68N
W2BeSBmGkXHfjlax2rfMFUHKYTyn297iwoNpjIv1C7FCMKdnb/jntrEVk0yF3ItMH1nQZlZ3w0s4
7C5n4+wrqfM5z49tMDdkcChF5KNv9HFqMoN4gV7X9DZghF0lRYjybSR+Ock6h/2s+UuvA+mqziv7
vlKSEdPpWOaLIGl0f0WKHgDpZzriGN8/qCEnbPyXo+h9uQvzkEyFq7jUq2+Q1Z/yGKy90cKw+mKX
c//vFX78ksEiY3mCkp52hlc3BcTkMGmIKEMTcw3SZ56kRDqpwzncuibl0XOIbW9JlwNwnSazTFUV
VecYEjrjm0b2flnM1iXW4jhmelkC3fjSob9yMaBHSJpuvzq6bxqtlMJy5H9BL88B7vClQSRvrvIy
CG/MKiuApK2iWnygHI165M4abeugfVsWYY9Br7NjM3MEzcvVXmC5CMgjHrA6EBTen/i6QSuRSqsU
mq6j85ajFAe6vNyTwm171jthr9yAK70tY4+K3QG5KQaRp4Bb8XxUS5aOBH0mOlLHW2FCDdUX1LHp
dpsOQ5lq90tFdA2PLsQdTxdl59LHlOx80ZsB0wDpPQtGh7wRUd5eG+Q/ZD33U2X4/SHpnfFKe2FC
a566kfJkxCcNr1lRr+YH2ZxW8hZv/35DE0IbAoAIUBqi012CQJ3lLhNr2EcyjrLl2sovETvrwRZT
RLJVpdY7j6WvIJnw5sL4M40FC4UuEN6xWwl2hZrREH/xDUkU4H9iQupr+8MqISbdqPI2fVg4vXsD
dnhMy1zjBc7QD5BnNunmNdZq7ItV34zDv3t+5zmZ48ku9ijq0e9WibFwkFXiCs+1ST48p5iy5cRL
yeNHLwsz9h9+OzAKzOCBmffJmNw6X9lI/C5rO9TY/KkBZiEhZ1D1dBb9/lGGb+D67j7bioiL2uo/
a3QtQWgBBeCSUiHROyMEUOiNA2TrJr1oX8ERW2X+Kd/6uacUELjEJFPNWT14W1Xj43PsByawZHYu
sPCm11Ku1QvijxAhGpRxs7BKhGB9pdKyJ4PmaahmiN66/4lcER1QQi1kA+X8YZybzrLk8LH8QcpH
v1AAveMURY2oQJZGaTiBFuHyPZXKkdo4EXZLpaRSCLTsx/+Xnu4IVWtPkQ61gWT1JL3vPl7Ss006
JAA+Xr6xb8xarf+5xIehRRHgcc5YehkyqvyniaC2aaY0IFQiemSYh56+HwpCRy+g8d9hgH6a1POC
Qsii76YGXTt7bQb9b9HPeKIwOA/3Mgda+Fz2gJTzMNiEOmoRjidnIHBkkRWDc2AdO/p/4c+8D6kJ
iO2DEA9oiyrKkWR60dlp8zNdJV5FEnXzX5r1gqNCLzu0EL0gQgz2P9iL92e/MGiUcc5SVeSZmHo+
fC02f/4k3+WGwb7cD/c57NgKHdbvkpVZlYO2dgcSsNSQPomLeWTxjZuH3XUBCs1MT+3l5lMGYfu5
LCUg2eDoqj32PAmh/8yBpxCZK09O9GDfUgFTX0ArIUTJEfQDTU4Kx0FV2mtM+mG6gJ3tj3Trjmi+
jHcmMDvpEmyg6Qytbr4d1y3Uu7s/p4dw0DVtm7ZFXne7x30PGI67/yqtfwM9MLANQgmqSj1YxZAe
aZ1CaRiTOf8RgUzOZAMP79RuJnRzeklEZkUIkY1jpA8SCS3WfUhB4n6ixLo93dLhPCMZO/ezKQeb
fTccYxxVj4G5AjVIq6g+G9xriYte09OcsJUzCWCGAZwYEwvaiXklsmsPP/FMJlmTj68ZIpalUsff
yoI9rlcKZA34IfZ1YZRNOCanLEXYWB+5kd8T9RxWlSBBFDfXoO7mCe5Hj5gYjV1/AQ0PjuSpFKmd
L9qCTYbBThysXJdPAn2f4v2AanAQRH0PFsH42d1J6hfhjNhhYTBedcjYxoRrrxtCbs6ukg5ftQOV
7yLTXyfM4S4JZl3DcWzmfv++zB8t/g9Mp/sSj7UDJc3Kt5RjhYg7yVccm+eGFB7Mjj4d6/WGdt+3
QBqsTVkpENt3HwzYJPFfTGfG+m/090NtLiq2eegw0dGmA1JlpO16RK7PFUabrKrfZF4Hwl74Tsxa
OxYu9BuaPrUAW25iPbNdqOAwe8ElWQTLEtMop8DBaReoArRcS7Cw+xTQH8ECUD5gqQBuTWNzS5zo
bNoqAZ9T3AtaECsOKO9WK1xPcCqCxARVnGwJUxACRbTh25HUeD5MFlprK0KvkNNJAYasd4NV7Dv7
4eJPyv/+FdKRv73qD7meNT3NytqoW3m06FrdOJQq2acbFxIngetoLepGW3d0HjcDlpNfplMTLQDD
zWhTswJmKJRoD0laWkpcj0pRw38ECamwkfCKJTD2RYWqUUgIO39yygS+7wfgMuHukZAanfT13y2A
TuvKA1NkVprQFzYks7X2G96eEE2DYuns8gRO9P8GGbAk/XKjBkK/87XN7EcypwBTz2NSWzrdrczm
VeRsNqZbh8ABCb9lS1ycU/HL93I51U9EpYOXW6TVDLEhIBqFUYctsbpLF76H+6xsquiYUp9BhWUI
oH+hDa25fL8tby/IAHKglxOmRoFTFU8Fjg4XPw6yl4pYlnWvrTd0gnxAiLgoSd7ezT+z/TGSyO5K
WBNsCPzrTrnVPwBKX2fXicxTtbuQqNB022myHDuOG2akUO6d0+NHm4Qbg09nT1SeTGat6OSneXPY
kGhsPX1XEVE0o8IVRLC/T5BRlCWxll+Bw1Vg/4mi+0HPZxMQefF2dvL5tgXo9ihcBK6YR1sRnFyN
polg1fpDZjbSsSGb1V+ETrhieBkh3UxrmC5dwqgq9d1I374P88qLeSh82iNLlGdlw8OzI68UC5mA
SosZ0Y7EjBJXaNlxU73ETtsjV7XR4Jbhc0QwIz5jImWLaXHRR30NlGBt/vfXBCCgXBbtcBMhKkfL
STztRR2gW/bMrWaT8lBFSY0EwN3fJvca5B2Z+5kgE+c9VYEMkaL9Ti/V2Y2LglPagrkGMc189U9B
8FvW1sK2aR0rByFOoQHX7G9KppdVbMSG5fkFLbOHnCinn9JiHOvaX0vtigXoagoqKE4oJXoafdBv
ZwZoVrFhGBE9WOi3nS+RfCOAUCTUupvTQlSkRbtbnE3KoZXhOuskvF5TOnUk5JpSHveoH+W+8nFE
AT4Hv0vkKziwCkUMhoQ4ShK8aUJlKUdGTH+zmTyXTl6YWzChF8prJ5z0eaQKGwFQl4I/SU8equcL
1rvJ2bK/puaDm0Amn6Ku3uF5KikyOvEQ3DhTfJVQza+cl/ZTkDJlzslT1ZkAi4mwNDP6vwpvFym7
Sfz7Qi9IG3MUohpY9PBXl4URnkFkLZlXY7rlXb4DHjf8sIT9rPSAFyq3XkxthXuF3I7ygJh5IC2o
R1+4mDON6YeVht9sYN449lfpN1gT6YmsZu49ryUCg7nE95pD4oYvGda84EsBvOXdZCmy2VN5OTsv
AQusxeTp2p0P5gSG607CLa/AWz4o+x6BgOVdk5DMCqkdd4eFV3K13/KXZG8rHGHgEIvVk52OvaYZ
Det8BnfpFjHt/LoiWPHity98TpTd4vVfnMFJKEFQkepOuEmXaUriOkIguO1HmN7L/qtrm0wVn6ST
eJnkEmG6czD0EO1bwAatzMVor7SVTp/XaNsxcAzcdz2sWUXJ4woQ1PgV//oc1gD4Y2w3S4chVkP7
H9awx/aKaZQfov7Hcr4faiIyfYkY4hUFNQm2QWAMP49cMaG+CviQttngl1/RYXU6mrRxE49UdLrs
jRyz+I0hpT7drlIH+/syi0HLu0z1bKJ+xC3lMx3WXFrvs69Mq3plaTr9mMugis/z2rXHYaNXaN4x
SatE5wMu0Dfh9C/x3SPeU35cZIEh+RFXPD6VN/5Yxr9iiU/sOiCL/kzDZC4SE1j7sUoOee/yTZub
KmmtETs8JQC1VgYorr9MHbI36pLhNt1MiNoijBMw1JmxS/g3bOhYAaba5fB4XTU6z7FFAxVSMwUv
s2Z7eR2PY3UcW9374rsY3h25dJAmHsMdbumhN3fCVVCENiwmAmoTCKL1R6wUcvQLjGgJWIUdm8Jz
NJ19qjIsgeS/lz7gElGEFq3R3dxPKnuKwq5DO00hlEAGMXxo+2/Dqb7kFfvM6ufi6aM8XqLDPT9v
5TkOqbFhtMwu+HSPeT6tgMzSOISPCTj4+JYxj/gnd0zwQ52w5cFEweSgBnB+rpuYSP+pgg5fVJdh
2bDV9Qxuw5EIFI8PWJztVqUMlSHQ3Q6DFxujG+VP7NPkyROvp3oVjqiGFOMbv3yEXKoJZyRJpoGI
G7EoOeN4m9S3J5lremNjTtFJNNFPF0+T68+7Ph1CdhdSSRD/KK5DKg/rnf+JLAz5WruKpw+hhdFP
pf9cYlFTd8v7kycAsuHRCBhTeCFhmn6m+3HR9lOtSBhu7R9Z0XOqwH9aa8v0GJXj/XVd3HOsCNw7
8/ipU2zZKGIllONkWXTBOgAZ7qm4J9U4OKCNp6BJq6d+C3rN64KDLApdagNFJKZyIUadnYaPgWmH
AMx6IyUZx1pZWIhin309ZhXSbB2ZyqXU3GdI5bi28eWqCqFEiv9jRtYkSkY+8uslcgWF7r/1rIQo
vD9k8edZ676astSHKc8rKWs59QQsoZs3v3M9wHRRp0gcTEXMt01ubsvDIB0JR1qcXd1wE55CGCT+
gmugS95HIRVxjGzyHN7AWxkaD09/lREROTeuC7jHm4IL0sGiXd7ebTFou9ZuStZwmL4W3haWQt2e
0OzSRJsHHOKuY+k/oVShOqMvw0se0HC5bdteXNs3VcqSUyCtN1RHFsUMgmxEZZLLsje92l4RxRzb
7OUhqzbkFft3PQ0YNdGHcf233jMkghWOsEJ/URJvYCOYFYLuCPPGUCubSdmvfFrjAPLbWBkpfifH
7XqU5EovQ7mJsmmlNUjQOqgpanOwxZfi9X5yiiwwqcPzBYEyNSeTb47O+Zxu1ykAnyNoO0+FyRGL
0Vnutwj8bFZM2ksT+jBavZFXI5ojy+vUdi8ihHAxs9rn2lHOxa0r/DvdpxHV0mVNEffE7rBdYSJ9
CbtD2WBPpeK9StB4lUOYGctFQVtIkC5GoI41+3L580j+mR8fr1bYBpul8Ou2IEQbY7PQHzd3KakM
3SzOy/nprQap7NeRt5bAciQkaCEZlnXdQOJrBUQP7Bp3EBP0F9wF/8SDJBemCy2s3NVPGukPAGW/
tiCI+rGn0sYn3RclWL0HcJUcCPGYPKmfA6ltjb/rUTQnIPKhcdBTFANHODHoq+dc+I3ld07BKZgn
jnwS4faSXxht4UqaUOnQ1fu7QyaODCrRO6Q5I2nPulh1SUE9e+dbulPHAwq7UDC5tXYXMFMFSySr
bxZhlJgN+zRfC51r3ryFU03ZGoSOmL4TfdvoyH18JIEx56KNmeejeeFCa6G/mDvUrSHmsc5b4Ygk
bpHnze1C3a+m7g7RVCr+egIoIQzicOhHfIgMCNp2qFNDBcJwGXdAZd+TxZj1w/j/SZlQlXa80gId
PGe+QvMcXj4Gf+2me4i8gSA4nqy4EkgNpf4CLYWgzpovv7gHr5jHTc53unNk7XkyNoVl4fI0yby7
DLXsXuqJlKvaxjLKaT0igrlOaIN9/R25NIpQYK8rnGJOWYqKAy6DrIbw8PLS/BalauuZHum6IZTH
/VVDpekSMxxKthe2t3PaI2k8PqQgGmlxsoWanD8lPfEgdY2LUuV0hXXtF2Y5GiqQmtz/nO40gTKK
SHtmgOAt3OP87HKIHSln4vQnmA11Nr96mUZAduFuQk34PLF4EOL+AAs9p6JIQA70UupCKdJygxg0
ffK4ttsLK0+lgHbBKI08bODZtqLnHRH61wZCTQXfF3Er6FedXKQo4oIctrtvmhzslmlq+4yKo1I5
CWPpX95w5HqGJnG+y0Pt/htu+CqEBrqqLKu6XsxxTt5Bw4/+wV9DBPQVp+QMsBOnLS4iLbZI8Xt9
xjjWB3c66TAjIR3m74WDzVncz8kfecqaqJGhiSaVv6XORoMFQeRTwOoAjZQHorE2w0J9UvSIwe+B
EFheemrO1qZMHVX2F/1U8Y6x+xAHcfCkD84dEQEWxsB8QLDiUhz+oSPez6Q3/XIgVrN/eZgfdkdU
x6Tq1LTKwPok4sM3sn11BIFzYBowxHvlkaB+a06+ygh0/zEH70JT+ZD+x72VTvLQeKuPifCbefnP
Y8R6aFIQy7HxTQ7h+lgUn+syG4kxRbwCEfQ0CrF1AOH7+BtrOfbUTJ7uxUS6cmL5aOha0XqxVGkJ
MqQQ/wm7/DrPA0N1K3wnHjcFsjr9Kxi7koIPs23PWBiGoWTsvdReeAqKgifMpY9lXRjoTJWpK1N2
55qcd/YGN+VOVvBnKDm4Z0i/dKs7IwBlMTVMJMABCTkmyylLGgT52gAitEbW72JcI99kM83sB29T
qbMWZ6iBZJjxieO/xhC0QPx9GkeCb/BwKPN7QccNV4pKleWDTK6VgCmZqrx2BTe6H6sqnmQNtz4U
4tnGM62so5Xz870gVbVX9HcHrmOYtZ4zDcJValFI/K/jwZQbKeWNUojCPS6QVBQKMZIaDd/l+w9Q
ziMqgaz7if2wZ7QtV92ReUKvEkpb4ZlaXd6q4yIOm0lglGP+JJfawNAj20NYNhOLegv5+D9Y/FCK
ee80cBk5u6g+f6IA4f9clVfrOLXDWdY9qKWu03QIYRTsmUxkvfQ1JDoETOhFnj4yb/Yln6b3JDx7
S43eCm6UuR3Brbnb49HM2DgtzBrzL8yaB8W5x0OVZ68UplAR8CvDSng2KMvjPJguCIhXBT8jw8ga
KTC/qnKv17JprXR+KUsnuwJdZNis7lgXOOZj9K8xS+8x7m9OUO2asJG+hGPMu2T6D3fu+sLAnB6S
6hwCfC2N9R0qsOO7cpwVn+PZsFExOjgrpvefUsbhPuTpXX9Fovhlf4UxdeNB8NXgHLRiy+EooiAe
moNGjsqDSI8UmxcpfuNxKRtEeSwUEbaw9J4GUNV7uaA6uxs6Zeee7d4QzJtN2Dhxk8I4BO2nF7RI
XYoai5Sg16NiBwEV82a2KkMpNMJ1VP4WjrCAjVeyVFJ3mum2zOO6aigmZ/I7cN8oV+FkroMTMqvy
Uj7Zyt1UE06JhSII21z2s7wSKGtyZk8zfSETBoA42dnY9tMBGDubGFFDzWS52eZVoMM1hu3ZaK2c
WbIDHPjcFtTXO6pXyLWDgH3vdmpkYYNcNVLfubbx5WZDfdQR57BPTZm3nZH34G5d0we0qvSSX5I6
6PgNPz0yQv9d1cKkTrr1PTy1ueoMLwvXn3HZ7PuXil9HCPzGNwGMSlJ0n0Ts8x+6nOXvmPoHzk1T
qvpj16Rb/GT4YJbNeiOZVNQML29WGqr5sUVLdDBpF+caKrHx3u1lVUu/v+4VH++hK6FZgXQG0mAt
74pz7cIeTTVVc7bkgjgCn43+zuv88eDsGs34Nc4pkOCK+pptIiYpSEa29ZDOEitPDr1c7p71zBu1
bh46ow8jm4bklhkFZzzKbidoiTM6Eu2R1d88qfheRSlTD5BhZhgHXTsAKMRDEIjpXFxTt8DPeagO
Mt2r5gmy6z0/NHkDonnx9ZWkRUJHtaTYcSMjx/b+wXFWgujsEyDALcXTeyy4Ve5ZAnmlDXWcDEIm
6spub2UAAVDqVB2T2SuEX8PhEmqstggcgv0ZtAi/Y7OAnjqU67iXpjYmaPL8+6CkF0apgEE+MSZz
vQuuWIKxdnkEHpb7Q8HqPT607y8JoFsx3oZtntx7mMtbD2L5hAq90Kl/N65+RhT75pVWIVitxcsT
+aV9Zw+T3YWg+Ji4m2od5d16oRM8OdmXXWWr8euT3fjiE/yVOPO7Ck5oZF/JISgVXeYZF/yJbbyX
ur3nZ6kRGeZ3VZflJGzFTeEOkWKLGNVOlu26fsOH5KUJPdRLf7FvZ+1Qb+i4HCWQnf29MymcxFZm
shP8ualt487tQc0TPfeuXr2ccJFuHo/bFvor1aWzMgiz/Pab/3fRuGALX26ux5zHNmAORwrbGaT0
cmCK80qzjhAHJ/Kwntmz1zy3wOaI7cdI8MNHZHuJX9YbWxesYhUd5Yu4+8y/PCY2SmzaT0S2/kw+
t6K+lQINomv7zkO0EuSdp73ZCg0k2sgkm7LwFpb/hu6S/kKUpT4AAdhs+34fz5/NZsuv7K+eLGtf
z+KICf1sD8nG2OWUJT0LsMQA41uQB4jpzIUszJ7XZEKmC1/gKihwWt0aogmfMwjpQEpC5PKgFOx4
TsmB78fPzpPqROO3rRkeeW9aORdC204cSHRnhpxxKERrFhIzdB0ORBwi+x1Asnt7DWez6ujMvmP6
Pux2s/RgPzku5ni0WFN0DIKaKPAQdhtzhJJtQeIPbsXWgRdkKdDRU+XAp6cJcSDOIOF5A0S7R61U
3JlwJrl5OKi8a2hrsZI576l4ei95lZx9kKnTpy2dE8NnR2n5QJ2sTYOFZWcmNqjM687JKqCV4YRF
CZkJxuR9TpMQLE0W3c1Upc4EoOi20vsJ4oOylGqJrdWSv5wUHNKdg19T+DZmmS+51gzJNPFdAP1i
O1dRDktZDf+kArN3U2BaJG2wOgYS0D+UqGtLsc5+acC6Z8d14v/lQeH1swD6gC5xtAsAHgU4iK8U
tyo6kQnZSISWY7g+8vEk6eX2GHs9T9wmkg3+JE5kCzQMLcUE3pCfk59QAfxwi7rERhFy6OeEwiH5
HUXaWhT5a9Q9LGm0CufbWshvJyl/O8RGlCFhcTG6cebtX3khUiABoCnlvvc72bWFct0metwaE/yK
TLdMXEAPNFvptlEnXpX23RCSAmA1wqiqTTBsfe+j4lOI1CRsFJvE5aLwne0MtOzI+g5a77u8Z8OH
Z8KJt6TY9CTuSiuzgtH4Ea/bXFeqrKLIsfN7uCRHWxCmbGHVt1slz4k8Hj+Wl5eacuquDssZgsWn
fLyLrBjVgQ1UUvQfSy9gPeUwH7pA2480bki9roTKAOjtojmwLQ68FOSiEpVI3VKj0whIRw5sl3Dp
kdm6DDUeDFmvZ4tcv2X/fp0PiAsq6btSzXw0C+e6YfiXUSpZtDQQoHCo3X4XG6l34bU2Yj1l9hde
JCnxPUV+FWREtmY/BbeqZFfHu6mUjXCdkfJGqQg8kIHTZuLMrSNuNQp06eueUVOsa+mUNM6vOqYe
j2Ia7LPhVPmELDoWli7+u4T2gK/zAEsZl8bLsuSFIxiogP/ZjzTgap4q8VDLfkTm+9x+DYmAWowV
GLpKzE8QtF/Q4X4mxSk/nvbgRpuOstFd9cZi5EWaf25SyUDbYvWTfcl7Gyz3MpLw74wc0vcL1B4k
NtNFnz50U2WCcyQlpoITZvxvsNX19zTuGTaVMniahanf55e4+FVJ0pt6TdN1AkBql7e1IlpyIN3F
0UeYbPr1mQEI1wJBJNy8fFqT3YEPn5VRtt6EsJ/YYmwTYndmc/eS+8J+0GxZiJrkCP+ihFPnBGac
xH3PgaqK9j0GsLb9SWDQrVZSKon8mZ1AI6YpB4PANJdPoV2bVX5PbQv0U0YRpCV1XEwk94AmKIzx
cBZ5ZCNxKuCGtFA/VDaaV+9nG8cYehBcuInPFUEFNrQvOCqizCaBkKVo1jTT6K50zqexs/bkSbQI
ZCpfCtFvhPQU2GPhcTOXuVRQfsBsAj5JSVgwXPgaBA32mXA2JguJ+mxku30AzXTkdRDJsD/h1+Z/
6ufMlpiqyVjTJ71j4qpsK4u/umJJEI2wzyuLAZoKFiT+XNL/p8brjOuH41S1GgT2zc/58odx5q3f
2rFOGuTXTRaRzW+n8z5ykonRPWKSW4FyjXXb4g8FBPBaJw9lS4PgelQwzqg+34qkPLHAdR0cMt7D
qGEeoy+5od/nAgCpEnoRUFPPWKEVsvO8em+88Iov4OpyrH22MWJk/KPY4KmubMSgPp5R9PuQEgJX
zc9xgX2cGvLqV8l/1n+MI+aP44zW3vWaBqIBlxpnUvjblnjqzm2IY6Q1znMPyTckgQVPaVq2qRR6
MuW2J5o9K675+C38fRKE/JVdq/uaq/V+kEg8vg95V8dFvy9su1bOHJDLdbgcKQZqh5/ZnevYw8x9
4j6htQJdTgAN3oHpcFGlNehGHALSlhZUC2mvNuYB0S08EzPG1yokIjrUZANXahdEbpLw7Mkaynk5
/f0nW3ZLXjER3yjXChx2J6tlkOhp6ch6LeFROyBYV/47N2Dt8Vj7ktBV0jTBD9lZ88Feri2HOAMt
3ptRP/gllPFBseYZElFmC38a0HSDOZUIuYvVlQJRQUh9/Tjfs1jDDhp1zmkX86WfIQNuSariF5Bd
Nx4dTu1gFFAS86tNXw/3LzuLgkeFgqIZHvK3fFn6qvmbUS0xe5turN2bDPTGeNbF1GcWDQvnE/WJ
nJ6Sg4XdDSUl8TwofjgCrQgAG0ViVFTek0tUeXFb30nZvgqaIZtioKGcIxl0J1EiEyJQQVfgsCMS
79PgNsGxYyeoVL2N3Z8ASpm5+l5MT7XmRjxiQ59xph8Wqysaq5RzYwdyBBFPoV1VHW/h9tFDWLoy
A4v0CxgO7WxB17sXvJMSSyGGGhw3mheu0+j6pCt3g06Sv7KQnKIvC3PeHWSG8GYq3OxBx5UI05FN
pc/DE0R6G10E3efIffJiaH26dQnQOLqS8xIHmdlpCGjYoUW69WAYSoswAkqzPjmd1BlQINcbg3b0
n5uYcbPfRz29vgSFn1I/P4gnAKVsniAIe642jhCpZ57JevxM+wRjGYONlANhCKHtcVZchsjrlgb4
+6AEjiUmhoUDQmfMAOUd/9i/bUFLal6khv/X6DllDVdTOZP/k2/WZk32qM1WKtXhp2qsOToCEgVx
NaAWD/043evxOKCLyFor9ncUPqqSQ20AajHzbwv+yxedVh84gukF7VgbelsZ0SD73bE7U9ttXv0C
tON1+E/zaoJOn2tJF56JMz69nqosJSHENY2qZVfz5E8EMrVSaj5tLzTNPEYdb5UmnmfnVW43fF4I
y8wTTISYxdNMqn2GzOFg3KWyjRYUcbmcL+JmHK21BXB/71/7+PmDdfZWNNcT3QsQqEF3hWQ0u3eO
O/oLbu4zdCi2A0asJxBvD6nQqQIKhRuhSjQrqtHivISc2ZOE6bjjBhhYwcu00ALgoXNKNsSyAVzj
0oIDXngK3/34qnh6l5g4bZtfsSsxnngzn/x5j5UTgkYrkfnhDxryqCupydEggS7DgTh7CoiIYFj+
SgvQJxwT82mI5sYLATuADsaIC0M2+/Yf8BuoAmrKWFAqv5Q8nPze2stiathWT++Wi1Y96qXBsQ8i
JZ+QatXMd7wuaf/UUdELFhUEH5MTlmC+WDizioRrjHCDwYCc9fOzIbJ5MbdD/AxQhGT2GxtZDvz7
zSv0KkiVspkm68Dj0O32ynpfg5zr2dxb0uG55QoCYuGYZgOBP1YYTIOPeRNwdHSnyYJUn+v4FACa
ebXySdtR7peUmvEagyGJz97KJuqDRzfhOy+63KUnGAwwshsbU2VpOoCCigcEyllp8mcWlT80+Ig4
lBCJ6xAA1yEqtZUKdgJe9+u+o10l3hlt/VXuNEPXV3/dVsBgz9aPyhJ81gL+Iogir1Z7QhtHQreo
R87QbiQUvIqhotOhvGu7smU1mmjIFfO0DrSNoUUpybUZtAgUKBrokm4LE1IZZm9qn0cujMZqTVxv
zklDeCZxbcc2ZEi7SGDqMzE2fRZ0Dxrmh48iVRjABIyCwPtm/dkeym1jeCjOW9t1kmwIsWjMTHKj
dEC6P04zcsmT3XJh6Sv+VBajPg5jnF4yboHb1bM9+01oYo/Du0QQnnLVKMSccLAL0BvdQ+ex46pM
QO1LAIYyk2qGdJEF9UBxhP2sNCjry8BAtgWEl9LEfZY4QbAuJARL29r0yA9b94LLGRmGFq9QQyNK
N6ICYAcQhcCdROJ0jwaQAeBBulCXT3YXd8XmufZhGPdQnAcXVecfsWA5FptJV7r0/4fq1hHZpkJq
DyxQfraIaiNu7pCnx4X145U9tGO+DRJKkIoA4amphPDbPT3tL7C909Zmc3a0SLn0VvJ4fwxwhpNs
iyErndTETvVQBJRLjAm3e7AKDkaSKUh63VS1d/gJOa3aeahNibie/blGd0ayGy+5Fhps1HqzYQk7
8pseyDbjdTL8oq3IrmzaYD5ygOyYxzxMOU8VGEsfgyjAMs2C/qtlqYywVy3a+Ii1CbM2rrtsJXrs
oXid7Y96Me51DAJAv7sR6uXVDCQQjGGF6JvL5/mmRZu510NO5lZyHTCyoU9VD83henerku+Y4n0o
8Emp+mrBHG3qo5eotdg+hnLeig/FD8Y/mP6o1BnIPmoQ/N91gcElGPZo3FsomXSIt/RkV8OHZuod
doj90yWAEYliRrxtZdANza1fVrShKnXqobCoW2dR9UsWKPxoIkI3kptuaKJ6xkUfdcy/4WMjMf2T
v45uG5OuN4bYx//NoDXh+Ka+a3K0AqiigAmyMTDB1hLcOHP9zKjFxtGAOL7bpPhngMKEhyXZ2eD9
lhBh+0rIN10c9tJmvhB7xvCNGKciIgYbLnd7zHh2IlwTCRu5sgmGwZqwS1tgnEETCnajmC5tglhk
ezXlGKUIckp5GVty39Nf1Dc5xevIin5+gIJbGnjJ1of89F528gz5tu/Ax4SAiJI9RfCa/KZnX2se
f/x6c6kXeSAS9e/1M66nUX+b+AJhLzH5n+ZD2tWKB3zLR807fD2xcjqIRL8Gi2zOxRLQ59DiSAUw
0SiZRd2iAG/Al7+fQ2ZZg3UIIRBZt2sLG/h6bMKh+JbiQ70DJE6FY5OgF5Z6k+iAoyGbPPMRxkjU
vN7/SxEC3DEJkYVNIUBsQZVc93OxswLDJ9bb5zay3cj6o5JHDKs4dgirZGO/gAIywR5kFHQYGJ9E
ew186Tljqj9jrDPaCtkwRQ2yQPDiCl22aWA6amAzvNF5RnliRM/4cJo5LJZ06C5BK0cLoPqYn+Ql
E4vZJGtvzKLdVyXl5/Sij6fYZXJ/Sd3YJ7+PNL9/rEmLEQuvMUyRhvc71GFLA7U/tg0T9fAP5v34
TD2jnktjp7Jg12yTi5aNpmNh2vZnVwvk1nmWX9ZezgiKyl6Jn7tVbRpV2kWieyiWPabPw8R4Tvq1
J5L9Sdr8bnZ7UuXCUkhsh7yAPcoUHp0bRvf2hrHfMlpQC4RVCEwX9RwSwiIoT318shxBHoADBhSW
xTdZVa3g+uWcprHclV/jdJQbpx8XjP6Sc0J5DIhNjRIMar/6I9KNLikYINN71a41kuq4oZP3SPH4
xuiiLUbdiRqsKM9ZqA4ceL541/5HBP5zHSx9X27myr8fL4zctYVwchItoq9JCGp2boUHCP8f3OJA
lmOoQAhoNOJWWnUr9XODfJjOsxgDygZHr3na0KLqe7HWDIgJv2AjE4gFQTcHiwMiRkebBzbzSS1Q
7zsViJlXVpADpM/K+a2x2FGN3BTXbJZfIwEK2ABBu8B8P/jAhYO+N2rOcYGY6QZJijJ1XP2WbngB
oAdLo+5UaKDCTMYhI5J5k6rCJc9hZKgidCb4UHYumfuwD+b3or0dmIH+8H6xBRsLsBgkjcvAW9wS
p37wnMzjU3b5Z0RbJfrOZnUOewRRzgt85k3G3uG8jNyKZWpX9Htn4eOQ5OrogV/M4/L4Fi9SsbmU
YIoRm+r2EHhiFeHoSTYHDiI7+/dNMb/oxDKFgklvMO5b6q1qj1Qi8037Y09EtOQmlzoyQaw0JOmP
EMbAvlXxDEOTlyX3D+PHdgvUjl0c4oOILGgKagchYXesHxZvlMvonjcRPFt1n2NEpXlEAJFzsWDa
haUYVbHFvjRkmok+BLXU5A3OS/PcKFeWw6E2H4DKFO5fsbGzrixWARJBCnPl21a6oBEKT+rP1aYR
kGY3U8Wp37wg5NA7mhlFYn/K3Cpj0lBFMhaMu/dirR883gOGCYRwVQYDxebdSyVjMAMSk9cnhGqu
AWh4ahS0Y9HvMOGaxjKFOfhum2pvj5qARTG7m+wKorjQLugrFszSUtZfGaUIceorgK74cRWqUKEd
6ZoscngzIYzptjZi4fHYscvNeC0q9HqSxSJ8HnqUcby8MhBEPePkubeTAD5i05TIseOIh5b1lRwH
lCnviO8vLAvKV+ghZBqIS6vohtP9cgCJzboWpfu9OXj4bTT5hMSA3kpRMsICLJCwBgxRrzBjn3Rh
nkI0WTQ55Y7WWa04uvgrFtUXBfxTA2ulFQA/PvhdDOl44bwX1GnZgB0SjbvGAHSgbBIGPxtqRXdq
o+FzWppPqo1Bqr95ZbtKqITahngiThkHNXD18P92dT1dYUf7Rtmn3IIP2cQn/7eEc3lC9XU+EMoZ
ZR+UgDsXVo2aFTxMZDRGGMJ2O0xCNERGz8W2XDLQWMKueWTxR5GGFCeqaKZ9zU5AFMkyVRya1lf1
Sxe7zet3l32yM3QbID8qyE8NgS8qriLWt3KJRAvKdH+J+lHHnotUYMAoJla43BTdaCVMSpoiosc+
dMDYyn5EBOtAXeMtWWaK3J/BxCd6aznkAOXYVDgCVsTOt3bJqYoUCEZAlbuMt64rOUZ7AfK2o19b
vu4SoKhtjPeAz9qTp6GOyoGXxoBU/Y8oy6URRo1wIe4ydSFkF6PutQKDJn9kVW1HbKLFqOlfPBh6
5kotaGC8d4i6am0rZUU1SV49oUeGvyjp3hBkDT/MReQHkxM9oL6DtOmgC25aMVnCFkqpv8KdqQTK
SfB3zatNIWjJFwpSkQyqSqkSvnaq4klCqi7KRRpF2VY7AeE8fHAA1rqkM9XP2YFAAxPKpRV6LLAe
Xo9UJfKgeBpzCUthYk1onsdX6lphCHxvtQKk/obpf59einOYs595aqCgKf3/slSAUX0tjI3x+wkF
ZEn+r1MdRob+wepZzEVgje/+2Td7mTVkqrlpXFMHkPzmR3GrYofKwuiLVrqh51RNkddTkSfOgxXT
ojduUNj9uQT+Qt8QntQYkcz9aBBe2EPtyv95tEInpahPfcBU8VLGgKJhfRLQlptV3qgVN2I3DqaW
R3PgkPJb2WPGzb5CBUpc3MppVJbNwti8nrR77IjYBc4PDOFV/ooJeDqxiv+IgPJQWYIBIN0ux5sa
jMyRqXTyc3bFqGxhH7fWF6ovKAkI55qcLaZDSEGHRntPKmdOmaZIY4uf783ITSzxDbkdolWrNQWJ
zJcph5M/nEi3n3kbI7q6YiEQW+p1OEmPYpqaA46zIo7afjANBw9i3qF4tlFQLHFmOoiLLStVRyDG
5Vr6rC7ToETAxrYIEDFlkMR1yaeDWNNHR1+qAFKpXKVHbO4D7r3duahIVTWvuHS2QXU1sv88N3+B
crShPJWroG8xB35RFHj2T2d41lxKtXQoBDAnstPp0hxcqIvVlY0jLAEKtr+eYPfQ2KzQco1DTMja
QEgOiCV1PphoL2HTky+yIBMC8Rp/+Krxu2K5cYCvXA4BkqbFuWEEpi4ZdR9ZYSp8VMawIbDFXXks
tm/ZvScFnWRxZ2axO2syJWFYtXGElZykAxAsRDpEFmQ/oaZXgGvm2+hOeJSaPZtRUroVPuCqvUoC
DkEdVij0Pb7NbzDvkWJOJvPCiDMphYm86Qi8ABxd1QXTBgY+wKsj5LxFbq3rPhJC9/pkLlPIjmbr
dZdvr3zZEhau5ywKD9HAOD3mmjYgtupdySktjWKt4y2/wkvLUgC06M62rCcDWFO2Kja7uCD4SQ1M
aalaQKu4h+UwYORDVu6H9JIj2zbuz6t6qfpEy9is90PpyaF9dn9Bm84dytjTnkED2JZDPfR+u11P
H2x6FH1hmcA8om8YxyhyOIaN1VLT3TW4VOWor+TWRGmYYPSDd5Q9CEjGH100UFz/6WncKkpZSYc9
EsqrLRW29gd3GbfFzCatCOnjsbVmo9mRbEtV9Ed3XNN7T34kLFvzBk9Y0isnJn91rqu2dil6KzHY
XCU/wBjppwEo4zsMq9kr/Q8d2QC4dMXqC5J5nS/ciD8HXKRmgs+MaeQiGUhou4G3GwKklt1JWXmM
OLZ5FtpgtXk8zUSasG425P+RPwhUPd67Jw6eAxy9J45PmrK8I3jVwT8nLT4NQS6IgzSvd0j86G/a
rckPzpCVQ7fCZ7uVL9e2GYwPREN6qXcrT2Ud46sxzBgAWQxoMZqjWAqR1di01Z1ccGVl1H5OpV3l
IajODphMHaKIZHJgQZab6U5rV6yQwKWYYyOQ6R0UyVsfY4VSXc0qEtts+RSO8fnYjxhuXhcg4dq5
jBBNmVU/RMj9UUFy7aXjO4jjz5Tt8pCTFEGW8Jh0hZEPKm6XHR8DCWqZxuRk64F7vkbpoH1ftaXj
b0Zooh+DIZ4oesOLxVont8iF+NW0HXwgfOoIbtGCzmA5Lf0VlrajvSvP5Izu2uJ8BEwzRkzOdp+B
mi/OAcE0etmLCtwMDR8++zRb1qEGYbR1qe6ZljxVwN9dp3ACuC+D8FyTH+q8GBgUqGVXZZjQCmZ9
XJ94RDMPF4AFEITY1gbIrr7Tfx9d/pcNB/pLDOB3I5zD0GpDpV68iHZDPEUwNMDiI74HTdvJlSsT
dgUAha+aDC/6fcjThDX9bG9BMaKkAv3Tz19XF1T0Fq4q9i0YVIdzG1wa6lLuqSzl6ssleWLpTD8g
fUTLAWPqmIlVLFNr5sCVILQK27Fuu6fv5PWIk/bCETJgKJ3n9EOuunWmriwCJg8aAb+8F2XoG89i
msAI1MiRoixdoSLJaO/QqCho/bNt2MNDluskAxGWSavep5uffX/eTrQ6TQu3aYykY503KCxbj2Y9
uTn8c31jNx5UQIJ6O7M4p7geIQxJP7+1DSrn5W5z9SxCKBTyadhH3QglCNYpi2FMCxKl7ZgjIj0x
Ulkph14YZsmTXEDwocpfXUypvunkA2Wxz9+dRyhmn/Nk+ejdnqpPjPQrBK4Ipo2hO5jaN9cpMiOt
eZRSDQqLKrtV5b4Z3VLhFtefS/6SpMXb5SugJdnvO6aa1nuSYO3ju2wDkhlkYgEfUhcZZpdyT87I
q3oip/xA8n8iOgCdrlL1xSrjcgm9HQodf5ynuKBI/xHAWtiyQKX0ZjH2zFzii7ykx7zHgPGMj/qL
VTExyotUBbRMvq86VK6YXzU3rvZ5ME0cR8Ed2ujsNaDMFR4Kd06k6lCUS9F/msse+q8T64R9LbT6
qshFnSJsj0bwRcjOCrvOlo2ibzh45juzJmJSx9Y1DnCZiJjPHSSvb2ueDCnmcAOvbPKEF3O7j7ZD
R8nCs+vli3oneHWXGH2f9BKCptp1uOrhOADsgN1539XhhfOu2Wkyfpvr2Ctb6xOW5A6sO3wSk3h6
Ug2wCkCb0ir1lcCfukhC+zbbqhhRvXYE2lIoIOe80giTsBOebcBS6t7uNp7VcUDkIOSlPNeJUXj2
XymNBTPvuinV0+teUS0/BLn3CXaPUfK8EnaZRionxS7gT+vEr8jcECAPNWGBkjke/u4jwkoiuKnN
84Yy0M+rMUc+7xoBypCyUyXE9xm6v061SkHxpcHmqY+zbxg9kP4R+SfabaVEznrUOfOFuUSf5ZFI
A1LLxNI4DgqOKBgPYW2iKy2e9oJiTJ7vWIcFL0HOc/qTIXX+DRwX8GHctmmhDVOczE+Y7S6SMYK2
Tm9pgxrWA8HjJDwFUiGviRv7r1nViQ2VfVKhHO4caxJovkrWgZOJGbMVU/LoaK7P1CFuKUWEUNB0
hFSu4YLo8jDzY5kYvek/k6KsWgIVSCKh3avbEhZc/9hG3QSkxhuHwgTuva8MMtRH2I/RN91hGsfS
EWfeXBWz8su6t9DdF3ZNq56oUvnV0JeyQ/CeRpe1CDzQimlbIwYwbYqncm+LtvlsqJYR6TOrlvvw
VIkARxwTu4dmfx3cCaZiALasgwDLXhit2JIfG2j+pHoogRYIqL7l7foCnPvR5uycXwa6zx6jnol/
iR92LukZv7aIM+S685LtnLyQrMXsiyCnoWqSDdhi+JzTp2Lcj4uwHqgOUdlnadMRQNyU3BoaDnB+
xG2xyI/4UTOqa6LC4qu86q5n8dT44sXbNX3A0yHnt+BcRum0bFJ7o4lXnuPHyTFh2P4r6QNzON1+
BDBq+jyDDClndtYZBGEuLfsZ1m0aanhiGaTFStBRtv75B2b8qalt/bG/S9oAfqvnDn0TrsTHbqe/
gwHXWpjXhtydG2UCDvgd2yRccdzJ6dv5j/jZ59MHzgeaUd0Q2n6aoXRCE2SL6ihT1SJizekFvSLC
lUEwSpXLWusnHQCRykMhmFC/Cfkj+js3bl8xS8++k+BjWoDQBTSfv6WJ7nWTI5ou6ABDjy8Xfv+U
jOBYVCsv98MuHOongk7mEA5EBp05K9nesi7vYEhayHC67r+3F7+l5vXjQ5UazPTkSmkgFr4WB7cT
AHRH54g1Y9eM4yRGJydl6pt01zjR9CYGqHoefqP9JWnR+HePzHl0KlIaP+RtEHwaJxeIvvT6p+xZ
/sd4fgylMztNiAbb82WJBT62S7W+NgkaoHi1rxgyVa+pEVJgPPQGdIuxVQBtGAzVNF8mFDByDuFh
oEXNpDC17rH+xH6u2AHW1BomeVfvMzN7HIuoLMim5a4sQM9sCxO+MqoahzCln8DM55KKxFru4e6H
Tzt4oFKRJFi8IyB+XDLntKsrHHqnnQhMTXkmkgJqW2v9WF0LQ0cFbGUoyCiFFV9tVcGc+uuOa1BV
+wOBp+RUz0/XJVNKMDG8R+ddRxI+F8zCv85zoY2jjg0zPiAzfr5U9C7GAycJeE5wiEZIqGdyAsdw
RkJzyX9uHIPcgz2cgQw4Sgd1Mll6c21brvOsS9T9q3ql68JWCnEhsmmRV6ysGYSE5V3k4mzK5dvR
Tn3p4eBmAtWg3sMwb6Sis5FXADNJw6YtuRY3gJYPKwU4k+OULRDwyUQ5vA8fUY8e9LqUq+jgU1xg
uFAlzf8auklr7idlNOjuGaiCjh60GD3W9rQFOcm7bdvLraGatg4myyK+Z8L635OO+f8nIPmzqvjw
vAv/jryGyjJ4FovQzVyhb/MjFWaGWE+IzkTq+funKin3LuI603+XjWMnI0xSllm0lHOdMrbD0kxt
Yw4dV4McIA4Z2JBNhYeVJPidGuOTOXIAD1SidSbqWoqHFLCU17yOVXLQGT59AA8dBzReBnh8CiLT
LdXlKDaAGDd9q9LcI1mnnnkrLBik43xhSdXHqgw+CY0kFmIQPX0e1Nq0WjF0I5Et//4Ih7fHNagw
qk+mSzAT98X8jn6PKUJLI2aWrx6xB4rtk3/eF5Me4G9BbM/1pxu/N8Bh6c1oA9CIzV3uvH5KjNKn
At24R5SMfghZ323YtBOGBiMAmTeXKxoiau8NcrPGYZa3VReOLguiqWG/4uqYrQamJopVtzisKQWl
abzVyQtfcHLgmReX+SOD04/x4+sl3Kf6NXsMsQVWtGTP1Jt7Fjm3MkP6OJ1biON3aOAzu44qTw1R
FYGnvW7Sbp1A+L3LZ3uEKSxz8Ts74vvwQvnSHWQkx5NVGdEClBRYD1nM3kxiznfkFTLNjEE7rlgi
aRVHiJGuZyN09dPfRxAeq8fquP9qg/OPCsyZzL5LyLL5jPDvneZhNmow9Xk2ERz3Ihws998g55VN
IGfkFOkzuriFkNxV1J6Y6g7ax9eIB4JkUCI+kAGfcCkAbg1CMKso33aQeYUp9OYtYYOk6sIHmfBv
dLaTBTbtWxKcLM99KngYCF/g8h9119ipFuu9+eD1BJqELQpLZDy8brp2r0ShrCIiWNyviFpN9pKH
LyJL6GphKFM77Y5y0ycb3Vjtqrs65sTFGuFQ3uNanbVFenWPE/j0E7YbVDdeUUJ1JukyVkCO0jGu
3+K1ezc3BNa2GJbcION05G0jmgeOS9E1DVoBDsP+HyhOxtVpFjf3huITAY8ZQplAiMadXUm6PhpU
68ylegb7sUNSQn/zMdFHddhj+AtnjG3JyiR1h8B5Z5gukqFpFkWrT2lGmnnB/Y7xSiAWKBoFucZu
pE64nzwMpg2yKnjKShQVf2s5tb57QlWzNyyayug0uMRNk1qInC/rjYK2hiaHfo8TpiepdexpdtDX
t9IW+SlJ2o8dNBR4gCVCMmJT6OamxQ4wpCx2UTAPWOXmLXA1o6N6XgGuT7TiM+gxxNvgEbImXTb0
Ei9yzz5drKunn2q3AthtjTcZcSCRYiqTrZBzADeFXstDQ4732Q0Xc/a2Yt+TtqwCywArUyOW5xct
TnaVTZvmbKdsSLLtNXS3s/Bqa5B5mEMWaJODKT/JZR0E6tRJpFUEkNFkd84WkQjtCUvVb0bvdl3g
dlKRTTZZ4HWRqjsxzzwt4kbJADuwOCH+cnSOFXStEHah12o08GUxnxiywZg4BifmL7akdT7HLL9E
6ZpIKNcv/XmdAxQNsQrrLFwbsw+LvG9RkUz9Spc985C02qa1EzuDnVPkochkZSaoE9VnWVESg0BC
jnWcT/Nk+ctE2n/WMXCMdGhj2i1+r58L/MhMk/ByDfu1zegZxZrOPOFnnv2Et/KXtydMaW/jwSSA
n9ub6ePLU7x+fOjTV9ola4ilrxkT5Y7YlmxqMCKGSDaWkH/7gqbOE/x8oTXrknfdQ6Amavmjf8Ld
lj3Fp1w/q14nrd4ouIxwPWHsL24MwH5RpoEQOfckNKEevkJZOnFifkn6R+FXy/G+Jz9Cf20vyrtU
qXW6/uynAcQMkLJJVANEVBF0O9jbYvWN2ZuUrM8g9y7xMNRreCcRlIqwOpQEN2T4oY4F0qjIhubr
qnMGk8vyKRF5bniahCkCNJYOA+nsHvT3IvXV1tP7NUVV/PpzF+zCNmolJkC7DGLRPZzaLtV2WoDj
7tN8R3v+7gdcrwuFTflUpx00rgC5Zbhp6ocaTBD/6mthXcDEZ6GYZ2uwvA34mDluyAdmHIikJtNL
H1Q1ZcvO25NUFhBnYv2phfdeBHuHhUvRtDLb8FjcpWrN8qDt5QVy7fWi8tXanI+o6G+1CadDh74x
WbIu2VwIKQiEX/g09PDFdA4k4ijS/4gZUJmu9b8F4POeBvtEAn+TniOKw197jRdK8viwTLLurPvg
rVaByLcZI3A8qvGOYnAJdL6MJ8txd68G+EjBYkz7BdxJ3R7/t1d4AqmTjkvIANEpkzWghT442y7n
GxFPIrPTwMuN4QXyXq34fIAmJT4OsAA+QZ1cGm9FN8OWoLa+fQym4HHCi8xTpjIuUA3JxfA6t60h
+3WwssJ3YAydfGgvj0pafDZZn3HInxl5WpZ6qe9npLRad8Wdnvhd30AiNFQ9V3j7CUCDl/7kZenO
4VyRwt2RBNg6rOALGZCh/neFmhzpcEftgjtKmlTMfSy4KSPs4EO46DceTvrpTOT08RFeg7EoQckV
WZY4Crk0RyCBfEmLhJgNuixC79TQWNLP3MRudfjKQzs8P+7Canl2HRzI9+cUFqi6TXEWlOayKcUb
bjtU2aHeqycvSUsqIYWvAGF9LJmxj4AoV0H3JvpfyjeGE5QOt1fG++2FqKm/tdJ2V5ozW6kPTIOp
igyBkrpYxr15pFp5F7dZndpPy5XAwSbH3v+YD3E512J5FNLzW9q9ggDyoxgObYPwvVT/v744jaJH
+lGlmHzNfuSTNQwYpTWeAY5T/El1RlHZG89bXS67XwJB91bkz1ziP4zUEvav5cNEyBpXmfp1J6ul
W4o5Gli58duO0dO4d9twW5JND0009Zav6kZaN/La+VmMsJaSMy8LaD6N1GvJT0KqtP74K/jNvI8d
qdmVxGKCHSuchssmop0ZMb3T4WGzJX0aYM3yVzm9d3St9C3zRZMta1ntM+SKC2QctQvXN1AUKrU+
xwT4uJmJT9DDFkrSKxf1LodkczA4dvj0jsUC5kUsjXmfN5LBqpt5lIXadnp4lyJFnF2PSfSR45YI
P5yVbKCeSawbDM/UnSQz4nnirvjVXlCJm8UQLoknN6JS93Me8IRvNv6U0eIN7SlQT5xv0zneueRF
cDTPf56VOgniXpSUPRrKYUJMHK1DXMHh/pQG/KdEbX05GnrSa4+KWASdVrMt43neYcEqILE5FH/N
iOlB4mhSqQjJBfKpurnK6B8GrVISwtqYMjNpV6V5aVKm1y59hS92x31hoyB+5ALgQvnRKdKFjaSF
DXGAH/IBsW5cVq/C+64PF5ubNPrQ7imI1ZbYa88wGeTtwBf9xwxA6d/uZv3VDKDB5LDYk8DX/ojn
z9SBhB23bAreCLC4ZHkKyEeCmQnPtsGYoFZLLMe+6uXWdn+j9rrNz7Xf5s2gHs2otY9EGpCWhRat
B9plttWxRBqnnRTHgjhAyHbAmH0q7DG5rBG5MAC/0TGgGDYyoJILW12GVAEKhIQ6iUdSeVlfzr82
H2FBJT8esoZXVrW+PzLmUnRi+YDi94J6d3OEbqY/S684NRzooKMTlVRoXhHwuI59vgcePlonht9A
hhLwLQXJu0d2OS+dvyEFtOnNuD1+glWUXrpM22bhRP3/1VMRzUjCyassNJIPibYBp9Xq1xXzxrP5
Hs+m7u8YWegKpuegItThaqWzFxl16oSCJ33oqMutqNUSrzvgpl2IKDxOiXtXP3KScReMArUchZv5
WDTGOgwzfy8pDY2wwxe/wc4t9oNac2Ze9RULk6q5Fhx8OqdPdGWzHExezzPUHPO2hp0lEdgCEtP+
haYdIhLA8ynb6+hTT0LO0qZmnLHXLeXwC3mXioo4tCrfGVMefqJm3FK69NSBlUzdVkfkmZoRnJ5+
zExbGWelPCZGK+Jg9rCG9JdwwA17riheO0Jg92/bqUJnjSDAr1N5keRQdqEwzjFCgNrBIc439Mle
GN97pDGwjqJbOjYPvbIpvmsvvA7hXcuapqN6dB2zsL9CVsAIozl9upDGAWVxSq6xretHbt7z/HeW
xXrlIClNT7aoO4grY1o0PDkuqdojcPpY9JvGr4GZ7prFv0EemLkYs2WqNTWmxWPNal5ayjga5Wnf
Zj9DzgEkKWYy+ht7P62S7rToKFo99El8BFD5HU6QxEI1zXk6LVQEQ2YXosPR5ZoqlFRGdIBhiPxm
sGVbogZgytLsQ+6kNwoPJbeXP7l5Fibbj+he0LamAo4652biaZ0MpGbTA+c+jX/erau25e2TZ7Z2
lq2cSMVmEAi293aTOnfnJtwcmeZ5kddMdMY10RLe3WRX5NnKPiSfhmio1/9VZs27/2Qp5iOeYKHo
2eXAWQrLZBV7cTGfRmfrP8XOP85T8hdBppVi8zR0963AndWf2m6BPH0X3lGLEu9jb+FjiRFU9Rq7
dNPGVKnixX/U3pkM8jDjS77j+pst8OIwrO13Up3ia3S3td9oEh0X2KGCXGLlRjdGxi4pMf9XhWi/
Mj+YMDO2c3P4txsWKxZpP5/x922Ly7xwaLjURIcEKhzcAJliLqcnlXB5USkpOPIF6rfkRhufJNwX
Ys2nxuZ0mWNPnSae8h0n4cRQmS3w9EUPzP6WjG/a20UoTNaVUJTVWXXxZlxj/JkjB0nbgFVWpVud
ugpTEV5FwqxPiCTEuAm6VxPD/nz9JRnhn0HAO4t9kRdm/pdZirDJnBDK2MlbMs0Qxa8ulhHAxApK
aaHjfglpZajJ/nbyM5U2T46UrQGlxiQ2vyrBd9x8XlBsbAxTx/FRX9tg9dehl8PoUH8qWa5KAfAd
a981z7IWRX7IvNFJeeUh0hvaz97KCXTj+K6V/sYlmiT+HLdbDawSD7WnNqJbnzY4GQzI44GjTRer
KwtFR8aezaWl1KJMvxHA+BX/5zi1l8UOiW/QLGtXo/JjkP7k3XTxO5SFKO8ikcNBBq9fhTZoi2EW
/rv2yaP1GNGE/oAKFF1HDZD0oktdQ6moJidxzA3afFj0+Fx0vWzd8baGRFGPIlJRSRc6yuHLtvvq
HlqEBLvrpjYwA/7i0X9e2cKCJyLHOmiysbgUGBfHNTiBP+4+SNJUX3CPj5Mocr0SmBKHxXzlwTwR
njORI7j97ZFxge5CSbPIQ+CTucpGqmyNCe22lVzsSgLT53yV7RRaCjddr0tkBjFZPRtXzQmr+4NL
cJWS0jpskIwgNJYNQN8c7ZV67B2LwPH0Ir7Wu2c5b60/wSvfcatH+WvINSo98LDO3A9Rp49zUckc
C+nnr4Ucfzf2m96a29zuHlsONpRBPh2kwe0l4gJ92oZlRZGusMvuILONb6TXAP5saX38PTvjoAbB
sD5/dmn8M3cZEvpF9Yw+6tTL/EuJB4nq5ZjMdWziIWdagitqSMdmeyi/9pGCvc0Wn2fucTnqJ2AD
/a+WuSGoVLD4PiztArjsXDPcPBayPWvYIRLH9rkYrZUsVRyj+8LcJ8lAvFpXGDI1Hjmr/j7sxnw2
kwR/BnkFuY//prdqIEoXBXeNx0VtnVau6JFXbbrr6ogDidgFfgZwsfhIsya2scOsaERtlCQWZp03
yXIJgGBdS7LAlJoulg6DG4FmBT2J7DflQrNrw8s1EjCkoYQa7gkpGoi70z1ojn/M8mQRByWkftXH
k2eeepvBQIxUYELDU1gasNivz/KX6+B4jSvFi4T514sMsRiPjB/6eW3jSuX/yI4oB0qNc88y4oTz
XdUORiN5stgSAyZxP2suUkyVgQ8ZiRW0EGm72iyiIbQCjTqAcSR+FXra2VXNOcOlUw/UbLG7bwnt
4jQtNYUCBKtDudewqsIW7nZ33mluQ/a9sD0ONErNeuL/k2I3U0uEXHUcndZsW2+DcpOcDaFaG8Hh
wRwzjkI5Ou57oiUbxB/aWtnH5TlOXOBJ29UXsvZW29nYHtpipMbSXLs60hMT7JuGvobE78888l5u
6jXKVJUYrcouErRFnpHhdR6ZnVFCWDTs5wt9g2xeklsKxzoinBV7tpHpATGOyKmuHiSUzJNRmR/a
coo+KIGi7iDlvE1jNhSBlI8LxtZDsc8cgRTTIcAp2FlSApEOc3glBBE6vZSgEMYmHyMCB+C1vk+W
VgddkjRpM++ToFSE0phtAYETTDDWV9ZDKM+yJnMGVQlkETtTnMW0zFtuMNpCnj9/ozFbjxhxkcCK
aYEIhdA/L/8o9sU6EnHwKBwSx0cUEa2gq+4/TxlIDWoxJQGQp0AkAEAaDopwab3OpOmwsUfrXdxO
oSPg1D5iac8fLt1xQeSXKbmMkTUEW/GJ2KP5uMJX+Wx6kWAUAnuLo6eUlywCv0tduvB4mvUpSagQ
5RLANha8OB9OJbDZwN8XUZ7jCSoWrrhqQzDgbWnoKXOPSiYJ1zAnKuMzWQ5ev13H5m2eTAE0gmVR
tAh5uQpXu9q4anhKlo/6sc9i2NtdmexoN6jQh14ibkDlzcsg6acNyG2VrClnFcVQltNFJkZSDL3I
dfrp7wCs5sOyHFdX3uALNASCe3qX9bzfQM1ncA3L1UZU54db3FL+/iEweTgN5go8Yhp3mrfNsrfO
qTvYjMNpWvUlc6Kpp2P+ONq9GlsTXNdlluy9OKVb0NaON8BKG/DYZ1o2FXsHCWKOVQRUURPPLWa4
46PkzV1mFBzmq41sVAfpST0CT/Lb/foljVh6dP0tY8RXcOhP6R2SnKHSJ9NQauZ/fmtg9pf0IYrC
cqdvL4JDSV/hHZhlL0XZBrSRDpBDlZu/R+FA6T/oiEroOkuxybSInQue1OrVh0dZLxx/GcmdUP9Z
/7k1LRSGDX9aDqYQMApHZ6KA7g8VSuUmxEGom/2i31xDzWe3G2y5jWZ6m998gzh3/WcAwcuPDFnp
eNIcWhV1AWsxY+3V4Ki6yKNH1L5NDE9T1aUb4heFWch3WjXbXQQ10k0x4woGBvukrYpTidsjTiXN
ivXuxiDWvcKEGBG8i829mKKdTpsSwWK0eHZy7PdS/21Q/ZFBk084UaHsvVqQ/ofMMn1j3IXZk8bc
hpoy0aax5puR3wGk6klLx59AgDYTm8S3JCpjUhX0coZcpYF43LxJyYS7gD3+agxiDL+CyqzJSAjG
dY6cZEvr7WF2rZO7ML90xLCuV8YF439CRpK57/7jEIYBLuVUbSng6p9/X4wJEPRfkCvAxgv4I5HN
iam/Sdi9pO8m9jkQLYVPsSysdDJK7oL2kHNyh56efz4XLxuPY4v0zL1GZsfaM8cy/5ooqBLHKN5e
XC2v595fWlHnIWkhHpjBxJBI4URjk37F4Dv1pMrWYBcfgzbW36RvQrY9JPkbzzAQplQkknr0RkaX
yE2IP3yXECxymdtD3Xl2+QwnAulTEhPzgvSOBCyaZ5Fd7qwGHsjVkPHUD92if/FM5MKgtE+8wVmr
p1NB37DdeDImItcXrdzZAX2NfDptmqU8tstu6F60mj5wpAgSR+WIdJDxYFROnfA18DERn5VVWK3Q
ThOC63jbl5FlzQ+6tQgKTwoz6cn7mWyrl9NhfeMcMoOZxt/7H7/TFUI+BATQysjkU4M9ejDa4fnE
c7vAGkebOEffL07hii/sGs/f+EWXDsEjbY9r2TDEX1qlzXxG/5KMXaxNFdB2SZRNzQHDyRvmBj5M
YI2GDDEcP6pyO9gUDYOfjfkBR9R0RCz3LeY+suFh0dolp7m+Kcs0cpZ+K51/0QV8+y69+ue0GrDs
HwJK/VUNRbD+9g5zgm8LiEMA6FWNftcHIXnQuyE2NGly5ukEBwOeqF1FzwWtHSveiL9lbwTEBF1d
hZeTwnCA2POZjJLRBME4YfxKQcPQwbNf4lDoTfdSrhjdX6wCFIM7uk4gyk4KL5bwMpYPaQTmy5QO
VoXWM0IAAkS7fipNiMXabp2CqyA0dQ7SzKgjuxzaj+0TLXyB4DpwA2Di5pE8CxFJvXvDcFuxVny0
LLL/pvlOJwYEQXZ/VHMnBg10OnAtec+/X6P1xiKockR1IQLTHEn2jnxVALvgVv4xW17xkgjFJcj9
Pdtt9LoqS58/aOaqdvdzyn1TW8NibL1TJSUGbBoP6bZavtoiuxOmA15p/FziWMgCoRLLZWFnTE20
f4II0ZWKfbGzloW4/1U6bTCFqIivQGKBRahxQjghUN3A1VlJ2hUls58VsKOoaXfUqLqA50hh4slZ
N6oPLtEz71ICvqjwdElBkpXfokss1CFjd/Yt3/HVhijnJYLA9srhnS7DvYGb8NGXVvCFPvtmyC6n
kCvJ7426A9B0mIwtlylMsDuJou6TwghIoEivnsZyGlhD49b8upHHOPI7Nz0NuHrlqMIpSDCvSOih
gwc9GZ/xyaFygN7c4LKahWUTAcSoR7kONeqJ6gBPwUF6t70PpxnqwzQND9ZMjc3t36lEZNoaLMUA
L/URVt1EFw39w6Hi0oBn5+gVGYIuPRfHsapN/fMyNnZhXQpPvC2rn6wJzL7VxQ3NqhMxmxGjUqve
YDWiFNQspHcYkCIkrJzb3r09od2ekDJoaNv5KZt1hmx4Y8P5Zl+4om270Ng9qLLZDSOX99kNXRZd
qUQqMF5pColxjDPztcqRIX6diE3Oazf++gOhH5k0HV7Qp8V//wqM9b4rJJknjQrzE+Fpn+h52UhF
vOnlIves6B9V+s6AhFAJQaKrrxxpsMyKVuzyRjJoWdKUj+p5lYklKeLRN1mcdU0roYRdSrWP7Xg4
irwb/wpqwJjfVwXCqQy8gXJVO4hRFM+OZtzVZT08HAgWPeNRelAlNP/nQzQowUuwdetBzPwCfZjO
bZvp83Ur9TbytHKDuVKvX/3KO4sDGeil29XzNTGiNXC4OW5mULTTQcyPPh6mi8/aNPvo75Wb8wfp
tVEj09h1gBIEedsMOqKQaaPyHQmq6nonr7CeCml8bLPI70VSSHWiVLZXPCREGv/xxjljmPn2GjA3
e+qs9GznWY/9MZp/A7oA9Z7QrfNMWBS0LJIVdnOo28QhJIYKfZ0hVwl2goiXjRspbozWCoWhY+I5
mKVv6Zm0lessZnLF/EBcuzHvLy69g4QOzp6DUda6BQ2iBrOVDRsUxPPYr2AwFiFvyetOi79T6yVj
j0Gm+x9xLGf+ZdGZlzeKkbpHYUiidr4F30m5zsTaprIJrsEauwldhDMAkVz47N2MG4ZXUdxWe6j9
aiOsi2WE6PstUMLaiEXkzKSikKzH4/Q+tI4AgeZfXGGwGJMSgfSR3rJYqxU3dLdOajP3aBk/pU3n
Lbsd9T9ja2XC71zhwlc5h6bKvDWeM49jC8sWVrlzVmAs1Dpmeq1ULxKzGBP6s70Ket5hfG9Y213U
nDDW13RYZcJXSELRkkL58+Dkg7/v5APi5VYfzTb/WXsJeaRsD2C3HEfvozbbRUJ20UA5DwJj/VUu
aWw542MeogtXRRML55i9R8A/7Zm1MP2FOvYTV/3Hp9BCHVQEUmNSEVCxMM1FkwQzOpTD5g1isIZI
dkbFbEfmh28u/7Cygt1z2wf8HYPy+iuycGqwjbVGXdoeMy1Qgi/hw9uzFQa58LSUJrAw0ugHjhEQ
O/y1KPx72liS4uOhlADozTFJL4dXdF4U+u5/93RBwldGCnwThW4irQ+Ty3/nFx1o+VPTWgBzmdsr
0DowyZXDUt6IGDY1zZaIEoJRU5Iud7tGXKA2Nn/l9kmzgYiZJ66MmJetClupMDXmxVr/neT71VzA
QwjCf4VvHr4nk5bFiTsLKonQv91Xo0uRoqsOg+LBB1L8LbhNWRwEYmUrGYiVKrNHVQK53EWuyHMj
kT2vRSywkOVtuhxngDHM5ogLr5meipFwUne6ofwt0BBxbXTdXStirdlNK63rmzh+13sxGXc9k6Tv
9RyozN5CQznm3JjocF82YQsKOcNONNdi3CCtQY3sfwjZbkd6vhrZjY69+7Z+F+BnFXxaIawPNZok
g5UzIb2/LiG+n0Z2qJh9YfjawUXb4KOBK41WvbkRXbRJi0nTreor/lTvPgPXoxTEcADAISDZ6CJc
71zg1DbAhCnBqWaLMDvIHWZImW+DZB2XlzSRb7o4n9REH+TLy3I9PGEIDseJDBRxIxj4MNOYftIr
Au9+NLUkLMW46CgXa6msTafZW5oQi+K1Qwb10IDmrTuNTcp32ZMG3cCrLRHhNZz7pWBLhczGcEWh
x7fNsMII8EAwfFZafgOtyCpk9O8KRneEMlTMRb+gzWZdDJPvRFMKd9Qi6RquChxoVSsDcjmd2htw
Epm8boiaJaU17vGe3tqrvjWrIVkJhdmzbRBQCu+3rHXN80l3nwOlJD4N9EoT0x0bZcpKFisGpe8/
EG31X5pW5hr1tIK/2YMUttNnTJupcl6XHBXJK49xCHqACeq92qzc5gpmoPRMj71hXLOzacujl4Ez
g2N9x+qwh2kLbg9Gyhk6S+ZXDX+3UKVGhxTOGBd3w1rdQqzeaNLl5dfRcKGR4EG1ehoNrqCg6tnk
NjlKqnBL98JMxKUgFYEGmKKw6Cq3Y43EQmR2NKV1iLB3CeZZiwg4MPXVo42wWmWGoP7/2BTmo8TL
oFtv4gtl20RVAh5mjtcuLazLAPtUskxQvcWGE6gONx/TCx2T97IM9oyTyZCvh6HxUaf3vep4Ghsw
eg+5LwuMErcxz0WOqSoxY3w2SL26IM73bPIznaSxHN/g5JlX7KcEH7ayIJZMsPVNF1dzWT4dVEf6
dSvg0fNBDvTKmkxvcA70XNBfWdcaVCbMfuvF5QM9GOwQ+ZJdjMZmBIOz8TcDZ5rN1cRlgIg2EsH9
fpGanTZFgzRHp8lQkcowXKpvfCXO2RxdLlrVfhRT2RpxigJa1hbr1NZPJGuZHH0kF7VNfJ5zda0S
P99eB0GrSCejW6Vl2vvQ0ScHiG+Rm+huFaJo95UWOopmFVbHB8GkgQ6oOZxHsukxNQWmP3RaL9nr
z8BWfnG6hXXAW8Uvr0sdKOwx7xeVUDo9c0ahLAjc642+GJsjq535SdhJmHe4PtVdsJ+mZJr9R22b
lyI8JrOYojJcR5xwhcb7enANN5MLSOdw8be6wFE9gCwD5qIUBV6u/r9Dj286NIz1pfYy+bIP+hsl
PoxIfu7YXtS24BybW1In4go8hf8LKySlNfEeYOJcgSgEOQsFOeeldC8Pr+oYuKlUvj3y5iXXCwyR
UxBE0eOq6oe6lnKzmI9t7jI7n0VRVFrVN6ktS4H7kwEhFuWFNJUHWvRwka5AaJdOcguhjuJaKuM/
FftufYC/YZjZN7QUg8VgOgEaodp5WEio1cknzymVeeMf7iqsSI9uOMnU7iO4zDQjFg6USulXbuq/
Tr1BuHJKOSjhNaQKbhPFoqxxm5n66IkSFGCpOB/jrmIarRRtmH4bJTlFgahK3axhtbu9u43GU7Ci
Ep74WoEfwCEj3KLMXkxKslCLfeg14KIWa8K9Xr0RpFWeILdC1U7Pli/DoGs8Np0gVXyllkPV6Usn
42eXlZADzTdzmToFVhHtY0XT6V1hMRILypCmQ8YHOQD4p2g5dAOVa15POvjymjVdSespaFSrs5qV
fuNY4ChLbX87jF/LoV4VdEs846fml4ZdABx43htuA/3Ud/CgJyolcMVqII43DJEQVHkTvsdml4F+
1BNpFhuuPzUjShxN+2NWhwTyefI5wh+cnmlO7jD++LO5SxaGFF/jjcfAb4qXGxLNCf5Rcctl3tjJ
SwHl68LyVE44Z/HV35ryxwSANGOH8MIfEetbmamy87LNb96c2m+t/gc8GHs8HJf9gGHoLTHWvmvn
Tw4chVfMXxDEtn3kfYFuDzDVme9u9RLHPGgWSxtQ7zHfOr68/aCSCA4OCP3gafOAmPI3dcsSgrVp
uwLiQyj9cB0Ehl/PT7A97t7AFAeqOYeoQ2nhM1ZVDd0jVZgbQpYhxIUFqxMrh/HNslgZXIgonWiK
9XPunw7irl5Ni8RkbbjEdTZjzSwZHa0eL8Fgyd2bG2gHn+fytPxRs9krOH+zEWanI9YqVoN5HLC5
TNoQx6Of6zI2qdKwsuQFAr04OTC0YKKvdpEy9n4gnCgWOLal5owSb+4gw13WkGJ2FLJjyzRmUn5K
dD9m7+xp//AIhsNQM73qI41JK9bPMoJ27SmhJrRRpIRaWR3aorpVX095Zqf181hmAhV1CheAE56m
hoQ8TUJmj3/fjD005ySKyR/FAoZ7Z2zpiXn6Rq1vaXoczWq3owLOW+GJOL4n7uDwsewdXz5bHM09
tRFTuT1NbNKFBjgeq7vxwCoX81Gc45wFVZD8pwIwanVlkQ8AdgVSJOvowiNt0N59q1Yh6C2WGxgi
PoaXB2ajNhuko0bGsWWTlRIE6V5BZJ1Cz3U/aKjhnBe8cl3G8sHB84AdrnfzRX7OxXKR9g0oMQ+h
dOe/tz4veiG1A5bul4jZQ/+5FfZ6iW2/VEYlslylDRXzezbFxv+Z3qhSidUQSxzjiVHxFNYuE9XQ
nyrb/MJeJD/c7YeTb8bIN5qiH3g9vcGcXQ7oyeQ7y6tS/IKMhaUVuS2w9ghJUOvFssZ509FST9eA
jpad3I6bHPdZ/ZdY0Nu9CWhjwvLxAjNLdBZCifKzJn5JT7X6lNhFUs1wNpw7QlLqxXIq/hMicj0N
33bFseK4IF06NJM/R4rqFXzAo/vZqyT9PiEQJA2686P+UGwerfbhvfq0lE31N2SPlyIhGYfo5AnK
zUEquh7YgRTySFvMVoza45sQKer2fHpDnw068EgmqfKkeOhUPb/XwD2CXhFwcuKtv+TlOAV/kGz4
NZYkeF0yqlsWpFtc7jkQFjtpI3qOf6R5nXHmWcj1cN4YN68qWdTtNsm9fTDgmbaq/uK8jsfPv3d2
3Gwem57OE5IMUn/L23F3WSQaePkPFF/ioHg8bJoJnC4Hd0skuXX9OLhDzf88qq76/7QWWD42vnJg
Ut6LgzFMiq/yiNz4pXBZBHHdSHjbqiGVR8Q6Y5YFutZoLGuXne/eZwxx1SMEGfMvmp3/MaBWayvQ
a+EFwzmC8CEBvCguEm8sXljpg5lkG5tsncaH/b8d/UXejwryhZR4VQA9v1WI4lRgxwBmBFwhzZKa
pd8NpX6ekqdaJRIWNwcy+bNW5QE1UPU2CswBqTSORVLo3noty2HeM6dv7w3AAmrG3FkXbQO9W1rg
2wxpRqZnqOULhamt7IFIhc19r/Hoek+7Xg139qdHGaySekuaSqldNOTQ4hgstM8snt+AWxsGyB3s
Y3psxFgjlzB/ZwLJWSC2wVh4FzbX/8gEXobYfvf6q5l5ZesWJW+UdWi31RcO21wfhNQOsu+Ly9y8
n+H/dsIRzkXbCgaIXq0xPlJuBQZGTgxjPM5R1m7t24hmcOUNghOdJPcQ+dZmW92QNVAEjHkJ5Vub
af9bUdbU5L5zRwtnyRSHi0aWffbiMyTkKdR5lVtxrSS+CPI5PYTrmrB52fkSPf5aM4Q1bB6DT1JP
iRkDNuYGdeWMBJSLUYjyP/dShcfURc5WG2Tg0Uw9X3q6t/I/oWNNkisXUi9bhXCjSrzoutistYkN
y/yochQIWqzSgWmt30F2C/KAXnfCXYFulK6pqcOC7pF2ha2xV9/dblgSZ5mcn/mgDjNLQ+LEpaHR
/I3rPxZcUZ5/edLIk5W3iLcUatn5pS9XTadEF589Svso2TUEtmbjCviA7PB42aXQoQQmRBjbnpgb
zW1nvr+WoJcW1XdHkIF2aMN9Oi6yS4gSOH1VNawRfH0mNJUPQ9hy46SUJXjIAelBh33f2WiTzcSf
aavW9Ixfnh4NGIf04Oy5VryerG+PO4AQPVmbaXy+bj1WfqvRKFul8VqZOg1wlLuMe8hYRbKJ70ah
KRIqT++eKga4RDPO/JMoIwuOh9vqPZJZzmNQWfSqZPax6tqtd2Hq6gXocjk2fG3m+T3wYXMIg0mN
uGN+PXhind4pGztZly7/KV+RE+zY4kvijPJK9ZXfUFbSQC1Zya0FzDYJD/8ZfZLU+LfmSgTYonoY
HsantuooE+HY9IMTVydBE4VIIywYqHTfe1H0ALKI037/zudZiwUu5VrBvlrbfRugvYpTdeygeZlb
VMSOQwe9BxPR6NPM9XzL461R+v4SzUzuXM7B+NUtbov2P2h0FiWF3hF0KoryWe7RJO5g83IW0akh
XYTa4rHBTAn05orbZA1B+srBNBpp8ng4RBkySG6a8qSA76E+YxsP/BhP1j6pg6bohNWpGYXx4L3F
KVUa5ZPv+UXcHlFFIe92oROcOL6DYFXtOikZ5rGEwgP2m1lvac0W5lKTWMw69HUISZ+sY1hAvj/p
AbSgm73STcSgeBSlqtANap6AIfvtYz21wVYPlcIDxgdPNMIDC43bh52FYlrDwOozSCgLomT0xf+m
ZnL/NOoxL++D9fuWWLJ/lyvwAA2SBXdx2dw366vXIX0ot5RqZYCIlCNincbHfuow+JDYoHex4cMk
66aH6fMpS6AqJjYt/Elz9Cw2j1DanV7T/0zmidFJb2IELQM4UI0u7tiXyec4ZRsqClsE4QfYcgsw
ktl5ZfRdkN72i1as69vbks11Gu1zIG1Dc5NTYdWnRRK2tvVZw6CSn5+r82XWok7TKmwPvicZWL+4
xz0MkAF5ceh80rn3ityGhrBSDGSRioAfcMRh5XBzN1GYNPZ5f6deKeUgT/M44GmLS5Wxyph69f4a
DQ6NJz/AbGeEByLdO25Tz08xuWjdv6jqSH9DDGjqfAx583BuGkRVhu+Lw8aFzZ+Szl8fHYiWmk+l
/AK9E9MtDisqflisaY8OaJCIOnrBf5O+IV6mKz7N3H35w+ESYzWOsdUJEXyQSMXmUfQ1/fHNEl19
LxnDcdifIDUwj4+zzK1YYZIh7y9cpxmBBKDZ+XX2zL/pLPofbOlDSP+/WJNZKGm+xV58a/GUm1f8
4DPP+/2kZU9iXhHFIXqpvcTBhNPsivx3nt1G1JOLzpp4VpjfjMbBdhpSg0BfxuIqM2BCHMMfKAAq
ivGvUhdI4CKklxUSyKsQ0haDp1JhuzHofIkJCxqIEXtGcTFBdAMQUPejgDOlQvuemDQ8837GXr5i
nLeJI8g/XTc/n8ADq803bU+rKdHri0tTkLrLuE2AmreC2rCC386D0S+fKV929wVfec7VPwFLGqSr
Le+94+K3JRnsSDTBK3r/qh5b196TjQUuY0mAtLYxRM5yQZyVfQHcSW7YR6G3snsygoIT7YoyQDNB
pjcOFMjgy/XwGWAWKVMQdEmpp9jLYRxGFxRjuRkkMVVyoqdRzCufizUJcnqVF5vxjrsBcXKbGzt2
rACv9Q3d+78OH7zsj4W5hN8WmZdFHrGMGV52ZYojtCwSIVZMW+LLuRRP7ds+j/Wr01Wer+nCFLqA
Tv9kxYeIfTKGI3LTUPWxT4QDUmVyX6gycs4ho3N7rhAU2dWF0oI6IfqsQa1GFT3n4i3d1yKlL8g5
XdNVzDm3c2k/HluqBTO4JcxxR8MF5jGDslC67nrYP9wbutfH58deDO1qRiPI5IRaj4u7NHIGfqQT
OSgtABBiOuZBVzoLnN1e9khWzPgkoV2cLHXuVtZCRgrulz2qB2ZsPxJY126TYylIpTfVgCsaqg6C
6hApGY6Pl1v5RuE52zJw2sGSsJmrL8BHYu6XvTTDsM2HQASVVSh80QE1MayXtqCBnar2O/1J7QUY
uoG0Glqd89haeTkpMCulpwyqNPTR64q9yB/YGPSLbht5NMr5dh6Fi1z4I+ZrXqJwO2LXM+mUzo+I
K0OUqG/BlMYcZGLjCn2mMsCkOpHNwljSGdF6zSvndr09Fm44BmEkJXD/fVAuP8HGkOgA9QyID1uZ
ryfVnqbeI97sBTWQ/1U2BSy4J3wW07vvrxM39YenzDelSPC6233mR8BBGN7Wnlj1mV6ybSuxl8Qa
qaHsBMl5HV2WF4PpKSChbw/lmcegred8dfvUq5zNe4zMgx2Jcv5E+wja92D5rCrzcNf3xdKXgHcQ
jTUdvVP770jG/pUIa41NDzbZLAIMG7uP4dYPHr7eu6YL3zf/tMSm3AmHo0lG8bViCSdR30DmL9YC
IdkjvWciq/SrW5r4VVm21U9w4YqbFuCly/X8cYo1mjrp6p0HmHQEWW0MKQH5vNMXyng6NGOklwks
fxJ+kuCkNcmNdPiT2SE01KD+y3eArDuj+b0ZqEx7AcaDFjO4tWIMwvDEVD4rXce1b6pEdJfS4N6v
zu9GpLm03/xsXBYSmT9qeLqGWmk8LZnVbbXReD7UMJBjq+qkaxrMtloqwsbekfxk6hScfi9IV7zB
+aisZphG5Z9/LyZpF21OJM0WDNCtjkYXZRHZ1AYlQdvTmiLv93PU/tsu3+TO3GgfvltaapiFZwlu
CpSDp+8XyYZmfgtpyk/lob0dLwhs0QgihfMNvHEXb8YpIwStxtF8gTUjXDTHSvRhbZN5GCQX49Ku
wGv17CbVALwRyKRuN8h3HLqZDjFavx8qzRlFFqX0srFT8COpRRjW4NZPtcRYH7z2e0a19IP71pb0
4ewOXmDDXRGLDHHFd2fvYz85QHmtc/PBeIg2Y37PTUvDiwP5NcTJ6+uE47cJjQVpy8/O47O+GtUA
WZy1KSKvqKfZkM/tDtI3oQh0BLh0raA7/MryQuEdE6Xya3+cCKWfrh4v6u+KieggEgHcKwI1E6Cf
Fe3aYmGC+v6bX+WzdroPae/xeFIpDLX9QjZLJ97nZ+7Lt0D4J0+iz33OwhNTCc6yyggg/Gfkk8GH
PN2IO2FPPJ+Nv6CEsOkp6B7+rev/HkCkhlnmn76S/xm05zN7lHrqVtWL9zNb0E6N3UWq6zsWNrto
MN7bs0Ofca/IheYzPNW1LMT1jJII9JJ8fve5PnmjTXDBahRxyXUS9HXZGghCGntM7ROicTJTM2cT
zLlC3H5JcD+G7KbammiorZBXSTsgZ6hByCuFZeNab5mYKCHTZUv+UlBlv4cATDyXn3B+FHUJ1hJr
o0d9lwJXMPSve2uCacrWzxy6Vaoucnr1x9hZKQMn3A8xuQ/DyvDGz8nBUqk5b+0vLz3O0rr+1+o8
L8XNiJU600jTGEL0A2aB4dS/mBCUNBg1ZRtYzWZkN3pyreIeCuzfJRSMnGFnQGm1ZfpD4BPCt7/j
1VY0zKTuHABTd74QCvZ2vyoqC8AzB5LD5BQ4ayWg861xNlnlf6puRadhXSVYbk973AZXrmvuAbFg
lQfZWVoiuhQe6ExJtkWt6Q55U3/sRmVCvkpxq/l+o0gfCETaNlt1wou7qiLElRxoZx7R3uVRGsLq
lcOhk6MnQABuN41rqH4ioWN0PV0Sb4frB76JVsspI/se07eJtHE8Kq8EUfBmlRtnTSgHcelerR1v
CakfbMfj/O2RxEq/y6GE7gahWNhiV1aBPZv+cA5B6MNKPLtrmy9IeQE2rTmo/zsOlcrlVXsTUvR+
Pq6f/yDWoReBeb6JB45nGqVPqEV58sUsdWphVBTlJ+05nY3lp5zcJam5FbLoJiSrVhigN6A50cYt
j2q6XDBabug38AT5iSiEVM4Ob7c6zmSAZunNVRDDhlx1qmp47cWmP5Z1MLMlxTEYoz5fpp39hfUr
W7B7puePvY6BUAx9SJ8+8+1sS9OMLLGIUD8KfyzsHNJrMW1AlsgnEhNUVE8ByIDYXns2c/0dnNRx
XThNSN1QpKmZfQEXK4ai+7njWYJBCLQ2Op1iKIlgenHlE15q1YTAzjRYf9h60uV6Ckzc7LscgD0V
KDCsjCpT9kw1qMT0/NEeQM2oDrh80MxL/fJ1tguS+LB/fYGO/+X/OrrqpOzQYkHG6bOPLNXgSwT8
Tud9Lw10y4DlDOyEBKlBPPPsqoAoPaB1g2S60nLwsTatoxtDrqq2AhIuGpagQDfyQWUXYs6Jq9a/
wm/XOCd7B0ijbN/sfuIns7M7rXsV5Qc2e5hN1cuq5lfc4ebMWv1Ib8NZ1vcT0yuaa+R0xqgx8Nfg
phgS7YRPjTQIQtX+RroYNQwgJ5ymwR+bvhFi1sg8NMZ3G7kPiztmqGQbFN4s6K4lQ5oXsrTliDE+
p43QCFkRCGiUEpxewTFqTMnOSCwjspY2CrfYN5/ei/nS/tzNeh8akIEPQ0BkGMxKkPqtuN991cji
VnExi9bs7fqGSN8sPok1TuyvBwPAi3eGDcoKCiU/S1tKcqyYlWbWbyk1VQDmtH7YlRXG1ohhvya0
+0e1ke7W72MIwps45suyi6NVWp9ltenTUpaGCe7SZ5tei4i7HRbDnTefekaDlqJ4axzMuOfQT9Wg
zx9GuH52HRUYTjA4qtj/tFf+Z6udlgHTBEUq3p8Jyc0QnEEN+OY0s6vuZ/Id9FGK5A6IPgILo/w9
x11VomEuaFiMhTBwBPrZAQsN57fEw07Sl2+Mt2NwS+kxCwmqZt9MtNEuzdWpsaY31VTCN+Xvqv2c
1hK9r5YnYqhlD/+wXNDSs+v+F8na9Xj2oFkSmaK6RbXea+MUN5vDfULaOdGruYQUe0layMSTjeNM
dGvJTpXb+tJDT0VDgXuO0xfb/i5Ghr5uPy0wPluhl+yX3K2F2+Gj0URNppWAVqgerDkdvplAwhxt
04JCvRQvZMiUsRGM30B/8wsalnopcEKi6yfRaxWIXy2VV/A3Xl/7YTgsORX/M1FBucJrqwcdkFLs
X/5udTzarkWjG16it/Cyi94t5JU5O+Msv8NSANryZMxx23jz4ZIX+gT07LyFOdkbFks/HPGIEye5
Z/qDnXzfh29xUA3BROl/i/gkAMzshTh1YoSwDAO+Sw5dTly/M1gdcZM8g88DSgYa0qC8ZXDjPyC6
CPgJW4j69YQmg3DnJwKGCDYF6yPobY5ny6+AsuYRi1W4Cntk85frlTwsKYNZKf+ybpJJzHkVBJKW
19twVhTPGPNke57KQmSq58AN0SAMwqtt/MQYVnNriI13CsyHr+bkngWaDzZZsxu39vxLdHnHN7Bm
Dd5kGjMRLf2J88DPFQVdVgmImQzbNX5C6jwm36CLrhQESlboRH7oBG3e5nr36oViq/8/gKTwEn9a
lmGjF2wAZ5f+CmY7xRegq1m8/2sIGYAsM60zNK/gzIikKngTCR9hzyb93Jqjb1XtuM/MYSSQddXK
hm3Ok2UAxYJv6YYA5oQ+6zbhOumkOVUpYQF/ywBGGNTSFCqHvHUAxrFgf5N1NOw06C5isG3Nrhi4
FZa8ZwAV1GAhud2+ppLsF6chp/TZhmUYRnsw5DBQ3VHZdutTPT65CglN07Dq12u0ol1bIjTIVtGY
1ygyj4mkgWgLC/taCdOOXd3c6li8mE2aJuSXECsHaj2wORAQmyVO+WNRJrDrcWQ6g1M1Ts7Q7B1+
EOu+M9KB/MA6TUHYwo4JNfMUp8ycjLZXcjKtFDUu1KHvhBgpaB7cnOlyd4/5l0mlfK0PhXa6+15V
XFX1VqoYm6vr+fNhhhY1hz76qx+9614c4fdnT7d3WtZKwYSmcunZeDk+tQ8KNtHEWv+3g1Hm0VLF
vcnxCfmQJDzKOOjHHa/zWOy2Y5mmBUTk3sdvduOfI97fd6embs8O+uoQG2SrwC7MtFwlw7mvfH7S
MIhAcsE3PaakJ+uPpMime0bCm/cJWUGjWBPIviR3bKZ1MNwMs+oScrO6KjG8rWLRkZwFhkdVTur9
aPRDymh5of2uQuoCu4lQ4RtlMTTxBi2ZiTmcstl5RCCaF7bF4tS/gxQiET6WvnSPCE/UcfFzYdU6
0Gd/T2ea/6Pa/gJB08WdTVtGaRehgvAzfj3vGzekAk6zXi95ahrQs/8dZoZ6XUjtOYaPz94BtqIx
D16iaBfJ0L2qIe6uyNUJwM2DoZ91yakSgoKZfU+vZU2GekgqKMOoWAZnvEImJ2WsbjLsC95/Q1vs
4AZxdhWakPTAp1aSoZYsxy5FQjwe3fZJgTTQI5y/WvRFic9PE+6HZZqIJGglJyefhCz71F7WA0h3
ihRu89Obhq5r3Ftm4Uvby3x86BVYSc8RrKFbgjQI+HIdbPS9m6kpB+Z+XedtzQbeJzqDV3r60xl7
pLffK1zyCw609SOhYCM1yNbFCbC34miRUs+mQl374iFYxTmSKUGlWFP5pbXCmALacHrzDKMaIW8b
6/PFY4fcc1qf+Vv8jDkPGjsHcK+/HVM4G+QFcYmk+ARc1kVVUEUSfTSunQ108INjA705sEzy36Ja
PLuuKfyzqVNsSttOC/PXgrUQiaR7o0SerPJ81KN4s7GLH26P5LDLyhEWb/3sZrmLiLwsxexc3Ag3
Ae36xJ99KCDQ7LGuK3XMim+guimsTcQgvSSYo8I4MH136SYt+78mT5k1eEPY4FvMWG9RbpDaUeSC
ibYMVTfnmXnDKBwF6ykGaG/8319r3dqMfb+44FkdSqekq4XjT+NViw0SFe43uetxHkfoMLcKGX1+
rGbcl5mRtIKZgsi2MJX8vvmcVLhmHts4XgqIvtxQfAXKfvTsLgtkqmf1gPUSLDGxIGiub0wahOFh
PPBYYYjyQMfNO3DbPGHaPeA+rmWyt7I1YpSeR5pwDaRMXzku74fgd9fmu/CrwW1Kjg0Z/fNsThZN
M0JaqTTud32hjpdfcGEEmrdfM0qAqNwlEYcjvZPXfYLebv+G9qFqwByPufm16w9aL0wOrCpZf0hW
w8jVLDkNctkkeUjl7LHDYs/3ACqIucitvmyfkA/jlI6md5sOGA0QUJtxXSqSCg0qTNcYx12AZJK0
qPIUun1BU4Rd9tdcgEUBvbzu5JO/lX77ehJ+SkJ5fZjaPuARZvsep7Xjrx4XnvMnHkP9DHq2HE2j
NHrnndpu6T4lwzXmbTEepbajTJ7us+EDIblvEe1MGwlEPMa5mUmiTza9zzfxjjEouE8owEcnDjcD
89L4sqGKzk97bbALBaOQtOPP5d6d1sdqVd9weqgyef0mNbXKedgGqH+8Dyg10vOI3dYRo9ncE3SE
3r7Ktq6ceY1wts1xJALS5N6RQJjbHlGFGiHR0KckovMOgiHVe3rSnJGViNv7v1KeJubkAfgL5pNx
4ewUAESANtU6QKCcCPz9bb6f5eEAeCcuW7FBigxZe2flwpt9Qn+WMqj6Ksvp9IdKfqTjvVlZ3sCS
3RPTi10ajzkUcIfB0tbIuu1YDD221Me8fmnMfeA4tWyXIHGKCf3jJwhfuqKVRhxN/86jK2YrlgCh
ngytWF0JoQ5c/xEv+DQ/ZwmbXI2dwBbAH33jEfwrEEUknJLcfPpTNK9bqrMSLLKCrSWJuERVZ8gS
MhvkcNaNLz5p1qZWWRxz/Fn0Rn7+SKfuJW2aWZR5VB7FLiJnLCz+aw/zb1wfT8hF/21+OA8mZ5f7
kYk8TQGZm7H3ZJIlWjax6z0VXgeTbPKBU5il+KIo5tfKAcMfv5fnpV9TuY0zTqnzNA9p8GPlqncY
xQ6B4v5SnMTI182jDWLzNASWQ7AqWkeoioMoXjQeURXayA3jx3rz9QkMz2lM4CZeguDIEIyFkcny
FEWmGsdpi92vBEkMVdz8aW+llviD8J4Sgv1Q0IqFA+hvP2/xlfH+BrnKyCyr5ip7pxx6tr4T726i
S1tbEC5iVxf+s16Uln9jxsTt9YfFmZrwDisUx6zoGE2CTH1TpKxsEEKbpeIyIeMXJuxrZlSxS7wm
lLj/ZjToEVM5gXw+G7A/E3C11cymRo/m+VR/aQSoNBYL9O3DW4XxXdtNSDdL2l4AWAl48yYgiRx6
kqcKvwa0saPMY5OsnkDuWpoURFBSqQ54pm5EEeWE14U+iYj9lwv/dfPH7f7qmE3OD4ETdfgMqpmt
MgC7KyX2HlzJeeTdo4fkU7WzRoEk+zH5EjB6QW8FBL5ftFvNLdnYL3hqxdd21Z7qbTyJfIce+kFS
RCvc8DQ8hOc++xQ/yAQmRxStrTuB2U0eu9iE3Sf6yughl7JbXTMnqNXIUnPxkSXNca0qyR3JeLzc
LK2OPGEZYuhpb0O+JrZtmn8vW3MBZSND7zdHRtt7/KFDDPhOiuk/oRD81nXVGCUS+3cnBaNy+BZq
ZDVYmhgG0BQ9vbrpNTCG4UArT8j9OQGxag093Nry1yxuzrdajP9Jm0ex+Wchf7kqnsEQcqtgoD/q
wU6yw4d5oIkpq9oNRmAIn6I/FOfLbqr6uJipshZEzuYomaclLRyoCHSQzXJFFyx1CHcZJQpI9w0I
mC7aB/b7Vxbl9eOnT1xJGBgXp2Mz4Bm+9zsbOkOR14MX/4eBG4mHSzFnikSOWWij3ZnU+0Nt1Elc
ssi8LnAeSpmveDJYa7bD1jnFej7nVhMqr1foaA37PU4EyGL8bmOGypOu4TuezKY5Ms5kQEt6aYrN
pPviyFN0GhV54Aw83ML8/HXU3jVQ+To6RMCzREdDx0E/Dj/21kiHO30eZxZvCJEeZP51zwLz1A6U
rmxGH6U5H78eu1lLgqaPsY2MYiWASRQik/yiRbjM3Y+I98fpiHXRYMBUXicPqZOEkkERqrf2HGaQ
50u885RkQDmEIoVviDS8NycaHnlrg8nJOMdrN7wrmzKnvcTO0HyqoAQPaK7UcNGd31J3E9uWXbfo
5nQYIGs/rVLOKtV2x+nWkiJqdhDE1j+va85FFQevXulcjIQZ9rYZN+Zyo5obGrO8JXDl3EbxLR7O
H0Y4ZB4nC7JdDj89SVfG5Tus1l/pnixIXiWnq630c12aTuDdv+gMwEcNYyyKVGgHBbaYHvs6Z4g6
5p70vey0SVjNJ32sS7LpOtBQloRZQtn4Pt+Ng/hv7xGprGPNSAkw+GhKbrdiHwhOZJQ/8mODxxnH
fFIEHsioQxyekM8R/DkRQ/fhin1EkXR4XuBTAzK7I0FtCiTVkmVmGdfSgt4KyXzqhzG+4Izdg1mF
fesqZOTL8JpxMp2wazXVOi0lmkcVCpsY5J12DR+8O4m7Gbj0suoPDwQwiM+Xpm7Aw/uznc4/+Pho
g4TFOyIfRxQP9YheZ/M3bK5uj7bRqwD/vyPqqd1VsjFdlzd8xlp8KKBZnXE21IyOGAZI/EmLE145
m7so2iEDYS9KZ27BWSlBCGhNnjB4xrsViBETYmoeawfmHMBI9WtVFJ8BYYiJGnTcwqunw/Q6GoQ9
FI5vHxOJLhPz+maApwFR4L3pED1A3i4Ck8L5K5CTFFffBYz+ekwygAKhdzKWKr3C2Xapyrz0t27s
Bf8St0/n/SVMSaQhi3/hppZ4W5fbBCy5rEqiL0kXebfuaNvmRL3Rv8VaLw9yQoxEg1WzTzCqWR09
sL9TOgtCraOnNpITSA2hl4Tdo+tenDMHIVAxRKl4o3bsKUuJCZsgtnfXpbRDf09SQv1vGpVXjQkz
EmaQuQGAoYkcHOneghhkaewdSTyfXqxEPHW1PSGU8mJ6PIqV5RveEkQ37NyrkdF+9DtmmKrLCSSk
hC9CAqqkZGgr19ahoH4tq5BIOtl2WC23ZStXSRiCjHUAGYsCzPTihXG4NoHTcC96Hsgrs0BGA7Vs
OegI8EjMX6buDsNOMU+DqDL2vZfj6hON0bLUL1yS4FwyhGDND08moz3nDauQZnMxpJJcOTf/FLy9
5RMZpDWHVjgkJSg0XN9TRXDIiLRsZ0JHH4AwaOBgaSlR23eCPNUP+UjvLNz0mOExvYVHY8pRurMg
RWm+cZs+dxzNPXRk8tAFO8vaaHi0gLmLE+MzHNf8WBjusWfOalf3wiwR18RVGRxKc3rpy0Ggh98I
SohhAuAodKshAx1V2g/+OO4SrG5ns5yuyebyUzttCRAZelCdymGWs2gl0HmvXhragNNkihxnru5D
ZOh6J7bztfeGIUaMda+nkqml8II8u+8kzI+f27oXxAIkYtgW3efdh4PKtT2JZ2jrmwiefjm+AeT4
9klqeLpPQ38pR0kB+SUn8z1QEDW6dXodj8G1rD17ejWe6JfYhMdgVCjOFN80KlJ7uMOVy6Kgt1VI
/fNtEnXCkHDE1LfnyJl08LUn085AhAQdCKeOWF1D1vKv4Mg2ZAs1Y67VCCzaTscKtiTwxYkFtQOU
r1LE67DAPv3Nmuv9ycC49nb/HjhydJKHlt1WB6lXk0l6u3htrCL14zSzr0QRJwro0dOhdoa6cpcg
BLTS9FOLip8BCwXRTrznOxcnecIbQcU6wVp/OwFTYIKN1/9chkjGXDqsdZsLGSvWa/LtwgD19mav
3hi3hXsDZqjVcJ7Ix2590PY1Xh6A6Vx0WgajiHWM03O/tiCnN1Yb83hnF9aEmWUQWEXIjqBnqeCc
Jo/ImGv2COAjSBpl4w32C6IFpKBnDPgU1q3NLVa+hs3NHJENBvz+l3ZJXr9ud5v4EH1rnOcx4Av8
Osi3t5cOjfvIgJepjMaZl2TdkSL0XhD97mchzu9IQ0boJvwI4J0RYbogeY8lt6y+/cfZEsGx5jrX
dJkzQcnns4ADjcHijZMs16z3e17ne3ZMS+qyMJMLt0FQHiO+m16JeHEw7h+Yx2fESO4IjhUieyq1
hHWbb4HgeUi8fou4+9RfMUrjrHEgioUU1gRgTSeMMDPzHV17rsKOvVdzpPiQkkh6Mxb7ZFm8/u9K
Yu0C1TyrhqOFs3c2sku/iPXqgnSbidv1aVMoy4wLObkUv8ZV29dayjdouIAzaBMcFRZr5oVOrLOb
kVA4oK1YCJ9q2+75u8rB0CtOr2K5vzAUUOYMeiVQ8T+63IkMKNODRe1bk3nVjAIX1hcaETWZlpov
R69xqAYW5YZkO27LgzHZPXKumybswAmO68Y7VLB0GR9SpYqud08XqBdMpMDazlksv8iBUCHwe80a
Y8KigBjx9huglgxwB0q3aMZOkgfm2xF3Ta03fOyLtBHXDnEnrN6MlEDlBjZqAvSEikeDsTlVXy50
gTfNIBUn9UtlZXoUmCx+VzNm4E7/eN9S38ESIegv28DjKeusSiHAsa3ck+zjvDIKwA+hDr+XYXqW
il32dBjqSgFFjr2MTjIXxO91ngVnP3chzZm63HZfoT75hcVaz2TChfJa8/RkDJ5QKifQo+ydLum/
IoDfdsuyJtwbh6n5O8kxaqhi5V/Ko6bUhHKSX4m/6mn3X4J/VNyWthTzLFZyaVmFZeUP/0RXbgtb
ecpj7oew/rCdzPCFGBNXBAHWg2/X8Wd36WXtCcwVTvK3Y0u7T9B/UXtV+bcOaVqmXWTwWKF16fkN
TTKMeiHovQQzNc6Hfe1a0VtvM0AUf07x180rD+tWAt0LSowxldktZ39Fa+5sr8fbPUqgJ9lXy17E
VeZ8x0kv6MXqDXOlswrs6Ck0Y5KNAKYGZByI7drEM3x7/sbJnqWmpJJQGhPQPn616OMp3HVyG4gb
szhjn7x0BiQf+n1X2ZAfB+Ctt7OqmA5OjeznY8vQt+v8dDjA/3O4WgSiqMBSvnZb8aCJKhl4H3tt
7P8o3bVcBrJUW4UzT4am6xEU0Dq7NcNVK9tnIPZEJryE9hFzXSOlvlabDrUUQgbR0n15KZCVRX22
jN8WncSzL1Q5SNPhkY/X/7zTQXWdcUbgzIBN2KEzGd4QWsRXfVtALIOEu24OyEB9o8BlvzVM+Q8s
OejeVr1/dPVd7p/vnlfwN8cFuAA/P3okOHsVJqCQHU4gw7ZXkP5Yv0krogc3P1EQKD4jHJO9n6QG
pUJIuO5jsGCtiPYOQLfhlpGbxV2Mn6PKPrPHcDjpdVIQo2Rb82jU9o679lB76JzYaFLOJXVjbe60
WlIOQFrMDQKDEh0pO2xue+OrvpwPS52cLoxhj/b5DFKK06ptqaGZ3b9L2SHAggNjJhVIzNAxksSi
JpuU9h5UW3QnV1YVFGa/DKSQI8e8NP9Vvp/jWXyXA84u2ZWr/cHXCIJN99WETqWeNfq+EBl9jSL/
MdcmgQtkr8eldoSFmfsUB1psN4wL4HzEws6rpElVveM+hbFuQ8MtFZBRUESOGuGFaNHI2XDNvetS
8VUyaMunhsaz1Vv328AEG0UKJukbC5IjwAXm+wzBNXno1aqpuO9WxBiN+mblFtLptNmz5PmBf0hu
o9HZVQDzOo3ffFzkpJsfaat62Ht9ySSs7tHv8I6qb0P7YXmh30VICD+ZtfH06OxZWUA0vYCWryH2
Qi7bWjV/c/hA0JGWIKsQZZZGRsuLkDn1aF6hr0MCUsBAIJXGxJYG8ueLAzL8e20pdxBJEgGYDxuT
NKXPDkQO8ShMdb5i5+PI1HmuaNwa4IZGKy9hhYIfLoeKK8D0I/ojCvv9pJrMThdhryzBkVcQ5BDy
yV4JyEbX9WKQCru30s/pb4XXtM8OXe3A3RBiU3/XisyLnSXMZBWHCKNB2rjrdwr0tVXBAi+jPE/K
ouzzkzZsPs4da69GrVzQD/epdJ+xfhFvEtM2jrZy1X6HU4v/w7wqIanqdo8jvzMfu+wABR5cl8au
jMGBK1CDTRJO1HNOrE59miZXryfJjqFy/8Qv36pm/Uu1cBHI2RTKwIBp6x7h/DqR2Krp5BA+62d0
6scfuFOFUTr6rGvj2uDpJXhl1IXbA33M/0PIfJC1i0riNIPH7t9k0Jq8+avxDm1l1TRMpVQx0G+h
0PajGhniIpaLsg08XwyBe6Be660FpS6+JEHlWQi1afg+ahJlcm9rT0DqKfWqBgWpRk8twPU4CaXA
8p+JEPBdlNK7Z6r5wx3BV3wfPwDp7OHC2gi02AYfe/D/00IBdMh2MTsNY76Jkbgu8S7GTZH4XEHn
kA2caUW2dxhcugC47g5iRAGBK6C2E07SCzCDo9SjrdU8l6aevPNnkN6hu8QxKaRosJBu8bDxR8Jh
FG4NLRAQW5dg6jFJqiHs5H8122tMglX2DPt4QxlXxD8MVytnpVDHpG4gj3+Rj/1ioBadjvRIOED1
wOPCU4amjkPkUE4qi3Eb0/ys8ozEm5FCDVTU8yC13lf/SftDbrq/tLZdKay0d0GRc/jADgnlnkLU
t88kIfV/PYNIPYHOqKLrzSsWf9Rc0yd+jQuafNBv6s9Ydfr32C+0cQ5pFrWqu3Xp4DIjuB9IOQzn
Op2r9BI0frJ5QtmnuoAxQQB71AHCOUyKuv97FoyXm+KzK23UTvy8PtZzW+73lauf6E2JA5t8Up0U
ac4nZnNJiL4CgBce3zRyL7Nh2kGreRX9TwboAIG4s70aX24L7Slhy7YmEyB5jU1bPadjujGRvTsl
hRA7Y6dzARFIejBmc3r4ptyRD+FdG/WkjTwrZs60rgcWhvhm6a1mHypVoUbnP3V6EeReCmGLiUBc
bIRhJPqHwA/Zw8QXeqDV0Ctw+bGXI6BdWFAIzkh16lxfV+K09RJRmrb0xGnG/8HRMcJbVWBasK62
RYaQOYQaFrsEDBLb8ycOUeM3IAdL2/0Z/fB+jz96VQV5EmIaGKc9ZBV8qBe8gdLFlieN+a3qfd9y
EZ4IfyMR3ewDQQDatje2dlQO4LeNmy4rHk2JZstRiuLasCk2CnE02HU94q+ZDjy7SkTnJ3oCrXvk
3yvqCln+6eLSw4WV9QcUFlA4E34fH9nBzmhufDvtQ7jqcsEKQQEqhF7SE1JTiu86kEQwN5FMvk95
Ql1c2nGrBK7o4ypf98grNoV+zAxiWIWI0K8Vg/97PP3SgUtDlHfOA3hKiQjI78duzjpwFSRMbahs
p+CxRswMiewBT/p5QH55BRbeKivB8DyR/bCWKN9gJu9yG5RdEPvkyBGR4m0fzkcpCa4e+VxIsRxb
ljIucT1009fehBLAnWriIJ8C/TZyXqT1njGsCn2tpr0UDxP+KayZ+T+56uC2mJUwUem9ZoFVAeJ5
ORPNCLYcQ0AGHzAqyz7rftiSaG6qW9VFeOWlyxHh36r7pUmBHhBcxfFefL9/j1WzCTYuKX2gLRxW
sReNmoMrAis856bI4VhX/wuYCCN7s+Co5R9HJjQZKwr+1oFYOTlcg002bJHapzzNoNIH243dTOEg
M/mhb08tihVhsJWIwncyDcYIMy8W3nvfrqi6JvEXdL9KoF+VyaLp3wH1Pq8mrcyXFKV2bUbEW1/M
mtR2TUoyqraw/C4Gt5rEogEDHZKHIL/UIPXoPFk+z38xOxC+Pia2Qpw1vDbEK2A5ULecGraxLs9u
Wrb1cJjRa/s+SmlHKxI5WUgyaPcxBPuE2KRrIESOkf2D4YPQuOoEbIrd/W7OSQ0HHdYSdtWwjt+O
mLBAF9qGQBA0Rsc6vNx2/us1uqpZS8NSaT5dUFJ2NmcPrvaWbt3HwbUHIAIQdKQy8IAnqKp+8tvu
bu0ne8DeqtvJweV2G2QmamhciUcEV72VLMR2X6Zgjnbu+D7FpVUl5ThTmhIA9XeLmqKYn/Cuj75/
p33ZnIkqZk+Tl2mh7Rc5E9y3WQLyhQba3xjvyddKmDOEhztldoYra2HG5T0vza3XrLXm9g5GtKyF
CFSEbDFrx0d5NoVpN4jTmFYrurSJMap3IreNMG5s88hFnOPvDGBVAI1UYEZV34iuIw4TS637eb3E
4iDt0s4b1Nia04SDTdkw57xRgpn02dCMihXZ0V7sm14sNPWpR5TW/YGU9oHVPrSLcSzX6eNGOwYe
TJmH0h4UZgmlLJq4Sm0o2q5JL54LG/pcJYRKV7Dmwz/sGee5vwdPZpvjMUIHKMvLVi2pB0PVaEq0
6CXQmwRLj97cj4FqasSRVfHkgXHmxsUhYZyqJssTou2QJXln9fpqrWuC4uVSNJyh7afc4gzjq+G/
yCZv6+ipIQPlOoOWMmVX0HsLAXzuzDhN1z0h4XywXVolLkKhLtDGpXnaOVXYBjsglk4cgRfFsPmy
RpIFwX6BNwHUMrjoUlVG+Hi/ISiujZSg86K5gwKTdahN/yYvuYXoAYvmLv6k6FyXPFMMdsWAYKTr
PH7h0r+3AMJgI2f9ZS8/1teS4ozThybdGCM3E1M8QdiKvWKn5+ZE4PELPDnwGwEipGVa32FLtijI
OG3Bl8VCJ8rD7ZlvH55HpmZIkk8tLr+T9TlMKTQerMEphSZOWI50Zki0whYpHvpWY1FUUqcWMBEy
xiAQyUjHERS4N8Z2BBPWmXEcLxcvhpnJo6rSW9zbwLH1yURpM4tJx3mq7rUdm3gvIbQt4e6Kh1Fb
KqSBDwPMhpIftwJLP5Oo2BLN64PQOhAbwLODPaexa/0eppDGA2O6UmRX9hIf2liWwlK87B544EgT
4TQqa3eMexxEf+F+AfQOav2vhrgn6FwZ62fZLhh2VJnGNFQSCad2u3p6kWdi09rRuKiA6PEJvi8X
O1fElWS9Bt8xTRCAKB1OVPPqhK9Ve/d/Y1X0V2g84MkAaBI2V5hFuEi74kwodloDhTH6UGqPfgDo
zUn33nAB3Xa9dv0DuXIG5YYOlPyUdyNN/+vYNw1sa2iJ3jQgbHmD/62Ob3Y3xmzLHrJlxQMh1nFQ
X9Nr/ksE6oTejjQ5/Vl2pi+d84l5LecfvtOzm6qICGiQ3e4JzwAvJ6qKE2yBg3sZ0rPLDoP5lp+O
QblWLJOl9sVZVShmYhhmcVQC7DcjyX3rhHi2ozP0OfPOESub8ZLX6lhG2D9VRqg5KuEztIXDk7mE
CUYP8t5XUAftXRPX83/lQL+l9aDOrhgFRLh0/bCWJSk2NcdUtznVKNMjLs0aEquxeWbe3oU4G+Wk
Pa1EKxhJugrdFiJaL2FhnV1OPvNydn4pVB442xua6/ldaNjg2SNQm1Z5HMxzP7+dsXdfeDOAWLbt
BLrMG45lihm6XlAP/b1fuIFz4CnLFuinFYeXjokydYigLNORz7Agl3FARPW9ycxi5V3BguT/dR3L
UEbop/twXzTbKu/Qt1Ove075LsNOXnybuMx5ZuB8WZJMLl0wrtmk0FZhi4VajRmIucQKwlTa3TcK
ebDXk5evb8QTPT2ykDLSHCpDrL8TZSPh6w4OXZ5ZIZspZJS3UWq3Ugp9reggcm7Enwe/lgMIY/KM
r5DuhgR8JOl2RnysjaqfiL19hbdWtutwgR2mhHB2ihcsgJjN/o94JjiQM++H24cLF2dCGPbuzlJ3
jG+Tl5BMX0+ax+IIzz1giW1ywVkQAnsBNWK9H9rUd7FERIHSY853GZVXSP+7h+sixbOZl1wGuJwf
dBdnSR1GCWBZ1guWAneV1ns4NXmuwCU4iMwjrANJgqmqJni+xQhbjMZszAQRhH0PYXm4Mg5Sktiy
gI+Um0ALq8qZlyCi0isVll09e2CYKqMJHs3sCB5OxNLXlS/oRIeb/dQvPR+4wH6PxkxqvYWeaYwN
hjqre60gwGJdxjzgQdS1FyG2Vjg20+14xoc+RC9Q11Mbkc4jDvoOe1j4UNpniF0XJ+BZXjTl7za6
BO745quH8h1KXu5q13WQHd98j72R5TH85lwkEZP6j2bt+oExB9Abd9iNC6dIr/Qs2yxPJeW++mNr
5qskRmuKqrhjm/ek4BkYeK44fj0PYiZpmGIEWbfMHSDXi/XRG8tmjZJsMyOPBVEHZVBgAuMgGQ94
hsSFM6zG208tyMRdGAD703PqQ/HwophDhEveNV4iyoExflf9U1w5JU+7WUf5gvMFCKVHZ2zKwdYr
/DdV64AGSpQP9dd3MGP6YH9XD5McQHX2ph9lWwgaNvZlRYUMknYnalvyPrPxIR7x+KqPRpx+L/w3
oOXSPnSH82TBM0oMbxzJov/Y56HW1+I3HJZ0Ye930FAYWjxjHqMUa3cxAF6OIqOr17RdImwcXUiI
vpZBUmnB0iGwe3i845G+8l3On1k534I03ZowQusU00BNv/yJgQ8PZjxDiSI17ywUFUYAWe2GZSjt
53Ae8K+OK7J1FB5HwtMZui5tQZgoxjchaQm3tEmony8Z50Xl/eYqI5/vZp66kIUMcRkOY0qgqKmq
KoFw6OSMPm540zF8lUy/vHk7mgoNtr48sf79+CQaNheVHNHz8Vrp7sy8jtK0oH4pUvJ/hleQSVN2
4mczUnWkjvgSHAs9pgN6OZTd7baKhX3Aycq8yK7618LcO4ugrLV/4wcXDwfjL4FaiCdagsQVJFs6
bqAjraLeYZPRfryNHHbaP1rlGGNNQ6IZTHe9Q6sCE9D8KqUpnvw68fsyC7wcUZVDSpOnmbThoeSA
3oNfEde955n+VlKhmF8GyO8mc9nj92gKj7sqQwAhkKPKxSD/ymBTkH4C0pzYxjVs3q7WF/rTXz0C
juJJFvdFiBppC87eLWF125KiPWro9c2k1b7CfADpSukh/IprCPqOPs0ydpyMAmWH1mnqpqm14eOL
g7kLTfXg/JONhPmlsBpDRC8LFrsd45oYp39nrsStloc7ccgrwo2s4tXkAhTb0Xsz1/HyTLl9p9Rn
bV5UZAnuLz0pT3SIJ/Kcn8u4Gw1ZOQcHQ0TEWx95uFGKlGKUJqBfNEJMJqIki1vZnzpzi4moC4ik
tCDY66IdCaJEpV9NVUGoaGYKCP6quh9ixfRR86H0KtnWNOqz3E/ruHI5yDm73z06QPE0bAAd4r3k
dcLKVSNLLhpB3MPeFCVHCSLuOBOaDm2pY+ZrELcYDzva9FGdZjNCZSVlcNVWePsmvovnAKfwkAPn
0diExSdKyU/cxG+9PUDmYLcdnvME76gCUAhpdXeyuTXbsV9xXdsmMt1BrES/6U/x0U7vyj8HSbXU
oIonOQB/Av/nqnvXfDh3qs3uy67qeiexcnAVl7Z9secbkLvhrOASUQI9q6Roeu/ZFC5SCcDmZ0/L
xi2VUZ9BlMVFKXzpohbJbzeXI8BkHxUkBegf1AABRi1YdFRuUL1NFI8jz+piy7JgtW9MzeZoerlP
PwnG2TUsAmFOKWJY9csKHK2KmaK2yIGTQ8xNIzQipKSBilweIu49CbE0X8k9Cbnmt7TXfiSySkNT
1Gil1RaS+QSGSxqob2Zh2l7ULC3powYkMI/DNebncg0NX8h1O944QOclO+dLc8e4VuaXabcmBvS+
XkWs88jXrfY3h0qnLHZYgzPvV2Q9+jLhV2pYqWVrsYRJwa4Th4eXQ0C+725vw+6QKCR0AaGwAKbH
vLmgK5kTgYadbkCivwF18pb2KgVJ0BGPD/DqXu2C2A2RmJY6Ail6HkoWqNen6fI9yNEfhs8NHU91
z+Q88YeX3DquWYB0RF200yfSXMrunXHpDhBjVAvSoHfRORyXRh6y9O0inF4vcLgXYk/09Y316qLs
Apx9MuqkAIRAkbpdm7jAGuxFi4o9K2H1jRNyQaNlYrX5SBaKgW9LnKY1xQWLAZXDHrpwl7WBwip9
XYjwsiW8mA0LjYf6DCt37HgH14hxoaBfEQdILR2t5cgpDuLvdx3MaFmYjOIV/bcNwukqP1rsfVi0
moD4gTHKsWI/N+O2uQzVpbEpPCyYbHsBITsmtTkkQvRpyHMsde9tcRnKlLGnqzwcrOC8kdmqZQzV
k7/DBuLWi+OuCtsEP/SWIAZaZe793eob1NEL+Ljg/nLbopgQB3pap8s3c1UyV/AUVlLQ6bGy5okH
Y2ZEFOr1UZWlHb5fxHFofCf7XNXiu5VRBzb3HwRAQPGt9v1kLmmlWehNhOFc2aGTWlZh32maB51S
17QVLza+80O+/VaBuv7Ck3qqb1Dcsv1WZjVJexz7TvJwPsj0sQvuk/LmSRlvj7kDaHj2XEBhFWLO
B/+oNWFQ3sgTpGzP9s6iVrr1tOPyUYgLrpGK0xffRYcBXfpGT9lpJMeORKYqTTLNW4TDovQxPNKf
7YVzfqafli1ZatJiNRsBBXbyb3qjqYQgzAXhEVKHRXkLXhsEOetbUn9Ckf+kwt9q4u6Irt4dsHQN
lbEW1KH69yJIJu1dXdTF/3vAul0KqRh0E0bKgd967CNJxUQ871fmc00BjaioatdQNP55n4XcRDRx
nENnGO3Z3coo4Y18sTpJuq6lAEZ2WMkKsRkZmM+mi9fBlliZnWl62M3HVKCbSeQ3pf9En6Di+4fT
07Ym1fkmE6s/rz0nVAkLEBIRBMSMAAouEuWwU/9GYNKIdhYFysIsVdHz8p2bHi1swqFdyhJXswEJ
y8MTUDECF/42OSQef6u17RIajTxjN7Ou5LTOKH57/rg6vmnuNo3RbkqkzZ9xSoHcriCz/p9MjYwS
3CldI0PKGdmSo/s+U/sQ6Ug9/Axc6ayZnalmhM9xW+OkdC5AoG2rwA6ZKzzX4bP6VrntDuBRctg1
KXDop4Zb57bJfhJ1hhy+w/cJqpJW7Y+CXQsBstziWdLcRW2iFzQyDkOcPSJw6L3Gm++hgNDubZC7
pGYs4M5Cy1iemfyzDkPGCobxeoYrHgmmUKK/LEq951VjnMf8nWrI/S+BfdVt3Dsr5/W6jCL4eaz6
XOMOIJvy9rmUrLsupunfdxsX8YQ6zSIytsDz+6w4H6XyU6keHA0KndpxKKIxANePRFNxyi2UlDG+
HJB9JqosOCW2aZ9duOw1ZZ1TWExhNnkBgkFwwRcQmxAaIYAzy5A81LR2eETcGhOdQ1AzjRYuF3aO
sB/tonCBTKjhO13GUXxrtoHdSFiGWx4Hr+JczCISfDsl4xe+ElvfvoYVUPIvA6dd4ev2P9yLC9KQ
5WvK/6mPXRnjw2Nu4YFIqCEjVJh1WjMHGpJO+IPGa570GYLk5kBvIYG0wqi9sZ2Z/U4MXK6SPa9g
6fGcvLa47PZNS74q93rt1Lc6x5RVWd64g3BuQpOevCsi8JnXj0sSrA9HRtB8H8v13My97FxBQ58/
cxo6PfeRzlj/HissT8rHl0ljqzqaFbDM779ZP4IsFW5XidHe06RyT269HVuZDaVO1eMMNnQS/t9d
1Orjaoy6A1izSq8imkxMfzk0iIiJt08/zyYTk7imRQDzb5A4iYDWw6fG+kS5mS1bsX/PDnS0CVqY
2R2JMaCaF27o5A4u00nwtld1XPEQ4d9crT3KTSdp4WhbZVS4+H0FDCFHU9oWOV8ueYQBgwqFsAsV
CY32aWLVpDxbGLFocQwPjNo2GW5/b+SW1GEZYQaeE1UULYfw4h8b1poVOF6GDsmzDw+geUrsTvRk
STqOEOB8GY8FiRqQcJJrVVnNECjzUeLCJxKkIpzMxjLV3hlSbnVTd+dI9TcKhSBxYRnOZU19+O8U
lvvhvLJASpRBIDIAabUJddp2TdAaVq3fwdOFJqX9h1w1pOf31fGktdo2JwakckP8FAcqenDsXvBE
1WBTuPgpeXOT1oJzihjK5KQHd9+DOs+lMsmDt43gS67au9v+XNC1UmBFdWcVpWx7D1dSLkKwFRSe
TIdzlQv9sTjROQ81FJgTJwe3m3mcgnk4vRGACJEUk1BP6TRDTSsp8PazNz+4rgwcDrXlbFapqx3Q
5bHJkBvVIRQxI03VIYtGeiTgkp2MxOvTZ9Ql1Jm778mvx1O74I/JKeqAHCuaxLpHIfRQq+AM05Mk
GC6QcBKin4GZaqGFiHAGBWa7DDK2oGmY5V+Y2MAfJSKnRpXE4Ceb2cAUccmCZCl/w+4haIi+Kv7f
lXlsrgZrV7vteUk0mkkslV7fxDRrmVEyDvzbx9mK9dEg+iaq9Jj8cNgkgSoLv65f/xj0px2cmizf
Z4bR53vYLXqXORTN+aQZml9bQ8H8s4Q40r5saTokoiRsR5sbiODOf4r/P5InUoA6pC6IcDBQuScW
tSGwFK4Ws6BqH+rJXIJ8Hv+DpZdjOPkEqlDeEaHGjKnqzYqLi/RYO3qW+7ighMHfYPMl2h37HkHP
Taek1Tq2NFzIgwSZVSmU1FVo3neQmP4HRLIuQyRMa8EGXK1r+PhUIsyO74jNuVJf6zIcqwJPxfzY
enLnPgMz6zb7WhbjIFD2oVZvqaPeaQxJTbDFTsag59SG3T7NQybGqoGgnCy0CK9Tdmtz0vvHFI7z
NKBjMN7RcvpNlk3klIjlWnwEkHAPnW0G4h8eLnWKrie5m+lKLnoiBeE1OW8r6QElm8MHmqwSiwRC
8EQA8TPgE2dlmk1NHWEz8L6WkHvvwU+vSSkDsitd1Gw/TqucoP2kmghjTAXHUaPu0shn0ZXdtu2h
9nmEsD1GluMG04xGlJ9gYDuK5jGgF/EIFlv4TyJNnShQNvBJ3djr0ZVLbVpKtHC4xwMCbWZeKmrS
WFeDLHi+QHrX6kfMlEzZJYFl4j1+a70rUIYFJZFt1ePDi3s7OKcSg0DsGwuvVsZde7GQu2671eG1
VYNvhG/YgihpP1cfPMCrXPkep7hqQ7zk6Y2DidxmVzGA1ly8Hg310gs8Dyccmz2JEb+EtP0N0+M1
iL4lzrPbYkcbmc/L2muR1wFYVOlkDxPCX0/Ij7MYnXgEdNKaCCkBTUYD057QQHe5+Q21s4ICTPkm
fAAnNSl3qx15u4HBLNOSQ3HWBtmaRerzu2deaGnvxKK+JyeOmTZJCvADskh1QqeyfJnxPC/DcwD1
dz3mdnktDvrSKU37wjvw3WpXM6ou8f9TqWq51oYieHf+D4ZqiYM9qj7u4PhUKXts51ZzVxK9XBwN
6kXtY6131STDBjIQ4qicY/XE8ozI6Xa1s8D/kpeskYa4F4v2h4TeuHcw1uwMyGr0nC1q6FYydzu7
AW1szF0j8Kor/VsJJMX7J6oAumtZk07b5+I3ctbJmUDbrBHH5J/SCj0oIeLyyqlqcPar7ZlTYHCc
DEm/19gH+Nv3Twsn+Fz3T/N2oHXXJBJ8XB05fYW1srtj0pWAY7tbTcaVyxr1KxIkZaXMeCYElGVs
0Vnj8d15Ws5Fpnb1pTurKdBgFOpbtRmIyCqYyWy9VJu5jdyLt98iTHPBrt8hJuRhkjzOAYokL9tk
jnet4JKeDfcah8DlEiFVOAuR1szKEMfe7dxczby/eN4YMxuqUqlaoCEMYJPCgQm7wRzJP/mTWlRx
XfGbaXjQLNG362SGwfOpWhVTuRJzpehXBFcj+yw1v19a4C5158G8tdExOkLk/f1VjmfLU5zFslZH
5KCDrrPipwxp/EPy8PNxjoHDjNaQPfYzuDjfE35j0sbsUBP0fGGH2wNKsmFsR1P6koGrk0x851mN
K+ocORUP2idKsTItDXsJeCzGk2dVm/0vR852QcKXJRsLQ/2jH7T7QgcZAwhJvp0zyOK4DoYVnxcg
uxGo5isth1AIIvuUw5RQInCr81dmOPd3qdkGMMzaxYdfADAU89VB9vX3Vyn4rgpfcSHy47WS9sqX
Y7b6UmRRssqOmSE6L/CRCcl9RI9SqcfvGTKlOX6BiJouz+Zmf0gn38mz8eKG56hQR0WtfhyOx8yk
RhFN9gWnBxm3PPEX4ATn5b+dovxqFewblflpw7ola3jHDq7KCtmgfFu37Hme3KE1dJYLDgsz1Sar
CUMHVCE42YZBew4SEayZ8OpLyo2/VvzOCwSl0GwFvdnEN2MD5WfBlDqCacClXcaxbVIz9h9jw2yP
MqqvIBxlM2KAkFijbYmPZwvH1ahSRCV3j42qZs6Kj/64kI7L33mgE2HveWWan9f95fKmJ0lFWDKB
U3B93TJy9SXgIlYr6FacsyQ6g9lk0ZszFyuEalQpr4ReyWDNs1RepM+F1esFddDwv7EEV6QuxFeV
VTl2+ywohuayc7SjY8sLYOROGm57zTJfS2FzFvcPH9FS0jqY1wPV5XK6DeWFCgLzFJQJoHxLliD4
kBH2yjLKXIw9HIDiMy1NhlyKvrG/a7gShT3DV3sy94Z9T3I8uz3PIx7GPLa8y22STpqJ26a7mhft
YBMNj4Xvk5nQVHj0h3Acq5gUk0AGP2xr7xk9XFrF7V3xVbICv305oyn15GuLH+RX3MGuFUWJwwd9
SYvo28usU5Pi1wxv4IfguszlxNSWBuGcPCf764mmZJDo3fcQ0V63VlAkFNyRNDVOY25RMm98J9DV
UNhOi+B45ttWZLQ9CwvP6PeBB9Zkrg5NRZPg1MQZ6J4SMhPCTs9TX/J7hDbA3HQWO/Ky2uTD5/Fh
wrvEJDS4Q5atI7Ekyqo2dIkMf8TMFlBCM8dTZb1xS3aJeh0sq8C1TZNHK+1c3+f4QxpioQzOwb43
lyRN8agfpEsjO+k7CeYAd6hVln+mwKBo8x7eUSxQ8WQjV5uwp++ZK/jfWDLcfGESlhXF5SsoOpe5
qsvaC8D+X1CcoHuoZr8y0Il4QyHCKdCxiDqDB3imL/3l1yEIMdwyjExM7IPnPZTlwbF+BOneaAic
1Xz8h3kWGgLTRanH7h+GeFwKOfo8EFWVl6APDCsX77KJAb9dtg+bnWvnEER0Jo/EmnMWuVZIFBIe
M6cQIiBYmOiZuMe6hElatuAq4k/nutf6MChRFkQpp5IgmzADFaPvDriU3BGKfuLyHf4BkZgw/KmA
c1obhKN40ebk91ielBWd8BURzrjXNXPYFwqKtSc8wb5HXs86ff8oRSPSu8mu454m1bJbk/dRmU9d
PwIuURjEahQIGVRsGW5cVB93dOdAY6LrwCGt5Dcvt3RuQBHtxNJOWVEKm/yR6jiEwsMk0wkeQHv5
QQgOjbuoNMrEymmeiBuxOF4PCj3pkFsUopnB4LruHs5515r/DiD4uHTuMojl0cEiOsIIfJAktryB
jYEUVLXzAzw/18qfV8+0vyhU8H85G3YSR3euPdr4/8fxIy03+m2GjuYivWgeM8Zc7PPsOlEX/HQM
MrljnBkjp79Q4WgKEHQJ3dImKRGnA+mjT1JzCnsQUdi091kvQKTE0FyiuHD8En3n6BvTtg+r3zRu
bJ0JoJS9BbNixi2INNqw3XMc4nvBbbjyw6xRC4NEGRep0LltMlQ7sUYSAjFC9xotaynTPozWYJAQ
NIK8w00H1CZQjqoudZ0mXQJXdwnPDtR5MMlZTZI3+odnQmE+hTH0CTvD6xGJICQ7vBVliR1vrKYP
6hIfInpsrgLzC1H9tONu1KPSjq+HIpacqIoW77lRiUTwi3TLKReKdFb4UbRGVxuLpUGduhUWn95U
9S00VF0BRR9ZC37+IyX34M2+/QWtF+6tqV7nQplWc2851y+xH2J67Obsn61Un6M5yoTyGjuFKZ0q
EsM6Yk3D+/H9Ckx+U+FbcXxtd0VPK/QxBxI6ZtRCfY46Mv/LYpWmdBWJVwvO0nUBtdHvNI5lkmdE
YSquk41JjeMfXjFJw0KM60qfjADl94uAgNaBPmiFH0mUd0vMj2xp0MEjIcwp950adNOhCHs1P1uu
Nqpt+8o5VPown9D71lm5aVLbgimgNDPjEck+hG3Qkl6Eqmbl/ly8KParJPAlDBbNDF4sqagmspND
auuIcXFrCFnFW26SnRgV8MeGEohPzMX2ON/2EEAiqdcf81lnxmvnYodQS6wvx7EFxbJsUHKTF4gq
TO0yHi+DC/p7n0YVTU5czt5TTI0ovpnf03pkYCnv1XvzHC/5g78jif5JH8MvIyFj7PED1SvduSdu
dtG/IS/728bk4NjjfPCw/obI7KIECYvVzv0ITAbwuHKhsJwXQFCGm/H0nEIzdRAwPn2dhRBAKWQ4
CvMR5QfurcTuFVrSSxeAEPM25BwKqcydzmUzleP63kMDnb09WqaIMytyx41W4dV1ff9ASYMWBco0
7/2mbTWWZ3BOPQwKqZZpxNk13qHxAwTWdiBm/6p8vk+c5iZG3K755iT9LTt+HUgtD5NChaSVLeTk
F2UOu/VRUA5NWR4gcDpzQnrHMIKBuWfy+ilTY2gP05ufexFtuBZdt+5uas9nTF6+YmTWmIEIff7f
HWug2xsvWun5BeEuFVfU7LpLWPIcIB6QbwCfeF9kyUY58B7TUkVu+JjXpCqow7ZqBbsGRmgRPwQg
8SBc1INmntkY6K+ynwacTGKidearsZ3Eiswi1xLC6rVVUrDHGUXQHSH62F8hOmAw/HTQ17k2PNyu
qLUKhSLl7Z1G6XHOIKv7gwR4lE1H8vITk4h0Aj6ZzlHrVx9nXz6Y65u5rzSbmH4LqZrx68oYDzD3
vlGyP1mGLJxHWhxIVx79veEPrNhx74pJWX5XMKPSCCe7ySxuOaQS8t0r/w7TjGQMKnWZyQzUfC/7
4rIP2HJyMB6Z2T+xP4QpyIxJxOZgDvsPKbra1njNe3yb2Yf1H191EtpwIA+c+6wf5fPTwTT8D4n2
nyMZcs7Hw/oHUhahVsU9V1whbPwj9peb/a9uLl+LUDwIl8IUMDnh8mqjrYrbKC9GnUyE8ElCgF3y
LKE77CS7jLcIQ6sWm7WQHX/iBBS9x5r/hkygydbdLvc07Z0UtSrXpDbpmart+Pxst016zy0HXZea
cgj+X0ZIsTckTZ4fXzmd2gG22awU+vTNgqFgoYRwjj9N2zITIo5ADxnnq7PdUdJMx8E8STkiqszQ
YA64HdX2J4qjNV3THW1Hr39RC322oBT9RWcekkYGaJkUXUAqvbHp6cW6xKPZn0EiJdF6cIjehYuS
+KCGli85hK8MOuvbdJUdnvwXK04p5CTkHHI58y8dPJH0kg+Bp0h/IWY9oYCZh2G2n7a79MVAm4G2
DPaJari2Rv4Ul90eYkrhFBiaHrmCi2Pyj913ogDPdxm4AK/9tDWZR9fisQEeiGC49SHOj3v+hN8C
W7upBdWwNamGayTzBlzWL60zhrOjDu0To+pTesM2WFD+mkY8WGGCrnQX1zHXoJz3Ne0GYRJdwR4E
BeIWSApxX6rYq86TfTyCFJFCTq0pxlClGDWtqW7ZsjYemJQaFh7zrfOiyHskSRKYH539MifCtnT4
VO8iCMyRM8KUZWmGYfN4FyovQKH92woaIMkwLbVvKkKGnQTxS997veYfAKhu8ZDuXW8KVD4tSS0X
R9Cv41C2V+fMP+iOWbySRuQ5EwWUsWhtsrMNT+zIHg5WXKLTRoOMS1gZf69jdG/QtQYDEXHAyH7t
7wZd81VRJGJM7iXNB6iDow59jsUB23zeHzdPXQiEDzkigibemMuOIPnsE4uDu5zJcGHit/KzfkJ5
oktJk8zBFwB1MmVABQNCnT5dDCIho4Cvxkz9PwGBwvGFgBfFYlH7+vCXYCKvqO+44Qeu03BNhy8q
tRVQAAzqz3cb4EkuP6WqmaFHUtKmX4FkHMCmHpNE5g8hsRaU5ssnFuA4uMqeJuGh2XdetLHh16rP
SiGtylkqmUH8sMQ3gCSW7DF3EIRWO375TxmUqr2SzBkM4PkWKcmVw24dZTdVyfo8pZyvE3Nu95nJ
/cdUk/daIcVPx6MXnVMHVW6v02F0SQIgAOfjV4tBq22IPH06khB2hiNKFrz5mNb7h498PrD2unc+
WWfkqcE2QaGowUpJTGXtACPUB0GVEUPXt1bM0cqMTpHHKS9sE1t2QnwsmZdzGqpJbgqnXHNfOY2y
nsshpG3PwLJz7Iw4FJY3ClBtqBrLaL79aIP+BY6Y9qloPXgImcFIKHXRp8sAkazGWGOX2Fo/NT+q
85uMt4gkOS0JX733W8gAWIvjCvaWKNiXU7Omd7ZzpNFIeohJpvyfQwDx3TPqunfsNTfgK9IUnb68
FutaB5ol/wYKDyk/M2pEeKbMNFruIsPvOM8niybjmlA6e2u2xEFzxgnkaxCLdmJnl8A4QQa4iGrx
Un8SfPWAp6I/UJjN4Lo9dHXIVvPZg0qoqdxdR4Qi1DkjFLMPQ/PIt18+9cwcGoVAb3oViRQMy0aP
WG0FmBJ7lUCW/6EAz66YLJZKmujKSTw/QF16jU/idwD+Ypu1tmo5qP67j6RPkLHYWV97Djv+S5PJ
rYmb9IjqG/Jn6LcypzCXNW09d8GzaAeKy6JKvcmTTznIN+vs+eYC761xmMVjikACFWWkiHkD5BNm
lp/SKa+xhzcItOIhxrInxWzQ8uFmCY/M8ZGx5Br0LlbXY7MiJiiPKS8+xhTL++WvEjeZNix5FNFH
1cUPJ29dYphTN9O/YWrLsKU0rUfpOtpHca8NFxoi6aLH5g7TBXlW5N7tyI+Xp3uUXtPuT2zyOMqr
vu8yap+BKqdghUu38BkBOwEoYQTzVqEtoYyj6pBXcJLZpNIn7HpCYE9zZcgCWTYNR+yqsEsbjE8j
64ng8kN9XbvMzinW4f0Bclh+yuOtKq24crsJ53M00KQbWOzjJmBDyGirJdAqUXBrBWoR/P+qzVXI
mNMI9ygk4l2zz+gh6f8XutvgxSvHqKFnpPMoIvTH6J+iNYeWoqnFzOz6ZVc6Qz+Xz2qNuB3Ld6fY
g+KESfBaHeU6JZDsr01NeuChDzRXmP3MQGCpUQHqQ782IerpvdqOlm552m0FJ1mXAXXTIL1UPRjX
8kdI5VtU/KTc+Cbhr5jxaT8Zuzut3guDLC6OGBZPxi13BqGaAEwTp/ndc4RjXPmboZ/jmPgve5rW
a9PDAC5VFhOT9jXoW+f16Je+wzrxL5CAAviAcrQyryPPp/w5ZPi72oIjw0WfejDNu1g3gRoczT1I
Hfl2YylBsAbMG1lgC+ZBxjhCNxE7v5qBMZasQhbjW7lT26bbVvor/0VVrK4UjXkn4+c7eSPd1Utd
GXCpo57/gDb8CaEeCYdFSaqxpWMCI3KNja6hvj/jyO0pfCpJI2emMtIAhBjAjvxK0p1Z15mORPGz
bU13oXsh94Nj6SMFm1E4EDvMxL7MUc3NASTcvm665AiEokrMUyRtJiv8BmzEiYbzYtWzCFBT2Y1z
6cDB/Db0EIPi9Nv0ol6pFgrIb5z0Apcih3Dp+5r8ye1iaAvXYmIZ6GdStuBi8JOtZNLELdI5POgu
osT4sr0jOC27NLYwi7/hj7LMBEX8MCvHae1vwJvvfbgPCEavAbAmb1Or/AoCGerR6aG8Lgg/GFqY
rE99pld+ZMatiQk3F3nYqlnm17xuIMzsE7ulkCPuOKv92KKGN7ezJRwif9NqMqHYlDR+pN+15B4R
pi0ut8M9c59B1dHFxBEUAPfVJokNHK2XM88GTLCezc5IESWzwoNedHgkwT2KRoZqQdXUjvpfxQnm
UxO3LftpoINfWH1KBV/5jOvH45M7YF9W7Wkr567LPzsfWffRZmhVFArxnXpS8Vc1eEK3weH1Wv9z
GlMXAr/FRLH6ZzNiHHtoc4cO3UGiaSEgh6j3rk6ghJUjNcpg82z+N8axVGnTkSuW3RdKlKYK/w3X
PU/8+SCj3gZ53OKM/9Z2/LeCQfueAKzrzo9gdic2Il6OQUDYdViNZnX/bpJC4zxy37IFQIcxxGkn
4i/Wld0PC+fFeWc6JK0IfAYMllqHszL9xJY93+NMURlLu3nm/3qX3lHSo7NUIb7ZoBRIV1SxIqIz
rqSSMyClJbxsZSrZTQXrng7+UDOQV71yb4HimGzr6F314tRCuiZgbQZIz50yAjxq70ILksMa8xCV
L9B/drlS5v0QuUQOe2amT9vVoe2A+GdfQMlEEvzezWY1kRkQ+8vDCs6sM9KhHRBl03YW2TsFan4z
byqbvM4f8i6PD8BedQ151XveGLb4/De5KqM7mRfd0bkTfTo4xBl790RalPOnYG+GXWsxJWyGPSrJ
BZQ9X8hpsIiE2R0ZhjWj0drsOBGjzjy+elknWtXs1KVfUSy6p4NcXznK5C+V/HGYpzwivg0SXVY8
w2BgUkoMAS79CpvJPMoyOSsgG4Wu1XPiEjoSgscKIe+t79i8vYLcuKThK/pwG3IVwCIl2gqENC9D
5LrdfUIUPfipSPeVnrel1VGcIy8P7m/Pw+P7zA+Gw4rerSubu4Mec7Pv58/W9hKmacPtoF5o5jri
JGfidCoBbzYhLNmvzwUGELbcoT3K6tkF5wc6ACXHyJ5vRP+lXUUDye5F2JjHrN0pNmimLehuQ3B+
tzQ4BeYvFlgc5/N7Z9CH2YI6O/YjZLl97beyET6EgHm608HUlhbjYlh3oYqyxzaI5G00y6CSYA8o
wPFNIzsNtahkBciYewaAZbmVU0IeroUbg8wAA/OTHFn8dq1CWVY7xwvmEfvC9X/k39ZRlNpol+Un
TC6QxeM+CQq3YT1S6lsO/WQgEZ0B7HcoeUMtujOuwmQMjEDU6ZpbVQLRQgJJlFUrg7Be7Ql637n7
0lqyAeGw1nMjV8ibBIEH2U41Q/PAEMBR7gkq2e5evBjhqsLozAV6HCQdHUXSBcwUxyNgLYSZT+lb
f5HqGwm88RwTDZzhvcn4KUYHuB/2CmCpkQLMTvrQWHJIx/mozfJ9pHVNP0CJf8BwkBMi2YsScr5j
LzhHtssrdp6bYje6kL6u4HUXwJsXk2m29ez+VlN0MUTAMn+LBzJinPSA9/V6qdeAMf4H5ZEXzOws
9P/QAmA0rJ0HKj+zp7GVlpFBSmuXSVhQ/rQUgsR7PX4H/X5MuD/sFaXnvhD6NOCB+UEIUfSYmbG2
KMyrYV7XjH4qrS9rrEEZSEUXdnlQ8rF32CuQtWDpVsYHDN3QaE83wsuS+sah1kkh3i7diyH66zhY
6FqxyhzVF9cZ5J4KCQKO0G9BH/D64ac9OVZjUMsRau4i91CH/hAUgnVWVEvLwdYWE9vJA0Drd7M2
QmI55Bhy+H2p04lIJEQvrfvZo1K/f0mWHQhHjQGhd2MNUOZLYMtXvcaIEup0uNejwdJzM6SD9m2l
UuCALMyLFV3S9iS5PoXqRyDzGTEx8phRJLkgyOKlL/48NwESh2s4KUQh3ZUBa6kY5zAPLIrceyro
/T41FYbXCXEBydkdelohp4fzH5Y6CzxO4gOieLXo3ZyUvWC4NSeclW+ye14L9k66Ifq3G/TbpvZj
a6IveUhnLFGjRu8dp3sEgTfwdzbs5CGMBA7RDMWiOPsdVpEoFSv12AtwaYei9bzAAZ3M5fYK/M8e
wKj1Hu11ifM/khnh+v9Q3qXK6N5/CdpC3RDMaG26VqMnHOnQuinI+cfvVkurH/CJZk+UhJJcpmOi
XyOb/wMRIgAGwRqB7HmIQTWu5UilvTN8Ij6SDvEUiSE3NpjOZmlE0sP+3TNYcjAfH5fiE/mv7qKy
d1YA2YoJCj2Jx9J9fux7SvSI6V5bWg6saJnoPOl+mSiiAruH2bSUjw9mbjFp1Ast+unSgDA3UweW
lD766FvX9m2z4r2VTSL47cDvcR/zKpulC0z8V4rRlq8uhigRK5r0EFzDYHx+VOmP+i5Y3ROssayK
5/eEeD0jVDRs3jL6BaYCPFI7vn4ogy2oRYw9tvJBbjMeaNYLroWXDewfCfopxq2hXmTLzL/p/KYQ
lFMmcbQYR/pmDrcfcpFOIMX2gGFTSJ11tL/S37Xrxb4aVdSHi0BRllW9DI+QvBjPIYOShqDkLj3X
bIqSCZNmyIWG8mE1x/ho6yeFFDB2CDG66oS7zppNMpXVRv5ef381qOyutJA8fdztFeQV13hi6NSI
LUPXZoXad+bLpfkCV4zZhQXXDTbWeV/BLo82btsQ0Pu952EjoMYhzS6OSTERM7V3tpxP+A1DN+TR
3ulS5oFy7f1nhegxLTr+57F04LX3ELHOFSPhzopmhDOiB+clq5wCqZhl7234/h7B60zebptf3mtu
M/wgQ9cedMCQ5QYJHXGbiLyu7Hw4Q+IWT4uRZh27YTT2chGxWoGx6mInhVPuR62I8jic/MFOm1+q
KbxPaOoxHUiZ6p+9+x4Tqm+GfQSQhM36Z9Gl8w5eaxn6KCZunB9zU1F7kIMD1thL3HYZbo95aD6d
QFcNpRP2SAHqolg/rVGyO/Q0/suWqlAFxcyI0aHFEnhpNuRufytV9TyBd1THuK4BHdTWb4UJQx5y
1U4sU1KLdGfyIjn2jmtGERVteJoChGm+b2VOTdlVX5W4z6nfVUWefNpH0AKRYBd5h/sq4pHxNR0B
N1f8fMlU1JnpOow4qidUSn41VcAeaeRs0Xxg+JliWcFR5z0jdtTQEHR+x7YOIf3HottoP7/SdVLD
KHEr2VpfNbcSXaL3xK2lxG0APP/d4NZMw+OH9Egk0lRJqHIL9fSKB5VStPbXWA+gGFyOkBPAVZWX
xrMp2uw1DfkuELtGhTZtvUOJoL3XUbzWkBQm/H2hY8KApR7O4HXy3SU8HB8pW+pG0rcWWUUhsP7T
e1HRhL3FQ+Zk7ALnimGBRAiguGaklNztO0DKw+MjXw19WBkH/zTrTRR+WRyXcaVlRrdG5Ujrw1qH
wSXM/gklXU01HT7IoigeXx5K1DScdNgu2s/XD/vJoVdlAW5DnJ+KPAQKYQcYOVvau3cO+0VQrG8b
jtWXXPYSl+2gQS5zdqOGsvYht0tHk2tfAYXd8vOX2ObMQ0IXcmEj4gYr533CebgqJ4qvz2Khgw3i
DWdBeH4u9be5S+Jm/3ocOwHjigppR1lpxTMpRRngCJQoMWj19ZRlMkgIGxwYB888J+fvABdOnjMb
6ZnqahmOo0P23fwYoJZvh4bY8iuZpdoRlZTIa9oxdHTJyZx2qbpOG91uoO+ktUziMAkpIMaNLFVC
sSgfEuCpQC4nk52XrN2tfj6hFIpkIGzdNYk2sZi2kZjzxsGzOKeFDz5jDqeWK934ltr84GJ6LlI2
f+Edqs/du2L/oHI3MGarrTQp2kl04oNviXadYWr1NWkQYSu3CSgwHs0C+Y55uo85u5370STK6R1j
VlsA0JkZkD/ku4Za5Nqw6y0NZ2hbOSwiPorDSpqQfQHJySTCOCBc84aUjhjtQzzFh2g9uylR75Ph
SY/6qtH9mg/4IPVC7B0DbXqpECArmNna3wQXMTwa64mde4g1vvMAnlglx7D9mL9o1CvIq/c7pDJM
jmUavBriHyMeZqNZudQTyMD17VLAYZ+UDaidC53MccnTKNX48eof6torOH7gOEfPyuwyhMkfapNh
ENUG4099bCAgBWSaR5VumWCnkl8zG5O83A9x/8PBnLDxmf+xsKu+CmrH1q/vtDjtyVIthLyxK+jZ
ZagnWO9LrHyqxtUB52UZFchi62eMUK1CCWbpJqUTHfA4ugDo+75+oP18CxEfAaCSOhyVhAlG3XcD
jnYrFnhSCk+tzIug4LZFLYtwWVXDNV5a3NAWMlsKzqTbOXgq9eTA3lHikERQFmBoZuQyjs5z7okF
0PA24R9YWLjs9N8GxQjDc/u8+xQKZ/NGt5QVvMhdWCQKgQ1DVCInetwBxq2CR/Bs/yc+Vimda7V6
GozP1FysN5EOao2kmhlDLXwy5JRgcsSiW5ux7Q4BLCMplNm8u6VCL59PCQa6c66kMeeZCflcn2jL
arkyR2hIRTbYv3IDPYZSBLXNAn/PoiJ+25Lr6ElqB6f0IpUdJKDAa62t4vtZEvfNohyQ3B1IovQY
vhGSQ76WDhh54bZeR7YOuQeEKuhE43xFnSZLNmXASOdB6TlIhxyZJO4U4U9lelCV8pKmGXFHwU2F
K/ISFTvLhwE+roatFpmdiUCDM2rTOhAAoERB0QRFzHrH5mvJGb+zWGCy2d8qhnvg2Lkcs6Gz0J9L
6oO2SPN+2EyovlztyNo9kQ/ULVGBgfRbl/TH32tTwBOJZw0RCMzxFy2bT+Cj2b910pjw7c0TGq3l
swd9i5TV52RZ8y4iG8ETl9HEG2XKJN3Cv60j62PXjyTrd6YrnYqE8r8eLhqkcZy3051u9omPNMG5
s2TQeNoMgf4l0ldmY4sYMo0jlezcLW4TcSQrc9/hNPNBovkx2CawtY9D9BqajzBeWspUhbnvkk3D
lFq+MfGdaj7O7W3UFXsFxol/VJbZV/EaPvmU5M2AwoWz1oC9dW95veOUj7Q9TW7vewaZYrKh1z/g
ceFJAay3ALx5NwxTPfOYHmZ9nhqBoU8V1/nl0fwTTKycNG4X3DaCiy2ytaa1/e5fzAQwkbb8JTa7
gT05Lgq3qBTDvEg/t0BCIFTi0qNXKi/XOEhmRuWlTbKLSjHDNA4pikZaoqKXfNgw24Rv3o+LowOx
JmcGiEv2kj0nd6yGuDEBY04fHH7MxaylQJuvcjbKQZLE5GTM8j3AzBTrww68Xzb9FlRRJnzozHqI
DiIr7KuaUlOw62+fwLjBxB0TDPN1/c/QdKOm+jRaoP59QMCNmLO2YYAwIUq1Zf4Aknp1wrHaVpnn
8RJWsduz5ovfXqaBTq4OQb3kRGCdDLPWya32DxdfaXpPVMdpoc6Eh6vSxAsBu7mbb3DuHZJGTrO7
tawH63KXfKyfa7PjIoIHnCApWrKDn7J3ekRVpED0x2MnP89nFr4Z51jIaMx5bD4pv0xUmywnmztC
jgB/ZV+qMQrUM4qB53XtKST66QNS29cFTzSsvoP4WVZ2cWScf1l1TItDV//wPUeYs0j3+HTIsskS
rtSnK0pajS30dirsGNKk1P77149E1QAY86X/lWmqCK+SJ2VnhdYO9KqCI4piowdpL1NugZ/XKgl3
16jVs7Zs3wbR5C7iQXtZ2Doae/Knx8yb8SQ1HyDotJY0lrWVuiITOwa8GjcMoHzlBOHOJga5DEcH
FqGz53K15s5gleRUVXdTdkrj/qjHRJWnxjmQLz1LQy2998da6WJlwCsdlVKiyurUBPTtZnmsaNhQ
aSTZSW43dqSy7b/9xJbfUeUZz8ubgcHMGzUshzlPL2hT4GinT9BcHwtL4BZRTnkPYXMEq8qkRi1o
sCuPcigM92alC2lX70XvR/jAmEcUaD/69KVoF5mcjqLnRpjWAHZPHTY6SRO7yYigtJWh2G7Hc+Lz
uwe2VJBKgFlBtBdVSwAYQ7ckG5l3UXF8Fh8y13bNtu+ukho2bYgwoAsq6XEsSUt3VWSUKefrCjkJ
Z+77qM7Z5nKuz3qo9LnFl6xhpZEYA7pXLP/NQAr15w3qVF8e4PMgIADNpnk3IgWshYII4FPjqh6O
6tXS07UORHidqrN4/3zhpA5qQMV4pUasySJvifrtjeUcdfZ7cSWY/UnXLntpIeSVGgYnm2zdGLfE
8SUthnCiWQ+NoqbBHCZOdd69IlyTaVHy+AbwCn0T69dR4NBrQXlNcznnV0FdqgPFi/KdfUo/rjar
VZfuspnCplWtInsE8UgEc0uhaqTU9JYs2M2mUIHrYUGjWX1Ytk0sPlvHoYBk4rj/V4LP4Wq6ywQr
z+IMEmG4fUxjyxVVK5voyjOKmXruu+Aosz4ZF2L7LIPWNTuaqsmCncjAFAjQP1RsqRfgBj7bgbUZ
sBt7wFX7R1RIRLDz8kSrczB4eA9dQGELRgfAFtrGx9xX8ZNM/OczY6uaxJu/rSqGMKMGlfCuf85T
UnwvCj9Pd/x1RdMtPvtllJd/VVNeQVWs05DWaAYV+aZxE8Zl4T2PvlTb4ps7rx6EDWZnZ8WiDn8T
W54hNna/YdxkwOxeXkG1b4+3lPs+lkxZDHej+l7Y7g5jepnz/G0iSaGc+ApIVY6X38KmUvfKcpMR
DFpVAXr5OQmWz/F7XB0csO5YPEpE9hxprEH033SkWpf0/keVO8zi0QyAwnhDtje3sLiSGfqqhC96
C9J1XyJwiYZZPnk9WC1+snrtpidcebt52PMNlM9U6xl8laGTYL5zFLShmI7iLGbl4BCJhAF8OICv
y64vyt1juQ3xsiBguRui32gklgtQGnn2dZMjUbfiZNNH89gSOgezPWo1nut5Vc7hlPrONC0LtPm1
kkiDutdIEvju5iqzegGeWXewfBOvscmUViQoTI5BqsE8jGceznREUBIEqgtRm5vROztPE2wz2kuL
Z0AUPGuyYLKu1v2VM2+5xhUi8T25ImAA0d4QB/5EYzVgZMY9Cv/+cB1dMkUxloeIf0Z2iC6WKAgs
5Jrve0Gj8V2VZJT+/EkEGxZ70PXjJL11p3bPWtKvCY/omg2992fAxA5abBZvkBgUI/3OjS4wqf9Q
DzfTRDSUldXJRuCHA9qkY0s8OMT0SKgagocL4QZv+z6jhhEJwwGnuEdTGl+F8nQ/Y891wvl/Qrqd
RN9hqtsz/MhvGYgPRakg3WOUNttgQfEQazjNxN8zqFBHgXbAIvoBQCuor53VBVDKpCIthf5BMOi8
8jL9UF0Vu1lGmHuaF3Sc6EK669CyFVOAhlm5sGfXtSY8FhZGuUsB4ju9rr5vK011qpyjqrc6qIIs
igxNnS/futLsXIt1OBxXjVlQf6qNt4LZdCPeArnY572wZCCBVX0X9nUyoDY/fCrvsQOFoilB4f5x
lH9z1TluNTBE5VPpIQJEwGZoOWUrRhSmYv0CjIhsKTR7LhEiGMYffSdWJURyhpHGLSW8i6ZzME5q
YjNBYdHYmQagRGpspN9s0unVa+G6DTaE3LFtimR/8l7PnhP/P/7nGvUsXhAMfXGHgvggIWu0yHrx
7BJnwi4xFyCO6F2dZz4xBxvJGC1JYZhT1QAAZCx6IBYboIS/safKCZY8Lje0ckEgv/sja80V51E9
Y1y79PuqHrTq6nkACGCudsc5ofm6A6Ij6m+RJ99iJlJRh6PZgJuGx1B1mF3Nh2jIgJWabrdZF4Uq
ZZ5/Q3hiDTtIqG9KAI6SME2wkg2iMm3ckQaZrjKCbsAoCbnTEwDFm0Eg1pDfoSogOpgk/uhT0xG2
+pxaaOF1TXboD+0oqwU1S6QEG/8AGpx5mlRv4XhnY9El8EW04sxxKwfnHp6V5RB0G02nmdTVMB64
Wf8XYOQSpal/JT1KXZfjgapHA4Cbs7Xgy+gEX7QR5vc2yTZm5Sye8yNLicqps+e/nGurxFXNwwjL
MqFSsmUe2J6TzeP0Sffx1wRL3IBbpyu+iTG6wq5wqdogAnA6SnF8h8mWiZJpmaqCq2IBkE3BF/Ry
p4h/HehCOM+Z7Ab1sB5t+hzRl+PsnNniJMmzruAbwDnSjucfhZErqJFJbtjToTvnT8Sz4Vqcjjgg
enQe4Q8Oqw4vk220zuCXDV8b8zn7e5XoC+vfNXRx02wvdxW8WYdKC7pQ7oCuX01nkdXW0xm8lfi0
HlQEKWNpQgsz4EXFcKrypnom1I6E2/+FdS33AbM48OrFd2Ta61111GbAvghuCsPFc2YxMZLCH29P
i/To++W+2v5y+/glGqq1aIstb3DfefyfZA9eHKp/4+i5rmABWHUbMwgx5ior1gxA25rE6FrC6iqQ
kZjGMKTHgwHdcKqnOZXxQuYzT6hq1jdYKiPmvqmtsFy2UmyNda7jbZ6jPUF01WwOv3VXtvjjr4lw
thX9iBfL/VoqXodiUpBBhoFwD4l5s7wTAo4hpvVLDYx2tWY2wudpneYxeEcmxnbTVwWYxBELA9e7
L0ENhpdiIzeW8fowvIUXiCA1SRZB0PzodSRa8YWri0mCglf0Q8v/zzDeB2jTYnuiNSbiuWgd0j5j
V4s0sQ5dagzO+bZCYsVA7Ovx+/AuphMUHjas/UlBZVFIgOFd2k/NbD5ArPTlJqnHJQgfQ3XhH/5/
guK1Z3ctZ5jvxpZQbN/A/X0K0u0ZTswZGWp0HuH/ldqbyyy0Z6J7aKB1TfVb9+DXfw8uRlGuEcEE
CGLpz/m5G4CLputQ4+tb0l3gGnM+ncZRlbR4YRXberNMBUYW7YoyMK51437PGFadQqrZTrZpFmAm
HfNlkJfZW9AGgIj+EG5zb9018dAYIc1JGUs2iMOEr1b79C82Sj8iIiz1HAQAEtI2GfD6tt3lI6mC
+LgLBDk2jMMMM4GLdMJmdrUqvmg4pfV7kqcZPC0+f7jAOTFwugbeb8/SALhndbxMkqGz/bEQtckz
CwMzRjK+mea1KvcQFNcHiEWhhulWJyw2vp1Hgm3hbT1x2SGg7ZYjJTsPrjp1YFqeon+hiuR2/K1L
eo8gjuu1edGE1e59EL9V9OYNcwrRqcay1G3KvbR3b09OpO7EU60OTz9uZKAIRXBDVbfNn8JQghRg
SSwKAHNiAkHUdRkUyeczfuLwUDNg+2zKxp8aVT0XCfFpXHyqS7EyRrmyS9O4VOxd8sFhvWj76ztP
tJPsdvTJ4IXZ5NZtLYqI/CKrHG2GgmniTuJFO/9dM9A1VshE9w2+rZ+ijGD5TINIK4rGa+XH83L+
1QfqgSz7sJZvIiKH/u7yhBWFRAOxLIpTKcKMA+UGbrPZ+x9/l7i/8dMY8K2ojoAyripXY7TAfiv1
yYxo/zm5/haCn4xH+odcOzDhAOPkjXWSGqWcP43tbauvPZ1viFA/0WBOUf+xMUaUHN+Tf855FEB6
ZyyPLtfs1397qIv78aBoI7TTYoVgypg4Mm3Br4rE8O8iDmsFw99vR3ttUFKcMzGip4+al/gzFODX
C266erP7nN+AEGKZli4l9wE7/5fDMJ6GruFUQA1I+xwJDb+Iu48/8oc9zbW4kU/STWgiXpM4eMLG
unlFfQQPBBPnzMhjxra0mY0UurVN+d2Bw6VGzvMU24D332Di6bBTElSBkHe/QPsl0snXQPCaxK0s
Fn84AtGSVCCCUJJwDHt/yg1+rN5+U32QFWsYOndEJlxQnChNokp+a+ZQvYK0i4yzi7tjc5tNneQB
iov4rEtCbIPrYUquCZeA/k1W79VX5dIvm4qiqRcnoG0f/fFx0t5WFYn5yXV23rjWVS6YNdz9a1Dv
nJqiifcd5t2YdgzdRLMLNLjtScCjXULcrCprEygdbFEKiINnyRE2RWfR5NagELMGu4+8zugqp48G
nXzvtSxiFCz00aX3Fs5Wr+RuOKahulOHGAXWW0SBc36LEwku7u+PtDHLPvu/8CkaOod5bCqrwE9F
t1Csgw36WG2TrupPetjmIIifGYDoZDyVOpOzQSnwHLQwZ3UNkzJnLSKTt55jaxEVvqu08B8QaOSF
KCsPVYZfft1OiA66U0slrfvXs3IfKaG4X9gx/0ZlvDiViqk/7Ni9z0USsUucAz2KUDhhS6ffGTty
9ZWyDrx4pvT24mAbfqkg3DhZKzLdEGVmeHGoCjV67FHDl7TlqFV0twO/YfjWuqtboZ1hfC0gPz5p
zY2Oz0RxVIiL2Zr4EEBf82NbnrDgqpA879vxLW3byBDubCQDRU/rU68El4M1/fwX0X+A0n9EJd9K
vh0OngKjdC3JLrjBbtM6twerblEEGT3JaVq3N+k1Bg74tGxAOu/3FwcxIh+02hNAZVOiCH5/HDhp
Z7NqJAyKNodytZV5xYJgV4zLiDMhfxtIIlB5hldgXv04K7MZzproFdjZlXvRT7b03MS32Wv+xKrP
z0w/zI8ccIGjgln6c3R39KpHlaZi/KM7i5qGxWsS/4HJL51/Xoi0oGBluPat2J6RyrsVvQHxodZs
vmVbLdA17o8XX6ESYQEXxEASTYx6Qv296injCU19pOE1XykJgmaEpFi6SWxL0np8CP9XRIokBjQ/
j2bSCpHFLrGAJHiEqeJ/G3Nb/CkwiK1La7GFp0l+Sz83cUPGEczF36TX/VDCB+yXfzlBtTlt5cvu
8OF7n4M2g/U3p1OIYGF4fSCWjtisFw5naE04Vlz//LUk6ap3czZSDJu1Q5KhxRspbTxlP9yUB5gF
Ud0etgagT2ZEbPuHC4AcEraHjfVKIUQD71MGGR0RVGDYVczJ6VKvpAmzazaq8uUZxFMIaPeIjf1u
kUQGTbB9LX9KxehMjHBC28WLLb0sc60RQ95Ss+wNR7NJY0TFhRz6lUzl04Vd4ANn+L4ny/6SbVUU
6DdM3hA+58zFU2FqiSGlHHCyHFrVBqVBpORHXA4/Q06xk8DJOLGE081c3bToyfHIXx0hxmD/K939
RsF/Ku+P2KvNd2DXxfrolCsMBzFHcTp1oERmLZr4aR+x4YhwJCOUm6rAn3jOKXXG2M935T0W4aF1
/cmzmnaFZziMd3xG0ezTWzQYwK75bTlHtjC2rMgkEsk3R7TJCy0fGGRFkk3x6rmCnHgnh9HnefGM
+XF8T9Fcy+GcYZnDTiivR5CEQCW83Gdwkaovsu5sXgLIwJ8t9qodvRN/f1NkQDJMIJv5i24F6z/a
0TQPUJHFAa1Zapa9KW5VzgIhHrfFMmQM8TImi0dt5W64pYr9OdtXm10VK2jpU28PqV+3H7vEqaMR
+E5BfH/dlM3uaIoYSMwPSG5ClmA/8mym1EGrh2aOB3jBz/bH87TvIeJ8+lR0f/dRtHFcScah+iPZ
CXQL6hgJOEKeESWyZDaskd3bvlQLrVCWTNdMTpegA2HxwOl8IRS0X9vFClsDsHazOBHQnOB0cn+a
tKbPk/3J5pzhxebnkpK2bnuq6yY6ON7WvOCkSkZCDeCUaXqoGMT3jFVnwgNMqiIE71flR4R1A6ac
Vqg+yYkuvC+0Ei5qSul+9kbbn2QC+wolpvB5AyFciPFU4R9QNzJfMll8vwJgWHcRE3s6pWfEhQMO
4Y1GqxwMBu2wwitkNcnUsBtkkFLTQG7MWw4+VU4BHhn0yK0KqlpKXR+DJVQqYmgxkCSCPM9MbTKV
MITCvoM/EmtQ1UkrWavp1SxL/qnz2GFtlq43pe75LVj/115xFv7wu/Yv9PjeoL6P4zPswUtO8du4
vfMBF3GreDW4lzWQpaGfWVrLlh35GpOXJlaoKpkSDIa0uIhXVScH7mVQzVbplzglKUCWwt4dWybl
g8PgaIbTGI6flJ0Bl4YsnfArC7q/d5zOncC0uX38r2Rh7RZ9xIbOOQH/betBEBQq9KeeOyw8xaHL
/OvSe+cFGAJf4UEYcO/Wn/Mv+7BrB3GAWi9RhfKeOogeCgnDfFYCJG1WWjJHQ2LoeYUcEVEFIbt5
z2D5BfluYAGUWE1rE/A+3/JPmDHfKZbVv4uAI9Lw3VJPCqg6I4WhrIXuqYQ6h5HEQR6PHDmKVSOW
c4ENHxDZ7xFoBy3BJSAP4wMjJZcM/l9IL8bODjYXFY6269a8Od6iYbAxZ3tsKq9ocN846mkLQWtn
2KpbZ1/9IAfSVEIAOTZGQFkkznyHoHYIu/Wf1d+3v01Klyq0dY6SM4bD+YeWerHJQ2oHAoKTGgN/
nyLdpSBl09MhKaRxoqrkO86s5qxE5KXxWgmeQiXdGXU3Vy63LrM+TorOiwwq5w7aMwwcJibnwVAB
cz+9N4z0VeZx2bLNW26z01xtakZm0IDJzbwx9fZjiAagie5OwCUvoFCtV+PU3kZ3JJwknGjvAscC
15xcfdpvwQaSC8bxWWVoqi0TDnJDFPta6QKtnTggxpkZnCx2yaxN7ULjHJGZfrQ7Ln/Wlp2k6bWr
a4i1Vr5t8DE8C9GN5K2uAf2cIo2EfdofTiMPl/sZqwRb5G2yXXoH7CHjq8KVMrMUGAFsI6X54dPH
NKJpKQlsyAXk6kUTPZ4P4BtG1Wr/Q1YVYON8RQYXkR+J7lg9EHpWHl6Ir1Rw7Mo0R2SS4ZrbjqcP
+3AFQRUqrNfseO3k5Db1gi8lbTHriw/iD/t3HN/AOFUq1wKMmnrFcM0qmRxoSSTbnqE7xg42rtaS
zN4nPXqoExW0VNSEmd3sDlhCWPpQR/Ejry62aF9Tlsdk3eyFFIVUlKYQA76iZfA05a++vL7Cmyiw
A1grevOBStD53hdafpBu+YpQ4mqzoYOnqF7RCGAsBoUBfJS5SqdlVgHayAGCPjA7mmvOVed990uX
oA04LU4rwlR6Ug9l9KBahrypL/hmMzI23X3UQ+iAn4N2chaDOm7MnOTPO4eC29uOWe/yRI2rhJuN
cq7TV/ikQkWtmziEQLSdphNFqUgtPjpnUBmSLE3pT2Mmg7p8m7vMSGfSonqwZwv5lfS8EoXt6pgf
rrWIVQj1AWRtvCDPyDW2aCpdoIrRLa+/lj/QQus3nRGrkXhHqiGBZDPvY7TApO30gsw+r8BRK1iO
YKwU0UU8bdG8rut5KgawKdMvWy6QOrVYa0xlRUEu+mKXKm8Q3BlAXqDGk6FioLAzU+yGX/gKStwF
dIemYEUTT7sciZPDvJaJ8YLFHtmgxTEbr4pW+twmRfvwOj/FUkjiklBAPjUoioMa9KvftNy0nK5R
61rhQcSqQ7AAzsUoDkO6nxx8LTzQPqmj3GGWmu4fJhqKLdIvPAgu51Zq/uCjpvsH345/A9yLp9So
OKVHWAQuAy+hn9QD/6x/09UmDr2+r16dpVsPAA7RilmPi1ljOcStxK9a3lE8gXC8IQdmgZnt/8o5
rM8KwxFsrj8k2Si1CZRZ4W9NiYfaDfuFmAfDMf6wf82dZ6K1XUT/t9eQBgVrWY4w70bbcAz5JRFi
Ly6HyjR8++8eLd+EeNgclsrEhXeLz5FdKVKUV2/jezcFvwNfCqt6YKNN2aShP8fbxOCRBaVvQ1cD
9RFf61q/EBiVR27lA3Prfu+BZzTquGypg0rbpShKEB+J2m//RPG0caKrLPH2YxBgYZFcB9zkKgSl
p22CUKA2/+h0gmJhaFMQlEjqdUTrxqIV28KZMssBETh/c5zoqr42Kn2Ec74ssvo3dn6P1kVZSxxG
7m4VjZPKoQGqTMq/Co7CBaX5613Od8RWUXlOzjjdoa/Ze0+JheyOc+aH4lqGMJA0L2kQFcLmIHyJ
O/eyuNhbyy5tQmuM6bOERb6rHWF+WRfdJCSrrkywNuS6CGYdPBpLhAiNyhbxMptBYk5kE4bgiGjP
4DAP6y8Jmxy+Vlkv3zAq3Ata8tywER9E8rA/55OM4xEV/18K4oFDMmQ6GPCi4Fe4K6ogJbC//TTq
kCOHKiuLB029McHwjJfFRR4ym1UwgKUNV6Ke8botuG4OPM3r40VQDzKepCX0JTpBQBWxXLYMC7DA
+kXkaNPa9RNREHU+6TllzDH9eHXRfacX7uTjwLsYH+yMx0XnOxcT1KmI1S5Xd7ZQuIV4ilfSebYZ
tNGCh0m4ogyCmB27Bj6o592SJTxgVhcGNfyQAhBXeH439EKK2czAe301rCcb7RsW5NlOtCpEkX1J
mvW6xvKWNDGhaoyNbNWQ5D1xk8ghcqa35j/gMq28zxbSItq8d9IgJLc741v0RhEeLdsYEH0fBer4
hDfxeIsqOHy8AVqnqanSyzioZ9eo+YtNrMDx2IlOo3OJaBQiFfaqWYJO8xVTBJqHsOlMk2863Tuw
p9YInuMgn4keT/1o2NbjoZehEp6W5Nc/5hA3bEtUEjY9kL2MNYiEuS44LFQRo/xSf2RuJZkoaRAR
Z13bqHf57fo49huIDS6wYCc8kz7k8HqWOV7DyamTR48ULoG3n6GdOusPZnUUolKt4kaE58lBBk48
IxTBgKsoLOp75wZXGsshzd/a+plVL+ZDrxVujpS9GshfMeFRrJ2sF61lMjmW1kvJW5VyOKQX+onq
X4uZC7alOzK2RpPLa3TNl07512L3ps+y52QbPHDaaSPJkh3B+VhRdbGit/GsLK5xshsg4Nhv+YpS
quwUwg06v0e/hoJA47ss+MA1Zyv0UxKGrk5ZgWsbf3vBNUns7Y16/IIjPrJuv8DsUkEJHf8RPui5
hu70kBETicuepT1pdIvVPlh4Raz2qMynMSSWGDSI2EQh04XpCkFYsL1tOPTW6xX82apYqiWNXphk
dWn6QyZrxu8X8EJHy1IOc3OHRxHqsUi8EJyHVNddErLQ8//2JYPEp0TkEdRrjEB3BoK41oD06yso
FiGWdWNHVRkcqq13yErJXwyGmg1dz9dJ8XxAz7v6M8oeTx22yUTblAb5ohRYOm3rBr3EWjqojjK0
IiaWrVqpKgnHwlVC5HIrUYu9w1brQhPtsWZq8a5QD1BArZWK/MUr/nSAi7bK2HyMUOnR8Xhtk6Wo
gdNkU6V6C/U++7rh7nefcDQ++XoGSEBEtIr+NIdZh/oQzVTb+jwl63xiNkmtaQQlldaJbggmotAV
4EZ3NX5MLgZbSh+w7YXxLsDTaUWogOwC5yAjAuBu5SjaUIwZNulRBgOMONW6D+vJd9H3ZAevImjt
UrUn4dn9NI3aq8Ga8V+Nv6if6VaQSGB5wW9ZLvFfYcXt9In38oHAJbobAhwSvcQ19NdnkcabkxpO
IB6rbD5k4c7iKuZ/Gs/clzekI6yClKA241SM94GQpe71ltk7aI2oHeI8QgoEgCIqCEwL7my2qvi8
oBM8Z4robM5fOzinPuPeh8PUEx6j2m/WWtP7J46WQcsYZMcFRYZYDUcdl4RZWiq2pTqiFTHQN8O8
Wr8jxzfn/13+bllAL3G8sSg4a0ebQN0Cjo9/wjURD5NPRCZbPlzxNeRfXPI6QuUltek/SNvNWSFc
fM9lotxHJbWdrws6FnfhV8K5MrjlBW9b8C+Y3Fvg0MKyCT9G8i/rsMgMffV3B7chMyKyWE7ry6+w
HmuDk8uDXB6wQbsMErW69fyYutq0H2LmdqrpXuVjxltWyHOyjK7MZawvWwkyOaBHTYKUP2McYxTv
JNkNbKJp/jwWdS/Xh5y20Ah5493gXJzdVfnOLDF8XJAhrUFZJos9Qofa47phNp/rO+9CRsn7xLyZ
FO/8cNOAvqc/Hl3vmj7qHHbw9+OyfpIynIRUUmOVWzqB30KHLnLA/5uqo7ccPhPCjcEthQRoATi1
M0dkn/9ArrGTyEwMluDbSXEKLMwGA9V/pWH6t9xTTqGDwCuyXz57WFpx+bgvdQ0X+aFZRHzFR6TW
NWMF7/UR7JWuxR9+tPpTZ+V23L2XEIJe053al6Hk7Kf9o7zM2ijVmrOIr2ajN4qFCZdN0UxNVZ0r
coJGzm4YuKO2VFgbQ7yZoTvQ2mTmixd/as/vGChHHUsOa6QpHSBQFoE/5Z8aVkzPeGLPS14XTg+O
OvWFMLVe76rQjMeJeffcUlPvTq7tX35gcTdD4RO12M47lwi95Wd5Jp7HhqwfTZDyrDRxMBCoiW38
XW8wfikkeA5ivJczbo1/Tr9AmgyXoG4K6YW92fs6bNl89fHrL0M/aHB4zj8uuQlXK4W2vmqLCAki
gqTvjnkLw2xin8bFawxLXgnvaE4gOOiz5mlxDnFHjpnVNf9A9rC3DutH3gp5jlUd1LnuzcUKTKeC
pMGuO2eXgGuAmrKk3ajOXlrQJaoe6xaMBJCxgyJav3Do74PRwERd9ohubI8ebZTFHVhiplRoPn5d
dMGUe0MUkZM0e8tLikPfHRwgChJCGMmHzxmjq4DqO7aCir1JtX+lZkim8MqZqv89UgDcyuF2zVnM
6NJG9iEtQt4hrRJsJHrayZRohH8UEDTGWA5Xu6RnzpwEITZnibweED6DJr7OafIxFlpCg4gjWRCq
sLRzn8Mnw02ziiEm7gF6wS8BVbkZ2Hm9ST7evtaXW+4pZSV2JrmD2zg7ynMnnv6MMt1zwtMpYZxO
IJCYLShvcNSfcpjUKbcl4jHs6ILrI0L0rfrt9Ev/qDrtus5rdeVI7k0vfi2ihRbd7SQSNAVD0IaW
+6CRXC/2zma6ggOkIEDFdtaGe2mkTfe1/9pTwDGSW1zNzx5dkuh4qbIxYT4XvWRY1WFsjQMJNaef
W+JxDIskjUzky8IsbsUSLp3Mc9AEecuIYEdY+tjq/AXFt/YaRW4QHpS2v27/dxz25DEWe9XGmv4P
q69bSsenSO9NKd2vayznQHgfxenYB4fcVkzUCu04BUCzI1ysUBHlqUZ/fZiftg9CjXbEE7bMYDGO
8QGdbsS3b4atuoNVbdmGDbX+lV8O9NtWzabtAOC9Kar6k+EGPpS6gfDoh/WQY/M/HixwW1ScfyBY
eWpoGuUvFzGDI42cH41g2pVwmaPSTogLLCqHJsxsLFxmZ6YnITJQABzSCaRQnxrNS2bKTIYE5i0a
dXBBU1j0lszm9OQkN3wduZKYOHrjEZumZA/t+gz1+w5ZQSAB3oS4B3gVGFcQztJBdNZx/kSy41s3
dVQdhnQF8RuUZXtThPgB+p41Jo6wYHFl6c1g1OkbZ8olDKN12pZDy/GqIJq8SqvbezJOKdz+SZSw
x60RicBVFrZ2xrb9dZ69fmn7UjVAcCbjd/DWKD9Fhe7O+cLNRxzecKStt6rkFZfoNtCLs+roGcKR
SffPq8LS+ojfukpe5iRvph2gzGQtMFuzY2iejrMHWiWGmMnpfNPDYNW0B81SwT1zIeGfiuUJt7Hs
kmFP4WYPTqmtuwjAd1UaWz6OG1MHDTtwBqWnwRgBQS3OYwyt/rw+cP4vDnv4GQh8FbI3t/x3HgKF
GV2EJ2S/TnY3XA4SY2AQTA/OGTpoaegxleMHn7iw7QyJ4h+jksxLqMGhSpHa6/J3Dqf7KWLL9ghb
itjQYPkjNO60N4iagjArxmqEZIohQUJxhM76ANOkl/cryTvwdTzPSp5Xh90tgWOcYeAo3DCwpfvy
QRLvA4vnZqHxfXLghpsaglL4KqxQkJJiKQBGkkMokr7WX3l6e62n3qPmXi6vb/Q3e2/wohjcbBEh
/zUBxzU8moxR0c+KVQvj5xiLqZNHgkZ80tpoi36HJ3qH3hSm5c2PYoyYDyLY6MRwyoPfQ5JkNDDR
0YQ+MP0OjbC580oFh+yfNErMclXKTQz5U7gm+Vil9UzluDm0+KVNsGvZcd31mYHjjD/DqgaduWRo
GV9SyuIOatO16lKBe752GBnfxYglFOzTiGPfI7r2K9Ytq8otup9JRvahJM7cF82lfkLzOJoLOyCY
FGO8FyYzXtXTK56RaAmxeaITmf4PCpxlyDkbWGJbn4E8Q/kyn9T2HtdLg5Qjfbym1WMnrYxJgHVk
bj3fP35djTAn6zraBwg6trolrgpKF/VfLkISCeC/fZdppvX25T7OVPdo1sK+/94Tu+BDt/iPsQTp
gntG268YgZeqA0DH45PpYB/3VAPASILWw2QrBdxISJXEc5VjAvzIweGy8Nd2JGB00edpPWiCcDUy
ZtElHsXLLLrXgBxHCQ7jVNJGmJbea2Igt5g2GoMp3WgN7R3EHJlierhVqIKdNukHO1GNxIDzBAg7
C3Z+7gprh8xoMtxrdQYJd36580dUnPFEXlqMHkO5okvEar8U6hLn8cSMZwL2G4Uv9uESVjajKIm8
GHOA2NMZr12QgiL13DF+O5rNNPNREmBZh7MvH538M26VbhbOkI0Nr0zxEQXpXyhUSUuQGTycDjIu
Pc9M58pV+y+1GPLlT+XOQAsJvxMZxVZyb/ECUhDk+t7V7F0iKUzUkGJwwd6mR1trZKoxhi+yIsbs
RJMxHjAhVTW/R28EfHOCIt9uPvAEAGiYZHVLEpUOswCLUV10rAXB3TrKmeetu2S/mj7k6mniV/bJ
F88j2kgkptXjeeXjrppI9rILfw5Rg0mquvzkPuk6gczr13E4LpTYCd91UTNYtuJbqCuOkP2D1Bt3
lQamUzVwu741RJgCehG75V/7C0eS1UTZNXi3ue3UqlIHT0fkEDe5DAGxxO1evYZVmQqTtED8V6a+
qUCIgCyX5bND7IkJk8xI/AtpGGe6qXZZ0fzeI8LvgMOQf8C5aZG6HQN1/QH2yyZwb9XVtJLicnOi
Im1pOsKBEZ7bCLjKURIy/k7MmAYHGP186rUWvItCPHSGkvU0t6sfYOL/KF3H7J+9tQEL35cudEJy
WnwChSCHdswb1OmNwOl8VrhIvdQWbnRABMn6dgKMifQhoGU+iN2BjLdeomuZrsJGWAmKP8WnTcvl
8CpvvvbrxhKse6gVCRU2CQ8LZ+7PjjX2a68ApDpNU18RYIFZ0+4In+fpTNmSmfvjFkkXXp3ZEdv6
FIgKeCYcY4riywK5A0KaEbDSmRg0nuNV6LODIVzqk2ltQPNkQbnldJRAwY3IeeddoFvwOp+1Xabq
02Srp17bVoaGXC0BuxJXTRC7bND8G0KP/M3OmLl18NpNotQIb7/LJwIRL3GSPKwcWdf+FHSQdbGl
KMp7skEJ/J93A8vlvgupz73s+EPq+hwmQ3jnSQUBBGzIVD8cH7gy2e6MB/6deckDz8E77jOdw7z9
V0dQldMLPnzXWa8jpsrVoEj4WF2ytckB/3FJwx4XEJlwTg6T3FTC6rzst1tNLnIbNtgOY3s01NbG
tQXVETt1/jpHgutM103w4SAe4oubbgGHmwaCTMViG/S7qrwhgOl24h+byeRndG6Z+5D6GGC6crsi
OQAq+ZSvNu0M2UgPMXXII/46mmGhibpVHyd7GrBv2AslH0AjfThkGPakz+06WpDUowuwCdXqcXEX
lMPQWyvyoKjeepFO5WCalgfGa2xat2w8Y47tbSO4BssOFBNYGYl7qKcIim3ZhD46B4/FexA42LiT
jhBaJsbGbPjuViPEHu5P7dv2B0mXJQvqkryiElC9cySUpKN9oh3FrxtTds5KFKDuRIUhDeewHSgh
CxcuoR/1ciGk0bOhQ56TQ8u5dog0JWVgy7GbMM5jzYL6T1dIXMpEZHDVsnx/QcYPPhNRLtgrSbcW
CGA9P9CCSFKtj4WeqVUn0+STnVBjMHoMxRs+KFaMQ0kjbtiMSLkzOQqsRZ+tWoZrM6VxCQovndRF
ijMkZdfpX2OgkbH9E2BCj/0Axv+VmvXmQo3YXecGUVJF0UWuIs7mFw31t0hp2S1hqOeBLUt88+mH
YBw35Ih76Vvt/fvSJFdYjrN4HY6GaT3xMO0pjbzlm3i0HBhfnn97mhmkhceWLU3Dagh9mSexdV/T
FZFdmRL0VXAZf1OtjSRN3Cm4bkoqU1CekbSkaKXd81SVmpOsYO2AAoyAu2rigcYV2gkt8L5gvjZm
92ut9BWfhZXFn9rzGNvqf7VnSaJHlODe2ZuBNxv1Sreds/I3TRmekGxJPe48XERL7bpjgrCO0Vme
hSLmjiMWJEgtp1dnGBvU6Qhjb7yg8goY0WIrGyx8gbqzGfwxLp64411RB5rkAXQhU6BQvEcjvrCv
5+TEHIJdP36+AJLcgUgn3kT6bZtCfDbe86CejZOjGMkQp/jH1tKQelsUPPMLKbeKN7361EEAydcd
iGCgBp6rtT37+XUrV27EwKUwT/ji7P7pl8HoqltIqCi1XIs2WJVumMtWG/AA6OfJD+3l0iVWhkD5
yWIKcDDzBN9P1KhoYRK02iLMVJOAwHvp/A5/HXzoL3NyhR2RfWw2lhBCKmTg/xiLOxaGX2eaNZGK
j92TJN6YJzVZlTG4CtlgRruU3bYaCUDA4JryuH5OV1bWgne/GS3ictizUj1w+Uc4nMTU8ilonEsO
8dPYVH2jdnqiqqajAKxQYIqSGyhMqa+gg5D2xTaXJPI7FZN1DLaWt6lW40+2dYsVUS0q+g0nlcwy
3G38uqdcRDde4GqpHGcOEnPgWaZP/gPDemDDpUeDqB8jeR5I+Kj1twk8OVf/Y2040Zl9uvjmibDc
NwIdCBn/HLcBoFutiRtmrNp0oO4AFQ9KX670h+dXjV0L4FA/a0hyGANOSmfjT2atYYSLs5ajroru
lZVHckDvNdnuybF5uPtw5as1fvrtf4iKwsaICpA7FETLSNOuUUtTARQQQjrQg9AKcaeSPcrzHHS0
ULUOpJeNWzu7rAVbox4TGI2fVdnV0uKrZj8U9/hWLbPLkLI2D02rPfpTX0gfgnMJMY4RfaM7rcIr
uF5P/23t9Vfw0RRRZeYIliQDcRKcKkZWnSwuHG6SYXRI9AoxRCrAuzWYhCe1TdIsVVgQOALuI2bn
mtt9lvwx/o6cB4WKd2RIc0i1etqtF11k9zIn4wxqnhG/yb8O55QQ/VPXOTzQyw7FQAUQESvc8twf
u01E8GqIcdSbPeFnKGYvS3HeEOv6AUZgEoRvm93VtdzprM+d0ivxLLfb+Ang4JMzOJmDn1GTLNWl
uvFnzIr3dXvAFQ1AWkeUuB+ETBSVFMMC6Y93EureKfMboG+WfiU3HVr2VVGu2axfxNmL3g9tRQad
vufGRe/FASk7cozLZUx+Oz/2JgdCSd4z5QiBQe/OKWkbIQ57PXTUQO5FEwwwVh330ftPR2u/5Tug
KOpKRvSgUXLff6TMPOFjLVWveumex+kZ8wm4kO6Uy4k2HW8ARH/qaRX0etdk3VbS8UfZ7MkoR/wB
SGiGdpHV4+bGvLQKrMdFBA55KyofAjCyH8vFlrQOT8PyVJA0kv+A2iiIqcz2+6AWituKY84bxDmc
GdMpoRxuZJ3QBf7g9aJBW8hXn6JOLC7JBw+P5L6mAtPwakdx/BdPYcK5qx9K/aSts1mOdP2C+c/Y
XqiaAY47MkBafW9+VzdgnUj4umDgzp0nsfMa4K9/edHE46T3cYsP86G4n6gtEUPHMzaD1N6xnt+7
2CWryfB9vShvwr4sbSjUmk8idfxCKZp14qibqSNXdRAgtITeuPU2bg3QTy6NBVSgchJJ7ukRwViu
3+3dZ2JppUhjpYdSUVCy2JhHnlynKUnYXDbFkt9VIUeULKzAxQ3VB0aB/6pb58CTaAoy5XYDGNvp
59Khxke/cCf0M9dzxRoFLlz055NRAta3t7EhAB3Pz3jvmtYbxeFOhxGo0EX1XB0nzBDW3yRy55xd
UF6csMDQvba7RH79Bfi9a2IlShN7CCkvy2bLCCD7pWzvkdgdn3E3Wkh47d2IblyteXdftQnp7z0i
DXrBxDRMdwP9e3gwN3M+a6gAxmzY05d9CzncCR7vgXfjk3K55qIs0hbRa/HvMHY8oBMJN/uzTY6B
OEUF1bSNWHKltcLGDBGRYxOuqSHsAM8GF+JbD0kqWhMy+C5Qn84T3AYiTcnguszcllq+Oj8ojsY1
P421zaYjT5UzGVCspPpg770xJkaOxp32U+/PqChe688Ada7gszHgPj3lk0u6bzulNMBJCjDYtsKl
EDWsb50yzJvW8Zrk9YMGxBc1aoiyaqK0O5l+qfs9KuAGYE6Xmufj8nqchxr4nzEaWJVyqu217/9+
OAoMK8yq/+KMitQv9kNRAjZngciowzjHB0qISvWzkFjT0efPs0fQuXRjJCU80RS07UL6SEUDjQah
E8CDY2GICX0xkoBnrb/U6T+8BtdfjrkqaPtxhjK+MvIb91kL4Eszn5G4Mq6snuzpxZvYtY/rbjOT
QIFo5rn4Pi3tlb4D2zZyiSbSFMiBBULK8lz4OnBS4DK6SSmcIETt6/DknYFSH6b9mGsVFyd74Wtp
gwRpihBASEIsnwxBnQYN93MQ+YGDZDZTUwdu2Q0m1RBK+zf+Dtuvqu/YLCrPMKRjTNGbD6e8xHNk
X+9gGxOfnMDXC2lQqEwa9QLI7Yb0xazOgwWFZnpHJo2UYF5QsL/LVLs/aRuX3g/r4GBnwMD+RqKM
bh1bbuZkUyeDzVGJDrBXjBbZkN9lJwr9vtXUT8gAUPLElQnT+aAbYvx5Df3QU0MzQBEtxpxnUlaI
xng5ZM14NURR9sGZtUZEFojoiIPh0B++RnLqmQy7TfIqTB3295E28HJUB8YqzJ4nFhT0Q/F3VpuO
GPgN1Hzd+gR73gzZtn/lc8/M1JdxHfUmFD0/26MfHvK7d2Q+gorho2oLvRD1Dvf5OBPklaYU3hKO
GeChk5E7A/mgiQnmk+sZ1lJpThLavk9hsXdXAYMvKErVoSK8rAGZzqg5Y+ZbnbMkggho/EWZOKv9
pkO1T5hxG4HlfZpuz6scJO/ftYsVz0pw9019aALkrO6tHFaL3whjnvk2DgliGzZrcmZpumVUaQCK
sdDSX19KENL1MoT2cRSRnr3Y+kuMQYSRWJbplKfUFYedYxNUOHwMWo7Gw4M+deEeBJ+2YKVK4MrR
l7L9EVHDECh0sseGd86pybRY6bHU9fzPyaCIaBig6zKEw3Vn3hKRNHGO2pUTe1ASH+ruriu+1S8R
ETwTvznXn0f7/agtypTt7u1ACHYiGdMIv/PXJ3Ai5upoB+VqQSraY1TdV4eNKEPrECK0U6oIJLOZ
12K59u0nS8pAo/2lKM+2Pdz0zIK++PT+bxASLfNbL+LteLqRtLshds1HBtkCe8ky46TUAwSXQhLe
bZDYC17WL5UfhLTEut2SfRRPvu+koLSOXdGafE6YKJGCqyTQBXRFYiuZOosiaLeMlnFgg0vW0HR0
s56/PLqUuPv9U+dbKN6NupZ7bnkUl1lY/9b8XyyaakKUBH2VZlpX5fUIUgidxlowMYZVM4DpYi0w
I9bxKcO2M+3OxYeItppKLKHc8/VPYdL9lfN4/8R5D3lrOh/UqSM5fhUiw8Trfj346lMSrSrhQ0aT
A+iVg6US3p4YB+YaWDnszAQAUB46oE0iMGzpDAu/JphBBOBPFZ3Tc5HKWIGlpTn5/YF87sd0lJlO
qqLYNcnAnza2II9VZwyq3etWTVGuPx+CWW80k2x7HTnx34wCOIYk4iK28WDoRKF8CE4KQlxUjh9R
Vs6+VcQbmCW4st3Ypmn0wz9DKxKdAr9TM7fvl6kZJQLuc6mSwTON0dUOHA4Va34CkReTM+0QY47O
sljdjTtgDx+HuIPs/axtt6aItPf4jFkZ83woU/BQlQfeZhTDuSYmh/cv1QNhN/VnYFZybxc2HM8Z
+H4Mt+A7y2FkVmV4NhfnGOBHnB/8qR6PIZ717QOzNHh642RTB/fcvL8pCPemZITP0cpQB0DSTSAs
HBHj9mL38DOp27gP9Nl59IK4yD4ffSz92IZpRlX/T7jcQdZc97PMQ7Xgsr5zBu590o73e9trQmxm
Q36MtfQTCqrAmrLGUOKhVtNxg0ecOBisyt2aIqEy062jxsnt8y648FtaCG9XR0JEXghjOHDDNyzD
hL94coVELebrJi/wRJsHaTZf1Kh8FLLOLAcxADHH+tKaHeBUlK9ldUn4rU/zWZVnbxE9W8ZDAFa2
zWj1YSdUHu5lWxp05ufGXIjx8e7YF/SP0RnLRkQbPS4X3Y86ANnccnSkJ+gZfBrlfUYZGxs7o3rH
ZbHhWpmCg8ZFFNoK5gXPDbyWmr9Atua0MQZb+LRHD8YjBUCIEXTFExqj7F9PJQjp9/kiSSDgRn7Z
bfy3e4eVxFLU1v8wXd4DGmBcQDRPt7NZKYmNc1ljU4FrY4Kilyp8BL9XVDoNt2y0HJ2pMDK9ojKs
8yIlI92l41bVjk8wNd3dIXm5Bm26sMEizh7yehoNeH0UZ9iBQkBl+TiCYKXUjr0otnVZAMipTzZG
NwgnfHRx3QpwYAQ8df2LTceI23FYMS51xnL7U07RJllHam8UuDvkB07wflnZh6YVbe/NFYJ/5zwU
QD/pNBHY1eeH6LqPDS1mFN5chdupescuKNB3Q0aQMRt2cho27wa7nEGtRxicZMh4FsVDi2fkq0im
tot+BQcPXR2H5YFv2OciOWaFfVvofBJXuqT8Or02JtHNEmqjmYLrShVWNrDCAciNFklwCDohdEbJ
RTxynW7SJ/6d8b5jDNEYOO2e8WQFeE0uNYk+ROlk2I3GOn8LDfANuTlWRZ4mJ+h7mgdPMje8W1GS
dLLKeoBeegdPdZoaBTO5yYZTZzEBFeH+eN2efi1wjpLyz9yz3LmK2VGQJC/6+edC3fkvZIfimUO8
GOA0S4NSBCKEf6gNc+iYgljiEVt3M831kSpirXRMm/GTqvNbk6bYMPmzqzpDzxtINdXpSN/4c3PT
GRoCPYpT7EYs2ZJaNf3F5fbT3g6j4aO5dz+/mAUnhlHCILaL1hngDtLM+beZ3vYO5cFxfACSIKXw
vf9s/enFaL1v9emE+6v/LGQouEAa7Ln3QtR9MA4E+XGLxz2VdBVr2TA8TJbmL208cyHLdVb+ZBPX
ZADzU07UgmLxXOXLjmLpfm/YC8HEb1Fea7s325FxOIxsEz98vz9mIV/j+lBDgsoOEJc/oO//e0jV
pQqMxeRFGSQOLMNfZROxEDwzo0POcScPcsXa1Sj55jbVweUHXJfHHYY6+jHc1dPOM+61kU3qw0GG
WHE2i+myhM7LxWzBPlrXV6LUisNxTwnucA2AWTc874cW4j8Dua4r5iZQ9zM4FVxz0hBBtw9m7R5M
VySotd+o/+ehaCJuN7ACvJvgEmzmtoyvBAzB+iMSb3b3r3ColgAwJP8Pvdu3ogMgoHIbStQ6tDi5
jOA8elTm9vil68jvznoFZ2o/oTHWwuz6DuWLFef6Oi+s5OkbtBNR7WHA6/iQeiH9nha4V0FBJpnX
cKJ3gp1D8+Is8Ct0U31uM1hFXu0rBAlObyTEqQUl7xFqfTYEnPcroRPNLuji+XBMk4u3Lr3EMSgf
71RSWHshAOtt4vNI2Z04FgTgO2dq49Oe2tE4snuTbF8LdbMHWRbz5Hw8cqi65nZdtzDVH/LdFyyc
qWLXaWbe0j8boUdQovOnYogHSqm9lVJ51Jm0YNyPGYldHQkI33Wx0rwivtm0+y2dQoN77cqWg5k9
V0DPN583U0siiSZJXWiqtvNsGXrGFc8RWw/ZX4X/qAhrhIZuNZ/Au3iNhA1e6l+HKEL/+GWwu6yp
wcrDwvaTD0K+lF69LY0fz4I14wtdqbOm6gspOdxFdqCFBs+TeIc6U2MT17AcWPKHwT3BcCoQwtDV
04bHY0wpdgYSt8GlfCtRSn6SJtW7S5mfkm5KvvmFvwC8cG7Lw8faxA3iSO8Y7C3qoEbS9mbXqjLr
i9S7APnL13a6RprHBbilLLTDKEUPbNWazonvgUnvN5L1NlZ7uDRqTxL0JBujZyY80KltX4+Q2qr6
Auxn1XnDxnKFCbJWELZoDiPBaoyzNPuHoL46wWQpK4h5UiT/yOExARM66xsr4iih7PM/X2vTEyjA
9ldlHzgq0NwNg3RjEOwhK7xY/+amU7MxbDAnOVuLIbMCBMCYY7+K63CNEoqzFmfvqWf5AOTZ6LRo
Nx9Ln4QqLxj+DD7cAwPFPNMPluth3ElCBNAIlx6QdelU4pp95U9WL1+8ZaY5NjUC2iOFrlfRdHVa
/m1cKAlHqQfLX331fhBsk7hdQ/yMEGa9KtB7a3PbP2UTZh4pe0yaUIS6zqvgryCSfdjQb5Jo4Unc
pPHoU5yd0Xk+6+zpqQtbjxw8fFhGXbNiMEU6m69xvEqHKsKsDDQ+T03J2DaR74f2FETQfl4CRRhK
dgH65JR3aOqMeB3Te3bsETq6VSXqwjacsrE6Fwg8yy4vCHW/u4kDujpdIbRlJm7BBlNWPe2sZ4cT
agjKFCFZV7NZZ+G28tY3polnH2nIGJYsuz92yQFfim0SxjlbXmm8X0HMPhACFG/UGs9fHVjGRblB
jSLHueVT36sWiRdvCUj/cjzS37D/KDy67x5bILvd4t/Qo6xDCyByXOd+aLmijS2mDlVnRFEH/LXo
zvYrU5FKrFNebEOLGbMhHhnNlxg3CW5rFC/2TuITTox4zhIPigAjBklQYSK+4GOPfZm/n/86hI0e
dgvoo4/9w9fxClbWZaNRoUdVgjnow+Wafl7R7cmOa0pt1Q669bEK/TuLGLjyal7emb98cT6yn3aJ
pNprkt31PXf200D4fJWN5WLZwCHC/oMMWmmDh4RLi9OBTY6mnBCZd3p79G+p/s+4n+1o6A9qH5TO
d7FjlckjeW1BHDdkRzpfTIp+GtEXHIeao9kjKiU9KfIEv8PFbXmG9jHGS2vRzGj3rA0FnMio1NoF
jOkfls5HZ+8JiIHPF5FCS9lTXD7Mq75nysK4n+Dfe0DrqQyBP7ubtxWFMPgv2deaG2cthkzN4oYC
FssYHzLWhTv7B7Isq1lva7S9AJaE1dMHSYxRcfLBuetqVptz84sdKLh32lWz7zNbib1xl75AkOff
sl6IHNGB2LLRmy0EeU5PrVbqw8urpa4p/RIiZDcPXEvMUaHhwBQ5T2zvc3eP6izWOmVMRGIWJcf3
8BsfI/SUqHJxRI9CVlb+ME0rRjKvupBXmB2BJ+JX8KQy2Br8EELUlfWojy2MtQrYOsmlVmKVm6lv
67W7qWjbl/kW8c2DRFgYQFkUK75FTJFpe4ZfZ+hw9wxZFf98gF/T32zsEHKSKWZ1PYcy92YCwLCG
KlHb8684EXxxEM4FM7YeNzcgWmNR6MFWHoBgabW98OHoaF3hvdTmgvL+0iDPCamkNCFuzumwNg16
ULFRlFPb/4u0SyjWSeemMq51dx0l1N4sIZLeEklNroChZw4u/kWVFfc4psUZ9qlkrUk1n3MknuMg
IecyMbi/hKaRhspjWeX4yvwdV5XFA0aS+WEs3N/cTWEX2ybNO+acYNUTFlJ+qybnIZOZTgTQuVbs
nk/xI6fXuiPnjTNmtZLqogIjNKFY1UHuPf3ZwD5Ygboym9vCznhiH/gXR/NGnZs5TrRuucs2fw1/
DuX7PxeFx3fgzpeJJ+eeuc1LMLFJRuTbPf5s+K7mjw6V1OcTpD/bK0Ul1Zm9d4XRX/wlFX9/bwYF
PZkxTD/gVUGmcS9GxBXFX+HYs+TY/GJr/KiEXAhbEKJCLCuLKrEa2bzvkZeGdxPrNNaCkNt/LOpd
XOYswMURZNPxlcltMgYah0WWhQS1X0qdpMT1KruREkpf9PfR9XLeXQeR5hATx6MAZcfTUYRVO7Iy
tbntpOmBJqroXTEl+C56zFNvs14j2upDRbdpKqUr6IW1bAPAARmaIjWCmOFNtLCaxahW4kZ3CmHs
Xy8WmDg2BRZCvCA2I+s3OrKWQZQ2s+sgvubBMkcUl5c50X56LQBf/AMxmgnneRNWdyGDkFh79cIN
qzFLIHNB9YSJc8r4A/QdPZnfRZwcJFbtdI4pJi8F3G+kUntXNxcVwakzR2giH0mkz9+FFYuBh96R
OOwvF3Er2QNtInhMHURb6vq93/7KKb+0iiLidyMshjLzzxo9XWChQndYHynjaFIinrAvff6VZyl5
2qrkgWu6pTXsBNrrrtE+I/Iwk2tsvy0nCJaSOGYeastde/dI/hXJ2pbTDb2mRglyLgWiq2ii4hkg
crKL+iKbvfYCfVVbE5WNTnFMqU/C3XjfZrecw7hE9YUmMYwo1FoYU9atnEH/bJFdhlLhDVRMIrQ5
rTLyEows1hfJBxo+vJVnmYuLyHKPFXn4bTPdu/Hl42qf3TPNNp+xavc19vs+xP+cxbgsNVSUuB+w
0NgaJwuWIgYuFOwykPbXhGm68dPwmtuCEP26lYkchx7tJHUJVvQTXPTg2S2EYwBzzA2hTwr1TWRF
NygqUPKjgKiMwt9cqoBos3VGBylv1sMstoChSOUfzGIw1iv3c7d4PyoO1Nb0jpxogeyp6r2RVabq
VZBs/oE65iYBsBCF8nRQxOfOl4iYmVyrSvhMtmrUpHRSPGSMoh0/Qqai7tc6Gsv9NlowZKivcfBQ
jZdapdjpNGBDY4EBsjr3RVsozOZi/GRAITE1ynob+TGppXSWSZTWzbd0KI61brDk1BQoZGx/9SWj
Jfr79QIpiqPqan1XI5qzloJl/aNVtoU8lC2s6o85rCOKNF5MD+Rrk9gVf+ftkprZEpD1rlOrskZJ
Abxl60vs6OyBLFisrnGrE6VyzkublZ8LWKr2SZQVUtwlTanNXxbLEk+yKdRmFBBdll7wufRQ6oqQ
9vORg42D3SRiPKfDk2cpJUdlfU2zvY75E+xjM367Rucb7VmqBe8Q0o1rIRvPN0qNRCJhP8kuvwYn
cTQDen2dtx/DCzj/Eg3DIUakc16GRqlMAudytPyL0hl+iMdJs8UgCMLmcHxe8PNiCFL/0j+7vgSo
zCDzTXxbfjWgp1BdIETzbhYcnGqTD1bLBiiKHOQ1cEU3hNeGypbucqsN5rEZ5P4PcDnydPHR9Boc
8/1VIzHRmsCmGhc3ZymXMs201adIAgtJKtqjliXo4d8FQ/e+aSi90otHpI4AL+sPq7mNWlblaCJa
ufPQyRzE4YPCJyodF3TRsBYO9KnKPKiocBRC0ZaVdEQoG+eAqEsUUKlwKWqf78ZIJysIP4v8jfod
B+XwOQyRLKUVI7gW/+Sl7Y0LCSKclbUWafAalyUJGwzaBRayu+jIYZ4DVwYJmfSFd/4e92U+WD1t
LKnhvmLN3pF0N+lA+Rjrwk4oAwzVUtbsKF6uzgOv/7FFpYs1lUPTzXcxTLbcmIhkb9IpYKEKDLZi
j8xe2qgFqW4SwGp3m5i+vzQ7N0fIZrmyP42LGGuiBCOZtbvNjSYCm+pXyYa2gYacXykkgbN83JaX
e6Cc6xsjoi6Tl1w9jdg7FgWVygOe1gN2hPJRCfi95rU+N57fTvbA8Y/fRiVyen+hQEFpcwih29dR
LE9uHGpun42JSvsTM0HFTm9gPuVHpWYvb30+s16QMtsVujRGVS+/4VzFx3dxoNYJ/fbdGjNtyBvC
qNRpj9lE9GBoIX1GPj9Im/8dIbX2q0FAIYORU5oyKcbPB29HTft4U8I9pXK3GaEO/qNrqA2F5E3d
+NXJ2hx20TtB/1QFYSIEDqtxcHUP5kFkRBMjxGlTrJmUDD2u6nSdEsu+XOaUe6yoMYwteIL5ryLT
zwy8ygr3Dmt1pzg9WYmnEqfoL6boiPGEsLxF4vhF36AduKtVppnTsNuLxz/i8scCqe9qL3+PmpCO
lkd8nVh+AQulNFvRVUw2AI1O6j9Gzq1zMaqzlI8QzXRUjmAyRKj/WojyhdntMgpB8X857GDlKfNG
xXHfAxcM7sZHl2hUrvfib6nRWAEhCBlV+KYAGbegDgyWFuGxkykjSDeDYjY2mzvnJ61fQcHC4A8k
IxIGdl3636q0Ktq98/e20ihHmVFhv8YKzskRfhiZQ0ya07nSX5HqNcZEzWH9wx6OBfS89kqw0eMo
jpUFAhXDen7iiCeL+sC7yYyUgaMeEZlWRpqLHRpGE52zGzE29vhxdUdpBQjm3EkUZh0E2z6GFZMw
oSSlEb/aY+02QqLGXyhUt+e4ksy+nzglqcY2Oh2xTts/NyjtnyKRxmSOh67sdftRGjVsX3EX+Qnu
K4V4Vw7OYwqaT5A72w61YYVydFEnkb4iKys4ieiM3lykR8HIyE6CpUM7MJ0pqqAy1tHza21+AQDW
nVo5nnSMozpJsXa0fdp/az4DvsC05JL6tQVJczcTua7ZIofjwGVfRauaXWv93GSaarlT8lf1jbPH
wYO7CQDtOpE+V3PHxNgnSnOJkT2HPdRym7hEI9RFwotpsRc4Nfuf2WwRYvDKZfDvirDN/E/N47VC
9IhQcdUfr3jzaGkL9oyC+TG50FcVIQoH9O8u8St7OYHNFoLkgjGTFBWJo5ZTDkukw3gInKXamGyK
kd9a0zne8aTeWB2inLO6/Cm1kM/56H29NpD7jd5X/rZmW8C41ioTTLvfhH3jdCbIpJSV/E8AZ0Y0
eLh0VTthNudzPecp21GwzZQiMdz2/Na7jVbQYBT/KIqquJlrneHEb3jIq8keGkVHXadc1/r45DU3
SO5iFAObs8s5+4gaTnQ8NS/TZisCJq1X1Nm8QqGZoKm+s1xSc3mcL54qvCjg/+lyw2JtumOkWXWy
Md5Pmvnnn4MqXq3Zq88IWq4jdv2t+LWiZ1Qh4TiQPOXvBnsutiOshLXJ7sKR7JcKvkUFyiCCvehc
x4jhrnJOiHvuKB3kWzgxp4Vrd6PH6Iez0ROlQmRCGu6nPfV2GXx40/rYoW9q3NEqV00d6CpvB6nY
1D/RRy1vEh8ROpQuzQ60aWFX+q5G2PUpq0No2C79fF3AugPvmCjbR/RcACdJbRxJQAnpIh8D0ukW
QuBx3N5d6s1jOYAie7Sca9FgXSFVo2yePgAg1NJT3UvNK6cwvVGeLHEZgjVwU6uTl2hMIQovVrPK
Akp5wO47aQ9YCllsKyAVHk2qb2JFF/4nekKaG7+yUxP7m05wWnlSue0db89bhrTPaB1WpGcRMR8L
9kZ2M18xK1Lyr3QDtbwCQef0rLPenlX4Wajb4UFvnFWIiqtQla/NAHP5GEnBC5q0+GacKBLlaemU
sNWkGTv5vG/P+rMn2mNiprov9WmxwBXtNs98ggN9M/hU1Seq3Pj6uuZeHfPcbBerZlNg8xyihrb8
kLSu9DhIMprKnQnbRjv/oMdn82UC/WcQMfqmGzeUcc+otddIQaBpQmFKldg6gr9uoahXSoHPanLC
QNnezmmce7Gaqme5Z4YCTF0Pu1zO0GJ9vch1FVwSczOunvoFUOveto2uaFCHid1DU3/B6iI/5xVh
2rHfdKBn5LVuL4XhL/BeOt+RoCwWmqtl+P+ngXyo8Q9/eUFahKOA11DyEqJAVhPx0+83yTTKEtNE
OeFbyuXMoObJYBNbY22MVrA76WPXRcYPvDtYahQ2hqL2Ro1Rf+QgCA1g7maeLDZK4LA40tWl9vuO
kUqha14D5lp7wtf8lNDZa/58Wg5/K6klxVZfJxEuXRFyiYVxT+VPgCFgImu5xykQbJ4cj95KQQtM
KaCaP3YFV71uGFdR1pdr2kQmWVh7B53VZcEMz62WTbKnY/bjOojmBoZ6aIDyaMR14rZKChZZP88F
+ovP2DK+u8PRH0h/Vf6DfusWbXVNn0bqnRqP0R/d+UaLbxdKpv17JxBDFRcGSYi3Xu7Hb4K173vy
8XWWcJeI57j/LszPUru5cr6bi/QHGN3UOeSSiFSaKYuC0sBvRa2wILXa1zHq0ILZJ+9+61kr/oQs
/P3psl/omhLEtZhqwYTaA/37rU+qWYHd2H9KfWuExQ3tAzF0b8SIkwXJ1ZS6Z01atHbyyw5oEEpC
VnbeVxJSXle3RitHNiQGpaLFWiMNQoAM5UWNT09m5ZVVyvNSHFzhjY9wRWqSKw6afkujud7IsBtM
2ecgk3F/rUGlIAepsJmb3/tELqnwAgI9AnnRXiyv1ZD8rwLVka+eJamIVHe817uawzu5ZAUQejmu
g8TcccRmTEUYWjjx4OqsTvrMRVV5dowpB6QtaaPSR2nGU24t2lly5/0UaUq4aw7koTa9DMa/fXxw
fRQ7IDzecQ77GRTLDh7R5Sv+JuOElah1LrCzHy4l2v9z6fcvOENLo7lZw/lUIpxKTQTx5dpowTPM
0lhu4zNDU9y49tnvCMcdFDo82V9+PM/TEE/wGgDu5t9tEYUODhAUpLuXfK03/vqW/3TLN/dWZ2gk
OkM1qtG/1dEF4wwUtZW3we5y3qviVOvGLL3yW5+MCiNFWY24fLpGEWRwKFityRRnDJLgsQ91nxZv
pvNOpchv9HkkZWEijGh4PMXKv2UeR6/qqST08zlKAJTRrKsGohCRx0HJ0u05vxGbIYSO4pupV/pj
WqXWHAGrlCro2Njee5ad12JZQDhAKuHJkwhx1EuMcWzi1/FBmL33oy+//Q20el7YWUxAznRRhqcO
OvxqUp9OCLz6XE1dsoCh8w/uo28Whnaz2naeoaYx1GTAD0I+iLTA9D7xKwnpE3t+Gqp7MYPjFH7R
y/I7oVg+FqJpPuRvsniZVqZRCt9qOjWW5yKdknjHsw1v4J/xrNW9y5jGEFM8CfuZRG3WvyPosJyA
IkrBRs+sdhnjedy2+vvJJ18UZYx2rFosDdMtLqA6BmhtQbuB2uzDU5IuHcCebGDCY6N/gdmNRYd8
2Y63dGzyHPmrhycgakB/rhaFpXQPyabE7Pt6+cTLS0zmUP681B5eywIk6C6inSdxbHLRfhAkjnDU
JJ3ZyLLB8YJEZ1JKaiYzztkPrkRLllgKcwwzOG3gFP7wPMlL/PsufqcV4+zOFdOmnhKocDhyBewW
pIgUpTO2kSFv/Rbwn4kEzlBHMfIfIygOVJkajTYFdma7Nw6hAMCNnx/xibTNrb8WMVpU8Lg3Zsg7
3T4J3vy/0HfxolAZv30QyBxGR2dLDQIVTxHI2nVYJgoiFIcfH9XiJ8i/aDJb8le6JpLH9vUdmmJf
LREroJEA2lf8QQV5ADoP7VZ4jjOEkdPH/kw3jnyCGXYoWLj74zIhCsKFyVV26jC38PAayu2qXh4m
TtJIK7WX5QPWaeov7Rm4oRwiihXylz04WWW46/+joQ2SYKaTc3THY0Y8pLDLgAuWLEXGelfJk8s0
RYLwTuM3hiSWNtODstSr/HwY0wGpklkgPITB+KRo+ty/9bMHPGwG1wUzt/8gc5we5vSXxzwOcmvh
8mZ0kbaDIIEmXGV1H4+32s8xb/Nh+RiEHC5JvyFaLhpNHDzc4ePSIWsQQLPp8iprSdeov93AkEM/
JYcFdfkr5OpkPU0LPN+ogQYSho0vTGpE9uDgqkry0oqT0qhS1uPvrLzx495lHApEVgx3Pon1Bl+r
weTak2F1jaEP4sZwr9y46dz8VAdmC4frZtgKrHiOxu6L5yloB4fzLdrYVx7Ki+9X2oWTq1ra6NoE
nqgvkW4Osb7xcQ/K9e8Y5oWGEiDPfd2EJPhr+7/Fsur+eSTOQWWS/KGfEt/V8QS0bi2R0lnlyL5O
oUE51C9F0tuKOiBlo0Szr0P6iXul7376nB7/yhxk1RxUFp6cecVLXoDPCsDfpF/fp3bO0ymcqBX8
D8MbnHh+5Wvbev2WSrEQAVf5yU1UcvfwERbO7BhscPLZoMB+3HQtxrQK+psZ+D4lF/xLJRuXh4TP
tYuMldGCkP4HagU3QuNQVQBBXdtwM0dZi6BwGzkui7QGPapjc4WqT5pU+9zXRDgdQjH89garRpxQ
+w2VkXyVKDlOsPig7T08BMe8Zk8xflBnTZ+g74sqQGlX7wrBO7sy5Fab2qNE8ysNscQs+qxjxRVk
yB5lQl3Euojmsc+UPZyBFyYdMJI3ogsxrimvBGufWRjMeFU7Fqh0r7yfIiDM85ofRSoe/lanThdT
13tnGHCMNB0vVNxyC+pGusCmu1eHKSRGpdcGkjC9XjszNPaTCq+8inaUJKIXQj/qRhci9iucDor8
dSChEMLSueyQDrBk95lJELUNruqcVLCBr7UUyUuVliOK3mmBsqWAcTa8NPw0/N4HWzDILfKV87Uc
ktFqM1/vU/gCwr9HC7UfTHL6hEQXecMpjcprswDjSjnHxYBnXB0/ecPeIj5j3nVYetQDdvS8uQWQ
nUajUw1V30W1bdI1zYkrHSwRwwMETyOf0gqkcg96OTZ7LeF0vwzc7O8o43wtoH1Aj2aA1ZLC9Iou
W4rIjhd77eBBZB1qef2+F+Pa+NwFvEsQUTNnd2M688sdDznheHwYr4koBZh4M8mt004pAOZTjADs
ZzH5nZmsQKi08MYjmO9dTHpOLn/Qe4zTNkXboXIT/hEmzy6yCY+IDlLrTC3UXTyXPpQAkdjrgH4q
o37AXZ0mHzfm9K/hgjTMPDIu62EHmVSfcCP9J93ISCtGr3JV7AGfPG56f9r4VqUWPnqNG8iPlzdf
Qo3fzjiP3L5667+Tx94I6nPKht+uyw3N4iiQSjR4Mz6hQ/oZ6syhC9ZBy4bdzFYwkEni77i/4iVz
Tj0EXm7PAe0P71pk2LhpFJbpkYTOsfaJUfAqTRkAm3IwS50vNj6cuCkwNWRBoxpp3YAZVVwU4YiM
fXkFhEoEmK2N4xOC+eH/n3iOlQYjjBZVSbGTPCalcW+JzY0fnbeTRPwSN0dLzfp8nkVq0TCViilY
HaPF7+/1ALVHpqSkp+h30//FJ+ePNkP5mcwHv0ZB9mnDcDZCDclu1MMdhq+lYxKvJ3Maku72gAXN
8czAIuNboChd9nDeNbldypJdfv+CxNVi3vS9+vM5/LqwT/THaJ6Oe9OxUDy+MnG1VdobC66LD3sh
vmDFBvS/HbMr5XTyUmtVK2Er8GVbRfC0fA811q7LtKwbWO1j7jLRx6LoW1BcFh8+U8QJjSKUmWN1
+bTwfvkocRuSWKUu2ZCVtRhkRg/R3QUWHJ0e+lfTiNLLeCBdeMw+SDx0UM7QzNdk5PfoD6qioQEv
QMbOt+zfyeSyUq505en0gXuWFcz6g3dwuDVFUuzR0yk5KpjKWT31J6wuOc4Ek6Fo/Bp4vxYAFhid
Ei2K3VDgWQGEtjQNNTSH96z5WlhuYsxLHTazxPXh6KuCQKYLpLz/kBDWZHr+HeW0vVtxBPyeRHOD
kzAJqZb8pcePX3SnR79oC3SFiJS6ttVJa5mt6I611dc2vPkUWckha/fTvgx+7v7ySeUNoJgkInqN
Hg6Sc2zHQw0WtYYlli7VWb9oNA/KMszDPIVIN9FAfZl3UWS/RFjZ2zTUs8y6R2TemlAEBV5vXJ4M
Gn3qE4RhurWCTm9OxvnNlejJ+SO+v12pBlijKfMh8WfR6qJVevfxZEZgWRh4QssI+bR38zOmTSoV
sFX+hnbQRzdsIXeI+ypBFijz24Xjg3uvhMlimHikL7hpafrLdMPnNP0LX5ykaffQl4Ms0+iHrNU0
Sx/b77chjtRFSWYwEMoGtcEIdWgYR1UGctToyQPmlGEh5Kj9+fdbEMMrIgxj3r7Q/+xsRgv42Y8r
O6VMPFnx9/NngSe10kWK6EVIommAIxaL9QWDyuQFLAfqHYRLi+XAINoT4BLvQO3q3FUVk8RKjSfQ
flJHslf6eMHqvoKqRIMIlXxj7ZjMHGRu7X45Z1Ko0Wvv11ebL8O0P1fS7bUay+l/QD2ENiSJO4dS
XAQUsSPfsDyGjyu7cJ6zcWv5zB8rW0Bp0iLEQ99XoXdzqYnrsdcsqaKAB+mOUWCCg9qAf31997go
bZjqhDaM3MRB8mzVnNVr02HwXSY6M6eR0goCqJwOrzPwFstWNeh+p21z8IrDHpEDiANmFRF/LEbb
v8SGESz1R8RbjzobG3U+uS0oEPpmOcmi59/XoUBNePMZ74uMeS46VKBT/CCkFguOxydS6MmKJ6LV
KrHQUuzGcOfW426YhivKq1E6kR13aQoxhNdTwBPqdrX3Mx/Myf1UZKiogKu3umbP0nsDKDyrN+UY
0O838kS/Bskng3QV+LRyKxbYUpAZhEFtwFELR1h6KnlKh3+PbeAgTdP1pqgBbsQmXDOu7OHWsBFu
ipfLrJGQMhpSnFdyBnU+1/0aKzwIP51I2HITSZBVGHajNefbu68plZ7z09anQluoUcJWLhZ8Z5Cd
Sr9oXjQ5D0mWoTAGf+s4lnf6kcBQXDvNdk9PH6GFgeY/2rQekHypcshJ8rkqU2SApEljgZoPDkGd
GfcKZZ4VRzo7T2DJ0TP5yGXnNaQKR+C4cpjQruuLUcGz3aW85zxDUTCsmW+mYxGZ7rjWiOGN9gdJ
ywQjNyiDI+h3CZs6BgdeEkXIG2iX67FpUwqd/yCTYSAEk8TMTdJgfX6o6T0kHjtf8fBlWFOnk+Fv
r8gpou1NdnyX9N5jIN8ZJancEZSGZAaj8FauOJieVpUNS/OSxELohIbfLJCMaI0QKLx1jGgf/l25
kALpXsSz9LPoaIXEcvRFSSX/0nxr5CC5pxQFTcHBjSvzK4I9BKoV51ViCXKW/90H5dV7qKuCArW7
UsQR44yIan4Nc7uc/1JxfUOwbGb8o0UlKfL1vcn2T/oUvvTJ9/glkhcmSEh+6fbNMsUUD+SqhWyU
3z0t36AD/q2QVbGvi+659jH+p96NlMP5zO0NCqntFbvAyQ28f2KNqY8rQGZklMLK68WPE4GstpeD
dIac7lOjMvnpHKNFH9HtrrCo/jAhOrLoEHFATRBJKee2cHh50pQWW/gCjf8lvwkop297TCooc7ah
mjRvzBbCEmocoKfO/mX2mld+shBVbtUz62d8GQzRJTURPhkWbv9hf8zlSlRWRsZ2WOfPd84HM5G1
aiPGzUtYWhlbXP1QKPOgzqG0IYxKyqbE0zbW15r7xx7fXIBGuN0zSU1N/RhO3VY3KjAX/NTB4D+9
LkfW2z4nUFfPGiO/lfaMX5o32N9cowZR6jwG4YqablG+rFOBM9frcB83sqVaXYgVS/+EwEeMY9z7
sdojP99fXgrcCYOBNuVH2qja3U8ik1Aj8loy15rqnXnwk+6d+GoJu24Tui1jA+mYxpSw+Ff25IDu
iBzoZIAeieA+5l8nEbU/FM1cD8Ej/ejq/6+cAU4hfctB3Hq2RwhvW2kpUtSVtZn4f1dIsAJveXmG
+7eHqhCUviDOberKaecfeIJdVhtgBktzy1sesqDanmAwmEF4S9Wt0sY4deckwJIKm6AIRe37ILAT
uVDMEvM073EAc97Po2y0YgcaqUTawkDEZ2OebpKL1r/Zg1Pl2mWNA9idxN14TS0oUHvImDEvvzPT
EEGo64QHGRRiZREIAuM02n83kpRcmAQXuSHB/DY/cbiPO3Z7A9y+RbpyyKQRZQGjcqiOa5SK3fSx
NQZqN3WUAxy6Bk3utq+Go4wGAOF8jrClx7F45RaRRe88cx/ZBHvVLzi4qjnwfD4nZfwsTUzAYDcm
PP5YcscGOcS4IPaL4+ZPEjHBJGiUDh6+2NShseIvCBMRJhY4hSiHfr92vs4hQC2nHgQAV2xPm2Go
ZFO9u02p6Y/BSQNPivgEYqwNCv5+XtPm609YW8IdHLKQs8k7MdX6kl3u0aAKo3MfRK2Zg8joSmct
qRtevAyhy+FNVdEGs3K+tpCmpSJWcG5fYPpaMwz0yuuLKxRkjAUSGGcTtGN6k6V2JPAdMP/68q8J
4end8MPKnuhnFC0aEc61e3F1zdaqZqygapwAcw2E8LlcNZae3YnQoiH9AH0EA5la7JtZ5Kt+dFTL
oJSeAW3Nhnq78mhEr4t3jNxeX3MTvX5gdZQfTsPlgWaV2YDgtgu3sC4M0gNhU7x8hK4GJaUsf4Iv
i+hupN9q/fe+V9hXzv61k05s6Bp7W3kc/VXoLGlQNAfXHvJwG31oZztM5iwZxQW8L797l7bgrr5t
pPMofwa+w9kRVb6mxIm48THqqBOD3tBVygjegvj7aF6EicCIOCvQwByuRmxG4iLmpVgfaGzOHEeZ
Wcnm5JW0lWjKHKQMd4SmwCv+Kv1DtaY0Xeoo6rF1lszUbRakxLZkMXwgiy8ECNurteIoDunccYzf
zQ5MQ44JmNaQ0tBJH8HSOrLVC4/CVzPqr/f925uzc882kvwEzKhIeyy9LaonCKfKTMAGwoUsjMCD
p5ypex7n9NyYp8lZM1W4zgrZancJ2M9U0l+Z2Jawq/RRS2o5IoYtCDJusvmguK3srxBVyzzRl8Km
feB0DPvILq8nqvf2pUQxxgvAHGqXhvJ6YKlP9H7WcJ6cx6O3Ktek0hgPW3Ic0GqCaDkn0av2Rcyy
GDFnvQm5h5ZNdLcN4DZxziCxRD1Zct0CsqjK+e4qZJ2y/sz46MDZT+GedIEDDtcsfE5ghxvF42lX
EbrZ/iCzm19YhQCqhEhfWG1fjYHb8luivMrYho9zed8X35AqksFYrZLC3DZz/R0sHPcw1y2+7kuB
ZLP71SE/Sfb/yTsNRD+3LID4sfRRpHadxT+f/dQ9oR2/Vb3W2gIwQP60PlWGNoy2FwNBaTcahLab
MUOl5yTVHDWRgyCneWB6vHbif9LWueofjsaNmpCRQfbv17dpunYvb4fvy522y3eE3L0VWfjWJ69S
o6eE5gc1plKp9dj3+6E8/xtmNXz9x/Kn/DMjrCxopIamHnNiydGQuELTsUJcQQ89aBiWKGj0v2in
aG6C+Hq1P4eJ9eJ1S3/blls/7ELAPrwdRlMCv5v1txrz9GAt7qG9HCRXsASXulbLIXvsN8ImrHQ4
7ShSonms9KDmqJO+NmS6G/jNLHB90VmcF7WlDwaOftpnOZ3rUuwSvMhcOjr9Qy37sJ9BvcwhSEjX
AZIX1j0g2yWSKxfJfQm5AHPnsfA8Zp1CnfnoluaRV9bvIq6AGMDvNkv5T6BQN+Rg2m4wx8rv08sd
DWVLy7S9KL6on18CSYVElPTxMysGgwFy108LGwkihTY3w0KTfmm7qTOjPpXMeIVTW9Vur4sp+YIo
DJgjTXcOPwV0LofmLIp2VvKc0cFIxJ9+g7a77axiZEe+CcpBcMrbMubbRRyASEF9AEGkxVk4Cmqg
ltksIvuk8QfGICj68jk5z9myPXU1z3dSMSZRkYXMDdG4RY9K6I0URp0OReuISSIIogDtS87CMuG5
0tLEiVi2Z+9uSIFJXcVJUNLcqBmDXCi4VgQbO5Gs2eKPC3CVMAwBa7Sx/EchhX0bpdUXYm0HeFBq
WYTomrZavXsRbdZ0fBSaYTG7NyQWApxVx+v8hvpcB7auWvtXfuYJYNkuakyAHb7oxOy2BwrqrsCx
U4Hnq0CNhAADYLdUl5viKEL0YefmT4xfSJyBIgBXDh3WDmcvj2+pzzRu/BK+RCbP7aP741AGEbCz
58dgJL6pZmkTdOHaz933QOhShHNu34SMlCzcVZgI2eGzvl53HdijSb04Qe93zi58/vJrEgcoAHUX
Tvenv46//+3sqowmIt6PRMzsL+ietHTcmPsNwFFeFkNBTUZQvYsJqGctiFcYxPhVhhW+2hUHvZoB
qzZxq6y4Di8Hcizp/KUQVO87Fyxs2wBRjAScPfsBkWAPrcHI+SBCZsT0HlYKNhGwBkayYFwHa/jY
4xghRSmaJh2Qxdatthkeni59dYkCDUV8AWskh+IKpOAsXEa9+SIxryIW5o+CEVDHERc2GgKo2HFn
BdH8EUTQFKCBIrAx7PzAygCtDeaq5lnUFmjxmdzhwxuvDRvOYIGcVGU3IO12cd1Z6/A+go788EpS
05ixzvtq4MaHycSh2WLb4dRWtZbTqwH9VGXifVUsR0Er8EuZ9MuT/0dmNmoQpHnMUzC6ZImMLccQ
M74MQtTysbWOkfsW/Lmf+xb9qmZcDIQcaSScPaYoqPBgy73jafKdZrqFnoabWjlzorQ8OErOgiOz
x6yLRJwd6HxrC90PHSz/AZBYSVl/hXgKPQY2pfi2jxVIGE8tR+nl3iHBBdAe2Gc5nw0zK3LLIjhu
HxgBiZAhQV5ot0uGv2eMpEu2IFdFbUeAQOiO1GvhIFow0GGG/OsyDHNNtUalVPj4vYxzfaFWNG3B
t6R9SGU7mnsIrtFss86iw5l5oZP9OrKgNI69DfQ/O4JNfukELC1mCfUy3FXdE/oGIU2/6bH2Ssp7
HFB7qWwD8AFT82bFjTSMfM7AUnbLP/A+o6t7W6HlkBIWBCAE5oPVQgYwCVvn1jzgj2Wfz01RdKcl
twNDqc22gdkgy4HhcUBRuI11a+bnKxlO3mJesnaC9HKtaN2fvlgRfPw4I8XW3vkAF24BoAAnOcbm
qQY0zsNq/mBJVSpwSE3eh1rFziCNhbZLPf4zs9qBs4WEg/YHSUx6w4lEevm2m+co0J+19qgBTWI2
LDLhe+M9M9tbtb/OGt593L5NRG+VOhqnqNBjXPKRlE9FKR8j8+BPU3hb393HDareeCd6WN+PVpWh
VdzK92/VRuNtl/NQ5PsV0oRtS6hNPSjzjeVTpK/N6TL6IuaBMDDBbSZbWxRHf1deV6HC5KePJ3v3
NDn1VeZXTga2CIwkC02eADutz5Ep15rAf+pELY58LD4v2lMsAZJTHo+2cQ5SzIRjicTVFcWo+5PM
antFHhtajPq3i9mEUtP38LqzInj3WQ8uJ859HyDRyeMp6OscwH9lrdUwLhT41lalc4aWx/32/77B
eq2MR/BdDLR6hT25Reee40gGdLNhxNPixeJ/Aoazbb3vt7dt0NK6KJY+IEeG6xBQsnXHWC02PCmL
fBjgu7+FHDcFH/kk0amyB8okxu3pkQUsuqErYIq2BTd+yYvrR9P0yDnQUyIa3d6cCDK0AKNv6tuS
EasSnUdV5QAacPwvIhYRXjqXfHf7Eg/7usX+qGH74Q11dZ4BiBiM/5fQERdcWNqel7474ABuK3Ns
oAdH4S+mB5kNUZ9SSQyZ2yIj0huGtY3FT+dyVudpOGUxNAvaBC2Hxi2zegMrbb3dOihO9AoxmgdE
MeFOAeG6XH/10ms6fEEM2i533OHleWYeqLjjb9QKuE4C9M/dJnSNSC0yPBJZfLcpSQ75bVqeaOvq
tugvjSCOY8HpOECoRQGmmVePoUTov+Emx4RZYkbqDN4cs9Mdyz3AmUUEeiyE9T625YNvukh/+fxU
OU96W/gGyIAwoxd/0My6vkC8SVdKOrplaR2M0zr3hhJJZBdzTSIPKXh8cH6KP10dYkmifroBwUez
QtIbbccdpDVLna+VKHq8BZ14nEA7gYurqm8HMDy27ydDywLW3blNpvNgDc1WQCOBr17h7Vk/8wSr
sYU5K1glb5z0qhDJ/B0dnHvRAbUWgQEFAvCBanhpaKL/SzWdDsQntNjgbVCOukJRqsfANSxOViAQ
cumVq5U6meOJ5Wg+G2qF8rgmkj4ZRCZjr3pvljgQKOV98NeueAleN+Xq6dqi8cZgoj+yrdONi2zi
wr792M0lND1FYRSLG7i+u2wWwl+6zxqIQPY84xUDXLgf2lyD2DOMEwgMdBlLZedKGIg6fE6KbHMM
DZdUZu/y5IsYRxUmW5AmocJ375ZAJcKmX/ksBRdGwjKDvHsKtbIr6/FCd0+Mp9yAyrXC2cfO6epz
gwwNCUsxL1yqBM4h5lS8fccPKU+pv/PQbY7V8tTRYH38IN+fnmxbPVi/ON2P99P3Lyag4czV+3jf
8eLjTBXhhocFWxNR2WvF33GHZSG+qwhAj3ILh3PLQTs0MPl6paLCqHsGy5sGPaki4s+2iOKcXG5z
e2y3qZZYrTTka/6UWE/oSYlb6me5TiiFfbxD0Ebefm1qygHufSejw5KXxLAHj0BU4o9lWM/JHEiA
GusVo1BPFaiTh3Xn7T3CqxWlJn2dTcbsptRpVgp7IyDA5m6lZhm3+pM3BlVV5G6kZGwqQNgIfpqJ
IjL9ISnfv917ffO+lrWaX9Z1rH4gv19q/PVMQAmD47iTx7T1S9k82a/4KiG98zu14LzAotSPO7sA
UCeLhOZZagLGiUvCgnu3ubE5+xk9YzIy85SQ2IXFzfoaVvA/kFFlReGUZ1nFMMKJ4hCMZtH/L7zg
4HnpI38Rb2C94wvjMPwI4rN3cD0H6PbNqfIKXsTblmziP889mwvf5oET08wirBWlnNCx9Y564hiD
MlWpA6t5pXrHHEF4BP1B4FyoZWSKYNI+2QhmMnkHyd9BdlbdjFgPLqcnlUmBSBMqO/6bRfbk+nd1
/PUb2d/IW4+tD5tbpDpPv3G0e/9NVQNPbUc42bHyxE8DiRGxf8++TmwZg6WMQu/Yk0LPvucko7xt
6sQEGfC64E887l8oFyNhS1plPozZ6ikscht08c9xrValB+3ByKs6rCX0+2yGEhWAgpwDjtM+12AG
3UOi2xXSookPEDFq8itqVglBwo5jJV3A4PfX4yTX/fHet1jAA5i+0SWQCwnEwuQcuDSWyjPVaawF
VW2KvJ2BHigBbNm9NtW+5b5m95Rk7aSzeH/6PSpHrOFQngM2tl4QSweWFdTz74Pn9RD7oaiQAVBg
HdOBcMglyVhypuQCzZv/4vXYXprGLgkgKZT52SMP3Bm0bNkwYDySh+3LiZKK84JSLBHwNA8D7G8X
hRJIIhMvY9TXCumZWu24EJwapdzINKvb807+Mii4u26kOUetweG+9CjbWFc+hbX1oMnK/QPkmQJA
wOROgoel6FGSFCxq0pgwry3dXmp475+kILlwSqIy1TM49gQr7b8SyNrPUN/s3B7Ax/aQcooyL1R9
H1rvoKY4gzqFz4E5ISp9qroD81Xuugwub1L3HMH4Qx+HR96jwqnKNp+SGsgvZFaPuXvK0f8mwYPr
BUUer3b6ItKUtGAH2rjF1H0K3TUMd6jDWJClULzBVPcSHmWU7duHxJQE3cwDBR74Hj2nv0OrYQ+Z
mESm0ZlUBSy3BF4i4682YaQ2IZGIWtUzt9CJhAOA3Qq3g/buaiK5LU0fLdTqHUq42SXpRf6cwAY9
v/b68oGRmfv2foi54rAqwnuhWC+HSsD0PERu2d4mW6Znj0Zo2z7nRfT6Z/S9c05wdNY4iDHgXvbE
v5ZEwFT7hYhblcX6SNFz1hQhlsegQj1zF4/FnrWQ2IIcgQycZC++Tr/yHoGrKui6q2h1PCP/P7MK
7aFbw1yWTtGfuXugCkOwEPZMWvdTufMFF0RVitA4y0H7gXwvneHuM57wfBKleCCriIRgrG7PUPRk
4sQ6Mk2t1mC5B9MNsATQ/ppmjfLFxHs2W9TLyxkIvdIhTgRN2wHJvlNe/bmOf3Ysx+d7gLDi3QSw
ByfZ1x8uYR1uKwpttB/YUqgYl2BVhTJMxV5YoaHa4EBZZ1l97TISxJuKCCZp4hnZT+OTw90/gVU3
8xbJ93G2plHPR123W9Mdf5/e6yEM0dgiU2xDaPZW7DlMOm2lmovO2rJ0Gyj4iHlewOR4GvopKBVS
cF0cOEE/by1iuXS5MmlhfK7y1DF1D7NQyGY5+GMD+aKtqgt1EFJbf2T+eKuMDe7hNAHGuFvm0D9w
HKK2k7TvoRWfWp/f569gPk5vKZrHPpqSUSxehwmN6s8el1VAPiPc9+Q1/YaZ8gmx041bwDG0eS8M
cDIrJU9LEh1TEN59mQn0YX3nfHyR4/Wbzez+nuEbu+/3QiuvtnvzhCPuNqyIPYI145I+rU13EFvl
0bH5d+O928vuA5Ay0jZs/lzxOpo2XdnVX6rblctmr64cTkv6ZioCIY3WVzRN3vRDp18NjHvBpDAZ
NBhm+ya5mFVtLJ2S48phcXA1O2+NVOLzkDthzY0l4bcQ0Mj5LKIxpMmtSNpv4JpPeW0T9Ngi2hWj
ECZ1Wrx2VOXvi7uLrdyFcRwo4w4w53laTyj6Qa5GXweWkjzGEYEQ15rp4TL6RcIv9gz2/hAftJPf
jZHAoOXDbgvSKmAJErd2lRD+9e+EGwxXuyb2dS+OvkqsOiil6x+brB7SSaBuHQkJhUEdriI71PuF
SYR39YjTbNEguSbrTFvGT8h50hAq8282FmgPWF6qNEWEpLzDMhvglM5R5H4it8Q9m6zuE+cJhI6M
fpYcP0WOSYg17gLqhgwBdcSCCqNtfBzZpHm50otSmJyU+rkOkVkUXXQYJJ1qBox/v5YVAKeJD1+S
RZap6rmlYxRfENwgOl92CQ1rCt8Zp9OsVGyHXinQY4IJJWu31ePwG5F9g2bdQOMeh9z4JGQCXhIf
YLKtoUsXrPVPFOCipw2GPzQv+H+WsgcRH56Px2rO3BgYE2yaVNFfDcYtIHn6CPVXo07+qH+Rsa/L
XBRb7N1qw3crY/gGR/5ak+stqL0Q5NfcoRCGYpY1MOolYKkfmY9yCTeUJfJ4I5OrVvGCwodBgJGx
VKj6E5vxLYl5mlFfAPW1uG9uSv3B9Xti6uQ7i7jsdAHiBKvepR/kV4AO3scRNQ1eDvlOZBRfulQS
irLNTtpKd6pEMbXSrqh/2ni7fzMUg729Rjuz/FqSjrsP+JBLTeEJLHIqZ/xYEGbHWieVVu0njmzd
oR+eAMm4XauEcutPi391vApeV6z8FErFHPbjtemFh1XVfvp3jo6PrQMFiSzT3yGESHjMhDgeKUMm
d/e3nLxIEbhAph247ax1Ao4fXXwpupDTgySfFyP8QvJxlfKuofBaRO7f6D0tM4fGVsseLENOx1Tq
pgWxlJ9M4hmJZy5NqthIcCXtqUifyRJ81XI7Fh4xtXhHj2RxXiNhxFUYJpWkrA1w8nwk9b1Z2qaj
d6TalH1Ox3x23847th2PzouXuk1xUZU2jonn5bnmljYSqQHPgdn+b5g3kH5XnZaRhEFW35c2mntM
0B9cohGYcqNM/+e0RUuWPa/GY4nMuMlFP8qBYLDAHF9Mb/W0lkXVhCAxuu3e6wEi8PDcSmdRU5G/
Afm3BcVC68v+9vShqMTA+wa5DgXqzzKmwLoZR/vgaNmyMkRpRrJqOrjAOh/7SGzURW6y4FEcnFF8
A0AAt6F87EJuAygkBfhZHV3mUlWYx6zJy2fsBemXdjZtdrKlGVZuMeulD3wde1PR2BT4EEyJaSrZ
l3H8Ia3FRvAYhQ+r3a2YPySfpKvzK9NzMlt/n55BzlFmJBsZwP8IPV89ufJPjsu4lbYThi4lam0p
Mtm/XdY01ArGJMPraa5+FAuANfW8ORNEVczh2B5q+dur4ADpd/qTPWXP34p4euXez5EF+zxDJYkS
Ynv8IMEi2YYUrNhmMweaImbFVhiRAWHSA0FCJEaSGnZeSQdUud+ZG0yF+MHog/hexUt/1C/qVDrW
xqxAXpnaFyzUxFxGBGBIMQFZe+3RQzAYOO2XSulKEq36ie0z/MZPQ2VhDmPlYSIYoB6NxBEe9SPG
+jMPHXjUxxyEZYauxC2DN6in+HjobmDlQkCh1CmiR4xqtCaUD9aGtKsu9gSbUCrPLdfbzJG4Py4n
Q/WOHoqqYRFFnCPwsIWtNDsSa1Ajmn7/7xyowwja7NIdyfrPgUDbdQT4Iv663mz9P69TyKseFiAw
m+6cPi0APT3j7S0MXttvK8Nt49GuoTFP6x6D3QhH/G+jBR3skhxUiBqJRkKTAlsBta00KOVjUA1m
O3WXW9ExkI89aF9bn4xFqes/8V8k/AgmM+aDqvLg/VHd223sXtm15OSd3Uq8J/W4aNLGA8gj626y
kvCaLvDyn3GKB1SbhrqzSShXuezdQYaSpQz9oN3TTsDMekoOdWM0hdZSle2cfhVOYuZKITzZWqYb
O43npoH7fDJkpR7XP3e4Qzn51cquU5XQTp53MwtGWvg16JO/9N8QBkYewob7e+m9If9EmnS93k8F
JkqybILCl0DOhAbBVEnlPf++lxHl4DScP6Q5S85EdTkXyy6X4oIEeKWxLwId55qDIUBYr5Mpfk/z
YWMISoPwvac0xJMCr8LSI/2o/u+cDRloXmo6eVu7SDInMBopNSgENrVroEQ+FSXWH3ETEJ27kXLo
/cV7Ml1w55MK4YgygM2IYLzhoqmi2t85grs9tQituhClLXiex+rXTSrptHqSTGq09NCQLA2B6D3n
iQZNuVe5toYvqfWUFjIc7K8gjEG3OjYrz57Bo5m9DX5dfFZrm118Id2Qmjb6VfuEqo5tkIx7BZBM
+kphLFth3voBsxA8mZkopXTLo4U6Qck1JrlQN+qmamyW4Gg2jHWIyBr20vpwKTJlGArIOZA3Ftnz
0hxQFvldccQYBEDms7fThXHNNlgU4MG0YJPMal740xoOszvG2Oq0Uyo/XYIs8vwdaXhdBLl/XNeu
0O27W8E1oFelFiCOfU/fV3+nG2vytdClR4TBmjVGzZETa1cHPaqqIjo6QEbdSdRTPdnvemCMjv00
IfizTZmNsF1dTqeJ96dhWUfcQdbVQ3/bIxDJbXoSV8QabVLvY17zHLkAPmDlWiSqh3Kwt8G2YvOb
FR5f50SzW+EW5fxfg3KC8BsW55qEbLLYkSHfMtDnWGfXFgpw32+QSvB2dRpH8Ckn+ux2v6k6/ABp
9r0jQJcUYJqvIAlyF8j7ixEyyKOX0F2VM2bGegmx6BapCy41sd4fHqKXFlI6ykwtlhbine0LjB/5
VgKtc2NAuuGP7cJ4pKqgDtb3N+wnm9NQkqRMslTv59SpyjOo8t/DV4etJh1lNRm1+eka74Agd49z
vSkvzcGME8PgfWT7GT4tcCcH1/b6OqQRxSz81a6yIshdSs8Xdsds1N3JBS80pIpL+lK9TxeqAMNT
Rf1J3bVmXguAh342Gw++ZPLjOja16Eqv2jbOPf2VHt4kWJWPlcgHGdRvCWGg4GHbsPb7+OGIF4sB
DqJ38X7/11Jv3k5FCrMdwri7sicVclD/4qDwDF5ZdUOS9jrJYBMYtGvxiI9WyuH4ikcqw2t0Ucss
VeAiBhIw00VcVMavKtDXKaalOGIOdUPxS/715Qmx+ScFhkog1eYBG/cPEVZEpnX6akIO7K/njL73
ZNRlrW4V2vlQXmveKeCWRYsKlu+2MKAf7JLd71JHMyapZBaOURCJxyU83kE9HfuK4eSWT43e2KPD
6lUd20Mf5Nk9ygTV5Jd8yMjsUhHK2a8NPDE0T444iz29a4ABdv0nlbwjyijr35qNqdhsQUndl3rU
SVh39g+ev5g1eHFB26KpMYYWXgIxuA0HWmdvt0VF4tGPdEUrMEA+Ti/Zw1LF7RhPVd9qiUMUhEKb
Yac+K22cAB7etXY0wOTONUvtmf4oP9sD9V4IJ7S1WV9h0ZwG/iU2Kr2TO9I0Xx/out9o+Va5h0pc
SKtxGEJib5YW5H9Fql1p2kZIKmPWXhtAdrUskGjyg3b5AaoAEaEUERqcuq8y3lRabsExcS0RmR79
MCkkvxVGlGjo+h/LIT6oePgktuTVvIJITCmfzBJte7IY0gQ2oYteDXhAAbwNtlByGpmtFdMz8TpB
v1BAIUaBGTnJ2jE/yGiuDtEPtd46mDFw0p4EypqXOX4k7W+L8KZ1jQSoQuQacFtRYJ78oxmxv53m
yvKDW6qAcbnuelR9kqC9SWTkQP9vcxeXEd9Hm7zkc4kktZsvkClT9IObeK+39PzN6ZeTFyaEyiAf
pusyIlNG0Rt+kJx2Q2YnEDrHwZxRcYY9hlCFN0bKU8JoaItabECgN0kkiK+WGiFg7ZB6I/L2HFrf
3u3VfmAvcpZn0ZOXWBMk6SX9SQUVsmJIiqvTr7SGUrofhTqW9yI85FsKVGxCyD7KXNufmrhLlJn+
m+0Za4ahLvG4uejj/rwZYLu69KL0VnxqM2OMwnUIByS1WbC+ql+0cv/q4hP3GqRpzT8iA822QxOF
WMylJD3Aa0rqXohQB3/25nY9R6xz8qNdqz+GZh5i+LdZcsHlh1s8UUBYSKtpt/lcYX55CEygkhxa
8CO5v/k5hUqZnrcig3ZjS+o6SqCXG77cKMvnTI3vU+b+emyCAiftz9yXDUm1ZlO+0w1LV+x8mKA8
JtJ4efjPnlpY0t37KnV3ARanj8ExbyF/gQMcsOwbvu3GmWIKJYEEklLEY4P+bMwC5VJLRmIv6qkq
vfZ47M1yTiCsarpuKq23V5aWQ5iEKlWq6glj2vbfUynNIVLAdTADNTb8nCN2ZtJbjKoy4EBO755J
f3h2oMHHn1ekuiPDELaeNj9zzXPX0KkpHDCGUAWEuTmGrmB7nwBz3DOAfloeAcT2YuXxugzKRj30
XJCkzu+m9/QVX+ntAQ7xaJvnrTQu+4fiElqyRMHQ+qqG/4o4bcaWdX2VxFcZ2noxv0758IQzWTGo
bSEls91wOhR+FXJhQwSpKOZXoGt3vcKDSLgJUHIBXNxWzgCH/UsYbJiO76uZsWAjYEGaTDyxURY8
3BDRLfd/ZF0B9Ca5Yxo6hkcFWjQXjgx/TDgzjKleVsLXnw3qG4RQcKo2YEHtreO7FBoBZNZ/gJIb
BQGtqKN9uN2RSALlA/TE6XdX7ce3ctyWS23ptNfUuesqtkRaaWgPlZXnDO0K3JDAY9J6HxLj5QvK
7iLcoe5qJj67fN+lVGx0OxVAiSXoFvGmMqxulEpcmrbgLTFx0j8XYrbk+jkxPc53I+jXKS98n9Iv
oSLZ4SKRFenmWpIHnH6qNqRdKYe8wjk3tEsSCmVudnB7hFtiXwyBe+yW/6M3X/DeLyxE7hZ6EAVY
WHoZi+g47atvYA97Rr4LtaUvwbJlHV45V6WjC8MXiPJpgcD8F4w5GtLPBYEDdrQN18s5WHtIM9Ft
aKFJNW0feVHvoG5t1GXunr3f6EhM/bj3G4Xis8lc/I/mmT2czfC5Q6Z5j1NsbPkZChnHlVKsAtgl
Rs3LK950LIpQcAAf14mwH6G4IEWzXpw5SkW8zS2lQoD0zxpaWlvOi3vZwfXmddlijbTJq+mEHPRB
vp2jbgeEn30KV/TNUxv9JfB93+u/nrRCUW6i10PjjHM3nw7gIfiR8jAKjSftt/1crlF2QL+VRJJo
X0B4xo/+v7kaPIPLPT88uBWBn0azOBPc4Qk4mjdJuPheBpAyqAU4qKXmMF1JqNJ7FdEiY7oWl/HO
UoGI9XGSPA/WWK0XAVmPdjxYjf6Q365YIBuN50/VeWwxsyEOz/y4eKgMlNGtxXVm2qfsnRNs51Kc
EEisSb0xEl/sFsPw/loEl/GP7OypjZwxuQ8FDtnlnzuNqBS2go+wSl77GKeb6mfezUjt2owZc7AV
H+ykLJ2/WSmdQ6ibb+laXXpaT1xAgG7RnSB12LeKao4ZeZKEY2bN+fAN0UKqozSpAVuLahqoHfxT
uH4s0bymCyvjhwuVfGQDE0lunAWNqrwQEzNOLL0N64qn6Htz9Nr5aomzO6WSRAQ9bZDCfCcnuHI7
NVHrpdcl75YTqb/F8Q5/e6Jb+2uBx6+Mj9W7dvx2fHWdC6WSPTKFDtQ+Qe+fucrQm53dunoNi5VI
cmsGCI3vDqSiSdZAUYIeSwvzcj8fNHIMYQh2Ur0s2Y/Zx7tpaVZrCQAD0W04wgtJo0V3A2JvlGxn
N6dOsk/lw8cRDqvwk2kkKHegcG+nB/w355y98yNYrQvhUf2ZfiDeNA8Qt91QvtO5v+1aTXL3Othm
uJ594FlytBwcMM58WxQnSM8qQ6aztA9/JxgGDhG9gIpZ4Njo+/LnDV2r2pRq93WXYtc8APytOZNN
hQ4BPbnYPBk84oBTb+BtvolEq6jbnDD4USHCh1GkLBLfdOkuB4dVTp8xvirOoRfHbBOXtykANh+L
0DSwynDqSN8PB9fI9m0F2zLPuLVKcwS+vAqGVN/zob4Tz0UtQ6jZeeE3uo3CnnlAeELqIrneaG7c
Rpc/bbRoNu2INqMMcKfa8zoYf5TUVoSRlwO66UReZkzyGVkz55TbW3pbbLpcjZArTcr34JX81nux
SimlgZeSWJ8Z/nDarBeS3+xem5Ti78fKpkKiVSXeA97XbrJ6IfNMHF/7Zirbl/5xchmm9asl3L9k
5umpI6eoSpcqQ5LlhRe0OvCCrQuY0ludZXw0gX4fZxqavP+rmI59rtCQftmPJiWGGW1o/ehasbpT
s1UviYXKUaXXIGkII5v71uwhQ87HNReE2EZase2czD0SLrsOQu6MsO0IXzwOcs5rJCG/Ha64B+nA
OUlE/WFmjjekZc82AzOD0hGHIaXhArAC50OKqHQQNdcSE1FOjlY8jfeMveAfNeU+wjhrnBc7tF46
M2mZiYB6g+fEETcDLCN1aJt+ZgnxZmsac7bIygsH7oiihcv/ns3ubXgniqKnYbdymv9uhPNJ6AHb
SO8oBTwjdJJcK7QenUc3Ip/VXVVf1QT0FESHQWFmoSO51LsktuFy+LMzSf1BLPMdvCYofPOjGUnR
in35OgSeWs9/ZKUseJxuOSQ0d6ygI2aoCHbaiVDmy7h/RJ0tg5oR3+ec0dFU79pTXSFHUGGpM67s
PDwMIK1K/Fd34B1Fg18zFOJU8ZFH9N9jMzY2Brj7Ssoj57E0l6iOQpD2bKxawwpTYGBj4/WwS0Q5
AxLYBMSACnEnBcV0X9diwwbQC1H/t6u/qzz2fy4hsEf2X/2hO8JEAYAave+wwSua8bqlYv37Is7a
ESizbyN6GVURGRT4jBfTNHDGBXxSvNq1vYGUdhnxPijvVwxs+22C9hZzfNBQ/1SZREONLXBt8BXJ
CChO33u67RxIzmwrx1vSTNcRShSFNfiHNqEnTbCVYAuMxEvHEgw+JUwMN2qoYX/Nw5WEt96hBt3p
z6TYnxgI6xB707Xmmm8mGIoKS8ixWJ4MDwD/j2YOkcHqQB0DvTNY3L3buhyfTlpbo4+ofwo1yuk3
HjeR42zrDTBjMJ4kQctV1XO9Oh3OtBANOeQBrJ696rXN21W7FKjsiHXYZlm02LzMHLCjB0YJESNf
WoDVHgii659oFKWcM8v7VM9T1XDTwIFHUiTQP1EQYreQZZ4fSYjcpR9/L0dlxVieyeKLtVpCaFI/
U/jL3pz9MgoYWpV9TuY2EoIrA/CfUN1Bx2wKv5BBeqhVXkKTnJG/P/cjjDXGYUKzJJ1X6d5X6CSb
LhAGGm9gzNMtaNnROw/TjlFPhnMOg3rTHc+cxohOXVgqAAfcpZ+STxkhXqGWitAAXz5sLqAWJ9RG
jffOewehdW8Elv2pXAdRnzVUDrysoCysrj6CvrUTVPxAvnRUZ16jh/xedx2WsFYSXWo4EYjZX87Z
etmUh9sDGoV3P3B1DYpGyZBPdj7MBuMrdATRpr7YGC4KFW+8EyzAwrY9c7cXAhLy8NHqbtK3hbrZ
e3GY9jSv9FavBs9DrfPumUHD/ut6UBGo75DNFK+/v+8pFL4SbB6YSLH+ZDiHP28H23NNu40iGKsP
eWdBQQQsA4GwBFMOqeC+HtgM7M+5RdPcSmTSebvZ2aIn8ucvFwBN7e0CRXbKZSjWa0wJQ5nLQubl
sPXyaQzfFciw1p6jgmNAwHJ8oQFH5//LI2BHCtuwtMaJnBwtkIwPJX3PrNn5LPAeB79GTviwnudr
Ww8GTqLsZvnz5PlmXu+Uxv0K6IVGE6UlkeAp6fqkNpp94vEbxdatyMya6FizRsEwtNN/qCCoUS3P
TrkiiDSdgys1jVcBTBza3bv6lzA70+2zAxJUiT0weRdfFWk4K5W0NpiTih6XaMroeirfhmsZ0Db5
aM4UjVp7gnH1Bveh/tisAD4555Veqjiwf+wBTHu1TRjFMmnwabpmnyLp89uK6EoP1M5s6/u11ZTt
cc2Nv/YcvJH5/UsmAiUePYAyXeugq166MvliIpzoqVaBqxXoDiWH+2GrsMVMnXjOEtctSdpfTJVb
qS/vEXLOXIBEKWgZW2Tqv29G7M9a21NpQ5qfs3MLore22OzU40hnS2Qa8+c4uBdQxqJeJ4LbPjc7
HFoN6Jyr/7+itu38N7/I9CImadNEBQ6QdsbvZjKrEFt00KSYL/awXASYUgYrQWD9z2VDWsdmqFZb
m459rrK5OzF5bs5NqpZhGk3RrwbEum5kubzyvGmag8deT86tphBWTfFkKdCaTJWlCFzGwTgJNqPh
hxfx8rFcImzDJ4a/Jj/1cXnt9daMMj5jcS88OQF5rgBTZUBXyVBg4d7szfNhHN/xGya6ia7Y3Lt6
JZOtwXjI3ilVRmePOTgoBLM4usz+qydgxD9n75godwAXdT1gQbmFtYFE+FEv7GLG02Z8xsrHtMOs
2TApyRi4jeDbSp/HH0xkaiO904bTbdiax0SzuLTkM8KzRSd7KiSoA8ECc9Yw+S1PoIUjOAvYlNhl
DHb9vY/0UQYEGpOqYYGh0hHlj1tlm7dVroORlYtd8pkkFNTQ0lg8EROHmb96lQZCkpV1453wT/ZE
VQW5JSV2+AEMC+UK0CWBzeVp5LBaFyCQeXz2Sy+yaqGI/kBTY+w9+i8nczLN8F40NgditA5fh/S3
g/g0Tk3qQfuD0iCd2My9Y/yRYqIWXepHzFFOktYrkdkfXQ9CIgJ+uE38MBKEzPk7EN8S88/+og3k
9i8Fw9y6HHqnynLaOrsgR9HMq6VtIPx8UPMx1/fGd+X1WbQkJt+fWSgrexcW7AJdv54xgrgiAo0b
GKRbSi2hPUkA5U7YqTcIwEbP1T/4JWhxRf4vjO/qjxJc/MA+/EBOy/7MfYIECgOF6YAPzZrp3tI0
MNj6i6jGH3f/D9SfxpgdQZXKtN2ENggI7VuE0kDzFLIgg6bWmkfPyqtTG4NWk3M/hCWYHtJoyWvA
nToLSQPpJqr7/dlvVLgSnkrz82o3KVKiBZPmrow5vFQSFRC4TcglB8i8TEFk/8AYqHTFJHazoEIO
QLhi0/Bj2UZrYfkhMp73iyLtQUzPUJK6EknWVOeNAo71XEnkHzi9ZFevwP0d5LoLDTJsZqVEtsKL
DKkt8wgJcBZUsjjz5/0qVmfaWcPA53gwHot0+XZREHITKjdhyZ2Y3gImc8hAfNBDAQEISa6bTt6p
ywv/tRn8VmHQYviYoQHrN7SYyOqJLTMSvUMxXnk/TmhdNNSRZFN/x178R3yc6dZ0wfgrP2D7nHCe
EtOxkyVAPFt3HDX6ysUsCP8QdnWqZsWGpz43g7jserHRFJVFkwayhEhUOMol7DlcnPIL7Qn0LCCb
9awwfCwWfVaxf23U/SD5ZjF5dvEErXO7anCWyPJafuYXC1/uRmipz+Ypp/D5Q12m5YdjqJxWWL9i
rN1cIkxv55i6oo+KrZL+v/v40qbQIrmq4iPSZDNVOe8E9cvWp5fKXlro6rUtJlw4ANkpPOROUQmc
7SK1L3rv49s2r8YNNOhPp/47cV8k+mSUkxPXLBpuH2fjFOSAsfoqhhkqFfBGtiwO+glrGa7O02lc
SYqvYYVtuoyTgxDN0ApH4VHqpwwHEzPXK/Fxu6MmRoOb8UwLTU8AcbCKNZOpJcK3NROOlKs9i/0D
jRPLn6/yzbB5lCFGnpdF4+iHthP0+X2+yg71NKe9fBOmKXeX+C23vVCQgorfQChunWjYseC0ItZN
UofHLtIifHsDFf1UHhvCOMWTNDQyB6451yoNiFwrUTFx++/1QFxA3E/MsBsbyMA3uFhYvbF9zGiz
e6KTC8qdn3tCISmdQb90TH7+OprntXz2zdmu6taGwa1hdj2cKLCw8oVtfBSu5CaJhXRC34MwLbFJ
HDNjoj2mVsvI1lpx7Nu+qDfEx1Q6GAcjHbgQTu9Ni1PVkRZu//cM5b6JD797Tlg3s8nljwTlMj7Y
pHhiYb6XpfEBpDUxzaxiX+01PL3AzCRI3cpF2nH0+nuk3r6/1mvSxEtlFz26pdja5RxdDFHvJsgH
8DyPjsCY/opYvakEbiRVxd06hj+gSP75PHs9ArwTvITB+ZlZnc9g+nOPDVO/rqLjZ8C9lCuwvhiu
67/ugEFxDwqf+uqwPK1GLjrfrzwWcO9RFveQ0OmEZRpBpE5musFlrrBdSyR+PdQkXZ+dkavXD57y
NMS060IR/ml8FORN5kiDltBHU8xXpKKah3EKf1pzQpGcg8wCuUOx9BFqMVu1YpuzH4BXBye2sfDI
kocMzr6lccyomjYYKNo8hAPr6eVy6GFtqBn18hZg7jmDqCfuvQhPnr8jBdqPFFNPr4JhfcbgXlEq
+R8ix1KOALcJJUipoqjdFF+J5J9O0c9ezA5iVmUyQTUQ2IGa6zmnlS9rVDX3kXuOoM1AIZ6djqfF
qvMHB2TTmvBvxGdtzSG/Ukraj/HKDOsrY5+H4h5Vy0Se0VXelyQCwg3KXYvdxaHLuMppZn2Fuqo5
Rd3QOqaTtkZFDGuRhXzlBa73LDhfcDrkPFaPJz1GcZ/9EtmoHLsJ/Mjc0ff7mAEtJ/nPi9H3T9rq
3YJs6i6ZcgymEKpqMcN1JAicoiF+mWrWU7nXv10UoCihN/dYiUocxBVFuoMdlVhiJhnL+aYigiOL
tKXTa6lhvw+KFMbAmAs9xgPFATgUMw4TdiX0ZlemqaAPIvKALSQgLac8Swkd0aehnZXkRNycmmlH
amOnG8ULtpZ1q/uaHWpRYNjeaIVKsJcnCxBnw9I/Rllgky3lu1rSoUbQFI8wxh4LeMyF4XsQdDbZ
qlIJqhq1eyE6q62F7fJJKbu8871bvwMZ7qK7wLPJkNXg+VRcIPNYDrV/JMf0EeVIx75py7DMaa+I
hFcEjv/JgfXtP1b2b2etm0eDNefKDMN6h9vwK9YroqQD73qvYwAOiqH8+v9R3xoieH4d1srx+SwD
7nE+lD11SX8HdZVH0Bp86wiPk48yPZATJh6yBkddWXbUglgQenlYVk2Xd92QGNACynbgkkdsRPFf
wdRjtUGnSCFSkKCqmsJRN1dV9AQ+1ugv6hwzz245VzwMX/SQeSvzo/nro5gAIElbl/sRyVyqlYZG
PfpJodPciAtmvU3SnsuNj70Z6sQNj7vBghIaOWChlHcs+RVoj/55KSJn30hHCghxp7Yen3z05lPq
6sTgm9L6MYb9WvTd2G78SEJbP18FpYwYyR3zbe/ZGGBk8VR1RZeiy0hOM5xggSRSxyABwd7gXQKu
97CUs3C4Gy9g35eoFVZ1NvccOHlyROU+EZoIbB1cIYx8mdCGMOF8hQqkh220r8G14Rqh0W4cNgCO
mW7xLLVJPwmbY7m4fDnr7gaFTjFdBVXxykl9yEtJkBvMoiUiFAMocV9hoO5C0z9Emp2GN2Eg39mG
Se6F20GM/Vm7LVIZJ1m6gTxsxuShaEy9nLEL2RZRoAxv3xhtGW3s+YUUjPef66OaJKEejBtgJmyH
QH13DbKB5ysBwdQspaSyZ0/pmFi+8Sxq2IaRi6BeDzXjBlLD3cJD8xBPWU6eAXSadPThEb4HA+ej
Gmy829FLGTXEfzv29u92MN2UYroXqaz8xnlSy0H2tFuOFUTRSqptJsxfkvrtsVUhiq0mLkKDPHl2
DOMbYmBjfr21v/i1jfs5YABNlt3dD/pcWyWwCNY8KtfDfTsFHaVDLFiufv4Y0uqoDc+e5ItZGy2O
buiqGLSM/MXvnSHIFMmuySrHGaUl/S/MucH9JC6SA3IajUH2eeq++7N4/KhuiG66vCUkodjzUebV
1N6fqkqC0WK2aeGPjhI0bXPJsPSPVDa7JXq/DV8UzPzG1VJaQKkL2EBZF2si35D//Vzyrmh3KJwg
GUdabmOYs9fy/m57WvbX5sU7jX0Vw7gq6tZP4T3hh7Mer2JOLgZQmlXxY5ZjD7RuWNMKLrGfO6az
zzOW2PN1wpsLIlN+q18cEnLtbI+KySbqmWwjjyL9klRjLhFWB2GOvbxXVk+M35K/51TUpTyblgzf
nB/fuZm+gMFB+AlreXlgPZMB4mksZ8LSU5cyE4eWRuzzRcMjs+HtAD+ayX7HZERlpxmTBD2HOumD
qPnzpsiSoUu+ORhfbsuzjSydOx3SrZabadrNiPBCYzjZpIh2O6ItHtLn5oBKL4e/tL8FAGPJZki6
wRw+FDIki3D9TiBXAZrgT85o7jmNnYMLAnyDEfYOdw8JZsKPvITwEZVEuNcs0XrmCBdje3YblNzA
hhvmxmdOudUM9H4fPN3SrE9KQ8vsBay25wJsqlVtibt7EYQfBvMVJqYdljsWJTkf/0XprsHmP4tb
LZ+02YzVUSRmzMdXI7S3uOsAakS1pf3wDKNnhGDDn5/cZwp3tfwpqYDQwwK12gkJeyL9LpYX5Q0g
t/mDSoRPOsusJmwXUajhiHpBKj6UzR3GTnPfhRp9jYpkJCrAA7IrOExqeEsu483ot2ptZhAJrkk/
qnBS9KFAJ3t8d6mhZNXXtmUf0b5trJc37laCBz8K7KrQ31M0Na1OQOVQZ6T1gqy9pLa9gtVLUhPE
TUEsUlzP3EaQnJF+FS5zoVYVJ1sDYsEBixv8aRZm1j/I4KbKHf7pEOLEoCCouj50Kn7c/s5USzWI
Sx51epL2yUDuo4RqH45183K/2EP8hRZoqbrIOvrt7uupib6iDh0cE6nOQkenWUEKZG3BaWmrL4UF
N3/Va8rpiRT0G0Zm1CsmqveYnMyayIo9UY9RtxFvkhnNTgU94xFzVw5qa4jJkU2Ks4v4jJZyFMil
+D8Bl7P8TnENgId0JAan82xtnRMPNzMBx+rry7fHZjuh4WcyKQ7ZS6RgMPwL5RMiUid5+y46CcqP
oCzzhnQu8KILBQQxk3dIm4QymT6IGzHu+OtdpyAptKIdaFFV+yy/5a6MOdXXN+3GlmXq9Lqt+ZvQ
CDy5yq14sAQAw2b16ZtyINehKVsv6QpDdBNNGTNoiFO5yaxb0iZtiFtTAPwvaAemUP6wXDKm1kjy
Jqap49Ws2SFOBtEpTme38Nilma6RiXch2ctulg9uB4m3HVzH3tfm4wxBLZPMVWayQ+caMTvAN/XX
qiZL+JQQjFFWwJ0JtgF42RWuOjFaC90ILV7DLzQmD+RWy6ySEvID4BSA1Mag0lz2HeI00f6cHCM+
ppPQvd6XrnORNiUZFHcj6SRBWG2Dn4tvUSN4z0M/09MYVPlBlMswIVJoOieA65tK/zMuq4yR9SAS
H7vEy58OQiDUgZzb4UMj0SM6CsEhXEgZFY/mVzpcl5/HK62sGXSCrIlpaKn/GUcQspbYzMRjSMHl
to6JTxbYpFEHRpcl4J47S/Yj+qthry7Pn4YFOqCURcCa4p1XUJsLxGEAtPCWlfWMWWcQgqGvRlTd
fQy+Br2zs17dsEz+aa7Oxj31gR58VwFDfX7ya3JXL6uABiEZrBRbsDscOT+RNUBnK2FhhX6OVHXa
F4e9SU3s4cI42l0IvWJ9HMNfGixSe0msmOPRNW3caHEGwz2QV2Qqp2jEcVW86HDJMe210W4DjlER
x+q1MbeeaTmjH7knwnl+tACAxNMeM0AOzG6gpxWDjXKr4B3vllSwdn4XsZ1z00qEe3lj1U+cbrVH
otZFOR3ZjG0gc6299cS1dfEpmLuivdM2ok9AhfS4vomYiI+0poKXGDAnlG7mORSO80cbqT4j8e2G
wT6ZfHSDsCBFkj8T/wFhR2mMYkF+tas5WstSko8j1xl8MEnr9S+7p0tvt8DTxUhNwZlyMv4LAA+g
6pUdN6uJOyUYk7thZExBPqeWxrSqGD70datQlkd4L0nhvrt9KOWORJ1ynnib3iPQAbT/cwjuKxJL
bPqAUMgRO4/o86fpuYiyQ9p60cC2HZ1Jy+4g3gQzzKbBXKdsRfuO9TgwmciCNofOMG+ruuVT2Cgy
Glw1FcKIy0GV6vdsxmX3y72z/JaMZJMyjfpAy0m5x2u4QvoBMBqJzHzY6v2R7dKI1lxl9/GIxwXx
kUmj3trvVzq6qTFJZMEXuqSp/s66vKLOgEpcYNrV/AKwAlFtKPQ6zaqnWSiVdi0/4L2QpPxdvz9w
z8KJnU6S8NfIuoHVkNkw+DRBbFvYfb931OqN3J8vBXM9djvN3MAYqF8DDf8skoz+57lROcMZDGvZ
IzPKDLPi4jgY9KrDc0RR0goZEqwwOjgRtwSNPePxM4ieM1CSOCtbaoXzKy1VJBzFkgvRAG3pMaoH
hihkszUPe7Dws/wtJnCSO86kcLLGV3ttubQf6bxmCdV5GBpbSYUvkUJXh9lEwSO0h9W4rtd0DDkL
udf6Q1t3Jja06OPZfx06TUsxeVFoMoPAOnXFZpOpW4XnXqMfwpPoFIVNhs7coos1PuPc+dSZWqod
oSauPtDFXPcgnLKW/FywXtkjQJ6NUE0Llt1qPb3soxx3PSlUrmcyWV+Lu7B6q8ms0KoP0ry//J++
6Eu+tesrsW9DV+4DBMEqmceynSjqH0kZsClOZxAQNMEuCP4U7DcJeZqvByUwQgKRUy+9mjOv/kPn
mFnoJRcAXWdLk8C2GLYsJbbS6ensbmsyILhcJ6T8AHscQaBt5ONIV3RctVETBJ83MWTdoMQMVQC5
PAcOW5l8zS/IreniapGl1oy0fMZ5b3fkMVVi09lCMvDLE/v0VaOZa5F3bo4mH30PJ/fjORzK0xGZ
7gK0nGG0xckinch9WVoqKXr3ikxjYLfq1d1aVLRsscTiChSYo+Xl6TxB1T7gBwZ8Md6aa8YIOx7a
r+wgX2p+GkakFPA+3VpbCLg+XeTvN6xNXHrkRkapZh5IWoYSDiaEmk+M5F5tGk+9P4/XD6SSud6n
5odlPAKFcAH/1WcwuGMsCbfKbPvOim1W4h24TKV8e1jk8ysZjhnNFidafNiRg+FCPWuq9mhfV1Nb
akw/2sQZ8bjNgdZmF68US85fcH+uCyrYsxrVzyVkhlV1kPJImk2LXMy0iMUvy/NTRFaxGIVdSd63
MRmUNtrQsgnrX5cmejcvpL3DRPlWedV3Fazw1pU9vlp50NafaaeNNHah+SaCuhOW5K0zW6QAEeYO
RLQa+YzVWNR8U7giWvpu+91mcUc3nKQpThgwP5y776bAWStFUdUb1TtkKdKd5S0cJ8G6OkTI+9KG
7NG8DUNLpjBX6APOo+t0pZbuo3/fGIuZDxXqPudxb7ImEACO3Z4USHV+FjP6TWdqOZgiGKymRxkm
eKXw6E5HX/KJzSroTpsElnUZ/ay9R2TNCAt4amHADMsKeEr7cV8h39otFI/HqbmZxcmN6XF170Hl
5T7Tx9+OE72nGeuRsBe2hvvOgRfR0OJNZzV9DQGhmHgq8Q691whH592bW/Ij1FAe0lKighpB99rt
GSYguTAfOTk8lUO0rYTUSyn/RUVDbe4V6FYhQyHzrO09A2jfelEMwNHntNbus90Bura+qZbuF708
NdWdwglp5yfVotOw4d4d+HiPc2g4bJPIkEWCmoNGRACPEb3xWpY/cWumwqAluCujJjUzV7RWI/BA
9p/m6dSRf3ciJoXQ207a2ThKMT3MJzycl3j7gWE971ootvtsVRjXlGJzgf1piMjHhM8s9Yr7mLFl
lSrscEwOqENdbCQNxlGI+S7BJM9n75QgsTw31dTql88xynLPZ7xRWkGZuErQ3wBoR7cbQtePQfg4
Qf+X1Z3susV9/YAkkSXjPzc+TK0H80wtfWA0NQuMllo4G+iNWR1MnS+vuL2wegbRXYrv/l5LOOHB
6oJNZiOyFKDpP6wS817CxgCydV7cguLHFUgFPTdMScerZqzEnhB0HopBswV7k7wCOb6pFOlSvP5Q
SO0gtgsi6JrNEc+4z1O/Yw/3PB8Qn+zBxGxnfdx9h9Fri4T2/Uyef0tM46I31+WdfgOqSpy7RE7L
YF+cjry6XAuj4oGrwkflevonPxEEU8nSgV1R9CHTIr5QnZFU6D2kZcd11H8BAb5I4FHB3PYsA7v7
AoTbSpjTPBiKYJadALHzoNP0k0vMbEKmxMNn9B6y5WGhPc5ep5HLH4+sB7ZCAWjjlNZSciIhinbF
7YGZMb35GZU4QcmuaVpyzQHz3HY/W57VOEeKctgDOOlmFWPnPhivFbvTQfxlBtSuJOCOAxbFZjX+
aOUImlxhNXo2/NK26mnsjHctoJHBiHzZdSTneTvzlqVHkNPGOD4mWPc9cF642x8Y3QpMY4kgb4KM
aMHBXETHpO8DeWnPEBeJTSTXzvslQU8nlCV5JwCtcEJWpdNR2C025J9Akr8TBYGqSCGTeaUzuxaq
iI0Eq6HbqvH6DpgIXf44TIMqfLcIxX06+raZgMUlGwfV/53wDzVL587zefOKMs+ip3bNEioFsXgX
LxAqI8l9iGVVA12AN2YkL7uMUsrjD9OszEYZqU8U9lhhxbznJCE95B0K+LnldJPwLIxyzyjka3qa
bhorowIz+kKj2b11xPtpRR9sfrFEQB6YEhFh2/2VWJtFilXq04lHVOKqkWdJJIuQXCDEgrc8cATU
r5HxmVIjw4do08nKQ6fjjHs9RWp5uK0eb+zIS4GBwfQWT/J47qlxXX9VTapWTZreJW/Y2yn9WNvU
ZyAzeYFQ6wYZpCQ2mYpmCRiAkuWyh1LOwjzKqXSfPxyQxcWZK8ntXRLJBJQ3GumXNdVNje4ExvoD
rPGKqjTkoh0hGAjECMkrZkfZEb0e5TjYUdsuT3H/I1DdkwW5smPqdA9Z2UeDMnYaibCM0qscEdGN
o0NJUmmWaXla/0V+ssucVBpIVqO0YRuBk1Jox1DObYNQH8+hbfBaCaA87ldmYJyear0gks1DSqGx
eSZdB/HF3ydkavJNxEi9At7xKQMkCF6DYHbW6dxFvzykG95ngmFelI7cQ+3Tq0a4haZrGTfv/wqU
PRwi7aLefTaoreUzeZtReXN/+riDfJo+Ah6jp40JGPeovBGaIlqMkQ5EZ2uO4OQjMYFSaCDqx56w
hMJpdhIBkaggNhtoOxHs/9DERenvG9SZQhTialUQJeZRWZbQ34UbsWsk9Wi1lMVU9h74RVbd9Mz9
THzW5Vs0vuoYYwbzLYLSm558olc4rKmPVqVY3ZkM/sEXCRevb+F8BMSx9V3cu9N/+RckL3cZR2UV
KJR82vxD/fFj1Of88npVnutAVvt+TUB4hPkDPKZ5wb0l4GoVft82wrG6hjEBslYyOj7m2IcSXfKK
7Ocidv+RruueDoDjvm9bINx3znJ5BaeXnLNCyd2Fl9Ui2X8DDlKKXzDW92/hHFClBQqtHubuVnh+
5s2OA+P7SdwtSV4rgs9J84l41ocxj0QAk0jvKwMiCUWQ/SqQ+SsoG7L5pSpAubMAHHsCR/32XmkK
/s33A2ygbr/hS+uBm6al/oHFPkCgqLIlnT116W97EC3kJHaVYS6yeraI9iNFG3g7yOCNpWjaIyQL
HIOCNm0Y5WM2jyJ2ZmWV7c0jGfaw80McZgaRCTVlYzqj0THDQ5l0vFxCIExuvH3eJnEREluEFQ0I
9Yh++sm3rWSed/gYQ84WrpX+fMLhOPLDXmq9ShjULMDreJF9Uh6pXbDzoUQXq4bc5Ct8lDYroKBx
AX79nLbmM2LG2D0jy+KgISMl2E3z1pCaiTr1/9JE5JZb6m22tLz9i/InW2tlFF4CBmpmnv8SdYmr
DJMr2oIbxWQ3PmhXknwjsJOYP685LGozJ1L38ugMIyFZWxxLLzs87Z9atzg6E/ipIDbx37CvTIkZ
ycpAQNlTxO7x3Ve+ZbGzk45/RF4MWmXIoNA6maF6b4/ts7bMP3NmKnqI7uY77pYRqCxXy/4CACXs
LGRc+r/JJ+C0lnWUJzs9AYb/o4h5/No+3BeClJX72THvaj/FvUzXKLq7VJc5v/E2B0AB06/TLQIe
EJz156jQukM9+44ebsxx5mQyL6eanxsoNjUoLxcF6z8ZdTHjUFVQ+buCDlHfFvj++wElbYrkb4IO
4WQQuhuGJPQLPA90uA0ufT3lSAYJz9x+y07e1U0PA90HipOX2KagMYtPR9EarGzpblEznXKS11Qq
yyG8PLf4EMrb2dsKhK1id0eXIYHi/EPh1NxFQc9dbhohTa74yzB18pGyyja/mMbV4lVCOLPVgmcB
IBCAk/zmSnZOY5t4CHp9bTu5w0DEOUZg5ZoqamNV32HI7dkvZTM7Ily1Q10oFKkXD22f0HlxurUD
GZle+rKmdVoJ0Iw+wZgUUsUb9tgYEtgxQNIv1XpKICV4ERPDABuPy64TMdHaWCRviDz091IhIl7J
Q0W0DSge5O2K086ZxncwOyuauPvhRv/EmEM5Ic1UHcELXjIRJ8uDc+XPSiWt9HP7KwCcK+zYTQol
LSyjq4OWuUOkGeXhe4u3jaEXPOg9xi/4D2+YDXV4KZ4vA8tLYGwVaP9LWkvy9r5+VEZCxBzVwOYL
4GBxRa4QkmmnQFmB+kvyPuPncMeoo7OvX0B6t1x1JfFaVhL3NNhzF3vR39D1GaJEH78vIRe+q2g8
F9BFYmaPUPOWvxUbMSTzLMlg0pgF6Flq927LK8aYHrINTUJFoA/hE6r9014iaLY7PVw8veiSnbgz
re1PIlr6o7YeRJOetnHUxfbTIyBIAnd9wmSYnwZaLqR9GlxjJGQblhH/u7T8Zg0g9v7ccnxRP1tk
9CUAySmaexRj47dXGb3zvKN73hXG5Rk5lQqL2TaZEgXbL9jI0iAozsnEwGlBivkIjaY4bpDVLCHl
n/O2cObmmMPl4S/Nil+WPNb4Alm4VEIcYMVtdyX8Lx7IiD0ma3JJIHKhqrpM2dqW+wDxS+L55v4e
pb4DXOeIufCsN2y3rWgLlLr+glxam4q8ICPBVFw4vg5di2B/mED2gY2xmZR/vvpetss/MTCAU1dL
dcrsxm/gtIipvcVU8Reptb//HaL4k3m8VtpTJz3klt/hYYpGPe+zpLrvjoOqNjygxWVEE0QMIjv4
A+3e5iOsR1alW2qFx0ITTsNMAd7hb2YNeByygHRmrqnDqzdr24rGQ/SB4McfkPBmZCl4p5hGlbm+
ceJqPGzQb+FO1X3QGltu3Sls7mjQHhJGrFkLnvrVgGcGKBRlo9VWF9BgEuzlyhEOq8TKZS7CtdrN
XfH/9mb3yIZHFJVKybVMTd+ak/CFyNSlXmgTBFirU1HiQnvUDgWQx/W1LmJgRzUc8mI2pbOkrQaj
EPQRktzyhf8YrmIGR1wvGN6D0DbW6WJI+G3DWFIrq98sd1I1uuBAGONCoCU7r4SuEePAF8ydlhrV
KorfD2IvrvaUqYKXCEiQ26u3W7H82niJ5HTOr4w0FL8CLanVMG14pcQqHJTerNBiuRv68+O8gFPN
uO0SF9aN9/vZDzHEtKSWtnTRtAf6k5UawCPaczhUcqdMozeoTVpCUkIfe89bBNtPmG+2QCAvy/tp
9J2BFYwvYK4SUcXsEeLqGY+ckAkAQhnHVL1oqf04pU3RzcG+/qXAzETptahvWZa5RUt5WAcUKXEw
b8lDHatXBoSGdQKxI1ZlsMzt7Mdo8QKmSM7WPd317RNWCdATEQzQd9JD8UPM7IKZNImSQqZH/Plg
pRPMrNYmQDxsCLLGK74Y/AKEa/PuwrGz9XDfOwikp9x5ZBx8dbLzUW4NtUJmvVVjf2ma9X4JxDSx
OklL4kElMCtb+w16D+ZOzMV/z2fo7551tCoQvxRpfvnmeSWOlGZVcFYvbfJPrDRbDTYmcLa1nHLZ
O/hfKHwUvLB3WHyrTVyr5II0dYb7dXlsjMS5G+IdFZB5nM1VdxYsSgf0NwIboxmpkv3YDXj9IFYe
0GRcZA3yS1cqxtUe/8cI0Qk1plWJP979mcCPr3TtAd4oTzgfuysXZmh2eNZHajC9kpiN3dcHVcoV
kDaK0WdcwGQQ6X+h0thnIfl6tdIVq9KryN+hbQNBYfNDQgNK0RFLlWW/p7K5czypanm8WvBy4MtO
ldH3GonkqYCE4h2pOGtDldbWkvl1A/LhoOi3eG8X3HkhhCSIpoT+Amm8XAXKJPJLx6KC4ZXUmzWf
s1qfbmTkultqaiVrWY8XqL8F1Qd1iCy//PFOtRvx2hDw/nu4pjN7ojn1tAxvkbwuoyk8echqfhXq
QlntI54wMIqLtGYBNFygzByMTBGS7bVtdIO2pyOVeN0ZK8tL4qrMe6QHDSo3LnIuZ5Mmty3MILR5
3pOkYBMdKC/suvl8WqYQWit8753wVRsGFDincIFzYT/s016fmAy19WZOxZ7TO7JwMdlflg0pdN7T
61QfPuz/qO54R5wUBNkWrdwn2UhzEiwtf/n09HXJ+WlGXFmVqlEkMpPwQaezALKRWhZLzjC91tgo
4XbXGFDPYt0/1UC2jioDZXk57qZ/93VJEsKTuHbA+PXENC6RtEMovSkAMfOkp+nU5/a5aXO9pT9G
LpvpOHcgf8sHo2XS3BEn3QOqsu21Mm7U+P+l/PZR/LMqZ8p7ICuCr0q9kwznG43AgfNd0hHGzlIG
GRYIvM0/1hb0Vbyj4RA3d5kAe0NzRKmWqWpPUsQ6EVoFgXyP8E1G9hlcXwC8329Sub3rQc8i2OZa
aYGGq2eVY3omzTBOrIkoL58oU4AyR4xCxy5KbUgs+VJOPOXq7Mr9n2PJaNgYhTnzUt2ZHgMtZwAt
i/HQ/SMPqUJvYhzF3nPQcy3Q92ZCTSxYi7QceEKWka48L10anGgLHwZLA/09u2wJiWPaMCeihZRy
dmnwyILF39vYUmZQjkV2+sA/Tt5Zf71Iu7hy3oQbQxeKzgD4T4z2LSx0+gNLW1VwJA/VTGWZfVkz
jpg/NwwJhCAathatTbaniZNVm6GK97rim/Fmg2d81vR0btuDSlMhKWQAbHKU72azAL6Erkd5kASM
/E6IUaoAlvgnx1EHc86tTmyDZTqZKQTQ8GbzhUZWNjRllkzGK3B6bd2T/1h25rpQuo1Sm0gLJInc
Wg5Jb6Zr1fkWXY4/Tb4KxNWuF86rixmWZtwW2XEAJKW8RZV1SHYzVkqdx5q3eBWHVY9gI5f6m9JD
OSa46JFOpffzlBeZGVTELdTNVfI792hZIWypUSE3ShnqIXBN9DpkdnNtVrV5yS3Yo9Do+9noGaEd
l2g14I7B07QU5zeQic4dL48lzYZ52ssQ5FXtYbC2ep73715QdNVazNifnWEbfTwSCQzT1x5C9zBm
hhH5LVJnM5MC4dRFcUbu28sEIfw4f4sOpEUkCYEWdf9z0k2ciV9idkt28lX27/5z5bSkrClnusnQ
1f0Agwc2xJeIWO9HdEIWk7RAvLh8spA5BB7ddpVJuuUuYYsn1vPwSaaHG4qcy1yXNd76DVQE/vsi
x1PFCvS8gcSucfPgyJHQehpgantfZYkXXq7iqS3KzjGWMNabPnvwolX0Z5k02JtZLLdo92llmoZC
jyjQPKGkLSkfg3rvbLmCN8cH2DEgA3FEec2ZNh2lB3YuwxdlLRDryKFVc+9XrXoIA7WEVQAKe1u8
zQMHmJv0N86BQ04aWtdRAhD/vAUf+Cw1QA17lVh3auuFi2t8r6uFEyXM8xnSbZYGxOWwR2yzD3ju
JyJT3b3C1fHo2bYNRrFLCh8khSuK48PVa5WOD3MjwvcqGl6+80ClF8m1x3ttUje0PDh2f/NQ+mkI
lZa8QGdPjOfXFw1Qd+PO6dUQCrdPnRRHqhwQOIRgNYhzuyjFaKqmFilQnkaOLf5vh/msupRrRxna
v1GuJtnLegcSZfE1Ao/h1iGPDVz+J9t4f99Tom5v6vx1fnEZk7XlCHT5XMI6VgRIKNN2zccgmZkV
jD4bDDxGrmMZ6rIqIjarcrtp8fdg/ojGgTd5UwZyi1vEHX0jaMHvQUZQZR9xV0vDM1gluuQ5SCtY
wv/zAQ8tYmwVVM587I+MxkfMrrHDldw/onKcyrS+6bnsGBMp0ZckVGpGO77GxfSXHmlL3jcpMEJg
hgQaTjba6UTIn3W9GSoR2SbBVm1Hhen5JN0Q6TKHRO4AZkxRW8kWHhruSukF5as56E1Zno7npav6
7qL14oPDxjXaNWKIwWmvUh3imbbZw7nIsfHghLOdnJnB+sBHYTBvKgnB6OJ06rLgvpBcExs1Cltg
ihnvxSYfuCJ2zM37389TQfrbaBITffl6wYqnfEiMg9o3SwcZmhxa6RYbU2z83HS/IYvYy3ixDTvE
XFL9Wv9e6JPCg5ODoVu7h5VToHyuQZ37qYPUezN209VVfesHvljn+vyUw01YDysOOd9DXNcXVSvA
PGV1BEUyV76fQ6ndXwDkkAlwmcUs022XTdpZB6CTkjaAl71/YMENaLLbaJkTPHf+bjEIlWgMn9OV
r4Gooh8BiSWxvjjIqRS5UtOI87qXaqdQl4v+PUKyN27n8+Ob4isgjGAWV0qJGV03FNkV7p+oWwvc
fkg/+NuK0hjZbueYaobIBrGkffkJgB6GoZnOAYh8nhBC34MHvWht2KMO7FDcLwZLhEg9Nt0ExIFm
Ue0vBOGqzKUV0k2IvMGRqW0S5NkTUIibzQVXb9k6e6HPzcjtVNAFtGz4SuXq3WbWnxWjQ3Rv1/T7
fRwDSCOHN0nNBVSwiBjeDSeEOrnO/kZ/ZdJg24fRku5ilXT4Y7e2u63/6XSK6YkAmYt1l9xi/1HJ
3b17J8lGSZyjNQnUbLTgoSUW8vwVUfFvRJTnfQWHcCBI9mRhFncFR8HLuFS55q7Quse+onzALIHY
rjUs7V9Bi3a/GSByNpiFSIsHFcI2e/F0EA/AF6cUnSATyQMrw0ot+R12XYQRPHsGK0At+TpQu2gj
DWaSuipDQ0IYyzjPcNDrCMTRuubL1wPmTrPjcPEdUnTrM6v5q6I6HobiL/sDXaj0SRUactO4cMDk
abTYjNn+3F50yMGMUqnbfZSu1rjzNQSixbutHLuLKVVLfnQ8S0B3iqb8K4v+o1FHVbVMDIi6txIB
MkHwmHF4NUuLhS8Oux36UyJM3YiwTp9veLJq2IzEEH/8jXJyP33mT2LyP9VT58ZBfSh9yMVnP5Ma
qACUPEqbm3GYFA7rJfFj/nPD0OJqz+MuBckMvXBN9Gfp2drUmZ7CEXrNjYW4LP2BaW2FlP0ZowgU
OX2aAr7HnJ0i6CqTMYxaCoenPtlO+ZzoafhQiH8a+RTjQhpOLagI5p5Eru79syN16duZnclrrtWv
HIYh92876CvZL2q+HVQ3IQmQdZhqhfRdtk9+KjWtQ5l4ZV8/Dkm+NAIUxXTVj6co7lWVxvnLT0M3
HTDYv1taA1yUFAVJT5VV+BjJNC3g48GXud6jvDyPQlCkdV08E42yxtfpH3oT/1ZQxkNka/i3wet6
c4m7InFUH6TOArEPeGEb66tx+G5J9A5EcvkFXCdmMdviRab7yfSDsew4NHMFeG6x3gPWnvkj68+1
gUfu20oHGniqlB4/jHinOX3Ovw9Guzlh1uD4/2sBm5nrkjmhtyy6ZHLvNzt8IfFFUWoNZyIKp7cC
wVHWLDIVLakUxHsHeAoOBsE7ZrJvsm1ghpCS3MC11VPZD9yNZqV6OTLOTvIHkOP/18mhEI8KsLGc
0ACG/RmL9drNk+4aPkQ4IO1TmD2/LDxFx7pR+UaI8JwQRqOcyyahOILzz6vCPiCqDnpUOSPDV/w0
V2iFXnMnWLJdWgI6t4mEQQHov6wPTsgAEOikE6HBm1orabm3499r0bBbimlFOY+a4srdbZGj5pvt
fAn9ldk28PKEHMqPRvjSaWVxun6rbmxuessY0LTIYz/LBTPK4ENjoE6d8ugDpR3v2qG4E+YLHQr/
B576uRuSaUovXPCmPgix4cP6Tz/sbrcH+iXFMCxn/JXPlpy/ZUzffJ0w6dhivcaU09UGqX8LiIJr
YWsh0AAZaNqLrWQUhM4mG37OTu4D4aDU9dxs+6/9vkwBNLpGzKzjbeX9MnKEAt90sdVifRfpY6IU
0yztjG8Z1QXrslBsqtLFAtLf/Euk3Mltndo7yXEMVVgu7fZciq0qGnYxLJsD2JMEunYeWWiXX3Pk
c8ctL6SOYf7h6JgAXZSy3xe0AM+R9YvwpSc/pIUs1XrFs9Q5qzDgkrASxwnNmxnrKe50AT++nGYf
q3YSpNCKbPw1l+s4Kv9aBjNdt+A8sxgjFFIuGzNQQ2HlrCa1vFbHCtFFQC/Ia436B4iNbe49l4Te
BSYith5vGcNk4ZsEWh10Ay4zW1m2krw5ySap+3hFu220UV/JP7eXx86BgWMCOIEAJ9Xq2OndH5RH
e1UTNBiQx14j69MUVQD0nzKU5yQrBbdIGG/t8PsEa4N6QeZVuW3S4TWSglnL7PEq3qKN5L930GY8
ytsmEWQRq3aVwMY8Hqb71/khn9gkCzS83je8iPYi9G/864T9X/p4DN0VfvIOtmaYbyebQMdzZ6Yv
m3U0IELZzyTLWGkSEvN2VoEuJoaw4zxq2QHSKOdS/ryMTE98EOXUraHiL11kwC4wGMJ3Teje6sh1
VMtDRJZJxM0vs03AMN+ulq2cY8iUgADMeLlSMqyqlqR19t5lQFfSGNyk+VCT+6n+yJe7YQvHm0qY
voI8jNARw0kQrf7yVqlPVL6l5k7kzrAxGwYbYC7xmzIRgt49jclMTh4A8J8yg4Np4rhPM0dfpvj3
BaZOtBQ5LMRFeR/XEumN3zMJXjXRnt2XhQzIV+eGISFeOF4pA5NI/HHEin+UOrS0iQbGV1EfXNqR
9oqLkG8BH0IWN+KrztfQ6Rb/tBrflMSNHWCPlRCZDmrocmcI6o49eooennSHIxZStwWmHy+CcLD3
47T5xti46KpurkShFl7VsBH64wZ2GmxEaXuuykXG0xvqr25vrYLOpj4IJL+zIdNEqBgLWbolYdk7
CtHqlK0vF3UZqUfeWPbK74fQHBMC3UJ5Cvmntl0aWn2KPAFPr9ZkSCLqlop69Ja58TVPhnekiINC
6SmM8aCYdki2z8hHrGwPu+wr3N1igK/7zwXz27dAmSVkxQtn8em+2+LgOXgPt+ziQyC5G59LTIM0
bkyedz34kMKJOiq+t4qmsiSOVLEeSU2I1U+i12H9E6bTuuDFUbEtapPUyJNs2R8/tjP8VdqviI2q
6/+kE0pXBlstvyr/AKlgDsAN5CHFjTHUC75Ri+AzZjaoNW/yXutnj1fIdZfQoT356NGd0UNGAEA6
ksMHQ8DegYyaYR+Ip20z0bHWjb8Yl7/BDtoKtSZUljEcIFMXR1+rVr/zTDpuaoNMOqPK4PYwE6cX
vxO8zWkbgYpKByAU0leVVJlWrqBi7O9Z5MpXLZKGzl//c7wJm4Ibfowug41N2En77m07GGAgICWV
klcTxIerQlZ+BOhDzJZUADnK2gGBZHuY2mUCyyMukWlovoIuGR6xvGhYhBTwAJ2/eJ29wJlaPVbB
25gUvqsDZ3qx4LDCaxZgyD0ZvTJALbycH/NdbTjZytVFpaMr3PLrAUmFC6DLfWOQ6Nve+CjWLOG/
gAN54pAVOGKm68rXL0pWInNwqgtsyVVBT6LLcAK8kJpKlgqEOCSa/huYmMNTv0zUtT4jUXZBNrRp
BUKzJE0AHZ4VxWFXSrLCIk0mNvXbYXTy7cB80UuiboZc6+nT2gEdi0GHwYaV416GJgf8uPW08sIQ
nESSlKgJoiDqKkuLWOViagCmUz8fuGXPF9BUAHJZoJxk32XSmcmfexvLjsIzWAv9w02kEPhxEuzq
aaMYL2p3PRd+cg7Wy96GlYM1qSnqC33E9+0xDgTn+kZlL/L+s5wk2srQtn5W2hdpo2ekkypmLnkl
Tu8ohhisQo0nvM1GpTcowJsd08XHb9xFAAPC4oWIzkKNjre669v6eGUw/Z0LVpRlPYGVDrIJlQZm
ocg29fIBC6Tfx4U94YjHHYl4rwo61dDa4Slxud43QInBoIGHwZqS5XWk5CATN9kNDvi0g8zCyQwD
L48Wp9k5HTcdvdzLEd0A60d/X3TVZxm6p9axE9ixyZhUcHZ2YlQAgiuHNimY8DYPsenaGkTDTVEt
Z3TjYpgN/169DJpF1XnO4gWU5qiySUg5owxXUt7On7hbnfPH3JJ+1I+ZyVyi3DJ6ltZw0iXngTmr
mnXaUCFXagsP+b7K0VX0+DJEu3moKnHAO5n3rslqad213t7ufh9N17sqIQr4SI03bMJ94jgVrelt
TimDCnUKLQdYhWI6n0MIIb2G9sfjHLNx0WCj5Kt9Zoou2DgYya6fV+4FLCRVSxWBcIwAPVKBQTJF
a/0YzTMhVMqxOv8+m00oEHa5VgTAZJjhLhAZd/BjablnQCcHe/aZD8qAovUVHPags6UhEQJCVYJK
SvhfeH4+LJMVaXbyroiawyafLinhOokTrtG3WZLfWsIgz2kTouWx7XpjpSPmgtsG5jdzZ8PxypcN
6y+FMB4Q/baPXGDVBwG4r9wNakoP/jiPXStFziY+7PpikZoeV86qwFstEqWW+SavsgYlL9DWkYBL
TlZd01GrBA1XCSB1CzC598uIB0NcDZsCBRjitYoUOOaXgYAM2QQeHMmAYey7m4ZqCQjmhR3bYB+y
SsxwNmw3oyTVCh0zagSI3/pcSXReAB01tfxB3EBXPmxPxghknb9nFC6qNoBQ+KTYo+e4/kuMxUO/
Bq4JVxkdr6x2i6PDQq2aFxRDuEoFhV8kneRYm8xnqG7PcMDXd/4LSckS4AkAmWEARIBYIuAKHMq6
s8XpmbxcoAU5xVhpftpqDf1+WJr6B807dsf6jwSyVRehuKc1hWlSwI3c45yBqzNH9hMaC+HS2NQH
4JwgjvQHDe/0JQ8RySzMmlfvGuju4MuMxfug0z98jAT8OY6XT9qvgefZbIOyTMILJIebdMwryJMS
9snQ4PbI8QZcvjkIUPYn57RUW0mgYIwAB+ZnX078XoSUW2jBttzzTD5o4LBLKksrfRZcjIH3dy5g
HWWSBE15cUPWPet+ajIEpsxzcZ1NXvbthZi/BlHv5pIwvL1YvTFXOETSm1KcrvmzLP5XiwaAT7Uz
HYvlSTFS+ZWh0XiFzp8/YCz/NZWOnO7KbtKWc4IVbewsuVGA5QaIuXnGKay9bV2Fl3mFXxGPAz3t
ls2vMx0wXJqMnGp3uBtQ7kEKXVCKoWCIGgDEKpo428stWGx2e3/bFA+hheDPU7oxZoUQGkgNob8J
DXtzLLdEHRfj02h528XgpwGzGF3kT2O6hn5OicEV1dzQu6VyfVVbYqDHxY2Qu+aHoBCQhJ+xiNdy
LPJ6UEZ3wjIS1/9VVmU7tDEJdmdhyM0ehTCGc2yR43MC9q/Soc3GTM6UDthr4xY10jPedupO1j4G
HU7/ZHP1+YKNPLDC3X7IlgUnuihmfMkrE9PCRSsUuJC1mHYA4aBOIgZ2+cjglVXxY8RdeYVFbl+V
6bxui/eZRheNNqbAiuk6+xQwuIS0UOlGDQ/QeNTHRmZ8QFI5lT9vayC2xksMISGPJGERz5eQj6FY
bYNwoHnyuFRKDpgkO1LFdNUwfrt12YNgpKupoR6IYsb3wkCimKj8q9RL+9fo1olZk2b3xap/YLTT
UOz83Uy6/AE7CrG1Gv6bpihmHR4W4c03DxDKUkg30gsc+6yymW9vXzlAqQmpAyhVypDsbvlwVlFP
480OimpimsOpG264UDkEYeOFv/eaNddwUSunvLEreLyJ4Ox1spkCeY4oSFCrvvfKhMMaLGtB4Mpc
TeAgsMuuWpQ5m3dGYeC8sb5bimLJo+1CB0aSJjZJ0o6/eUq9GbaAb1TDPpKJ+VdVlq5VlOEqGRe8
sbKNRr5cKvDZ1RSz/EQ7JnYYA3m5Lr52JJnDE4FPb5ZDaZJvYXcVCLTbY1qgp3hmh0T6H+4cf8Ti
VF3TfH2dYkN3iByO3A0ZsElRV3mR34rO7yqPoHFFBLrDmT+QoEVoR3tBRUYeIy+NyQv+YMmAStWA
IV7znNwad5n8G98iKLWKNvzQgX80E7JDwP6L1wY5qNC3fs/lfS1m55DAqYASEfPxQ6K95/HiPdIR
Z1RPN2fBv+Dytm8x4okepyhBUeVh88OU8mciyNMZQ/3pdXEuswyQlMfvMW0uaDu7h9/Hcyj1Qxz2
bi4f+y/JyxMttmHRQ4rAyYRQ62/2PP/LHkeqT8rSVJv+SkuwBtd5pzDVj7B011NpBg2bNgR+vks9
agUoB5F58osbZSOcG4pVYY8bFA2wayjXN52OS4SyF7SmoRCAS+l9f2tTgmSMJUkWb0ptsoMo958L
MIuacQrzygM0BMYD3QmnEFdKSnGKE8hm7H0yc1XMvjkiKDd4Y/oGJsmjJFUslcxKrvHBpKKoobtP
iB5zFLstxU2aC4ulKagyR5833XjqXT3INFc0z9XiZVoPmXUYahY1Vztw1gfrqGDpA4sxAWgJEYN/
D9/2K5fwb/uNWFK1+Ml07nIop5m25L/rXS/gwYgYlODYluBpIt7mqX0FcMu7kYhCO1H9Is3rAJpD
XtO6vRx85iANSOGMsXtwDcvYEQlUnhaWtoPIba4JqxM6izn4xmA6eibI79L8msKU4hWnPVkd8xd0
nJ/XATAj0oFRQXWPKJUZu0SzGX0VdXvk+51/Jh9bGLlnPJ9l939Z3+9SlSBlWfx+f5uc2ZpRVjwG
INzz35Cjwr628i3LS4PUiG7BTf2lG2oi2zroohuKf/xeRqhmJCZ/PHaZ6p6eL2UuwM4ayWdIfudp
cNOlcoavMm5HFCDDvU/JvPTywhh62ATWKG3W9650ST/aEyNzAIXud/zHZBAjUhggaV1pl/60AanN
1Ydef4mw4yE/hLYhuGk9NyBtBnf5Mrl2Wri1+1jeZPTnmQ5b3CsoX81W6mfNPbN3Kycj+WKmVkyF
WJTfOHCx4YnL3E3sHJI+H2rC/KfBXeuaa9K4TzqH/dkpUcJPLLxtsm0YjOqwRUP1t819H+P3O6il
mM7dTelEJ6OMKnVvkBUEmj1M5tHjX0I/R+fb35d8JxJ7Shg3ysTGyK2eRqnHPFm447nkqZag2ger
2/GB1ZkyMt1IGaazIaCbwCvgUwKCmERdVRUMM8imAD670za29BFNvAmprbF9gRZqfMkXrXAskIBD
Udg/vrVGKYlf+TLmW96puq5oFYATx7UNYhI5KI0ThSRxc3xu98wERH4pyE5Bb6mi391N4f1XI9S7
+E+LsVyd45Jc6y3rqRgg8mh2CI05Pcu4TYoImgPduiju7D2L8vGcA6gL98ppKjRYrL0BrRADHsgJ
A6epLQ4BJxurCKOPJ/t8AuN7WWT0MtvyhvJRIVSPzRubhoKVPbyv/kY/FlYYQahFipUdU+mvnHc2
pMEtYTKDJ58w+A5EoQct3p7g34SI1vUAm25omkUS5Eo1DDPt8zUHXvcl9xYiV01m+Qhh5o6taCyn
lPWGaISYWlcgENXgjUow3bNQyE93ZabFsOuR+t5WlN2t/2pfjJOm/E9F50jJeguNSsQMfW9DeB7x
jOlyZui++jLk5yAKxU8xvcEyx9uqcFXIB0gPvgw4lo1ELPbHJYp/2mmnMFyeC/lvv2QNYyNQ3Lit
5610oLSfpeEPml+HxNCPOJPIa49FgrGSgfrgjQ8Zp7q0EE/uZIWkPzpFqH+Fhi59Dd7weQTKF78T
gyapwyDfoEC4pT/26fsgZhGNnFGAdfvLc0PTw2iXu6oX4APuA5dOer6cCqY7uMl/Jg+ATppwBkKi
dsganWi3cinLno8ZgA2EcraYEc3YEHyaT/VKKv6lZFnGyfe/tXGWm8uY9natN9tC0HPJJwGLB/dp
U0ljLH9AsBHGC55Bdjg1cFBPH7w+MX0U2vx+S5+OmFbaJE+e9zpwWzU38qxE67pJ6BTPUHWrVdaZ
4vlXxf2wGyjmMU4eAgtbnM28VHOgZdJJ60HVNqLQfQmZxrvRKTIYGo7DG5x+n8BdWcTGk+6DXHvB
ELhEmaDT8FtGm0+/MQip1OaVujYyLn0Osp6PsR1+/X9FmDfQ25JGcPPLb01Pme+oEuJsivX+wlbN
LqHL6rw7hZb7TC7RdpFMyW9rWNy+nuHlQe3C147CEC4zZUyriajuMZsAfO3Nfh32aKQpDoDlHkE4
szFD1zBp0lXYD19ZlR9US2Wu2mb3Pv54j/YIYPU/JfI/SNcJb1INCiRbmCaQogMBF69eRf7d6WVO
fDEXsb9qAo23HHtz9gOUZxTh75Cop985mc5CCUYlMQRPyJC0F45gmY/h5IbW+H5TYlt3fsdvMtAb
WZZHoI2pPuAZrg9mXfytWSzPY2WvSIPl9fiVhPOx6K4UIu4Z9P4QsQhZjoxLkhIxkPTYXWd/sQN5
aeEZJSkyeC3kLma7Wk5ThSP2i8+EwlxwNfR5RvAH7ufsgvBsaSog23HTjrBBINw65mCz4QkBg2js
qBGxLTKJ7tTpNngJWTiVYuqZnjvXFL/l9KA4RBVwF4LpMA6/Kspj1+aOFcCdg/pc/pSwbUD7jqAz
ZIO4x7j8ZsiGfBWIwsSmPjBoYUATFM2EQcdDlQIYLqXtSHFGP87yrxvfunlPMogoNAX9/Dc+LQvX
vHIemjuq9OdpxNsFYdHPGmRTuL8MsQ6vjB/QbAznIs2w
`protect end_protected

