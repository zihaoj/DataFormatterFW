

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UhVeas6K+zJkxzAJ/XH1tiqQR+XspsoQJ3dEE8+NZ2li/evybvRR2CFFWlkn8VHqMN9rvRtldUOC
AgZ6PTRk7A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rz7+zXWBctYQ/50cGVEG3Toj4CInTVWZ0c4T7rfFyHGo1fa/YgddoAqsvH7qyYwDZcrYpT5hpEmn
cFc1YeIlYloc1EaeTJDtWuPiIlcMz2kYk3MBHTzU5MIkyzIkATn2/OxceutmubtSsvRoimZqpVhu
4rHEfrUXr4U61RD2nsM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
X3azlMHeEDySdNGo+NHRLVhUQeoDEhghKhi+IvY2MUX5S5C0HbXWISGVnlCl1zEfsB50hXL1G4OR
kOAPftYogI9OPmHAVfLAUKfW3/AebOq0Oykvg4+sU0VD1VoueDHkcct4AijoaqFAjdFhbDGl4pQW
DdiL7zN1Q9uXwVQ6Aarj8w0xF1fxyiYw/e32FnfCVuw5GVRfdO2e4Mabu84yq8avdSobdF0oBfoj
/oaBxlsYxSoVPNb4cRBubTrF90rAt7/lJgIHxnoLP+3hN36gpW9tkiytunSogmKo44iOBbKcrhIg
h2SQQ87sKJeTDGxyazeT+8OJho6YuMPNaQHE6Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mbIlGrXZMmPot30Jibhwb5d34uJ2kRrtfyMuP9COPO8/wvMqVlHAjEAFm9kAbyNt+P8a8ltkrgIe
noTjfdkgT/jV4xOK8Loi32GdoUncVm/i8mHnDk1HwVDVW4H6PgVoSZZnrIGUYTvd4KkcOFQX/TET
wouLW2mJLw5aX4PYJF8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TIXqnUNEqWbewR1mPB8N19YGlayBdy6oisZqLFfYkhOvNm8MeNH+aT/Z/okD6Sp1ZlLyCqNZtPj3
uWjaaMopcBv3dk8ixDHEmCttVJVrP2ApTlw2GLb1ZMtfCxABRbJPoBtZH1/84uFe6qY/4MD8eKuL
Fa3ZdP8KVYSDqILI+DH8OjyzIboN7OOExrlN08BcCsADH9MiFKnBH/FdCd7IEKuMiGEb3nNqHxCE
6yuvfo2DzFmniZXdPqWuHhYF4mhlrdggna5jpJMAryPY/Z/TAVz/dbVQjoZ6bsFSUDgLnTFwG3cJ
osaBYwPy+y+wR3KCwSlWSJGiq8VTTAnzFVzYng==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6464)
`protect data_block
PCLiHVfIAtU5rYnWDB7yFNhO7jZ1vbU5SR4qEvvtyTfpJsP3nFdKrnT4u3wPPVov80OLxuDrvR25
RubKo2QfU73+qfBi0qHVvEXY4grEugP4RRfeJBERgRapWkyznGe/YaXpkafZINZtfu6Ba3yK177B
ISydNkfgHTi5jYK7MaeepM4gfKcJicZtNL/N+P7PD8ELhf6zbIFjkLEYyeOkiZN2foFG/wrJBKna
2mSGSV1BWvVLYgOMZ/fxkmp2Ubvy2AwFT4XhA4shdtZvL3rrOe5aunEPfiIE2L6Igu2MDolWR5yM
HwT4xAL6di/MUiKoyU/iLvu2y+fp4UpBph2sbvLVGWzN9DtLTwLs6gn5eX14Zf5Q9tCB8m1CRxpL
QFmo4lMKThD5Q/JrPDmpUQ3iPhbgwaxCQ7FX0+vGM9Tao4GpuvK8HitA5Ahb/TIoWfLbVb6vn8qe
MNghyTBOsTkszBK7q/6V+7TL84e3NQ8VuaHYAcms80Vj+iqB6w1PPIFF3avQe8jCamjz40zGCOjI
8HEVEFhNL/qFSUsBkTadkEFjgAmROzgD0RyhS3HTI1qmsCHDp7OLru2FVck78+GWMcsSdOWbI5rb
hezsChZJ/9bnDtml9iSHnKRsjyPXfQfqE9WoGY+f/QG9DyiSY5tYIAAaULnfOey2mbgIpQ5F4tKo
nJZbcURWoBHu/dYZICTkgrxqfvIVDE7PcK53DFIAy3f7q599vbnO27Us2K/sXPFFfraDWTFYNKZB
qSB59UOpNy26QhBIjxV5cV4TQJOSSXouiueisfQfxFoH0VGDFLO8BF2fwH7rQzmDfYgAHFVxKvr0
KGBid4zYsn69Y70M0xMZABIbSwPp1v5bJNrhfZgaeOsZTOTB5scKoAUuk+72mcal1FeHpfnQaY82
vNhuXjnPUthGnnpS6JKR+HQwFhx0xwezbe0JcsLmSIi2LDJ6xvf/t3qoKE67tFO3S2OnjzX3kEPs
hMBZVdusULNbWPvO9tBfz7Hdm0aRI4+AlCwvErLOj7Dd5/14mJVvkCdNZPtolQPvU6WgI6RITTux
G4vM5TwHl47xCH6c3P2yMc38f8yE5yvn5a3ufbNoq/4vGmgml0NoPoCM5qlsiu8acJcUr/XGlVZf
ZFB+yfCPBBNBcgOHAB3rA6Qzq6mBzVAi1JTuz3/ZRigHHpRYtk63ej3A1/5sbLZ4COKJm4jQSVuF
p0tFza6Fu65U2uYo1Y4t2EQEy8DTaaY2L1PDdhoVD0yO8cHKd2vdMlX6l12WygV91/UYtx4YY64u
OijZqwEcAcEOmAQD46Q6emVq6dfJnhDXN642ayMYU/5TWEKoMgIH+8vINFlXQfYNBQ6qSVrFp9Wt
h3Kt4dV//JxiKPa1XeEkhB9vZ1sdLC4tPfYPaVMzNLWMuFFfC86/8STyAnxui6BkOXQF974/wg5a
ATxUpA+UuYNHVbhSJUeDI2X+qUlpGNx45BmcscirftvgaQR2LDKOETAzvQJWwXEAhTyjg7K82yH2
uc5sY1nxsQG5fIJYYM4dSP7QG0ofd8li5cKAAN4tX/f7eTiolHSLSPArqYB2l/xgxbGOOGJ6sb91
k06p3RPftJLyRlftcl4VFuqcj4XjfEmu30qTYQ8Irrsf1HTms63bQPabnxp2iYbxbqyg2nG3teYk
be0odjGPsfD3p3FNJKPCq7GnXKnmOI/4ZXfkM81p4myiHLS56V9O5pdTKa7xdMNMQCdlA9xgpV2d
+DagSHB8ZtpHW0r4xT8tcuwyLCVrj85Re01mvDalkb1btSM7VNgs2Dwr+wUVcFSW5XV2Y9uQkv8V
Qgol4Z/PJAn8f/0UT4ClFmKGGUbyISK90dUAWataV/2d9YvY402rFapY2PClCGtlq8XKlvHJ8HPT
ofpGs3cdoNQVU81Yy+2q/7jmL7iUyFDxIN47mkGz4IsmgfIZTZr6hXJa1/zyILUH+1iKKBvfupO3
uwTVq3S8u/yRcvempClIY0AZwoCZgNL+OXbX6u7y2ZSycwM/7zqN3Y9nstT99v+XMC15+OEx/HfQ
0iapzZFGNywtHHvOaQ6U7ljQwHBMBDiiyhWdWOfeyfqoF5aObO+P8pb8Ktfg/cX0BRDe9mWhSzpV
QzmJR3AvgL9EiPxKxymPf7ZQQtGPCTyTwwSzfj3hxWwlUC3kA4aPnP6ENHxaz72XxUfYVmlkuLwS
CiGuKQRZoqYI3MxNtDh9d/g8XtVi0rrQkv388Z3xpdE76M1itwlAaXrW/H3GnunIF3+1DEw1qLJk
5epbqA8FX27pEHPmItd1Od2R0ivVoAwoaV1q+ddADWkTSL4TZQBUtij8DBF2NDCo3+JiLentUsBv
8EFOzK0F16R/uL+PqHDL4pGmj5D1R+cOqYlUhJUT1IUaRNgsMQt+WOJW+T4SKeE101mbH/lbXO2c
uQlvmZF6aCyCOAnWq14t3IKCg9eROVMlVNeZHkKk263nJ9e2F3f3qXFcLZw6DAhwhLDIuyN7CHk2
hy9Qh62kH9LBbY5kyNNtDjQGjnGM/4dpKAoGxpCtso/Ypzq37/L7Cw3bXbvX3URo90u5Iv75cF4A
/I5YVc1yinHbceWTAPCbElfkqJwYIQ54e8JnyVYxq7zhLTTWjnKOhy/w+6BnOW3TV3TddnKIve67
hquQ+jO54Zl4QOqjtNYjsEE8Nvpq3bk/cs6436un+G6xZblp8KyLuPd/m146MRPN6kkMbN0ns3aQ
tJEDcksmybXWfXYvt6OZUXU17QGlXHLyU0VdBuPVGBatveR6GIX8VYJStYfjw08I9M4MezzQlYjg
QR04Pn5Kpec5QQKxevcGkvu2NvKlOMu8FznUworczMn9KHk3YRct9Ow6TXmVXaMl0cpPQBn/EBvL
kK4rvW3cC7p9IWKpiN3ps8l/bblpVVTNOCkjTriIQhp2Shjm4OtVIdWXWLWU3gznI5ubLDk5pJXs
fwgQUrlf8f/NEyZSOSevlM0FWjFLG7un3u/QGt2SlpAXkd6N2JONfKz52nUy0GR17j/XWIne+1N3
yZ5JQkgf7TwIyxMdYiG+mKx+P4mdVYSotVX/oj84sqh1rPxmsJhND1o50QOqeawCZxsdrAgw2K3Y
MYN7KMheoJKrs8JaFQ8J4eUMEtpws2a565SVAJsx3WDj8eMkqaWfwn3FFLndzb7VtnTIklhd7tOu
HChEEFhr9YcQuPX9NynuLKKXLrvTxoHYXM1wr1AvsZxLjmvaJ1EneM7KFH5hfzTg+orHJdfFcGeg
IWhnpFvH9vig5bE5JufDQTmHTNdiGMiBV4SKVLECT8AXPzFQvhr1A8O8wZrsa87akdS3Asn87iQE
6RTD7gtz+MmmnfRmxTtcyFurPZ/8+OhxExrzRmqANuqEfSAQ6tt5wkX0J/tshvR+qsDqc7jswO2c
USeXZRN80uYBOb6kFv/YqB8+ZsTCNO2li0emVvsQNTNKpoSr7/4dX0xrkV98zaNpWAaLefBzkKVn
TA/SfwUgwXQXUYdTgV5vwq6fM8cWUmDU1f253GYNk63FsoEW910mDFuaIPuPknClXpiZw6OUCF8y
5j+jaHtyPs88y/og6dHy5MJGeCj/OSGMbnQa0tVpexjeXwJZQF1tX+41FDPwU+an0k/N5TDvSZd2
OtPl93YosKn9a2LGDuwKA4gVtSBGevmsfnqD0S4FXIr569lwriP3luaukMczDjtbpdi/BZRj198F
pJC4Qn7oZlaZgr7XZBeru6ijuMJRCN/SHJyM7hG/jTpU3sC1NCIIkFKxC2lDJuStMUDxi1OWTpk1
0f6Go6z8Q2T+aBhR/BW2Z4wyWTd5JpJ+HDmuMYWJF+LWwuQlQow5d8tJyAlOftw6dU04JQUGRIGC
mM+TWo229G2Z2p/jLmfOALm169Vj5eEaWqP3TPJZYyrO+6hhau6Ugu1GnCXdHtId0S1XHGA2dBX6
453tNf2Qh/IFQgJhTkoGPye0W2AlDh7SkJeoFDrrNv11urajroLM3JqKU995Bz3Wkx9aCp09vcJz
tRtIVWtPfcxFfc++KlwXuSxd0Ki7X8WixuiPtfaZxA9Os/qTbkrB0kF+uv4g4cz0FN/1n5PpeP0E
ttTV4EQwM80s5d9mapf5TZv852Ti6NFGSwM9WFnpjMZtHcEQK/N8isBjadqLwwgS4Xali1ZUozK6
V4UUj+oq1DxtNTn5s26I0wdhtqHmGK8TKQd1+Sw9C0PVmuHLJbnraIZAr2Zp7Xtl0zGLGIQycyNw
fsSM7Ke/S1KgNQ1espvf0zV9tVqMU9mLwQ750Cf5JUdtIQM+nZ5j10KfbSTpuQ316aKdH/eXLWIe
0pFXjyneKjtx87Z8RBByoNcoEttyGlmvGgxkDJMqwuMZQy57TkfLY3ZFWzSfAWexTC8GHT0x+tJZ
1fxtUmAVtMVIEK/FqwnVOTeP8UTBJ5ZOjKiSfZmZaj+Ga3nxad8roslxjvBr0AUJlMfNI563jzDI
rOHmWyvUlxJGlLZ0BpWKBudKKWmN62psLeBk5yjTd/UVWuHX0SfEAgqlIQRIxKAso9iKhyl3nb/w
gLjCvWYmuQfvKSIhhwQcRiCrh63k46IVhJYK37N+SJiXY4fkwmiIFFo+NFL8yvXs0lp3S6ZIMsCW
kirdz2PaxPwkOWTetMbI9NZY43iNsrnejQOwQXgvNJqfd9/lJmQcI27Oz7j73FRagmmn4zVIaXuw
ecErNAagXYszrR4udCd/UcrSPrHcUrAwauxWMW2lAwOX9AVv7F69t4PZqRlcXT+nM3NDfpAsZ1Zo
Xod2gMd60MYPOYN2htdzy0kTVvs/1wnKEXjO5ENE9mO465Q5v2AIakddhYrhurQCqzL6q4gqdhAU
0OITLxwVi+1ERq9jtQTOq5+ejeT0+vrdRDJBUct0hMCYlHSfmKxiPyY5HyEDf/IQM45wCIWHN66E
Iq8L5LhFWxB9cLJbxJwBV9QgDdXPIl2hHHCWUQsVv6sCknS6opSdHF006lbcMfT+6AfdkjcO3pmS
7h2GWhR3lWwia+FKeuVlgVLWkNJcPKNWp3Ssobceag8eSAOcOWXmwP3llFC5BEElDy0Iizuzxr8W
HTBTm3MML7rHuzLgeDT5N6zPAKn+lpIsT4LvQG80oPHr6irpWc+eFK4oVKYGxFEJa+K3tX17ROgw
vJxVQt5voGwDV1gJAtOOX2HaStDyh2lT3TQKriyN9NX+oCSxDRyYC1lxnoe7bJqP0PONbjMbpPG6
vmhCVPaVJNb74iP+D3B77MT1xcktGmDzUW5MUl21WqaASk+Dyr+WTACe/pUpGwMNYovY1mo11j4B
MW67kdIqWUOMVA3LF2BwgbMwoDpVGMR+UjkRf9Hoap39bCr3yidxlFHXjFS359wrxoPM74yiipxJ
cGzjx+OpO6DwFz3CzYNLapQwxVZPQggEOeHl/zHBM7ZTzEWQws+ECSIzDre6iuMxcpVx1d0AlwXi
2aRCwLLN8M/75TeMe9T0XcWvLHEXaDWlq81MzAG5qeOSvCZch3fR79pIS5zwZ4tfC9gvMTeLg1o8
dJ2ZF7zU2BVcx3tmoemxmeGur2UMZw53lhYpyRRXLhYbEPn5STitlVhi2iM7+EjlDrlbnon/YP1O
jfiEjFAi/1wZsqO0weMHb4BlRks6Nc+QEB15MUu3RrTi1ihofqr5kEATlQ4vQWCg7btm+OCLFW4I
Wt5Oqavkj2B0SEu8G4+U+5k3LaLcUILLu3FVJUwOkiPoDtwwlpfsnj6DvnWGmDUGI/IqmOY8qdkM
cF7IogO9Yxb7/s7Sen9fmeL9D/w1/O19fU7uAhTm0yxIsVtToEEaQrRQBlmDfbcKcehofaq9zW8Z
gB4zEdbsojKNFSTDbw02OFso/zN84mWlvqAPqUITOkf3+sxYhxMCkOYfUFd0vsc1ZPt2BD3LrWgs
MMv1uxRImvz6nmIqzPsd4060JbrEoyi2dvQHO9Czx+RreFCsvaH3NaoAUL/Me1HiEkzM15jFEC7w
AXVToTfA6fPT9/UtbxsY2S8FoyroC+eVzaBKXRptX7XaAOX/12rgz/8WpH+kJ5y/CHxDwC/j4Px4
jguflHOPNyNWzpyNy4FVdLTeaYCIbM7sEuSVvrpAN/T/ZtZ2xBECkXqC2EsdNNXlM1dl1sBw2dyL
DlSa2wa5a95uH4SER2il/5bywiKvjSu0/OXx9JomSfmEDrh0DY9VprBVkGNR71m4sUAnTYcn5F7s
/bxnnT+ijxZVP2QzCk9CNOajf+A1t8bbMxmrUZlDPzjkyR2KC+Wt8wPFOClca29oQYLQ6bdQIdgI
kBR4nkMcSCa2R+3dQtFlIVWt6dqpYnYFfwc1J9MBEGAkUInL1BPRVJskLI2O6PDs1Z/L7OQsObNt
Y4ToA3ik1t8AEo2o3gBCGj/xxiVJ9HMih3ggOlVgfb1naaoibOprz+DXibo0IHz0OWh6iF6sGmMK
qbV71bIV0vvmFtOovyl4zwanhK1ZkTzyhG3qCij5gXqAfensrzhg/WAuTgqevnNeX79lWeMgUCzq
m9fReZMjBd8UpyGUvS4Y58sYGuXXqqP94ZSwV49+Pe2JmzRe5jHjllWLHy9i67vJL8E3vCagPnrI
X5X+9IMCOBmgvHqFBrLAU4jxRFiChTdz7aljEbCZ21qkQsRDnOZfxLe7Givz1mHJ9cipQOTj3uqt
U1woIl1QJB6YGldlzctL3swi5psSVwOFydm3frMW7dVoOyIZEOunRrYJ99tJrmZHaO3Hq45yEfZx
yGTKGmTGW/XTBWyrYJe94PQ/OUo/MqD5v0Y2NzsTLHv2qr6p1UNjvsp57TwABE0Rvf2VbCggrDMO
Wv5aHCwIYNx/cMWXGHo8ltInqZxoqstUC3ezISX1ZxhuFjcA7gyQGvs7yulXAyvUD3kgiKw95tR9
5LifvhkW1kPD6q8+5mOcNr939AjbrbSOM0KvXM2NHh3iovZpqEkQkNjs8CZx1Qw40CHRYIbShUyw
xftj05GbdvMZQD3RR2zOKnEcCOwsuOYPBZCyW+3x+jBp73QNWbkQhQCT+4lispXYpz8+yJYoTPmy
ZzPKS5rVv2g4URP6Lx3ve8WvVklht/Hkc5xNq/GdNa+1r608Y2Ddxf6Ppqyj+HeFTSMIWWW0vQxL
MYMUZkbapkosEYZ2+p5/SwMRgLoaIoOdMY6n+J9trOIGH2yaHiIRoV5UPAJhU5oroe7obmWF2RbL
ApcZxiSZz+0zwSNvQN6iVMQXXYIqTds7CJHU30nGkeefDql0pm8vAV6k4dWqm8KG70CXtdjc7FGh
gc2dPlGiv7x4Kzt2BPSjyU8AQe0uU2DlvClq4B3nouK61uFqUvYdXA3PJSUyB5UwiDyxsfkTKxHj
+zoX7ouTDlO09hK3JYN2sZHHyJk+r2NqxBwj74CUqet0Tqqubdx5fJ85Zx8ddxZCsHtT8uW5UCd7
D2YJ8wz5wYc8tOVGg6OVHxRHpnGR/I5rdjUAbRLbJGpOp+PyZwmMyYM8fGrmoL1360RbtzY57GNc
JgalKBLwceSFuFXynIF4Xq8khVMiqnKFSKyH1tOt8ntD9BNoXhRCqMyq3z47XP2dfwjYEt1qA2N9
wlWVYETVfoQMP8oSxPi61CUJtEBYcZ9+N1EvN038wGEBXW6Kr2qSKZeW1NvrsDmL3qTr4h30wBWC
QeLbiTwzlEjZhqcyVIqEnwrFR6rzwtx1cgRZjhvFRzqyCbWjPdbUstv0xLLtA5ABMyBSnedP/zqr
pEr/oW4SZCtbGbF9CUZa/eTkKo4Wkzv3yJpUuRX/kOLQYbQh1V3+VHR7lq+wTkaDXWJytHzqtPaF
PVbTqzaZyVQqILxCoxYC8EJ2d0fcoLH13cozIHcUuE+kWD3ssTUIpkiO1NVv3KaUawSLTR6qc3C+
ILWwg00xuR1xr+7IlGQGVXojEdAH379x84/+bcb4Jh7WFCZllTBr/SlrmqtxUJuNUyxF9c1PpjYx
LOW0uvlVnVsvGkkKBxBrvwXFFKOYcW5xDClir9AP5V0dPB2EIe0Op5OHEO6NHHWnKZYxHbaHzvzg
I7KsXaEnCtR506ivmSlPwaWI8ypAhaHk98ipTCshC6fQS67dA4tcd1IsQAQfhU0twdC2YQ9cWQ93
K2DcypdUoAIV9bulEysfYxXXZLqSYUCn7q5LQAUppWbLVzrGLac06xGi3OGGsyQrYhJZtm5CEvun
xRrywF7dH8xRqQk3+Cn/9XqyXfAtrSoz5zJqCUbTP2AUS8v5Ty+mrXFQ6u49vvsZWezZTCtbL/wG
x9KnP0qrccmZiu7V6Bpg9T+RsUpqS5QSFQ6Gtj6iNr3Dd4GXirigoAiAAyNlRye7MQSEhflHNRlt
Gc0P0H95GDHO+o+T/M3Md3q9hoHAkOq+9foEkDgV4nh5ej2RNuPYoF+ds1q/5BSWYKsPuE2WfcUx
ij15tE59QTbIVCWyFWXgiL9GvnprklB1QY5VFQfSALJPArWIdOqamQPkcHkxshOqE+0FRAK0Dsfg
JWUK6F33VjoXC/wfVj6ic39iYdlyC05MdvMVmlcPt75G+i+oFZKIqELA5lWVpQ5hUc5AHY4lOIlI
YtSvgTKuh5aQwTxCV5O1ooSV07nlz2Q=
`protect end_protected

