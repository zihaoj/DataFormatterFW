

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DndfBI7K3jXgN7GHRcECwyAER1W1Qh1PMsFelxk+HDT/ClV9Zo8izeECQIpMvK29OdY6SSkvB4qZ
+AYx/myMTw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CdiSOlcZSDfE8CurfVdELYArX3+TnREZq8E2Yz6CqivQQWiw5RGxv4Gl7Au5kxChzGyLzNLvpmhT
ppQfKBpf+XrJYAfKx28pTmAx8X2waXhIlI0DeX8Ov4RDfCu2fd87Q/1t9q5AVlYHTpz7Pm37oQMC
BonWIfylGOa+liG14eQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gt7F+PGAaFvQvayxMkye/PdntejydD0eqxluJporKL/eE7tO3gqhoJWrHr6EJ2JeFopjz8ez1QhZ
7fAYU5KG/SEWjH1mXWJASfakqz5iOx3/i4t+1xPIK6IS2CWsRDWrz7qcp4f25fwEKkNTRTb0kA3S
z037QRb6Gcl9T23pQbGxiebbA2gHBh4zigT1WwGjqx80nEVyADg7jOuLU2FeqX8nsBo4aya1AaGy
GqejeJaJ5IQ7EY9/zBAWE+DzyhN4Gv8mYP8lGSxa3Sth13PiRU0xsOZGac9yKFHDFVMpCjhoYAJR
tGl0wUk3TSBcSnsYqPGgP97x9w0OHGuDh5JvkA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iuUGkiCJWqD6S+Ivv2+2YU4CYQvzOyv4L6Khf5yoSOlP+8rsrITJxR/snSS95M2cb2SYmzGxjaxu
2TAok7Q+ox5BAM9XQweWOfuwovlgJjHrloEcnxbtYORZwicYwSa91IutF7z8AhDo36QmuOnZx1Z9
NZoQDVYrfJs8Kz0Yenw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
a8x2Lj9mmpL4v+zPKabbpGXEXECaXjvwa8IWoZyGK6gZzcKlusapcFQp2jYobjGuXoqhkYYp4ANR
/7TGF2cuIszd4V+i1ZZL4M5UXTQh9kLT8emsG5cwnR+Nehucye0a/SdOcbn6Pcg7yMce/+zpuuV0
ex4jlZMAsXf6i1il2ddPdtWT3k2AbR+Am3/f8ushp2fsmcGMgRVNtOOYROsCDX4KlRdas9YXlkq5
9d+ubkYzakIVQa0PQ0jQJQPW2/C1fKNsLisKy4kJNaDNwiXo2Ve5N6Qxb5irFP8wZ6iapscbnarw
DNy84LnVZiSVsU3OP8/S7YHAsdW5lukpeuJb8g==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oHWnYLE0J5rZZEnXMuTAQxu9NgUolVXZM5hq9TvCFq0x5b12/jzoW51moxTIzUBj2smQ/sB1QlS7
m2fDrJuFXKoj/HCk0KONHoXlaXmLeXQqL6HYfKw/j2F2fFIBmmAhAJ5qyyPkPnlXCvkE7fsc67s3
qz8a+KKsHGqGWBdeF3lAT6y/10HKSeR6oGugaujjA2CDnjVv5Me6lAzz5C8lRfbolqR+3RNm4o5P
Ra7RJtGQz1ANkLxMLrxpjcw7kXNTLrC08BCVAukRWzPhr9a9wfHitoK0WlXx9s/o5jOgg3Z6WSqF
sJxU74LBWwstEEO17Re4mT3AJPySE6IUwgXMTw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
m/K66vQYu9QA1BLl/gcAAPcw5OmdkIuCmtTZhP5ny0XauLusZmyQq2TTaYJJHp50enFL083AdBGV
cuGBtWI8p19fphHg/q6wQ3Qlnc2VgSHuWSi4yjRVixlUWUBY1q1xdTqZyNyBmMDJe4gu3esu979z
mbfULVfM642BSnFyj8uWkmawV31pTYwf+NgL6T5h/52TsYcQKSY9vvfjzMgLaqPRr7O3yP7UWd9v
wQ0Psq+L0SUg5ymQfK5lGJWKRuOiBQWxSuR2YUK6PlhzNoTUW5Czvc6IhRtlbU9Ld/xHu1RYCXq2
5tmCAPpPTukMzfxtXC10zZj3qecwvU/MAR/w4G4IEJx/TSFliXSZgG4ap8PkWQowOJu9iMBIRSac
seBbh5mj3+f0dZxMIUOmG0sGZoPBGAFqtzRwtuXG1jrb5h0ZEiqIbS3riOqXeVl5ZiCsOUbMF0PY
VF9WYm9aCHRC8JuHfTvTsDybnNUYQgWFGFWQ8TYMQCr9zEhvHQidrfPg7P1eMk/4/UEkuihOIyCY
lnAA4MJgNyd9e8ONr5UulaSgB8vkifeqIfQGFgAT1MtmWuc/98of+6PVL4iWzPwgT59KaAjDrBM0
goKdjVe0YCz9HH1TmVIrJvSZ+4sjHXQgmhDJkud8dTfGO403Vfhz4fqywPDi25AdNhCf4oZKkwRX
D/vGSQv1ODCybrRkI09OwWdaGt3oi7dogv1fADZM1yNrkUeVru9FeyCXMNGHV7Jbm+mHcZa2AJ92
sD4H2HE/lCfMUMnRtmOGpcn6HvvKqAIc+hq1tNF2WN7U12c+bwCmrO62EpbMgsaqfJv8+UMh2vpa
5dHyMjCQSUJ7jARmgT0e2lZGBiLAL9EOTaIABafSGq0L3MzpfjjpoAAIvNJSOGkoKCSvshhoaLGS
kXmGRGMyBvXMgPpldtlzK88DvR1HFhjFR+F2VMuQwQ9oDkB4+vfLCYeTsn/5nwMIk/fXGeI27a+N
F+/tAxmFgqTN2K9GSlG3EZu2/3XMvMHErjs4ZNvFvekK3q69Dd37vgapETyi1B6+8RgVcycAjP62
9mre2q2ZP5ewZpIHq2t4P2ZsytJopMJ7prdOjiQ1e3aoW/pOy3Hz1gqcDKqxt6lSESk4z9YN/ec1
TiPse1Y+8D1Q4QYyzXQviAo3gmAfAHok08c9D+RKSE+qMi1eJ7PIG/ykN+3lY1k03YP922kMRSur
VzL8/MDLwVnz7FwNEBzxbo5f3XDPymtBL7YZMVouXH48AHXug90LBnA/kAah5Qn7PKPAE/JbogQ2
BHEx1iGSp0x/t3rwAlhteBPufW4OuahGe8O0+kExMeBhQsbJgoGjf+Q2hKQh4W+NkvmzLEFODrQT
JmaaPE6jEJbEojOdjMcG8je+skiD6Un/tXELy7/tQpP56Ae1Jw/jtlBkFpR714PAUXlNqFn7YyHB
Pjjuwz979BHYrBmUhN8R0CLkTAHIqE1XrA+fkq5I9/TMGVFO9oJZzI82ds3epuIbqFM4PO0ltbrH
jCI/kUmofJSh4K+r+QtIxZDQeld/cpJxQK4OrcNmz2UeBXsvoeINp5MYk13JXJurNkdbDS/BJNKz
md8Fq511t86fgJOgPJhJ7r1ww9S7C5SN0xYQOpsZLkhe/hz0PpHLelbXaVWFx68UFKk43y/Sbslt
dudT1OwUXjkDIlhr/lP5sJ7nyQpFrHJ7J+FomuW3S3w3kohhTPM0IE68R1f5wAFLHMj254wRMAi6
vRGbv0Tr6ydMIX7/mvVCJEXhri0GkpeRax1phvrsuGweJmcFoME3tIrdhnE0AmKNtzeqDpDA5K84
+npAxR5fTguWsJ/4JS/6P2EHRTQ8xSTEvO5xLk0YUpsBtxnpLpDUDhJ8cjgcjmuV14TQcCK4FRpi
4Mtr32oXaANX7ES59rq7pE81c4My5rc85ryRShRN+svkHgtAU+bBUiqxbYiNSSgObcomLCNp7pbR
vXpIPtbHwz/I6co7kDRnjqRUDxMNSWh21cw0gp0q06//GyHbM7NJEVkZIMKEYfDDz8hJSSBTuCRy
ZUAfEomg83MAT/L4fUQQxrojP6sVMAvQ/sHMz+a0LM4ui7i+lKlh4GZH8nvgzUTgshLA3YHKAvBo
7ZhB0xwxglA/+mffHIgEisV8+REmNGbgx5BKCBH3IShVOuaw062CAC5BVngO7Ag11A+N9vjSOMeY
iyOJqtJMUHyM5TuI7OtfA0KBCvAMZf+DefvWxQlwer6J63RMDgqfkT+KFY00UZOvnLWWNt8xtp9E
YjSgba6wHWIUViCk6Dq++yRbwX6tKa2CssQBSLo7v2XJ0FGiE/hizk1scgKq5tl1QU7f8hC2NMRg
/rorXfAxVWXeMCffppzgo6HGR7qmA1DdtvTepQJ220brcxJTulpan5UZi4naI8IwO7a5lLXAkqUU
iEwzyKGIJN73zBbFthP536bGSTyMajm7znZobuITE/IXxSjbHylM4t4yuCJL/nSdzZegBEeR8IbA
32wwirPQNKH7QNwtAA9XYtk8CtdoO8bUV92GjhDPsrPi+VgfNlUJBd+OB+sicnjwXGjyU9oL6P/7
hXCynR74rLmz8vQgQm/y2ShFNNVdDH2QzDCdebYLXUQppM04JYQ+EzAjjPbe9R5aNaXs5zmpLWEF
ANXcdk6FCjOlXins3D2WB5TAcMmqZnWvR5IzbHTuYZv+cFm753NIf7T6+rLF6P9KJetFXiAei5Y0
fnH0GrDjNdpCAz0OoQq+2IGfb2iM961OXjxn1gVBqnCarIguJjf9EKp3GbuZOzKQiqAtzlOzPj7+
x5U7xk+xe9NmrJYdMKqfHmHpcUF66150FDQrahbq+VONnjjmznGYXaA0mH62BDcL+PUZUxPzL9M4
lc8vfH6WE3lnQqSXD8jRx5HEoD+mLGHCF+42pZsXxxCB1ApgF6mchQMcgt1jF7kkZiVUYmfD5YPP
iBXkXOK1bAiEcqwAlRxJ/Ln+mkJUm+lAe129Zje14VEhR74klTcq/Tp90BWliwg1kzaOQM0TmEcu
lQlt2H98evZYufvbTBivBwC0kLIHLhzQEfwK/gwnhg04ulw2Bpml1Q65K3VeSRA5WpQKoe4CBRPJ
hCE9gk6hgKQEMeKb/l9E12atj4OOdoTF6TxPQvdg8CI+hQyssZ7gTcSKgGblBkdeBUnCTiRw0BxQ
nVrsRgzyfMVW2AGRjZ366ASaa/GfZBEdBkqmQ3fAIL5NcAECnE1CYo/h9I1ErSKaq7vJacse35c6
9bWtFDOHBSWUVSyhB0CBvAmSWu26ahNGOfngBSqnmEDx9a9CrXHp+7wgXICzU+MpavY1t1yvR/m5
500+1WqRDAqgfAD1yYvpyJCZRSX3MdcSJiCh1WXN3BUXzq08MP0fS7KlhE7Du/za3klsVQK2hwKU
0euWAtbsNhGBisf0lB4D59UnCTB5SkFqM57A3nsZ73Wcr3DnNd4ViWCqdVzZNdRKGWOrrTi8Wq/p
fCm15kliZwwrUEHkAx0kkAp96PzWJhGgOkzXkTGtes5hfHYzi41wWWskp8JLQXbABhsyL7KZocVj
xFWWwEEEzf+1MNKtV+z+02lR4h4X5koPENp2EJbr+WCgo8rlIft+rTefj/Qr6XMgNY2nf2ASYolO
LNYdRyKOshrRVabCFmw7rbWzoKMdr+aXsRn7u6voJy1sdBDv8GI3/P+8mQq//WRRj+SLSPrI/uxO
wpz5fMfOVWiUn8tlZgnnCU6cysAQSYsWGhx7FlcQqOKbdMNs46lu/fLtsxtE9REOOCwVjSymp5DF
a4Y3XTNYXMq4kpcfDYzXGvMYFwJgLaVW6vwWkmsj4a8VpxkgcxzicF2DUT3GdybF4uGrr9JlAe7q
4P7R5JtJscmLBoWLcfczG61i3XSSWkXtS0BIGQnpCRlLdx7MOIA6ftXbufT5045btiIFNV4uJ3Do
DLViEUhY6zglp9TbMypDA3zZLBWEhZlaVKNX8P3K7TwfQo2n7c8Lebh+ntjvgf/yvPgYjCXdys56
ZN0uehs7mqIEuXolnzDbdh/j6RAJn/9BrERySOZPmS6teISWnJL3UYPB9apjsM/aCt6MpVW7n7Wi
sWCtOOFABW1/2sFzi3qI0sCP0frJozqS/9EyRGYTcuqMC+MNZRvJ9JRj306xGLhtzk2m8Ue2iQWm
qE1wdSVObrepr1YIVAZJsY5Yr2aWvGsaOWrURdlpeUjDniR7Hg/pg6hJdAWXxR4Y0UdReJbnlA8Z
tBOluw+zXYbAjgTFo+h/k+Cg4ilVC53g1iu8jziDuyEoTai36zss3AGUdOG29l43jrGzAs6aGu7W
keevMgnbsY6ziJ+G6W4zBSDuuPdpvQcAOn5vNnvAbzYB/GDbZWHU4mR5VDMg/HY6fcjYmIcX2Z0q
uvEIFElRVWaM0eUBUVbTHHMM0AaypspW1uORr7LvGukXUL7CGGpR0qCgrgLRG6a6ffbIvNqXWr08
5Ly09IwRpRoOLnc0yd8YLTiAfERJ+ps7c4ybDZEEnXphnMyFSW+gIl9nvixgsymhCwYpBWX/T6Yd
depi6cLXZrEYNiyxny9JFEA75Kb1Coe6wXdcU22T+7Ziqd9NGY+1pMhjPl1jyN6NobL1lkE/loAq
ktK/KVDJQ5ss3Mh/TKg0oG9fNWx+WxBVfSRDaF1g2hLqHK3hwjqE6XVYMtiD4BhhJACXWrjbDQ3Z
vTDDCPirUdnIiDEM+ov2eHdRdhYH8OnP8/vuUw5ulkRLQ8k5bMBdE5b84EltryxRx+jnNN2i3jVP
rnLAPhi5tY0YiVBnbhS/BWA17+/X2gWugu8tMw9mi3HVHkKUrBw552I9Lnn9XpWMhL4irHXQbBSR
1z/Uut+fGLS6Z4P6cq2js2FXJvy7F9psHc36k4btq3hRvuqrqLxIOCJS4ShFXntKIui5VSmd0tu0
S6q/vlF/5cvf7jmPS3aGdMjiuPV57bmAjADgOqMk7hDwt7hq00aRZXHvQnhdj0gnH0bg/WqS/6jI
pZv/SyTttPRO3pvRweaqYGQkbh5mQ+vONn2IhGUV/mKPuD3v12lV6bwMtXyrElSTWOJFPpYWg8Hs
IGdR7NL+wV63Y7adrJXt+YRRKpO1F29oPzNFEnnCvY0zmvhNxJEO9sHcV2v5kbswctigwjl6hkGW
OD6jgrBUnsfzrbpmzhbqNcKXa8lUw50xe4EeLYc6IM9tISYeEOPt1VepyvgdGLt+6xePRDj8/bcN
t1i9/eh42pUF7sQtCHxrxwvJ8CZOgx0KQkoaXk70esJoDs81YLl7AmCtu0UfgUoxhyndbSjiQXTs
bvLypzia6SG1MzHJdS+FFDGkXweWGhlttKKauv/NasYy4As+GOM32+DjTVv4cWZAsfXim3Xehoi5
nzJzxr6OMKGvxFI6AVWcYxj7sVgcsonivpfdqV/f6RSXPlu7hBodfE2xQFvczvZIuXSqbc5wT9wv
e8jhBrA6mSwRGyk74/5C9nbsJNUcFGeU8Chu6jO2dijpIGXBJ3mxOZfIUi45MoDHQG/2ZeaMaw8q
MtQOvwnIRX9dzks6ARVHFSuyRKu6j/5YaTL9dbRsv3Ft/1qlCR5GhYGZhmNgcERCgDkLcTZkDFWn
n9GIbAQSE5uPVpfikGTPghsFdmoIt2AFu0JzEHV7flNrl2nEFoDTcRXiQHoQvEZ5lhTybuDWkAW2
d+4W6wza/f/mwXSLUePgcPf1mv0N619iPEe25kRr+6o2HrBzzUfcjXp/IOuFaU+eg080eCXWsOVU
wtdWXb1TvVCp2CIFz/30LgDCp1/q7E8yS9CmsCdXaEW4ZKIJeFwo2g32AVV3oyE4F7eVs+TTkw7C
OgdaPTjmJLPsi3IMRVVWs3F9G5GySbwTxzu+lMrhoFtBVuNPpXE2mrk0O5hUVw87Oqdp+VNI0b3/
zt3hkmmCmkUix05dFhQXMVWRAK0hYR7o4q7CfSl3Df+rcW5gACGcoLt+wucCS5KzPnmpRmLyBQvy
AlAQMdij+8z1BEJj0YdLZv4qWyoo0LURf6uv1dAZjAYLkiObGZUZ8XeVp6pEUiT1m2BnAOW+XAE+
KLaHMlwF9jiM1ZRMZ4KOqS6RrCuUS+PwmVaPjc8AHOzRQmP359DmMmIMEyCiPLXyFjcR23T9yj0w
2NqgRs1mTVZdNcsrd/95FBPtw4gWNtp08cLIKz0axQ0rCynT65QhGp2eMyYts37rE0aDIqvOAqNT
coIo+G4tRTzuzeqUxhOLjo8KLShiCwwxDHLeOwH86RbRiiwk5fJpxqxPdztCPcaoe8q4ZlfMMcIO
p6/bPnU29CKydaVHPQ/6ILwQ+P6TT9O0nEIcFb89R9RCfIuTmgG2AsjhK0n+fwehsGH8tdGQg+gS
9yFE6kyxbpKOvNK5s7UY77l2YqQ9M7NVo1NYUmKNWCkDj/ewTQmrSqrb7rtyilVUfA3xx/VUGLkR
g+DzocS5vn4E0eJkFcF40bWUGBuJQvH8fAhdyH+5hKSwIWtuMX4MpCgmY9E3c3Ia5Y2uXDqKKimE
LHD2fOqoa473gzwtg1ybJaXKJlawbi+CC9lJmpxmAKUuRpz7s3QyVir4nCTUGmVCbwDahSJW8WUf
4RGZxTZ73Po9AnkOBC+ruo0RMp8kwC6tpJC0TKKkWBReARejtEKH53ZYU4HznMLZpkfgqKGqbi+Z
DLu9/Yxl4w9ROElGPp+gr3FiNTshcN1dgF80CwKBGq+akmhfzahZvPVL9yW5dFfGMYnIRwPDyVsw
eijqz3Wgo1Dq3+H0UuBMRPcN2K5gdZ6l6Yb7I/Cguug1N1IEMjpUSi7wkXMzbtxEJnt7t5QoEmSD
a1MHhXDnU+vk5r5hsyF8KIjqukteY1Wm7c9imIC5bYJV6tCZF851COwXCgrQIRR82Llu1iwGkWuV
7jGYmbDgtcLer/1cFLaFrw3ncoqntKEHXXoD6CcEb3T6182j3GtN78+HbK0PC6gBe85UTSdutNMB
PV+QLFAZyeArXl+tuA0yMSewkVo+DFElUCX7qW/UG7xWR3r04IMDks14EVfnDsKOk80gPAEYpInP
7PmlXHGka/noVjg=
`protect end_protected

