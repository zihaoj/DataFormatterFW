

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
O2XOryoxWHSJpVHdyGBaJQNdc8dOymHDuiuAfQsjyy00yg+Fygx/oSQcLoNz20CMTJ0oXsfO0N0b
OcuaV/bA7w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GVuiQASL5MnoVfjBYAuifaKQBYP5qpKi94ZTFg3hPhVSV5Z3K+xBNk7HSc26fljddtOPeyiQrh28
UfOI+r/9r3w7ch+EIVITv736T0H00tqEtDgqpJcf40ZaJFg7/DAJqa4bfrwQYMPPMtN/+LWpquNE
dRSjfIReTFFkjcqBuxk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kP3f3BnKcYzaKjuqBtrZmy5+UEIJ4O5AkfCZWz9sAHrlVU+4nM1IBXUAwmiC3k5d0krwcI3sEm4r
vt+G6kIqnFjoTn4NiQbiqvWYDmZzV+LJflhoMqNrJkRkcVVp61x4JZUlEr7e9p00rvVMbcTDW6Kw
nnCwqMLBkzM5UVDhuEC2tdG2CpSgECEGlLMMTk0DSKezGNtQXz+KtY6h+PnOfx+PFZwhFOBl/jB2
jTMtcKAeD4gg4WKoAn+7IIlgw2/HhJB3KvzLJpLw91PETbk4sabjQbQ8KStQpjvFK782EG+wfv9+
81MDogRQiFyFmN6oxg8ELCZnY8O9CQoxYornjA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
u1fw90y9ARra+4xSQeglVz70mgNc2urrAekaZxIT13N7fl3y5c7IkQ5+gaCLFemZ6U1NIJElw95Y
NB/VTj4qfRZU4t2hFTedbkAP9HTfBoQLkd5eok5logHyANc3ZiAYnVdPL08Ys63j5F1wjpsesyup
0l3zS8O13B+I+gzKcFc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tgz+QXmbbEHiuFJzeRhVhbQJi9JNitJrdU91eD4OUl255UhEJMjfDaR/UN2Kmj3daj1Y6N9XoIi4
93BpVsNATisoDDeAvL/Rji5I3h7VXyiH5+MTk/s7Sj/KtzXNgKZlWFjJ3fcXqt8NLD6Juh3fnX54
GPDGKSPlW9MCzzT1JtDTr124bXptK/drTliCAmE7pdznkO5CQgRoDuEMokxTyMyOhM68hW0orIve
hBJnTlVs0V8aXizs6E2X9cL1ipD/zg1cmKwssQsXb4Jo38wsiBwFRI72/29AenPb8DiuBit8capG
ogUYTJYZPuHqoOjMDVs+8SZ9yLvbdyM/mPqYbQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9wfRxLjHUbwfTCjVdZcUlkVYIcSGOY5nHZELBaw1c/NDgsx5AflnXGqVw4ZcJVPhssJ8DFS/Hc0
BI96JG0oHrBsT0vEMRXoqAsIx9uiqFlhRbqlIF+e7F7IeBTdC6YXEXctyyXaAZNLmebzM3iZjvNh
ALtVke4lfkxz04zLYQv0C6ISqIwI+PlZWuqgIkOTgdWEtdxW+zW57JrC//OTuGggYGgTTtrpZN+D
56aBhSpOLY6ft3tCy/T96Rbxc23Ol2kCLBG7e8/nHNSSDpF2k+L4dRyTkMYFBNGDcszGyu7cghxU
TRsP90Nwu4h9+YZrBGgV81oXDRYKcIAKdTl2zQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4784)
`protect data_block
oJeKqDGNiBYjPNbC+BXEn3GFQsm5jh/B4C0gQFI+sQ16L0vTb4w0QuCd2Cnh4desP05KDnk7GEJn
SnNsElht4Z7xEnm+ArqS2fSqw4FwNP8sn8fkL5iUBwhWZQMh5rmAxpTu2mLLQKLl77TQjOke28ap
0zDdzE7+rAg+mOdgMou8FXwjCUQ/s/zaFfkJshZBARzmaSL651vwV4onrfBsnCinn9rESP9szstc
1F77WcukJcukQkAHWDLY/J/TqAvCB70LaQIMM5W2NTXOIX4abFR6noLfou6gzFcsCprXuR9OwHgr
TFP5AsTdUKWHp1TXGsPerNE6/nlIrwNx2SoPwInUXgIOZlRnZH5RvuLI9Fd77m5+TlTNn+oO1E0z
Z1wPK5kD4n14Od89z1iIuTOus9/DbowTLITEnZK/qVJ3gQrAycUCfdv/SiwSNHWVpk6dadTNLA5b
+fZMsQFkJw8Tp6QryNpbuS0YyLQGLSJIIR7IQxUSSm1RfcMXRz4PdzrazztwypCDgoP64Y43GiyB
M8uNb/SxH7f8/ogk8cLU9yKlwiOqOBN21uuNh8nw0A332Cl/W413/NTfF1RZ7oRU280J6lAUNMfm
Nwf9ELSYD9L6ZT1+Bus3DkqYM2TwBzCMhBzFtEIED+/GkpvehfrR1xBeJJ5dy7FF8a4UgDj+0xAN
aHlpL4ZtRGIEQWMC8C1qKyHetCc2Z2Lu9+b9c4sDjbIkBZHZRbSZUQMzFcCCCUz4l41lbhQVIVDM
1aLKZbgiq5SnbzcMEz6k2jHeN+WfxXbQewSzgLENVS7mXPmkLV57J2gdCnrmpIxi2jifFZvgoDEJ
bq5gqfjMx0KQmF6FR0pyKBNiFvuCRJ5ezzoGQsFGxb5U556sUwyU7Pn9XZJV7nOVhNuy3gEDAPBF
Fq1x6DxmQ1Z8OIuGKy4L914Mjg6wYby0vbDvBrF5Ew3XG7u6xRGwfU/PDTaOCsy0F7WKbZuFHBLC
7btKWII3E5xQF89XBnFwwU6GXvmN6gWu0y2/SBHL01kQNUrTCKZlz0RAr9emfJJGIF/S+2Fqmrpz
NK3fupeCtUEbBawk1eIBV/idZORhTnj56rHy/h7wzxrJ4Oo4JmWd3eeUN5KUxVZ110Ge+ev2Sflh
gbro/Tz+NuLzBvlmsU3W0X00nHcEOTi200EQGggQ1Yfl2yGDJUx8MUxijxJ9q7ryeiJqpdlZG2mK
9NZzFwmqPhj5VuyaeXbc59LQq2ZuZ+RK9166ON12u3/btcJWejFMNqXVJvw0hlE6XTN2qUf2P46x
joA/QoTZzZ+R2SGEUdCuFrDDByRPkWgqfvstnnne9X/zcV8pdXM9DMkFdj2JZMG91NQz4O5UwoWw
0RRii69aSoIaGC6ZjwNMLqKJ66yhzFy5u2eOp+ed7+Ps5Vb0qFUwqi5mSgpW9NlWv2zW4gQ3KF59
O7SJ1vQGWOvtazcB/5Io/NByT/U68mLCaDAebM5ZgbKJqFfvkewI9u1tU4n9Bany1v13j6utOWbK
ozDWFTy4gtqt15ueNns5FjsouvYZsOFoI7RnJ8kyc6nze2v+BEHcx96iQdBODvR2riYMvIHPQ01H
7yJJB0eoFNAYe8NkTSVaRRu17zzGExL5ckVHLFNEBpxh5YgchDitdte8OyRmJqdrpYAXcQgowkTn
nYST58yxsEonAjn+Eeefgzpt9ZnzDcFwv7FHJOvrlxKoO9EGoMQyzw/typZA8jR566I8cuMpaNEg
UaDvNZnkSVwLdUajVpO+ji03QjjqHytZexGI8VSg+wj0k19st9QlU0/FEkPb5iRpU6ua+bE2WnCO
2nRvirpazHGt6JcbReskCifh6dlsoh+wQVj9vbbNKpmAh7gWtWJpaWMiVAkFBAbkG2WihCa2+QAB
jTz8RT+98sJqRbISpQaqv7PmGakE/gQuVlAmmOKH9mGl+PUW1+RdHRZycycj6he16u7/Nouaify3
GAtrgoEos7HBxbhsM4ojD4XHfSxv9mDINrPH15upam5dEC1CEw6L19Zoc8vQ2NiRlaDEIAQGwzex
f3UVvCRkGl23mZ6BfMSy2k0A2FnjryoPejCBsmxjFAE5IM+IaJvczI9gNwSTW38pga8YQXCF/Cen
Jojdz760vxtyZxwMX0W49n3YQUHMhCAa9swUHuzp1KaCj/V6DGzd7jf62i2n6NFpynNJA67YQ3oL
lxxyFbpoHrr0en5YFjg3Bs8iUmVIbB2NpBwEpozFwGVmINLyT2/bZObshjc0josBbsQ4JutNUnXW
6lq4I6vA4ODd1CfWNYKNTPI8FZpoYVCUQy7hO6MyQq4p37QfpsH7kLDK7HEJ5pEcjxbsaV3xKHFi
PKUXI9FJ7FoRd8rOzcY2pbhhgE/Cy7Up6Paox99TqYXa+RgV8a7Q+AdIgdBUbew8Lr+DrNCiz9XG
5kAvcoBFae4Ugq+NpzgsWfYTdGnX2TnzmqOFU98UPg1XSk3PJAur5YjOnAMayQWSWMCyQkKBXef1
gW5a583M5DV5IuApkiEmSrMJ4RI6HA7GIZonzn4giS7RACU2yp1tpAx5iJlN2CnfIi7rXh0DWxzf
T86740hYp4bxcPzUj19q2akmoq95w4Se3roKmaEGFGC3kufkJiGpU6eiMp5sUd/TUugRZyVPCQlS
6Hgy7ZiZ6HvtgU6iI7/grfZwkA/XfDocr9eJnzROe32DhnWaoJi3xyFJpuyNjjx5XDEuc5tToiPz
PoB5eRLZFzHJFyyBrtbIK5aqwJoxP6c5+88bys64dvdyEaW1ciQ0PHKEC0Z9AVf+kQtTxWa7Lp6j
Sq9mZ4uKWL6OeMyb+uycXX4yBY/AXSS+3+zn+p2OOa5QBGKeGiRklwBxNj5hImFs+fnTA05Ph784
LrIzkkUPimLTaSSjeiGyFp0kmrlW26WXj7Kgey8Qyu25ZXBS1/KTEgK5Zmz5SLYlPIkKmpudEr/7
v8pgFt4WIL2nDe302YSHZI8ZaYVD29HOnpa3ukse+S/dPO6jj3GOjDCPi20aoG47h9kHGzeI6fIi
XozGKaJwY6yCRYavUZKJ2bZvQ9Fys/kr24UJdeKEEPdKrIqOz9a6Jyeo296MuKze3DAZqWmC+zbv
1u1+Aiszd2NRdxd7h7PDxWNZgtShjxnwxuT4sXS60ONItZiof+HuRYDemJ+ZDVduegXdW7s5VQkB
JGRwOEI8nAV1UwMyKaXH3iGe2DVXgb5dXh3Phj1g/P9+r+UfCJ3PtkwpEPlBdXu0Sa5VtmMPb3zO
Oi8KRWiWJ/0Yd2JckO95bHB1n/06fxB5lVttrr6qpPMqXyYWaoSZtvmK4D6SeBi7hQSr7r7Yl4ye
ikhXFRXgk9LKUmDFpz0Dq4wHfIbTwZE1+lE1CXpUIoJTNWnCo5BHqKrECTylh3VG3plDRHf+YL4P
qOs7NVJ2h0gMGdFI/E9Pe1qzPFnxpZolSjmAStAuZynGRa8jBljVpXDvfdBZN89Kop8nXJLmMqYf
mse0S22pwSPwBpUVv0hDgHmXcP3toHoYyGwirsP7R/yzOOGkXEKSb9TgKZexzq0xaw16DMr/Axq4
odmlE/JcKdsj/qP0guZKWDiYOQvd5NQs4M7CgaOkPK1KqH7/W4oaqdm85PBIkJQ/1RdS5vp/LJFf
Tmnei9DwT3yRWZW9o1wX5uDL7RJqnAaclpbRqxfipjpuY68TMNqPPep46hZ3t1CFNSioPNhJrWNS
S0UAMbrC8lNmVi9MlDkXg2VSqZOF7YtFFbedcXQsyOlnfUTE+DizzumRQOGwzXf1+dxOTdpKnzyZ
xQsGWlXJQN3Vxx0mH5mhWRyCCdEYb6E55j0zPyIcXUTyiOR+kLQVIFloZI6bmwzEzlfJTmZyp4uv
Gx0i5YJKTBQxRR5v9nB6ULddz72I4PYnHzDP+kTziGS9E+P8HTqPk5wVDK6ebsOZEMW1a3q5z9Or
GwguVyzG5dNevHr5HhvLfRCcP98Rg1Cwy8rMQ2WLMWMz5ESfNmnrgYJjf1N4nGmL9OaV1o74Bibp
5IrHDiojmqKepQUO6nytaBtw0XNPvIudEeuC5QoGuGPKMawj29FIonfKC+C4lb3AZvk8iWpEZnNg
PnHX3EcAl9ulqZ0w22z26jqxcG/U2H+aETBUt0tsxxjys71sWWBwmTfC1coYdG3YqQoZadFdwcqf
QF9E3yHiE8SFKXBB2hxuX76jcNWnM8IT8UjrK/RP1eP6YgF1CIdCDC4/uKnpXryN7N0kho4Ha4VQ
qT1w9yfwUA6A1xRME8DFNy+BC7y/MUJRxdHmb8ZHSrIC1NtGkeqwrZljiDYGDRMzpOCX4widshyb
QjOndnYuVskJTcrHg86IuGRIgJNNxcpZ8Sf9c7f6VBQpvrETLBW9DxDVLF/9qhz5TqgiUtPaQJmo
vzajdmo8/JpDQ2AGzQDZ/OsYOaGqBje+rysY9UUydWHTUQaCTCm0s6IEfxIgKHGFeRdzs5JIUOQs
xoRHNThbmftpIGZBZgNih9HWDVUMvZyqnVsWMdbmpW6sJzNvltPBZzMBHayJpiWQbaYJ/bOG4jP6
CKinV2/yhh2mElUc7jJO53aEISf/qt5n8mxox6fycf51wbbN6ZturgBHf7iYsg3r0B9TnaWbEYC/
YjFCVtLyCq9yupk+PH3hCV4y3XueU7HihnevWy7CMI/K72wf4Ly6BVZYT1vx7KrFPv9+UPyHmtBS
xMcownHBJV9UTSIGCqrR19M/wFXpmXcxyaI+hkEI9c5SHtJwvuz3AagUHsQdsYXeVwJhJXIn8XzF
8AuEcSR2M6WZpnRzJ40MIZXS2+oPfqKDevCydzXeu1WjgxSWw8xLwbn30pbR9BW5FLucUIo0FxM5
1mukbcomVzZlwK+pwJpZLCGoD0TFjKj7heWqaXs/0XhWubWGBTnraN10628VKqFv/o6vUqoSajQk
uzHvTlomquf9pUTIoDoEXiP+MxdeSNOrzTa8jxKQ2nqNVot0O6Vmu2mZgrCmhotga5pL9yDR9020
UAoORso0ggS768q6Lq6VaVYOOHtQqYS9ovf6AlgVwNi59/aqS8geQlPF1KqRUXx3lH6hdgMKbmEH
VXpAaaDpo+SMuOy5rjBx/5ZLF5bsr82g2+98+JRVy9AIDAyC6Hzon781HXQuMIqZW1zoRYWCtfNd
ZLc7uN+ay16clGP8TWTnlVrlxYR/iyfghluBlklEYQACXw5ij8W5EdYKnxY9WFTYk7Gitz3kw2dx
f0D5iYylWJL+hr7g+FM6MJQAoJY5WMP0OEE0shEjrBXTOiWTpuNBy8pnCdV2GELrMpovfd97jnng
YIfu7YgcDRH8eb9RAg2hYsWnmSr/TxBYjZVvQBIwmhTbZZqcgLkInOkUF3Hw0AUyhf9RBC5KxU99
gfd0RqE9fD1OUkMpMokfdfIJmo3KnlvqvrGDof6CgsoVgF3su9K3WwUtTlTGfI/qbBFq0j6rYFeh
Fo+SGFr9rN4xGVIV3SriGuFkuJDeFmrju/OJ8kUlM5NQ2PAeh805+cN8bP5vNAJFaK+jUtj93LUp
F47B4wYq0keib9J16DiSf4N0K7Lwgl5TVu3pRRRb/6Jgq+ip0R0fc/miYjn258sEH364OKPfXnx6
wDGj9XO7n8Yv1anFKMAwhDza0EISRhHNKNkmra5+kPxx8vQ7Hx9yt5C/aNmIicmz4nw0ZBnrBOmK
aZDfOCkfYe0GK6z0CPXKCUPyXf7LPSbJLonsYkd07DVa4fxKgg5YwStbllCoCx16eHIZrcdrK178
uXmmMz6F1Tdi+kXYvTXK1jgNPHGA1TshskHHg/aAaGC3kQgeUbBb7TnBtjWEH4pO8e7GcZpKmu34
JgcaBvwTvXRaVZ1GOiYB3qmnGvfm2pGFcFq1Tr+6a07SO37e7dvPzBlI2eoXfeYk+RVkDFPhZVbA
fQnqejPSAQEHToSS/jKFaNQfKM1jgm+12R3xPWqzRYlq2GYddnXuQyl76A1rgtE7tfpJr283+x32
isoGLFYpLG0O3FjGHhY9G5KhQRlroM+Snl8RoELc3/XTbvHiG/bGbArQtqe8UopToqkJLxBkhnvo
nlJfqGdJTRRso8XGnzDdfjz2nUesplhb2UD8JGpcIPyeqqTw8vhn0wLfAx8l3qguePW75Pp8MjdE
cYBYH1oZlEscvXV66940fenCFeva4lZKkGswu5dERSqSmH+i/UryjVilnqEBpUC19cyUXHMhCnP7
j8zYY/1E015V/xvKGNtVCd2SSClKpQFBR3O3Ien8NUNq35CLO5QHh920+IeeCCqNmXMH9t0RRutO
vM2keNbptRWkRqKWf/mmngCs6pdRibGEmaXlfhlPcI3aHDRUEYrPLHOzYkkSvVT9lWeBpW0=
`protect end_protected

