

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
F7epTRDP+ATLdtqtc2nC2OSZczGx67L64fpl++a7vO0NSC8K2cMxcWhGCXTuSyruiKkI52pC0FWi
92USfenllA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZsiqUgXk28+FPYFbU84A9fvO2iyXFjc0w07TvmIwxayLYCVtgv9t1adbrr6AaWzUmo3xaSIj6eCk
8rm+ZDLPzYTB/jH/1iWDWQzLame2Gf9aRTNr86ypFcAb6rfUFHnWvxFiJRW+Y5pHL0QNq7m4YRr2
vI0X1oFIhf3mcdGnXLs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JvA3K8ql3Q6rhslV1z6HgDs1h5pfPDtPPCkAbKIxdLTkYl9A9jKaKmHnv0pWsZuRjE58tjmEmw77
1gS34IhfrxmJwWaKxLYOZC6ux2UZkJazTZ9u8pKgEp30O3v2mBmEipvUZ4YW0M3GSfQsD51a7gFB
81hLGFgshyi2sg0oMUz0V/K92iDusX9rLgHCMP4Pt9VoHoW3DcMvTwKqtLbLcEwqF8IIbruKRMHr
4fq8Xhjk0YMZa0faXAeO76z+KU0//gF7PXOmgDYJHlPqO+/mLvLI5zX//CZzWCNJoxw8y74pmWCk
U+kzgiVU18Te5Vo8L6H7fo3bQLAb+c+zHQNPMA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Nh1ETOQwBM4Ffqo4RPRwCVBqUPEYVk5ZWX6kJzP6bReiD5QOtE+DxmVrcoba5SvXOP9Qd4ratu8y
FcnoIN1ham5QuhZX+86RHkJISdhv1rdmTCROj02Fqyj4w2r9z+hBynPJkHFdqCJ7h9dq2Tr0Htga
UTl8YN7DWZasu1O9/y8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gt1D1fJqX4gbwd6T54QIz+e8PpMNQxpsFDicvP4VA5Lkj1S+RqS4TAeTTq1eN1DHhXXHpB96WZER
daGiqWoEx0b5J/lH4/YdZ2xZQE/EG0+ix8ikLhMe566K9ZtBE4SF+FXL8NaOItARJNvNnAsofd3v
mJMleeqXC+Ieudo54/bPv2b4LBskGDPrZIR+V79Jpm7+c+N5pcyu2jEI1QJs9f5P/l0JdSdtG8XD
Qw9vz3OysCIcZAzQ3CcAyYKcm1B9o7nKtRW3nt7BXNpOTpBQCeHAjteNn7EAPz6H1kKqZChvv1p1
s0t7mduDI3pauCmDopGG2XWCSkr2tjKr+kVHZg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5312)
`protect data_block
LAj8MyZEu6T1bxFaH4NfqtbEjGngjQ2P5kKdL09u/zEsLNMs0rdDSSAlbJ54cmmlHuhYAODlNFIk
DieuIbCO075MFzrpYJ5RmhARr7poqqa/dPs+1N5WFqxI/ynIRvzuoOy3RjmmcAohIQl3sEk2BCV3
JPaBj8lEtL8yttAH30tVc3capa6OP8qtzivDy9pMSoTeMhqGwNcji5pSBX6NlpXDselFl+ZX6VRK
zt0qrg4BnXWdyXoLNf96/vvmb2+yRL3ylW3hsbWBGI/izfGFJb/IGqqvrjxJzSyLrSRGdZGr9+LA
fofczqFqRfdpHb3wMlJfYNHHbUl/v8YRsDw8h65hCeVuoA40wYZcC3HVZqkM1NQbZiFK8CF5+jt6
5Lrg3cApgIB9vIXFAkLUgj06TAFztc9/KQoq91l5EOvRr/qMjYwo5l0tyD1lRtLoxDaUphKTxhsg
9reNmKmHiAkm6LDzJt5v/HbbpqbD46587ssiOD+QSe5/1TncFgbV2lbGF7bB2kaN2826kUKY3Djq
tDuhipHBj2UKjyVUuFLnJlR5UI9pDI8Rzun+QBJ7CHaCa0nv5yT9tRQEE3w0G/Epy6V6O0WKjull
VmEfm9odmHytsgNxOhlwqBnHIIqOPcsxAZ1VR5lOW1erG57mAXoqy3DAvx1HaLNMrmPp789ghans
E+UbNC8/APrSM8SDUtaAIZwCzxBatPPduaQWZuKF+9jZXkuPfAyLHCdrNxolyAxRTb1oZU65JAHa
qfXOWu/Rk2PboyTZ+LyqSG3BriafYLaEltwWIuu0TQ/FTaBPXHSTSyHLp5DmrRwAzfhJ/EDDFyMS
kdnqqkIfhxU2WTl3OHPdBWNV9hwcsVjaEuJrmJQHei2ZeOts60AYIv5AG527Z7uDyNEo+ei6nycv
jHO9cCKBZDsRj2/VHwl+oO9lXyW2wp0Qx7jZ+hjEcB8xCA+zbGFG57BJUtyYdUxlj6xgn9JolaBA
oe/TT70r+usDLVayO0H4b0rVZBtrYaexAATWidoFYdk2YOMJ1dBbLfEVTtcbtOzw0AWJ5LulZ3wr
F506g+s263D3dYnblsXk72XP+3+FwL+HNQqHJCQBsNHhKU42K0HeHjAd226HfntGQDnDdX/wgVeG
CTxHv9O/iGzcxxO9PUZ31Wa644yUaRzkyVfXzzPKFiC1REgqNSiLDXuZYfvxNEK7dIubKsA1IxgN
1OqOCLc7vlji6jbJ7QmhcYA531vtiEN1tDptPOOvvwS+r/plICWXTo79VJxUq+dYuH2giQaJFsKz
vU1ry5L+15klUvY51zt+Kjv/baxMjGwZJKtjudYjOx4HRDtravxMa3V/8Z3oE4yyqYSeTSAxNmTP
rZQCMcybRA6w9AV7eiYlIgM13e4YjvXAF+TRIVv3E8pgQx0G/cVyov3tEVTsseqT8EdxNuYEb5Xh
GKF+HKXXRyapmUxKP0O3unAKaBoKquqjBctvvnAu4osU1ErLN7xVp9bwMg6nl33tiks1LtOFBK7N
rIEw3we5h/5eza+7AV76wy+7LHN++vC45PsEB4Htnth2hckI7Yt72kulDyEPBSIRjKQJi3vohyO8
YPysS3d3wbCpmCw5fSuIKUpwYhKB0vtkdiQXi9IaNeJz+oERCZQRYMSGlgvaSHDGouSzTuKeobpB
xLvViP3GMKNbuTTsXeqcACAH74AmURcggBJOxWR/2yKu6WuRD04FedYTKt98Mpm+sdsx71kqNPZe
Wr03QofRaHkXJUsddatUq2fci5iGOiALWktDkY69iGpVc4+79UwgQNanMcyikVuTTS162cl2bfhR
2UbQerwxIj0HPKYP69TeIEDdJjUD+DWjCrxvn+GZRl20u9dH2kxVCxUdjKiAuhEs34OyRbHU9Ayt
EzWt9JfWPkwS5CDvZVEaeMD6qIUZQiRoPuot7t5ouOXCQQesm0bZQ7Dsf9k6O5j07cJubYkPS1Dp
pxP8yEwb+rBImWTpzTR2bp3G4OQyXXXq+foCFiIteGxjxHgXeO9b8fCJcsghXfgcC4YkDBTxy3H7
NisBnQtqtNyx9V7QhKJrUgGf4GkrosOW3pot7lR9l+SiYOuCEnU6vdRDkOy1V+HODwMNYSM83wwL
KlyZMBl6+5DhFSoptVxU7hzE3vbELifGF9MnLchj7h39MaJyFZ90mvCkZZfqhd7dtmA2GvyQCx2x
TYEvf7UAGxtIFUgCOOL41fqszZIRMsXp55WHFG0xUunCS0zRwuopXTkR0/5ZhU0Fo5W/kHncdGiq
AhHs6Gg3/hYL2KMqiqebiEt50mIR9UngugmDxesjv3Vf+WYyBwLmAgQeXFe+PwUY7h+i05smJy64
r7z3izFp8Gcv5xDux02W1h90WaIwB0wahr9DcYigkKT3Xja1I6Tcsx6b1Yw8tesgBdNYLxIrdV2K
U597QEXJEI9RnuR7KvBV5u6C+j5tnVwxlLpQci0npYtvKEgzQManaQuBDWgiGsmDNClrJyH3POT4
RUSnSKaT7lSoNH722W9KvYmyOk7zrjHURVmtY7E6IJDZm4qNNlYgeOeHCFkr6Zb9DL+1mgsHOxdS
kdEURYHo0kFXPLAQfuRrebsfS7pi05Wifp8U9Qk0JnjhLf6gqNyqKgp8j4Tn3o+jJ98Dcs5eZ9Vh
R0K0b8QfcHP+d8mZK4YNhyuA68O8F793rwc8XifQFar65MKBo62g+g/CDhfFqkZoZH4VfKH56jsM
R6VSORyMyiQSHhONdyL6GgshK/xvAlaI9q3mw1pLzg4eL/gudVFAPKQGTKxWpYZE0CB1it9H/DKl
CkzHfD2xFFR8feDa78LA7g4q1ncmMIX/1amNEYgX7iWDwRNUxEWubT/XivyqT5cOIKFwdKMoSGaV
LDNx9GxUYpZv92irbPL12Orirv/yC4+HojA2qSMj3HbKj2HGdJ2cTVmrCcc5cpN5MKs0uFYcpfNN
vPKrVWreJU6o5XmgS90NvYKTGup5kH2sTtGmd0tm7ebizerHEFuWuQl4HNzN2WVuZtDjJDxwV9at
wkuZdCVSuYa4ZGij4o8qs/PVz4LZ4K6Fy1WxDZevB/IvFXhm5bcHj3X1s4tL+EIRzRAGUCesyBFq
M8GcubM18ZYowjWogx1Zigg737vM6M2a89rEk49BcWSw65UHe2GJt/t0mb2QTdjzSfSei9ZGpocZ
AWpIF4t0U4taYgiRDLMBH26NBPEBDjUk23fWrumyu9aAl3931rdDNCTpWtqYBfBLKefC+6KbGbns
C4p0MAX3Qi4Wh6SZBnLLtke1t6Vvf8a3MLaJxSObaoBpbraY5qL8ZAxlCHNGztqv4t0kPTZAgX0X
2+J+IAFjrWJKZ/f+i0hq+xVmwpaNN8HPZ6srSuAkwfravfbxmxxXaP4MAZ0OOehrjmX001Zy3384
4e0Eq8frf5LMPD4B6P5cRkLWU7Oazzp2gYGzGBZEFKtrovkL826mGjJv5gIe69opWbM4zl3IXZpg
BvsyeJpMl3T2nI6bxbhNdzt06cnzC3bA4jFNcxNlYEpf2RAQVO/fRWWlfccDMtoBW3RPuPFUc6vr
rYBktUlR3MxZig74wReocBtZpmWmA+scXU6tC5vEiM7S5pPbMC6tKtXDXyIal0ZDDN837cjyA1fK
GOt4vw0eM6MdzlUbo81+Gzz+O8SZtC+Ita3RZPYUst+REwYQBFHMjnOxiE1j8QRhDcmH4hzQlEhl
U18lFQmSX+8V2zBJMH4q5GTOeOjzO28xDDX/gSMM430Fug7kQGj8pRj0WxZLwwba6B+rTvrYyeA5
zosNrvp0FBg2zovayEvgb2W+aNZVXX/f0HDwvQ+GOiKwuayUeQO52yeslowY/mF1qUMfNfdJhSDy
s8CEmODtwwKUY4g/Gr/26/QzF+nGU1PTmlQHydGQuuaHteOBQY3EvKj6MD5ON9R+SZUVYGYw8b1w
jrEcvHcqbvBoJsW4n/tbqhcvQKikFjQrd0vO2xxh9QqntN8UfO3gB3jDrDGW/y+L8Z0lJTnYQEhk
s634kc3bT1RHyWLnuux77FvnodgAJl/ux9cYiQ3riQ2YBCocUo5T5RuvdwJexIiZ0Qyx67blynyo
WRUD8dP3agtJkx5sh/9Z6zrSUW3S8Nzj4ldVPqnEIormqIkcg9LkStlNPKb9erVzIEs2CCVXEq4U
ykYf8BPZksIcNY/It/ftFw9C+s5Ruo45kQsmceq/epwbeNPvk0p5pMAGjYm1uDOHDl8IpgiVIfzN
v8ETFK46E02gYsBvAE9wPV3vkILP5b63Vra9IH8D3LhRsveOjizF+N976yWpypVNbANPU6b3H2MT
NKx4bZbKWGpWX/UVtTZp90HRnPNzElp1k0Ybb610hWzn8Nf/d19llssMU+OjMRvZrqWDoexpI2Zb
d/6Y54Jc7ShXOJjoLWB+33613dYSLjmKB5tsmyBEguhKlnFQUREtsoSpc+85B76ZtsVpUhQlVTsM
Xr/DXNrmQAdFH/yncXkl3ZkdHNZ6Pxl4uTVwQpA8UBHDBMqTN8FayNa9oYU2yB4olps3S/vhk3yS
mflMH/NNeGb7aDxdy2LA7F7NAEiB3cVc533nMpPImuqysVg3dD0Bofw445Y4KP9qE40u21DlE5A1
Q8NkqoBfeYS26OXGRA8leQOIQP4Dwnhj/eVs3uanerbD1hjm8C69kcvhIZ6Vx85FwsVZsjXpvvnu
O04DNkyV4IcAv08QVWqN0h4flWX/DErOe49eXmRib1KsZbLeXoF/WGeW/kyxMpv5Q1uawsy3ie22
/XJkBYPIZR8q8UAGCwMHgbZWwFKlm5BlF60u+NyT3Ns95iF9Bt4mlGJ6DKtI5iCYtDn2PiKcCDBX
oSi5tKmoM6BIjR9YC1O5ncSci7Kf3FZPPkyhSj0Xr87kQhro2jvtB7hUiKdGDnzTCS5LzMLEOJMA
1d4C7MTYwTCFOCjKnJv4+YCxZqYcMIcH3czTox32EmYUeMeZJTW+00khI4lZKUM+HzwW/IYvbiw/
xiJvieX1FiFPbNJHvYc0IzJnKhxRmpYi+/DOXWCvNdsBTdoFtIaWRv1fylQiLzYx7Uj/zgGTX0ne
Hg2iFyJzkrBjLO0cSJkx8Q9OT3U8NCqeAn8DRGcoPKK1P57mTE6QC8upY8HQc1Tx7TPaMmAvOBMa
g+7gKaGdqM/6iZKTeteBq2pcgi2wt31ZY/B/87VYQZoZPl1xJ9GGIThBzppjXUlX4hFuunDA4ibw
PnT4RizLuKaAt4NdCNxFCYdvmTKrLoSuDoP0MQm1SgooE3b6Vs5TLam+DeSR/jgo+W5oEIp253Cw
sV3dV7ejUNWZRjkG6XtVtPLVJerLdlD8f7g6DiH94ATj8sTmvW47VH3DznTbN3fJanGdUOVLEeQZ
vfemProNbxT2yusAYCZcOL18KvJYnvpYC2WNme9Gruqy5cIOe4UBFkpB7KC3q3BODoD5c+rcOURT
PreJF1fsKrfBU+6xSMKFC5Eo5GYdVV05TAsDAOHC26pcpwwD9Mt8mFrUxfnTGshSU8qE6Ty67mm0
icCFWwYwAFixRjkebk+6HVSvXh72y3bcB7XNaiqoW3/H3WA5hwHlS4X4Rat3ImMz1bCBZIs4FL+c
/kqSHIpnUiAmXkbELSK0A54p31GLG6VO4VXEKY/nQY60RqibMc5cXFLONDcRB8hPGFPEDACW9jZx
K+YI7KhWFD69o49tZULk6IFJWEsuHarRsx1+k22AE5Vi02hXMBg7LCTKuEMPJ7nZ5TxSwRV5hx0d
SIOC/Zf6RdLSgsikaIdSQPSy96cVKSg58JeotXM+utM+/lt3NZdwx19mF4rBJb+FrREdnS1FH/y9
93AXSH5g9ZKPaD+KvOA58arHmqkToOlbtSnezRZ/nr1v6HKXgrYEL25ezUrY/h22RDmI6pIaWoRK
ziOJauJibdrx6npu1xpEiOgbQPe8qv/YyRafxA82ULWhEEKLBJC91CCcCfpGIMkASPyvmoT7f2uY
PVrGrp67WN3za/V3yuOV+rCh+qZnRoN/GqzInIEsmD/S+HKnzrAZmzBpmf5hQB6lrHOUv2zsQQAl
yPf2DKx/3THo6n+DQleGCdkCcjHOoRX/QIIQe7KFbcXijceydJYG+LEYREQQK9313zEi4fEPKBL2
rD84RMIbJYpn17iWUj8r7o8CrDlUzp/tEP9pPo24sjZxYQ9ncelm9KcRzaBaAMn+SFbuFR2dO/uB
RsPP99y9O/SPfHy8+dgFkI0d/8kLGC5o2XdI3WVZKDKxf40mHvK9cfhqBGLQEycRVMTWKLTP4haO
OSYFJFsMgEYdImuiMvgrxR3RTxCUhF50ntNJOwpLNvIaGMQEtOYSY93uQllId7YDN8ZJQ1aIraya
L3Zhlkj3N2r5k47NjS+vLlR1v1qF9F4GSD5er8M4/RG5+bSYXdElO0OkZ/53E4SrlmG92kH9ABQn
jrG47eC/m4y7TQYBAhzj+qm8VeMO5kmI3HeU6VL8kiBRiEfWvVN5XrS+RUuXTqaoCLwnsWio5nKd
9oUHxyRC9SFh87wKUVMrLr1+veC9Gum/3mnceHDHR194I35qaG6QwmsTvDNOruiauVLUS37PJvFW
WAHHpgEyHTimb2tZQeSkbqdXX+HQ17JuZbfvXU05S02KzNNMMs/IR0lJiB4n5l1U0z1Z7iwSLSNm
A5nLzBf+pTt1qVG6gvalGz1mkmRC/xVtiDZdWZM4Yw/EuAW4qTrIVpVOxlcAb+1WklbqHrWr4Nh4
PJok3gA2ymdPWgLh5m+lqpyoylYd5Eo3JrKhEEDWVV0xqZzYm7BMArBXoATXQhelTxwcsneIIO/h
WhqyJLnuK2h9E3fTHH7YU1Rvyw9N2JhoFASUytt9Jpd9K716tIDJXA+8MDewg1fbumZppWJLOwSS
SwlX+oilKrf1XSTECxhhQe5c+CnBIwCwU7RMRx+TkVsUVp70jsF+R8xaaaOYdwFCt14HCc5rWxLH
+5I+pLvJzG4QsUGHdX9KiesM4kBurdDGQ5/1Ty9nInYIuRy3GoUMINC3OVt11dS/F4sZ0DClqiXT
JA+Z16J72H7phkM=
`protect end_protected

