

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Da6prWG6T8v0fWL8NF7XQlzf5Z9lQnxgJ3sUkKkXMXFutcTC9QwG54nILyBlgRJpX2LoriK7YLo0
JdRE/dqFiQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iVzamXvV5tHBMicRNbj7fryNs9zvashabKNqrKCHODfCC5UYFevaqScmbBpMVqiKaOOUZOVbPZos
XYYsp1eghASEmoG+JxH0/ZD3uIeM7T8RrTk2AR4tONhB71Yi4x2vV1KeyhRY/Ul6/0SUrP9a2Pp9
PSpSD+8fGPC2tg5QwU8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
USDhd/cRLcXLtZzdotLaVL9UWmxPCwu7zWPz/WclJffb3OzDPNQAUbeat++K38XRL90D4b0lt8+N
rxHvntitiy0G5ki7b4srtunrdoAwXB5qSm8PXREuCwkxJf63YT6YF2Om9jZMaF3KQKwb9Euxz271
QpKZYFrW0gPfLJyPs0T1+yL4V7NfojGmqd1LcO2SSkWcP1VeT4WAPog7y2TwGoG5gUJlAHcLSgbj
iM/Htz9gATcVUHK+SCR1S1DUJLdDofR8sFEiCfig7MdFzPulujKK5JobwEmepQp/5eHZrleLC/I+
Anwydpsx+qkl3dDMxj0uTuRIoFTrwWNDz8K9eA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cn7AqgmMaLxxg2JaS5yD/MkSl23E3n/Dr+FpLXA+JTuFshzxzodBc4KGpFSAAX/mfX6u/6zVTmZq
3oVrJVVUTChYDkXOe5AftUTIpcOiwwe/i74GN55kel3PQsAFLP5K0a70FGxM56aEmg0mry864TSf
+7aUqC/t5J+hftO3N/0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gct1L0hVTPfsgjOxYj0XRzvBrEP1E9yXonvta5l3fS8lCfEiaYr9Of80t3EItFsGzdHneFXRF9A9
scSOVxUhVO1dxc6RdnrVtA9n+txOppq6iwoZJ5A2KAS7bDquD4GmJlDGjkFmZuYVXuQr/3R2w8mP
yFHDUOKRrvwsGZZUPfrN3sOL+EI3UkqGQq7b0unUUI1q5j0LF+LEbBFNU5QPS2mEVBQ7wLynv9r8
EqCh7DZqH1MqZ8hLMmktUq+NfmeCQJ65165/C+EqglKtbJY5MAfUUmyUlJjmPuQAgn/c5rtNYH0N
qc2bqKvmbJGgzFdJPy9hbeZvOuq78Qea1tRqzA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17008)
`protect data_block
1KAaN7vL2RjvaK0PbN0Q9Muz0b8Z7eNnxypEQmSLee89Pt3T/WKZ+sZAqYca6hVmUhvFImLqDRTe
6LYbiaYHSvNzZ6p+l6wgRzNQ8FD6G9UyvJVhWG5upwiIEZYq/kOWPJwRkCxGTVkpCZrz/Oh3oHr5
a8XW0bwxhCbaFOiCUcTOSqNqdTc2SyIge8VgLdD/PQMqZ7YdWex7VtekttbDTjyRcEcBjklfemwh
m7ssWlsuCRyX/PZWqKjj817DA35rkyg8yo4T8pw33oMkbE+NusDxeqdWpo7Uv94CZ8QWjVx9ltjK
RDOea+cV62Ptu5inffTNUFmrNK1EPRyx0e2nu6EMo0/mcqZW7yOgDQihl/JA+FQfZPHMB/H8FXAy
Ye4jYNp9OZGPB7IqlFR0QiCB7jQRMmLtLrp7Dz2dMFeQobN1GZ690W/OfMhbRSGf1ha++OzOp5Jx
RvZ/KdoLqfeYBNRLubrhfJExcjsK31xMYw4Xc7a6tUxhO8sq79r9szqx+0Egu2TZZK6HD5Okwevs
6imr10m381DhInumB6TcdMAGoIEyZozuM3TtZ5vrfhtV8GuKcGb6OEvqoh4F9FgywoqS0Txghujj
+7+9UckbLkEiwmiCax6OC8Nxj2ekaIUhy9enIoM3+aMHc34/SEKw0Wo9wqtrAv65zIa9I5xT+Wm6
l/RONY5oh7mC9QtUkQ94UdjpnQCVpq2AGdIjvui/rxhrH9FsniXx/wLVJJx3ujFsZYtkwjn0aY2d
uKUjrLLCmjJzP4lspXc6HXIqHFwqPgDOQQnx1OLhkNKKsqvFoVeUW24XQMKRfUIdzVpabIYUdoS1
SKPRuIJxe+NObBEtQYlGCjDT6X7NN5Ei7172mmLunLjF9mefsDQs+fe2mrAlu10kvNTZblmAxAxi
57WwfUsz9sPMLuERLUYkG43s1sfNjEf6nrIEroofvAHTK9T/G7/HuYWztpHZ7jjSSo9VhmMM1Hpi
Tklw2EptkR89352tAnJHQxzAB5rp+2V9kygSrTL5Afrsnmr8gIgV+/RP3xNzfsMgXaKYPYqPfh3r
4BSB++rO4hwwUTD6j8jMsJPaRcFqaEO2rVglGjlcVn1DWSeAoS++hXKVL2jlY8hVnwVN47oPbLFz
Pd/HLvJ4AFZVS/VTpWRSSk5nA1pC3SXeoKVqWZuaa/VX6YU0qFHrz1rRej/IQZ3DcMV8bIIvw4SM
70RXs3aSmRr5lQhA9VJAUce4chLH6GbJTCIOjJawCSIwHM037QohU1nT6B9GB/G9Qx5WHDBbPnYC
i5EXvLSRfIdt0v41/4kmEdY/mcSjb9DScRxQGjBKbBPS0gjOFUqVzGVfHOrEHtieNNlV0WA6CpGP
3DltrsjC0rPLdTuVJMEqUcC/uOMu+lgAIgV42cpxBaleAgoU3wA6JX4p2Kvh/3bh8ZQAJIsWz5aR
8nCsc7ApQGBMTmSwzev2FTfXEl4QQhY1iCwDvgRtNDt6+m5Y8ydlt4L4evGE304yYhjrk9nyXJ52
gwBce+xmFbVB1mjkK6Je3/+HCMZXDh0FdgZv26AUwLyYL582kxGtxUws38OgpK977l71ZYROp9xJ
gc61HRDfYdUeEet923OHB5cLR5kn2sNujnWpo3ZG7tIAwN8d1kCiO/l1ikYJM2Euj5xC9KfR1XIr
OedpP/sTG1XL9A9fLJzgON27zo6egX0toJR0RzKRLR23Zw8G+uHx/PlFofclV5bj339H1PVpyrfn
BcvMhnSBqLX4hgTdDTK+a5TIim1RSGOKs0SMwnp+GftFf6YYPWtPc2+5nNic7wwoPkBJfvfAqyvH
w003DVVmJdFvBfENJ1kDx9JYHCEVx0VzBBBAVfUOSssxYQpVyoWpbqWzAXssNilZBgTNMxSqmCCF
22adHgF963x/TdYK9pXQEKrLWooZSBT/saeKOI797zJdw8zTgHufGfhby+OCJu5blS0MBDL4cvRR
yZfT+CAxmSAs7oVhpNbx04/NOSArD2FY5UaPwGg3NVE0dCz06A+yGu7RP8RTs48ksqrsWcidASwY
/6yIRPGjTVoCjqsPXWHVsqx0BiwJZdyzIVjlNVwwXVxsIrP1tGIU1xnBhgx8SpOMP7BHi+VM+1/w
PaIrcm0AAQh0XuBGeEU5RtMZH8gPLWW1lk5vkxRTsC7Eg7TXeqGA/j2hLLuFJN759rmDQ96ZJ2YM
uJXZtCaqwEcHVLrQa16WGKoQt2hYx9jcjen4ll1djdGm3BRpvoEWslLKXfoRH962Jg/47sNUxjtA
ouREtulaqUpZJi7Yqap8jt2zTp5tpgTB5MJXWwNAj+FQn/P01P+epuCNfTSAg8YQdNcK+5vN2OSU
jdCWXJKWcFSkI3CXG8CBgzpkkLm5MK/zl27KkC7AF6L3sjeHNJYFUbOwVOfR/3Bhx+awHUEpGM26
3jhaG0YcuMTMIlH4+BaAT9E8NRiIucr0zq7Q4Ci1lk2w+EJIPs6jCqZBEnelqEIFbcy4XNW7cBKx
Rb7vRn+ygp4o15ZsiHFz1C2UFaugi3mWDYKlmTv+EtewKApZvww2nHg1T34KLjwgKhNVfnb0qLVC
EnA9QtfwZpp9wJvd0dzfQnzZ/ArqHk6qu4VaE9rn+vT6HqxULMFvbfMeiDwrMMBCf4rYcW4uU40h
6by2CY04L+yzU/qAekWIU4a/tKEXoc3W1C2/JBBp37QPOTBn4Qazeb9a5wOYy/C2Jds0PWpcq3f5
Othlgu5XTmLGwuTiZnE9W8ORQwuFo3anQyxWrB4qD1KaRyCylVm9myeVjJnwa8ZcOwv2VLbxLqAn
aAeb5nzXbmnC9b31vHbHsbgdsbbTNXtSpqQl/2iRgc+3NSTTEHQBTqHlNdWgKcDabVq/pNM+GFk/
ZXHp6lJwVS42XfzfjG8j3KG5TgkYv3PspIKxFge6phoQbhO/KgLUR+fo6OZjo/1ioEqnE5Rc/QCC
TJ1OLvXmsqpTd0Q6BMcyQL0MRdJZYNVOfWwo+n4rdhl5yHPV0EHBW/ky5XC4usV+prAtm+SbYUV7
Zq/3edrTGKGjUEVXhlY6+ceG+ujH6KUvI3V3QVjD3TVP/tbkEpy4quoFYSHoItKRz0boXfrMyNOG
ca88O5QLkIH6gGRa6sVEtwpheDwMv1QgQduYtoHtanvOn05nOLYnPt/pGk+eVIT5++3lzA+0A/SI
IYqjC3Yt265mDFm/v5J/gf+s9MDb5Ju8Y4Fmt/UMFOnhvtXXfMcZy9tleDUibMv9MvtJuKIiJKzt
/M4ZsEvQOHzRrMhQNT8/7GnbPQbL285pt4ZCqCvZR7tJO1ChOo4ELXiA92dAU3HVdQV1GhWiGI9/
QUv7j2upUUsYOlBe08csz54S1wRPD2qPQJk5MBKp0xDwkjw46j8y3WKX97BjQ79HIHVPetmMoHUc
n9+6VKgUNwCHZzTk0GK90XjkpTJ5o0hzWrjVPhHjxKYlTwzdIBQPTY7Mj1O1bBiKtHtjxvJZOk36
uea114TZa3s0uyF+JzN1KT7mtA4QfR7kYUQO+5EryjJisWRaoocNQfIQ1ivm7SInxjj/uh8WdIGf
7iQQ5EqZlsBRZpkwzgT8tDIdySBTyqaBod9SFyw83Kta/OjtOmMCmdY2Do1skRRxzpykOFcMXHo1
DIYrrTWHdyW/46EYmAlLjqzmIaxylAZFshz8f24OMONAMD+T4pOuWQDUF+wZ7XrQMAM69th28FNP
F7L8CPTKbiMXzuot4baMSP2PU9sXZRHv1mzvWdGsk7VpmP4VdtnSL9YruDvwps+unqn+WY6sAyPJ
N6vA7ilSnREqUATyAcNWRg2BpMyiXu9mLLAxdjueSRzTcD66jQzKUD0sb8B5GBZmSZ0t6cFJkK9w
W26kyGKErSAbK06MrCLUZliyBi1aQA2lN+6PbrXRPkFw4C6P1Qeyk6BdLjEXzyuwZ3sViEshy6lE
yhoA9u53EVwnwhqtfq1iJrEiMjtmp2squCHwrZESal8yqtSst9IGmBKR3nnsBDhEw0FaptVc1lyZ
v5HFPZ3I4MingMshdajtDSO9/NTxwnU4cDhcxEv2XCca9yYL08B76SIe9kk17EcWIauBy3iX6Cjf
qZkNq4XcHevCIwm2pI6izftskeMaZthqu3SJLHAkAaW9hf3QCvELG/cG8lx/3SLV4gbMCEOO2URT
mNuGXxm9aVY+kPEiZFL9A4XhZVOoywU75o2g+4McesV9qnd5kHDR876AgUh23brs/KwYL3UagBaf
PLEs0l+0ydbKRLXMHIC4BAgJDxR/CIiCzpP+YNmBKI1QwNJKBqwhrP0gHI/x4ivK/X7chB3oPxB3
mlxFHZdsA+oTQ+Q4TSbaJWs+vX/uFaO2nHQ9rYJmz0cM7YYYkGeu+IZVqhICAuGiCtHHRj2mz3nS
jipS3s8k89JxolfsY+NiLKKSuBxYkQtmoYvwxhxIt88unzOJHtchd4gv12Q8hpf5zw6ZSIhQtrJW
n3NPvti0EKW6iaK5EwWhpqQTm+8XAvYgZrnZTIYoLl9CV5n9+nyJd+/ceGasswPl4ud5jyk0cPEa
dseaijbSmE/HwcWRimxRI9OYbqMpSu8+HL3Vnka8/WUss3GdeBUK+0SEdVPvtv2gdBeDspBcUS/g
QykVbQwnR9OmX0ScE4tRQUXtEcG/ffeXuk28Dy8zfRxlm5LJfzk4+nZMOrUw3vwNV9/ATZaps+ic
IFomVUteljkXBi1aNXePkb6C17vHiu3IXDvJSjoQaDorfCSxouYdgtfQx9B8vqjYpOSV823pD/Br
4avP5qdwqCxSbRGxSa8I07cvgMr4dBdeTlJ1TBQlTSRBK8ntJKFRBW3ePtDMtUBDowoB/z4CxmxO
skPI7U877MmJvNOgHBW1Ndk8EAxPNx+zT0efsOYXUEgHI5QnFkUFCenEhYp59vuIk0GMuThV20os
sJC5KpgMdiCvfiWKcX5HRmqEVKggXFd1UgVnF54PmWpiK2Zyx4XOYbwbkpEIvMKvrxEHLAVnQau4
zD89KIN10auY9Q1hbgBYR3Y9eTGet0vvoRPvWNzk/i6YGZsx3soAA/yh3YI+ZoKQXqnmeO4YxZ+P
rsesM0xFxvuS/hMcRc3aWo7RjKp6Mvf18VH2cV8nMKGApUSvd4l1EZ4qu4Xg7wX+JeNrJaVCfotm
diS4DYZJBcpXWlhciR6bhPC8o6CkCfC7lqo7nxWNArGDiViQ1FiGVTz+S1ZnD0c8ans8ZBC/1YDp
8CJi7O/P3UkoDkEwAzzqTEC4BE1+OWSa2FmYSq5bm8+yDm+09NmMJHb9vtUsFZeq5fgYbqG77/OE
0AbU1+EWsDM3KJsBdR1ChyR4TYTh9CeEi5mms/mfEYf9HHGGefGdLMmcK+RI8NjNrpWvuysQViIM
ICVFplKi/fXm8y+OhlZDI9RP//xskbafl21gel11/EhGjh1BgFxfHgV+s4xSch7lL8r3gUOy/Qk3
DBGpn8zVp7KZME3LziQRvUcH7SM6IxQJUduoq2Phy4agUbPpr8unJQCcKXmhw95kTiVJb3Tvtcbb
j+vrrWvZ9WKm4cHSPlDlg/xkrAGY/aoF9kACx1ECEXwd10atru7bIbrITz8JgFDgOHjA5Tf1pjBY
2gu1LzAc60+rzOELmbdFRirHcxfTRSmtd1So8WsQnEjjoICnjG/n5R0mUdmEKJGXkv3j/0bMM3Sw
OcMhvWx6PSHaNGAc/NTMEtubk54TsbeOWNArHnuVdYt65Ah8Zwv7oQTAdtpk+O//ioQTZ/3SArrW
m/G2Ih6+CNONwEtcEqhyP9vq/3q/cYA7K6D7+SpYdFbVXic+/uaI31zYt3Zg2WPHkGv+DjvttXzD
Nb5h/1f/fJ3xHN+shFwpFP1kuZOdqBRLmn4lKrOxlBAPPrgzyZ0VLg+KjDq9plPTpVjutcJ0SdKe
DnSVEQKRYS6S1rIGw7K4ch3rBaNeAZifafbpdYb2yBVFfLdFGH7UJ0XO1Yulr0p7e3G50tYKrfYy
KIoowswNVN1LbqBdE9EU5rjobxpbN8nww6jcmWj06popRysopUfHmEv7QAj2j4PC+kZpbbo3oRNk
qQ2b7TpPey27hPaFlAdHOGb788SwxRjzRKyYB16vVKlAmYJYrl9ebLrqYtTUyfWPujPDemXJR8xO
RrGCR6AQDB80HGUHo6ETrLRarX89oim3wb43h2W4YHItKOJ2arxgWQRUO3C2282MYW/YpOhtc8Qm
5dgOL4Es/SVn/9my0Fe2HtmFrYe7UtXRZp8h15bTC6iKCelX0MtEYCyOujjIpIBxlPyCWIpN4Ql2
5YVJHLJdfDYqLxh9LOqJS3M7B4pzwW7piSi3ojIk+DH0EJnVIMVMXtqHZypWbOZFxciIfnL9zwe8
nBWDpCXwQwUMU6nOMjh9kRXWWOMofz49ZtduQkSERmWzi3uwQ+lCXo4xHTzVg9yabN+j8CI8V3K7
fQtxLOmTE7uYaUAXyflR4PBWuFCvnmn3/B4xuZ9riGCX4DlkmvG4x/Jvw0kBcgSVzaxNmnBTRAQ+
LMExpEVwzAa3GEUi4pahbBa56WL/dG7xWaUfbcFQ0GuxuXNV/xSDzvU1iiF+bdzdkNH5CrftAYxh
AcCKLF2eP0RbCk4V/OiTwg74B9FpNpa1dXT7YWgPCdPf75Hn/E9yQM8KJkxKKCsh5F6PatudwNl1
4r5IzLJPCwtfBYyxOkjshmZFEdRHj5Sfa1XxkfFyouPicHtiRAbSz7Tz40LcHDW21nH/zTMTzLho
YN1slQazwvh3afnr7MkTmpB8Na1OW10t3RdOvPxCqJsByWCxtT8AF+gTqFZfw0gZC9EfyNf0aBdF
r2otD1Z8l+wVK0DyHF/5T1KpzXapkuuACEKBdZGprmmRqUMapAQ39CNdV6fmbMBdtHZWpINMEIx2
OBLXP/3nXWfnif2P9EIeUHspEzCdlX0hAMtmV83XV5+wLLiPTPI61n+6aLKkaF+JeAgQRAFz+fG3
4QrwOMsGiiHq9DtUgiUfvEG9OpLhvlqDgyMn7kodk7HPyFEnUwkMQHv9ikhTtvy2+nm9ygoBzW03
t/3Q/VtgGBencDz5cru4IVUF9lgxJXrdK2zUexKsmYwLf2ul1VWn2hvYnhF1SK+BjIe+oQt1OWAL
jnt9N1lU4b9/kyfRTqzFICMC5z0Z/Jq+r9V0+dN2BHKQoBKmO7eeEGdoselyxhtyyUwBro4SWF8l
nKDFFc7RR5gDOB+Jod2NeOvlxfGpCQrX5+zNwuQhTGi48p1O4aNbRdWLrqEPo59GV6WQ7uziTmgV
XJv68mjwCX1V0WNzicAWT8qCdYv81s6sc9iZzE30FMskxLfvKIj06ed5LImrtk3soXHdlNbYmLtg
Kab2ySmOxkL5dE/tk3FL9yn7f6J7lnLpW3MXPO//xMnhY/YbBkAHeK2QNjwo/ovTNlgMYPtDyHHU
LfB4fgqryLT9yggv5uFc6tCCGZDbLcJ+jZWlnQdRw1BphtjlfHsAywkXhnrF0ZMp7AVwWkJZ4bg1
y1JqVHC0McWXwZXmyRO0qMmZWdMm0iWDdGt7EoJ3lc5Vg7DPuz+3tciKed9PSIE2KKkbl1VMYSwp
2JI/tN6dsYyrWDR1DK1c07rud4X3Zzq+oBwHMr2qhg+c5o0EsN9Kc7KxGynqBHIMDgl5QD6BOFAH
AO8zZi9DtJd62m/g9aQU1wEBrFL/rc0sJXxg4wuDcJGH1ef5JWaFEAg9bMpcM4kLzsGr4gojITHZ
NF+FhLECSYhKYirNWSUuUjAcErkZGLdFBCXhhh83JlSp1ZWDTc7+9gxPe222OMBH06dIHepAS1l3
1tHAIn0Ouu1lT73R9x2utDB5GvPDf5m2cHYoQfbE5o70Y78B9MgOVCGl0lsvO0npYrdbi+J+skt8
j0ZIDrHGz7+bvBldpiv8t8wx0rU8mS0KExE5Kp3JW91PHzgzRq7ZrIHOJEB12TMUFX6HF9dGVGp5
fbo2JlmU+DL582dQSlD1zQRpLnLA9CGBBqGoiGaVPsQX4jLmw+wNFsEmdXNACJqu9GDVmeRoyM8j
HGHFOfHmxpBnQAMdVqRP/BKbdC5JSPfWnPGEYIJG+MFgopDxl1/RBIvGbW8UJPd+9/Z0ZsN0NR3K
tQwP/04P3cMJAcghAdSjbN/82fT1Qn6aZcbatD4ZqPoLZabAYOH+AsjRzcH/4rdFmUX5X8P9NkGy
Ll6GQw/jCmH3VZhNNRPJurMtKh/3ipJcrPKzXwQq4G9SUOHIob9cEfNJBEYgkx52LYrBR6qASuDy
4Cp2iLbrpFIl0bDidN/gqxFzDbophapGbwBaBAW3d2XSXH2yOdYqpuz6aoz2IwPf2ljy1MmD2c+d
uhLNOkux8rTZmZAtmPvmjKeIh0Lvwp+m8ADc84U+cm54DSIngACKvKCj1R9qIKDK0K7FA+O1GO9g
uTugTDyVHB1OV0ur5+Bkaa+Dqz55ByZdM98UVzyFuJ9Gn3vC30wfHylgRq2yDimamSKU9DlYSow7
8YNCcI8914yITEbCwPU64AGW8xIUo3Slwa9chrp40hcV7RoCNrbFg46eA2rLEHX+nNF27JcSVSEQ
FfGGQ8Iu+KqNS98Ztm/joj/nLUMZs3RTj9SrfMc94/1yHouN/xBJwICLEq44enen0RA9ehGEf1Oz
mTLRU3fRfwudT/Z64GUf5xLIa/GTxQ+0WpXf0T+Ezz/1UTHdrXeIttnCowXu5+pCWDy8xOb8AZMi
QlSD+TQKham8D8H6UBpoG9jLPz594Rkrv3dbfo7oBWcgG6DROJAsw9nn1JVu0svkp+LEUUjearMt
UnmEGuGmSp2zU+AAXPbRRAOPgPhjxXJpJ+dvDZyP1R6GI/4gCdYAC+BFEcul3lX9UM/iQEV2lNp7
Q2Cy/EJsDix0imaaxEL1U/1u4nlAwIY8lM1FCUwJgsiZvF3nVSJRT9WqgrbYKuVCzoTxpfoDMduz
wk520TGIqT/zAoWgsIkk7NAyphlntYeOOq5nvGM1Z18F2n4X3EJEzg+Uyz88Fm46nRNWtT0LzNqt
YloGv9zFxO7UbKfdKUwCcyfcq45lfclqwKDDfmXJpsSivTeDdjqxiEpNYFGrK47zSchK6OQMhxXy
dO4G9arcsZSBTOaZyWkIkY+2R+GFv6RMllW9XSJ20qEUDgxPz/lXLNpTDfwrr5/zjulvuK7vd7iR
6Hy+6Zm0FOb52JT3rvznBO6LDe3/1++drGXjbYVdoeEfz8zi0QWTPU4pqaNlxIk1MNS7EWZVJhis
8sOu6OHPFbtuRG5dBLNYWoA0XILRRZEf/2OiGffDlC08M3KrulaEQ/tjicZKE10AuPmNoSq//b4l
5KSMmdS5CIwL1sdQgO2uklroBAdf45LUYLc9sAMI6IoKxo3Xbi5c7EP9IJEtDJpX6f/IIK+DoqA0
ZI3Q/JuNQqR1lJfkMA0Rw7+y5T3q+XhAv9RDQngKxctLeeOrrh4sOi97cDK0qqd04CwHFwdjqFNu
dU8qJmYkPQMcJh8JmJsSHB6y9xz3HP6K/560Ku4TwCujqzw52ewcB3vKtJSrQ62C1XWConDXTl7w
CMnFlUUtdALYQ0pAbPm53CMwYIkdb/hFKaIGE6a9AdUtWmg/w6FwdTacPad1bhc34n9REkxmDSsz
IWlNauHwTFDhTKwVBbpzA3PXv8RvSvQ5g6RGYPrnmhxxA2xRixw5iQd5VGlwWhk383Do9u/tL2sN
+Wkr3YfiTZCsBfIAqGrw52JkpuQDK6tm7tR1kXVVoc5aawtHZqdak6zLZ2Oj5PZrVBgf6qFnOfbf
0hjOcWDhz3dgT2KhIeKV0eUaVkGYa+lmHjEz5698LtHQ0TvrKSczE9AJj9BnYwF7kd/QDYqjBs9D
VP3WWik49C/KvGr2gtyrxQC0LdzxvELUf6IElWmS/2UfbNjSqigl/oY7jG7yUh4RXuZ0Y0ZDflQR
8A1ALsnvfaaLdn+t7lzAnUzQFoEJbf9CANnHKN0PKO6nyqAvxSr4DBw8e+gaVu7LMiQClsNHi1D3
mJuCPvHsH7AS9t8cO6JW7ylRkmE1Ulqo5CWN85are8eH9EqRbaPVQfep/Cmm+BV25JtYtFnNCg5w
4/kijw+mGe4nFYYnpEyp6i291VFmQRHjGyybb8jHKdiRff78UO4pF7anzPwpN7APWjbmZy+QEjEz
Tloo0Kr0hqhdB7Gv6HKB3Recy8k/YOTRaayhwjMdWIFZXBscs+o1im7zzWXSzSmt9OtxOLvYqlSq
W55BNThnU9MelwIChKUC9qfuJRIb7klEDfKAKEufnCW556siBGomH+ThhYd6DihD30MW/6mlbQZI
K46WBmyTudMn6BzL8wIwp9smoL4UmJ0rRp6O+ePsam96XQ0spTWzwT6uZNBJtYfg8mA7jcHdMlgL
IjVfEWHJDv0tq2VlghRA+SmaAN8OqF8sMBYodm+bUgwOmkttI5ZqP/MncqmgzeH7TXmT4beVriaS
MXQnJf12UMm6Agb7+mChLbptU0mhYlERawpOb4i4dS1ASEBs6I9C+H02IJc9/Xk74qzNvJc8pf0+
4v/36VAba9GbtjzlilgV4nggRsYeVLOZF9rnlU9JMOuRTivxLaiPYAZ0+6MvsJOgboerSh6WmpK0
2lFJo1ZriqPnMDHjrukMsLQ0RutJ7xLdOYa+RiP2vpRAlPJ73idVn2pkGdQoc52+IFgCfQ9nJOPD
ibH5+NHILtk/FxNtYAux92fp04PEBbuTD6MaQjrCD00KARkH/loVaWlwjSE4FqvNXTJJtoZ2PHGr
WsUmsydAIpDz+mT8xxuDARLkqvQOGSyOUO1XK+NWU5G7kkKmqpzLo+PTsQJ9RDjSsg/Fr+QIB9A0
h/rUgIYI6xu6XWmXPdDYeSp6hCKrp2iYaV6QYJ+MPer+pD5U9rcKPgcp/xx4bRBfY62CkI/8cyUx
eqYgmxwqn481VnMjk3sj+wgbGj/IZsDHmV/2wMUKay8iiEFYz3g3suA7khqXjObqunsbWd1xRYen
7N7FQlRG0qNSl7ow7baHtFrbvjvZQqnwSmYxWG6cBNYkN+VBjPmtNpcA/4h5rYrLYCQUNBBAiPA0
C6RPmPVdnZngvAOgwvYo8aPmVKZWqPjEO8PhiBjv0Q2o0GiTl2jb/pqwxSALlLnI16AEnpgezOp5
OpAo6kCANLLgGFsDshK+IbIU8qB4eBryqAt5qad/YazaKK8o9tqKuPu/q9FQMGgdNXowUFZV1Cuu
VI8u3C7n1x7VdYmBx6VS52JSHSPI+DLPyK1BFxIMmiMoC5LbqYXHnJjIpQVhqs+dc9uku/Mt6qjq
HPbJEsZaGx+NYPkcGaCi1/nyUMjo29cvxi82UO1Pg3/Yw5xj+uoA4SL5DJB3W91c/JkEn4JqVhlh
9IckMFoIorMjzN1AhFb3bsQ7iURpAuIjy4SeYXD5PshgUnyDRIGSjlSfTGFkpW/xjDpP/zu8JEpM
lMpAQdriMtX6nIgPialf94hV1Bux9y+nnUxfYbLJSXKmnJ9H8UxgcWHdzdHLXE0dj/UVg0SN8A/X
kVRDosDExv3xMTMMxETlKI4qIqf7ePg+JOboj+7iS0hNNVtsXk7HWmTMY44BbIXNQIZWTJWKlIuN
fXJxKMATWqL2nI8Ers7qN6Am4oDzB8MgodMR4aYbSPr/uwXIjbDjrsZ8McOKI3qSrzPsrmaWx+qm
j1dSkrZFrhu9oz/7wRJe53hdW0bdjPgLQiSDsbpJXApL5xyAePei6YUJ7oN/sQ077LGvvU3g/y/h
x3HClDIu82V1W2+GrmODcnlxQNFQNtAqxp+drEObKDOt4cPYIKvRuRqKVshaIyTIzKeJ4AqB9VNe
toqfXjGWCOsEvZiLLL2L98UrxGbDL8PJMiI6g0epZDmHJhMUIsW62KsoGrsQzNMET49IJHjyIJVm
2y0NWt0nMH/DJ0w8SrPCUXVIV7nPGQpo4e4JeN7dp6cQARzv3TXWJkK1iRLA9b1qOHYkpAE4GCvj
ELfA6H7d8JutWU6Ao0qEgTDD/rVnZu/HlKYlM/3L2WCGWo3w5y3psjtIJAhP/PDAzEbJOthDWeI7
PcFby3voSahEfELxJopbba9ac1A147HGmfloq433pN5FqEEfEEi5ala/pJ810SL7sqCI3eJ2PYoo
xV1NYGQMNTEBkuVZjHwG4/84nozb3Gw407+uwdhyRkyN+zvzFJzg0LboP5q8L5xTAavIdEc28yu8
xuYL33Y0vSVqut8kj4Upr+WFnDlLjrxfdjxGRF71JjxyUQU8RNu7fKmE31G6J05FXlq3/MhCNqPu
/NWWmpCobBlSUM1gRDOGoNtODNpobYkGEF0lagzYu/Ekbex8fiph3nn78NnHzV/bP2BHGH0GjBhS
UOx4WjK40xBWz88+UWvL9lcp0LnIe8D/va1mUP3bpGjq6+9wHqXtsHizYpOg+LTaGfezPEBmZguF
WQ1Qr/yulV7V8DrRrh1YsoBh/Ww4XbYOidTY0aa4uUb8Fj81ovNsOWZpwrh2Rfy8LUUkBWW6CWVe
CSiYcyO6BEf7nmwcB6i64/Lg7NHBXAlOMEIEhvO7pnFpkka7F1c0IPh7jQqixSq9Wv4LZlnwBrJM
fYd9a1ZrmRvHPCs7weM4tWoCP1q1528a/AHsKywX7+NiKSK3eaQcp7Ii2r8OSMN189dwSMKZGCzw
u3IAvxw+rcIYZaRh7R2QjR673NuKEcFtm2Qbt/8Vm7e+FwJ6lE7dBdkeZwFoJlKAxVDCWSs+wX46
11QsquUpM5IIEOkf7tCCW0bHPQZdBkD55Dum98X6PioykqOOxOkSevl1RqkY2AKWoQEL13Bzxuhp
eFAYQ244cmlXay82+6U9IioikX+Gjm3yDpJkpIfe+hoJ9ATgykv/D6hK5CLd6mIhe5+PYlBqdPvc
MmHF9DRe3kSEInRt8FBcRtk6ZXEZvkSlaep3iOu7F1E1JkTHMyDIPA6c/2wSXpO+rIwzKBSEkBQV
kwvcLbLqGFbNRuvsDs5HHYaBLMf74dk38kQID1T1Wp+0y2ghQC8fvHFVs3kRNOUkOfw5DcJdqzVI
RduhXLK37BFN9t4Y/7rZScFQmcHNVfJLLk5Whw8nbBWPTLtQy16Jl3H1T4jYK6v6hfJhwXO0wnsT
BO1eEBF27YRAEIjRcb0iTEUphM7O7z2nlnw7jQmoHy2rjEX/Zu3s0D3+NueJuPLeRYohsEoRS+a1
9Jop81CHotutk3A7YA1Pp+Thr9ezQ6knfxK57vDp3NL/SFLDQeTQQl29Dz9K8WjmEo5VDzqXgnnR
IvcfVgQzFwNFsh8y3UEDPdRCTis2cDL2cQaqDsZeJTDKmcxeqhXNk2KtYSOqWiuox93Z+7lF96dN
To99CYsBLBrr5T2Ca5PRk9EvyqoIeUqzBzVWsDvZcZrNQ33BieNfXtlKYKNuAYZ6ULgAQrtUfeYF
3Afso8g9IDM5rXZjZgln33EASxNiSz/NmwFRRsIY4jEabnxFBadg1G5NlqAkOXMDHvSl8tT0V+JV
ULbbpfp70vEs4ZObUB8OzWNDcprmmRukeoOAw9ApjxA5habDh4tJy3KZm6f23RWLnysW7FtzJrJd
mYZwDLGTQix+R8o8EVpzqxqerlMw94QwbA/TzgTtdgoAY9TUUso+vH4OqTMfiVUjiIN9zdPVa49r
UFZC//cdJImdTMkLpp9H+cCqat8e3msM6Ezsln4AwL0bMZQyeS89YqdzTBMgycF/E6xMDTINX5n0
6YWNFYsJiVz5QJHUsVdj/JTLSqmNuvDtUPGeZL/nRY4MkXPwfmMRtffvIS+u9EizsKtzbQihHLVZ
CWhvMTaYEkTgsgQwuWUjgC55uNe5uSdEhRAa4zG/NsL7IbeVnMMMkA14xtgKAijqz7ekwH7DxRPq
2dJ0aPkbVWQzuLvkIQAKeLysd5IPB9f1xkYHmUMQ2CvaUKeXmt+n+MHE8GUoxo0RQzKaLxtIPWqf
AN7z8J4hkmwWO9WlwHruxjjLRQzVrpfDEPg4YCRFs4ZqWOCeNSOMF4WulfyDSLh4t/6zQiDMlqY6
dsgD+t+mO8Up9WwHE+3l0YMTUvsXXk/tkbXvmiRgyeBRYuqDPBboC6ui7AkrP6cNatboKxds6Rzo
CsSb5Y6H4gCFDoynCxNy9qm3Fr8/lHqV+u2tgY1Plzp4HSor4tKWnzdtzBEPKgompHaSj0HexaZx
FSruhwmiYArPG2SKRvZ8r0PzHklgZ7DLrfwItwb4b3ZJIeCQuA4uB0LOpZBaHUIXdmUAPJpfZnYS
HCO0GV/F4hB/FyZJIk1x70gUlRFpKgmBxMW8pJHk90xQKYxaZh43HXNL0uogBZjAkYTIAFuVDpXU
VAOJxMiATcisELodzVlFzvGxujsKuFO5wFV2xlDhwq5ZU8VpxcbD5oTgllM2+9Bg06eATq5xCAki
FIUrqlNzQJFLF3vLbB5dm4JtTk2sbtZVowk0KmmJLfaEltu6tvFDZoHfe9KKqzfBk5tfPrzld7Pb
0gALFQpMwHD8x59irvUaLOFZaokKMVwQELVeZrJx/uQPQk/LzUimIQpvalETzl81PhVqfW8TQANF
iWd1c9PysmhgGDMgOS3STgPLxMTwSVmp7nS5Iw1KLheoNMRL8jj4lW9MBhtcD8CYMbkMER+80p0j
1QNIkh2JZo6VCxKfSc9G3CNErKdwokYN5B0K6oWsd3FITL+WQswKkS0iw3/VUpoe3fE1U/AEAR4Z
sd6mjGLc7pYchI7mxC3/JAMoJw/5WYl1OPctuuwqfkxER7YsBynWF9LmaromyHoVKVqN0DWDtQxO
sQlN+FBZuENFTgA3unnaOSbZLYPYsfsMHLPM6/jBokuOA/82h81YH+7Nff8L9ovE4f1ossKP3SLq
JsASAALkVHlAq9K7E45wnU4xEBNSZ/fZC2I/zcrBUWOuyAijP3QuB5xqzZ7RW+LO7eHgVbEbGFta
h0SZRtb8i4KfB4GgmZkU9g+imvEw9TjdGtEkQVmdYE5iOA5trQ+f5jXKwXpL9GOMg2jX+2zbRMwv
C9MAxBdklj0Fn112h557Z8KVAaWsKx9Ggbq4MEploY7+qu7A2MXB4tW4fWbV96m9IZDEhBcxrVTz
56YQQW+5IGNLNrGBUvp6LiaSdajJ3QJQ+97TEkQOA2enVqw+AMM75RmwUsTsL90p5iLRHGw/NZOc
Y8OjBK/rH1HYstsosK/9XNrWYdYnCJ/f95DOBf0NSR1Np1C3VP5lF6X3KsZSS207vLs/c65hExkw
7oBtvsDXrM18q4FkLa14CAtFyspn3mkmSfvDZpMW1LOzlBtzEkH4rAcWhhcKreB1Rh4jDOdSj2Jm
J9UwvKFyz/+72mPKiVQbMvzEbUqJ9dNKyG7HttwW6tKUoZ+bsGBn36mQzinoZ29hPYiKKCsKyOIf
Y608uwivOKNrj6aeG2h5kH87gDjxsWu3zSn1M/dXiIcVISJwV2K5uF1D7e6SlSwf4R0Vb0DmJRf+
BqYrQCHEuK3btfE474hKEjOErh5NRKaGWzpdihZrRxpJ8m4IEOYpoVBWWAT6/FR/YLUVTJFGBVZK
kYFsGDxRkGEReHkGLJWNxubyzjF9T6ClTi2Q5+PAkJC1nZiT216oOcA9mOBiUmCXh2YadP5v8CdS
qMFV6ZcgKXHsUqvBGIfhGRQ1E4wcWpuv71JWBvAZbhxT4gYsufnM4cqrsDSBlxoKn0kk+3GWsHu6
y2NgyVlfn1aHVSH10bkKcLSjOosINj/U5WM7RKbNR1XYNLOwdlIrSzgTnJUIzW6Z3oMB8+12KVOF
w+slH4KVFA8o0uwVCNDuoiu5NqRfvRLgNDntyJzRgzoCB4vopkRmxNgeiqPsL0JcWXn42fdixB+u
dkd6YURoS07htOrDcprSP2zQer73VqgPIdi7hzWKvUH5MKpBBePX4+eivBRx1JI7G+48hcuMEwCj
tNlgs2TkENeqSE3huGutz3J8cmEohbo51SkumubSw1LIm1uy4nHLMRCT2r3anPo8HmNZ2dryrVl/
veQA2wfKO+CIPOOKzFXmMb8/vrMFG2X2EZHe+y7ip442f/OJQwvDOufaqW7mmyJ0jEaqyAyn5q+t
2YRqlLqh/IbCLLmTXDttBOzl6WORG5hIieHEz5/Z4GcUh+7JS6bk65aHybOszz/H0lpTCunrc3ub
CgePQMPxD3JUzUV92iWsa2RthOqOtrOE8nWbYKYjqLWjE45u369azu6WYgwZDpGLQ6n2ddmzhtjG
4mR9EaZI09Ydi6DihajZ17ucadR9DRAbyRHUygkvP0HFf3Jao+Mrkb0O7oluiyUcTZfycFC1mgXm
fsv+v6lruGrd+sB3H5aPswhOf2RkOEfBUtAu1PZpcQbrog3GchBsg7DBq0bq99pvLeDTvqociY31
DYWIEizF8dD4M9k8KCjP3dTMi3QiD65PuTUWh5FPhej1GTeyLukYBipyNEQWTolFBOJNH2AhHFkU
T+fsCNpezn82cmZvdEvOfrVM5WCneYpn3HlXaZqb8uckEa+3fMBNqejQNHDWxiPnM9LtKZtuclpV
1os2+jubC8L01GTitH8k15UEqCckEnXMGRAEm7Dhryvylvgm/RRjge6kane5WvIJVt1SXkkrsn1D
SGpEYvTy0dBQYbQ48DZyKPZWo4UYRHlNGkAxENUVkzVcvF+Hv6FmYeEXuqtSlRqwqdQzDFvo+lus
5CQFouynLV3czOEed2YWpqKfUtIt+1rQnOLXrXzaXkmtEPCIbdr3OhRb9Z9kb48zyeob7u7x6cAh
rREz93sVVehDh8ymbXbhZk5QoyZEnv95MFM56yL8n3/ojtJ0cIPHXAGuwGQB37Gax6/FsO2NgAqh
o0AbZdM4FZb4svZPi4KmuNeVuWis/KjO3aoFg3I4opaGHLxB3CfUZQ1IH8I/WWBjZOro6FlcEFEs
5uAsEKQD042a6DA7ZOI4vHRHuvR5cYHuk3dBpqIPDqn8rqW5aqGvyAR4nAgBUxqaW4zQqyU93qZl
ZdUS2dsbsfxrPYsN3fJsSBEdRJVhZzNPBDLLgFfd6bDl7mqjbGvebEcVzmm3LzSFs8T9Ozl/Awm1
KDk/uQGi/iIHg9WBik08Sbd0nMJ15ykJc8l6K6fdXMwz4KrEHREjoEX7jTwf5QFFfconVSpZ2nmW
cmuEwR1aKV2S4xcoTrhuDUL8khodGfFasVvlQrRK/tcrI6XOdO//RiCuZ+KNEmihaBfG+8SbkLZJ
+d0uHzWexoJQ4UDtERPPkvm7gmWDbRtUXiE2Oqk7m+cR5jeEEvqOVdmBRwRgX/a9GNH5ONBdrxZo
s5YyKwpCTf+j1rgqpoLHqhOGU+7nVrgByQvXtyYdUQgrLdfCUUMGSZWMEG2FOuIM0JjyudtOdI62
5HxiOcINQPXmvuag92wGgsjBuGH81vJdraQNEV4hAYA6/MAagPGdJMYAeggAgOQGqf5+sEsRXd3O
mKreHWaHFd2+209+gQ6ChGlisbgy4sJKjUlFr2+ec3XjuT6djuLoT91ZcBSRr3dSmHXpddHeP/8d
wSVDMWw34bZz4mso8NkF2jYTs8ko97Qh5nyYYArx+8G566DTUn6wjYCwMCr/YJZzrKzCsPnkUfXN
tyvGb5ZehFcPffar2qz14qJmWMf1M3YOcDY1cqPwjNw8U+sNNDazZVu9GHUCVFePRw6R8KEUL3lq
2KXVg+pNMMGvywRG1ixECUiOx2HawiFoRUpRxjal6JrzZ1pI+TlzyB/PdyMAJnK+sMsI5S+m+zE8
t2FoGhIQXbLvjhujCedvEhokbk8nywXTz3piAH+iEvLItrWYBWXkyBF28Aqy0i+WT5X7CVrqtZfk
KS75s0caw4BEmQMV1Eng8S7cs4nbRV3OSotU8cyYbfPWr7aNL9D+pOh1MpcTPz3KzwmZm84XCkeI
8xql+mdG1GYc93rgh/9w1zOIaOpTmF+Fc2H/YZ1kdULKzkU58hUdeoVcXCIt5t8DtMcZndP0GbTL
iW5NSmhMm6ez5BpeD5QxET9XbZVJvl1AY8hxEvYyfLpE9AIzVHsnvfBSX5JKHrK8jPb/Z6/86Sw7
cSM7kOGofQHRsiCnqMMWW0xeW33qkQZNbzsGQY18Otz3KjjHRBhEUMUBc51VD5MjKKtrGluaDug3
6LZvVI2a/bbaA4+3EJjmF8iSigdJxBU3ykDPR1vOiUhH1yrflDa4yQe+Ke26QhbH8CEy2HxjV4Do
OwhtkkAKa1XBRTlBWb8m5QpTGAfXTLJm3QcoUvpwghrIwzVBm6yfikv/IyFf0BX9wHy/RxzwFbhQ
SPzHGBGQg53+eWVIAr3s+fisI9xPcAh5nZ18vfvxxFn4tbzKSxXIepNM8RSiRF2eEv8EDC58Ao2D
5jsqfWHFTw/pCntNFNxruyG0cED93X8rMNM5Q1LKNWeXpoNDALoDaUnu2vtCIlxF/Sa3wYr4vt5Q
CAP1XrcQoscaOJF4nW3F6YIB2itKsxRJdFbIIKLG70xFprAXMELa0NPPK0xA+Yjn45hYUYZzYF/L
VqU29RVXZFDJsPoBKTDsxOGD33TQtcN3InhCvy8hx5X18TbURfFRffC4rs7xGQETgceyyKXwmQ65
2dubkDqIGG9lYrogWaf6KQx2tumGZPnIks+48V7dUq7ri5g217nVNzcpBftM62jqo4OSTFJjGRzZ
L4x7mXp3XpZft4npHeEN7jGkx9JUI8yjJrrDCmLE6luf8PsA6X7X4wY4fuURqnL4Nr9OSUmdG9+o
IWQ0iNKsAL132IZULRpZgqslkHjaVeT3uotmU8JVrwOR8PkwkQNTyE/F/RkVK86UQafKN9bwkX3c
zvM7O9eCY7veR2ZiqeCd2k9tZuEU/0x3in6J250cpEmqMmQVPsjkauAH+7OEGlH+aeEC5cZjN3fg
yDIwjbRYxWdXgHIRH1+LJPN/zArPZ++Qy8YSsv+39Rb8jYemizNdnyeO+DQ3FBPA/nuDuO976KwB
LNhgSwhTIVoDXNrZ4VTg26WvQcnFUn+g7FZftoaUHgHQaYKVnQ1MaHolCRIDbmkI62hsrVNPrzxb
FpIYO6Wht+P2jir4PQD0zRTeNBy3vBR+UjCo0yaeNtoS/jnYLFyj/SckgE0ED2enu2DnjZSMh/Ii
P9vWNuEWhVglI0Dg9VBuV+NTkDNtkDsmvQoFLqDf7rt+SX68lAHJnM01Keo3CEw6btqKMnz3XTRt
CMsC+Jf5WVsVjQ0lhKsegkfL3ShPlsWqTeVAw87K9R4HcDLVmCzzdg7kH33JSTAexIMytglRTVtb
0bGkOy/UDwOiScH5jZkfFieula8OlpxPvPD2jYvpw/W/jRzp2EqMAcBIkVeqA6rTRsKSqCis+8Nc
XibDVUX0is6NJCzEO88/gYKjnsiJQEBCbzvQNFykZNX1xyeZYU53H6fBMeLeOzhPwNs1qRmxzscz
fKfB16O8v3Em0zyGbvGKCFvEcW8idczAO28qU+y26+UcNS8BKcQWR6UXwBsJQd3WKKp8vl2qr9Qq
ep90bCxEHrUK7oK2izgPSVVtuP7F7JQx2TyD+jwVbBovi8RowHKW+5KC+oaZl4Tbco6QEGS0q9kE
mRConx5cd3uXIk2rI2cPes+x3ugyTJPPd24ybrvnZIEgWrcAwxuSLVAfXl8EFqM264/VQPhyi3KA
+bjH7vkt0moV/hl36Qo3rfs20tC9vReN02T0EV+XzSlY7QMhEIrqjNHwyemw/xTzttVDAoaro55U
UtGe/3Mh/gU5tQMD01c9/ay3BFrNLGX2d5TaYFbUHiadFHLijlxtL2sBSEgB9IpJcWcsrAy/UQDT
T6gJGiLgxSffUpuP//E3r+UGhUXs1EXW32UoSkh9f7KfAWeyeE4sSRxoVn0lKQkUAlUJ/9Qs1DL+
0dDRZhwBD9VH9GI2y+dxjEkaKBOUBvCtb+M95r8dvLdZ3D2HzSo6tIGChBitLYB2wZ2aMmUPU05T
bSrnvPktriTGSGXM8OgspM0OwZlYoxrwCeTiNIMEnIkrYXBkx74LEYzem6YHcwQupQG24NFARsn5
RZMPo/zOGkBibvCzphI/AfTMFAX+y9MN4HDhjAnVcu+C/CPiNmIBYPXaGpzUE6B+dpqKsuN+2mGP
86B7SadL+T7MNHa3a0KZ55wAQj+6Zq6ViVOoECVq8m8cGJT1oyZwrVJ0FFPysQRWq7MWkkxXEyPK
8NNpCXuP4lpYCs8rqBwyTumqZffCJTj5kBgRNoojgVkZ9klGBo7OfH3TlI1z0k6uK+Z6BeFFZBcg
47PkW34NqUro5s1tolIlkhO8txAZWAGL5jaUYwuZObDA/XRrZQmvNsG2VMdjwAvpl37kpo0mO9Aw
JpVvKctx07I8ULhqQNmguxeNFjtTeS150SYUykiVQMxcwsw/gSIoEzitTTXPvNWqDz3SCLRqrWje
lySRvB9WWHFdxnH8x4Ib4tGudUu1RAPdoZCj845OqjusiADyWL2OgXsnAEvobfqErmwG7KoZ7mb/
D+WIuCDNTRjj7Hw2E7VkwPwNyNhfMxEy0JZp2JzRbcV1l9MxtGjkbSc76pTFUr/aBabhpfvVmIhY
ciMO0ygfaduFk7ira6mNGAAl6WTK9345+lKFf3KSEi/cjb93qkGw2Huut/FefjjyaHXS6EG6UTj7
QVVzpkdeIcVY00HDu2ScpBoxGuHZuy5KrGgzvrGpWGeFteLJjL/n3GlZn9XpljL7OAols0wwi4Pb
i2wq4slmudRCzzQA2h7tagI7oal/bqZCEdTyiN2rGowN2nWa6Hl/4tBIldt5x306zD6f3e1lASQ4
Cxhb7WIbax53n0Hb0yCjRqrQqbP21/Ia60Ejdr3EpAxwh7grHtYgz15PrVkBeaXO1vYsMexjrEfV
IC5GqPwjVd6kESIFJ57A4KbPLUH8VJf7giul7rgl7skpSww5KZ+SzD5y+HC2Tkwpn2TT5WNRlVLf
xs6iyBVpq/ECt4qhX41UtjFzUTzr+fdf6WZFJjsdu6hJxIfnspsOTkzbpLG0ekD0FOrXEKC2O9qi
tzAKg5IVlXPmjbDVDrtcZVkDZaABSjkjNG/yLQGiILMFOfvZJD+eoESlGAoLmhvbsyynho1y7p1S
vzGhDPHqqXIQKDanC/oNCNWWXC/ANR1Da8N1X6w/ZZHQVqyd9iOwWFyJvhxTdi+JrFDR5TMSYRW2
xNaJ8TfMaWzo5L9YvfNlkP/HnfFm95W5+L1AdZnXtAuehMWDG/rFRuoGPmwgAApHmhHBbuU1igX9
62+YFCacEFztBdL4ijywxPNGtaYLag0qljQrOAsOd7mjuz+JqPpKdiL/FbcCnnAQSN/ZE4nEZsZb
hbhf5FEw0TdSwedVZbOzn+jVeqSpBbV+roORQBKjzQYZjO3joW+OAEfNr3jgdgLKQO5lQ4M5qrvq
m8uYiAlH3Pn1zohFrQWa16YMvqhPVm/UuYBIpMWtWNsw1kTcqgeo5bGu5Iw9hQ93+OFSsGSs4z60
gkL/2USPjz6YsA5ai5LsvOqlmFoDEK4dpf0EnQru5WhhvI4pwIrE08gjzvq4WJoIY1TuveUuq1Zf
VpWFWYixCH/e80G2C96HRobQDhZGHt8r6oBTC6isoGycnVegDiMVoFUMFP8cmO/RUjU1aPfO65UP
AsOeaGKWRcSwNZRAGrAEcQ6W8uQO9wla+9hD3eWCYNxQ2omlBRYOwyPxwUns9iTaSvYgMqYk3ncJ
1amzRaxm+0UoWvkMswfr4JQABc/xiM/26KqqTEB+CibNXdZKrom8NEGkErbeooKvrjXpMPG1+vgr
+9SroNZRxT2+JznB9bpfhPOtgB+aRsj3M1KYZIZ43B961x/qeL/Myfvy0B188ugdKIgh8Je4Gr6n
qUq979x3xWik6TFHNS5lgt6PN8mrJ6C1VfScWTGtD1eOyjPkX0lHQHV5XN+pAFZLtzIonT49ma3X
BnwXBVw2UELXBT+4ngk/pJiwNdEJH/eKG292bWxhxzPXPQF1sdBoDzScxauESnSYMujuQgpzXXe/
u2jaZhaHiT45Lqbx9bjlkYaLbP/j9pC1qgVHlfyUrkMxBzaVzrVkERBmHRRS7iZ3P0iCYryjRyO3
OfNPT5B7joN08hSLGaKqVWe6xq/OJnCTSUoPhEvrmmzo0m5Lq39P84Mh7p6OlGFrexYR7hOzdujN
XUCUlnPHHxDBqdUxF67reQnJ/Ldtr8HWHpwwtEiSl1BHxlLQ6a23lnD/19h/27D1LsbbtlMwquBA
ig5dbnBNTPdUmABRxvny/XjxhALCz6Ljy+IL1eBS71PTDUw+BG21087CtE7PGK7Q/M+W3epYOFmT
oXRZ0nKtEcCZKhGtJf4c8Bl+cGJ1OTLimQ1WzoS1gEGBkAaYdsusNXS+1aneErtPY5IQwIqPPIDv
ewOpDabtztJbr2z1FVhZ2v35F1zmXeGT6eALPI2xh75DijNpLKq11jzXHhu8aVgRZnRNPZmEocwb
ycdkVCQ8YEOiA8rwL/cxenVBbO+JePZs5642MWIXZqRf68sfmjXkV4SMIH6U1h6vIIAxd6cRxL5M
l3WcwA2HqS26xb8AVIsyU4aafaEDV45DIB529JDGJn/abjZOl7Go+DW1jzZdOv/Kvhw3zx6+guKg
gjHil7u7dufjkNGKzfNwebMJm4AnEg==
`protect end_protected

