

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
n88cX2Zddo9hCF/vQG5gWA2CsB/NxhugEioGwy8vzzTJfJgiYR1Y86uVLOsAU+Pba+vR09EA8YQL
RaBliT9OxA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Jtj1cMyThi+61jTvwaox2+7+Jwqnbq+rG0oyrMcjsRC1JqePCsMiI3RK+BFu1916onjQHte+FUqw
jzujFKMzyT+U4JMxxne1LHz0EqczECDv7WM1X3Z+/RRil6LAfoiUu4oPWKBkqJ3QkI7FQHUPjKOm
kzd4a7S7+cGdl36HArs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qEMOOi9K8amNroFNIEotb7n1RL3y9sTnhjv/DxkUSKl08KG35V+4EN0nJNAP78AeBk/MOP6lhyhD
yznQaWWuXm1lJgaV039JSSPrx9OjtMlRSRTt6chBS8kr7bfVWcDWaM2CqWSwl9bYv7FcEzgfKP+m
vX7lMhbUgVc/Xj2YFeUFZPNoqDi4TAiZZVg/BE521VWCEVBdaImZB6yZJIckyXcsD59STVUMjE1y
fbUs1lwjFxOYliPg4TmJViy6HtGYwnRs/t9Yuzd/Cgz/aiAvFIFSF8/GCIBU2YXV4nscpslh2BQ5
BzA2Jsen3nj5cPNRyRotGf1CAIloSBW2XAMhaw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
39sq6NKmyKkII6Qbee261bw7jMeBOpNoVT0bIpXXKJzbCgQKMwSkepxPD81RCujIZtWp4bsdl07x
ur1uJ4cPwQ3WcCDv4ucU7LlUxv6uaYSlCGg5sS0R4SU3q6AtD5zMxL7TAdsFgLvfLtF87pmfHeko
4rm4tcnCZhZ51dZ6Des=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
elnbtgEnpXsVV7zLjWgBzK7HYuSsQI7qzjANqzb7pnXcqXyXahPugn8SHQNLsSeNObhctj/PMapX
HD+lI4kth/BmMBwk/MLL4EEASxIuwfg2w+ukfZRWbuRKbwNmbvRGdyzn682foBeHLjeYoEtLRFz0
RMNcMFUJARCbmEyWb8MjHP22hLxzQEDA4xbq4Sy0Ik5/lMqTVTffqrlYA5jLXPboNcowAJGzXseK
nzqLTNQMaYpaoKbyDwpKdbed+c9HWR/FX4oR18IvTuUqerK95/81b7zXrQQPfjI2vdakTQf4WZ+I
GkXXmIfF6pmA6mz7wXdKA9m7FgTY6FdGqDgO7w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 158432)
`protect data_block
zWQVhrjE8HuqduSlarVPl+TiVvgTWpGnkccHbwVsyXgi3C32Z5yztNWkdujtWLbcGfGuZ705em4g
Fuf4xef/nVVCEsqDkZt4pnbLqR7B+a8d9RO35o/eG8XctlCwNXTcbEfhahA379DmY+p6slZIvBtE
4hDz5dRWC4UnNrDn2dPG1cClXokek5iNpcy7tQDBQ9elLsgoLwTs2jEHbmFyxMH3EQIBNooWnfw8
4HGG372GVNMYPsCbhleXe/tVabFwdCcFY1EDN+Wg8QJ8aW3hHaEeH04dq7B1c9nO6LG5Afvl+A1U
R0true3KxBgRe2R66qDSKWSIQwohn0OiCjqqbhUMJFTBCiwpEBcyE5CARqSqA9+jGFs+OuC4tQSC
4FdE5056+ZkehrFLCL32oqB7+NY5Xsg2z8td9d5FN4igbN5waQHC9dCubvDnNPVXkz7u7fRd3Rww
4hQJ90wYi1C0g50EPnRpWOhcY5FegsI46d484N2W4j8o76WKMA1qTTC1EpOCjm7pgS2eN2PBhixF
kIGbahp2iACgYt3iyDINYLFTGx0BcdOPb3kjlNTOq/PDg2RvVXPSuH4ECnQJe8dVlOLludgaSzqS
mikNjGLDWTMNitNvahYMfvbv1uvYzYLRgFssXXWar0uKubW6HiBCd73Y8z+ZW/7uPOZ04Q/I33GQ
Vyx+KcxT5e1M0E+99dInU+i66wCwhEHHy9YAFVmOXG09vDBKsqtiJtSW8JdmPQC+7R7dy7nZg536
Y9kemkjzIaZYwjTHMmmcJXHHlKhqsrHVmXT0g8/zVMd3nGi0iJuFO+f1+oKjMwA8CIY4heEPqfLt
9/KzF81F7apjrDKSKGUErR+me5A+zpu9A2xCoF8dsszzEBtIR7tONEiYRVOE4+Re1aeAqVqunvyK
YqiAN7J8tWcxPsQ3T0ymo8+famqFUteYKktiZc6+SjT77koRexVRyXvqYodh5qqyXNoO6zO3MSAI
aaXIZi5pDIWy1fvhdPa/QRPeU2IVqRh/flomoG1Vklglf8/OTFCxE40vgBXWse454Hw1i+KZdMVx
JJu+dpBYQbdYYMbiivRB78YSsUXklgtOdaNo3GTOg87mUnro3Zmb/cXlBxIlDs7FlKM5bwPHtXIP
/+PSW5+WDD3Xt+tTUZk0jyLrPu61hV3zTTy7uQHsT5C7FXj4KcpV3iMg5g+AQai/88/KhSvW9eVB
sVb4qmArLXrfg6JfJsNGGlmJ6DYUWc+Eg+KKhKakahIsA80Y1hMz+oFGS3ywVc5KzSLP7CTFIzoP
io79aBSxCaqXqkvh930YAr7+XFsf6uD7gFKJW41U8f9JyQ15BTVOVUnwhkYNg0JYv75fmvqWnlV+
uFbxBoGUGcVjaqzf37PX/HFikfJaGE1n/S0FNE7at3LTs+oBJiwW9CM9gtTpz9WTJdgpmnviqonq
JixANOJPCreRbKxEeSDK9ES0berZIMO9f++bpwUAVWqqjHzJStSqVtmE/ivfRdi6lrpujc0fLzNJ
5yaPrcwAFLkp3xBoXmj+KPh8eZ+WwihyT2jFIkgjIcsTnzbaYnorErgDZ/97GgDPRjn9luMeAERk
29BVBC6XK0Q2tpDod+N2HomJwpjdz/JoS+mUsmKDGFcE/GIW5pEWuOKBQBBL/f9kcu0yq1WuX8fb
d26it+mbGo1rp9WP7pmyrAdIH9b8hdgeG67RwK2uppMpoeRetRcG0gq2n1YSXbT2tL4sB45pH52o
uXY1gJU00grhVFBGI44NzBtOwrgrKhzqu5R/Rsg/CF7A8rWJOOZp6193AMwWWl6O3fCbkIk58HbU
qzBqmfdvrA2IjvWFPG/lLyRzKo9WCcjtA6pYZIpWnrkaosTFLX/R2Dp6D+qyueI9dldCk1rRjPHp
otFbaAmmkyC/k9jmU325k4fCyA/GJdT0LxoGe7RoGmFd1k6PqvTNtMYPSsrChSfXgWWw48UOxXZm
0YLJVEJiBWs4MxmsfxXHnT9It0OkAggWBBwH84r9Y2BnCiEFlgNah4EW68yPVsyEqWfit+4i3g8p
jXqzlv7k1J8Wb76z+fI7GQzfY63ml6FBhHm+fJE3aVDyUQ55mbYsOrriPeCeF2MFAxlq/FNi0und
TUSDsIlaqsKXwlOIGzoZo5IUv+SbtZ52buHBcaDNtDP/1QZx7ljBrRgDWARho15qxfwpj2qjLpt+
8Xn37sp89bdTt8liIPulU5Ndh5adsmcOsBoBU7WX2lLd52jYBXo0/1+hAoeTZ/XKnwwogI7cnHbz
WR6feeVLbPOCBUveGXI5zReS4AbAkGKMyio+qtZKsJDR+p1eHIFkLBh+ffIEhNE0f4zVzuti8fKN
sUHbHFN3iJ5PCzOQPcZWYu0UrkJDYHBGcw4d7a24kj+Rkr99rzb7Enj9t2oH8jgmCcr3zRqNv3tO
uUilBTPtxj4u+RTqExlk30CxpQLBpQ3+2s1VnGqwuAKWNzPgdezFrv4OqS+pD6At++cP4yVzlWgv
R7VFd4+Xj8nVPPPbVMCsT2gdFbjI8jhvUvelMFjUwse5JZ51xGwSY/FBCcDCaSCJxOx4SyoqHFzJ
6OOOysINANclYm1c/E6KjuqOeJIWMgSU6jFk6r84JoqpnVFKPwkRAjMKBbImT0mGbE4srAiHQ+5f
BDx6XZZDOr4U1n1Ox8ijodsGC+WeUVIfH5v/Qq+ZrLOPqyuMv1sMy7A2r7dcYNRmBoCx/um+5MkG
c/lS7534E6hbr/FrriwxRam8dV2tw/b29sm8TL0fHULIm3U2QwqLByIKLSsQPF2wVpOBEEYstBxH
LAU48i2WnI8SVVKUgFPjYYL8V7SpE1DY8hPPxMtzZ95I34idhqcYeHn66xDgZ93Y0RocevU0aoLi
wKzpv4W2NsLe8/b7KSgTIj94gyWBKBV4LWQ6KS1Vg2BQE8cYMn9m2bEKQH5c3OrunPDMCleuaVle
MymxGfb21t7Clh7F4KY7an7qnEeObl2ZLgozFRzHbwkpV0tNSAFveqz7PwYb2mkZdR5GXCehSHiw
E/Vi93KT/6C3U48IdCucPNkXqCmBw1sCfA9vAEkE2yudms7xoDNgW/H/vXcaQ/jSStKtDsvT6shl
8OZbYm/w5Kr0fWz+CQTVqsB5pUTa3BjF3bPSjsXxWCz7zaO3/4rr9sj2mzh8gP2s2dFnWvfI9HiW
PhVLO5KuLeKjnsocKDVaX3546jdUXaf5KgKCA8TNuGzveP8LnInQ2J1cA32XE+PF2UEVrK6Tm81M
D39VMdttlGz1w/V2yWiq86Q4wMkg1W7iMp5GotUWitUFRbSmVT88IWP5lw82Dm0P01i4e+OYIXuq
QNpx2qJH+JHeseduzURYVQzAMJHn1a4q5RiVHbFh+NOXX/DspZ/TQ35gx+GARxA8H1HEALzl3PWO
e9B+LZjkn1LpqlnmgehGNfk5LdIKrSuv2g19jHUz5eJGUyF9p68H8HEgghou+TqFVAo1PjkarV7R
B0r7G5VF0JX8UoYkncP2Xyj2Kaa9kz0OcyzQWnShm4Xrl0Ic8iClHRiSZRZMWSHpUGva4ANYI8M8
jQpWjD9oCT368MsCMwLIK47Ols81pfwmvZBkj8ilYcoqgLQJGddZU00JDrjkl+RyluNUZI1Z4ZZq
zuaFOGiCTRwWOW1jXvCPu+Ze5BcfCTfXTWoqIgl27H0ae74Qju9AHzjEXD0Rj0m2B9EzvJFyx8wn
O4b/aVpxKEtXLJeb1OxW02suCyeAaH2qmEvz6kL4duS+E3UROc8v3rvgHmgVmqgofK0nwKypx/pQ
SAGrTKVWXMzCTwSGSVnr8ZvXjbTuJwRjrY0rp0TuaemuhWhFtQUhyyJplFq/X8egvkqB2bg/VusX
juSyz9vb9lAgV2FOJ6VvXSTYW2jAFuJ0B8R9fBen5UB3jC8UxyGxg6r3BxW26Y4LfX6zocz9Wh6H
gczx7o2Zbm1eTcoKtUh2JpkbdtQ53xtEtMlOo410YQtJnrrQaLNhjAYQLsAvR1nn7X1/N4UG2m7M
yKe2in/hE11H/HyubJgOtpQXuFLef4zPo+OqM7rLZLMZhzowYMdiOAyOsT3vYMxZ/dKxCezVwO2k
WcXno8nfhHlw6Wtjw+1z06mLNbOhAWLlNuMdrAL0TGSFwzrRwwvUqy35JVleKYbc9vQCUMw9uDw5
6gRAy3elIBIZbXxKe7MqZO0+EdZvdHf+FO/UVeTJvNTWqRQ3QcAZb2Ig80blJ26xGEyuKYv19ESj
nLsgZBxThxi0TNpu2Z4Xy3wZcZgTDMDH9zJOUCwbEUm9Nu4IifGh2vDqRtnZQd0hCl/kOlUnt5XK
bST+i9mssbioH9rlYyc7z5EcSwQKdfb5btmeE8GDunt2tLsEi6Rtk/YjIdBdQUpZ3DCzYT6O90zr
/ZFzomdrDsMC4RBM3yjStDAmJZfzVwGHomwl7/RwJFDuilwkAYtZP3SasgAag4Ths3c3Hh46DPrI
CWLtB+vyaALH8IqVfm3rKaqm2PA5+m64Cwyraub8Pf/6AYUjylWO53Da6UbBskzMI7J8H1Zelbwm
H4nGlsRxpiP4FOOJ+miPG7qyk3EYkCGYdpIBXUTFegFVeFYr2oDGzElbbqah+WAdExoBPFwZX5M3
2hFZKzTc7w7DShgE2Dvb346QlcWAdemP65XelYZIA7VvfKnt57gck1xM1AsSxWRVAn96yKEwlABp
TIlk2s1zVJ05GTLMgFu/G0a6o5IctDElViwWpQ9LGdlULgFQeyJM2HF3xQYeAn4bpzJIURgiWUIm
AWYxghAA0XA1t1OJY20M2R6iDXQEeGouY2Uiu81REWUn4eFCY2RJX7PahGK/7Yo+jMqrctan/g6R
pFhpICkikvrtAN0hqt7fUfkZMQTDi6kkjhm7mispKhjmJ84FcqTCfuvzzgYxXL75BJJbI5SIXZlE
fdT1X6HN1SB3uwj6qI4reL1KLj9/Wb0j+0cgSIgSglZzYwD7HsWeq8beYaYcQc1lIEEvXkw9+Lfd
oOAYhHUO0U4YQi8J5T4jZ4SD4ZYxoAxoUciaT/G4+7b+VlKO/AfqvQBmPI9g1RUTJfZhEEITx4VT
7CGmxRTjokWbqWC99TsrnDNF59RwMFJuczAQpT8kLbw0zUQpOvjWGV/e4Bz4F8ppaYKS+fQFBgfR
OrHD8yL+kqfk4kChsNBgcVCxvaVeLEYiyxEPJNrSL9HJklV2dSrHx3SkatCPcc2vjIqgUB5+cLPB
A+fVpoj84rsqsExwPjzy5t1rY32fiYbBeDgSgR+QQ7uDQWivqgQd2W6M5lgsg1qLSjaxG8zmx/3+
mO0OWgAZrHEJGzV58kjrTdlgVa4rJYSg55UjmPh9OcJPrWQAVSOkgqD2Up+yr3vTpV3Uo1vSxAls
z+H6fUu8S8FtPLJ0urg2WE2XlsOvl2rcOegyc57RYlkS0QDelbpleQjyJspHPVdp6zbN+pVKq4ak
RDx4hJuWWm24bsFl1B3Cn9+5Q39VEuPge5PR+HY4NaWXjfM91O+B4TzH/TVEzS6E9sY550AjY79a
O9N0F6l2DyKOWB9D3uUnfVh/FX198RFTB1Er7Q3eubP6TNMzj0Dopq6XFsk7AXItMPJKGEhaEVwN
iExhMgrAcP2DChmmeD3+8PIdcd6DL5kfiNd/evCyxp/s10CFqhD8C9K1BImwch4T1OTN3BkN7NGe
N0GjHBXoL2wVnHd2ielyPJgPjUHv3B98wSrh9rNyPoOJDwL6cAio/ifnx/lIMfNqJYlLw+TJpA+5
OPPxfDK5/wqyMmOJU5m9SE3WxhSGZXxZ555IMYIYSbj/4nO2TFZ3ipdlWQCWnjJPsLsKPs1L+YCG
yx+2a/yYkkBemsfDPd8o6k/1UkbOViN5Lt8MaRgY3R51vl9coGdossWH1kzLUG4W/djTVQ+rNjZ0
CBUcbK4HsE/pSXOmI+ORH7D2wFB1xICQ5DfTnHhI5ntNW2zgzT/bVwP/P/KlL0l+zfzHR+VugisE
67hE+qal6cHRlmzzQz0sf4JVoaXJhRUk9ejELOl3uW8gjgeVb3K3N5mcNYcIQIUmx3GQp0zmylRX
w6xs9wjjEqXh7rfL6kCgY2X2DZL51mzzmRKBCTfIsEGry4FHtijP3TrZm/bJ+mKBcOnhJxjzHD2e
b4q7vIOhGvD7Cswub8OrOg3aBfzNK9J5cTUrsIoHOIAWChl7vWpwnZbOHmSxQ0qE3pkrs+o02NPG
+mfZ2w2/wq5A4KtHsXECLNvi80Au444Kl9q8Tq/sWcwJH3Dn737JTZdlDpYGEaBzCAUWKHgS3jmv
oe8IMC37PZiDZKSB3O1unIrf0Q3D0bAA8r3HBo2QugIX8v9Qhvc4/MZUpQP2M+XRWjvl02J/ZrMj
f+GYTuf79+2/mrISA52bcgCXmJYmf/wwwLCjk7Ubi5AQrmr8FeanQa2nLL5Rwo22cFaq+Zy8B5+A
csYZm6ardmy6RHj9EdC5vQnAaiY8R0PIaMPt+KkZI1C7+1Lm2lwrbzz7KAWsYRbvwFhGzeBW+ZdG
XFqym0OXDHDtpFsD68cTphrX1vhmoE85WG8a97tDGzpxXr+s8Xt5uPavnglfRNXRrF3lZXUybC1/
LgpMh8a0IrQuvTPT35NK2hcFi1CUqOM0I2vxuoHyHuaDen9tFoK8kSi47vb3/CaRMFXa72JIU8SC
O4+eTjm9Fv9W0bCqo71SscNkhVDZq9Z3XZNHMtUs6SphBlITTC1oJa2oF9DW5puq3efnR8M3OEnX
ODZQe/7nYjMucHQsuFOdZShRLjoYicexffanBVfCxpoXCl0jylLWVDIfms9MFzUfp/6duwY99ESF
WbliLW5RIMPJe5ekgMQQCKdE/qTkrnX/uqJGkOQ8dhtjk64WLL7qSSLCrtDe/aA4Ww9EnK/213bO
010GZznhsPkSHv0/wwqHwqX68Rce4B3UN/MotP0u2sNIsTCTgsNfYia5rxOfFdk4i/dZDM7tRU+u
c+m6gWyiH17DhzP02RNmabqNL6N0wBLXQQLmv5QXYZLFM/ta5wMMLmySmDnHeaGP/ky+1F40Q6y0
YWacAMOFU9ieJtXC/2JVgdBYsg9h4/XCajkiX/PvVJNMUKFCEZcMCEy//ev4+HogrSBam5YGmrXC
a7VaoKMtavr76FMX+q+hk5B22yNdJ5gc6kDakeZ/2gkMMGbRRlGPqFrbTVRu046p+MpcbDq1+/Gx
MpZpHioan3I/eYXBEtztWZVyBlKQBCbB+2naScllYRZRq2fwDdeGUyIjBYRTSV1sFKjwtgD9PW7H
Ec46I985NOmMR+wD9rkSyeGZI7TNVEEkmyKyKRg3+zqg6UCCnZFIlMvBbW7Aqr9AJJ/wdU7NSnHg
JDyoFEnpe/V1ZtL7nqLrJqQOO2XcgNdpOdObWZiw4jmoIrKDgg6BCdB94Ub0//T0XutApCiCxA4K
RpU+wbo60i0NPXw0ce23SYn88Mme2j2hnNmPQnjCzSrfRwfTtZDpnZ4TXY+zA0OzZSmnh0rSYg+W
eRnBLKvr0O/lyVPR1HcBZFfV1NDKkWb8Mj4dZoNeFbltQd5u6IFpqnsbmi1DM/4UksNv3XEcJHW1
piaT5C10hk0DL+e3qtR4bP+nHfDBgQ/K1Lmk3kbEgkMWGCpfSn+g4ZUENwjxujTC/w6dCJSTH633
2MODuy3fRr8YESiOtgrALtw4cuKJASPkwWIHyXmaijnXLWe3F8v3pp/3evFMDie6R18JN0gst5vq
C+9C5bSoZk7OpKEFVNAHr1V3oZECHspmnxjH+uh1s6m76O1wHwcZ1So828YcxCbxXyTKaolDCgHJ
aV847XzZ/qaluyIIlODz4FBCFENYZGiVHCv7qM/6YllmFS/sfUcPT8vWEvg0bO+fuzUorR5vjNFD
8hcs2I78tMcogOBR0kSAVxh57S6cmPVkr6gPA49tpN94YS6ngr7r93IRaFgHiMKeBY1jEHL2HBHH
w2MkNsf8ky3eJ90YdWm0WA0l3mCMejzeoj1icoacQ1Ojk6SN4IH7TrGdXJShaeHGc+3mrchfJHB/
KN/bq1JRn6qgoYezPZEyhzRXeNBvpyM8kJ5LqxxIZep0ZDUXUJPaR8psnpJLDKnknr4Mr4P4JkZT
9Nqb6HYb9OM0iq09U74LHriGvRo2y3gXrABqUMXgiDjJXjpd+lg8ZRsqamhpNH0krzGr/gUg7dSv
TUh9m4+1jIik4ITsSnLeYSyd7Bq3vXVBeHNlw9ShyxlCkUMLPPG0h+EX+FYm+9qxvkgQuVEJebQA
H3i0eY2g7vIaHCuBZ0MoS1nhm1qsfIMrmOoKpIaQ8gmKk7rYmcJExSahno/Tp7zaC/BWBRaL3tej
2KlrpWsKNtZMbo+tym1yG3r5nwEdRkjN4JN86zrFYTr6jQrWPVGugYuuR4V6LvELAW8BwNNMSC9m
hNx8wYLVbb9tLPTRqHVqoWlMnxi9bhSu0ZFyT2W9N/IhytMML8Bpco91sAT58J5bbr6eg4PB/4QK
yKa0JvpKx7r3DTzp6Pycq0Hd3z9PlxzGcBs4M38UwJXQtkoW2SKJQ7qejLHvF6FAwO0H4+ClaTB5
Np4pNYzNSCpFepubkUXbwTbDDcx2k2q0tUvP5KLg3CEb9bTiGUIn7ua+CAJcg5jZv8bX2Ce+xWRZ
avUaaAaWbF3oqar3jepY67ZzBtma81rqQOmw4e0xHxOgGcFdRw2mggbre0+Cuf6y4TZFPUUnAEPf
rECGzk4dmOEUovFcLY/foiWYTtCr4jUXVlYi3saCGXl8TkjFKsxu/rFU0LPCvgegQkgp67P/Ysg5
4zETwpvsi25lRJqWGlFPZfCUW3iC+GGq+MT46BqBLI8K94hu7/B1o+Kt1V0FTxUfsBgxlg1wxe0c
KhwD1gHcDMHdJqgHiOZlq10Jgjv/y7Ep1zA56rueD+ScAvESzKgF/fmybo7euDnEQE6NhJBlKBNM
PjROoe2bQI7wDOH1A8UV2pWgQWts5I93wywokUx2JIJjFzT1EzaJz91v3LG93JO2AicxMU1t/py5
hHzBK7Fp5SV1XnXFIgGx+46ljNfB5B0ndGxFNFy90PKc0jXtBYZtrKC0xaNW/z9NBw0GHKSIDP8C
bdtpCr2gdRtkyO0RVymFgJn0iJJ4BMRBQT3mwucNdguJr58dDQbEW2DpZy+YG4sWGPEFvg6H1OIW
dG1YGU8NHMNyTeBb1q9CNyDc7Ci8rdF3a40wZs0SY1+fseGIXIzVqODGmmb4rqHZNUL3GGxwuBuv
EgW9TnpTS3xtyPYao1sTtyYvTpeCHqjrdmiSsm+FpMDKtuqY6x7IM985LiQo1ru5c/QDxMH6PZkJ
o7t2L3a683672ud/uHR5kBF2v0YZ8c1xocBgoY+FpP37hd3o0es2ieTpHsFkJEk45iJWnITaYlSr
zwmaXb/UdBq+54bkjNq3RK1NNHB4ZNfjo9EpSd2JVbkJUG5POkt33f/5WugMVryeTk5w7NR9tCvB
Kwkvs+MOyclVotpAgKng4pQo7gFVcaLGxGxCgn8uIfqmiUWuj39uJydDHmUykAb4UJtVESYmEMMv
ErL09AhB77koueqjLl2xeTkkC6dv41heg4YarXCzFumLItYMzB/ZYCSSQi7fIkai26vJSpcNqT8W
fVVAVQ1qoRy3OrZQiC5Ny/d458SYeiZwFWH6fsVE1+it/7bvs3Xl1vd39lGvOQbYU9NXu4vSC3SI
IENROmxLJ3oBWDEUKF/ie5wTPHXUf4MVdk3KHUq1VmXQSJTuVS8n/4HPPe6EagVppR9Pgqo8n0oI
UEnQ2OITIPZy2C0lOMfE370YAWREiQBrq7pQYk7I5N5bt6vMmZUNAZ9ckHuQW1kN5nWz7Dm/ROgw
gm3/9QFUmoOTsJQWTAvm46AsWR53vQeGRp9ASsF+fl9hub03WDjAC+iYzcEZLWuOGe0JPkppOw9Z
FFd/d9nqq0lXOz77CQlNus7/vZ3J2krfWsPQONVliFMhiKYF2DOHytBd/JT4gv9wNMPaYYWo5kld
+B/f5oJwhgfV02tRU8r9egsg/FTcCorF9aHEsxa7t85rIi5XLFNbTyJlehYe7u7cot1mxfmSYseO
/UPZ2Zbdua96mKpPWBUKnDsmPf8Vs3dSRJK6zbd3rZMncojQY74aKWSA3hdJIK35CkcgxHxUhyRe
4U6YltWHsmfiiwuLDZFVqCEwtufwsrcSHKPqfgi85re4Zv5peah0kb7SCzPZTnAcyXTd/6Ma/LKZ
T3kZFJ+eXPFoVk7f0f0LiAuxCtok9Fwi1vVbjhEKIV2uKIMIfXWllCewFGbsySXHPQl4rSbPBgbp
ch8BAIHrh9yzrb+THMSE8nFoCbArJrQ+d0EObUR9YTJdidnrqz5YWRdYQkPn2hCZkpPOy29xR4s/
cIpQ/OYn6OQISGIi0vLK56ZCjBZZ3aMG7FEvF/GW226wmncu+8EEmW3aEOsSMXwb88+w8tZ1DVVX
nIwXFDNCfCV2g4tXcAxUk9TEfTgAo7sSZTxjFgpTLu1qQo00BKEvZmbNFqGoSZRjXorKGoZWI08c
l6hmk1X6MLpMtThNGAPcJoQ2/K0rK0UW8aDTF6U+zgvqLfSUfePjPEPIt8JdsVpvS1gwPZNZXM92
E9Z/zatRMot81Ib7aHRTjfb8F43+LVx697srR3W1YEKhraVDLQA2mAy0MLLwwxYxyeT+GOhWfmoB
LDX28ukMAjQkq67JIHu5djHmKpkoJPagrCf7OWlUq25PPOvY6Q7vavL/2W4YFp+GjUI5utan4Qpg
K++vlJPgDheLm1M+XqNr8vOcMNTM1+2yNFCBWVTrzF0bnU6kxwp3BGEN2O4yqs5fJplD4RpuyD8V
JHyupWS5sY1jHQ/Liyfyly6lbKsCKjwOi2kX6aLRrb2b1hhENktgRw6Ygj0uf6SwB1BTq1j9BSbf
fkZ6IFfuhQlQsHhsXfpk6NSdqZQmgC++rHw4lZ1c9wAmpOvV471LxgdLey9JB5fE+8iiLKMEmbJe
s9vAWMqWQp9NAnmIq292aBvDQEPnSG7l6kHhy04h9Xukv3g7aamPFTXTJG6GqJGZKdk5F+0VM9Hp
txTaXhwm0yWTH5GLPPQRprjMxPdvRnRjf0O2kD8OaOL6j7erherHsbsSVwBL7qHsFmtzNdURvpLY
GeYft7+Ql+RCAocD5B7tDOxKLTde6cGE3SB/a2D0ZWP7ip1PJBFCmQcyNL0ArYxNUGdjFG5AuBnZ
y2eVlhNTsUz1QenLUAMf1OsjCOtPX+Ppbn45DYYipwhJTYTYIi7bP+Qqagkfb1eTxbTq7q9bPPSd
6etiq0DAzwKmY5YS5Yh7fGouA36ipCvXIiDT8fWcPq8m1O4IQM1ZNrOQFWWu2Un+aO4IJhZCfNvb
v7XxHHowu+ZHRhqkzgTyT5JzGaf+inBF0nAf/4a4O1/6b/hlMw6sFkCYnVjXMN1R/B7ndBCj50yf
eyitMuJto39OOKSi66K7BAQ5+7MZOjOkzVS6egrcC/byxgn/S8m0mzmLQ6OPI/+n/mouaiefKzVk
tPdCRaScCGctKZJiaGQNvPCnIi1T1rE/ccsYNsCejJqZiZyAQWACFBtsBMxZqLbUAyD9qO4zS351
sSMIr1VB9GwI0ORznW1lE7+QG585m1XBUpukhVtraCmZNaOwZuZjKm/VG3AZDxpbWs7/ug79vAKU
Dr7CRfj7TPuTG8lvW4u7S9SFQKz38tIeQ26H0yz/As8kpHg8WzUvMa3A+8y7lOaFYVvgDYMci8qV
+GGQsFFg+7lmn9aRzTA9n+DxJbPVnMp+B39+bak8BLojc5QIMP9PTMYVCKcMQpvGmB9qW2KGHFgY
jdffrz2PEWrygOTBFHWsT6ajOjwEdJ8CKj/6V3h2u9n12GaAITMC0EpkzfknhflpAD75F9cUMNnl
+LXLOtL1EF+k9V/G28Qvz5eCZ/WEzvuaIA+MjV1elGKCztE6G/NklPvv5HwSjAyIq/teQbsc1OYp
AZAx4Y9QkUc7GoSDIX17GryFJWx0Y9O+T4uNgLdRjAHL342tVZa6av9Uce07InzHta1pZzPO4t3y
5yNMagCwBlnGoq9T3vengfV5GNqASd1B0LtWVRz093x2MeeQmsAhKUfWDuBlBLSETsz8O8OlmXis
+58pbcdHZeB5/AfIc6KKq+4AhUqU+bkTjYtuyD/imf5IF8xKgmHZpCWjRC+lKPerPXLkql5usCNM
cq4NUKjXLE9AfXOTgGrW1BA2OtAV0qAaVEWDZiTlDVP5lAnlAH0h3dxfDlQTVTu9paI74dQOBodD
w0itPgnVnQMfbeAxaMEx0cFS/o7Qu3XP6GAC5se5SFt0PFrB1O4wtTSwM3Cxu6QHg9LCW2pAaq5z
EcUbZy5HzLNW0jK069M+G0/yQHru9ZP2JTNgGZUraCzxcaGwaDdrAU0rwtX8h00e1zfsHezf7xnk
GoMSaMGukiFNuzFJtuLbkMNVhdW0wmRcbJ0dvN7kBwTI1zterS7EGvJJzAfasr5+IeY9s3Fn8krc
f7ehMzJ/lV9bt4sAjewZpqH91X7Bbrtl1sdKsiteuLSIW7rscQjPzI08CIyINisdMAxHgOPY/y9b
gmzOIlTNcHo8PcbP7VjxOKVkNgDRZvQiR57B4FMh4nNq9TO5xE+k1FK5bshPjthPrMhd0DJV0R59
/ki+oVTjogoWqwyrJx7nucNXqqWNf58cf3dBT7IMGL5g9Ro4iIfEnLCPrmuL3nGsBbm+ipXBs9uG
iqAINUaPHzvzQhkeSZn6C1IPVgN/ZlPyB3ZYJziCN3/D/+/i9sCTQzsQXIF/OCbGirh1aELI/QEf
FYKHp9g50LdiK/DHjLq6WDF9yKTjmR941LIaTjTRFdxy67JbQhzlraM+UW+PP+dVooBa07GqONXM
eVPzGUBBHznkKLWYumJP89UmXxxBvneXM+MOLm8f/mteEg7OGECDgh2J2eSVPkVbZtH5VMdbnQzM
emsqcUyeeikPNY1jbfJlqOl/xgsR83BzkqzJQG7Pahc7lXxMdkU9qT2uQNwwNItjG6Vu0+wX2iJq
d/QQjhtvFzrcRCByKrDU+NZhJvqMPhiooj6I4RNLYaTZL4s6HUD0hHiaStIrWdpc4+d/eE0690h1
6uK93JadLdQyzfhW3MANfr08KKGXPVAB+HeQpx3msv07P9lO+dzsKpIJsU/mBgOmEwn4FdB5p5Fw
JMgcKnKhUmEyH6jxLxUFA/QOKiiF0Qf/LzZgDAHeftETy0EFE3XO3txdoBRrF1ZJblKIJ0YXY3pw
X1aMyKPcrhXBxiDzJsyoK3ov2B7MCCk0oVPWFVgr1jRJ36aE2MxMf8jXpCG1DHwzY/vN26YKyEyA
0IWwJR+zvE+OBiKMDQZFpcBXkw2lx4xXLP/MmTvjPN/aFQGqYt79X3PtNoOo0hP7jPn4wIBCWK0W
auHRM7cNl1clBuoiquVfz2FnTvH+CBkzBvXlqbiveBJ3YOgqu2z0+ekndpLvBLGL0WQZJ4GEOvE9
2iEDq+5Hp6kaDla6kbfT/8vsh7kM+oZ3i7G6dOClM7pE/LrPhUoV58iq/1TzqWOxtXIs3qRwFBlS
TqX9fqSZA3hvNJbNKiaHaR87x02Qk8kVskY6uUdxkTNB2UwvvkuJ15TPNbUGB7vTIIHicKBvgpVn
9iCURiR2AvVWJJcFgcFRn5xaKI1T5yi5eAAVdRfkYKMv28UoIPT3/Rz7NkhXXPcl0dnTcndz9lMb
82MFa7nGweZ9Z+OnEQA/XkrqqRZJqywClAloAPwrRXCzFKK6ikzZ3ao8YQX49HPX2Qywvzv422C4
Iu/8IIWc6oZNqPY32RiwncN+oGs6W2XSJ5xITHQ0EILHyO9oEgx8VHyK6kCHLS43cv40SbBvRZo0
TdKsEoOOgQeHreGvzSTBUdoS6cHrDuxkZ/b8g4IspuxL0YuzfJgonlXGMSGm2TB1ZEarbfDSaSTN
yYxhBd/bN0i8cOodzE4kZ55u63RQr1cCXpX455XPeLANWu+MbqHVBTqbkNGfVCRRKfvuEFu7Cr+0
TIm+GEKqOZiNkiNdlirkCBYLv4t+tjG3PDu9T0JzRC7w8/0HdPR/Bc4mZxCq473UgGoktoMI7fJt
udWSS6Pva6pemK1HqtwatjJj9xEP0LltIL4SEfeocAB//zyw/jx5o/Sv/J3OJ0FuEbDijeruttom
BBuHSLiOYpVDEnAESaYDJTjkDczHMi91EMo2856+kfcgZvz/AzV+JrTLohvXU5oEGsWOgbgEgnIl
u1zd6aTBnQZuKK0tcsfRD9sarGfB5BtEUec4tYwzTbSgRdbqOavuaud4H8orNEbZjTVcf/0mqFnG
4b1oYtxehpu4vmm1LCPFo3ZLOTYUEUNSEfobg5TLaz8X4gUuPzdJRWk7cb8e+xZcpatl9YW63LS8
HXeIiNhdIPwMmz/I9d6dmfb3n7hK1ve+A/DlUXcgRHLzxDGo1j6Ibg7ajEC/spzcYVgrstSUPk+n
DX632sA2dlJZAcT9M83GPmMzN7sol0lx2HNNmfVsTxkaJVoM5k9Hs0J8in9JJ+cdV7m/g97D9lG9
3LJI6Ypmd5+GufzlYJEQt2PZEh9FhXbJDTVe+HD3HJqg90WyQ04OGy9iC8qvIGb3DnIUKKabE4MF
Ka9BL9yDYSW/YM7IT4LPiKSJN9zkgSKb0/yXz/ohIILyeZzi2bnGM+MiFl7jrmRVo13uobJU3Ptl
ejLoSh235jC/pSYkdPuSsR6W9lfhoQ1sLb2fEp3snvMpZwXbqVRSXahIO/r7kQNauDfkNrmF4bxJ
cEtzuVB7BwTvVups70c8CHCB0aeKtGzo5NXY+iMByQqvZSxCheqN1/csyYZjWowAAMOlbLMED5vp
zUP9g3YIWc4QXbJCRpBd61FFAzdTXk6epkcZTVzTI/m/SqTABzaNX3ZF6WqCZC+2ce6c91Lq+CQF
Y1GJcbaQgNB1Ft0r8QdPcB/2wWybwPnOhmhXUlAdx6oqPahmowoMMHBMM3/goaabTP4/hl58MzeV
ck/JFSvRWUDCZXNDxFy+iGwV5gpOLwggygQouNARaoBRrr89DxEwX5yBYTAP+VPvpktwPWU9SuBs
A6xGpadsPse45Z7EbinT6f81VDqnbbkkCiEp4mBgSVR2wkRwQPpg15IFyy9/YVSTHHy1kLBy4tiO
Vu8DfoP9nmeVw41nPyjHO5976RM3YK8kIRZieK49IXPMa30wCoFGUrUiGkNwkEv9AAhep9zJkETE
OdiCx0PpBNGfZfZhxYPzuSV1NR2csl/shbUKxzFBKH/d6RXplanMx+j2+woiRPc1Q1UAq4z9hh6V
xwZmNJbmTaQvxSJuchygGY5NTkeJMWeEfEgnmntca8Jn1yc96arIxHUIkZ8ueSUpcAaEk54CECdD
ep25AfgL0COrhpcpOYoeObWRf9sgJl8zE4YQAPTgxSuyKb/Ht/hShONEKiE+jlO9qIUPi2Rg8fQz
c2Q2RSB/4gy+gDaLtfFcowoXoNchWxkaxR3QsGy2FFlTXPI3ZXuMvTAXS5T/w2NH0DV+oAB+3iq+
WbarIABRbsQJochYcP0c1vkX+3eloLm0XVMyp5f5umZMf24RDo+flQKnaOUgl1ra4P+68Fxhd25u
nUhUkylv9hxjRBt3NHEIV/mWtPAUrGaPCtUDNqsM/2SEcX1jk6aB+7+FNh57ebZkuj+1Ld/BLQ16
HjtR5hMT+dm0Zt+zcj5JeoLg304Fx7a35QimlNmU/iq06NZj94GlgmeLMJTEKr6euCXvojVnb21o
CNfMmnT3SDBPFMQKTXUGqusI/hqicAByTlcE85iHsl36iwaX7FUsJdDXAa4FFW7WabAlWy1T2tZh
1Gebz7E4WITYMEjKsLvJTkw3sYLb1RtlNkpNF4Y9m8UrPjMbpK9WDIO/ijHp0WCFAX28br6+uIPE
xthr7aoJBnTRiP5I4goV0lUkX6RsbOmyXP+RrKXn8N+HxvPhruhnXHxCixYVdrykw47qYkiQWKrd
L/UcaEo9RdosGERt8Fe/GYu5aAB0L3ecw/p1b7WOIWJSmAG2B9rnM9IMRSN9URFJFkX3ZLAghag3
MG0ur5ofglFcDOagOYlpSn/5dAf4GzMy3jAxjjbOn5RhfMUibwSR/RCxcIErp/3yQGyowVHUjvas
l+EyCPvmZ3xxlm+47wMWmvMf4blGZOgHCBNpRcjNEC8wfZXr565JtC6w/ISpv1bUAWn+p4IJRe/4
O+fvSA9uucPx1DjtXZsPK8tqobYFoS3BFn+IZeBuDegyMwPcWghiDS0iSLEieZwAbLPvjcDfTnR5
PUqhsW0mohHobrTWTY8v+DHv2+JgDSGq0o6FBBelZ+8mf6mBnL6dqtP3D66zp0bihDS9wI+MQYId
vfWQZq+Jbrpok7/51p+9SrXwCma2/W/URI/y9bfoO+C0ymgEIuPW6l0wMPNvJVkDKQViU64e4Zx2
QvGKaycjzOPbv69qMkcUqrgBV1BFpfChN7MoPPhDs0K4nM9zmUTktAVolLqRejzFAZ1gHbd+jBfx
rkthCpbhQKGe1Vcd1UHwxnfgi2cRrZ7Vdd9SeiqafAcbfWZdbUX4AZgRXNncb4fv0l4InRp1PBHU
tlMo7ttMuAk+0ChJodvV8K/JbsM757ji46ZEx0Dnb7feCsxlANMfKBnJSmH2N8Ob4ru0WgcQwpCl
XiWo5OprWgFy5ZGSePeRWKs0gAJJDr1oD3TOpELdYLr8d+r1wT6VQrTHr/F3x52j5hyS8JaSdWG1
A5Nnidm40FlLndJ2a5neBxngn5UieISi2B0DIV/x1Ji10wGikS9H/RFC3z79LEOlpwqpZWGmAJub
GZ57G4ZtJEloPZ7sqVKeXoTrQhvirBVTUOmhc0YrvMiRT1htOukzHWMEF9FIUF05S/5HPHX/031p
JOSbbtAXeQqzwOuIIZ47FhwEqKqnN+QlvDaS8St+zAY2ggWqsYTrD6rRph+ldqBH6V2eRaDKYq6L
7W0kcQIgb2cdJzbHjfJxCBiK0AD8oBHirKPX4YiM2aP/C7TRygVTA07u85HwI0GJyxB8zgKNVPRP
yHtVyiqF6AtCrMpuKPBixEEFOCTCL6Odhz9d6b3NpqEzlWp2/1EE77FC1i7dTIuXTr7hZIFPLeOS
4b/y5AJtglARbPIfrCqkDmEtEziAX92klZ/PCZgoRoFBeAL0Y0JO4wM7V1fCxb5+ajp9XS2pLqZH
1rC8buCo33hhtXH0FbAUjdM1OKXqcO1qT7p9R0mQyzw0/bhdrOB74jWUwKngt4gHWosrwPGZzDWu
K7Wx9jjCM3CSAbp3SSqT+Sd3aaVQCbLPuwIDO89TilINsZXe+X+kqqaGU25XsZMu88UXs4eKMRld
QRHctcAE5XW2jOyq7obKNvBy44M+IQdTZYFiMq/1FvbjO590gCSvzftXfiKQZg3sRcEJgDTt1zEO
wuVeekGu8M6wqAu/y7zEI60rcoBQ2Y1ctskLyFYkWwMdtzh6Ng3sbA83DxKe6OqcsbUU572v0cWg
6VHoIKRJ0hg1DoKCiAkPQw0mwLJEspvFMMCA6pLwHSlMQlDMaXmyHLwE6MUYJ3xk497wWtAi1zYR
iCKb/qmJjKAnCxXwnbmyt9RXisACuGFqipHisxlCT8Q9lc4UxDHGAnPeJTv9yYbew76T7U21op6m
NDbuNzc+m0XEQRKGThc1K+uqrbqgvl2MYS7vfZnPIXXhi64FLlzmlJO4Qj1cx7F/0PIueOgjH9gJ
vlrrSXrHoLmtferUNv+U0iP9/yiWXwLzpCzfmIdlDfhrcTIH88rpLN99Qi8IajQ33+j/8bSxWNqv
K0JndiNKW5X96kxb2nPdJ00U5mUxJv9Lew4aiyAsbBoac1AFWN2u/NyEK9HlvW5jiCnrcPGBhGF1
WZ+AtDiZDDzF2v3IDyk2vP9G+5Utgwuxn3sO7+FAUe3R+RZ7/mCj0WT/CCL5WCPnfUUreq/4AAZG
9BLFeHnU8ys3RYpyhFMT2KSVHA/3PgUUFY0G2rrhMxsVcZBXSMyjfxlvVSMAgI3F912VJd+ipd5v
Tbtpvm2SjMjcF6xFihGLTim3qFszxM9r6unCrnLeNaX4w6BuOUniJEVNgVe/N3ws5ftaHhIVKc6Z
4gO3rrVIQYLlGr+QL+FjTaRcD7xQSZOfZF2j+U8DpJsSZ0ckGiHiUZ5OgPZLkeYjE8cYATyg44Ds
am8U+qgRIzd8+npNE/q34dux6ZUsAouEM5+G5GOTTAvoKQ3fiqKwYLCbDyB23luyWecAFxCMXhI5
sFZyMIhptbsQSpBFfDQyQZZ+earpNtednd0v8i4gH2jVO/feSRYrj/7z9e9nEabwhrVji3CLCbLY
qa3GCDDByTrqmMpu7jHQe80+miSZ7Bv0HEDTJ3oYlnjNNWot2JVgrKOPclKa17Svk2rPySEZdqTV
ZvKOKrWR3rQwsh3DKI5bL6jTu83YjNgNSjk905utj0pKdsWOfdJQLpqLimCLBQ2SOyEU0yQx/qLF
sXzCUX0j61H/USzDWmNj1rjCb8QdOArtOQZ3OkwMmd4rda9T2fggwg25kLew6eT+/iramNRqAyrr
kc44d0gTO/EjRP8/gCFcxaxApTwQuZN2KQlmYncbPs2iR0LmdIk7GRbQunEzZP7RnKGp06XWIimo
NJ+k2CzSbmbsrQZPubF+A1gpJPlN30oDPdb+U7pKpYTXJ8nlzJo2tcJAuZ305PydSXy4KALdGBTi
aclsv3Vl8D3+ryOvXNvA/ZPV4adr1ZJpAJBRmM+k1p4yCbsyScnYhRgFjOUjnjTYTLH1LapVVf6E
mJfQqjJyCiXdUwROiT2kLJnCE/YjoTukYnvFh2Bn18QHx8NfNkYqOPDfx1Htz/FEo20oqihv0aJG
dzQesn/Sb0sb3rx4hcD9MTS83TSmB/FO05OkJW6bwddFbzaoCTLKtHdV50+KQ4+QwkNNcLdzL8Tu
E254bus7uqICmOC4CPbzeT/7FqAAg1l6R9Xx3ZqvB9UVGlgZO+y8h9p/O4VE7xlxPTEkLkDfiFXp
fWlAVV9VbyLu7N+UGV9HwIkaKE9hZf6TiqxsWDMe0vK9Q57kJQavp9W4RDdcKF+2scMtzXk+rhIL
NXrFbLEBWoDJ344rsWOPwwBI3Vib1MWAFe49q5QoDI/RJJ4kxCD85Dq/gu+y6pQycsrRT0If7I/L
k3e1eLSsAfWPE3Ith6psNGm7BSEVmpNNo98EfAMF56pChZtAXpONxUqQl+gYPwja4znkFA+r1d5i
EUfQ+jEoReJhIaeptBCi3KATtALrTAvov7eIq7Dt8aCa5/YwEy4gLQbv1BdWcmxd3mhyz0CJrKRL
tWpAG1ud4Hr72JYfCkhY5wprDoDWvF0+JO2VD2foUAgcprScvRicn1V6dP8cWc6igVSWnZDtUqfv
54yl3ch8XA1tjKunUxKpQUusO8gECqjz9fRQykvBi7HgY0UByHlNF4bIh9TRATUlOfmom/mpN96L
DpWbA21ux/5vTfgM1Tt6KkqNYmreHTwwfOsFBeJp+T+MCTwfTkSAGwKyDPXExaZ1yZRIwOt2EN8T
07RuYAc00Ten3COZkSSbTbZwxDFV+Zadosd2Y6h/5pAHfqfCcmQQfDxGizFVtbyhl0sR/PQCzwUz
TkwSn45P0HjVmOX7vleZG5Bw2OycVvEB2g7NQT0vMYB3VzCjAB6g+s8LUtpcB626Ivmb+4iRkpmZ
5WWbNPyXmz/xyQJEQ3RYwmAtJEpvzLaShGNtBtzwG0ZgiVMWtXgh/XtcQLh+GTWUfq4F09jtCpDY
6rNHKv4m3njx/mZj2UM4xmMZEGd2RD4YYYngZWWpYNnTb29fFKxOGYjSeHU6UztccuxFwkTCyJBO
+jy6kSJxPEHH/wyQeLTyKg2P4KliSbcgeCE7tbHEnbyyL/DwoJ65sUvE46cjzDvHofc+Vm2b2JwE
pNuAY6KHCj7ECrM65WbcMPJdraDVnkHno9k23FypJ9FiKxYiba5zFaLuGpUS455Boe9pqoARb5G+
/Fei20yRLcBbffYRMt6aoTOI8/INXGaUVZHaUA0DjsbSJ+1T0uaUYvsoghzrUsG+zh2tOwmW1DqU
RxWIRTTBwlT9+BiOc7cryKehTRmNkUTWJeRWSxmu4/WtOeJVyT9YPrsBA1wqj+jIC/E+DIy+M+ap
Wk0M/510cFS6dga4iWG0dLW819x+lvfvNQW8NaoZI0ANIuSdWXCXfkEkGsugK6tlui9IOqlSRKeK
9sn7/7fyhpMeLehstMtaBplGoyqvjJQJCpNjmqqNK1yaKpqn9126h4hR/DHmtC++y0Sdb0zEC0Wn
cr3n/6jD+Z5t2a/+8PEBLf3Ru+Vl5DxJmvluQ8/ESrppE1wnROVS0b9pg/CUuZpk7eos0VM6p7LE
wej28hwDuSg9aLfLlEfRwMm1dDJALgVqyZnt7YkP025xT/OFz8Z5ebX9IDCAty3TNSgfvh+hA9Im
QsZK3ROf34oPtMSFG4Oe73ZAW5+1nAMXAeGlFmWRYj/pbevYBK3dQ4VnVliRjhjyyAQ6VOMXZsJg
1gFjHdI+UK07B+6QndCwQWPs/+dzV7NsrXb/7hB2yau4wL3TWe7FAtE5Ov1Ll9vtFYc/yU198K+4
WwpXJkQp3Q5hROBO32bV1ExO/JZT4mQQkGRFoD1GNu5Uy/enWsxzSKULV0XFbvWYp1U7iQ1m/SJI
debpX8hqc4v2SaxDy7YXZK3uRqCx3YDzmWXHzzbByQ5mq/w55PVFlpvftsTa6NTArd742mtlFUfc
S9xjnXb3uE0gK4/RiFoJLtdN3wjQIhiAraHZCBXg2PwUVH8IjTWxMdCgF7/07saaD/Yus9GZxX8a
aV0/+1b6J7OYaqvPMjnnye8jisxusbT69YauTppmKDKQshO7K9S1SiJEXdcFPYO4GTAvoUoGD+xa
pKa1jLM+ra+2BwUUhnYLRlRBTfBZ6VwVhBkbUNbAqvluPUOQ3UGnh1xJNGnR5LIMiBLz55cjkeVf
03kStz6pPIcYd8Ft1z6HMf2V6YoFo/YyuVXZ+juXzP9O+8e3zA+3XdlS4mSFX9MejJeSSjlhYKzP
j5231kSXvq1g4Z8GuSuqsuyoEsuvNYaOJU9I3rsBCRqVXMABX8xC4TZ126Ixe0iWUaJ94mVlTv+S
E+jS4YIRDCdFJq7qr7OpnRweih8twE7EqX/Q8IZEPaebhX1JRGxQc47sKmWk2KaWvgVa1LxMZn2Y
JEW7j8bkZcJAhroCwtMuMTbkM+iBgEpOPEngT//f0QC/oybsnzTZEZQO6rcIjmF81U0cYvQf1COe
tyqO+dvIMiNwkGFbjqGNRqKiGMqRbPhtYT3ROWqOrMvo2N0kPHddeYoYDvt9Ck/xlJWp/700QZMK
FyvxQNU7LI1txLJ0y+/+3uSTDIBbocwg8El4/DUog5WoeadVKJmI5VtrtDdbJXp0UOTxjGOBh2f0
EYXXF/2DHuugE1nvR5CC0cDxiD0aPCCiBZHZ3sa3PuTHhrDZSoEpVpiQViArzKdviZpJySHxULUw
2QYqcDsrev0H0LodrM2LvCB11VVFdPB+zLtVK8P7FIyAKeS7aU2mIyBbAvMbRd23fnYlho5M9345
Gtr9SBlIFHU4XTbDMX9/BYJLpxW7qcpAN9gZgsuQQG1DrzIH/1r2kDT7ANsd98j16ySuaG+UV4uQ
afwmZ2mF43d/HOK88C0SaBruhZMiw+CjbZzoNS5jN3nSujPCfcFhnJSx1EwGW/a/EMMqCawB9S8i
UmwnHiRVG6Po8AXrYYD4uAo1hGS9Kyc+K6Du3ng9EcGDKrSqC3pMfLKWYLcv2V5L0WyfLGNxNje4
1ZasXpCLeSHiFJpP/QhPl1plrutMkApz5tCM35eKr99sOATh1b/F7O5aefDkrVm8tm3x9xvD+iWt
IEB14KtcKADdZVr8suobnODD1xoyc6p+/mUTdUPCkPOJ1PZNPo392gvhSUnGRFM9EZ5CCKzNoceB
Q4ruIlnVP67J5nIXiJ2RAbGwsOUwocDiulvJUiMmGy+1wPQJF/sW+1yPzLP+mAnDVSDJdlTYclfS
2IsuD2BI0nHv530MEqhBl8ydy26VsGoPty8d8EmOJ9dPDpe7RmcAv9JmpBfc2SGaJvVi8ImyHOWv
RQrEri4U2PXxFgnwVRkEZmzFD3R3+wasJ+THZGjI+R36Thtx0F4jLOE/NFAWdRnnh2+Q6an90g5T
Wl453N83NwY7pL8APY6tpkgu9i64dokIC/bhKdzSSnX1GyWaZ24pv8xmRvWx1SGn081MW6vVNP6f
q2VoIyMa9VZkcSlATnE1VsnbH1AfQOmtCWQz7QxaMDUT+pITSEZ0ct2RjoEDaftkE+P5efqbvcFv
4qD20j1C0gU8aGiRXUl4by1vTug8CMTu/wI4YTicTGnyoup9D6l2DYRZk0MVsHginhprkBi6HfMU
6kjVHMlB5XPzEdu9DmvBH4m2ww5QrqJMoANibzsL9tsAHvxIBmMSebilwae0IZrJmV9bqUWnMnPt
yZgbNDOOI2gFZJLFMTe8Vfemw/UizElAm+WYXSziJZknombd5sIItraT7E0k8YlNZGHjTPhM8zC3
KX1Bsv9Bx6grk40EIoT5DcIYioc2kPsHP+TQij8M7coVb7swDM+3NrJOGnqVPobm9GYLAOByPlUF
s+GeN8FFHgyTlEXD7J9ogHJdrvCw7rxnqZIpLqZ5vnq79COqdJk3rlO+/Yg/ZTzWY1FI0sTDhB5v
i3X4Rh53dL3UtexjQl/iYx5lpsR+/ZLm8Yn8oRY3ZcHEu+YbWCDJ/pJBj6KEP0f2h+GfntsF3Qur
zQNjZVgsDswjdRNw7nKy9t1H3Au0CHGY+Nl6XVfAamDWRf08WoEgvV/1duTnGAfARGFtBZ/2tjZ6
ECYZ8HHvXiEdDygfI2wHOly72zDI7mRKU+CEe8h4JohiTaYN++99S8u+eFR8QO7aAXl4L9/4QoSN
UzOFbopEpWEaX0s6GBnFJjxMqSIxUik8+qVTdDRuHu2n10lMtV6dXPCA0VoBOyXj+y/C2yivjP3d
8wubrQCqcChVr2xhUNWMAiD53+xpm98b3KbxRJWRKitST2CEVEn9vP1p4GkFKwy+9OkVuej9RNt6
6AZ9ESQzQshIcUk9/9m/wyyOE4h1UdT2F2MZTfYU8gOLbbxfz6LVw8jNHbzgxOCXZlBNSqW4GJtN
dAu4fNBcJRug1PKdxZnwPDO56id+5KCsKj04KKBJLcbNwQ3OH3xJ1IgQx/qsnu3m+g4yRMjGCAaz
25s+4iRPTKkVbdD0Cwd9picaKnz38xOhI8TDjhBJBqvpv2psLLwvRXPvvw8kZ+wH3TWixdGqvGFi
cQdHwECgYYsKqpSfAlkadZDoVPh/LwcCRcHzSZWSP+T0DJJnwsT/VhIY8ffNKwYXmt6+TJNSF/zK
k+E/tA6qh0PWt7hRdSD4rFP/djdo+2GOWkcx3TB+nZxwZZ4k+CzZjV6xjM4NgEDZ5Y2z4GhL8fE3
Tgnctwcm1T0ixgOASySFIHb+HKjPFQuM0dyow78PZarBeqK8Ri+sAiW8dgTqdB8nJEHN2CzWtPJX
4xdAHCy/PlpxDX714zSMwRNoPSt72G/DoxBvvrqH45kZi64tecT33d8AHuEb/tCdwtCA2BQCFsrS
NBOaGhEZcLhc7h7jDkvQVUI8naoTc14AQVhbr9a7YYzk+ZTJiXp9AHU71N4Ah7hXtZEAPDRSQ2KH
RSdAc+9EHRxNQ3MSPuv28GehW8nJJJ+1f7V59FrhaZ57Lu0CAOjIdbROwuFDuMoued7C6Mz2m7oQ
NG5BiJ/O2yb3O1uDbNji9wUj/e3lV3UvJ8mDTg2BCTGDm4knX3iBT6z+Y/fVwtxTiBph8BiDa+Wn
j+dgzZ/LcC2Fu6d4MaYL0dLDgNnbaANLaoi9sX2fAUEszCCws72UwJNitml9Z7U2HvEKeqA40upH
mMQOsiH8SMELVRtPZQk8eTdHOExlsSrwoRRCI48zcJZkxdqA14kmQcBMSyArv71ep68fOEXm0D/P
s2rxeu/6r4aJBUI3kBvKZtIvBNUbKu30E52Cg+jdS0JM6HbFEKhQStxjpu24jhJi2je6B5u/p84C
2XonX4b90jJZOte/H0hU6tHx003rZ0PwJQ2RJ3QxWUZkFadeoBTfVxBI0xr53We7ZHKr9mOKSz2b
4hscBW+qKv6YCLlK6F4W2F5n1KFNqtdlRd/VEUtjZW749j1hSNn5E2Po8mNx5LtM6mhGbeyMHUul
JReJ9lAIJbBL/Ww+eiz9BOFxs84j7niSbJ1vbHMd1I/6xWdbzcyds6sIbRQ4OG5DojZuAsJL34Yt
jO96ux5TzLBFwORaAE8qSosmAkFvQHaVQ5ofY3JqfIbVRAUuyDuylELoD9S7w63642AcmR6MzEcX
gWMqz/MA719KZ6xWf2gAkcwQ6vct7w7l/bYS7uaNahXixxvjcSd0i1ZStG+ncqcoyodDgAgImYwT
2Chpj1KUOS1qf+PjDSs4FsKCSiFYuAAtNIWUt3nZm7e721TPZ9XnU/jdyLixe0694l2tcKSbDUVo
GLmzYfnytsjgdPFiU4GmkcjIU2tNNjxhxGvOr0nZvLIrTn3Us4EV1Nq/0bj8Os7bzZkVlD7MuajU
iBzeocWaRDDj0ERv0hB1WO1dI+yLtXth7fHVS+c/6mMONzQIjXPz8tWMR1YAbfLZGIZK2V8IiS/k
/DM4OzmJBe/VySR11d0QT5zOENfpsVsdcW5w3t9QnO2ty39kvc73JAQ/eLNT/Vucysgiq/X9MLr1
Rq3AovgE7RzqGkOYTCrTv0/5jPKi4KSoEV/tv/Iy36lPvQ1IBEfXOVpbS9ce5vDSkOgR5udp06eK
dGdMQrq6zJ6535j0Roby9dUOJIwjnX68prYK0U9YOCuIRRBrsyrzZENE1Eaajb2Cg2H+1iw8OHRj
xOF+3AL5hifv+FDJf0KAc7R7QIPnZdp60irzk1QHb97HzT2QOdq5E/lkEVr1JyD5un9/M94DSDR4
Q4FZApugR5w4SpTt5xmCErnzhgmh+CRu6dO/DcePl+CN5IQ9eO7SgHI8v3Gv7D0AtKLVerQLSgPf
sBRwTWosvWPpxunskVzzAD++CeBSvdm2edVG7QtflaqvzJ64oDXigEK0avSF4O7eA+Bt59wWtjJn
Wbg7HM6FBM6BlDjXgvJ6plMzx+PALNY8YOUcMsMUDYiiyqmCM2ggfnpPrEKhNS1tQnrRTCBxjEjS
5ioV6zac3omkQboHgqzDd9lDgTTANAc1cYqYuAzZmINAJp+N7AIKBTeu02gGOj4sNcIzyaqSbGaF
4b4SyCET4Sw8tl6MXOBrUr+J9xIicTVF0oeLp4mrKD6HbvvFGXxTcGzXGGjjrPPXtS4bMz/8tqpz
amPeSoGsYKHcrk3A2Y8P0YF9WT7G1p75TfUrl82CwV0t1uV55e2mN42Vb7k9l/pIYDAiwdUGWQ4u
Y+sXpDFdVASKgpLc/BZS+yiodrT/NH6kMAJ3tNXooNWyp7lda1T48x97TgovCQZwTQ/Sde2wTZ27
3PF8bO+tWv9w7BzWAc4ZgRl6+HiBzFntdOqrmxddDG/SBKpxz6eqBYjKizG+bGrHvGj4a+kEeqTL
awV4DYT4UX0pUi7xEBtIXh8TssYb8u9iS73IQf/ZsJVlKVqlm21MfK19+8ce2b+JDWmHTUT7q196
d34Gthg6GTuhtZ6H/wRGmbxYoZPLdcZomVAHlMJNUO4ejSLaYJoR6no+gDK4ux/+SEM0x6mDA3WF
aUixLl4I1w0kB3lA//VitNoUC79XsyyJZ3TpVrv4Pt1zyAFZSWsVFzyOSSsWuzYKO8RYiMSymuS0
M5pTVW8LKTA+CAVgiwfYy6kiiM+X805ij6V0VoFEk03+UN232na7/xioiRf/YaKj1jgEKxOdNrRP
7bYJKl9LhWa6PvZ6xtxCUI6OY0AnQsk45dKCmDDJHuQsIjQbLvytyzD7QLJwAsQh9KVi4HVV4BIe
NzrlOBRDZIKF7gxovqdhpBCB3N1gpDPNy/7m6dOS0mTlSaBC3hWDSl2qntaURaBURWGGuSIRH5Ui
9A4Xeq8n96DbybZhNsE4Ro3kakcvyPuXGqyiPdy64AqbRYSxjmrcAjCvIIJxee6snSYgmeoCYGQD
7yxYY7Q7qubZ7/dlh80HAD5KqP0z4ohKHhNx30I2Lvblhyr9Bzo7o1tgD8OcM0SkFRNFJuDPhuZu
P4qaLK6LPvTR+Faphm6F5VTE6zt6E1+LlvLJK7ZwFmDfk3aaSbvusu6DFYzO5Z37LC2+yQsLbfb9
Mfb3rSJe66X0hUnwl5Eu9tlCeerskJGv+cHyKfEZABKDQRilgNuDTA6A96QcdpHgJSymaBM5PobS
nBcWA/jyMAK58ftDMNYlAz8ihZ6o1FYqPE00cCQyJZ48viOjmKR1W8W1Swxi7OwxwKRLuTruVeHz
PpVt0jMYJgzJ/YAT8Rre8ydMfp3UzisWUUV7IONGgvqXgZEMyCOg4pFpoh37uhSPvp6dYjBu9E3e
T5cXa5RF58684+EqeWTMKTt0cg/ujscLU6tItvVVxeGIlFrV/xc6lStTigKpTmIPEjoj5n5GGgTX
QhflsdZHg9U+iBWsNW/DTivL3gm8DrQ2WiMMk/Khz6G2tZo8z/fREVaGMF12Fo+jAxZ/UMHE3al1
e9rW2gcx43IhMsXD38wargP7ym2DjIadQF9J5RabnPMfox++qwalDWYiv25f6oY5pS+D+MIMbj/W
eGWSrfEVIeAkb6nkOJEn5KkF0aXZdMLOpEq7OJTcTtRPdd8hKbB7Pqzrcxgr4j5t/HSWpF3ae5zn
aeLMd0lTn1CpvAHsz5Usa/wmmAj1hkigppyXQi3u6GQ+RvM+Tm2204/70vhzhG3JOnhGogk8ANr8
0GXyJXrYm/i28V4pt+/2rTVPrOyyzzfOHpS0MPH2aHGUl+jFxwC8mjI3tkqXScWt8uJ9Q4yaaSpZ
Jb+G/61UmoKws8BKtseiSwILIYrvtuGfen0PLQEXG7ob3hEDt96DJqAsfayEXpzkzb9JzxGV9A/J
bnE5/aP3zEdHzmaUAwdbkPiqVOOcPpHunorRCmSGvXfSD0AT5S73tldVEj/sKBRmShg91M2zEAQR
6VveVyBSvpCNxszEFzGa31bzo+hR96tJNHOa5A1Mt/6mhSA1lePZMaukW/RljqaYf2QolfEK5FcU
SmEFh72j0Z+X7BVrV68QMmY2xFGtu0aRZqrNJS+45E6kJnZ3/Rq673qrw4OCzPekgqtT8apB5m8L
WamV9i0fnxKFbKYia4CFVtyIMTC879+xlHU/arJr1pwV5JmJuhVUaPsjus8yO/0FFnLsiz1V6I0n
OWkkHYZ9mTnCEOTafMhPZKWrVzaGUyRLqVk8MClNiHxcVqH4+4ox23zGIE9gWWMSBAE990jK34s0
7JGqJMQpYPPp0VgiBvAeHaJxoUOUZJn4b3G19LHkWRNlTEVsBVzb1j0qoYNGVyKHi0pfgkNgjKny
Mqyj+JNycKjOwvwAzRX1PYPQzFsUH3cwtTyTTuPrdJCUhYwFftg/y5i4tSOVRBVgvZ+yKVNgEywA
WY83QYiQgLCzOkC4ViW0hSOIY2Z7gOpcC9/oZ45J/8W50y/W34GS1tMC9JbOTPJmcys/IUtDpIlz
0N1nP72wZsVxhfvJGoQCDvRWski/jqhkbn6vnhkcyFRHk/pjirkJMJDeFt+8t4yp5VaLCx7fEmD1
PicausNmOuWc1nfymyh88mJev15+V9zftlNdYw7AkbNHC8lMREYro3U/dzzgscM925+piXYcmwW1
5TfiS2+YJyM0QFNI7RvGUpb/difJHor+mWn/oyAK2Q53soRZ/1MuT0vNpohBxR1IqY4JHx4kaR30
K95aMmC2TIP4VH0sEI1pYX6jrKj62yzdWVlY/5fnJyOxUrsmG7N1kUsOdlAILMZuzjDwMaYVHiaY
6L7LFbTyTiS2/mDB1unuBppA1W+j6XbJQo2CXi7pk0SwnmtpSUJX+JdG0o9WWwafIe0o7OHekrH7
67ec1XS8PgWj3QUOODXm5KCZ/kmKrB0WAWBw1hzBtdar54wlw5R/HYpZ7R6SlKHaECu3VWfT3kB0
0Ebx1CXQW5GNAXmS7qDuuHh9+foUFWyD9OqFdxo11evnSREs0qLK308d1bU2GBSWCkPbksrIZ22b
HHdx7w3rDl3dI2M27hMgAgxXZue0wm3Z7IVCgCdWXuByo3gYUgc8+5mqDWXbxRIoia8w0oFHsuLG
l1+GfGmi7wgdQKvKBGnKV3UBh+5OR/jImdI+JmWarr/k6OsJiO7s72UB6M9PhycgOez2i5B2xpSR
hNInw/YMUw0/evutouDyxKMt5JcnW31iUAJvSeDd5nl91dtNoH6neK/GHuolkfHyyL9f4tu1uDCH
8B+M/eYFNydFJ2xptRo5e0ODoSZ5FBwo5g08JsH+Sn7N/PYmXX8YM1oKgFgkUiOivehEVREOHwpN
OQ2ka48z3aTDM4ZQmzPFWOKH/mcfhH0ZevWF5xz+saJ/mZ/B8axWlKoxtWUN8qAFpnuOzZqknWgs
uQbtMTVqdGX2n485mHxLCi9zELRLV9DSYhtiZl94fB9VFWCKt6Kdli/HUgu1r7SuJU9kjOY/kBve
ZWzOTJmkCMvD9ETmPd74c4QRIq4Vm/TQpDbYHhn9mtS7GgTvAuluBXoLCnfCoGEpit/NbrNEitEL
78JI6DQjEKH6REWLyAW/twUmu5+EQHgbeztzd5iKMIHoR9N/v4FHyCfQ5h8FLbpMHsMOdNriZtX/
lX5AwyhTeSMqapfKax1AzdfSAYaDPA7oQr21lw84I0+gnAh4nSd9/J9bJ+an80OvIHF6Rb0SdG6Q
PiNhXkulu1tpUWFaOINI73znORqkgwGjhPf/WoAqPgjFDD42b8Iad63GWScWKGkNbq2isC2f16o7
h9mwzNcsL9CV/O23AJL/D2RCQMbFbwqHSPn3OwtVP4yfamSPvfMJ0Gd/HD/FxZ+hIiUNyrIReJx9
jJA1hb3bPCd3EmemGw2wsodVY0hPhqkPdeHBiccCYuBHnlwCVARgI9ZtbUndomqZF7q0YfEqntd/
uMV+dfcGPQoLlyoAkNlebQaFf7RUf/aXf5IOY3YTMG2xLh5Z1SZx+VJbmjEsPFHIlvub9F08FGWf
EcdsBi01X7RADbcT/YdE257hI/QKicpXKgFXxPvdzPg2+7G4aitGCIHc8g7IGXPUaByCkEKyzYuU
n5UgWz77BNnsVsA4eWvInnR98PSRnExsnvngq2cmWn/NJ2yLlXFIAkZvmmmOUiSwd3I6kJws8vUY
A+JpxakvQGci2empMYU50rJUSPSImfstAGRhYRAldsOE/IgNgx2GLWH8+9NCe7U0eIvcxCaB+UIY
ekUqpbdG9BhmtD12D2YAQFztLQKXzwXexOmg1iFER99gTtO88khGZMGEgKlN/luCoSFUmYE0hXy2
pJ0zN5HKFIC60WFnN4rxD7/yomBEvyTUcowxj9NkMs91SRgc+HW84WHWdZg4YOASvvglq3u1ecbc
FyMtxdsoVnmQz2umPB8YiQLC5ScqRb5b6q8vn7fGA1IVtKF6RTeDOnKQMMp+0wGw8p89Nj2qlfVA
wcYvZ/JzR2Wvu7HQ0z6AzFJ5lF8huHZoWo8jDAHoc13ArI+2h/aaNS6Cx67K1Z42Nxu/BVJ7NRC3
EOmP76VjfFjoFrXFrXXtHHRXVBkbNa8JYtlRenRMFgPP7AVJkyg+98FP2mIBAlKUUHn4nI0zw2EF
c+heLlH0HMI4tlcLU/iwS5bVD/rvJKi6mbSVtVeo+gLcYmW2d6rjQbm5WfBI9UoAnmjD0LTJ4UAX
N63TOMBD/0wyf7fWVngLPz643P1YvjHAOSk+R0rwGNCwv1N2196qjsHbADLY44ZP0uT+u/MAAxXD
26+LeXru57HrB/kTerw8D/LWrv0mcFfjkUUEhDDWq1SYo6jjJgHrDa9+j5tnWa9TeqBGh9ILEb7q
vny9ZZPeAgSM4bAyAyoR6EDc6QI3HIxkE5iPGkcEMFMy4KiV+ij8Gxeh2e5FIIjrdFrB16OfhjTJ
bhX3NN1/vdxwO/e0UWoDiFcmRoP9wlMg9Q76iOaM8g7px6KtB2enuRnUx+inmQMDySkDoQOzyaXp
Y2w2OPBj0airtjcr+00SHxc89BuZV4jK/YwmgOkpCPCddL2MLjgJOEYKDa4zXaG1pLXcDbuJtK9d
nV97CKk1GwO/CkLf9SD8EeG6fKg0geIkoH+1nIYpl9CBkNJoojsKZJ+uV8dylRri2Mx5Jq9CShH4
rakch9SeBqBeRNl3ooPcFDMBkjJVlQLHD8uUcTOiASifo2Y1qJ2cF57/JJa1gqSqzi7cGjUqli2A
BVAh2paOhGh2cNh7qGK/Hp884payT+voyeB1xrg2d3w0BdHX6B9gfO7Zdz0/2KEKdmBnXoLYQQqH
SUzCMD4QRuLrIOSfY28/abHZPq4DZ6wBQ+OzEZpxuCDQB2NhHjzevxMz0I5DNEB+DXRMpBOQ9mLH
o/cdQ4vZq5dMnoGTup4l3dg7RypX8TzN7+Q6AHi13Fp22f/rdgm9RJyb+AvXnrp2XYe3LXjbTj0I
wcp72DEMUQIrx14f562zIzWpQ88bOj1MGBgt3u/zbQJoXMQUsb00BdC8D15Fzj44BWxqE2Mq96h0
J6nMjp3zw33T6y7A3+2jsTQmyFo5YdEfVaoPMCne+tUtzFrs8/DLI0L1T/lnnUg9TJxd35Ei+e8a
xpn2VEDoUdlonsK6k1ntxh05aY6fSnQ3cOmMjgwuyXCzDdM7/kiEw/zZf+3RmdCkkCnTl1zY60Wh
TXK+rCvONrIK5wCgHLEKAZXAHz0KEmxaCcbIcZziljjeWq2SBO2pfTs1ymYdWHCf5TtlGMeqSblr
+SLZq8S83z7C9PfsKQaFH3JJ+w6q8oXMT3wGVt4JrWQxF8p1GK3lm1gpDTL5ISzHKHbCDsIMe58A
Z/zOVRadZ4GbbTr9efaCP6nHnf5uNOuMoO51kG4/PfpjR9UO92Vf7eqtLXH6yONroz7YAqBl//mq
vaFmhx9Moal/eouSwf3t22YlcSbL4A5SrDaZwyO1felpn+7nWa4OUBTgINnQ0qm2LFqsInU2pIPk
VVPVw9uH7JupqGFi3W+4HTJ9XOVzEvsXLjc3qHrKRK3jvuYlr/3tkVZsenZXXR7OSX4A+SUZGMTc
suJeEBcJVdv50fQ6+3unN4uzyDzk9FMaMSPkSJUtK/yhGTMnYehw8MyzVkHKw8QaSMASRAk8aW9z
bWKItRUDa3iuVNQ4du6q0JLXgl7ZOIfdwKw4WOY1y4BAIqvZxnazbAbE0MY6g295ZClU8LhNl0YU
rKGlvGU1e5ybBjMKGHGdZKMouyfHD/l9e4ifp2O2J5p2fOSuOfTIEo7gMSSP5oDNpeDMhqgUm0hz
1C6f6E4G/Gq2i0vGGmMdc0ztogXxWPBRzm1nA8hpD3Kd+VYQbrAQpkvVu7Wc/BOTo64HmxwFBady
XC5nQTvYZcInb0jR5cdB3yF+jLWWBhm/sDvabsAqaixXgqYXzpqM4SHUIwEE+bYIuOrPha/jeDvj
p95McPi70CjoTmUpxJe8NGghS07t9kt1C9Ly8Akt9gscBWsF6+YSJ+5RHp2RHeuymN7IlyDDNYxL
rOXyN8IQj43aiIUGsdqYgcW0PGH7FF9Pgixd3Ebn4BenrVdk7cpNzVjSruWVqz+I2UOf9I8vlxSm
mGRjXMzYQS6TQgBglcPR3FBc//bjS8ZWQwPKcEko7yby5PKx80F3jYH4aMcMD8ug0bijqbKAxxp7
/3nS9orE7AoSfmj72kP8EqdcgsajRRbrMVnpbz3Y2Z8qPKkHEL6oLnYKqsmuVUT1ZYXxzQGBQcwo
+lDCGwQFTsZAy/9hymi0TFRIh4ihHC/zWUIAKc84zJgzRdlUxCYTrXTT59INbl6699GIeP7Tu0YJ
V+CEY897PNCwQx6WPD+BKGFZzZC8AMyIZf31XPD0vC1dqReljJsBfD+b8PLbqAZx7gohSSgqjJgm
KBYLHR4zMGsTUnkdoM7TWoBbETsX0VYHEiPrwGq71JzN8r/dUtNjNlVaxHTpRveWgM4nloR54wCv
c7rGa/QEFjInIVh7k1KjB/4+OlBURjDVSyZDUfpzJRKC1nXceDdK8HgzVh20g+XyyOL3lxTleaZ/
LB5EY6WVK5CdoYUQovsHxrjhctsA/kaF87j9c+I7IaeG4d/QelDpzKo5P+VcSUK0dznTk3RRikyd
U3t8yiy3SkrStZ81kTvpjZm/JjjWHAInb9IOcP5KW4GTB5nehllylufO/XeAnTg+3eD3kSCKEjge
vNWTRRwlaCL8tUU5xIdMDTf50s5hdNJwpcq4mnPCS2g7PMNB8iiJZrgWXZFqfnAbgFUqRYogPTvg
lhlJiWUeSQKtbIhF6H1G3K3oRU+XAYHGHQ4VvdjzLvwZqS/p8N49f5REJV8zUREYJvwPmU5M0vBr
5jk0DIK1n6rHNirsxuW91eX+SLTADK+d5+lChyzz1gGABFI0QZiQY5wibOcJ41nEpYXSRT8pPjoS
4O6Rv+pLJm6u+RyNbIPDhagZv1A7wqSnkG4udAzMqvI80tfrveOhHiNyNilCtsLtCq/D3EjU/ALL
0k/71JmC55XX/gKDEA+VHeeMOTqrVZNzSQqbe/AecBtcbsIJoytRZWKU8COGyRDT42unAIdV0W/T
/rLu5A5LlzlhWdC5QPTJNkz3b117VLGY3ip1YNELa8oFhpP8QOO7OoGQzThIv2zm+8yGTYAkT0HE
C0YJhogSnoq4lHLDy5b3DQjaSLEvhBTlHnlwNS1X2qOODUcxebuZWnvlzpwI8wsomN+w12OgJo7Z
PlOKoJYofX3o4sp9o1VVIaplHOOaHAD5LH9N3fjv1USjkaPVRq4ul+oxxED9sDymqFzmjaNXsDYT
LJ58Hy8fxzLayfSixlGcfMIBti/0Qb2wdtQ2sUTNMDsmnz7gbzsTn9oNpJvtql7GHS0VB8fgyPV/
jsfLFcBdr16Bo2LYezB3ogIK1weZ7HsCGf4QU4jbiQs5u+gUAdzAFNfcCbPKJDag7LY6rUnVUjyv
tmYSKJIhizAXAHhoPyydhtl4BrgKePCGzF5LwwO5FbRhWGqQjyE5kS/DAneWkKxEqu19xE2RRzAt
yh7mqab+FLrL2m018bvzXnRLUk/NYckGtKm4hMWV+FGZ7uoRIeqV7DiaXN05U+do/my3DNKG9hCG
EoRg5Gb0gk0SR6x5XBETSRioiphkGwqAAViafLu0cSQijs4ZHwcdZkUCnrnEQbtsYovRflRAHRjn
IdXOcqFVjQOY5ojRWQzTHJNh3IBwdtUHVsSJ+Xb4V6RUEPJ6csjsP/e0In+3IzDLCHKsSuJDmaJe
JE2ntAU7hfteUCCzFisPoSMkOXNGys7dnmtWxTaPEjNutKjv2YnAfaTWaL2vRn8Kpy2QxSzz6SjA
zwqK7AoaQsDlDh2eHGwOE5VHvVLiv6P862Gxp9y0riCSxqNPOm439Av9U+boucAN51cY0x4O1ZBo
l+oOz5ELxICnI55WW2iy9+zQ87LHT54211jYCo2f6fzyB1+tOVrq12TGos7QgDacC8SRxx1cM4w9
z4g4K5Krqb40Bhdm6wW/mJA1lJzzXuURZZaddZOL4kS8xHt5xJ+7W1SlG9oEiBana+WKS1OetEPY
r1Ob1yeDST9qsibTxEff//ECClhZRyijmUi2txL4ufAvz16hkoKSUAVDSc3WtwR5o4y8R+0Y1tkG
uTJvfRCHGTcMmdtQ2MoBqsv5Nes3dfrDOW+3gNhSzGZCzAiua5VvMoZJ//w26SAtG68kgC4Mts+J
TMUeEojxaZ3xwzbTZf/trhqK1kQndUYN9A985BClcMYsOZledAOIR9M9f3aeF2ZbNftT6YmsCSZX
B+9PX3prKNdaqTR6+hhkchcmuOIdEcX1TF2+OI+x4kROlTT36/9ccvFqoR9HDv4R4GZmzeC6EZt+
DNUoT/mQ784hRgHGGzpt9YCk2bL8b4XbioPmn16tuOq3yKzMPeJ4X7XdmfJeCJ+7lXxUnA10t6/O
MNsYaq3Nc0X0q56fGkVYZV+24BjXi6k5bsgLEVIYba+keijs1sh57JyLvC1jwaujd9TBcHWJkWX/
IbKG1UavIwX8Mx2aPn+aij9AVKfbRtheemR3XfY4sW1nnHmYUsliMah43BzYLsIr03nD9e9nWADv
T+bU2TuRQlOEJlQy0lip4ZBZl84fPDtNBWdLiPubODJTsSD48zoGSxAwZ9X6f8+u7MsJXKtq7nZP
dGWRjtkiRnkCw8St95+C5hcLvsCxoG1pKUz/y3gruopYG6MaNXHmdV5Ub8ucenMPkLwpxgqwdBlN
Zjo9vsSgxnI/0Dh01HSQdZCwiXqMT3EeeWrKUDohOq3xdNY4mMK8iC+0vA+uV/q3saS/pwv3RD/9
JU8/7MoFenlglhO/rnnZ2q0ZavS2ZXTwqjdVhzFgkKm8XH0p9gKnJuP8T6+nfekfy54xZKo1Gtz9
NHzrWl8eKePeqx/BkeeXh9XMHywRqq4ifNiWV1CyiPkccc0+/LK2eSjfdEboRbLtEQYwR6Jcucln
RG/zv4e5hlWjw/1QlV7o8OTBa3NLFa7RsPukUQ9937fFsA5xRCD//CZgBIbu6WWzRqocDVaOzdze
/h8ObrPOOACR69eLdsdxGbHzaxC4iRnICi6DeTQLDluHQnt1ZryYjcVxWMVcX9RAyDpjyRi6Mc0Y
uanXgQyBqc1vPt+K04hs+tzFAXLeITPA3a9pyyqltVAfjsSnuZq7zbFePQ70/tS8eL+XfNrKWYUH
9p9kSNPXcLAJ3UOOIQqSkiqVsrgxz6xzxSI9oD657qCZ2260FSnrJu/9qH+pRL/pIlrUBzFIMZil
FOHv2o08ie9G72wU+OUQ9NykMcP9WX7rPiQu431IOIQJhRxGwWX8QRKm1MK8SzogAyKy3iQfe6a+
6risIB1P3+kYFH/lAtwgR0dIME9ZO4S/TWzjPANaG8s5ZitOEWfBXiUUVcodTH0UuMdGnsyKEyV0
qgZ0AOkQiPnxEL4SZ78DOuIKRZ3xwsB679LTzU3H2R0QMQx1Iwm4yembhFqMA3POeAZGfOcK7IMu
B8Jsc8egs8lWGMlqSG1CeGmul0iTAbnsc34d8GzbJK1t9rT4hToIPRg/z+IQnlxWUJwQ+tgc/Rjd
akxPxfZ3YIR6T8ktjVC6nIcOVssStpiqFeUfXaD6VDrDP/D8dFHjBgkL5vuYH1BTyU6/2JgTydIf
a+dvqgWJH+JYCKHzU/QxANHnIXeQfdpIF9iOUSpR0+BgwX5jTKlSkifg02TP+UBFY/v+UX1rAAYZ
r+Ih2wr/LX8q42z+5lbSODZYObSDCgRgbC4biu3LHF33klAHgEw3c2M6DOdac7JceoRttTntYUv5
KdyMjy4WzD/G5zKOrm6jOe2dBKeWy6uo6bZrebbsI5mG4IE5JeNuKguFkc9OVGyAMyLDAc9gsqLU
LgBfVtmQCTync/2HzK/zU/PpzlkxeUyoqRB9zjXdEcQ4TY/PSBQQwE50SZhgLEaX0KHDalJdgJY5
MT2fGXiSrFlt0q/Nxvab0BqeR37Nhf8YtdZJYpdACdFDhcec87wg0toO4NgLojiAtjCqhBIqqLG6
UpTMlhrqkFQ026wGSiVN8ba0JQ33TrKHsKOWFfmYbV6s5yHveEs36S7I7q3tHQMzCc7N3/TCLwlJ
spicUdgUg/R1d6/oIrJ0R4GaQ5FfamRBt4NrdiGvy2HmuDKBG+81dvL902OSirbZ64VQrNU4qMGE
DNX6002CnowMMPTN9fepIxPnwS750x/llHAJdB+8cFJ4XIz95xgSq97wWUHcjtsDsbmuFJLZ2Cio
Sz7mmCkMUTEiGzjfB/qSlhRJM+8hawFhCVpe6gc9coY11UyE2WW2ZM8rJ5iYBpJo5lgYx+0rSswB
Ni5aNgDaeNNvkpTtMTAvflQORDCVdpFtjTNvQ0q2wa5QfQ4XLFuuKYQzfeD7wm49HthMPKPewOZj
oosoTc4CL4bBWbRvlv6Flk5MJYVb5oiTktG70PQmGO8rpzOAm7fuGwPtr7yDD3z+ISXx8rY7OayX
tgbc0ayOMf1bOi8Bdcr28juB54Bzv9nxiSrBQjo4IQI2nFR9g6hEvHKcT5S0iC0sr+eGh3MPQiTN
9lSrqqlNayKxKj15y1rzXQMUAl9bno6UbKwXbXK6FSSZ8MlBTbP9O1Pzc4kG9ft5km5rpIOjfatc
2HN80bKys4awH2Pjbt+EBJYuoKygg7fiwxVH56tIre6wR9PQrq3IKdGPR3mabK11PYg4Ttvt33To
1rAbEAPIn2sRx9HAKlNT4RXOX9F6T25rzCKzFrasF+t6b8mwGFQ7ZSpYC7/bY9KYjKljmH29dbeh
ata/c5wbbYcunhPF2hIj8FJzstJVwEU0RwWE7m8aIFlLTgfKm4c+/7YStJEudZWJn3sUQ5bsq7un
XwcdkS1bsTXSk6QaKoipIhDItfjc3ysxdLbDGdBCMgxkBnkWuYpew5AZ4Yszmf+Gk5tGmpjC+5Ol
7wvAGT4K0G9ROx/mlOv5k41YGKPEcCFPBoLWWC503KVx/GTtC0c13Vq33UVDbyaS7dZZay8UbfWK
5HlstN5DptcTVvVFqxlcEKCrviiexebx5MX66iR5MRIqDRvseeUKmJHKRPp57W3Fzzpgw7EvHzSd
QJ1DhXuY+1Vcp4mwkwVUbeaXeMe9H2V/qPUt+k9Qdk3cSgpW2WkmQql4X+EQXG0xoycUDGkHMXXH
EKzTKKTelBxk2IIdmKsI+KXIu47Z/oiWEi33xlK/bLHcuxxVkj7bmv6y87f/YWADFmbut53J5GGb
fUFd58roe0xvKuDDrM3ehVUiZ2O+35JG/3yZwHa3LWbFk0cPHJzd2YQTrv/RIC7Oa20vzSbarXav
OlAaQC4xC6bUTpZ98ZsjYNRl519uoR//j8ygf2FoIGg9HA3/yQNAk88sw56nBehHT0OmYwqZDF2Y
ktIC7VypDpg34ZqoPKUawWsuq3sxpDhHxhQWhhz0jxLmtsxuVHj/0bGaXP1hIQFSBM8Q0iWeDb4U
OsTY77XtUnI/L3rKt/UC4LBj9b18URuxNrFWzuHIZ69O9mgu7qOWbaM/ijy99NuWl094xjwBVLHO
5YsfaTzc83cOOhmmRwRF8VJrKTaXAUt5/RY0nnyibPIe+q38IaenuuGbVESbIrD5AqMtt9sFga3v
4L4aIKqIJeRnMRNdWprT4WtpNDZT8bddUcCF3aogppnLYVnQLBmeKIWTkPPhi5SLbcDlGNyClw1N
0UiEABqKplsRyvXe/a4ypgtHGcIY2bdnWUj4bEKiHv9T1SP11eDGgSiGFArTTCvrnbmQGk+IZ1E3
jrLMOTYKvhBIgWW8zTtUrVDReFa9AfL4zY5rz0rsbwjFoM21QyupsxnIP7cUOELGFcrvnb3LXtaK
7vprzDPWnxIERhMhvKaVkNcv/Tp3Ng75F7qSIBgsEAXhpUFeVnvgRLFBgP9SioV7+G8MqadtqR2d
Dpm2o7yuD/yqmIt9DsB9zvlnVZBTWZnLTYAhfx91ueICvZnzo8Qt6mBnvrSx77oMx5tpGVu/c1H+
oEQxQ0NIPxI81Owz8q9WePzmrsrQ67sHUkulLoAiLS6RBM6vpu2NzYZ74xfGjFLQtGCaHtrNAt6k
RFZXYmk76gazh25qNNk98jq+GTei9RzLimq14dhusy1/ZBuzZvm1nOBaZiPYIMr0cDhkhoc29JeQ
Q8J5ugU27TviHfa6MDqLM0zPwcJcKHp4gRsUVsQA7jHvl1d+Q2DQVHWvYOyTzdz6JajHJcOysCyC
HJHn3FKHj5MPa18NQdnvdIqgZnpRsczcsW1z7LZ35l6Gvv9PDXHYFpaKTt/8StmRhjuL5g0sU/wQ
xMyCCG6Xyio6wkYoPzeGy4X9hWPPEDKWb9QI90ZG6xiDphQ4PFX808gcuelil0eM/KLgUjfSygzb
6CMc7oBfFh+H+DRr1lQXm1GSztvk3+P5a6FvuTkgEPEofVUu6qIDB29+YZ0tmQNGcIdoXU+pgdNP
Qc5qP7qc8yQNqE8QM1sQCG52/UppNvE5uIoN71MXb2Iy+4vTW11nj2kuWhlMlEJ7LTHCq7wovzlM
Prb5oeUdLLceQd7EC8SroOocVdasOf3jhZ0gXtmm6HZaSPdr++FInqP0XhXnhD5w/J53c2V1Aqo3
l78DAWu4Oq+gapjqljGY5s4GtEfXrj//HMQkYqxS9rxG6BHGUf/0KNAGwgIMbZBMvOIkfjGIdM0Z
sJBAlynNxzbbjzXFp3VR/Z2vONotS1ReVPV5EHEcJjliQSmH9MU/LQDh7KsrwpQnhwLDpDuAiXqQ
dJezD9jOTANn1KeO7x6kpOS8vBEWoZA6tkUEl0vvF4JP7gSHDgmKiuAFtezS/GZ+W+B2ZDZn91q+
uogVNpQdJLbzc7f/iU5tf6GBcxq0y2B2p0EPa8ZOvOAPf4GvT2zzu3nPZJX3jo2V6Wm48hW8s7qL
fXMY1q51AhH8xea/OhXfkzITBIgNYS9V6QUMT3jklnoAPQUcNSe+77+XFDvckbjnGZ0SBjXcLC4w
AnIJuqX3RdG6BgnsoOx70sXHJHD2YPzdthztPkDrvuTuQcRybcpWVT0AjGSjjC0zdUuYKl+BNZ7j
TJ4H5rKPqx0K7IImfzqLiwFDUNtFR2GMMA5l7DxSBJlZwK2jx7RvE/IJgJe6Lu4/FFSOk0YwghtC
WlB0HU8VTj5thFoSLkP4zNhX0o0vFHV0oH/rp2dmbsUgB8hVKu6eQNA2RLjQAM/mKTrrm5OkoJAC
rxRRUwUmc9mghYlNfcYTe6bRHfSYVEyxWuN2kDqYwkIVOGMXwgPAcKqdf8B97Xiq5AcpBE+ZdefR
IGjEQnQH/eDE8dFByYKZEIfGOc8LqT5PmVc72Qqvk+6pOUr18dttUuAnSOPihTzIYGmy1/S0QkXU
CL60RXYJl8Si9A2cl9oR90YQLtb7lSnZt/0NMXiv8dnVnUd6Oadeskf7HNUqVetWrzny8Amay0ry
RX6E7cn4rt5R6I/QweJy1Vkhip7wq33vLOh753Vex0s+S22aWy1KNgYPAvwENe9hMzS+gzzx0D2n
Hrr2A4rLQmABfJbQMsXaA0UDSklDuquGA4sMZ2Np1y0SlxshqD2AJB4of1DbrBUdFpb9kirmI6hQ
Dg/JeOG4tgGzX244j1tuTq5+ULsH04r1WxeCDgY7H7UDHyWVZJn5l1A2ujblCDEhcXg98thFsq6+
tOlur1GWTGdXz+l9Cj7Q3jfGYMQN8oX4hUEpJHcsmjLhucNHIlgH4qpvYDcyP5/H8VK0R2tm1xcr
PILkMaAIpDIwaBWIpi+L3/B5nU6g/gKCilNncT3GErO8Kwsx9L+A6+g1Sv6EPzEEe3D32dPQEvzu
OFR80luMiJrwqdmaIKtzfc9Mj6W6jzUrMkAbKLFr3ZtoZjxbJC3FRVxgnf7eClj+CG1OXwlzyMYr
rQ1GRl8DDtZPmZ/HCA4Y7ZUMna8eyVlK5x/eJPprLK15ycHIBuNUksmppit8Xb1aNWHomGVLP0HJ
ZyFupRU82AUpR5XfqgjzgpUcZXGWGmOvhh3swWPVxh20PCE264ZpYS276pHR7cvu1PrWLjcq3qIC
QFE3cWsRPM/UBQhQ2sNfni5goesu0KauZ7WQ3MRyCoNqqS0iwKvR733YNf5pR4Dv2uQhyzDwDkMq
cE44BHibOATsfCini2o3wqWGeDtwld4B0E2pdjeDl/r+wlj3FcnK9RTRXSwuzbNOYOcXswpdKcnb
ducWnasCmX+nE0FGpvHinCaB8vPZnlCmOhr/d0Pxt9Ug5MBcKcdj1/ww110HW98zvyAcIzNUENJE
bwjmQb1Kx5bpVqRAzlc/lo3l4rkxOijIqfqNZ3hxeH2d3CCAFtv7T7L20ezkOKgTY7XGvX/zWiCn
PGFNpP2NGjycm5mRooZfkREuzJWzT/1BxdvbvUIGdoTYtgL7FAFvP4ktboi15aRDbPn8LNlHL5Db
Aaxrb0Xe+QnOhiPb09tKPBnW6JcmixGu0cBsuzI6fOOZDga69thkMsz/89waJfBAjORa4PydQOb7
aliQjp3JJUxGfc21GkpP97fE8ZQ1WXWUQS8VJkc9X9sTLwmefeDNAMQLh25Xi176bZ7Jm6H/LUAJ
WqZtvxgG+Xg1AUDw/6CJ6Jc/yzhweWj29DZ9PtGIUstzOE/3bWqHVnqXGB/Qls889CcGh3HSc/Ab
DGcFbjZNoLXge0cjrgqgSGkD3s0QmQCaI5VhzG19CAidpEOgp/jDcNi8WLJiTtmE0zjNvV/KEpdq
2BnBCwDj6n7JKEhKeotP4Lk/8xhDsSf0xyEmyyebVIQOTcYloSmi9aysf66n+thhxYbByRT9tdNN
7PG+gX3UhMefPYtzsRlJtWk0qj3d9IOQzxGd6zIaMRse+SljDelozSyz1motnH44ztKS8p+R0zGj
jvm3g/+lsQbfKhqkqCmq4QXGSNds+OnULQIV9Z4K1X0o0uNfywmC8ScjnIUqAiwSkZ1xnOuZDjid
U//k0zssnpU2qN1phQaYTdeVPym4TfRLoioEDUSAM4HcPTICNd7fnYWEmwnHQaK661E6Wpj9yUhD
0TLyQFnQUHt7Ah9IriskDIjb9gdqGiWRiGqwokBejRqefVxHMqqS9t9Av5n9UEdb8sxpgFEoAHmC
phtLD7d1skYBPRrR4iuqlMvDa/KNZz72aBFK/yxk1HxXqd7XFNMIcMJB2x/dhPRvE0lPBv+qLeL6
PgfXoLaxUyuuk/3KqFNdqh6l1beHx7/INv2Sx8SEUTF9R7GJV09nqICHYkohffpNU1dZEm7BflZ3
BA+YBe90PTXi5Vz1m058IQx/jPcfBdRAgvKbroxoLilcjQXyvkDcOF0KXSTK6U3QC3GabBdhoZwj
Vu2x40FlGPp/TADXdZuS9k0oC+KGT3RgXlAvA7ybp2Q1LxhVjXegs1whcVnanuaFYJtjsB7pKnea
g0P3FH3Mf3jYibBxv/SSDmVA9LXrN1hsGCPUjFnr7jxe1bdJ5vOZDLDaxZZDnyx82d+bpaeIDEo/
GTJD96J6eU8Iu8AkLbI7DeOoAIS2wefSyufzNtPpSd1MsbDxV56v9V2Vrq8JvktkWFlaGR81fXim
Fy87OiGtXdkJ7GhrTlXYX8HN+ftHgfPHgCobPa18bMg2L9xByhoxXRp1TqEbFhkTtyShJqx6K9B2
tXSl5+w9z99mV0AtwAU2MIzzaztEw1xcizrON8z1GEqMqbeilxxuSHbPVeVkg1+60SOR99Jfj+D8
PTVzudTm1aovreMq2Zv5P4dBMEArsQlX1/x+aPPHSf/QgeIzxlG31KnyIW2ABhEuNJ4JSOSvVNvQ
hrmukgfyOcxhUwR0WOqi1qasP1j2jPri7YKon3MxFuPeDlNbd1qjRSCgc3SsqHxY6otvgPulnckx
G+27hRpDZT7rEo+Ni9xXTx0+K19dTTqieyWD6O0XcmIFkhlByZjsNMBNl6/krDzpuRHLYDsQi44J
zB0urrLVlJ4b9X06DKc2irV8CzyFwGjgJP1x8SrQi3CCZYldSyr2REgaeE5MCw4fEN//NwtN7UQR
m4wgoGWTYyB0vBbwoqYDziGE0y/lY9wkwwmfHeaRHLOq4lXzAGBoLUb/qBmMmUJLt3/8FEGYwr9/
PeT7MYCH4sXw3V8Zj5e8wJy1uERy1yH8FCFNe6hxC5wR0LprlLz5PQerp28dKcDq2DwXQQ9GjpHt
s6L7JnZzBW54zv2k0jDlxwGJChFFtRSnyRtNwZ4hmLGxsE9x3nAFxEZhlQ36b5KEm811ADiL62iX
uDa2yRm8D7ev7BlFwIpwHuS6iJX/gj7Dn1eTFUAtwBgvB87vAuLTrC++ChQx2+maqNqQnOr15gt5
TN+mdKWpyoroAaf19dH89I8DIbipm6l9+B3Gux/8IdOk5m0rvBi4sdRTkrPI5T0mbdufknEI2w0o
jtNeDU6qJEJkKfnwT5FC5zK650+8oSqdkMDyPaJdqsnm16g8pgTFr6A2yOykrhnjQzvm2BJavoLe
6tC8Tq0f9ex5E6FjqQLZLAfKNnPnaqL+p7qH3OX+g8cq/mTqx+jRoP5o6Xxn6YD9z68OFoCa0QYs
ggWNEe17QtL4XrPc/wSbQQNYw8DQ8HhjC9ynV/KnwX4tGD2iEw49sCvLj090ORvpZMT585CdISUe
lmIh0Q5AVm71AhWjRr3u8Vebsq3aNqjicW0RXqRrzqttE5M1vhASD6nHGNmeuoOEMawpwQpwOzTn
YexyW1P3OCnGTEMSEe3/9aDD0ngve2NG1Y43wjG9l+NgFuLwypP3y7RPh6MYiY2pkRDSKAg6Wa7O
AArVe9jnI9A3kPXDE3xlNa5aZl9bwpxdsy/A+ej7Hm2A9j/FlWkaFtcLtiWyI4Vvfvt1C3y7ukNF
Lj+6AdfJ6J+7RIx/1dcaiagiumN5e9IXNT7z5C56HU45rF3cjX+A7LKIXzwccL2KqjXPhOcS6ilD
880KEKRpUIE5KaAMRl3UzFvjegKHyA6dICEmNu31IxfdpvalFgBcvleY99oYUuX7jUCO2rx0odW1
eK3eRGpc6RmosyEOjxjIFdZTMo5qR3oZPq7K/IxnyeKFsl4bl6x9fd0OKf3Td1YwIcDcPK5t2seB
ZvrW+argK9ViYcW1GPla03tv4cv6YZAtfYElt5ptiNz+OhmZHEYLbL34wtHQ3UuAUjvL3cz0hTuc
6D2xp1WXVygPL3RSrYHCM4/Xe9DYp8wofzgVZB4GaVtycrUzpN+MTfVBGGdxYBBaYCC1TnO2caNu
OhsJYh81zFHZG6vWr36UoxDGaA1GVPgJPvn+KKiGYzpbz0GDAGi8octWZh6gVldh8BfJUorYD26w
xzphga/qsYmX4fFKWyEEOxXYRuKyDA5BVwk8Pn71vRMVS4QKBhumEK17QcLa/4EKW2cVvGnAaUww
6QiSaBrzQOh6eEci6diWzp/7RrtI/m/sewofLoBgdQ6og0D9fAQe8L6SeOoj58qtcqHmJ9HTv4oW
dqFJsS2TOIgXWgEPT8ax7RQBtsDke6WbwRdRdiEQAgtoC8ZF+PV7HsjXVJvQK7RoXJkTHj1gVNTB
Zt/yDxwatQ2+uRJOTx6+pLLW9cBimjbozCG1Yt8gZaZBCIJxgzUhnORxuNaThso7+vYuVV+3GvKd
iXJDE5oWq8H/6tYxy7D8PpgOjPNN4VhPeb6DMeDhKhZlJle/ydRppl8MyhovQS6fblnC9vZtwMpn
Z5ZkI5eFOtTQ5Rtr92o6jI/4std+cj65Osxedddy3AJtKvuwvfANRwFBJ9wuWPWaGhHSvzgwzUSt
pThCZSkgbpreJ6dUjfOjLDMxKMszAix6+sEz2OaGnopGVhPb+PBYG1QTlxwDw7xP5nKJ1eNHjqXs
/CuJVm9J2WunZIUxiG6c0Fr/j1JXOAhbTXap05eTVmJe8cXM5hXtx0DGfi4u8KkuLlSR0kKl3MGz
OOVupxnKK45TE65daaNmIq4DniIvKSGW1gO+NhBig5FhS/Gt4C2HkFs0UtzN8NIUS4+48odnBIfY
UcZRXeYlvZQY+M0BShKofoAhlI2TipUhP/F683cK9reg888pQgYDQS0+IK+yrLCYRzix7cEabBb+
caM736TRlzC54308mkLRNOGEyoxSOufu2kYPCoic7vfvuhAYsX5+pPX7HYXMmsKDOhIsv+95kC8y
XfQtwW6BgFNidzEkzscI2bUTznoim3u4bTpCiA3vNlvPzpAkMOh9p/tSti3I6ATj0myaoXeSDw7l
Xxb5Bs0WcUtDGpEY6ZCN/sWHSA399OaFR2KQs1Kd+4mOrc5D0Lz4haCO81MN3NSJNkEWl59IzUfu
2Lyk3spjo0h5uCDm2JVPMAjDC3LbtI7OIbPnGZEgAuOkdPUGSk+S9wIOgdRtU/y+XqsBweVPsmy9
3APwQk3OwZ702DxEyce0b3tRYFLsKgwrdLYtB50O4hjXZk8xipXprEXun1Af7lhB7O3YFw+lyOar
7y+wmtvBWykY56D33g3+n9kNxn4Fyjnt4PQuAiHOv/P2904eA1QSSAVXW3TZI+O5QtiD7S5M488t
njsa6MgBu2IdNuJnRwazwVDpuA2zDkPeAIebAD0WLpEQs1MetKEXmHcyZJDckOHDJblVJ5MJw8cQ
R5T+zoxMaOcrF5jHuvOy1t8gRRR8avixZZPsHAia5bYoxCKqpnrCQf1AgS+x/5uB8LO9MeJ2CMpC
mGCRPHQmPy6Pr/xwPFzdBs3DjRGl1GCrY9zvmJ1B6xcK57g0Mc6hEOAWgNnu90C9UQEu9aYEbWhG
9ubPYXjRznKhapPGYMSiwhYXoIQIdilwHCKSJtXdbGsjhiqARZdBzog7DVI+1GyE0m9YQA2xNgqn
jk5Ath0gYLlMvApqGVvWhXaN1eAQI+q2Eg3xoUedtdmFNBSsqC0VijYyqTMT6xx1Ite2Ofeto1Bh
TY9O4GqpahkYocoBrlSRqOAlRGJJah1w+Y1B2Ntt2W/0PfOemohJ6qjTyz9GW9klKMuY5Gp3Jot8
zHBWda2pQjHDVyrhC767ZTan4/Hfj7yTIaDPBs5UJVvkuR7RaYdiqaZ4x5ozMJjMITxe0T8FuN5k
FMPo5nC0r4/qeaPj8gK/f9Ib/PLBAOPcEFRRwOAtc5dLIKb3megOAFDAS77BtOooWRSIBjogCkgg
1ViBwGmqbvDCbVRqLwjXKFCfD/8cFRw5dQ/buV5dIlIMM1UnsyYr98c9qc9iwrb3SOWYQo2no4Eb
W2zlanb5jLf+GCwksSwwWoIlV1Ymv8W36vfN+z/JHxKt6BRXBc/D1unPkwv/xPMq/qL+AWeSne8S
IJr4aAYH330tk9fywlHHXvbe4rk69H3kXDtIeVFVHchQmmxZG0SbMANMZG0N+1vk0PmpVcJQmpwJ
M9uOFGmSLlPGPpmftQpKuAl+lC4VqmiMs/UCLKoqo87gBFmgdsdVcKnWBl4o0D19BDJN57Lkup5c
zb9cQbQldHJDzCOwhtIyOXrKpC4EmFcWwBCfGfvkh/tMwdn6Rf6Dti24zwB037p1gpRuOhtKyNbm
PdEvanJPD2Rh9wgKagFJX7Nd01yTfbWtmOKokqWrAztq6Tg5TlDwz6D05h9mjcyWPdUqqkCUxE+h
/Q/qweA4xUD8JqigvptKiSRysNa943+KQUfMg6PIQJ1PIMOMjjbkgfQ5DNhLan61QL5zz1JjE3+N
t75op42goChbxyD4Ynzt5lFSq2MoIlQVuDagDbnduMsi65/3zRqnaePP/FSDRxjKSgfXIbQRYl0m
FGdlU5U9mNdDu74fR4u/TlwxxOsF4kRVc4fngI5wTGcn9n0KNzdOVaaNkO6VoFEERhBDJigdIWrQ
AdyKVWd9bAEYye9CQY1E3e/Gm/lr0sTP02K+jxWkYoHSwOU/vJ9C9gPTeMU4X57CCaoM/xB3b1o6
7pLjew9MQzJdNAZmYC49mpsOQFTDZGPd4rw7Q+ldPz03B19/yscU2wBBBkZ39moJDUOcYEu9mtuF
+yjTSX0Eumt5yeg7TDpzKPiWTnoYa9aSO9iDlHGmPcrCyqDqsfbFr/eBEzKigULJK+FfQtgpJHoq
oRiH64GgZ8SV2vkZmS8/vznxDJban/pe4iHNdkl19JcNHOkOLfI8c1G/aW1/ipOgY5U19vwZPWUY
3Z47eOX1I0K9oZGqMMQmG+aL4GpbZ2hegujdomlaKwhj7GACnHnSgCiap2Ov0lA5c0psHv62o9n9
uEYPgJb267o+wv+GtE1vtxkubUgcA7L9pXRPbQxG2u3QkkWh8PAUsei1Ay++Fzeu2PIV8YPGLfQz
OKZuDWx6+N+h7g1ar36ha8EIRhkBDDAlfwI/i4numd27coNBalO3eGIvEPbKm4Cup/xeyyK2FMTN
LYNg8odixEB5Gn5MiJKgjPwt9eE1kQmhPoyVQ0nRv7kJMOusYrijQ/+tC7pjBlcYaBWv04CSZ7KO
Tin9GGr+16PWtqhvG/TPgUMku5wnTyT8hCLHXTSJFa9ZEXLEg5glPa+OKCb9MshqXRd0Cy7nsgat
H2GEFlVpoPREMh6egzRblq+xRElpj1OIcQTLNjVSA8Ae/IPvIaw2EunWCA9IYk5iLXqVbZRXMpPB
ZeQi2lQbLeHn0+aIT53EkWEl6eGHmC+Tm9M0EcEuzJM7xvVcxLKY5F5xo1gO2pdlEUPvcw3Fb/qI
5R5ieuCeTDhUbaHwYXvZAmKmmEG9FnJHVABHD25ffn8CUscdDR7cfv0K2vPiKxs7n/7mAMJVxHyU
YfOIW5HolyoHpAjbLgEOiIziwyN4bqAZ8eOjAumUgrckUH0xdNb/W/TSGOvELxq4XrPGqK+1vTYJ
qD+50zh+HnwL92VCvwPkTEGdsXAbJNxVAVkzOvWPhhAHxa8v75bQhOcHpqbnmsW4vN4T3l7n09eM
+Q251wbdqgvpmk23al5iHLL48c5eq/5qsydLzp3LmUfGoZsaBn9zA+yxHc59bzXlGc4mdwK4TuC4
OfjOHxSkBlWY/xHGMWwPn76kbk8xMk5RYPJOilnZ83UaUuVuG+mc1gUyXiRuTP5D0c9fEFDRT28m
ypfj7DPHKeKTQ3416R21UTZFKCq1u4zliqHnC0W8Wn9lj2cqqQbRAJWHepMkridrsLF/Y/U3WXtI
jA+4HfyhVuxA6jRZqmjVYnSvjZUGD4f3qz1lgMYYIFJuO9NdZ6iRzwuqxcrWRkclLrbXG1Adkky8
tajNdN/P8JqeVxu9i4AYwydaIC3Ai+CHbehTlU6NiBnMbT9XJFqDCRCLC9SAbvFLfQt75wyNp7xN
ZO5Jl5NOUDKFkARqdiIyw4USQ/ICBsW8tzlQjoNhyJEidPM+297nKDav8HzHpZQ5Hx2ei6DRpd+X
DgW3qlzUvBC110dEvDES04ZWhxMZWtHKBmatLm1wpg/D+i8RI57MyX5uiyTRhKEZI5qk5Va/Ba9g
xQ6TBMSdNfN17pOleUVRGrZU2b5qZOF+xGvePxKJlyD7EpJRjJaq83aAmtDtOwvVk5FlUu+ZdQ9W
hvZp8Y6d+RLgYKekxc4SfcvaO1XBOCULNBtoEPo7l936NsMwYTRck++uapj02wYtEzt+n+F3JDNr
iVSsddok3LrqwqyuNW3RfX+FNb+EP8sehLdQTkjfHaoURXwNEjxfxi2q0vpBS/NR4vioVEmtNPdv
26AP79q2zBIMA1oLOiKHa8fyYVQqXTrdfcqQy9ZiyZJtr0pOCj20E3L/m7rFpHDeJPHQe75lfZ0Z
ROml5uvwjyPOB4Rodgr3JoT41KdP2hX22vXGtktEWUiQLSagwdo6fKUNqrk2NZNGhzlL6tGqMmIr
ljB45XCxPVmitsB1vlJ9mdreMicQXfUDfALVxokY4fNMRyCnzbrv6OsGKa6WTsvGuNXj51lvUTMf
JUamC5EXU6oaBw1ETpVabGxMaq0vgNsFrZiNeKZMxX0eAafxG1USzYEs8gQnMzbDaS5LTkA228H9
yMpHQ5XvtFApKKxw3vqEEDr6V1xtzyM6K6o4B6kNH4Mvpe/6OtdBPafBji9Q1q74LnCqveCPPFCM
BqATjZdEZqelz0vkP209dcyNFkBTOU0DbCqUwZz8TZeNl1/I+frMdMmOpJgV8XLZi1RZedLhcz91
H/f19Z7w5L9Z+HomLFvqZsjZIHKzhjQy3X3jEZdYMOq+8cbly77l4fQ+F+m3/PTlYvjMjr2JYzQ5
Wb9XPpG2PDfRsY51KPo5hbcsN73Tpci0Dg38T5L3E4EuyITEfCWZRscCGsLDYC4zw/jkmL9dJ/Uh
tS3E32vi0SBB1wJpLxz62lm7rminNGtY5qbx8D7YI0mdLoLHsHZD2bv4yh9ipSFSrQJqaWcnpoED
pFErOotKhvTNv9TpVpgxxYRUUZYM7zFxw3AInQiyoaUX5GOqQ8p804g2M1vc0NKY/PVKTNFlTLvs
nSBXU4u7uWxO5WP7SLQ259PJTEZY71WPMu9ZjdmvbWQYWn03jWp1tiBSCtcfuuQZtyBz9a8B6Rdf
QBv3k7xu0zZUTS0Nxt8R1bEPShaVmWc2uzF6EaCrpod/yrnJyCcvY/io2/N8EykbsXCGFryBGAvT
lwhYOEGRGlYjrnHf5A73QRaQKICuXn7zLNTvY1CiEGipNiyM1OhLJzId4n4vA9ui5ykgiH0yaWhu
nZ2/HH5BQD1heOOgMujNlpP8igGDdK8bMbljROECvluM/koUXm7I5nUomeRQtNd7V5vzcoyHtDoR
6+CXOoV/rxTCDNSztxTx1QvlB61vRPKdRMYfXOX3SaDvjAh8Gwhs07uuJr4mQwqUhul++iADJwJG
YBwWaViPKMk3DLaYAaaYopL5oFoNYaFBPIDaPzFWTORPq3X1w8NNHcHjr48S8mRS11jYrYQb1aVc
O/beL6jkZS1nJBlhrCZsvaq9G/i/fH9/1LgJ/UpPS+gMOrUOgs00Q/us1GWs6qAaKT8nnAuGziVs
VJ3RSAdZf2N2/z1ccWAhK3BUazQGtrcMR/fA+ciPO0D8UM6zyysdNCoPZK1p8yPJ31wOMUKpZz7A
Ixc8b1NuRiW7bwwKlTPAcbeIMxWW890XAXU1vwzF4QD1HuecOrQRVVGvgHup6xQW7PsxCtQ8bD9o
kiKnEP8BKvdQh4xSKNehOPcOEAX8OIsu97wGVtR4WeZn5twMQ4odl2Zk6cqS0/M3icKx/VAixG1i
3MOC/BQis5uqSQeOWSVgKcMipO4Wlrgu5CVXPcRiegxUjcopdL+y9Wb7RJV6F+ClSSSwbbDS7LAy
R2sobAbKo9CWoK0UUIVmD57o1fQiALYk3SYw7cbAfhCA+HE+4OeGOEe9R7wIniXii1M/XhnDg8MQ
SUK/0/roiOjXutDjiteheVtRl/6ghJ+TbKuOzNeVNIB3Mp7YCpbsvm+HCEPxAm5DlSvskK5nyTGZ
UXXb6mlthVK6eeDXih4TR8jPUNxpG/D2FCSj1IOpeacNDIj4vQoPzf6iaVcdZcRofZ76b5rejLf3
hl1oIE4/UQD+L2sBWKDSG3cCMO02mlVSXMo8O81l0Tueekodig5kfd7vjt4WX8facLC6RSulB2NK
4H9htfs75F6REhfQ3osm3aSOR3K6pvqVgGvSGUKAvh6/vpWgjzwIrT3pygcbmhDoWtan/AZu8ahP
TehWzWzgLuV/2s/KaQssACi4E/mOVdR8i3z/JBrrgFvLICud5GYWD6kXKw3mMn30PIFq5nUGBb6G
eo3zE21ppsCaCdtxJ5m42uy1Y2JXTu7QzY9I4rcdTDuwNotv7ZeEHNehytwX+fTGgEKkbfYLjG52
g/bxqt+Hkosp3MHOsdkzSWECnrS7hzAczvyMBnBwufwAHpQgP/LQDcEzonEF9HheTge1TTql/+0N
jrTQ7FLLlc0RZ6YWN2Ks12GP5Tp6LPAtpjn0BN891tVKloFfhqCwCCSCzEoTC8nBaT7l9jApv/YE
xwT5Mcn9wYwJbuqEIg1rl5kbmx2LMlLuQt6tcAQ6egkkdXWQQHK/KHc6eNzzJ3QgScefCrHrmixh
IbnYwTgdcyg/79cn/cAJaNNXTe8J4xXHAoSpbhj4RKTCzwkf4Ivg03o5jK91vpZWNzltf6wBKOy8
akosNrUh5SXeBLAriFYlbj9emPoueVimrZ2CIKyErAzF6E23jTeX1nFio9qRJ4JNtFjKaekHBGFj
PkWxoQRp54CIg41dcaApIPUWkBnmt1IVIlPizK030JeISsU0qyBmNzCmvMUSgv9npV3ddENsKPHf
JP7FzapXE/gwAL8CLkSPku7Am+lL3yyMoP8oOfJDYREhPGl5j4V2NDdZV78lLOts66D2dMoUMU2y
uzFFD4w+1sSfXA9zL6IXECEO52T+Gm8yUCmUUv+J/RWTDY3W4vRU4uOLsRZ3CJJVRPE+Ei7jf5v9
BwBiQJq1oGHUqo+LVjSbk/VkGyisdlKmEoAXOUkiSDW8iezIJLYzqwN9TRGe/Uh1PrmRIQrxy6BC
ejN4EN3dQEQfZB7ILWoEWWO6KjJfN0Gt9s/idXsLe7/EteUaSBF7Szd3rwyQRQu1tWqiFk4Tj2qw
Xd6K4vQES2nmv/TYe6vNBeTlJymCmcmjOMHG1LfPbxwUEpER2MMVsIsqapFOa71IHnlkwkDCR/3G
DgWAcvbqzMhD2YfarZosxsVL9RPhfFQy4x0dJXHBklX1CyXUY7w28QNEQMSpXCX1dhSjKWl2yNcQ
lPCZA/Y6ucT+3T40Qj9sk0+G9Fl92D2ZLZ+9aVMRu5nNGeDH9tBDoBmBLEKSpRoLNDOJ71QkvBO+
I0ICIwRa0hX9xWJCrElXIh+Se7KI6YF6+8W3M7VgwyGyJM+Yj9kpMrsuAxXMSow0rG9fNzB+JJZ7
tvUX6R4s03dTBCJXIVEOXCvEZE3eW9rE5InSp/cyVceMI3lmBA8bR0k6d0aaJlDgh+8oUryM2Zvm
0/yaUz0eqSKeVooqrOB/TsHDLWxbLJnckQWzlBg5pjaZ2vYRoiMaoRmSxa9zPDSe0QzcTUW1pwvP
SOLfwnfCjKZarx9HaZ/7hBrfsvUArKX3uW1fFEjYacHq0h65yEs9Y+3qqyEeqvEDzJf5qZ1SqgL4
8wBivdBvCMHWQuFV1/u0YMeVjKOgdiXvdFHFZgHG5MrvmjV7gw49kh83veC+cjFOmXEKjjhaWK94
81+X7kqcyay5XSYH8xXgqlYeWBi6jYFwlyfSK3GKOCQm2o3+cnKyRP4rfw/yeC7m2jqXDGjT2N9G
4ArHnPrIUmmNTtp1HQs34LGLjiGwtKO5Tnq21JubWZpT2Z/HH9ALOocx9hKJ6m6wZqrQ8w7jXF6E
z9Q92dgrIPiJBbeyjFR0ni41jo0VlBs2G86ydtqfHT0UUhXbpKvPFvYg+r+m/hVa+Qib81qjCgze
2+lH6h5I95OHoccKjkFxrNLbMGsxt4odIW37RbR/JLjxWygJ5Wpnue2uIj3MUS046kLB3Bd2PRaB
1yrMdE8xwKH2MzAxRW3nU7+XabR1E/rBzB7stnKfdwKX9xy1G6Ek7BqgqWnnD4jJH35ZZyzsvlHU
/hi0KDUnmdA5kY2bvLHyqZ3eCXDfLlHIsimVZhBMY5UWgA0iohRGIk3luXoi+0BHz6BtnRPsmiD9
AUJ/0HlBMioIruim97JsBi9G/Ab5tk8NJbNdN1XYUnmBDvRFpMaX6xzOUIo7+glJfvVXjH7IZ8z1
WtLXH2ZM5CormbuWObL/IaEcmEwd6ktuCRO8jO8qOY6U9pKnyMq39ZzshVZBf/Sb/wdg2EQev2bi
ARHjdxecv0NLKwBsW6hnEKmXZoZ/XkGBADUIJIewYVOvRJf1aigyAt+Pcnj5LUitrM5R2qohmo+c
TiCv6jOlHy/T4fyXE1tFntB20L0v1O43GslQ8Oz4HLBCNKNBHEugS7Tu2W6bcwGwjkMKjz2Ij39I
jV4HfbgOqfd8+uYfIxjdM6KVfI1ZY1vWmKqJAhlTMPMGRw6MkQUfJIg87ds7HEy/9DcoRax/g5VR
lDTjoelwZuDJz0TCEXQi8hSoSwsaNutyQvZa1L3DPAVaOkw9RL7XetGyy9sCuTV1BHTh48BCvjcD
wTZPEEd1HXyqxFZhdhsWiPG30hOFdVlvIvrrj/Vq9U3INjnK+QMwhq8tqoOjn9jg2ISCh6KxjXkD
M/HOCB3ojY5zru8xl9RTtsR6ihDaSQ3VVFT/RFJTQYcAwhOCinxrdJt1OoFNsdvq1vbAsgLO8lw5
lGpzgkkmsk1WAUqjRYTndCI/dLcx2z3vGVebFsLbZvMMNp4o0ouCleah3XRozDHj6RzFCqdVIUtK
hVxtypsAj7JiHtTAfNvmrzHcqmgApXOmQIVPXZNiM3P5fgw6yYSplGglHAsYQUeLXjWy7sCCoq0Y
nl4hpHozid+sjEJuhA28UgJl7unFmDACJH7k7Gv0UiGwNmqRzJs0udN3YpoIs26YcGrQoSP7Zuw5
PInbkP2rv18W7OHYfSxbW6vQgbBL/fOkupjf8zNZQVjenNvVR4o5ii5hES0K79uiDc1rPGpdwN58
Rus5iKRT4C+KFSMKDiD1xR8AI1fbjZmcEVsa0eHGJaU6mh1DmJzRN/bks84krHqBMNGeJ8Q0BAxj
PRq0Xc6xKNtiqWHRoy39D/03OGRTLtcQjn2Fh33zECQGPkGlkfrjW6DbmnwEak/M/ZGui88SiY4r
pie5gUZBl6xMUEL5zTDA43G+ZQKi4ef4gmImLsvIEI8vTA/1j4ojW6F76VvfOGv/Kd6Fhacm4hk7
31LzEwE4CBo0XckOIhRzGtKfydnR40z6b7fyEzHdM5UIVu8v2ZSJ1ff3Ysy87Zj0fztPnTvBwpmA
GfBisyw9GAvIqPjbXH28kEhlGp+hAs1q9Zogen3loPpd1SZya6BRnxLoiZv7Yd1vLZVKpZCXUKyg
NT3vCS/dL/blHQDXCEt7SS1BEJ+CYxDGe/PnQ3DjcjGl1lY2sVGe/Tq7G2WJnqhcukqsiZE607XD
j9jKnHTF5q1j/eOlK6zt/fZIC3sQIeppOcaP23CbXMOWodGWxmxACHcIANSjsXZIrLYVr9u7K5Lt
q8lOcuOldydK57k9//zIDvYZeNYiY99KNI0D4w96/hbvMr9TaV3h6Pq9kOT81xKvCHBa8o+SQa9A
DyynmGIqPbApBD4O3yJVxzx199uluGXJJ36A4VTUy2FRw7jQEsSsz7GRUUM5WeTrejXtgCjynEB1
6JJnfOOhLidN4pKAtWD2zJJafzrvU+OuYj6TSFFkbDr2kWX2eQN8+Lhoj+1eQI1/6Fc9XZVYFsJu
2+HOZpd2pfAxPsDYL/Dx2I30yEekowvUhL8ENd2ed3ZY+qVTa+hhMUqoDPuHz4bC9ljQGybrN6ez
2Dm5IouTtKB9lfbhXLtGAejl1+k+HUd2eEyuhdJSPKFvcDB+Og4lzbMIeX0TwKIHpY6qs0xGl/FY
5gd1UG89Ypq273Ka/oVt5JjwGOYzr39q7702IJ9whf98fTKMK2xQmtqHJeZMfFIuYTdVYgt7IKyC
5sfgTCUy2bbCgFlF4rxv7HWOmym+Rw+0ZqjdO53R+Cgmu0TI2zf06rQyZpMSenurRbCw5ui8Dl6U
HwIc3dwW0ecSacqP5Meh92qjLQsHA1N1DSQV4OkEX79ediIGCB38293kDDMnjPpPx8H5bz8chZxw
XRFusWaLRW6W3RU3hVMW1jMWJdM7yTbkHXjNC9kShWzdWRfYdA26tzIPo6zWsznVVfTfPeCCwJZZ
aPC3TwfebrE3Fl6nXb1VB+bGuJNWKu6p/l/a0RIMDu8S+OC+UlP5bVh1aeWxa+2ZBO3OUhrwrUOS
GNC6lcdhMZv6/I1/zNEug28Ac3oQOEKsWCWb7hw1ITkSGvy+xRcprfpDSHtf1bg01VXnOKPbKUps
R0n3LTqd3VAgSXNj/Ay/IPhc9g2klP1kO+rbFGYZmQzitMtXDLjY8Xqyq9SwYm4atxdh1Ktj712Q
ZjlMgRbw7pRqg8/jzqYVtcSrvvUaiinWnzmVlHgp2wVA6PLxrDSIXoHCqdGrNe2OrBsbWuikooNR
T6HhQJjxjHD7ZG21bQ9uNyAcuME4gKXHDFcvhgfVdiGzsJ1fBJb62P5LqFDs1a7+/3oZASdG6fFs
iA8F3qCcPTr6tYIKFAcsAlN+093ezffAnMKG0WuVXVFVRTHoBDqoeGXCgKu9zksmjwShxbzwH+IC
WkCfQukXxaIdtBIRaYRD0om5/lyVM/2AOBtar27WVe5nNUvQent1EQVy8ymvQ1LjPeKrgN9CMG+5
AuaGkMxv7JNjmbZ5Ugw81+V70XPP6cttEMdc4hdj+1M6vTM1Eor4xK8GCx5I1uNdosbYy4nXlyhx
6q1YP0suTPoxz1IW8hP7Wf88OBGXERsbvE00g3km473k/dOalgzhvvLUV0qPhnqpBEjk8eQhzsJ9
nZ1lYAW282oe/nknhztixdXKw2Sw25Ylbq3no/CRve7UxRMvj25/ithgE1tjIZ68GehwLZ3oCYIW
g8zGvtgFezD9Yx3YWvtOpvI8kAQXnl6htH3qhvcNVJiU+DupUYks5+18OrtRKqKRT4RME3rkS71x
rg9GmW9I+X9ALPayLQDwSTGWu/Jq//oNPmCyaEoEHRkW1MYWA27FWZscFCM6uzlW0YDa2ZX4+b54
JxbljGglzy9RfdIMS1jAZB1pb0GT1XR+FUrwR6OwjVeNc7rLWL1njE5XODGnIOWFpgc1BprSaZLF
YCfa9bcjcc0Iq//1X0A/TpMurqC/iBr3poyyla/2azi1QE+n8VY2AlUrOA61OIhWvN0TyOng1YBQ
2toIscXp6FTdxvH8yCnPrRnYf0Bjr6YJPpPoyAPCcv99QmvnwKd9oXZIeBA8ohNzPFWUThLrEp7L
LcQ+pz4ocHwyml20cg6TXeQD7kqe6Ec1J01trBaMUh2708HnjiBmQbeIs4xNbuQvLB6zV61P1qC3
WPQxQNu0rzzjCA33R7mZK4CBdxgHoCoC20iJsnJOznTy9v9KCdbixGoDmvvx9NKFhRou8gp/e//V
tT0kCgTPnsHmqyHl2Vsxa0W5crLC1/Od5FcRX0OA7EBIMyox4vDyOw+D5GVqTrSgM+TzYneTyi9Y
yeEGWIkQ/P/1kJc56T9e6O/D8u+valOdCfZ0Frwuoc3ykGf1tHHY5lxg7/CtiGDfBSqOUI14HI+i
SI7fFp6v3Jxy8f03Vioa+NRv039OaGcnWfniW/UzTmFekNWsFrt12MIUraYYapjsMBGDxNvewguA
0Hw4m3bdpIbqcxlQ1/ECORiquBlf3HWkTphizgY+rpodQkEWD+E0ATd4PkNrHab4dWKmklF6W95/
ox6gXaNGiJFqdLt0coxZTuitdVTwzZIB3fbgQkp1V8uYR50csSa1I8WNE1FIYGszWZPGNaDQTXRv
GJgbBAlx2ZpZIK7UXLO+ZbO13vGJ/Wb4m7UgG7FsGFEx2XlOtc6fsFuxNa2P9V8HzrJ3WZcfeOec
aKXeIWACNsPD9+xdgmGXauneZwszGdEq6cO0FCX1bjrtp7ba6lJ66rV5gBC81y2mjtS6KG+XDzLz
4Yck0uMLR6ZjXwwlIiORRD8HS9cwBPTtj6nTKdoPr3heWi3C3Hu1hpPY2eYsGm+scPJd2kGnrjy/
zPwq9tyar47ptU9K2nY0kJsfqcq4axhTjsNLDs3OFS4Bx79MTXdH4gXOKTUUTxG4iCp0/EGwZWfL
LI52buQb5bRQmNLkB07Ey112PdIkium1cXaDi/874XYsvdx6mWQPs2ffrg699jT6zyDaal6Xo0Vc
rMUgHkh2HfiC9Nj6KHXHqF1QmjVSp/tYa6jpWW2rBiaQwS6swOQl82OwvWFm8aEMfoKLY331FqJZ
H12Vo/kceHlD3Jewy6rYwdg9yEVl7dV1z9ptbLR7GjFH+xtG/iNLwBu3DIoCaB8NCu5qejIjZsAb
n1MoaAqsvyk8boup4cWAjzvEnr0bZpm2wg0jvOvxC7xGb9k7Ay7fLkP946/bnw7tsJpql6dfSU1d
rMYJwIudSVsAc5Sxa/hmGY/RB+qGpspLMxEmtdUEheggQjdxI1W1CFuU5v39h5LLIxcjcr83AveO
+qDmAWbIagwc6ZPbDDwd7fXW5oTt9uyj0iSZuv4xkPw4BgOJjUCl4vBSTNp5NB5pPpVt/7OcVXYR
cEps2i5v1mzddoaw/izFtQr0NL9ysVDgy1kVwOhdx3oCOhfdTePJl8P6KkLu03w11+7KDjTeZn8y
OhWK3hWHsEV9bGLM4ByGG31aHf3CYpjyl5pzpF3l7+QzlbmmSj4+Ok3l9fNEFkCcynm3L3UnEQKf
wUElCDK1lfGGjt4TyUW3NfdeG0IL47AmVZUJ5lfhjZCUGmYYiRPaE+FuQ9XHRBSaou8H8OxKj7zV
Klu2Y6H7RvdOhUNAPvVzwY0YuZiTTqx+k7aBH56rIu/ByG6t5AZP1+alhlKSNqlx3Fpv7xzuEiMs
lUQqTbOX38Lc0FGonHscXtfDJ5kcsNvCmy3+3nAxDxrhtg7qWn/g99FZOC4o8mnY2Jo+DZWLnVha
nd/4mTFEo98Ehv09xLN4G3gYjfnHxp/nqL2UsPsFflrSl1OoqAMKJrT2/tsPiGdayG+clrKOB/fM
f9esCbWeKtOMBLzmmaj+D3eTnOKQZxXaUML6zuTV3mtnkfdZWrCkVks4vIsVv2HoTYv4DaUCw7nu
jQzyPziPginVnK1LjcOFiDWZP0JmvedVP3QTXWvxWrOdB7xNuC1FpmhGGREqy+kizpUDl/1sjonn
NZcREFiBCW4jjU4pTfqMrlMwWaIYZGRsevAmGcZtjPDTy1hQlvozhWrrtqydkKL+cBIikCO21oC2
yK/K0VqxbwhVZz0Twai/WMUjJ6+zpwsW3NDEoYTpIScubd8V9kjiUQoOkrcpOxPbnBQlvlu1RF5w
WvbEjHQxJf8FlogQV24saVu13KmgoPHdIfnIfebF7aznlQ2rX8ok4DwUv0kptZS8mEWJuqchMmTa
TSNV8Bt8ft5Fme7LxCaF6sMbNq0oJPRItOQU8LcaJ+b3aTZf/mYk01JoD/Gwy0A/FlycGVgGzAgo
k7mciwlkPoea3AKuHOEkx92PO4d5EiCr5r7lB3yjJ2HuysAROvGPHVmsHkn18MsXeaRLqAGgOs8u
mAKpXrgxWZjQ70Le38LKbjOd/gXYnpdrwSC9wljuAMN5YSNJPqdpMnGmzPcUizNXeFJr0vhjacxh
hw6lfGsaOws3sIjbutLJ3nrPknjguVGQq3CjL8NMoZaRnVrn/G9jQkSybYK37dyJqLscaGX4pM5x
2vXPBntQDtPQwtP5JQLf0mZmW83c29L/J6hrEsSXdWsbjz4T8SQHgzBqj1ItPFIXYCcdZYnqPLAU
cfwQa0ZKdkWavDw0w5zq7CA1Ua6lfWVXUMqhP3QhSP0/PiZdn17x/HRxGnUe0fZTq8c88x9oBSFF
GtGeyIvER2LPl2xLdQiFFnJurAYsKspCCKheF//Ovgn9KPP9+5eCoerQIhgzxKCmsyqgr0jlo89O
Ga0YiwwbO1yitzJ/PXvq/P9ROq8+GN+ZG9v1Em7tbp4mGVyGgf7adS4IPjDzUb3A/9k+flvQjaV0
sL8hnqjyKWU06lpv4YtsAPWfxfdQxmEuVaCEYQakgh63bGjh02onhlr8M+qyZO4JWrg3M1Eb1uHI
yXjZAhEJbnOmHrDXmJwjVScg3AQBDniDBPk//gYXG2+9MMw7AtRPzPYEzV+fLY7FeEEO2p6JgHGG
Fy14iys74RQcd4w1IEbqolkG1xwyyG5ZTSiZcQ+K+VEksGtUKSG9Xv4DsrJOuPz8ZVuMITc3eD+9
L93adlex5/fkg2UJVzsC8+SQ4Pj54cDOqNzIsp8RL7PzyaNeDPBOGdDRoATdLZ36AuDquCtu6xJL
UtnBkyGCeWvcm4vk5haCfiNC5o0TD1eFIn2RwQithaKgiLnaZJH6XGhjAXvSrwjx8p4FqXvuqFjw
8dA5qInGEnVL05foN9Dcn1I9mQGwwuW/7r58p91/1aLNh3KgPKWPVYRLP1iFXI4A481bN4B94BaY
4bgfgsmTb7oK8dmD9xOT+rcsr7ubdt/0jC1MIfAKP8zU9+5hx0esctscGr3+Bcm9BIBkqLyySdy3
eDggv1aMPpfrsSehvJ/7V+9LfaQ5OXYRLks0Dv/HVk9fIwEgjN9zhTHkdbuB+EAmmLVohUJZDq3X
Av4oFJHs4WN9qxsfMmEpAuD69d+ffdhD3zi6JazvVpCQev2Pp17QddTmybkF6wDp+f5nBbUV/0wn
tFs5yCIiHdAqUfkrgVKBFpSnsSReU8zqyg82ndG9ESL3a0ajRbGhToGtbFiCOeG12L0frMtErbXf
EUscynCjMLemzrGk8G0S1gJbL96VUjfKwTBBcbbX/OnOLjIE+X+AJZlwTlnYJsziGWVaHhDkzB7S
aIYkM8ERt+VdhQoLxOTQbMkpGEobhVrzlJSPdAuBvBLKfyu8iyFtlabdSAVCi4eyAcrN9IWZX46A
YgZK/0W9mB8NnQv8w0zt4k0uceJ9ztVAQajaaReZ8hf8OcX6sS6qFnjPPZNP/ez/wtZsNM2Ky7VT
m+VdB+bVwyI/Vga9Kvtm1T1eAuL+97xD+TAL6UChuO+1OM/ptbt+cmYViZjvlk+M08fP/eohPI72
qPGwRI2Qo4TduNfjLKVfKnzp23msa2vwtT2CmIpYty+h3YCQWyK4OxDfmqQgwNe0ETCKiHRFTxFD
ZLFXtlld61OQoGNc2A12cMMdQfRv0Z0hMuwtQnsbheAsMPvCd7QNdHqvob1mMzyOZhtplnxntx7a
oKz59LagztAA60a3s7snQuXcsr/HbDnG9bchIjho59o08rjghRFL0JWT98AEjCZC4UHE6UwE2npk
xaLChnC/BWcO4k2V2ya6JoCsYFlUdnS9uAXRXtxw4tZg7JQBB7o+AUeiUBRPbLh0E862VWY8ZyI6
NjpNv9chaXhh1yva+SVNNTsGbooBgAgWStZJi3MD6SjhmdHaN/rDj9YiRbE+gf4tiPKqWR3/DO4C
jIY6EdER7XRJWXIN+DuCH4y4VZ/XiGENmNbIoqKyjTX5MvYpl0/w7Rup+9XwW5jV/y1hyf5LBVU0
31NAp2saB8C6w7dYWZoYt88l6V07TuTujPS9yuBX+BmrhDkElNZCE3WN4FcuIGqhI+/vv/nLMCnR
/eyTAs+j0fxOVLhXZ6cRrKuoPgfkqBVRZOxM1tFJ9GdFJf/s/2t8o7dZSGWCdQqL2qbFRXrOnUhj
59VZyhXssish/0gq/lanpSs9VA1D9PO8tSGD8oHl7leYAf/DKyswVSJgKeINkHujIcgRbb6qkhGm
juPWVR4aKk/hQ4JIq1q8FEyJn0xL9ZmM5MUsoefZRvsxgbp8WQX884e+Hg5WC1oO3YOoQJJFhd3f
HhK6//5lDwGQQxQwiF13HCYwTikmAsuM8RLMRAAsLZh7yaIrUosdiweVUfd/Yq9wd4h2BQUNGs02
G72FeqV6hztZfuoL6ZPJjye+28WOY8twUht/DYHJgt+0jP7Cce+Mj3nuMB7TZrCqX/Uhbfkf/ABd
wXCA3nmYbMbgjJuz7zDgepM4ZaPVt3h//KEtFHXiFXW0lp7YyxTT1oxECnu3B/Kn7DuhgwW8qHAC
cnkwEazy9y+lGKMnQTJeJWxgt5lmoP2q/h/xqnB5ENRVOhgp5ed61/33wmdWIXYMfy/T9UmnqY++
nufnwNxT4TxmM3daAQizHFbIqE97AVX8yyt6etK8DwlbGePm0nSD1TXFFrjJIFD6jE+Cly9S4NeB
8uEGbDY93pl4FL6nBrh/1Rp2aX6vojFCulD6UlKnTFnZzJP2KpBZ3OcNaqFV7un7otchH6ATwcQ6
Y5t3TK/yjxAdywsICfgDb+i8JvmRUDyJfoBtBru4beuIwzaSzLq2NFGl87dDqqCNbCHPV7QFPbnE
miD6ITMFh/KfqnPZ1A9I3NfFFaG44U5bJIeT0OOw/Z9HNMzvOB2mcwGFusLvoe9jKARhmtdfzVV5
dIK/xPvCkTIwfqEPdCF7lv7FFhwi0mJ/EAc3/m71xC9LoNm8DCdqif4n7bP0pc3JhnyC1vTYAXRn
jUFJQr5wX9o1yZeRre8r/TEYI43vc6miDnUEFehwAmeRUzWYxccm+0VINJKLacRnxdbbfd+ZuQYn
9BdtkMiVYZtRiEI3Q44IMQ+L6x/7HDc0/Ss/+ta2SYAmNJej+M8Fmo3Te0dmBm2mfmAitdHnI4ZL
Yabp3b3u7S/RHIFicC1AqYge/IXAg3tZz3kBl6/lcsQ5+udmp43GL6u6vP6unkhTThz8IKPCilSe
NeRGv70xC4qvrmBNMeACCmw8dsM+txYED45uNyf+DBgpvA9SMhsJojWQxRNLV9EEZwUKr/q6mBV/
dIn4dWtkaDr8UeeWAWhtPj17B6NmxVcPeMiJ1ebXeLBEUXhbboUMdLV0HyL9zmNpcKVUWbDVk1cL
eE6HoIfxQUbO0nQ5viLRlte5FpXnRTgPn1tVZzwikHTdlVnsgzcBrVjs09131UUavLEd4Uqzyo8E
zC4zewT2nasue6xM/slvp6IHKOduP1pIIhKvXSXXbEGDB4Cta1GbukCVVPuoc5FGxYTFGnqu/Eti
+YTRw5Bh5t6Ndim8vc5fS8esDDXR/Zh8Z0vLGVVt5YSw8yddTDK1s8Oh4jX7yyEEVo9AyQGSpQ2t
GOJ3pIVDg9cIb5jC4Apl5ceowZacz7fa50ZrwSFGw8VrgIAXkI84mKuXfdGNeuSs0jJH2MYHkkTB
u6F8ONHPMKMoeBbxh8MaitC6OerQt28Chz4mQR6+/SXKOTGVPN1NavNSm9Gwu6Bp9ftLxur1oqF/
pN9nl+8Xot9stP/fBkFp+EKrg/FkVpTYqxpDQwSZ1Uk6PvSe156AA42wPmaldMEjhAVVuICGdz7d
tezg4PM66DyPjmlkPuUnAqLQx4Cns6rJyWc03o84vMQ2XD+YmoOZIG+Bfuqp//2WVbwaI8JT4uzk
REIIWz7NvAqC9AREn6E09BhBHTMPhGtpzxMzRGRuFZMt2slk2o9d2cpk2mdgokaX+CKTo39NlWAr
UVbik64pm5Kd7UNpxd4zR1tJWGaD+XByEFOOGB9fqpr5wsNtTnNBK7IM5fOF/T22jmFYu489t1dg
JzwywNDF/b/EnHBgZcroCns59AFiEkCdmqzJZVBhzkbAfuCdjJ8vk6PFOPB01Kfn4j9/bm6Gv+cX
f2gjxMa3njsJmhtmYEwPUpUtcnb7ReeXpr/9Hr6a79j38KSWfBGArxqz+ocI5go2PlSV7YBwsNu/
K8flnEi19PRRtmU19DZ0kuwf1y4L8K9MjjbhAqR/DI/W1fmHrFrkYlGBuTGOoZJVeExDEaus5mW2
bFHicz4uuLSBwgFs1wN4Sz17C2CyMkKBFFMOSrsGhLhwEnEySVh020sk7gezrgu0g1+Qm2+PPNbd
EgdZNxmTV8XtYQNzRXzXi7+734anjjygc3hqLRck541tbUwn+Q3Jcz/JT+e0J3LmeBwIre4MCJSY
JPB3fe20vfZRFItjGErne9unzR+iegJhAkk+mGBx7+npV8M50B1D9JRbn+LIMTM2EX0hRypJB5r3
CJ7NDP+hTk6s3AfiBulAufw1UTU0O4WErbl/GB3qHDxaXYqgfZWWC2zrTzaT/YLNVXTTQ8PbNUN+
DMvoT/MuE3jCNBVi3FWYk4kF6WI10wKvNs1ncdRDxriYaaH7iERPFOzgvECVR3njlBe97CWB+0Ii
rfpIUoZdECIyVZsd7BWcTe0rkqxsD6Dv5KlVUSOU+EXHAsTgtuLoZMnO/6yLOJLObwHynJ1lG4jl
J4tpNrRE/jCLBX8O6Gi++jmczLsml339JotZ/Xk1EgPLMMR5d/GMVCt+1aTNQUF8Tl2jdLkAGZ8u
cml9GOeBT5nCkoHpyoDtJryCr/RwWTwBeJzzp40IvyccVfBOxECxekoB6aollbf3N6SaO431koio
82jsG0z/y/KrmBBr9jgg+KaP2O5mqVOZXwOigATlcoyyKYSuZYOivhxvh0Tr8zp/FE34cedcQ6s1
6NxxEfCuHB5iy6qEH5xhIghOlhibnfnaCbpHwUyjyC6mY/sHobqcH67KJDG6Qw6BpJ41ccGMwEbV
ISGaG+JDNDywhMNb+R48rioO+zSX5PtAwUzXog9nQ069VsM3iZ2O+ytTKXaD3djH0905LTRdO34J
3nKmct/BbRlVNqevVYTsc9/xoe7qT3EQZDVdauLqBCYwzCDdU00ulTAon5gtbadQEIOGIgYnnfg+
9OlufVxgrfF9K2JE/VlBf2xvHBYHqqnyzHpDiq9kkjh2yqRCMko/LKGouAKgmv9XGaHs7kzD5MFO
WTzMeYClg5uBtxx0Eu3FnGB46DoYK0hMYu67kJAqcDzzYyRaSzLTPFdibfWnnzgaRwDzwv3EtiK4
E/D54vWWYqTN5RBNPtYQkKPKB6vgUAB4iLSVREGKK9WyNq4jNLJfMpX6rxJvey9Vx8cDgCp0i0qX
yvgbrVZISesUVEI8RMRHdVIoKpS8EmVcEwtDwQcZKh5J89qWO1OEQjxKomsp5OYTkxHMPi6FEOKn
gzTMb/IUCtEBXxNqUOEszQvFced9nRf1MA18U/+V8QNjaa6aTeNQTLRAOY7pTo7FygPONKXXM3X3
5ubKcOW2KzSU0aVBq40mLYT+T0S1J8AKOqEoj9AJIjlcvZf7n8q6/OVl0w8uWym5kIcr/PsX5thv
AD8RkFJcfg7SNh+6EwKz4Mij7Eame30PIQhhLMWuGJMPLeT09AdUx8rF8s+aAhQi9ICLq/UAOisz
IDTyQkpcAatbar6jb2AX6Inw/92SsJm4DkqOe1aYEvV9XWhJXsY7GR3Clg+ucsRpU816jeAVhuJU
1b+GfQ2UAMiLi4HDy8q4R5wi+qvLnn3qjBDsbFoP6GnN6Vv0PhxSe3WF2P7M9mSVU4eSNDd1MYVi
mCiv+PE+MpUWzMNB4azNH6euFj/1VPcHWtCOv5ig8vS5HZ890y0VNvLT6SLchfFB+N46cAXVkUZ8
DwtLRiMCSZDq3x2g4uDakNYLTdFrGHJXXwCa/QzlZEE7F5Bwrv0A2Snbft3Qp5RUC6lCzJmYJ8dZ
LQnnP1aKEZluBQviLcqxQ5x1vvEMgx7A08iyNSJ/QKNx05SYzqYWXxH2ZgUi/T3u3lZHdtFmwkAE
0YWzU83AU1o7c9ImAEAsjlGgeojEl5ecddTzbsu7uYD+kThLbr+k9uFVjZWulNmJ0cXA2r+2aoUp
wQodkZ6aQyWSjY4h3HQ6Hk/YwloFsj4C1fVUXpzCcBuVE2hCK250RdbxTbEhNFP2MeZWeiuYCsFT
KGHa9qYI2p0GrqUkTketV7M/4uBkQWehuzUHiNPEylb52zUiHc2BA5pizRHYGZXlV6l5PJs9M8YJ
KOQFCXbqG3sc5qpT7huMsgisi6isNFPRG1aGk+uxTxWl7GYC2HTy1jJ9l5Fy6qmpOIYcV4Yk3QN7
VogupF4hUBsJLlGpxsU44HNI7+EKQZGUKukskD8WpLZPGsbAGmvWM5IaLcjERxyM3BMJWKcGYvYs
bvDCFAsZ0pWEqvcuy7jsagWA5hEPgUvq3riaPFk2JvzqG2DHSoCzfJbphYWOkok8V6S/Q5oU1gco
EjAmeTcSIaw+CPey4cJxJ2YZnz3qMv+g7ANikdFsi/749SyZig3PJNsxCNaG76vKOJF2lwlFDUkd
ahHmdzCbJz+GKfjj1OR3+3euaRB8YtC6fJ36XLcoN6pxeTQax0HRoRZna7HoaoKs5iSofiCjZVvx
jdx4s2sOOuho8Ka//Oox6S1Bpij6mMQuiT9Fsg2odeSRpgzRKZb+ERMxe0xbJzyZUMM6sUhMHvDI
+ZiZB5xAMKvQ99t29Cd8uvE+4WfnFcfRfI8bRGlJ82t5ukywJSKpEoDSJrF1OZ1NsuptMSLRlC98
76SUVkjbdhsFCJiRdZiVpJ5L+ihq70V1660RPSA8eaJB3wkDcC85J49JWwA3xF2jkMcm8evIwzSA
qnZBJ+ZRgjxclFyOvZc2mg6l5ooSXnCmvsao3B0kYb1xDi5sy3sdWEHJOd/WlIqbNmwtE05oxi8F
LXFZqOxeGQ9iSFuqQIDuujitlG13R8FlLcI7gpTodGi6/qi0Cb8g5rcXGYmQ+6vYVO7xQlaqGkbU
J/GZhB1wUBu24J2wcKkIn5AY3meqTFYlsE/+S25pLe1dZChLXAP7qW2AXzCmypPXVlojL9Xar2Ul
zHmg1qbUnL0MxtGPrM6pTFxjpe3e9XQ7TRKVXPStj9x+1pZYXiiyPF6PI6GEstyq2kL/na5pWT8N
1bbEjHx5mVB6Dq+s4idF97Vjw0HXBieSXVo+VVhN04CMvs8qxV+U4JJuGVWYeerbDw7C29HpcqDG
py951g4XJl0ey8r6En5KJHVpXebp54moaCpx33m5mNi93TISEt/odG5RCf2OkFyXf7pWEebiHmLh
W47XUEkgyjIEgKRYrLBM9dIRB3zK2/gA1D+LGT8RxD8Qq9YcSYxKaBZE9U4FFf6NElGpu4Xqmjpd
etwOyIb+ntydUWLIrScn81Fe0uOCBFXfIACugXnKICwzyjPkssu+IOO6Ix5byScXXc0dajF2dqLJ
O6+ZSfAKbFJO20BNf4juzRdhF3sq4rwlC1WCmM8MC9OT3yQh5tJxinvoQ+Nlx7gAsoOmz8axkDnz
UW0AiUnScRG4oFhhHIjL3IZMOlryvvGVH/4Jlxaf/RDgO417wakKhOGWhbixySxVB1exNuZQEUZS
DlCo2Xj5d6RoQjaTFHTWWUkDwmd+luOFMVs6hYnvpztE0k3ibziRdXq2gMf2X4JJ9RxmM5j9kKAN
OlR/RY4R5zNrIjfQ8VbCsSoGCsFBXCUcri8Oc7cxEJS2AcldEfFiv8DxCAxvqX/l2c/VuoJ1BDRX
WTZgC60lA7lk0hfYD5DEzYT85dvtZm3k3YxLeioa0vifpA1dzCv9B7OqzXhSyDpj6XW6dgDane+i
vCcR8xiNx7nHZLABfeUBDUXvykW7Zcuuwl/n1KfQiVUn2edIpyEUB0LGyMIbaxIzsATBTw+mQapV
d7NDdJGGWKREliNR0tCguY9vHfdlN5YV7qE0/oeuv4SRleoWUZw8Y9iMVf/uLv34G5L56q8fvzEq
4pzuEDs435xHAD+jFfACDrEXlgls1851bLwci+aYERrc3rcIt/Ump5x527ShO0wo+yH5ERxICops
hP8oIk5Ar6MeQ8VOcNNjqXJ4GOlHcWNVqnFKTuxi7CeQRAkV68Sug3NxAMRQ767VI4mNItvK6rU7
rOacRDmI7wZ1eNNlQhih6WXyZ5EpcOEKTrKdsE6Z0+9H1JBYFWmugC1eBqbAZfUZoOpKE3/b4tSQ
EWW2C+RC0mZrLUxJm360q/sq7HKWqi9gv1AUkhdlVFuiUSYyUOO1bIBaH4GegikycvONTk9aWb32
3tplniv34LoYOmRzXW4RQ0aRCkaoMKqhzc7SeTshP3HE64IpPOIyeyXtyP3t9UBn5fYXldRAE1Ty
6r/hi2Uod/M9yx23aySnojtvXbZbinNoBUXgBzHGme4Ui0upAl/cYBBanBrxTjn+xSAyy4KurRaA
l/ZVuGUH9YfDAKqLWvP0VSqPf1KHLuMOuqRgVjLgrSWnk6Foe/TpebUmJ3eR8WDKjYscA4MuyjZf
5LnzTKCYsgjBhgcySyUrEoSStgYuxQQZlEzNYaN+Ege5vaIFmgZ9V7BstJ3vytOU2sOirGH0BWYN
N5omcvXH7C6DA3XuoYbBnAcXpJjFChPqGqeoMkHqd33+b9z9JOLz8YTQ47gHGkdxdQLC/WE348Dq
zmiY1h5XJkKbybnMlET0O4MmcWgHCExNs3fCRaB80GMc2i/rTYRvo4mrNN8+KnQuMdiLxxcuLVJm
GiP370hZOzjZ73ga4VqGLFgfoc/yNs29i0O3THVxeDvYDKzcHQmQ8sVHD/ELXdd1h6kw/ZooEPcD
9Y64ZTYgUeMm6r+nskXDQhBH2HfVSbo91CP/MDnLONZZSyPXt50UkXPW/+XCKE5d7fDKhGvTScF3
qgaan9xserLKu01ftgXMuXpLkTU8zjFe5m6GroZUy3obnqpM+7tUr1CjYfpAtEWUFcz7O9bWKROl
xDGsxCoy8j3qsJyPBF5zruOc80dKtj1Be50havqMDnVqzM0vNh4FiZAz7dIUGKAjNEQUTuJLcCpz
jncL5hbkjNQpZS0VOSsrod9aLsikhEqFAj3LTNh/WssyVbfbxireslmJBkaqHvDcq9n51K8F/p4b
DeKMY7vfiHpMf6TPQqCoBG962ILfYbyAdQHAHbapurpn74PZj2nDCAoCRXoavuBdf8ieCbLxGK8T
FI93g1jgzao2AwqF/0yflwzGqFj4+GVId8TsCt5vsQFffeI4OdegJehMKH93bGAMF0GUXHy50hC/
RnqXQMr4UtOdaFaK4HO5ep/F9p6rGXzbTzVxKY4kBy/o3Rzc29rgbCrxgN9a9vDp8boieLgjVVVD
PSFZhqV9Z5mqIZ/mUyBF/l8ZCrlzpnfJL/a2f00AFAhM7Mzyu3QFkr34InSadSLSrxcE8GEzV2cn
K+pfSfs9N1xjRaBAhSrQMHdFGRT5CERnB8oHbWU2YA40vqL4q8qbuQJl8H66hCE4yzTLJi4CTEjo
L2Klfo245IuOtkihKnQ6Mu+yyeG+upr++FiUir/K381yOZ+y1SC8M0E6yoQktFxopEZaI43s0dLv
d4/vwtEnaO4n2knvDml/hnF5I6IK2aeUaBnEMTLdXWKURRNSuzAalGPmg7lAq4N0xC3e47wt+rtV
l/w47seufzxVBYRNQFlGfHa3k7JiiGpq+IR9x+zaGUMRlch7MhT1+ozhhDmt668Qw/W7yp6EZqbv
cRnaOifdRuWg8PPhCBXRdzVcma/bTylVkH4HFL4i1ENhyhPJ2jhbi2tl5eIKZ3by3OOopgQ7Z9Oa
agbA7PfxlWOODsyyCLMvHNNQni/yG1xkm+hnEmQh9ocoQfyYz65Sops0uMIL1j75L1G+pG8H7QS4
UW95ECpjR4qKTJ8dLIh5V3bYLZfUQzUUlHGEIX1VSUZhtvc7AeJpRhr/f4UmSWF6u1ReU2WueGJl
Kct6bMZhAswHTVv/iPPhgX/RN2BLONiqbFt059q7Gdt+lNRoC1/N3AUHE8W2q8idFRiqwBuONhjG
/1WbNqfwAm/yrVT8mIon9deQ0QE2loYO/yDYACx+vkY/7AswUTvtobDzqIwVbF8n4jasIj5db5sf
IoHlCmgzZMbYg1DfhioVjB3p86zJqWmlmNl1y6nMnF35hMlPkwrFeQxZ/hjBf8mj2MBRHMbO+tAn
wmpEHQI+2CquXjepitS4rye3HNVa0du+wYLX1IggyXVfWYBAaocxWVy7uuVq+pU/m6IcYv5Lw22X
dT08ziVPZ5Wi2JzJjWNNeOOWoCHz0RNfnPi9B3xeExbZ0j6FGlrvaFDUTJLvDNUJHmsOxoAsbYty
Sp3LI2rkFP4TJpklDN+PNmaOTZKJ8QRRC4kgde/I4yGpUvlKIbg8A1y6Vk0tXxZ4LGBqfcEkCnIV
XOlehrNSiTPXROuXit2TwefaLCCAqwJGDm39hgw0hDL/vvNKg3lzaCOl3+fu0YcJR18dbDX1Loym
lklUiDx619QA5b04lp/cpBoQ3wbXmPKELV2BMxAICw6fuu6W29LSn1kRn3F3DajppENjdwmVY+hV
wmklqZeguocCWAsYkgqBogBtkF/lutWpQwxwAbn28I/kFSECLO1PxzlbDGV9Rb48FLKqkp7wC9ya
e54eFnvHRIhAFydtRxigp5ZV+xWjeOYmVN+a3eRSiTQQwxc0guUlkaKBgGVWccgVl30YOrK+V5w1
2j8KGmucMPMziByAyv32qjJEsOq8S57NHkGZDXQLoJw11S7SFPc5ThHQlk1cQ1XqKlxS4JtLBBZF
HA8hdepwgZ733RjkqFceG56ng/jhiB8SsPpwWLOo7jzLsBFvExpWauA6s+0xsM3WFo+jBHN/4/Zw
zsyCiNjT24rvsv0dOJzOhEf/p3awoPhyh50h/GvPzLyJzov7dHi1YYoWWwqgBEJnajk6SmUmgbqc
H0ipxq9mNUxxd7+b+QLDlI608H9O5MHRVVFyG9s6FOMbbj88250CSK/LyizZCoHkFN7B+gvd1n29
+SOadBcg5ejpmdIDA8mDGOWPgADLdgKs0Ok6bFV+i2f9p5srtAjwtr2pqUYIEE3Kdx/XNqmOCrcc
AcRwBsvHHvvLBZ27TvaodQxvDkpju7tklNxxWRTbppXbvfr6gkHHyggnBDt1Qy30tFy3j15z9Af0
TR07c2Y0ia0RphC2jHM/YPpewnoZ03gLeD2/gPANx102p9atBrbf1mRLscfzbYaSasH0zii9od9X
CjXQ8aSOyFOlMRogJl9YO50ef8C2LxZLbBcCM+Z1tBOB0/fXBIS0u2xX9Knjy7xAfmhCIbtnjXVp
WvGSQq5n6BZFRvCNvpoJW7iTMi1mTzbWnwGRSuiLHKBY7rZKI3K4VLey7BYn+z13CkWfMz/w71gD
S7RplTRAh4wlkzEqbliWj4eD+J1f8ZK6Vkkzyst1wD74scZBeMmQOpaNZZl2nHMF4wLm+fLaJ338
71QFNd+hWFQSA/K06nzAYKYA2/TfceNkqpmahSCx3E4PM3hqNV+UzkRdvm3OWtfhF3QpVbsGq7ZN
NGIzaBqfkGZzZ4zn56WPn4z6i5IElaXN9C4eEE4VZ9BPcwqE48up0k4GL3OCfILYmAd8PofMLvss
KYh2zWYf8CRXDws0h18rKfB2tzLxpcv/y3KP9USxVQdW5ay1am+wNblEI4fUced7Rg6b8tSPqcMA
S5f/KxRY3QwH2OVU+7wZ6DNDNDbFPyhVxvJubgjUGv490qirxGxKenUji5R5ltgM6M9vUCA1iCXL
/ZaIAEZYh4PkZ6JrgXVLtXT7iEOhJSW2sIq2ev5MFY0IfrJKpuUHv4qfhqJL6VgsCEkUX/AL7lEj
4PF0cFmhRV0o2zGfGLWZjtvGLOrK32gfpYd41b1ikNcLfXNBei0OthRsyQxYtvChqv1tjl9lxcup
rXqFyuRP0Yu4453h1nP88BYixeEG0iy7ZaF//H5Q/rgpFya3wJmELM9210y77lKIrp2GEIDO+Zf7
1I3j0MeEjm/hW1/fM5JgV2s93q9dHDaNmmz1MUAxvus6em6ZQE7RUk/nn/yoI+hiZ57i3ZIDnOKu
u/DMuuM48C1ycAjLQXzFQ97bTjeTUqwsc6H1YcmXVxjsIZGju5fspcXwhgWAoOfNHVNAW1aqhs6E
nMtm8T+/lZgCiSglptVjzQrCKwAYyI+4k6/2LVUVsZlGZOpX2cqD7g8TNB1KCFet8ABP2XBLDrmI
MyI6ptAcYEqaAdUzh94seeZ8p8k6tXoSvfIJv65gc8xN9sWAlTKCdwNIn1tWb81P6WcD+3j/i7oE
QhHhgu3Va7lXB/pIoZMpQSKcV1ykSKQ4z5PqGpDK6p8R2Gz1KawAh/SuUeJ0R8Bcy2vzFudP+fkp
WfJud9L01h/l+R7yKqwNoXClK3c80ei0RQVENXq0O4h/ZraM8T1p2Nd2eMuHiQFccFXVpy7UxAyN
CFi+Vryp+f7zqtvcrrQZXUJSYWLv12XLpERoJcKk0etjaiyjLkQyCWT+aoljX4oM79k3OBSjS24X
voJ/sJA1+2H/SJD4bj957LamJOR6a1DZ39BhzEmsUBaGkCNyq7yhQdlLQNifrVwfKuxdqtZQxzZy
NtjvqLCyhzkI6EyR+EsyCGgn9X95P9XY3gNm54CCvkm8oqm5CUZCG13TSxhLRz7N1wl1kFdG3i8I
+qXnx4bgnkoV0HF4BR0hZMtHW5H1NROWY0DHCyBrvHo9U5wHdtbQgiXhnRV9s2eBJUcFITwmFmTU
7xUZUrzbQpU5h9qY1zMmYH4du8FKxIdS0HvaPU6i1KQSjOtjvc6volU794i1e2H7WnJss2qq0zbU
NWpBhq8iTlRL2+8ujtkVUA0FyxNsQqqSNYvrniGRUITV83+Qwm/oF8S4Qky6Ca/FfH6oqK5N347u
nriKZ/dvUgxiEpV2R8bLUnggeNX8SPNKApogz5yC1Bp4l9GhQm8mMzlJNp/fmC5AcZubSRnktJ76
v2p4Yzn9KRx2RFIa7PLsYcSBYsvUjKjGNL4OZ80ikTG7Nb0LmULFvYe2zt91IcThBFaMsX7EFqqD
kje6SX+MZEH+jDkmBQ7TnUvuTTv0EbD8TvRD/CeNh6cGR286+dh9us9FPfb0Rz/RX+CcO7Vdv4WB
MLcY9HrWxte+zsEfKwUxebSCW5hp452QP4+yuESjG2gn9+sBEynwxtQD6yA0E22OdMCtI8OBKFHr
D2eDcCowzdZ/rTOWti/5F5dE8PVf72uyY/Tl0G9irVKMIkD4rNYEU5hksEWph3TY87mLakjui8q7
qANaOVo1LSRObYyz3ypByZcpn8esoJgTTWNKdnVm/1xl6Zr0QcSrM/ZnC/4goxifakHBM84MVHh/
DPhOoNgvHXEJsMjcFbl6UrJj5VAP5QF0kdKsbmAFk6DvMCiXDLyjQhEzn63WiYU85dOsgGb0cw4u
2XQZiq/pCV5ipgjWM+BvsEEclIpmXL1vry5FpsOZR3/wPv7UtfG/TU72DjNkB9ClB3cvwWlZHLx3
kIWd4Hc2DWdb3jmZVKiR+D+W7THAM76TJnA0ckxVdjmpayO0qKo/XOiD1PgFqk3FZfqkXyAS8aXu
2hJ5kncoyi9k6YH9gbpLsRqKDIsduec7IO2Q8Ld46gvf+/eUb9U3yxwEY+N2uT78cSyq1HB5oCIg
M1UgcPX0i3TbGH6u7iiqn4T16sksZ8N2ec3Kht8zWOLiV4d9FJ4WehC1ivAMUrhpPdCi/jfdE9k/
Wji1gzHuz7LMKodnypG8v9AUQt4W1JaxCRsce34uXwDXljRdNZKRWYgiy7fsnHEKziMn+MjoDUqX
6is7B9NsXlkTPQs3KlljIeLOUU+gwg0Thw6qWAWFeYWuC1rWwOZ5K3GtC7TjyOrp/Z6Ya5ZkJ67k
eFx59o3s+IdYWfdM7+NenSZrFSr/DDMfD0ZkUmvcSaAES5oBfQ7jFj0ePrD5f61LgmgUuHXsVQHx
ZmXYk9b1lEyvoVyr3RN3/z8a18udy023j0XTuc1iPVWlKtRNlsiJqWPaOYZVm2NklnkHHwfjN1mK
oWkSBisddbEB10GXnxrCJAmqd9LvJ1p4PPJi05CYsN0KFG8WfeMd2OH2OOS/Qdj1/9VZrgcEuIAe
qFhCV2wCOsh4Kx0XJN9tlTVnsiE3gYLXnA9LBFLYGlcsHjMn54AewcUcCc/JGVbITDXMOtjt+nJE
2MoeVsTqbiB/Pct3iq66AxXfgnvwjecM253/mesadj2CxUznyh2QBiSqxEC574ZdHx9e6n77xiOd
dEF1Up9D4+e8hIRz9YTVq0ssJv3xkBYIvYxrV0WmNjEGZKaQ2OYU3vne5+6rLkg+Gayao8A/S0JH
w/i1vqML356udIQ7llKHfellwuM5PDpZRywB+pMpGHASZhgSQC7cPc5xDb8paYpPenOoc3cR8JN3
oqYg7yupjnBA6PXCajDrNL0+remIT1ix07KKOQFtztB6kRgbIaMoYFuo+QwhClxtxmAdTW9pN5fS
ekpeVASCTuKLBqRYADAUSh51yw4B6U1UR9gG1jcSFGBB3fA/Gsv5VssEseCZanZZ8phos6kiYbso
Wv2VZjkY6N8HxePdyIQj2AJagD8FQB2U026+ruQaLcm7jWi7o7N989icfFDQjS3SUOBMeCSbpHJv
ny4lkEybzo1TzNFWAWcMD51bEohG1GY/h/xvbHL/uZBqDGvhcJofL7StxazyTmfNsRdm45gaV1/j
yHS0EldWxfr0aCsBxt9/h4bSE/YANWVyop5qNyB8mdfTc+lyrepmfnEMGBsWrPqtd5s4AEmKrBvf
9iFepV4nk4Rkp2IlThGrnqAUIDNVmj2pFjla1r9ypfI9ru/pQudyEye7FkgH40gkSloIyzy9I5Qg
vcaHARXKUbFamyc8KRD0z+FX1tliEHSipBDrN5IpfYTLl4/Qt8gwWtWiwj6uL2z9qmzfEqaSU3Wb
bVvR2LbCVVQQceSXOnr1mtY06p1GpNaWCSHdq79xqOd3oZGsfCKp25e0vFH3hnTo9Fjke9bAiODm
CVIVkptTJ7mHjMMDaVqeETWvc8wB+bPzezXdqs4cgICQU5Rx1QSLz1GgN8SX/tvwzU2ovM2Ve1r5
3RLET6xpVk8OxKUTclXET9GtKyPNXAcLRkbLB9SjamfGuHXosnu28dH0YvgXP77/3WNBkmV/xXSU
HLNz83y1U+4dluEvGylkuYFDq14ISn+wMvce9niWy6A1aFC7RJwE4rLKIvT/NmpF+6T1h01F69Mu
nz7Yg6aEb+vg5n3mXGfHJqqLT1wSIi6Ki6uFWi1YfkXKWtxJSkTA19kSnS8zCoU7W/ZY2u28290a
RkeNOC4a3kZLgI4WV5EfTtwvMBMiDsOV9qbkRz6bv7IvgHeTMzauP5RAOs+qsaoMAZ+QysOJGH/h
p1c39Q0GaI2To4vR3t6kiDZaTFj+WYXiYtgHKJlDZd7TvBUnWsgmy66JWafUfO1K+5lg1YZJJd7S
VgQXBRCRu8HYfkvl2quKeM2vVXD8vDhGpK9uH9iQpkGl16cOuXCxMEKQ85q6ySX+WEM9o3ZaIbXF
IwO67y3snHnuhousUf4qdMQxEMTOuh6BbfcWCDjDT7AKHAOgJYGynMep56Mbjgm+XQWSH4cTcdbw
3pYEuLDg0I2dvHqdLKUm8468GsbYDQuFvxiJXMHWGVPT3d74RxhQyDuwhn2ZgtJ8+N8FUZIQFiz+
TDdBSTuRa2x/EgazSrrXHBH+v8PVsWV2ji353BqEE7l1ISdS+WREBjUabxuTNwDwvRwxKqqpDSYq
e6tM9j2FW/g6lLks+3H9nomD+J3XYEqlRROU47vgw3v2GH2Xj3aIvpnYvfq/+rbNcavFOHTvZNeY
AlhjQ/vn4gQ2JfmVoEebqGrjU1D8FL6ltEXjiXbWmi2HA/zjsQ+lb2PGlrrYrTE+5ngq5EXwlWzH
fnBoFMXVXrfAd8/rdBemz8PHh2D5kmtiPybkEf03dAQPZar/ioyNOTr89HjlrU9g6upbj3XkP77R
iKhBCos1v70DyMC3YYfekwV4z7A9fjIAHImfTPkAfebIpxH2sKldFxiTRtNPxOEWqEGLqCG9Vq1D
4vzyMxWHbq7ChF4sD7VONsz6J7AbtubGwCNwJSzpr9+w0lcdZpSyQb5GaY/pXVDZOAsnv4blfsWB
KE4o6OhMz1bMKagmUzmZcK5b+toY4wHuyZoz9/v+Md8qka+nWnmRgvERwILI2FoO7vKEoIdrQHAx
NnxDe6PEhM0H36dHSQjcOOZraURQKwNn+y8DODtRncMSGrprvDN8VD0HtPgXlu7ZOs6uS6uqxwp9
fktaRzLt4OFXkZMDLqGpUQEbF2fF2Og9GZKygxW715U33wDw7RJmB2+9QGek17Zw4UmqrL2bJvcf
ENbheopDylWd767FpUweUnMW+txdr9LB5TEk433AMYC6bANdW3vOzWNitaMJBYn/sq7fCSLGiLsL
lbvyxEy5DGvzk54M5h7y/5psbg+g/uMMX3O9PA1vaaKOkxMHOWusY4IQR3Pijx47xNXrdaTVL65C
gHjgsr910B8fFqEF9zMydYTcJDSKPZn0th63RMABfvTIQH4FX8aZSUUJJcxfGDtVYVCTZXw7O1Yp
Riayu0lhDB443j2CNpEAqIhWkvl+/7PfGMc8Q5EdB2RxCfGLd3v2i/Gp304motgMXdzI+PpyuGvC
q53DG53e3qVHrWweFZd90fWivLcz+hHVsMFlSZ+5CloPNR2aZMPwwZvfMfnRS/yHaD80/vgtg71t
1Dn7/n1Db1Y3+cbgGxu7gsaeIFy+1Imu5kq2bSVhQ2XolqhKbRPJTGglhsZxnQk9/Jr2txSBveZN
aHrz9qVtRBEWghuPxqr0VRwdW0+6Odf9v+KR5I5Gei4iV6bd0kEVths+1aMR+OafDLstHBmMvvO4
0KYUP3D9ClsTequvGNl2IubAkG3TGEuPJsPFR7AEyztaPrnMrtJhkHOnXzQogFVAI829Aq6QNz3u
3Z3pakhOAH6/sM26E00kKkP9/16YnTMuV5cX42fyJBqGHZuTJ/2oY8B24VdaelE5qkxaRMWhgjxE
WAi39LMeZyyNMbCe/pS9KHdZHbtEpIJty1h3wxdGA89aP4MDbhrfkVyi3YhQiCv5jm0dMhChvhc8
eysI963P+f0DiPSyCcWF8Zdcd5uW2497V81tkESGXOmSUyWWVedDZRn2Ip11Ns1RJUqPKLyZE4Z9
D4KPR41lgWWxtgM+hHINuOrV90d1p9AMznDNmJboeyys2z8TjSnDbBUAQg5Jq8RxxiEU4qHoo23H
Zn8k91EuL9YzQMxn6ndYyhysB1dGzyzYSBVE0AUqQseTr2I9J8gAVm73CUvsOr2rkSnfoC3hAsxE
SEiC1kl78rBeNmAYYEIZZrYDnX70rTiwZHJkgq4AlHW03bPFfQviDN4SJItlBfRFJXvmsQ0vhEHA
wFhV7T+gSVqCdJVYty0XkUFkmJgvxUjCPPkXMiIgLE9NJ3ucIcjC8MZJF2AiljHrIs7z4xev2rI8
Lyp64++Kfy6YICplECOTzio/P/74yIhBW+flKkB8x6OzQYTIn/MvP9iOQAnNsF8/idp1Sevnxxlb
5cb2xaD2Yzkmdr7Ivg7qmTGF9mZ9B52CF9lp7zBsxzXkyPg7eleZRGgywsMcuK4id9UcurS07b4C
O6/KtTgdct2x3eLWHHzpG6LvjOIob7lfW4Zys6vyagQSuNf1A4MlV42L1q9Ie5eC5nTklPUwrjlW
fZ8VK0y5+HblCrz3wygmUcw6Whq/ypEUOIw8Gdseh90A8BySJaI/b39iMibGncGgcCdk9poQ6qYk
l+vUhGPXeWS8oqeHJvpKUa3sgxdM73fVy7sWciI8V8hATOXzO1Is3kLIRS08nt+yDKkiklqlYvVY
Frw1WW1lei+bmXOqmp9rkL1hu8wrU05HsR6FovAcwVQleh+FeBBoqn8imCm7cBUVUrEP7AAMIRAi
rYqEemCmcnB3H21/UKIfpgm++4yioDu/D3QG1ruNnoJdB3iMRa4GC3zJR2PvpWWxT2aig6aVO9yR
dR4fUxVTDaUDHYuRcBBQ+tfuQLG721qIgZOFRfv8T+Jce9lQVGd8yaigIT/awXc563x+9HpouZ2t
fAA8bqCldQPD1fv0osi0VcfOIFj3YjRiqpIlOnXrNvy45LylZoQ/V2hIFWAbLoF+RM1xQRFQi/MB
layAtiicNrUpCh5RpMfSNa/1a2dRTuyNSZzmUcQcPM0HBEbTuMY9ZTL8GcZQr3n1cx/fvULMI39I
pdOwBZGpH3wl//E3mdczC3ODjMaFHpuMxUVLx2wzHH1/QhURGi+j8sLXse3hWDb+jBLq6wjd0scd
G/LqGGW8D//01mqrvwBHjl2HIUjdRJNbQ2DSquAxd4tSsn25s/mdNlSl6hqwygfP1FB6TvPxvNC1
RKLpOoFuQ2uvEJJS2dw/oAFp5IDQ4pIwiUgvkUiyY0cJ6DQDeyq83zsNFY1n0BO6ZNwHl2zGJ/sh
Qw9z0Th1dy/foV3tnfSA//qiHg9JnpQ0heXzQug22KayKTz8awqTgzefDxiYbuolqaFbBhjy3nBE
YqYPOMgma7ygwL5xjptvdNnmFRG1eALP5H+B2YRNcjo/fgZiu3bfIfzMdBH+KelYUUZ6l6c4hzzr
PqJ1wgxigNLbgWUP0nW1DnZY5HKhmCLYXrLvQpXy/H/ET6n31JiV8rc6G+5/ad4R7PYhuzXwxaN4
6hZd3Y4gAlflCWj+X7/H+stmeFlW0IZtyFoJ5Pj2wUkrw2zI33NyBDr6P99NJZGa8D3UPopNeD5/
W5GAbzgVKx1uPyL5D/9rhRZwIESQ+zxbWqNadCvHIOZchs1t7i22nZKMovng0WZ5BM7uVLMFJBuY
L778oIHGO9IenKbb87c64mrDXvd+4ZW6iWq9c/Ux6BmBqazX2kNLMR6uY7BuVodB9cEcNf1IrU7v
j4mDF43mOLa7EqDYRkC2nj41liiXWS2eM1o2trBj8OwDNQwISG4Y6ksBbBER/cXNAe/XjIGyyhrJ
2OZ9YqWNQw16f5nDBNA+/bg2WE+zqTmqpFMJEsS5Z18tDMeS3a42XnsH090PI1j0SFHiY8BaHZI2
ap+mJIrDwdzE8KqUZFkm7jRsqX6q8DUah1JhSoua7WsbWuJXTX9KGYmzXr7p9XWN7syRtbuUbU3k
f5XMAH/WSgRZq8wUugc8b8Y2iuu1q87lejJaU17rXrZEmHyIxu1WnNF7eDGPyAjadp6cGcnrM1J4
6SbT4tUWF1AbY1J3/ddZocPVPHwjxPPxsS4jcMJCwOunq1byfO5KzE26KtaN3y5+CcEN+8O1i3v0
Kyhnm2UWi6MD+HSrddRRRF3DAyk9NOjxgbFSY7VPjZs7+++i6tgGm9z0dQUdTRlDtiZaqEFz8Btp
412M6U3DOXAo4+qJ6KRgVlBs600/+CUPfn1XvztiS0Z0D6GrEHZqprmursSZmOSwhh4Lv6rVXV0E
1DA+A/4pKErwAGsWVvLoa46D2RyuV7owNcgruWCf4RLElp9jbSkmJxpy/0xCVHyy2LNkSscC5gyq
1kMGjACPOvgAOkrA+mF58cbTRpztWQu+J2oDvblbQQ93htrsmEVfGGINACooevX7POgsxVG1B3KM
cAD5BQc9AH0TsGuqrXZzelsk+wFNqGWcPE1DcH8hqL2IEvvoUy9949u6P2IjyhfSB7MFiJ+GJpOn
xnFAD6zm0uTLL+LM64Nj+eTCSW5HVW83Y7rPJuvvhZKVy2LBlU+/r+QQWR4H//m/ghFxLle0Lf84
eDYbLOQoo8xl8dM7uF23qNgrhjane2xxZaNJ0EW+6yOaY5GkWse86UH944AWOuwL8sYiR8oi+4zb
VK6gcuVWsAwYc9++4vg1WOwgIZf1voeE4luuu7uwPdgd+2569BJN4EdpFzeOgazaUox6SlbMWAls
KMKvQMh+e/pXjMA3lCSZLHXUm9mZ/AfQAOdxrLnsJBKkc7Ejw1SJvD1Q5TU5uaM1uA3WHyvkxelK
XzBRYnVDIQO97bLEn1jRKj52TuRPOXvechG/Qxtsen3UvAtTXNkYGHFhbENp3IkX2++uwkjOJrrM
tPYOpPnhOnZfdfW2Qk7j1OY9uoU3wH7zB2580D6vNC14rHubEXW9zpA0CYelClaSraPtl7ELtgAG
vw6zqsUwYi7hPbyE2/AozhRxlmo9SM1ziURFF0RMufyGKuQy8z1txATtYB6qioCNS/qVKWzW4Ki0
vra91lTjfidAnqK/DotOiflnCXHYZn24K33JHcS60zkVruYalf0p6IFo3vUaOc9UN4L96O8+TpYr
kAViZeqH2IEjd93v0v2WeAFH+HwOrnsT5gwBbQu/8WVimR1Nwzyt+hCOyp10OQuE+El0+0PsyjmV
+X+9VXmk8oKJaQCqVPu3XClODzzlBXkiyQqrT3feC/ecSshMak5sronXI4zGcXga/ZIr+2l0RupE
ZAm1SAok930hONnbOVd0IY3PYhSPvOemWXfoipu+L+p5dUgA+4W/K+SS44IbO7MlwIAqSVB223Pt
3lX+Af+CDrUS91ot8Aqf2S1jLnqqhTACL/9eeLm+UOj5VYdiQXVyPpoKDvP8/7VHN2M56o8mkNof
Y6thBaNyq5Ii1Rv6GOdvg81V53xbrKrsOZPXarQo5zJM7UqLNp2NoH5jlsWJsJondQ8t+EJ/UvJq
Qd+FLlczoHu0PFT1nGNM6O76/z+iZR4liENnxD/xX5xUCqv726HMXaPbOJak/vJ3DIJ1QC+ge9bQ
ZH1CaKeFDDrKhCWhUFflVWPEodGlWY5xEuCFsclWcRuLnAic8NHwTjo+KNK7jNCIAcSSPzaIEK06
qUr23MBttS65WYK7XPEhyu6aF1QYvcI9YkkqQypGaNxbvD66hYsqainVe3Np01AaHKHjOpUo8UFF
rb3lhCf2RSASsauEzvZR6zFjHLzGiTYe3cXDLu4cy08yturB94cpMAiHj5AMMG1GaD8WqbcbGf/4
2MtcpHke+85CSyfLHPkpejn2xhQa70Mhl3F4WkTnhqUVLcmbuPVKgr7mi9ukImIzEPqSp3r5ERjL
zX84SpDAwoLmkl3JEN/+2oP+RWN9K+n/o/T4DjM0LvrndD+NmQQrm28WiZcv5sLgumvBKSzgz+ic
a5e9qdFfjwWMb+3XdLemUZ5OLnCpFvpcYL2PLSQAjGDiIS3KNgGaNYebFwAwxx/7iFUvNEIJnVI5
SOr9U44IKxe9zp8KzYmCpiIO72I6nAkf+lZtKCJ+miuryOQw9dVMBjr3LsWYw7V6LJx6TLu4R9Hr
zpt5HBl63V0kwWL74/NOv7ii0vDQy1TxErqK7Mr+KWRyZ00i8qCP7XomzyMdCaozqvA2G+E+aXeq
aYzQ+TAL8e0U71ZOyeQ8Mbvt1yV8m8w5VYEWWYtC8VRoJQK8tHCek7XsmyeefS0D6PExQ2GY1j40
pYfS3ez4DobF4EiqwpkH73FZZHIhJep1dGQ5TGT6FoM4Unn+SsoZ3K4jq4BQw/UZgfU7tvmjbvv0
cwVdOaZies0DrOLYEbXjinPOy1TiFYHeZlgr1mIxElQ6SkJBby5ZUdk8X+4jqfXjceHAX2LMcX/B
oikrTE9Wq6alJn4FOMxRENqLXScNKU8c0SddlSlR7LQQHax22cg2moHlZyBH4Y+aFKxZIbJd8CsS
FbRxNPpbqvWJzyzyY0spPyy+4SUPjUZ+Hk1JklvcRIS2OUd7aA1ZHlpgO8SH6cLtJUqwkx9GHH7H
JpPN2w2bGk8Eh+44bt7VN6S0LdoNGWNftqjwzKAi4lZwy/Gj2P8OzqsyREJ2QLz8asgbR42um3nP
YZCrQh0uCB7ofISAg+bJyl2CsL+Z1cinmU1wVSp49QxfgszIjg97kB5PRTps4JoAw8G2t3Rz7f22
w96ONzPd0pX7yQ78tE1FQF//SR0uTsAUFkfzLU2gGa6WRrUydpcKYVgY14sSZJgwPNs3I3HU89pu
m9M+LIlOhWY7EPx6DwbhBzB5yF+XhKn3nhYpXaY+qfK515l0QErgoimoc0XJUIcwm/5dWtIQJ22k
1EeYIbVk7oExUNnB8X7F6ZhgO1AkUWILHvicGFJS4W6oXXpgJhJhiolL8f9ubkM9gvXWJgkttxcv
4VSsOi1DSQsApSPtX3girI4TQ/G0ktKrWDsq0G/sWN2LvjoUDmhk3Glsrvj183+TIuwOZJnlCiiP
2dEdfsB49hPZdDXXum4Ja4nSDnEIYfQFUCLC3xzB8vmqcU+npQSRqvBIQ/BI+5Do1J7mYCXh+mv1
i5rA//1E2ZPXV7LfGN0MxgdxxlHedFHyk5UyQCwuMvcRG98AjAtyoPirQw1jcc4asrcA0dYzfKmL
ReGBh0+/pdDbfNt4MAX/GA+fI6Gk/xLCfwuxIryzyoI3knnhLroRjstMYnHnGNsfrr2z0xQW9Krc
5fqqISiOoipweTLIUlbP1oGuAhLwXhqcslr1O75vc62FgweeO6H2ESs7GhtlcuT5mic5Og43koJo
HIjgGiIOIMu+c3+9rfpVdo4PWJ+HUO4U8LJrNL6rVnq3F66FwByHB78gYSPq6g9U8Rcb+2o7oquu
0TAseJRC4yzLT4TtOQsrbQD/ZiQSphsxy+UhuCsiM4N75UpxnxkSUinIItl1JlJdemAc1ridz25p
kHV2LNi8NF+UUymAiV8P7Z47If2kurLs/+TZlI66X7WcXLPi+WZsMFCie3uh1y4pn/+piTLs6NDA
yoOkFnxpLWlIBrfR5dFSEhZVoGxteNg6vOhOa0DloGGTpA5lGw0zbRMC3gnnWgbxJmSWSSJ5Y+ia
uYGFClfIn8Fij1USZdM4AdPU9BrP60WuUJkL2i35psTGt40frUyq6XH8trWgwlzaXPaiOtNclL9P
UAM2F6m+SA9LxVhDqIpQMv6HHa2CBuBtRVRWDnpyYSuiq/uLRgSYC41+QRC3roUKSH3rXNBRlNAX
e1Lsugj9jRwQSOZH7QYAVcu0QWi6hl2R6iHEonmHXdHJx059YxTa0qaz+yP1pqaJdoLjnYHdrkuA
A2cnGVbOG8BM9DHDmtLHh1nXN9sAC62/PY89aJ+UBH7cduFbxkJjKVJkBuzzwVb9lHQYcYStrcnP
Rg0l0lvlCX1C0hHK+HjX4J/Dj4MjRJkoq/a8bnPQudJWYiRxsIJP4r2/gEmFSMT5lEE91By/DcPM
RssTRfsClVy/x/xh08E51ZdJOvnDQVCc1NP0QYdCTPQSbXDDvnq0ILpVnj9of1lmsHAUDvCvR1MK
lMsanCs8GOoo+/EJz8zRR+gYo5ZDyQU/0ufgXLzrAEkvG8eiRnyHY0d+vCbzrM8kpLi98qFWTTQh
uhH55Jp03p7KbNfQ0b30TOg23wTYo4KOKX/b5Orr+rTSGPP1x4amABYTd2r5Kb14v2Ixmas4rOeq
5RZ/QnsTXD/stwYaF/MenqkYpkCGDIUUppysxXRHf+mQaIEUHGi8FIWNz2xymxTuY+Hn0oDJyfIk
RxdRj/PJOmwqEDA7i1SyGg3ar5TQDsGdSQ7NAaZAreIn0o3bnoRiavy4hGU4OSrfzGuAyhrglFHe
ywZNq7r2oD//5tgrgZ6/5cziUJy+u//lPLxtGyDDec0S/ZOnT0Y005BJEPWGHmSiCIrIV4OAsKUT
88DmNHSRlJGa2GhMC/hUS+xT8SzQcHqmcYKT5F7U0xKaBZ4O+nm9T57gkg5itswFWp+p9vkawnY2
eFPSWJMvKgRLo+EG+DijCAgSVOw11okugt8vgi3yjtm6dMj+iBPIae6ExokIriE0ygmtGNGzwcGC
3tRGZE5jBG97OQRwRRoA9WOGLy2gKvUQNgh4wdhF0P0z5I9yZ45hUumMX/FodkZhWvohYpkv47CO
/QJgT2gZet29IgQUkPlxYx/Mji1rGVXvhnsYb3kGkOivdOSkpqUCQLRyUcT1pduLZECjRJELDcKP
qlmrRRibcpDcxlP8Z11RymN28LfQC+hWb2caqOW3jISoz2317H6AiEsniZACliQLjwdjRTwoB7qx
MI+eX8+y9LzqfB0qthrnPN78CNmIAKIDTS+g4DtpKmf42vPVRAOh2U5jNn/VyDyVdUHlvShH6IZd
4gtsyO3MVvdFwyuy+GrhPybg4a7cQBdCA6AaU+wxQXLZKmD1RIeMqA/Er1oEubTd26KrVxCIx2M6
rK9wp4lBFVIcAyTui39shBQZxUMFEQxqpjJDUB9JV7poOedfPQesz2VSXKm2iuksiFgl/7ScLKyM
Tv6mVaPh1BRpXqpDqSBRXmiBablY6ZXVPmbFi0mFMYt37t3r0fs88DSJZbzvO7rqgCe0ihvSWMf1
u3UczlQlJJ5iVDXejyF9qQ5jx/NXUCZX2PuxKVtT0eTFonXe2aElSun0gU1Bx3C4Zg632CJmuP1h
v5DaanLI2+aWcC7udOiykKySyN9ZCbtj6RhrhbGcpzw04vSCJrcm4FJQtvzD9oEFr87IQZdh0iAU
0g4vFvalxtcp1xb+oIcoaf7eOCwKmOKxfjc0ZFE/JTCBqr3nBd+wZZYNLVTCpijQiwGibE2rwrcG
sl0O1AncsjTRfq35UriB8ZU3OZ8cF5pJXzTS9ge1Vyp+Adpv7fWHdyrsvfX0ZUmhPktgx+QLB8pR
cY6mO5gVZ1kkofgjbeG8nKUubO+UEFpEQxF9/bgLTybB1f8y1s8G/XjGQEBCM4PE/vwpk6Wea00W
gc5M8MOLVlUZ88UGFdvFthUY1xFHKc4KKSHFHdsoUGFsYuO9QEavaljUPk9rph7uyV/W0kJRMBEG
MwvbHg9uCwSszcTjrAEMcGkYpesVLe/SvtGfDeXnxSVflh43uwiMtxXkHfRMQ7xUh40EaBF9DZ/u
5HLIqd73rqI78KV+xEIMyEFpX3BfgqnhyfBgsRIikvC60xiL7+9WTMs79mVubqTydgVFlO85xzAG
mNf6PS4xsKfyRqX3qoL9730WN7d/en20Damg2eelnxFpAA7zYvZ9B0vmOqjWoAo0/NkCn7xTLVQj
TOCFJKiVAsVqPja6lfjmDDLonvMDuEZrAifeLjfQgi7vDDQ+1+TJgqRRymICx1q/HmYIassAyXs4
FzfdaEqxIxjUS9uhB9fi5Xcsg2a8z+fU7BQV4MsGZkO9nVEy7Edb0S/LTaE/AudhZKOuVVTvzIJ5
61Y0ZVPvcFagU0zQOR0xav6bDrQhwmJrrXWuZnbVF/sV6WSRmKegf4eUMpurQAEcfI9OWApA51s6
EG/4mjioR3adnTw5kE3bjTHieEcSvlRW3evj3eBjwHCa/sXxrwzq0maSblGqFvA58EfMptSY2HgO
w6kon5Axyqzj71W/e96Q2axtc3U2vb9XUx8lQqKSPQqj56LlX19mTkxizFHgSDvzGtrFdpOwm4S7
zhvkscw7+kUHeiXWNrUP2tA5ZHMUtAydT0fNLUBuLLH80sZFf71O6e1gJnsTvSJgB9isHy70RWx7
H5e/0fLkZQ1j1imFWm/OaTDEvtdF5OWjEpUT7ZFaHw8FYf9FL+GjnowKAykntNtkULXKv4dj4mhC
+t96qqKpF+5lnR4JUoH/TsKjvyPFI0hRU2tPxp0HTCf4QO5Bue6FuB6vRpTbVQntLyUipT4leI0S
pLl7qJqyMnCOcEBFk2GSdqBTDcUVHK+9iSz+A/xEPDdJvNajyg/p0qcIuogZti2kXQvsTsUtHzc/
yEs6An1RadNTTtwASaDS/CLBUKDdXUtKlO+AH51up43vH2bAira6/0+MtV0Ui32tX9NHIhNR9b7v
AITWs99D2e0hmL+4oMOz6GXgZlerwdsY8Wno1RIpwWosv/AYrAeQ4XUXP0biEjIi7Qe90i5WJbzN
PtwTEbg3dEBwfYIEETBizLGGUSy851BGKz3XDAUL3SNYj1lN1m6PXkcXH2VfLUsymGwr2oS5/pWn
cYE34M5Z7v+L0YcCI436QdrMFXcpyQc8SLt7ZrFHFVWSNuNpvoSIzmSgMaz7bNnqhVOucGC+OPca
vukMAC9Gg592htMs/P6odf/tEwGERshb7CiRXGT5GZhNnBJFjkbEvwJZYA7f1XLHV9uU2MXgCQs/
FaElBnfLJN6zYVMccEvWDnZkMWwM4R8PkMljiK8beyz9d5DKlPP0Le108NMCFE/Bk+4IPCKZwprS
/wNyr6nQokWhal7EUQAHimK9WfbR8KQtevY9sUemP2DeYzW8wp4zTdmh1G5TvIeisR/n/85wNh2v
NI4Xhn5M9lsAz12zG+LeYRETdELA9m53Qjk2SmEZRmoWDCO1W6XW+hDeLSA4IRSswie4Vemeq8Kj
DcDsDS8jaUHOrff8FziFtmhvhTA9KSNxK/Y6YwzGr8KKExmRkoMvlslQM50uA+p1We3LuTUGkRRp
zHtrHoetN/2fxKlX9ijkZuePBXDZllwu6igYeGkngcb5FFn0HSyhydQxySX7d82W/Ct6V5MhoXk2
q5VwkE2q3IwAZa/BR9NE8y9RJewP9lYpTVsyxgRUXc4IetW/NEmngvBaow7ftdwHsH2z4NLpNKqh
twbsxO14rjJm38aJ3oR0y53Qc1mXtiCW1RtsPesG8Nz38t/bvfdp1dUv61ulML72eTEdiN/3gZpe
YSSQ9R8BeRk5Ilylv3RVywA5f2j+Eq2u8y7L6M9JJ35Yt/rN9hh/GXqn1iE2at/TJhoSR/nrZVhY
p/irWQYDMa4bTbVn6tayUlMIE4gmxjpZTb3931kzGUJLfQB7m/QFb7tKIn/U/g+NBlu7d6cl6kqP
IOpJE9Xyz676IpLvHan7GaSRamutuVrm+b/cOyrCcsfbr1OL17wtn7K5qt+QyHfQoRqbGz08Az6D
pTTeYW6qP7EkQtCDdttBuKS2eY6uRmmhZIMarQ/jxachwBRC8rYD41qL5eH+/Y88yUI/SIr/3Mst
58F8HsiNJRAYwRjKlHKhUJvKzomGTztzJdgI3vAsKul15SBuo7kOThfCin7JUwtmwil/xaPevV85
8+8YjWzfhKoRhtLQmUyY6g5Dui7Rz0jT5rKXc+PoslKc4+BKW966V143DNICYIu+IdsB51jO0u9p
iroUVmQLD7ytkKVyBuTZb5rl9wwNf1KqhYgyDA/1LJcKMOpRbsu40JZEGC1f91r1hkZxli7H5mdv
g3/WNn1If3tthYaHVjFM3doTCClwt3RLQdYBHw1D9jClQwBAjgge+9EjSnoLvgYz/NLLeMGgy/4Z
8Xuptd4ql0JJf/yPSRkxSpujoDvVeW9O4PhpbqsS0MXsw5xDDKlaAL/ToMy5vBh47Wc+1If+2Qmr
cGUbg3MnZBvTzEJdTlqYwP5i5IDeT/P+d+0tTarIJ8YoPnawlZ+/BSeepdK7dygF4ZQ02n1sgByU
qIl1qYkzbumYAxLD+WFPtyYZyQch1Hz2xU453PWXOGuQDXqMFtUUqijVxe0ve+NXH7LUnj4NGVvy
VNcEUCSMqJ2KGSrKv0HJKrYV328pe8NSf5oRSF9t3d1daPa5Hxq85lgJqzVoNgAzQHkvQEERayow
KbIzw4kwhKUIohatGY5rDGDALhSla5sNTub2Cgl4IUdN4fEAaEfLQ+o7o9Uq/Z1gVLPznmaGhpH6
JV4xVZYkqzMowJ9eLyelKIvfqJOHBx0jjYWALmzTXE5WvXltPqScQtJkL9Ygqkc9ZjJfWLkQOECh
PsM9C3bta1ZCbMpYwyZtED5ZU9QhKuJO4lzlPmFuBLOp8m9+Y6UmRY25iEiduOZOr8i+bta8UjE9
lkl1hw9YVggBiTngYrNMLleTbD59A2jxkWID78kFtdcMPqt9ppoU7XYhsGrj0VnFyPch6yWL4Df/
v+Ds4zklfMfZSYuhHeZy5XL2/mkLowcXl2Tv5nhAg8EdR9QGkWyQv0hhOfQmgKybl7QQ3TIsV1ZR
Bsiwrg9lF5X6ekLZOC4K8/u/xQk0ABTx+0MVWrm7xIGnLqdNUraFWcayBwru2Qt2M6bkw/kNV6Ix
vomgcqIM8RS3dNFOaKFRAt5P+UVCEHpgsFHb7cJu1wVqpNl/V3nfV50WLcWEAoj/qduGtgvaB0hv
Quwykx2m1Hj1fGkd3ma3RktMw/iXdfAGa3ovmX8B7+e6XlsLk3WHEA+zpPZnFhTgra8QbcabPuK2
ZQxO7ZZKfH6kULXLoX8F3Hz++sTBf2ZUtmO5F4Wb2BUV4La+Xhs04ft/jsuLlsCc2zrMd3ojrR13
3zd2qI1sdxEJ/dKaA0OL3ahf7q1Vz6cVNZqCDeIgO4Uaq08rZ8rWaOl347HjcH1InAbWEMk4xfvP
N7gQ9M8O8WR9iVCQgSXvpJ3JeAKvWS3qeFo4Tfmguo3aLkevm06zs7ZJ5OC6s5a4nh3u+4QA7kVH
Ndt0+ErIcmJ1R+o8xmTzvRJh8nS1gxJuv6ELsd+TebEzFjFfwED/K2BRKM7jq7XwoavmVA85TjtA
Pl5x2YwhSBnfVrl7GJP3PEglaCkK0te2NYKSh1DKtAwjYmXQwSIVInsgytKPhsADdbDaSpzs6BGw
e2dOjG85neibg4gvT/EId5WaQeGp01Zx6279ED9NX+/Qxn9KrchIW0NxwdWGMmqpV4KCLKQSptwo
48JlkHXYQQaMafyQJYsGIU/rQKUddXW6Xnjou0rdv/slxZldfKw4rp4DLmKHhrC1/YVZrTT4AUGd
1mjH6wQoYPyrPa31nl2FAsuW4FgqTbLUdgqxXxGKEO6RNpnFE2XdrhnGpnpgosebn9q/KRTV825D
442UP13lP9NpkRaBL1oSs7t9YFeCf3TKwqMOZJRfNQf81UOY6uaUEmk1o27V9x01fURBSDOVbCQs
r4JIs/f0hKRW0d9Kvm/cwu1//N+vs3rLLxde1Wj52L584SMqBUX5D3GbthqC3lX8lyb4kJUNLUex
6VvEDspBkiEBNbXEnY5elHDXwROhQkHOdcecf/bn6CZdmU9qI3KqGcGXX+JfhinbwX6Bc1xmHPum
zinbjVyE/c528YVe8LygNMib4pdigV6Vmv4qhjJa9HEVZb8ugdCyvTKpo/MkUoAUUNODMBl/MmmP
pHG0c3xfvTfa+UDoJacQGc1JyPQd+JkFn/BzrRBZ5nU6vQ0IFHs4a2FoLgevg1fivEqXoX68elwu
NDer+Y2yBa/wh/PtpQWf9+QpSrUuJtH6+awPyTK/ZSHMVmGj202vSWQQqRuAHeEvmaOk+mgoz7an
cP6Fw1WXoSUG7qGzYAyDMy1XLk85iPmBK7EvgapOYZjnTvua33zPSjIgxiJlcTnADj5TNXeIN0F5
MfaXR4w0xYP9ZD4qDtqGSVpGLSuqQU82Qj00JYD+zuSzBYENXB/+et5xCZc9pppuJb0CmRrarhyk
uVK5z7S53zWKvBMM/7Z3c9+TwfuNhlpUDZixgFBahciuzsiraYIbOoC5NPDanORcN5UiUbJHbYdZ
T1padP5eEUvdC0wP7Y5Qn54mIVeAUYja8buZ4HqxE8z9IFKFEM5q1AB+EiaC/+HLScl6H3ce5kYh
uq92nYi4qME/L7LYXwzeiS5rmajbs//mRGvaT7Q7ZopBpX6mIWFJrnr+KdHsNcO2o9bx3xVjRpRY
m8XyggBIfrNgWrWfbw0u4h9Wk2XlB15DYWW3COhPDBnUTQDtzHilSHK9Kq8zys6AlGT8ZVq3JZg7
33l7+Iv+OrAJBspTVQJ/3spmQ2ZxVOdBMdScSoL6iPTcnsHWpj1Hz2o37iaNnS7+wFOajM7KUXso
JyqzHmQDRq71lxEumAxuvJ6YiLdrYxcg5vynln/B3IzuVVIuhZShmgom9RUG7qae/k7K77MpRuhR
Dqtvku6Q4iaK6Kd6mzOzd9QrVGNM5aZB/GrKvzXoA66VU5N+G9ZauTFrMBoMtVqJ6HMlplxrsgtz
7xp7lNABjLwv66rnx5WxYC23Vjf5H9Q0zelAG0Rl7q19tXOKvzcHilrS0wu/NllVUPpJqyerG788
I/tREcg21GwmDM6jBHb1wdPSsSoVKce5fIkMb1g6Jk0Q7YeM9lv+vx1lGJnHdPtnzLz8NDSiTUkl
FK0qO+wMumPhhGGNaM8BVWS8wKh/DiEB3YvtOwJLUPmr5Zai1P5Yx4Si6ZOO9kubTkblIJ9cSv6p
GhAR1prPiD9vGf/YSmM9qqFWJXFwK73LmMf6IaqjkwZ2KqMzREIWWLz3EMT1jxKwr4ANZeOFiVZt
n7/lWpQS60QyzoZq4Zhv8bE8b4P/zwGocth+cy5BMdfMVYOHH3u3C4Y20axSQiiJXZlRuCC9l6Eu
PiPpFEmmFr+Kj8hKTRwp0kVyGt/v5VC3kE+vQWa52HWvM6Ypg5FpeM3Lnbb2sq9X4vYctaHZV2Jv
die/4CuAtuxXIK77PqRWVdZ60b+o5qJ3K1ceEq3PEZ6dTys4aQEuskSb0RFM0gvsFvZf4qF5vCmx
Mx6sCNb8xQVXET4zrOh3Y/xMFREO3E01PRVRiQf30x27s3HVr2N/4n3KLX/oqKz9BPTohTSJewMa
5023WlSdptSwkMskMFyaYQgSMlCdM7dV9jIIVw8cOmO4kVGIolSuFtFV8K1t2kGnv+k91f37pn5L
q03l8ATLcF5GT0YdJzfcyTmkXyeSOw25YfVapcEaIrYxTPHgurkYbMaP9OeEZtS4qYD9hkJZ4mde
spD/dUgZ9F+OSk3bP2LRbN1/XQqzyKN2aKdTPDv2wnIqYghlfdeSkpNjG0p/SgSkW8oRMnMZTOoG
ttuzQp3Y9gel+ZHIfnN1DyHMtmq5dSd57tD1VHJke9RFjR/zbBTcwzuQCfCfao/XvkQOqdzg1CIW
oaMZrSZ8AGVNph9xCP4Pt2jlE9CRnDdxbxeX6nM8jzX5pCEU8xZ4kCdOgcXh69Mw2yvXYIGRDuZl
OeJTtMNHnJTXcMIwcv/A8blMDXdqojXTiaMFBmk1cxHFVONdZjEn7ezAf25AUM6Gog7RQBPNGcqN
eavGqZ41W+ALC649n6Z5TlNRfRDxQm7DFU1JjKeZtMn758HYaw6H3EPAEPDdKb0fr6I3wR6URVAm
BubSpTJxM1Zv14Eb9yyX2tMVmnrld9ZnluXyTFs4YmlnYFvjDzhKQi2yfRNgvZJiEUIVMxR5kVcV
sagrhW2sucJdHQBUMHScAVwK9d4fYEr4A5bcb1CvGoYdDUyGXy2i945XXV4+pUomALrqSOhQGgLr
nQu/G5i3AiebuaqMPflAGJt8VYzjmOfV/8y/mh4Rx3leqUi5kFkjX3yLrZbJx1YTnptjIYbceKMo
UXSPVcypxvfHCB9JGjRhGE8kyK+rddQYu7fB31vYSrT4tGZtDHYSu9vdWnpNt4ydTTdj6uHLGh3/
zMnQAo8wY2W/aybPSBzI6qVlkRTM2UxQjNkO1uV2KknF5J+TZlEnqwev7aloGQBStTAB7hu4GzpP
Gmcc0Wn3Bjn+VFPEH5Tjhfj9I8xzw+fMYK/qH/BXiQvqAGr/DPVNfXbrNPqGuJUbF4H8sQfrD3GM
voJw5V5NYGVP75jXtaFcm7hgS/ZHY1w1IIsMrWDX22sltX7/rFE9JboAkEHZJkVBlfy+RMhBmxMk
bXHo+gz4pICZ5vNhfRX0E2AXIy0v5Ks5E+sbJiWoozWO+E7hjbNOV3Kjb6V2Ck51NMG4nJXIHKZ8
VtPjL687W/nYgvAcdVdY6nTJiuVe6oHyGiXNsrDnXCRW8O/3OCy+EIxnxGQ1zoi7Ceaq34ilKdnk
I2AD0K7VKq2PeDK7DuGOKn0wATqSSxkd6foiMFENsylgiGUrDNyTUJoX7CEAUrDv8uVGHyX89YvJ
L8TmTZbsGC0/itJtZ4RbM2u9Hrp4WaiYEwrBKJZQmEAyL6VXF/2mcTe5FuqSdarNrm7ap4NARbwA
bjZKT1CnSmGZX5BLS3vYN/reJWTpavT7Joe1e4OgueecZBuLZzBZ+UTjO9LVYRCWEWAlrzMqdFyV
f3joIne2I9zwrF3eHuUxB3QWrF0IGnoWaTaCAsze4dUpYvLct91cinIq//capKby4fCPwko5yAog
uPfhSy69Qels694BZBSmYNy0Eim0meKus/jEfjYd2AnXsAhIIUl44FHR8z4mIoYexTRaLk3Xl+QG
1SHOgZVWZ12MBAWT5ESD1k+HQA8JHsISfuh22SC7wUJ5+tX7ZOBJ9pDNGp2829a+rHvrSSVAfL3h
0rPMWKupUf0zTfq4d4vPrGTR8I5dfUC6r3R1r1zOYF1df6aZ14t08zZsJ6/PRXce8AbzEwVQ4hzC
0nVntT8BmT8g0QU3wkz4ZG1AghZYPtL2HBDW5LGOi7WNHe/8OR3kNu3CwrBe4MhjgNrvOF9rdcTW
ls2E9W+hW/XL7RcXU7EPBHAfP+WIofGsB9258eK/6k9N0LjEelnTtHSvQ3uNcp8K5t44OKYkmz+U
JwzxdFaGVTfhRGQy9dGXwfRXNlwM9/O19KbD2WFAUabSGY7ErBCY439AX+Q4bHpqmop+PP9TCilu
61shlAbwCX8XmDRo07ntrMrDU7+IzkooWLzr2sinOOH0s0hAME9Ms3le2NqVR5aZ88IIMMIwj+bO
hkbnXfob1uuByqmTnFPeKJy+W/+VXwFsLLDjp54EYEQJyjb8RILRu86LLy2foNBNLdtlLyFcV4+z
Mro/1WuMSLLwvzyUJF4z0Qn+87q6J6L7FKOojhdlIO7JdYSDjAFDToaVrwYnspPy4cZM8VmU9tIg
JZOD7/wI9X9j4ReiX0IFQx1KBByKbfy1vTm8WhQE10WjRjM0wVm8qMDXYF9oo0Xv4Zc2+YAEwq0I
uehgizhfaq88oToAppOz3C22pGy2xogoGywabIStqR+txtmM4xW3tw9Kl+Gj94tXQOOR2x0h7QBe
QEyAuWVMBdl+Un6RnVmFpdyDmS90fuw520Ud8jOLO3hH4RM1mOJ2YHcAmNiZom3TzSPtHoOtlzy4
VpjNfVS/wk4jeCpOYSPhS5dVELYiVdB7PYA0ZwUhRWvI57oKZwS874bj+VgIWHULfZIo/i6ZnzGi
cV6Mb2AiwCDuJuItnPi/62Vb8RyqKtdqz6TUY3mRjZc8kMVNMgHLAL1mbeqSY04vkT0nSpsJMXvo
XkJQqivX8s2fzY3xa4dJ+tHhKnp7rF5cuHEw26OEVEr6aGUyM2F6qxTsFtnepZzimZLaYTa/QbnK
H14soRQhXqfQfOeBFPzNVZGo+P7sFUXb6Xfzy78fjkY2zYCnVHs0PzXuSIoh3WGtPywCbxxn5+Zn
YGdPQZOENdLaLpO8LerPDojeQA6fNY3wcFV7eEOmy6/gqq6/wys1apLVce8PzcZI3KOtc3cw1QA/
4kDd0qUmv8Efm8Q36Qu4TVzIGvF1Rp/bbL6icqnAk4e/HTvPF0nK4jmvACwWcQz7t5hHlGI0Vpo0
e6tyc8Tn0V53IVEXVKtVzcOCKHSxuv7iawX5MuN/nDSE2DDM5KD1Wb1gqM8H4Nobh1al3ixjHULC
5ce/g56gwr3+BePMS0x8ixsF3jPGDo6MdZmum0pCGMMJZv0oKTKbAgQUdI7SzPXKbHbKfONsvpGj
Nqr/7/Lnz/YeArDINhgCsFqnwQ91QXcz6mfUgvts4Ew6ZYpWmrWHmy+vnwfULLygIRSl9OEeGyNd
MI+c+8QhelGu09AciqEAxsO5CyYIbb8DccdSgKes5NLZ7Y/+Yny7vLwk7ZFOcB75L9TfAzwz54z7
qX3aCJZ0gnDwJt04u2JJ66glu92Ebsa55hCKeFUIQVLmQti9r/VN9LCmgzc+PmYIpHBJW1InSN9C
rcmp/eoKJSpW85YwH7sXd6y2E2+kET1i4Ej6xnYmjgbAFsTeQMZ2vKFCzkFGxDcHIADLBkUtIaTu
EApHwO+9ne5GNUW13f/IdbcLd3AAUitaLNk67WRciq4wNWUVz4mBV96cctBKfXHx4zAmchsXwxSJ
PyUXtEeDvQWBubDBFZhJ7oaeBSTXMFIUd/eQKmC1OVfskslTH/5y0x0Vfn/9Nplba/SbnzUqdzC1
+QGP6FbdO7EPB8SVnusKey5PTDx/pvGxPZKgKI/xQqlevOLVH19FfP+QGb1U5pV0lDS/YCuIdadG
d1C/21vyhJz2ZvofrVwRA0CFWxUhHa9JojIRTVbYd77eUztVve/ps2RiEtwXeG7UI/4SPRpiB7iz
nCL7O0vAYDxSbxS83NPH7OFdX4//hbnda8D7oTQuIU2iPLkTYf+9XRwptOVk355hmR/TxwJxF3tf
nSLEIxojbWjS1slglOa2DJDykSeMxT+jvM65ZbmKLm7H3FriMlKOESsOn/E7qSz93j9qpSre5xZK
r1ALUhTjeJipRy1gECJ42fyi3PkUv2qhs82WcKALCtU95xjFeXaySPczG5Bj2NE1kp+OYmw/+YS2
KZtnG/LQXYvzA8XuUB2au78wIx58j/okRzwW2lZsa5M+LVbGtJVzvdzavgkAHj6xYfeZZPVN79zg
oDMvplepD6POlejLH7O2Mv0+QqSZwA29k8AKTysdCflkiwFuIh9UVxZRjH2/Ss4bmChDbJgZcmgE
DkbOY62H+YMd2aR5olNL+r1uJiSLXp5/jz/EdYSmxEfZWRAzK4/OE1D8thc4j4XCbVEEgCw/IMAU
URIPueI6mMmLukrj4cuGcoaYGTKpy9Z4pewW+R1AbTGjBEx+5zoxYgjZt65clS+dQNn40P45S2In
VKDJNS04T72fQ1lRgQU1ob0/N5gcPcNoxfJEIzo+2lK0l4WD91AnSLNs0hEO9NjVJByc8YnCOFCg
RoeU7uhxHdQeQ1MOlEKL8mFhRxLAISlAyKh9iYUpNJB6Dez8seusOosKOsPo4TV1iP0Rlxs7JrHs
RmUd3s2xzfGVQDLz/xJvVGd+n/rcRk/5rHovQi0VOlfPAhV5YfPkHjdnc0DVN+VNjaBHSNq1LF5U
8L/m0IoXzxQ4oUO9XLKWgcYcQsxx2Sc9SS6MioP5BiDTGctVyeYQS1u4X/ZEWW662XZWNIHMqtTW
4ofb8JdIAYlYekNXieeJZ2JFpwLiwCLzIJ3dZUmawDpjy08tH4gQHnFpN9mmbwXOqzQmLl1n1b6l
UdtwL6GZ8R9yLwrhSkVOUAPeXq8FoEEF1H/1EhRqE6JEMrHCOdFyGD7Nfu4UhY53e2RKUkc+4idd
+bGkTCdJgdvwkbK/29Z9sdcpJw/jlKjSk3V8AALksGxm6WD+Q1gQOsDvoF3vivYXqMq+JM+oBW+D
Om61JrMVGDY7VHEarMktGUOBMVqg7w3DAW7s4dwffc9K/dlAmcWRgqyFwOKBwaM4mKYcn7QPboPl
RXoe/+F12DaMAVdXNkyhozTgIOeDL+kFGAMPkIBNDPeDD0VGe9dxXefx2CBABsPR11xJDlc1zvLu
GyQvWxVkMUYZSNJB6Cs/Hus9ndaCfeP90oNhHkC8a2upBiNhvaKZRWcZl9ytm6x9ZyrezqTPxXkt
cwp8H56HIwvHJObnHWVtMLMPnEMNoyHndpDb+4N0Y50lhLHohkD3PFpXZ2bVsrDLovEu4LTIYhMQ
JE1vDG215IvLlGD4NEPNrN3RSBN81FNbxx281xCu+/i/2mmYumuEtQtX8hVN5eM9AdQzObkIaaeY
nP8eXdL4Hu75A/nERLB5ABRMPaeGeLXIPp1UI172Lm0jccllQ7XArMRAp701nRdvQfNGgQdzmibA
OD3zDcnDLktA5H+DBeaTts9F46N57lddWNlNl8SnBw/1/G2x1ojmMQVycyHwv1op4Kjz4i1O34mp
gytiNSf42IqOh7ZJPyLdP5CH8sDtDh+nDVpH09ii1KX3PsvgCa1Z9EzZm2bXF31nE3gAML32EZ4t
t47v0idSiZLNjtur3uGtGX7SwNZJbuCRi5FahkKT+tkvuokzl17n/wnECaLlfquqhDr+hjwaL79O
VuLktt4Qw6hqOmz1poerrx7j59LB4VAs5MnmlbiVQFtyHfX/QXVGCfM2/qVOXUs2pE0a5fGXwYS9
lrgTPZA1VY0Oj2yRK6uDcqQSgQRyZr/dIoXLE6XnLUyCyRSv+IEJw1gRNhZqWbOgNI87VPEiuM2B
KmUaOs5lsR985KdWVFgChxiTxJSDIPJ55+Ai2747Bne65Wfes3wm8gPWZHzHjNY4v+0mdy3N75uF
WFHj7OrvKV65Ir1Ami07aCFLqX7RagceNJ7Gu0eI6xH+STFhVJThWmeOu1ccDzu26/anZtcCBiJC
tWPbbqbpP7ayL4bzF3yZTFbwQVExJncof6yGq1Xa+Dj/kDLPnLIqhsi5dyO7ykz3xSY8/Wjfar4+
fW+QXV5AJNwV8jjOygtbPYT/1bt4QP8jRjA6lOLXWMPg6p7htoD6b8ttG4VOUnsVH/kLDThwAEin
8kDPA45SmZkb5pB9KpgarV/4k+s7eGUSqeuvvP3C0OAJGqEAA6LL4RiQ5JpSqUJ/YgH/jfOWJEIV
51lMg1qjE/qi8d8ttjJhNlS09vnr21kv4OO4BlsxCFvG8qxjrwLyfaBYP1Xa+16CNOXpcqBzpfaP
szpo5yrEXbE+sLtbjuS46k2XN/8HGyf7BlyQW97obuHrb97i9p+tBzsx/O3FchRSrMbGP59D6Vtb
LeCzq6ShGgbPZtOkPDuZ5HhdrNfD7Pd7NWySvgIgBVShucPlVqPFufm8Wb0MVmeMh/TmZvJ2gUJa
zqjM4rE2CbPx7UBe0pEeeHvttJAeAaxxSg6ZK+lFuAc2vvMpOhX8TJM/mrEKaCbQUGNLNempDEAz
dvvWCiJtcx3cHuV9oUkaJ7rF2JHM51KxKlvrOW+Q/oFAZgqGdZM681rtbxncjgMLDqjydp3wCUkC
AkWqnC/AFlj7ymqxWWQ04M4moG+JMRJrsh0DAsjc763bMSv3T3CTOfw3wVzvolWp4PoiCoSExgCA
qo1UroNmBI1NNiyjoEzLrfJHoceA4XxRPBr3yBMWJM9+if/fTiv8szXvRLs53eMMnKZV3yarshue
MjxSNX0OrVXvCYYFCTBBwZqc9QJ3aqvuMvnZc/djjTXL2/0w/RLm/3l1OIEMBUjVNCcKNXnxWVY0
QWxomQPs+xKhmKVGtHg6TB6uF6Pc1HPzsdj//Zv6IZjm2l43WFA5EHXDJV+AJiKsc11iaAkYTjjD
sbYD34Q+F/Iju6kdmlocoRdI7JAJ/U1xR11yaOuHnq8/md1lpgzSI74y+zUaPzLWgxzL+u+k3V93
0LcDoJrqUg5JPWzsIC5WspL+/Um59As0AhaXIRx0HmWIusG4bblpezP3D1FdU9+vD2v/QRb0JcIz
4QXOKR8prNMB64uZLpvoAwz5uJu/HdCoz1Y/3ClANu8gysLYI75sYFsUR0bXPhHHMg8HMFwOgeAx
2F11+udqHvB9cxu5dfj5eoIQnbgiTqEqS+0bgLt71lT2S56VbwYkblw7sHS8dL2Q0IIicHQ/7bI5
rZPq/EuS482z+q5FxMAQc6REAJXucn5gtPAKozGSLXRopHw8Rq/9QUo7K0nD1GXANsqP/AwWKnhk
x7KA9rDIn2mbHmCU7qvj/e7hEscWw3lX3HDzX0M+go0nCzMS5KeYt/XZ+iWdCEoWw7UhHQjk3Whg
QwSYlX4zTVihKt8TQudN8Nd5cNSk4sFO8L7bM26uTukL5FBNu49Kq6LiSNRkz7H/SyNygKrwMEhj
9Zir13zpIU4pkiTZ5KauEuQG9bofptAwr3RaBg1kfomsDO6omMcZJR3G0hyR7avLenAa6gEGekVS
IqpTLZXQc77Fd3Is0gLx0DrbbNnPqhSJyoYvA+zqi9SkU11LbHehPAVrH2RWCqPgoh+UY3m2lSec
dqRwXvN0fqPfeOSQG+lvMH9Dywj/maJPBbYxmz/f73DhKVuwsfnlQ6YZnRrSaDaqXfGQqys01mzC
7kNUkHEua2zlwzc0dviCa1yMS/SyF1ToO6TtGgBpZcUfTWMum5e8heNz82LwMhwDqYLpT9XMjuF2
En6U4dl1uhoOhn/RMZSETJe/Rkn3CyfkSwdMg+vDcVtT+LPSoQL/HlpDorMGVlT8u++Jjpkk5OeN
MqWgbVMnEnsjfsqxdXaSCAZ9FNZsDOcRpcO+asv9rAUvxgWsZmmoGaEIw6wzYcJRULNgLQrYwyV9
V2VqsQaECvFMOMKmoclTIsmTWHHggxkxMQo9ugoiTuLHCoSAbQAeMSmMbTS6d9gPAX2FOcWVjDuc
+JmpdnDh1dWR/zR/lmZgeVGmmGgEB6RrHZfcVKBV13huV0WYLvJJxA2fElksc0IKyt7HD+YUIjTX
OYSjPyif29ctLP9WWxdHDPS5BSiGk8N4HVRDuvI4I0ukf2kfcj7itM4j/qlNwCLFBhZHEszEZgar
n/D0A7U4NxR4FNjnBVGVKPJT2tYhhHwUfWPmdWsMQLD1dcFXlzMP0ZOmlSeACKI48wFV9t7WsfnK
bJJRmJLiHCyrIc89UqVNjc3OsmeOSh+Krzd3qsY3zdHviSsTffxDjjO9SiXfm6azhRSLUY6GaRpJ
37xpzzJStRHMFMSP2Dpopdc256qTuA/aHdytOowLZFnCbCQGCr/94MFZq8f8WJ06wqiipnlMcXVP
uY3EOUjWcMQQzoGz5l0BS2IBETkw2tDdZzp/OMN9GMeRKMLALdSyt0uLVWnpkYNcggbzpROKvTRT
Qw6nqasnQCAdo/HVmCAjk0l66JfcHL+nVdJ4YugdYP/OZfqOgwHSPkk5qk9FmN1Wz/2Sv0PQW431
OHB45L5Om4xDp8PlK+Dbk1Unehm3q6CjNojmKV91JX38VND2WokMNV0fAR8xSZPyeuSWWYGDM2nv
b8Dpr7fRuWwjP1fpAXL95gtNF31HnQwFnDATauAaO7phDVPW354jnxKXSp6feKhnSURjMqQ0UR9f
xlRCrh2Ev0bh2N6vBj5n5AIHan2ciDOjXTdSCWXPYAFQ1fjJRg3u68LBP2wdd+0wgDcDh/HSK8kz
fpT/aP6S+FjUzaYMbtOOkHIOieYbnMZrtF1CEcO7roJw8xk2AzjYGSW6gqLN0+52ySa6Ql0s60IR
A1gtg/drDmB/PUjk2zgR5cdEq82g/XHvaAjgXnGpG/TK4+6HBJkb6AuGMoiwS+7ZBOCbPurRYa8b
/G9Ct6L334k0cK42QSZw0MyWAT3P58B8gXpRpsYYyWpTGdCg/ci2AnTa0oz20IID7WuxnkNX161k
n05CmX6FAvBoq87bmqlcni244Yo1wQqE5SbwKJrftg+Menxmpfu9/XIhFozZq89QmdM8PIzVc3GV
ZjhIYzh3qVVmzpbo1sKFPzGC7NGAxdYHx1vYgZ7QDUUSTzdhQsWvm3K5kV8ygE78t86yyejfkVv+
4sguf5VrPWn4n48Bm/z7VZMDBKc4lwEImtxxpjmOch7wYLda/3mX+WvF3QCo9w4MC8L+707THtuX
NgntK7qfQSZGeoYkNnhRmcND922lb6CJVBi4BVaqWF6gH10RdMMUoInM94thTEJff/YD+NJPnIa0
wUaOBnrw8+vtoLrHua4zR9BGAQT6rS1jKz77ZcJVdvqFgop45jglCEYC4dWLIs7PdxBbyTfRtzLH
FPyenje88lT4tSolA52ZtndPIPufitJ9eB3/VQsigafdEQEKSMPbkXBKVjJB5w4JdnOk9HY4Tc7n
aja/rMCZTWso8tuT3Oe8k+4fkF6jBA/FHKJEu1qDU4tjg6nUrZW0MPO7KHmvNKWW4YXFFDtkrSWm
pqGB1DJZ0JZIcKf82acXwkU2pt6DUknEZOFeTKlx3PkjYSQHPUGgykRmfo1n1HnoA1QM282yiPka
IzDkGRfol7LcCeZ9V3qdK6sO/yJafKJhGj3i4oo0oFkSmiOKXqVN0Op1HqLkLJPxAzKqDA1gy1r8
cDlmnRT/LDjFN0FgKh87bhbayantmxWGoLdQnQJKdl6C3g/WOGqnwQhuuUwhAkuHX9MePSfq+3w/
tF5mIxwea/ip0aZadCa8RNagz3n5iCTCKE2wAZ6g2oTk9UqYnKTjjb6e3r35QeANVJKAjH71NwLF
WZSr0rIxtgRu4s2m9lrrxLi8ddeizRyDHZ5YiJKihFr2NLn1jtQ0FZFAQZAxr8tSpJ/BOHH8Z0w5
5QhoUSwUq78mOq07GNGO9iqb/kC5ddqBRRahiVawBGI2jEqClqlsD9Ku40OZ5ePQ66F08+JIqM9j
X60nc26t1/VHHFvxL518XN2ps4H9Oz0Z2R00kK2NLcBYULtGy+mqY5ZB+axleDHVEEPydGhRByyi
hXevUe6xsjFTK1VVA6VINtdx6N/8vBOO3fUeiF8lfTqDyj1Q+F7CsXUYqWRx52U+ot2i9jzWccwT
af+1nxGhtYWQePKHyCU0oQ++E9aoF/OG82o668OKNJb5lqS39Ug3yMlHC0OwTjMwaFIpu5WfmsAT
tuLJbl4t0i7qleddxUtAJ1s22t3NQOUwoSoFbI5JSwSghsPdN/o7TUCoBg6N5yVey3r4PV5UwlSX
vdDhJVIAtgjixJBkbaoY9wT6wPrBu7MDAEGsPNAqL3HwjHMtfDV7k0vFxnyJxB3Rn4UsJe5HkSJ7
gNXyP1XvXz8TMvxxwlAd2hO5ZSuWpNzDmjG6BKWhTru5AeWmbF+/T+EmnFE+EPpw3AbprOprjXRR
HmYGrMERunj1wZbkrKtJr1lSM8l6y4F13co7ijq1khgc2bHA7aiTF6oaVweNk1XszxTuiOlvRscL
C1FId+5wEE+Q/Zr6zeOlz373S3iPqWoJfKPlX4GQs1lIOWi7zTRAK/zFFcZEOlTbKH90Z393SCqQ
zy8pImQUTsGyjU0GRJufrIUwGOKnBuabJwEacKpHhJxZ2RML4RV7EOCTWACRemog50T+boDlhCS9
ZzCVoFuhTzmthGKmgXVKWd5WzXn1XByEyMBw0Sb2zXyb2tKTSff9+dPO90bkBVQHeOoHOBNvxko2
bYFEjK8NdJPHKyDddtzE17YGn/3xU0UTVyCq9dERWCzpirhnO3lu8Ou2E2myTYu1+5xU1hcDEKeA
zoCAKZpTuf5xoGEcWuDl7ByoaZwhnSU4rhSSTzebVwe68Ymw//1Y0+z1eouKhCD2KCp7Xyuj+hdW
tgxP6rhfUfcorYd+L21o1m9yuCpbVdfoNuNsdrbrUtxq10K7/P4TuId0yGtd5MhV56Q2fIegRzfd
yEaOwPJOHffa6X5mLOiTIZAeuYMBKhlOy7wAwS//sGQWtGMGe5taXBRU2z1yyrGoWadI3ctroloX
8tDt66M+SqrvyefznqJrvjBp6/ytOcB8BpKj30VnN1kcDAupLU9myc7CWemAI6Dq2ybcMYdoE0Yc
QVdNJxw3Dep983tanxiTDob3t07VNdK8kSmEQN9NUB/P+2pHvO/rMvSbxFQZFPor6CCds2/Dz6Vx
dq7LY2iDx+GGFJPlnQbsUXVD5Fm24JtHJsyd11Gkb9QC1egjnw1+VJVwYFkgkJXKz/pCJ6YPygTV
Quy8rzSXocU9yrBzm6lhDmsnkMTmGDX/guSf8GGefqdti0O5mk/aYxaxTtE5pJfaqoArvLuQjW6K
Gp95Xecs7G4ZnyWpka7hEyVqC5ztUdHzMSLnjMNnha98UXcWTTUCg/7AavcDsVZTJs9/Fc6TN64b
1EdQBXp94lHEE9IrDIjNM1IdsTJTq1oSnf4dAykp1bziGwQvXKBjmp3AFj6xtqLadmqSPdszUhxJ
9oq3dfj6gego76bg9A1KNm0hHGVJNF/RDUCoo+apTj4QziNvbqPdF9BYrHhihOUShAMG1pi0gOxY
vHjqMy0jPvB7+H+CMIGqYIHMZ0Co8+LKLzIfGmfRs1b5HSjE8Ni/yxDrfoeqEkzRcR27+KQIkgQ4
fW3/07f/eb7YJeJdnxI5Issvy4c9JpU8Zqlz+AiZPB2nSiDZ9CDko7AO2c9sDjmxUef+mgHhIsfk
RtDC5ML80/kGtgeOGpXKocxdZcF+brEmCF4jSmt0ZPeEEyL3dmpG+pl2TELc2HKHdswTAyAtzrxj
IyYPqGF1FzqeOqk5R/d0M7vBjF13A3e9lIWyc8MC3tSISOR9MhgnmdpqicdqZm19uKEbkb/FmS+U
mjyRutbrspSotEDvIXdyxf1WwrQ9R1TIbzLQrk0ujcyrh3Hg0rfnYPjWp5wYSdeoFSvwbA6lHSq0
j6a325W7b3Ib9fvs5vHm6uCxTCg08OWBUk6w5kuqoApHOvwOMJt08irkWTwx0Adl1GkjE9AMBSp7
TzrXbnxOGze6P+qQTmKH2Dx2XUcbaFr/j5WDGYuztN/LVJEmSy0hcYnjJjLaUVcvCwN6GxFl9GX3
M+lrcHlQtz0aLgCQnMJ5vVP6YmtIW4c9AeHER4JVzNrEOGpIQM10WNw5kcNvWLE3vKyhP02+TqI/
4WYBisafcu7xb4ozyrTvwF2AshBoEKby2ng9uThVYWUcAfj+EjckQNGUTHwKcqM1g0WuDQEg2MsS
TADPX4jscOgVvvM4p+XaIxm0yBSoC44sQaRRj+BqJXM9UgywA/yvZmBxddN7+FlO57hdc6veFmNC
5izTNaqoMBVBdrMPcHHtcX+qcXbBq85rZevYkUx1CsDXBSzFwM/D5RTiBZ6ONsbIOFSRugHYiBzM
KA2zB2qJbzN4hP8dv4itjPgcHVqEutgYumL8TPk3/iKP+juChb/2nasBa2/rAuZQm/m0DCJU1/OZ
NjgOZRwxiy/kmYWfak+bUJjCVzIfmCff1AlZUZrcK0jG9KcboL0q6hCs1SDP7/HyPent1UZoVA3h
K7UNze5fGwSp5XnkOFIPy1fLiXiIHg9PRBFLBuKDEloJGTSlEz7VrfhvgY79iS/evL+0ID5GN0lw
q7QpNqdd+xcMs3WgECiijOKzI0F7pIqyK9ZY9rS0Sa+1bi9cpNvLHEqgQXSwxy/vE8KMdaYbxwuI
cs1p72isM1AJZvLiIGGlX6ieU1ofn/QcObqfMp0PyPqLs+fBM8GiXgcsvh552nERwQk2JHvb7p3s
huxFVFguVbMJuhkR7eGK+uw7zZU4XeXrKTp27rIBUJGFpvcW3orKAnmK6GJmFreZ1s7EKDEV+bZD
jBbAI4RU7cMr+VpZVmGVfwCxTBxGie3ayisQy01ti7oqZyPr5PFudIXvzdhWBr8nqjYCD0uxxS6G
NuTdYvxiF5sYuAyR0bTXWx8eBN9hJJCO5n79LoWn93P8uBFzNVnsLoFWY5TQU//29DuvFHycpnAq
jndrv4M3lYUB4LIhDc0v8fIYmaFmdLwW0fIHUEJEeQoZCfNxkqYMin4EEotbkXqQ+sih/oXcgpuM
v4Hctnw5+qQMmegMcLNkx9hDm/HkG/autRbCtbCIMq6RKX2Dbnh1IBEPNon+FVZeMynI8OumSc4Q
hRzlZUAadPZPC1nn34KZYUa9VMozyeo73pafIfV5o2aLfq+aS4dPCbsbumELdNGStPmZk/lmj1ps
X8BtAm5SHx1W2BKcVW9MgBX7K9+mfxkkVvBXsOfwlguHJlHe+Xftrg2nBNmemtvLsYvYcVeNNzl6
PQQgXBRC8hRhj+0ScYovDinszO+BS5c1fSa5rQj9B/0BpxU6XnHoUY71lW3K8drdsWejsHsysBdu
lsUXZ3A1riRvvbPUEpHf1NrZLw5wSGiGJQ9yYU6D+5ufxf0k/mXOhL8iPMKCeuNM1I72DFuwUPuH
N5vIVKg40tsZu3DcTdRV+9Rgvi5nvqKmatPa5rUSWPZcQd0z1nOdoVA3vuPz9LP0gxzGmxfKL4CK
+aAEXYs50iMcXfpMWe6E25VRwCtEHF4uw8KQFS2wjEXs57kWey5tk7HQK+nKVnGaeDaiNCtIgdpq
bDtCT38hfz91g46DBDW4hmnqwlgVrCUojFd7yg6ku3bb74yC9b3sX2LHnMna2KV55ajpEhef0qUm
1xHdIQBc+nVwHWC7KWWwrudZnX+Zrrd8AmUxTZOu/pvikLeFlK2sslMmlI9Cjrd+yAnjWzdSuRgx
G3Ie0XtB0PqO/uGFihVHjTufcpZVcTzFDuRSNNFlHlfUtcqq//6YAmsmLAcx/LCFBSzy2biqgCuP
y+8jHKtPt4JkwanCPVcuP3mYAumexDBCKJ0PR5kzf+dZGFjS+iskmGW31Z3SAARoJRpkJHgRhNIG
BmavX9nTySUXZ3Mu0+nOIHxYp6uoreiLkMbzQAfmGzUJ6BQffzJsfI3wSQceTcQu1zvsKZSzWC81
+/95upVg27gLV1+toz9RMEh7sLW6O3JxtR2lXG5ZJxbr5Yg6y2QPrwYSang0r6FHdZUNaZnq2Su9
uLPqbh7wVrlQEcimk/JHMWGw56W+fv6O4UovyTnTbYLDKWQVz3ClGlH9yiOrkHqjZCVQCSpjhlLH
c6IeLxDSr8e/RT4RTF8UCeX0BjATgWrC2MWusMsUn6SQPyKBC2MbhZpRkCUC6YwaM0R5+CbfvG96
qrCJLALosYbrfxkMkB4Tk48R+JhxggPS6sS7w6CwdKkv1PRpRxgkFnibxorPT1LlmDXs+5ShO63x
b/cLzO4KqR0BKO3iQmb8h6nzPx1Z8xSAXRnRIsus6dJuTQUOYSGt9jlKRg4X1MN/k7nplcljCIXH
6hP2qmBmRWOlQy/74Jg16m8Ptgn7krP17nw2clHA2bEZ4+3LNyeOiTD2HFPT06Y88u5ey8bS7Lhu
QN65KOZwrWWyVGumAu2t2AEDIAu25/MIxGbl774UMaRNUatNOwES8Ru/1Xk3XxEcyEcVqKMXLtUN
IbcFFSBytIQp99Ca9lZbAMkAaCSnEhdyyDatf+rS/luJa5AKqpMsk238kKqPaFBnOwE8utotUbiR
uT1+YZyYBuFNFaZXLzibBBZDqDXQtMiV5a6V6Lq1qmZk+j1I7/mISn597R9B/BwvYCVFnmFxvaRX
OwLRZoM+s4kz0fmF4tLuFUuldbR6m46LtFY8AlK/Yfu48TVB7d+IeuQN6zk3XQaEQTLQkMCp/Fr5
FIuO4XBFlnFgWkmWoILCwOUOEJbxSzt8hVootw2JDbjpF8SxdpValkTX5sXpvk+FN5iSgKs09IfQ
6/rtbsS4mbukjjqGGtj+NFCaV2doKjPAN5VGx0fuIxn/zuyclMgsUa3NnViC/D+B3+ir4u7PZpXP
b4PqxAJ53kbW4PY3k6PpMuiv5W43itJjvmfx1Xd2g4RjGq9V0JbPZkXZrJIfEACyp7pa+5AUQPdY
V7awkCwTDZ45jgfC5gD78nt4QJ5ubmDzuBX4RIRdy1aMgUDNrnCLLlYBUuOAaAMJBK+OGSn0vAoK
AezBHS1496MlKmmOj/mFrnCpjwX3HUS2QM7UWQEP7ss++uJDspR7E5SX4sFSiOmnw+Gaao2NrkQx
wLCTTHsvxUKOzP3DOWdm42eTVBdcJtk6YCngQx72xRZPq2Piu3uf7J+qzYCEsMv7rjbYEdQMWXr6
ntcaughndJmbABqCQC7/YPkHPb5g5+LOAR3TRypN340yEKyw5giIrJTXFNjSRBg+nfZbgBFgcAGP
Sr4mks0ZBUDT3zzEfAK38Upt49EqVeSPwA2VbleObAqiessbgSllIyQSTQJxm+BkQlbXzictIDkI
0h7+dMSRQ7INkKp4nJYjn7jrdVHahlqlw0M09Nn2sknqiwn/wYlER4WtMYivsqrfag8f3ouXnmhK
/nsI1U1Q7WhvPBvOau0pBPlk6tEzuK66kY/C5pG4qiiqWbsyBZDNzDh0lADdj8H7pO5Y5loD+BJG
kzWhgCYfqrPFxYzX9MIA7ulRmKGq7/enUPvu5SZZFtyNgtckK+H6YqqXzbIGjm1JMu1dbKAQRnDd
G8rUG+ey11qMVRsbzMf6Dk3bFK7U2KwUt6Q74KT+IFyekMM3V9B2IpQJFCVrXVba7u4OgiNIqCDV
Qe8MnvVdq+RKyDgPVYuMXi+bdCnoMuD7PgNXMUx6YLhN7lajYr0cTWq9pUE+XU4+SJzCr5THQwid
23Kvpj9Ycm3zlB4w0PIgsXxVRkwyKp6FOuHu4MfI94XZifAHme8wq2uBkfe2yvdbMFgL6dfOlOsD
nLIwy8ThIdQc9t8PTxR/iASzOreUCqP2EBAtcIGpFkIeZ4Ptjak9DL8Uqme9vEWn5JlhqwBjZ/5B
geXp8JMiW9lzEs54fWHAosDtC6sanbTdnXZ79IbAE9C0czoAkD0ELhnaFa1vNFf81nLEXPQj6XOd
EUgxpIL5wgHNbvGQ/9cCgiIS/bLLFgyYpDoX5/4kJQ0yrAVek8cHCKOtHZvEIOT3ylES9LF26kW8
L3rcRxcB7V3oQmKEsBnvl+36PSl9+52G1r+FPdAbDQdzMVIcTtfDHTa0xYEMBjlDIZo8rzzBPo9J
kY+PBFHUagBcg8KuGFUHllmcGJ1R/J14TNpwTNzS5rYEXlsR8if+ifl7CgQus5TKMMh+DhJdFXXt
Y8C1WFr1XOMJq7OvhNIf3ykDxt94emprUCOcRqFXy80PhJjmW0ndS6ibBO8X/HATl1eve5/P37BR
0QV3Y6Cf2m3UX/367QWpKJodD4wcQQR/KjiDkmWIE8gapCoh6R1+VswKn8JzSIR68IxLFxroIRft
v29GeXj2XA1q+oHucnZyaTEGNJf07YIL7P20gOIr+BueTmiK3p7TsbwHCEdd1LdMh5lP0zC4MhI8
DIKLj/8RCZW6I4izx5CjKhMVM+qAjh0oQq8LnVBWzacO1j6ER7uqu9VMeGD3pT8+i576IfwoWkoN
PZOM5Z1aGHkQWcEU3dR10kpgNIhN+qsv2fNaZjI0P9SStNRN3SF64QxOukK3ljFS/0OQzCEC8aoj
NUC+vlObzT70+q6KX7Qoqi+dnn9Z2jTn45RbB+sgeRo1r0AuN3TTPZzcpsgI8FrSWrzx7wtLotv9
aQ5m/ULNKpnmMvhAQCaFem61oNtR5B008pZxQYXXeCeJCtQ5e1BgvjxnjXvRXGeJ6PM3E5OAL9Lt
0tnH8m7YdDxtMOLj7jcjZu6K9axmalqKhl8hzTiXki4qpeQjY3pBeSMWhDNGKRs3ZrXMWOAwmJUa
Sj/0+IXmkWbwLEdNxdoa1lPusdrd+aq2sHOkvzzj3BFnjRtvV8KATxaiiPtPPTW3EWjVW/8AApoK
pc1ZV+latNaheRSCiWKfdjZArH8W5x4Xqwpx7fqkFW8U0+brYi3HRcquVfrnSbpCCoTG2+wGrf6J
e/vw0ICOAjADhtlWCwbxzP3PaAvaROMZ8Q6Q61uTEsEOjI+9K+1s02FGA7i66kerHyW5wNPl8Ube
67qiLCTIghcDC2NfphftS5wvj2u9098HGo3lV4sUkKYQ+JC1Z56cBZMtEmqgYh/HtvZHQlj44+4h
h2NguKAGoXB3MYT3YQGk0V4YPHEaKVpqB3hNqGy1Y5RlnRf68VUoVU51WOElwjc4+JWCpRE2jGJW
vAUex29RfJDSplHSBc3Xs2RHBhuk9/0sxyga6hi8Y37CmjlHZi/s+t+vLn8hR56noNrSii+zXeM1
DVNeMkLuffLOIfPiTznmF3NIHDMRe9FArA6uCDcSpqHmPSwHZyvBFcojUdyP13/o9dafRbJfomCI
8biEskKdNa7g0UTIaR8ikbLErMVi0BZ4d4awVH8pK+Pa8U3tzhFMPWmxKqYDmoxx7fu7th6agrU8
rfPxv64LovgSoC8LLlvIdLpgb7Th5qvd+wQTt9GRFhZgX7n/Vto1LMMkw3L4R0ZMWCuG8+ABTxCd
Szm7b2yyYujm4lXVshAvB6o8KTwEv1o7l21X6oHzmGbSdE/tkEMgCllYF/zaUvgxuy6XgVrUuf1c
2lbVQG6DYg1CnBkytAUc9Qn8QXOKzNvT/FobOwEbNzxBAJTC+6mkaMz9Zm+NOK8HyfBBjAdPUpsp
j/CxAoQSsdUe93sqOjjIvpUHvnpN4GxSg8NRIIkwDFp2RO3o22lhoCEXFA/Fr1t1C5ZsGeg3fyfF
sbAYpFMBpVteV/AkTxobAsPyiHxCT83Bdg1v+bwWWxSJPmuWI08ayEW54aHzlqT26PxFDqQax8U4
cVcUs2djjri/i8Hpl8pKxKSRJLiZOjmUo0PBWXdmjyZ1Ss8RAc45iEOW2kOGUSqurna3O08E/OFT
wiJvs5SkXl+1UJvoUTe3avsB28cNanhjjhcj0WM6i5kdKdGOe+v0zQlrd+uQfRBo2qEioD4RMrHi
2NftHthKln5nxmeoKPprk4ILEBodopXpMxBST3OQeSNz3uyc+WZ8v0WsOpai3aCyaeldQjwDSmBp
0mUcgeONGfWk23mcbQXoc8kYu63h1sksLadWeD5R0iCwqIU2C6vbOUJ7i7Y1nmRRAv6S/NZX/uUO
QijrHKYd+L0aqXhia1azehx2d0OkP8KNoWEu1STtSYbo5Jk3X/M7sGZBEUqx3XBDhUhdlThWLRqP
9SCGy50xOJcfq3i9rOukAA7KnIEduHPTjfOB8yzs2DnH8MMft6UdkmFNjltC0g4bZ0vrhcS+nDNK
2SRkuFziYZU3jpLLYj3lVxXntC9C9g88B3cKeBaODQItXgl2c0wi4cNL7g5Itp28vj5KIv5y89eO
A5pbC8bLsEVCMWX82URC13KXSvdzGqW9bXMCcn6BmXbvLkHmX/NUrIAqMIFaPBlsVyUX4M/abn+m
XtT4bwgoJawDbVfzklWT4nFf9dadf4m67Q7wp+C6bZpSiwRfCjbbNu0zsA0+876PWEv9gGzn2hZ7
b2bRZZGb5T6p8ERHrr51zopQ7tQdVtsUixEy8K9BhLVhNhGvzLw64cmDC7yLFEI4zkD3Ty6L4n7n
mWLjv1QBvAakbi8ZJhrROonhQPjO47xkr+A6Zj37eh6kO9vo9neP06qYdTXayXQ+oPrCZ+YfDuuR
AMaJCr6KgDuqeTTOxc4HPPrRJbWFyFTwjQU68rI+cqEGg73PyrLD2scVkM6P6xgUhpwxUa6DX3Ct
9+UVHdP+phQQ5XL+ZPZ1yPUWEXpMtFanxUbWbfnxIZSye4UJVTiw7hE4sSJfngvg4ILf1vOOFX2f
3YeNNRS/4vmlQ/7nTjyUONs+cjmlFf1t41/dUDYesA+LZozwUb+acpb94BYxHTNAMTfHHxMo9VFD
dZjh0xpG62WClzj88/KbHVPTANig3Zh2/C/5WvHQuzX5dSw/LHA0EK+498rSiS78BQNH7Zet9JwD
3fUUTLu6yJK0Pb+Zxku2mhKpSj9jLAmqZJS2zj8tlYOXOKBGlo+plmPcFHVitPdvVf4SesszoKal
VV9r0VDur00fPc55Z9IVQn0/fdXyyoRSF8Df/EZUpHTDaDS5VOVCTbsK4ZzRtRWuaQTVkgOUjgyX
NFIkam2VU5GYSnzc//XvsDath3fBWWCy+RnMKlfVrcEtXs1zHf/GpwuMh7fAiF4nQGJlwulQaWgS
yGkt3qwNFCCPXUnpjjSp7wKOtr26Tzrb4Ctz+ul/SNk6KvO4LlJ9z0iVJ1VUzbPrSTOd9yg4JYwJ
zSykrlGE8+5H0J105iAFqn9QW63sIpsNFpNmBU/4jZ3BCAmkAmNkjHotLDFUgJhe5x2yCBSNAqbu
XewvQZ7T/e4MIhpuMIXWxy1bOk5bCvY9OwUz8XpywnZ5THzrJmWzk67clWA0Ben/NgQcLgD1E3hb
UklFtTQh1+VRiJXuSUHcPQDFAmQiKrmibujvdDJG79XoGiPaecEbuMNq3v+SA4SSIUyJqhSnsdw7
mLbkWt0c6FPB76oLujoe88QACCJdpcLwdaKlQBikqjJAEex8uXPlxQcmCieJMQ0+RuKdTS2wJAho
2D7+ihIHCTQ4b77veJJjV1uu7LaOZ8EjOVdyi22c0gfGdA8VP07ou4CFr6X1xzbyYV1T/jqCVO72
aZS22n7WonkVdh5IbRC24tQNWxU5NRlOHqHi3tdwvyJyGWHCUWcfdIV7jX7zTLcFQokzO/L9IzcP
xCAG/HQG2Dmg7NbDVphfkMo6tHZjfrSnTRTs+U5+vGRryIsero1THoPKTTqOQxKYtgbpK5jL4cOU
9R4xVx/Upu6yP9x9FuTD9JSOZKZE6ObmnoDztFq+h+HneWgi5cHxIwbLr5XpYBHCy/tNxTCgQ0yn
SApEx8UXCyHgebUsYE/3EYboekSXzoGjH1gkmRrbdTVMTFF1Wc1JW/JK26J1zVphkYT6mVQBtViD
Ax+iimz/BdPnBd2RxeVtFXOkJMPyFI2rKZ7RjC5MATBfc5SNuqm9xqyRJt+e0CUu9JvVQFkAwvnF
vNkVNEDsPtRQDmIl+r5o7PhsqL4PiUrTCQ1dRjIhCupY0LsezopkJwBh37zCAhhl3maKqKIZ+xGH
mB9N6Kd118YWLkHKlwhN0ynhQBOUAFwfH2lvGluX6hT30gfflkwjAIPq/ozUnwbxCP8ZMxnsQ9Gj
pKyl3BbPudfFl+0fQthZ40AuwIGou/8B3SeZMJ0K9Tt8XzDHtdw11bq7HNFpd2VuiNyyl885M/rV
jQLuIf1mrPWOU5zDKrhQ3gwyEFrC2CWlqHAFuIXyamcLi+hpEkKBPlrzDWj+mJSKHNVd8aKf1u21
YInatLCfcVw9ZCq1h2DHgKdlTGJJ8kH5lyFxjsxNcYvonT1lxfOX4f4v5xxH6cdsHKxAkxfM8TdB
kjPFvEsZDYhgCKbqH8DKAO4LHTn/Dl+0yjvkoqHc6TCK/a5liGUZtXFHkx07YIocllWHiVmEtHSE
ybD8vsloUhYHg2PVFYjQdwqf5Okij6OrYK+KwIyMrf3b209re+chjvg0dkihTpa8R+BZ6e4hn+75
pxB3yNezJAG1QVG5LQ5WDG09z6wYYqtvQemeFGXKu2CSlOn9zUOxS+bVolxJzLd/Ge0mGqcWHK6s
sLrZzgg/lOsmgbnLOIKAmPSegknAW+/1yVfjEosZUhRbbgqCs7X1KVjB8d7fpcRkNkUjpv+Is3h1
0i6xc+nuy42fzKYGJM1TwHfwZadnf59wBJuo6XdICr2H7LhAJXbPhKAQb5eytwP8ccnpYmFwMCFK
xEYxRB6K8xzMgQ6TaiDKsRqp/hEYTPErMINYUwQrEHqy/nkd1MzxGk2vOsVOUBYZHYk+t56XctZy
sEJ3M9iT3twf2lAQLO8utQN4JRqjmm0K//hvYT9n0NcWTCaqyUmQDaT6gJodtQKz8OtmGbrhzyN/
0+HOLz8xmrY23CRllSX5AQLD4MjLwzC4gz/4SacPmMqqnz9FiP7aEi9S+Y1H12PNHfdIRhJXvKC8
hE7ps70nv9PWJJUBVnWcTvMx9BJMXyh4U1trwGeOFkH/G/cl15FKqP9XSIKMtNgIpMUiqFLzER7X
8l1YQ8/UvaMxFzfcFqOVQZGgYX1bhGNHcaOOwG+oyBgMd+l0RUsuNKCWavMQYV7EheATJJ+wHlCK
C+x5HMP16mvjWg05ilURU1UXqm85+m41airiWQEVNJjT7sQscMpDPkDmMQKtlW83WvIYApRU96jX
7Fd+FJoR348sTrF1jwulEaxspmBq5JlyJhYGrCBdVkyE+5hG1UL9N5lc6wFstvnfIG/wnHdrnL7h
IEPDJpGp3/DHH0pPmlyCvIxFJX46qQLdT4u1fSn0MfGuUK1YEq5/uYRxWy5c0Y8iY0LzJUj84Xkl
IT4Wp+t5+kOR8VSgfO6/Z+ZklGK8CLZrh/kfDgTnajTOnIQBYkP1YQO8X/lyy7y51+o4bb7cMh/1
lvhyPlZrruJ20FXEtOug+TLLF0mZxspaxr1EaImCXpfHC1L8+Bzy7aOJWUvckWMB4LirTQUf/6fR
IIAh3uSMwX7tl5eIy46Dc9Ukz2G3NbMzRKaPMbKPGK7XABIhpOr7ZvkSQG+N8NFJ9lUbE6KT7mRl
d1UQB4aXK+5g+xUHkL1z3raEtLfzY/5H138GnQZF/cj/rX8H50hoxYZ3+KfX7/vLC76C8FRi3cN4
kgISyHKtqyhnSZgcJKF4YBo1kLtPIp/uVPBeTlC6sNkn5vKf/hJhnrjj8/QME814wyiv7dtC1Xu8
EqHQJ0C/mzjCpdcfPN7RCE5YD2qVMf3Pk0W/46vaiq1pB22lFgyTrfBffcQxc5Y8jXcp52HVOXlv
ynDcSQMOauAvGd/VR+HXt2qjQJLV4xjLiGmFwXxGFg0t7vY5LsZhBdvsMJHNgn2vaA+orb8mq3RX
M88CtXWlx46MrZhai4I+VAdaRqWiqVpDBEyr0+n7QMqPDRtoGMOhQ42NIKDZBKNqvet7rnpqZ2iu
ZvvoKBUOh0JoEbB0u7mybOG0UTjNID1Jf1oAsHcsla2y/WhX6hRfTi5VzT0rY9dRkTtLUa9ai+zH
pAR4nyvFwJhMDR2XnUwHIIkrkonpxqdjfVjEn5NXXaRxS9VRYPyJJCWWtCEpYuLs4OvIpjYwUInb
2mEsVbuVR0EQUjXqoKXFO28SLQuunTPxSYdAYH9PPBDKfQaXWOh+WBUZsllWzoj3Lgj6pPGalesb
DRc6MmKrEz6794bl/seAaAuPR4QyjfL6hY+2u+Cjz8MCTSyFzSjTZsCMZDI78HcOcUpItL4EsHpw
Ilh/qWxaBMSM6wYb0EvMsL97A8njUVIHFH92VyDU+4PACV0bQpuCTBDwps2xGdnj/wb5fZNH1CPF
swipFRWPnmSeQI1fX1ntQ1sBxbsVlupHhgYsV8P/T1JmIINoYha2huWTC9hhB/UBBWU/ZrUhve6f
46wYv5mAs/6D+nnCIFWejc+KmEdwTtshe7JKF69oGsh07f9t/jTGFSl1pbOg9tu6koSeR5HXT3Tb
KTx1OY/tkMvpfjafzn5IhCsdMSwJ/VCwIl7qX18snSUsVWAFj64UlK6NRsqGNU5+uMm0H7yLbmGI
nyhCgOhytD9bywe5lsmdPrXgbCtSKn+4ezzcGl6D4FZt7gPztLJvgCSrCoS+z62cglzQ62pH5/XE
33mhT74xcWLbTudyiFGuhbyK3VyxNQbLCSZucaU+NmbosHoqc3Ab18LsjSNpYdij3e8nwmuRjv9I
Jea3z4Lu2FakjgdGeEcnvIyKZVH8Jp6biRDiaIVF69hy4WW02Ke/At4Fbh+j5CEa5N1A/AvpbDhk
wQWwZLHkvzT5gxRxSB7kaVYKlidY2XbmXeGT3ZT3aRtGUVlx9hWJUF9tP7RTGgEfv5MDN55WoiIx
cKANMZOzjyZln1oI+KJhqMIQ1sYxQ0pCtM3zu8Q0e6pqmxSFpcnKyUrzR3sTw5M0GiDJ5d9vwra7
rJAssNrP/mq1ZEIlW2T8InGJcYse4UjTbCpG9h63C3yab8WVqNem7+vw2bwY4D15kXVemgaoP4Ra
RrnrF5spar64wInzZqbaOpmouPAFU+swVq4fGOP1CyKgBfmFeMdxU3rNXu60WCjUamKkR3hh+zJF
I92wAXpe2JeD0bOrnN4UXr7N+0YKD6fgoeoU6FNSaD4Z84a+FRs46xLy+06Ur+ZwdoLIhW9gRrRX
b4V0+xWAzNNTXtv0VbW/CPJ0T4dhgPdWo8wvnL3UG/6IbJOA/kCphbkazoBTcx9KbPcSMokaqAhd
Ba5beErtomnVIWKT8X7T01/h7yzuiUDQyLYINS0b52xGCPRXmzWpBpYMeJLEk4HWEBXs4jO3EGOb
4zasJAmpAFboitPPjyf6N6baTECUpS10CNqA6n0Mwg8xG7/WioUbqO4nbkjSZnjudACgVgn1MsPX
1012Psq8BYfHk9vnQ4zf+K8sHLnf2mE7+DtQ21chSdlUH55bNZAB3KpoMjjohvV2N7mWBBN/+0+b
woW/IphLcwNBIATOUZKkfxlmOIdTWx+BTE+iuiM/BYiGJLHagMkPKMCQRpRUxbbn694lnHueMWLj
QgvgX3zxCyg9MO/hHitdzcXww8NpRHg3jZxjtU3vi5rSBxE7zIfa9mbS8wzXc2tKEocz89qDOdNN
ZovILd7lTcVZz8+sCIjCZwJVsriINYBepolpkhAgkNazYF3L9JRFF+zjLNqTd/ueRzLnSwnr3RfQ
0xcwGuerkxZfdsSTw1sIjwABtukkVSg9cbCKGjQwdy50eWNop16X8Wwf10mVVpObAPltChQf6qi9
ImZxAvGlDb+oQ7WHPfdN1boUkS8DsK8n66N9geF/ErENxWD364N2aMxjPJGOER6H8qCjxSwQlbsR
JaMC34dHgNdvwUYlOnhBjUnQZYdy/q67NyYPbB7HTQWR9tYNaxxE2DZlwVTLBZJKlP4LRUizbXA6
6qjHgLAlO8fRcvFNZtwZ9I6UDqiwocTVds62ynR40Np9tgExQt/dmoiskj75DB3ALGGBI7I25SvR
MJmX11B3xya8t3eVhhHP2WuAMwJlXfJByK/F2UkAJR5F+WZgP87+k+TrPcsK+/uaxjNisryy2Orf
Exzitn2CQPiNXXVYlNh4UF34aLP5IzTekLAmDJ1jnUHm3FquTTYj+Dq63nI0tma03/EdzhbHjLSj
Shk7AIAQsCqKysil8PDudWDiq9t5MvYd2lXI8EAQ05g63J44zoq9ogahRR8MEj/rR9fw1YDasAH1
JytiPk7W006pTZKr6cuNKJV4WooRpaQGD0rxqzpucH4oJGZkJ5XLIscrh5g1oITrY81GvfeSJ8pL
kwjGuJRwGOX6kicAO9RKy9cpdJlyLGjgbUsoZDkIO3hO/arso6ElBD70nxMxHmJj2Zwuq8CSCKPt
RqGLpY5zr1D+1AiciERogV2CZbThZBwNxXuwpJcL1THulMXL8muWFIZf16dLctrsOba9jprpqFNz
GoeAbN2Ia61D3UGXtjwnndgdYm5dDsfPpiGGRv87nehqPWr36Kgu8ueFUypCbWWReW7botp3IC+f
xj7T2zIHotMsLnmRRpCSBYi56ILN7iCWsObwofbJ0rxcmTWktoTLhLgEErTIxAIiTVHyJZmMtSSG
ApmRnm9ipATXqEH7NdPxO8Gm4OjVKjv4gPltX8gu4AekIPZIpw4yawK9yqlmvbNEhOmh2pgtWrlI
pes8pKISoaKyxm9aR5OMOm+slvNKLjJOQQDK5qPq41TOZFIrNEgY5R3DNj0BoiIXwJnjdCoxW9xV
8KDlSv3own/jCiPndZTtE+LIMJNsaapFq+A7FVQFgpsl3oLBIAGky8fDCOcdocgtde8wxBbqvBnf
pPlxNnoGZcVQtjM+69DnY+2OBDTnTa7VzZuDn3eLt62HbGuO7iGmg7HVqRNxJU6ehflDk8bwJWyJ
Au8AoQaWzC9x1e6gREANKBqYhp6Xwm51y6XhmP1D+o0aeqoxTO5qpOwSgf/rD7CGY98oNEUvrFhQ
8TQTPwHLU/Kd1b+wWnD68V036StzOjwW4ViatU5BLbTHJotpgH9m1hGhJCU6cDpiJcXrfCoLcv5s
c/ZbMVNNuxQyidaCPRfeiJbz+ZcX9kCr69M/gDjGE4VvhKM46yt9mmGGylo0tX1LZRaFp30fNnQp
bh6BzL5kXJZSsSfreOSFFsYcwiP2sJsnAQZHeHPtb7U3WwWZ4Z7fUy8c4cDMPsXCzB5P3qnUjEUm
E5y7qeWVCHZo6fUogjCO06HXQ3AeR7HuT9DHItwjmqQMWg32DqMpVuou4YwkmHPkY5FcD7uKmo9A
zrB324cO3btggEMw4VBDyjuxWATXi9EKk7x0B0At5QY6skabIl+toGypUImt7olcMweQWkX2eEpK
nWOx0LRAkJPo/J7yIeCiIKkJOxaeDjYzua350DdwYb8yAEBcXolz8QTXeQhCj6naxV8tTIWORP0M
g0sR0B0hVGmZNBG0sfg694ecH9LQEu9Xgotr7w55yUioKgNaf8fZklIZXxoLtmjcZt1FCBkanies
j+KcCORUkB0PwjkkF/AnMn0sxA4ANYw/ebUDsOb39gEXbKLjdoXifvbOBdRC4ct7HoN/D+IN7tRC
9IggyX9PUJ8Gg4MJbyK6rU4FaHh8TzfN7rLwislofV+YV7YnrazFw3u4LM0aCbkvweyCo68lkRJ+
xA/PNsx4e75m30UJqugX09EDhrYrgXWdIywojVrylGgzg6+c3MoDA4NwFFt1R9qYujf7a3/E3uW7
BTrGqqR0pYMBeKSv05FJ7Jy0f+sQq+XhG3qcjbMcEQQNnj0tC++Vphlke8U98ITBJ02CaZ+Hh+lV
64euuLv6AnK+bEzV5Q8g/AkZrr2N3edNzJAvW/TThWeIYfy4g5tO9F6DXQa4GtNvOlHc0/vrWwGm
g8UCNv/PvacTnkiAFO6Fpw5VPcTGFKa09DUKLgLAIJtixmLGjIrl32AFiD9yRydAXEn255rF2hfB
/Abkg46AOi0ZPItW/AHE+mbMJqP5pIWo3IXOo+HCh5yxZnJQT+lEH8rTJscztkPg8o8pdWypNAPk
xwaUm3ZbI826FqLYKwlC3CO1hWdZ7iS13CLTsvJuHaIvJXb7HY7ABpHeKit7bkshlq5HY38jWWZ8
MRSAhYVBBe0bHyQ4SXuNtq321IqdjcCsfrYyZWVgYDpnXZrU7gfpDp+O9ykaVBGsTZgj7qppUhVg
5PAE0KSBOw8omVn+Ll7/ldu5Sx5QaO29h3ze6mQ35SZ0tUOEvcFUXaaWpXc9IqobdwuRTpljsla+
lgP6CShi24EO0+e2lMx+O7t/tsVrXjSQ1oNM1fWb4OcFTUBdnDqdgX0xwq0UFHTRVH3i9X0TmpZa
d5xackx2dvA22l0Fjwqm63Z7CgnUmjerF1xjdsd7nlANut03aweWSV6tNwI82Byfjcs3on7iEVqU
J9SLEBXz6NB37wuSa0P40uNwPp6biNJBJNhlELFHBpmj9G9dRgmPpDcyliYv3S/yipGhuAynDK1f
OqEb0HMZrAwvSJe0FCk5Jug27h8NFJ3UDX3Ox9aTTj59b7JJ1kMSlTCVNqwjwKwho9havwluYoC6
GQFzHXYYckDd0cxPkPHUMG2S7DbWUnt1P6Hp1hNdfCBRJOwVwvbWgcWnsPElKc/hHckFoeqFYyb6
TwXKKlaHD2CkkbN7t/xxlUyRMttgJxBPfWQacObS6HwcTqHzx+9fQjKpQMUPDu+s3bUYlCdpj63t
iJbbHHA40IMrI4HGHXmr2/7Tt/qfTdkWWquurmQCounNtVY03AsuHu/7Yajk3rPUugwvHC3f0XzL
KumVD/hR/Uk/yTMq6rq+j0mKw7NV8EWl7raVGYul/IqXzy74VOEkOQrM7u7QY0PI/2kIMglsh+Tj
HHqFOAlNWWJHz/8ldbAe/jk9UD9rR2Dj7pK2FnOdy5a6OX0CqrLSctMUESnfaAdEvucFVYfRQrfK
S7/caC0o3pKTsrH3tS51LCS38Akg4ulTO6pSzxz520ohFS0zSYAazt67K5OXY+DUronkiLKAQYb/
DAYRghEhJDp9d1PpPxqWHOUHLm+iBcpAxZzkWjWAyxg8CDBr44qOF2z0Dy1UBYvZtN8l/3Bi+8RD
jHe4hAWvFtrH3l6wFK9fyL0EcUdiXvStyOOpRJfY7Md0dRtV0UhZSoG4xB/PUWxT2ccMnSlWom8f
2vOQJou7+gGieVM/kH+S1xW4RqJBHh6X5Vr+SmDXU9mq0ZK5Ezq9mqVkyL2yezo1DoOOI1MJyACq
rBoBUC1OKuxYMRFV4KSxJOES8cSna5HyXCfLTh9a/qL0FJYDqSINkbhKp/00EWZMWXnjo+HwEAed
80onPxc2i3AjJOAguiqznv5Np5K9EZ4ARXDJEIPx/CTN44hAeZzaCtr7RrPLkmz8YKkpmEcUI9jN
IYIw17G7BM32N/wc5C03Vw/lFLK8/JcjmbL2Pwi0EtA2TW/oxtr3tUyS3OzyyjCzYo50Eu5sX3El
eJ5MCT0JrRWijy+7vbI8QBIQwkf8Hw6mgK97JHzFJrTHYCIJSrslUexjUhMqMux9W/LHbOl9p6RL
P5Q3jtg+lgj7qDo6LRBl5C/neANwLGgQZHkCEMMKjsn9eF5ZYx0JAITo59nf9FzDtNeJwNykgc0T
7GIS+GMI3/MDOA6cCnOmL6GxmeAnSDNX2bdHtfpJpT0YvTq0akPF7Vk57S810JIvGIEd4IYpzVe7
RJoD8PwZ6+FxqNQRWRRn5ITWc897vftR7m91zPWKWnyrZLlLhvk+vlHWfnJgzio7msDwva9CiJIg
U0SzYlcTdU1HWsYpDhH6OrPH0gTM2JGJO8n4M4lGbNlWsN5Yz7SoehfDvD+RiVyFshvucDhDrXHa
DMU2w88+H12wh64awfF3KFE8DQLGrhkKeieGLf8Vy8/ZG/FczPBckfNbNd9CB+VeEK5ozsgF6VOp
JJ8fzYf/k5NetML0VqSsv9iold5JOokzzps45TTyCQeTbjBrbuigb8V5zsEJXDnA32xGKqgyxy/a
57ySTVq0vKGKna6bULV/WGZwxKq5g65otko7XphgVVqqYlj0QJAIbV90lQeOnJLxmd1khtHQCh4J
TeVGtTpcYfBjP/wfGetKXFtp/u0eaTZmVBiKpGBQYJ4ByCSBxp8tpvAkIebqvYwnbTt9cPPISETK
iN6p5OoWCowFOjVZ+tUMF7DUvzcp29j6lkNkV9AYqW5skRSvlrOwV2L4QJkhTrfQgU3OO+iEomf0
UnZgtQIs1kGmottqXC62oI20XX5oFYt1Leng1zovL+njDoFZlYin0Y6ybtA93c/xtee6v6TGZ2dn
7nHpvVRRXWi6i7kNXaEceKlxqFr7SDgw340K5bZ0nT5+H5Grc+Mweq7tBOi9a65nPnnSsWLGUigQ
vdmkIsyxwZHRubq7xEgTb6qQHuuQp1ay2rugzYhSy14Cr4FRPJWKR10jljIODpXfSakD5SpyzG+z
Q+25acHvpNtIGnX85TAgHcWTaijR6zPcuhe+BCtOzaiR0mMYU82ZuiPDl2VD51wy99PibBal8e2M
YB3qFk0KcReZ2NPVOUA579tkOImjs5wwneHbjTWA6tCL7mi4NVJcAEmNpN8EwEPcnRef+a7P22zm
MUIENCVCdOPEfOAq+v5umR/RhO/l2NPatMvEJTbzPIGWwYBqOFEoMlz3GmvAdrTc3jK53x8e4YWe
rgrCxyCMt3AAW17lMVob0RLesPJGQIa8pNqEM6ZQAOQUbDxF/l+TF4ut7fYtba+xXdwAQgbg22Vi
t7M37y4kZY1aCFXmD/mGsWr73IUos9VmTnX8QollPMpV3HQ3TznX7+JJHrydt5nx15ZSPn8qVNkN
pEtWP4lbPFQKoug1xghlEqav4suH1VL9arSOdQda6upbM340yVb1UbQPBR35JMX7otCMB440Dsg8
hQaDIqjjElBZyIGHXfzm59YXMeO55faFjsfCFR6UPbih3o9klOeNYBAQKnmscDZiSA4zenfissTP
Wkj2ozfP0M4byXRhEQfYd5FQVVvx8RbuzFaWg0s+aVlm79MzsBnppiwSfVYvCF2j1AuSFpi94be9
hEveU5XDGzqQ2FKnjgnFbIcsj3mYvbbJbhI82zKjevmAUFFWDIHXbhpGDQKLX/O+RcfUG8F1X7CX
QLYX9HhHn5G3tP2QLmb45/E6hx09lvXCKqMy9ZaLJzYO8y399OMjDFMY1el2Gjp+fIMGfghc70iS
IsdTs3sOo54wC+1KqfR/g0EUMg+XjBiZP97vZAqx/IQ19z7OcA7gdYKWNqMiwTSPwbAUI4EqDV9l
+QBRKe+t0Yzw0kiIF2yPGjqBwYqnvtS5IZncVz5aY9Np4pk+ooZkplaW3I19grdwGfX1qyBfyvzf
HF4J6YGZDQyJUosuqj8LPRer06iU+CkdsFhWUm7g9stItlJ4CyV24fV8z87EMiU+7cdIZReVnCd5
ihDyr3+1yoN84mxGYwIlgIZqkY6I0gNSbh5N9rdHEpYa3hjXKQzytQRUyf3h5qY3EWISGxvVhDKN
CN9ThorRNF/+aPu52sCEmt2O+9qIoMhCDiTYISms4izg2zN/UznpOvGylXsD61I0BVYGsAGvKI1j
oSDAXncWQDqg/g6czReWKv1JDf7NGgJ5HuW+HrM/OGhco9EvDSde+rG/vOpExDJ5zGIFjSFj4ygl
L9uydOeIY9qciN3fbhB/W3QBcosSWrj4AvKcJAYx8/vGs45ASjueWYQVtST1V8ntPd7zbcTkQ2Y+
SOVkhs6hfuIcPUIY1kCalzY3BB2+HbzWuYFcWENPBXLalR2bHjTrWeQFerzwUircI9LkZNuYvYlz
TQ0JrO/im/E0nOOu1WTsFnE+31ul8seALiB+aAsTnEziuEssbZ0k7Og6RgyQict1w+yXmpFoKV5d
8Ftnwb/zSME52Wej76IBjretcGuCpaSPV0P8Vs6z/Q9N3rk2D7R0SaZmuLxU2hODL41hGwVjWvnV
9RssOgSLrjl9dMtMprbSLq4xH5PuW+C8EUN9zxHRKNtm4oiKhbbzLB4LfPVh7rkTAEKoU51uZDtb
gcLx1LugbOcsm/bolJAtijT9fm0IYJ2SxA0H0RNojM205WpHJv+RI2q/yNXVGjkxfhdGoPd4o7Fh
fpG7UjyRSsEnh5ayzwL9lpSQRXoKXm8khK4KDflNT9cGsNYIkL8wesRg9fNwErDb/Hpw9hWWx4rw
wmIP1cB3vGM5dO15DuzlwTUN3b16+4A+4sx1VoIQfvh9Unpx9XlZQ9TZRlCCqN7Xsc2NIFHrrpzI
CjIyQC1vPBeMC5PclOcriVr2QuwrJA0XlcqzCqcaDpC2Tct1dn3n6cQPP+oe69k6E4L26owLWCg9
5TkWTVHAKJUt4lHwVtBds1qvZVbFuxTwg5rdeztPn1xdkrht0wCDn+wignBPX+puxw37epjPjPD4
uN49LCTeUZmjcy/FRWd3Aina9QbDNPgZrYMia6IsVrVCCz/t6vg+tQvzVqH9G3YG4COa3bcTDzmG
Z+OLecJXrIONEaNYur3DhnI/DcNi5iieGuDkqPfunavg4HJuOatG7q2KSuc0VqhadpoxU/PlhwL/
AikPzEuhnqVcnlikxtMAUvaQGS8O5B/nIiIGX0it7xEWgChxMyYULDcvD0Mv57ucYusXaznoB5UO
yDtd7WlQRvlgoB+Af1KwEPqu6hXGvOLwbA9NrgwXPd51qbXsVKwzOW/aa3Zh25/IdlANTPRuLLbV
VO7cQzsJD12EVyfG/rPkBe/n4cDTBxkSGhF3BOkI/ckKt3RPIC+woPNxv7QXXAdykqV/Upm1Dfqz
rTDrzuAi//uNCjSaczzelKPHwxtmzT6ANjHaN266VzJTv329Os24uMJUmDS/xkPwWa76mFflKK+S
5HkmN7nR0wVhPhQ/1BOfV6Q7qpQ6kFQCsAGIV2upBog/MZDOJ+5JH68U03UDewyMLlcPheFuxQBo
BuCXlJWYOTZp3mI040FnzmrfvwsrjJ8UUdR8UvdduVzRAhUSqSCH4fR5E22/G1aKVmQQmEWDtP9d
/V3WjDXSYQOxJU0popiiV4mAFdu298YFLrvKXdqXrP+66RNVo4grRx3ohvB4HcC74UtX0rmQS1SR
MjKu7CuDbB/hUmL2aYB7rLwPpTH/WA9Tb6YtMrjwckTX9eOaq/A/JQo32j30VRe90jRn+OP40/CA
JeBCd7oHvtNp9CRfILmCdVklCRw60NR6Fn6XZ3djCbbIYLE8/FxQGzXbCiWdpY8mtMVqn2oMlscY
74eaKEHOSPmEnnywMAPPSobV2b6xBZFk4fUoQQ9XlMJSrF1YMzWqb3QA13kgg/g97qYZhYJm0BDy
RBA1PfypoC2SSTotTvHs5+VEW67Rvl/72KIvQMn/nv72Aaf5gU5tUzj8A1pBP5wYNUZWTlrsF17f
v2Toi0FAy7qnQeemiyjdUQdzhb4O47dUUj2HCll6a91b7cL4KWmHtof/Lymbqy5hWcFiIyEyX8bz
MZWUgNEeZczuAj2+HOgellYmDbVQQrrpbV2uyUbdbQNUGUf43hJrLo+MsxA9rqyk2fNH/Lyaa2uG
2ZV+ODIAsPKM/yGRWfdq22u6PE6mIxecEKAHjSh50p9oPaO7Du9ibtbI0jJeCzz8RDc6g7L2x2ch
AqKqrO1CmMvLWLwpWpsJBuWDWcDbU36I6cQx4BBb6kx/y2VMdKRnetT3InLZigtuouEyGCVxDFvP
zRdfZsAVpDNps9ceyk0mNWpU7HPTLPebL19WCZ3TwZ4ccDG4ENkTi6JB4G0B9/LaSFrXl07+urjB
uKYItMxkjfZVS+2+/pHiDnwuXpnxBcDRE/O7P1DYqN5Q3R0Up6Lx26kMlpfsJK1nzmG646tCQzYX
iehobhIrEk+ytHBoCpcQf4/XWKq6aBRmWQ8/5INqQUnPtoPe9XivMfwFkzoTtqHMZGgRrbtfwIg+
aDYznLAdbwTN0utIQM8K2mL5hLwKNTqbx32Tg82lmuK5L/vyC+T8zT+2Xf4jYg7KtAQkoxUs0muN
W8wfR1s7KrV9KXu5k1qp3uypWg4kU39VQ3jGaNNUp0kOfQR8/COFhfKNJAJEZb8Gljm2w9XuFmuR
8Zdd1S4JNf9DQruRWXx4BgrzOY6jcr32mQK2UMQ3bXuTJ4Mb/abuSCPIujXKJUsFNfhUXPGlgF2Q
EZ8kcOrGAP92WAm9LTbBSBXlYZHH08grKKZtGtZh2onbYeH1wksYdWQGl+VfkEZ4XPdYEQMNpnbZ
PWfuIXd1KHx2PNUM43UfZ8j+p+OJ3FehQurzf9jXo4p8i+YsI75jGzF1YsNlOOqPLfBBpg6Rq3Oc
AoV2My6ZYomBBFUog35Ff6dccQba361RkD4We6Jx58Uo55175e10BkMzoPFvLlwfhPmBioo4ErCq
lmIjv2uv7ja1fAtqn2m05egO+2gXf6SxFeO9P7zYqas1j/Ydrg7ue+lUkC2pTmpB9nuOElEuvjd/
a8GETpN5k3KAxfIpbCuhrsRhDr2HrxSkxgOG7bsIzsrZbb298LIFOCrIj0tHiC0m0xHqx8USXTXV
zeA7T+KcJYc7+slDk5Y9d2o9orUh3gBxBwfeqWyNrxsjo1UWmdJspcdqOT/b3eElyELz8R64UEC8
ePIZHe9EvMWMkn9Yi4ERatNfmcYiTJ+cZHzxhjYK5iUKr3UsybMkDe60hBPsE8zT4+AOb5CHwRqM
DL90432BIJMM7K2QvxkUj/SN7esxquXd+xulHzOyrXf4Oa3OLKgLu2Mp4NOttUJ6wGOnPv2BWCL7
ZlvcJO+VT9rVC6XDka099JYqvNh2tZO07/jvXpdHeTJiPgLHHg5WH5YuO1y8Iub9sKCCqwiQHXxt
ROsG+v59+71WG6BWE03OJkWZelxneieZaLPBlohk/zJ7cYRayKH9N2kE8PMmgH+hs97h1CXR80KS
IF5CwAQP6dOZWbrQf0+aHg7O0sJ5SVsvH1eWhob/U/8elKe80p3hYFw05JulsI3Fbpb8R6gY3vBz
hjhGDk/W+UnGety6/dkhr/z+f5mKxLigQ+3gF5nnvC/6Pjrd1WpJDHWnr1rNo/i50O0KccB/smd9
RgUVpXMCh+BCCA4ej7sB00Zj9va9mirWF12yKLpsNi7suj1gwqTX/c2qRMDnlYf9Wt8OSBbNaufZ
iEvnMMLzvF0xvtVH8SYM6VDonMs2aX+HmrAW/VXPikoOagS7xzUyLrXmGjpU9irNKwzDv8+Onq9e
3GgHWmNkj2nGXZ7RmmGH9b2TtwXITOSAkSBR+Qflegno+o3zT6RkqXHk+qX0s48fNVrmQG/anSYT
GuPNP+DMddZ4oyqwRy0d3RhRKBRB/HIOun7i2vCps2Pr4Q3nSdxQBV9rUGI/SJq6UdMKAyRRyl2+
lNL4f7q2WUZLLP04FCYmVRaCBmqCUnEfcJZSxlwIYHzMa7eR75SL+hn1654D42kZ4DAE7J5Efgmj
YO7QlArxmUTXaCgafQ303rL7JUC/unzsFAj+n4qqgDqZh9QbJzjVU9OcZTDKftQ8pjWbQamHiR78
lcsMKFYKCkLydzHnJ3XtIg+kq4EtdtJcWZUOLpxR+QKtr+sz8Q1aN6uXmWUw6d4JGtMwH2s1P7WJ
xWh+PRoscSPwZqdWgilQ5jJNoT8QdfUf/Z64AfLW75xANG1U/n2nu59+vf7kK4xYfnlQytPHR3sT
DfjqAjMICqVBxOWDjp2A8RYrWa7+47GOANN/ZcqRtc/Tj5e6ymj/jefZQaAc7DCjjgx4lHkJrOLE
JzC5lBn2wZR+U67VW3EeTDknSISTW2ojkR+gYkeHmzLkPdufbcx8qII/4yUBexsCMcklXfJXjR/b
KdfLG2xIeERVC93Xlc5S9XkQNuNHf8mSakMWebIKPAc5kDInXWBrTErnN7KKUHQsE3n24wzXjOP4
TuZPrASoivzZALVsEbvxvVyo9kAOot2JxQDp2Yt8kw/jOS/e6165L4cWOCx6E5zxaWCVWb1lKTy9
fCCK8upqbfulNqVLHTzFfA2DNFezYgBBx0OIb3/BIs3Hii+QBPCud5J63TXvUmQd2etJpxW6hWP5
P8QhQckdDqzeGYu3n4NOuOQ7StN7Ohx5a9OxoMLY8kfcXqb4PIYeU4VX7ZfHgFa8OVFWBmVptl8A
DVf1NkwEqNDfNlzEYplaOBvgoEJNsaM21HLSMAK2UavIghsIaikMMk+6PIzvZzYslcW8WkXz3UOy
6dhGxXhFEhzzQX/QdfVnPnVeHUCTsTyNB1X/f89sKBfDDb8rvOEeokt9bPkGdARlOAdXX3rHSEAG
C9Fdgn/m4TCXv8M0mjeIM22DB+J+30WBQDz9+2s2ENmQUCQGswZbTnTlEUlu9qSMB2ux0xvukG8D
orZg5qLGIyh2sjkKQgy2dSwjzHwfA3vElGhQfWU/ORKaspvVKaWdGKb6lJTLE6YYcDJkGDK4H2m5
7/vPTCaggMCJNLuEW7IwkxuhjXJaoA0nVUPsiX11vVVV0QhNfZ2AII3tk0pOC24CbzLhhQQSJP+C
28Z1vEvgzupgKY1AYvB+0OwWfWty+WcZksAPQpLCHFD/EPwUruRu6eJMx5l4LCzKRXQ/RkalglHI
Qye5TfxrlvRNVbkNFnzo4qZZLzpJ6q1t1cbDZUOWTcgYbxZR0YftZgt/kzYvDmQ4dWsxLgYleyxg
VdUuTd9zMbgzJ2FshIMCdt5WqEIssLoEwoQemeJAgXKq587D6graa9bt2ou5F1t1TpKEjv1/lEvw
Rj37dKJwAzoiKvGkpGbf3DBjy0Mu8IJviMPUcO064R/gb1dH0PEiNFQNXY4pAqo08ewCu9/dqd9Q
pVVY9WnMYlMh+DnKld4hM9XxT9uJcLw8fc05Me5dan1AmlUNFpT12md+IV+E2ns+bx6vAdhSAlIU
bkI5e5kAVBf+PCrSSQhIbn+8Q0oxAFDKMULf3E7fiZR570cFnDPkBw4vtXAnuFvhevLC3RDsZ5Wl
l5yNETvyA1oTTVN4ItQZKjWMKLlSm8ESPLiWgVhKY2JJpbLmvLcCK6UZFhzLkycqN+cN/LszTAWd
cUaZ16NH11PbOcCbOBG+v/Pl6ijsC+LrS9IAIjDmhXzesXSyrmiK/dvg9aJ5Jof9N8fDxef7OSGU
de2dYvh3s9unk7DZxtiznrYNBOvoXfqrro/5OtYZen4y8jaRkbHk0B/M84kAaT80F9HoPG9hIAw3
JF7ys6ko1pbyEN8vYrp9LlU1MWHL3d7ijZN1ahg0zh1PPFckv1BQ1pxdApN651+mkDk1qcUhM+9S
NNfuIOkCshxUx2KPaUveqSJYHO9i7V4qWmUbC6UgSiPm5EnH7sJZsAhV0zblbCbfS69fVqj8AK2P
kbUxDVt9yx/+NTXb5J++kRcUlqXRCB3eyqRUDsCN372y4rzz1u7SCoISiBbsU1yNkf1ekNegRKZQ
XRuka3jafI7n+busoABaGLbj6Glrhl+7vxLt9fO2D4Kw7eeBSzsmczPgD276POq2YSgnypWwk0z2
/lydHsG1CW8PPhKcghLtucmGcE7M1JmgfptpEggyByVubFqpgEPMth59Ody9k4a6WLq7xlr6ZgGs
58POoAWyCrMzJXq8DBqWbnkuiIuNM4UOH3YxaAsCk8X3fJCrqlxL7Pl0hMqSEQPgkMpOzNRbxeY4
1MUZAC0AjLG5T7CQbYsoRnApNH6xIoPJjznywqu05bu4tfdvd1UujfH528AU6r7j6KqR3A6+HGGr
1hGX1+VA+QLO4zUdtBRoHk/qFZJ+ydo0DL8bgATwzCKqXzJkgAnwKkTA1PsnwjSaQuxqrZqFAksk
MY49c5Ub2kSA+bl+EX0tNvkeqyGH7spsHr0eHuHq1TQ6IWaQy0jyMC+7RrIgmwFnsH0PbR41JYNP
3fom0JdLuWPH5HHQFl3672we8DFBzVc5LzI4giMrSck0Fg3/3N5P32syOnvGFsxV7ct4V2UHtwyE
hzsBWWfitDTzAqDDy9wbkCV+5ZjJshQ2n1CY+GC7SlF5IWeGEOF4T8GoYIcslZT6DDSPVkCwuQpL
Zgnslil/CptVxwAmzrZQzqRL+yMw+mqGnUA356jMyrsDMVS7/yXEIxBbO+J24W4reLNXODSzjmvj
W+BAVCGCYz138JO6qHf9vACg38ceBwlFzhxQB32xL3pXBEFdziu3fj/dGEUGsKJF7zWOmSARXfKy
16Lq84Gs9Ybt8pBxVuPSaH7SYqaCrVTrqOV23T78V4dMV3s+JqzmhVhE6z92FkfF662GptbDTvdv
HrdEye0LqqbCHPa2Ft950VNofjmjaqjRCTuvTbU4v6qeivxICyugPW+ssIFKQWxoHKkW/TVPbXUD
IzYhLgVYA0Tt3zumDjOcugYhKRrWDfMUc89WDUfhjC1t6KwPeJk2M56aaJTAqI2EA+WgKdCZGlOu
Zaaq9mHomYOU0svv00iOTY6Zbx4KBvTDt/y2DU5ARwVbg3f8iw6PdE06TM9FwDZ6jx7MMjWQIShi
1xwRFiWo6yVp8DjFmcTW8UsvJF1qFNHxCkdkgkMhr1daiaLiyF7ENQVNbxa/Y25c/12rOh7LSzXK
uH4ALGF+medFQhveFTFXMPfd06+uUgicHIfWUCZTomSwF4FyFmFH2a+C1pgtBxmXXZosC+EUkJJL
K5rTk2XEnP5alhmaX3tcixC7NtSibePdm5j2Fx/buotcKgoQBcy2BKBaDpKMrXqSBd2hX8w7AgFs
JwgrgdwPxgulM4j/RVJhjGwZitXAMMOtAX0Iq0+oszbSI7hfEY8ezUYAiS7SwP5KhZY5OJzl63kZ
U7oyVz+tRHs7yO4KUlnjI77aC+pU5AKte2oSb6juEA7XHrAadHtLZA/nw/TPwt44sed0uDtKpKud
sd6w9Y0LSHKsdx52pE7ALu1UUswpCXReixyqi7TDJFC6eOv3uN4CkZM9cTOFDsczMvMNHuQG9vfH
Wqnt/M9EsIQiQbaF//5GKG/U+iC8azfJq0RljMfRoKA3oF3p0+TSgIhlvTknBGmvG/Drh+TzNNe9
wTrMNvVoPXMD3tLqz3Rw/iNxvN60mU1pvNr6Rr7vazLUMZPsfjVyRDzF5u2C/QsQhHtoojkTgSDn
PhT8uOaSDXlvsVbMEEQPo4bH2q7/p/6kn5VP0wLLA5OijRpXRlikIwv0gSVo1nvH938bmp7H/6ec
4yTPLfXxyhWpwaPxuogRM6DvNhRbn1QC/BSJRdBXeIAgfJyOj+mfG9s0HjODmkfHOzCejZuhbL2/
PnPsbMalSp9dwaW716K9CMuAqIJ6jHOvkGqlmdUxF0w2Rp7V0rt4JeeRi/m/ATl6HFLLtFdixj0i
9aQXzMC/AW7+B8u/b1BOl+5bqJl2saLzo1zHCiRnNVFVr4wf/vknvKIgi2RvRadCOFA7LTz8p5o9
r+Wj4b6/kgC6N+mk3w8+D0oBJGwpdJ9jsWKGYLKeb/9dx+ViZjkKJAyF2ism5n75TOhiWvv9tqvx
VBOfrnJ4CTX4smURbJhC5P7yQqp0W1wlITqsgrjwhmPlKOXa2sf9LswSNKDskkX0R4AfWVs0yCYp
sjUB+W0xhU9y6PXRJhwFiXIIkoYGkwYY1hf6AzIL9C0nXc9sPMycIqRBhNvHkkov1Z50I9jRsjWU
13AiJm20A9BShHKCN+AIzXqFS+O5UZYdUs4qabGivx20Y3rNnNlTzLtYQvTCqDEzuTRd6iDEgwxA
yVJl93d2He30qVpYqXlrbievzJ4Xg76LcyxNHJlG8E6QT9r7OfenKIe5zoI2qz6U0vrO9gO5aZ7f
OFAJvhHUgcSfn3crhjlWtCFpbW4HfnMOtQJb/iH8DQ9IrhX9v5uQVgewFtAWksUhYxuGUXTe4cpm
DW3NeuoL21LTf/xav2zjYpApDFT4dmgj+zEVPZ/NgyaSvZlEZLd/4xiLI0RbbZjjS7sURh5L+z7d
da2IRmuWhfK/oRqAyRQDD73hG+HBPnzKOL5b3fsMAasn5KiZiv5gk3ZPV462S0uv9zDdK6blyRx2
yF3vqASaJUAkycN5cjy4vuau0KcLqRq0JIIz7b6QYoZ2bMQiT9pgVe56HLRdIDTOQG5QpNu8XQ0U
OWWkDGwpXVORG5lLZQrpXfqZZ+zNf0WWDnfH+y+cUtbhk+N1KjGC34FoK+LpDbAob9fBGP1hiXjB
IMnN2/uRCQ7seIT4/KZy9JwYC3nBTzqyy0nlswoPRxs3wGIDJWcy1ObiqgMxoeFAaj/ACddrveH5
ViF2vIIQIXKsfaixibBJ6DC42upxAm15zstgfQMkANPHEeELdUGZr5bn3unswn6RB4OgprGW9Kk5
RgfgXsBGDpdMCdYkWw2nJf17iNs6g/4R/RgUpREL3JoWps/1OBuXYGg3toDrLprL5ugJhk0E3GWE
F8GtaVsFzv4kAGs+X2HFl85ouB5DuzxK8b7qC6a9yRsHF8UOPINrCPCRF1/iwdzb3t/a+cvw0ltn
cnd8t4igjZZ73ZOsJbapeMUPExDO/UpsBA7PeLyicZs0eQye60Ow8WBY4itx7XQBZhVLwldue9FK
UQGFAHPxuDpeSHkTqVpZyS0mmQa+E2KoX26NCdY640oj+eYAReIVp2trTU1HlKJvsdecTUAYXlqu
yVw7b6TryCgFvR6DHqBhnrqVH9DQlz+NecF5QBP1xKJSDiat2pONEE+UC3onf/T+7RYFQieUBlJ7
Bl4WfN/g/NvYdJsdoIw+rBz+5foBEBwb3jpv3YqJKqiz/Sef0INDIOZ8B1xtD9F2NJa0W6BFC5cj
aOg7xTfswpzypVyVSXZowxcg+ojj5Z1ysF03HIye01yJ5yyUnio3whj4x5PGUrA782A4nwmUyEE0
+ghhX74GreaLB6C7FWQ4/LIfjglPyVS4Hvzs0IPIPzFBv+mdJQp6fs+vv0fN+KygqoexHrjTXP+m
PotL4HHvBdDMgCVgtE9gL5vpS+RCc42qx/855GF7AlSvRtZgMFUQSqwUoQo7ShD9zYHcgPOgYwO4
ZP6HP/fe0UA8Uu0+mARYFgL+l/D4Tv5beyo8B12hS99vyOPdSbH/bq6Wea9YUOPDgfFBi7jtNK+/
u9HjALe82ubNCA0L2IH3QxzVWL8S9b1O8Ey065z7XofPGNlEe1Pxq4ibERRQjNtmZUq3wWs5GfUj
fxACPbsz3iPXJOO5uHpJzhuPdmq1BeL2/idFNDCfKMTe8UL7mnj280dMOYoFN/UakXL1PwXq4xgY
Qp0SOV//Ywvg6ONzTgpFfg9ApNSnw4aVG5gy8viawQZuzAV4QMyzRioJG445xnxxCtyjJ6PGwXfq
wtYoPRWZ8V2E3POIB3aj4c4mPQauHKMRUIj6GhvyP2fSUCDsEZbFT221J0GvY3WddddXZpnw8tqv
wX8rC5dPAx3UV8g2OMgLnzYMzEAqNyCycdsM2ZOEPBfSBu/8hpwQZvWcRzSE6ef4KbSFlQXughdt
Sp+e5t7n6TDwUilYOsOyyaz4j3EG5onfjSIjVqevbbMvEz/hamD4nHMU/wFAcM/eL5rJbAQfZZk6
65dBMOazXm5ODfn40nvMeAjTrHbeQkyXRRreEeJ5Uy1hfBYqO5WsEy8R/DZ2aOxLx91hPkKlga6g
/Ct2X5Kn0cio0EyRapMGqhiVBkE8tVBBUYimejjLsppxwvo5ksUzp4IpgzBdqpRi5vebaoVagltv
wsuBjEV2Q+YaufheAZ1TT8P9MB9TAbjan8Z9J5QYIg72oo+f8xvLvbklfVaLaSlW6bcjZ7/z+kUp
U5HAOdhxM0ekWALEX2icl0zv5EOmIW486TW9TpXxYW5OnAOC495c6Ocg8wTknNT0a0wQhwtSQqcj
/mIWTnvx17Rx3NKT/8e0aBqj3et6UYbY/GQLNJ90zRw70e0GZVlT38HeWQNmJedUxecPPwu4Xls6
qE3yXS0pEEH9jG4hK2inF1/ERnlgq5yR6rmeBhs803DQMBs0F/vi5XzhnC4+WfkJ4Px3RqKPdQAI
gPyBUR/Q/aRIiAJkOtO3shIl9N8psgO0fs6WQklBUTV87t2qq7cA6UpbBI1hu6uZvdSD6Li4u33u
eraO/L44yYyTHk2fHDR0doBWwJwhEaW2ZfBD/672bjPbakdDsu5scN0GgbqEC5FdhZ43Fou2H7yS
NNC0kEJUN+dvaTA65yIgrMXdlqWP85gFgkZyBxdDdZp5JIwHpHTlqFfW1267INATufEE8vW3doC5
8xGyrhCYAK/6HfKtpiCUPS5jnD1YtCGFGkD3rf2P4s9Bk4cVwe5OJqydFPl1ktzAWpMvJSpZmDWm
F3THzTZKbgB24Pm2dvxWBRkp9/7GxLG/CN2E40evHxWLiciWhkUYYg6ptZPH1dxKLs7Aa5DQc4HG
NfTVdbrcUzCk0m68ylL6jSB8ReX1uEUJy1eBRZI1acYM8qr3ehWeaCOp7BjBT6y6J1kRGTa58nWo
FGbphDtCSTpHXItY9VYQ3+a/VHxwadUpzwJri+jWCrQo0dZ2Gmh10pKBm+UKbMt99d87j8cv0KKE
5/02uI8Mm3S9dutFtN4zdKfJPswuLcDmf1dyZxjo5YoDRYecex4AQoNBPJboskkKfG93+cd5L5JV
sjEACxkMLg+YMl+DMjsP4gshwDnBPKQnUyuiOMgndAnnV56zHBag8UdZwM4PofF7/WapjYYgARCU
YEg2Bsc2mtjmvt2/1GVRTZ2aDiLOpvBN7hVUhU3i3sit+rxZubfzj+fZAj7lK4pvdDz3zwUy3jrW
sQALpFLsZC0jxPw+KkHqLLaVGaVtGOsXaKlW4AQaMtchAkPzK3gUBgoMzkldzWF79OWrwCzepC3y
dEWPT1onjVbTXiTKTYKFjrOiTYR5EAQ8iPP1XwQi1q++h3C5lq74rNCd5/NXQsF19leaJ+G9EdV3
va247EfzHP3V2VpG7Ieqr02sezemTj30av3/whwDDIKWbJmmDEepNERo8+7go+x4gChIycLiFmYF
WKVmvLy6tPbwFDUuoJNZCu+7igue0EBunkL8RNwRp0BKc5/QXhMwNz8P5oIkudPKK/YLlYq+lGvI
HhgqjIfEdTcdd5Ddinfsq9lHypJvL8enKmqY+xjfcXIc4qRNcIMJP10O2h1WbTEatbboD1F5vOjm
vA9mcMuTqUnq850jyWafxPIawTKhaX7NxpTnHxltOmCqyu4xgND4LzPYgDbRN/NN5Pwk50rpWUCo
kdL90jnRKykpAli6/7cGlzWF0FG0nlw+ftjxaVFKZwMshozZlz53siC5YaAWNHvxXPXk4vrIp8fE
Zj1eRptB76UY22GTg0u8cXri+7fHdihgaKNoT1f493YkggBO8Y2gTfveNEwDgssrfpjTQvXsXOE1
1A2cZ4r8cTRricJrs5zKWpd5sR5prN5I3fnz0Mg0LHE7r/iDK+Mqf47CjZzIxYbgp9D8i/uGlsR3
LgHWk/fT2EHVs2SorRX8FlyoTnUW+MOyIhYCZXG3Cbl2IUZfs+A/UsBiPJqbZzyHn12Bc76pXTwB
KU9ivqrCzOIEVQzN9DRICeNwCJM5j5mGevv3ZVv3vwtNb6iiw5A6Old8eUTaMgcFlp2TaO8PL4N3
3MRHl6AlOEF0ZdfNKflJ921GEjP5L8RQjjC9frwjTIA65hqFXOorm8ldZRbv8u2EaHY6E9q09G8T
ifeDWmURTr9wANtCpfI5L4GHsmg0Gh3WGG6mhm0BcUw58tPYESx8kdYU4sPYQV+5PWte/wdoJKXW
JOLrJ6forPv17kQu03UlltV2N73Zx9EqXQTEy4iaY3jqOzIBpxNNeD19Fpm5TahPgX0j8QWqgge7
/r4pj07uB+GoewjmYtyC18drycVkLMTnnMBNB7nGXssC8U5gL8VJHRcKjm/qzBwC4HzkI2//5NgD
Fg2rjnbdNZ9tO5AY0HrLcUqp+mX8INrbMkP4ZE5C/H3mYueFvbfMMpub8e7SUp+0oIU8N8UazD3z
SVX5UMJihO0uOmbZ+wWz7Nrl4sixRFOmfInR4fD7Uo3UuP0CtR/POivlZ5C25hOavzDiI0i5HCdm
eZVp4QJXL5p07AGJRO8surz+if7DhHdXvWGVbI6o+VszMaTKCY2leBPBwczCTeGUkvsAEphYJgck
5EalFsOjXdPmANcErpQMLd/ibp/693NSgrMwOKjFfz1ChT/kxiLAXlrDJ5VluZyAGtoWQhbg6UXL
R8CRgMxm8XVxoKqLU67dsmDpA3G0qyl4018wHZRcPRQd4zAMyoMNEOd+8RyPMAOyipwJKeW+zp8Y
Ct1+uITN9eHjPO1hAf1C8od+NZ0JaSiuVOBeAklLWGoLg+HMPQyMX2hm6NutOZS5RYQP9va72hJw
ZvSkWHHJ3Cp5U8Mo+gRFM4Lr72b4qtuny55zBd/eCIA5LrKts+q9hLBQn+LbG7/G8tvAuZuQ1fsr
5acESx22M0u5Crr46QkjuPhzaFcUTm3NL82sb4nX2avkRfclPa0kdbQleTDMhxsXWmxw6Fvrfoid
7kBZPlya5utqqigaxi9rq+G1xW0kHI6Q4REbM8zfdjA2Ftm1RVCNxb7sghn/3z1FgynSYeTwMYMq
sdpV7icpBtZlkkoi2vp+akm7sCkWXpCJrJTpx1tc8MPLzqlSNfLvEAwhfBKRglfO5v3nAlmhPyzg
78c+m7UFa3Uh0pTu5CcGDcRbNp4+SZywaUnL78iZGGsYRNZ5gDBsghWqUe7qTtcg/2R7o6ZfR+sy
n3oblYrp5n4EmvLau+X8CFnIG8zDLdWISRRgcWTXlHFYyPnLseNHX1a1rmrBhflo6n7dH/acloSy
sAkgf7hQmO7z1ljWg77bhDi48aPXR9D9ht3L+38dwVYmjNjIosnJ4ahMnf1UJbvPFi4SOnqXt/La
bWMNqiXWy8oQ2fM+pBSp8vqElyRtnQ99jExDBjmQg4uW3cqbfGcU39pRNZvN17Dc15Y/XxiU+4XI
/WgdiE5znrJMRrInpRXlHnbPxP+89ywklT7K+PNgRxQH3IZuMCWg/GxbX6zTJWMW3Wp5wwPyG0Cg
gbFCBdr6x+IKDxXojFsS95O3+rSFKQL9mFKxXFdiSXeRooDZy+FbV58C1y/D9hcn4H4f0QmMdlrE
FcpvicNlsaJInDeWDPUT9LoyVy6QsYGjNBfoxoj8nkcuBkNv2DV66BnE/oqEHooPKxCYjv8S2Kf5
4X7N22LSpcC4skTEVU0VhmBZxOvdN9dbjNVO0BxZclo/vgKU4GpsWwcD5hIEH5bxW+DMWbgO6W1o
lgANAE3CBxgWaFiJYGcqTjr6gihwyXQP0jLqp/fZn2yNrX4asHLSbR54+xNuzDeJINCsAVR+Aa79
ezdJjjMYXZO0d3OEHmMVHfDr/J29ZxB0oiqnC2GMH0wQYdd18wJMIsCm/oflihaNT7abLr1ZxATy
HFN88xpil3pL7MbqYgHCG+1IpCe/wTjF0m/D1vwIURsOSUu+k44sdfRsXDu9K9J5SdidQll2hXKL
mbx0DwUORIWRTeIBOkUGwYc6zG9YCKmVUMclY4vvdtlHuaWOaES/cvwoO6rDI3BU6AnEHeaGlpzl
B7+fozGCZOaZRDyGd9tz4A1r71ezh8sbD5BBnGOGxXfLMyzuuk6KWpnabAdIJZgUcrr9Hili2mJm
iAm3OkH+EqTm0+a3yBY0nHF/7XafImM/ieBEnZ4rbolbiMiRaNqcc6c/SrV7lfYpo5ScGAWxsuz7
PoMSHZ+52Hw4HXUfvZmtW2YHGhiJYFD8rhi4fQLTWZHgb3qAtEmI48DXRgqHjI87IcY4WufP2DTH
xcMmTS/m+kQV/oar8uvn65EbfHgEnTYOfj2DZIv3U1fmqBD3J3ABK85wCptCH0yH1ml62IDFEGhg
wIPrLpUnoJx69HqwGEsphD05BHihSGIucb5W1AqRAByLpce2DeN1e0b++1tivvr1p8+UyVDOIBLc
XmkQmLUHG3pTyVNBRaSrxC6qr2GiYdwCyKMvBgYBr68H6g1/zsaCuFdelJP22QX2O9P9mrs1SQ/9
R5R4IXXtDuXyLXxCtxfegmb2CC7y1rYQ/qSs9fmJJ/mf6S40BV/OFkxUrk46uio1fURAsIXVBMVX
JU0KCDnfhdrdAjmUpRHoXefgUBmKXDSiYKeF1gcuPjMVDURR7bZlFVZKKQWUTnIQugR5MQnScrxo
JjQRSV341M2wcXsPo3d34pKOTl95hM0TfSXstNi3932XRpMWjRh6uNehVXVanOL49+b7V7Lvnwxg
hchLE6tj9hf4+HvOifnSjg5lkLm4525y/xRkZRkYnLOgwtircW/M3hrdvBC8ZAj3lcy+hHAJMErl
eCyCK2SkrIcnG/1kXLAIILL5zqapVAv1NLblVsVE1GSpdwKSZWxvPVJwT9CuHOxl9IsWULLEBPuI
76wcQQy9tKlcCIwtCiZjTRjw6LgRzZpVEJPxqEPYGPgeX2rY2YOb/ZcDwzpmEVbQdGmNtEBrIB0S
eDrxOE8to+XCy9XD9/jdxMFZX0kz4AOCJJb75QQwgNEi0m5orWee6Enq/pjoaagHcNNkegFReufK
7oq5cNXrumiG2GR6dgs5ot6AkKCfYIrgkQ9pXeXYpuqQm6JSDvGAXzNNFDTxIcR6svBLVbyoKpWL
7P/IgrAElJ92jI51ZiZp4iF3FhfM2zKEEX5LHWET/gUg8qc1tnp1bYRDW2sARHR51sBP/G2teq3/
uZimWZ5a7KSXjPxgLY+KD2BHGJdfhcoV2X93MTZPnSaJBRtQWxrCJ8fv8hOr4oUTjt30TzPZY61P
pPEgZOrK4yjVNX+qsukh0HXQ1dQYZ1dTQo9QRdfbQrrJP/Kbaqge2Mwp6T60R6Xmb+Jo5C7q+oLR
cPYrk30i09Ore5WcjE3FLadsrPWl4+ElaH4Iud7bIclYatmvelOSKd+nE6QLeasYC+M25LA1OB7v
4zCIxuxpHokdHxduAP7zBL9pYCUZfh0nE+3C9k0hY2P0EhcP9B5OlBkA8U4I6AdlGUTaF0UFXT2z
cNzK2unv3byNF4X1WuLs7Bl8ljO9B8WA7HDA5er3Ls1mxtaEeeBUlg8l1xybQPi8uRZbDgxA2aRQ
ncdnONhnKjYxLELflT6PyBG1wWyhe6lH2lTEnJBPb8Od17UcLJRlqsFuVqCO0liW//mDPrP8l4LH
f73VbzybLoD0qMdrNrfODJgJygmKTZczWPDT/CLGYbNrp9emYWbCSJ7O3ykWfdfJZMVu3pHh1NvL
Zc3dhf/1BXqXE3c+GdZZmD0akYY0tuUoYqME/O4upW5WOlIGQHXD70mpFNrAHAirc6gBDsq7mQBd
ZLUaigM0WCWQ8hR6D8GOPvy9AiXNFexvh+ADMgdtGnfsLK/zZABAjcjvmisbhH8b6Doy7ntMZyiI
dpZK9BNpFWW0h7DKg3Z8tJp1LEgnvt6tOi5G3Mcz4Ip/9MVMKqNPlTOpwF3U14nXhUJ5aoCMjogE
tKqEKtu5rYIAWs+uOjCLiP9jIWoyfMPNPBnniG7+fqv/A1mA3W1PzILSojlUXeJj7M6nTwu0TR5F
KUw6RtSTx78RdgQYx2S4ZyIz89zZ+Tx0CNvxY3wwi6HlXGVga17AwmVWfJqSpKOvLQLJ/cjOKq3s
fjgSL+9ZTx3+Z3z0q4ONd5dUrMjM4lW8H8Snf7AlwkntrT10p5iylj+A/lif0y6/jcMmpzv9FHMX
zz6KtpB5B39SjXEy2v3LGIjykfWl/v6lIidOZTy/OJEfmYT6bmoB+3LvvXDwfto8jc6LX/0ErFam
NAo6rTdjZuDB1MHQue9BBOPEf2CfR59r//wGbpj9w6y7W9Fqns3N/lG50gyk6l4uZaNYYzZ5o2sL
mtLNy7TGx7ZwfeYSvn4S2T+AOPl2BILIot/E3ACp7kumaMpD+9YUXCI/Amv/2GzC2VRn1DliK2Ah
3OcmCrT+DF1Zp+XRg9VA6ncPK6twC1QBSp5Jwog6B1eMtA+hndWFYIV6WkTfsRtTOjP4hKd/PLgt
TJl9f+urK5dHbSojEVDRURlqK7fW1z0/7oyk4NLpeWc0v5L4TfCzFmSogVSYjPtDtqeMvLBVCE75
ouw60Nq/c8+j7OSibTKceCmlgydVCOXcCPGvfA/6rFGioLwUVdejpdaj+jxSHeFvE10VKBDTMZCf
W8Ixa63RbosmJ1Ne1eMoItlSQHVm9GTL4jywwG5KAngbF6PABbTMHuS0+YLKFvHTODesPxduQ2g0
X5MlwDO+jswvgE7ZiiXHA3G8je2oCQmhBtOqWcA4CboEHvb/gCfOaUSw8sGy2JBrpBKIiXVbxUmr
hKWykCLOIEvM4Zyl2RYBBakvShfxJhvxK59JzVCHl324z8wTyzN2KdI5QrMXOXbXcgXVKE3ujj2c
4HNeIK/1bW4d7P9wagNY3SJwaCtBud8+NOF/3PFTyLJGDywAEpwD5HL/vls7UWmCT1HUc+Pw2WrM
ElwhrooZdH48/8uCV5C5pSQLkTT51e9dpRgLKthPpjdSwRl8e6ZMkTE/kgsquqouQRlQ81hkJ8uy
OPq8PGu9mmRi9PN8+jSlW+DH07gqCb9aH3LwnyGjzdsGbpgnr2g2O0Ox0tIabo0aPGsoLEVuOt7m
+x6wzG4TeBZpfa3ett2KrkOhKC4MdGC9iK9hkeRuyAYSaRu5HSDJYjdmLZXo748KZ8AH5w4boCiB
yNiDcCeo+UXxQYxHl2SfVduZ5MgvegCUVfLok4Xox63p1O+kiF1vg+tZFJU9OE15A9nRpsTh9K3D
/t4gzmu2pqSO30YebZYlqhz9ja7O5Fnl8IBdO6GW0Xh7OB3iytxKVYRIbwLri/KZHHhgCxKZmG5K
i1TdONRQ8Cm3x+baykUOEXYRT4yuwZcy8Vis56P67Z1ghHzLT670NArEFJxxvsVZeoA+cxOxDEZh
hlHEkQvDbjEKyUFMuCXZ1ziGGhXOyQKVLpRbc6E9EIZkhfDzPInAIIQeBV1BUHt1p384zbMm+Zmu
dUgE4MWUA0HmvRZq4msWYGgERqHTHhmMMEfZOQhM4Cy9CjURA5KbBlmyTfLXJiGESggzlrs4S+pW
aLgdUEYaTATLg21IPk8haWQMPAJfJDgfsQ6ASBD3gVO6hPqvUc6Pr26tzOEn56pTHJoYGhJxwJBg
b52dNvO21kMuIOzncqm02/X3jA6Bc3+/agZiDR+EVOh6yw9VBE1Hetsz7JdGbwf7Q2jE1qfXpPHO
92xfAlNHx0FswWqBsdANSEu8UvCoEfTqcXo63F/7WpJsd2wQ6qLl4hKXhDxW4joQSosyIkMZqYdS
aUSOSvCx/2kraA3So0VsxKaAHlSTEXXtK9Be5ybnEBk1quXi2pv/wgprqqrBuQJQkY1GZJJwmX2E
TLghIIY6sgWQ47flFgzYckhaY7DfFnRXxxOydkbdXmhQxRYnyolnguo4ZN7Kosp4J8lsy/zKb5pF
DQUxAxLwnBdfllReF7A38oHUYVriAafHp407KccYC030wS3fVZA19ZIwCRulbX4j1ts13Thf457P
GIEUgqAJIrxRO64LZ4VIru+smV9REo/pvBJwmvuOCHCip+Jew+1HUzZHkWtE13iYTuOAjKTABFzR
/L7TKL3qwGfVr1CBaCqqnj55f/NNmhnYCA1g05/9Sag65uZxxDgZVxbAtx2/JBsaRE71g8q8h99e
AJlEcCUh394OhmcfiZ4X660MHyAppx3y7YVxzTZ/XgjxRFDFAIUXKQV+Age7CHSsNYAJOXfB35F9
vD3L2M8bvJ7EAfhiL6kUaeabEST5NZxypXaY035ZxuRVI2StU7Y3QTrcu+Q+gfo2u04vBfygjCc8
cU3uTd1T5rOYgvPdyeR3GqB8e79h2FM3ikcNdA2Fund9N6Hz4d5ZYntUkkZjo7uK3BEz6CzkOzvD
2abDb7fPxqEzy3RIQiOIy21ovdLJy/3ennWVSwIwuLU5B7aSwGWS8pP66wUzpLmq42A1+kNwy/0K
O0cfgdwDZ8/0Cs3ItexqpgFnSu61YQ/kCFMd72RZlMpjeqh2QZpZB5DPyA4bXJX9mI43YlUNQc8H
i0KM8SxgMUA+lNcnEiCJi5h6dXKpCP30q640zZ+KMTe1xn41HrG2tlvDe1H+IPd4VWdYYOw7eRre
Uzn4UehjbJ+gI6h02k/SanOUurK/4qJLXmaShGdCKILfX0yI994z2X9eaiKmUvYIpRstVl8YiOZt
bfQxJCVoxmEJ8TaAO7OvO2oqqIyhZo04db4olJ/gNmqlyidMNbGrotI1Rl9HKYD2hoIyrhBHc/U0
QRpIM0PBbo/V7Vy6tvRIHS1PTtTZcjkojKBoNhi2RqdoutzbObCueLwWXjgNmiyllnGcvgk2Lfu2
4mzT9Gg4vzaqzk2QUG5sIU99ZpsvQAsM4sQt9uE/o2UdBlDViwVlBr+p6SHT61e2ZS8nNMwBQjf3
qBFNuqT/3h5aWWUrhkw5qUp3I9Gsrd0YXLDqZlAx8Je3g+2W3nSoCrz2oJMuqrTXEPggccf/c4HO
XCZp2WkRz31+poyaZ2K4ues2iFhkYFX7LSKTEtVXWUQvi565NduOvbJw8dxMNMusa3KK5sMr7cME
A3Pza7dGp/z0lDPZqruKywK8rCWkTA69sC5CP3RnJAWu4c+5E6M7w9+OgbZolu/Vg3+9Lo8zvSGQ
ekuHmPLvfpGchJL9oMcWhI+vrpnto9LQzVcIsTH5YIiGHNtDkj8wGvEyBci0En5H5wMrRuPP/7Md
u5szkcyuMqiTFLa+LRjIJPz0PcWOvepAB0ma3h+rJNn9dngI1wtxXr4Y7sILk0wqIcPVvIzbRJUE
hg4OLwuCM0bKSOW3np+4J/6RVCL5vcozVpWKISnQTy/HN5P8bQQwLizAxXhY6OSUYMdaiI0yMk64
AM71wNcKoQJ/KvrmwdZwkof4Wd8P3cm++7OO3pfpC5kV1aUgjwxJb0Rg4XSm1qmQg0adL9k/YiWy
OVh++7EozYluT7lg2QbFARyVcoX23320e7szLZXU9yd5oiLFvKlCqMPT+OIirLYk0zR6heE+ZXYE
SxqY25bY8gHqkwC3xTUbKHZGH1bpDb0RrLUL3UsYr0JGkodt/StiMY97YogB8k7xFb0ppm++H3vX
bAt0kVRep5zRD0VSO7EAz7iinSE6i2mFXQ/gWKGv1jIg+X5kIL8VME9419BHY5RN77pl4Uu7EV+o
cbzd7jnm6Hlc3TpYDG6MR2zMeKrerPicbxgsy03ZDZKDdToxVQwHZmXmeAyNDOM2H4CUc3AN4yKV
8tuWgouQ+ARQ4Ed8preWIryFiSBrz5y/enDy107Rbgyh+ghZKzrdJyGobJH13KA6Ub1WEuCAoG3b
+fjoxcJiqD1I0igg4XwtlbwxEXltDU8gzcbuDInVZE7fcrdx3v+2mpq+cWL2vrAnZL1hwgVdFO8w
2oP5SKZdC7+95fngNMTcoA39dHXGpO39DcZTAxQGEiX86H3L+aX6gKBZSa5ljsZhSvp5r/8lu2LI
ESqBIve309+qMxLWNkHIdWQ2Wzj4un/Xl9IA/KOlt0y0RcDQyWtZAB9QmKNBmFrZ1bNhukz03Ztc
GTRmSwNPfL6AYST0KykXVTEuOsUuF5hhq6d/Wr/ayA7xDYddBU70USjlMCOjdN9+NsU/mp1o7XAw
6ePjc2VnRgKqXoq8LmfvKcSaFnlP8pzzPZ3oAj1KhPvYrE55Hl0l3r5VKpRSnAJyc8HYnZr+vh+V
lDpqRbjWAx60w6Cl1RHhU0PagiDObAorkmzvdgZxRjZdaVIhaetP1druj7dW/zvpySQdCwsVcU8B
tJq2donkZiuisi8o8/5wH3XMawl0arYGSy/+RvayXMjIojE11YMnQb6jtVh8x/vS49yqrl5bPlBQ
TIS94NIidESmi9Xg/iYEehon2k06BOQM+VGJ6BUoXenh1pFieHGzC17BsCJHZSLyjd7vPRf5HfAl
PdWqXHr8tCvbxooHhaT3ggwZ0qRLq1mWxivi4koNs4SsS4jLWLIFWiKKtsW37VT8Tk3mMy54LGdx
FdiXsfNEVL4gT03iU7jo9TTXy/SSO1N+boPeZG12BffslFtD8oLON3QLWm2gR3nbo+SzKIXNDEeE
z558kFx5beKsSogf53xU+jMZBrPfR8BN2M9F4deG88xLepNOXnrcsOwzJlUlOBa/x3/RbmfbM0qG
vJ6D4A6/YmXvYr25+rZyKDbMquPTafbgPyZ+6Q2tDKsDF56GSSVUrwdk3Hia1I/uo6+AIa7r5v+U
f1G9XcAWe4TpnnWNxAhRoMRYZtyF5dvlicI4dEo4F0lzHfMF6KNrmRPkcw+gR/1k97KRu+CTTzhW
fDth9S8BAynRhJ2KmSgn6SNEbXj/YhqvzXqo3HfWCWDJ1lHfuYxIpl3OVtJXDqFaNv1XxNjCftYY
LcoaQ4NacTG07ehkd1Q9BbZjDW6BXn1VDMq+dpULV8woZd167XWJssvS0SHPCObhkZt5pVc3ySyg
FC+tW58S4enoEjggKqlD84f77gV9cZ93MW+OMa88OkU4u2M83WPtrZzwTdrzrHJxlOPzKWErxS3q
j8G0eXO2ovOEQmG6UbvZxybyRgIfUPqH6Z+g/hwcUXGScsb6BLU/ij0j0j7pU9VlIGAqsd3DIJsa
co05g7zaLXcvfSsi2uqwrch3PRiRHTvHs+daubwCYTzMMGqt3mabZIYZVWXhURo+RpJkbEo799SX
RjA8RzM0RLUtIBwcI0NoYPBI5yO/mGhwXAEF8tBKrI5U2qKQtMHYQjH+T+vdRyWjjCUOZBdqg2CF
OBJonIgu1/rNGyqIu5rGtODtsp+NbPcaBEA0z/bLKw7Ikyj/T8Gy0xA6GlHKnv2HDOd8vKGEroYi
svqx9kWohv4nlOyZCj5sL5dBDosI+A6dj79kj5JEkB0TvMG51r8iFEdyGuA0RajRpGEJ2Pk52Vgk
sjZmeCpgAQMTCaJ44Z1pAO0iiWDi1cuS1Co4pshZSshGuTFvxZOCa1VGxhbgdiP+qV26kjhzhaP+
z+K4TW5sgmJpjJAcHY1/icIkNFK7Z0qsb6CM2Jw0I89fHv8M6YNdOoMvCt0/CNyJ+YNWx6XHmIWo
ZRnCYGUv91E4UdTcwpvLMdfyaVOhHU+1DZdL9YF0dDd78cIHN4axeHMsRkY13rA5d+zdTd+dRdfR
6GpR9XqopWDCw3N9b9q2W+Qo0zIWqSv9hcGXBGoa+MI6/yb/sJpNIUb4CQZlExXrzlU8t0p6KP3x
6ls2eSPxGGpQ4YIHMcMiPAKFw1Db5PdTNCelbwEt7C8pBHLAxJnblsaH/+HesMrgxcfOkFh3Cv56
evDTAX2dZVezWVEs6A+0790sV3PQvgACjaQNDuE0i3dmWtKXn+mIOHQx+eKHB0dZI2CbgIGuQ4nu
dvSW14mxPOTZ80qqJxwUt5VAcF8/SYVOUQClfrqbVZDGZo0mQIiME/bA2xayZpyEMIn+bgebB6vd
O2cI78MDo+YeGVzeMPDk5jVoEjCkXaX231YrUlHi7421sTEd5YyPktuxy7Z53UOceZ75FhJNvZFP
/QGFw/tbkuNbLxkU60me2EXjcimepukZFzcoirxRmwKTq1lSE5eByMXqrGaAmBnVDmW4MryJQqZd
gebiZMF3I66IMM8Y3vL0xgKtdnA2C5WEVtEBArXlChwBCJ/7D4lSsHrCor9a212jIangM7fKoxCA
x3+oY2THcQZT+M6jTJrAiwmu+ZGNEGkihfzVekePXlvaoPOQxmPvM2N0ZW0Dyse5GqQhGyHfxHIP
m2jlchq+HvT/juOSF+gT4u5lZaa90QQHhOKKaetdrtfEZ0lun8QlSdpSMo7Totrt9CgFZfAiBA9P
GUBUCzGTMOze79h4mxbELwR66MezESrFcTdsF1oikIOax9Qcq7sQzZOSNedvCvLQU8osh3CWZda7
0fbCaQjQR1IGHcaMcJN1lIJNq7rUGvd+xD4y3wYMnEjzTxhtZG80WETf0kgVJbKE1BGFutS8fBBU
ARX9Qh9E0zAkBRIdEixMmuv3ZZTj1gnKtTXenSK+BPZJ9nNbVa1osnVgn7i0JR0vNK+DoT6PqZr0
nOeB7cWnkyJBAJqF5MOhOrz5dqD4YBK7XuGnB7SYgLFjaCQH/lGBGr4yPfNDhkQz0gmr46dYUd7c
pnnDTbDGbrdWV8iVR71sp5JIW9op25s6QVtak0UMGCEM4cvzl1585qQnqE3ulhZsJMysAequCDi+
RS/MK1UgI35xMyHsaNJ+SkXunnOQyCE3wSGz9QWUiWhsrEECvLUqow2l4D+0Isp3J/yBfLYCxCqR
Mch0CZQG58HfK/iDizaYgcX0+RwtaTjoyrY+Fezv07zdmd/sICFA6qIKxSKmwybQ40ANXkIbVVsa
zHIDezVywgFEOsnSYSzHkuKjLTuvlrEuWivPbVPAtHJ2QVCdp2hFrrT7nX6iSQqzKM10iFI3wJB1
mvuE10d5cQinHylz82kSnSiMey8VrFjD0ZHAQAxQfHK2QK9ViY+Dci18Gl+PPSsH8njWPGd0IVCC
pW8YTU/hu0hKgOQZjiO+KktHKHxjanTKRh4dpKa6os6fyTei7KHkXD6dsF3asGI4pinfu5xhuxmt
qRjbCVz29DpekzZ6qSJvSjQdEJA5Xiu4D0RvIti70LTjIgF9zCCgK/P8vO7fzF2JojPryqBBK1rX
AZ2NXyPrAxV9oT9jNtg7pYPo/pQWLqosIZuXpOmjQ26LpdTwGNi4eo+o9Uf2v6tMnijG7R7R84EY
jqgIIVhvP3joVcJEvat1bfH88Cr7wGvJREZkhVmCp3lRpf3oSbkxRtmKrj8dnNaFOuKG4wYTpQDb
hsSM9crXCzSahhtLZFyKn678ntWZw/yQiFLXDh5trcIOs+PC3rJPyn/4tsaGXoXxMPJBCsimMGaJ
QiXJkYRhZ4jqERFxIxXbyLGCeNR3Depz/uWigzeYYAUZIRsktrFIo+sTsJEEr9n2O6jeDuiV8w6z
6O6MVOp8HVCT6LKvGWmpDzeTC+pZ2QEvqiM82l3pog/bGYAPPJMb8xLVZ8SH4LL5SA4dfEKT4xAF
V82jOWRuH7Ewj+e5cUwLaX4qaUus3nSt4/orbr0XRmyp/FSubFu+F/WOyaCdQk8XXkjhbhEdl7Xi
mUvidpoSGQJWC4+yJNqcSgvNZlb+GOJI0e2pUlvTOLr8uzjAQ/x6fdfYBkpFcwqIok68+Wc8deyr
3TpKRn++LY1rn51/ehZeedRUhcQhJ1tdK7bxf8ya2LD9BcFHbqVq6Ay2y5OvIjMiJr9FrnV/Dlij
h1XyqQEcKuArfuUWeaP3MQ5KQGDH6av26NUiAEyzOvEsKcQK0eyasPJP4FZ6NmtykNAxp0MLxtGx
KlI1SWFXXBXppQweUJj+WpzJ/hXHRsusC9zOkifaAzNM9AZvHkZQnki9ThOs6EAOGXfqg6mc5XMh
IqV7zcDeypQV+PapWu4dxhliL6LNFk2w1rNItd7OYAOpMq6trblxL1KIo+5ssZV1lJICGu4EKqld
Ka2b3XGd3HlsIWU98XtX6Vu2v7YCPa1ThPmQMI9a4bF77W7eWmN4GAw5bnwvoo6vXBYGjgmCacDE
Hk+sG7fg7LQglHnvrPL3jtDPLJjCMN6QnpHteBCYIoab5LEM+lKfhC/ZbhFVQoorWhAhcMzdXSXP
KldUtDx6ZxbAFiWT21FmTZlSQHIUBaAQJdTCvn8LAOog5RIdgqdCP0dGqUY2CmbJZhU+/2gjjqHg
KXNLhwL6mh3l7+SrG6cutGwRiwq8aA9t/ccxi9v6n72X6pLrtZH7s8LOKrLcRolxspyJ40Pawcnp
pDe6CGjNy3P1rjlj2+NXCP2IKxJFnIC1vum0mYDibRN8fCZTNvtvRbeSdNTqIcpnzHSWDbL9vxi1
Pq8krcrW5XNEs2xgVB2s3v6erSad9Ej7qvRwpK56n6c695WrYrD2xTcLIoNjCzKY7rETu9+ICPLk
RfYWU2KgoE9tQS1N7COnhsg87ylI/rkQcvYJuV4NteBiIZHXUMawosjCq8kJJoEXqod79a2JAjaH
7NPoXHDmiE8ag4SlYHyhN3X7k/BF/0Nom7HoaveII9/u727qb27LwEKPDATYDCQAqPUWniNPYNSn
mj1KA4GqA27JNhNDLT2ZEBeJqSP5AByNKTbflyoVgLwMWL46eYqWCeI0PC0gF3z9W7Dw9LPVWe0M
mUZykkgMMF6gwXV7PYDOlxrkuQv1PtttZ4iA2pPoTzu5CXRqKJdU289nDymlT1cZuuxi69xxo+Lf
iyogIRCKL0F1HSlpUhneT/Bnn2L0puojjUh3L+ZAmuUfCug32ARvfw6Kb63wOFuhgPpxVyp8R/mZ
pegbkoRwV9ndy0nN0gOVV0WKdeUA0ObUtgEloyJ+DIF6tVrfrwPD6bDkFeaFqn9yLEAO97bhWAgd
yo6xEwHj+PhOAM/XV9BUjoYGkVB7CYaBKaZtH5P3mYtatwrHpOy8ELdG/sJLC9DFZZdD1sjqzqjT
LWMZ+78RoFatEcWKjBJ6Mk/w82oVn+d3Shb14yBFWYHh1dEyoe/UU2hz5EC06KgM4FBMJUHZDO/q
CSxnA9saPDa5P4lMDtSZhM5LhWpVr2cNATZhWgYSznHdWgzbZ3k2IHKcH2u2QYmEiffJJ1dBGfg+
37CVi7ufEJ7EY/WLPV38pAp3HC9UlLNgxkLt3giEvGYKGqIZtxs+y1EVWyv1rNN/IT/FpPbA09oC
p2g9QQ25SN8I6OI5686C3mgDzHrC5Od70tMqxIYGz9lDI81jkK6FCjd/uSjm9aidT6uHXeCXVVuZ
eEzMXmyLQqJuZWymVM4EqY2zI2qJmWp7HAvIxOPKPIENyJWYp3BIIJ3AJrHNAEqhpMei8lO2xiG6
30tL33moyu8ad7ZET/CqbOXSIUeQ1ScmYFarSbNdKiImY6/9/pNjt48lbwIiZ7xd1Q9EHxD/sIS1
qBuhJSrNLU+zWBusczYOerK2PXdy0p5oNd33Wqrd9gXX4uoF540mJ1tpZ1PRQgzAjf3Qi/2dbkRi
MKYIrbMFKeGaqE/0U8u4INh0AqhZITsAZvlEhWBXFT7uMZX2n8lKkn7VNccZjZ88isB8nW5Rz/jE
B6olRMGK59lrba/phsaLHf041/C4FxA5T+CH4qjCg2Q8xsxwUlvEU7jRj03imwxRZwK0q6/gTnL1
Zno1CxOkQGaCBY3Qt56F8UlWx6yfLDZZUM32KL0JR10Lxw0t88EYLn4vZreZszGvKxmy4CLSCag0
ZF9nMQSEgXvJsoacABqspk66WfD57LcOrfcHHSLTla+dh4eVph7EEnJ6kmZunlSxpAx6l3KlowmU
5lA2Ul+X9O1gXXURRskQV0iUdGCrpm1SHaakksqGI3OVY7k7aSlCsW70e/AFwWpUpjCre88ZPG6t
rPtuMeWH5jO0ARJ/hEBT9jB9b4pq/1DJuoeXraIbWYRl8ghK8g4h5vs4Z/AjU1V1mdkTfwK6Lyyx
bAD+C7ZnTBo2tt0qZ3DTajl9Xntg3/0Wxwu4wkJAnQ98byyXgaDLOcL7OBemSjLVZ5j2Uj1kMmuP
X2Dvy4HDGTqc8GLKccJIxpc2H6T8IZbFNGIGYb51hzupRC4N6COFPUSxcHT58OKRw7gXy/xuaBWK
qUaGRrd/CmeHxdMQb6NOQ+i02SFAaApicnDU5f91+FOHxEiDifMcSQTz2ieUV4dhVRtK4VV/ZLhU
N3QQFfOW1wvQJSYLXqNzU0kfbkZvU9EPaHBnwgi+HXycaiHg8i1aVHsebh9n+Xi9NbQRQCZadylp
7pRVc40+T+aCefPda93FIOp2eQrMCwY8LgukmurPKDxjcz6wRecKINObM/rb4Vqf5Yg8nOyJwvMt
4Tsz52l3kuweQ8n3Qqjy0cb4pMGSzo9kcAjf8S5Aw4gyo48+MHr+91Nr5+cZAcUKhOSQhb0f0Scv
15YSdqTfXqndcJl2J0PLC984/kcZBc9Prx+jfzAe08929l98xzgbxFui/xTWIctxUsTirRLYSBza
25c8VaeqDRT4IXx0T8rOkQg+YCw0Fj33nSf6YX/c4QxShIBGaGa3FqscfxqePdcLeqmB8X4dOd+Y
rWvBWD1vlOM5U+6C2HAP8NY1qiEl59KEusZuq5o/cA06i/wyR7cW4cHTzDk+M+poSWat02KI3a1D
CA155s14FOkAKrLT5DqaqdEFxmqNMP6E2GQCP4YGgPEa2L+OR8hNZZxweBml8QbzeR3okXw/zhWV
4iG/fQ+85WHkYw4sG3YQe9Iq/ZOGQSy+SwAh5Dm9c+U8Bis5MYAPgNW76U4sIsC795Qv1+NtWMbN
+1nOb/+p0MTYZKf9R5svyeMKgJNHwfAaJQH+/Jh7NjKQYb+iSRfdWnt27A0ajoK/+rliBvS1h2Da
h9fPHZ1+9Vf0IpGeyrnDuw/LcXae1qy3dd6fFUrOza2YGDj344d0mFqZ+JltWVdji2srRKlLoJwU
gFgXXauW+FRltVqKpaiFRk2F2B5cS24UwLIRpVlCXcb8ErQT9ZtUnMDFBGxbKDdzFaiX6By4INVa
kd6oq56MrNtpKyUou6X+nq6/0+Mh5eGDlyefO33PMd7u2sD22baLaxpK71WsLdedY+trpXI6VJDI
yT5NcEhyR0gEleRmPYbsZq/ykOeqWzpQM4eHsuvKVhxGtl8fNlIhYo/FCzh3CpaIpZwHs+F8fxYq
SmSUXbvl/WR4G48PjeMnBbbIbRgdS4NsQno7PGLnDRZhia+LN79i6TC/Qet9ZVtmkoK0Q55MNmC/
Wp7FuBoosq/8QZAY6RwFjjw/zxMK2wuaUcrNDppjNlhVakXp1oypift1O5dKyndxoij9m2hPZuOm
z+yls673UOnkTNQ3Ch3/b5z6qv/nslWiCQzdsV9rA/Pn/4OC/KihMwtOk1rLJtnzHm88GXG1CoWl
bMPjemAtqXYB/fyF5iqjUxIV923J67ZwEgfweHk1Sljq2n19L8JjAYcqCzqNjWXRxqnGuU3Vu8w+
nbKrdO0KUUkCsN6rohh7P/EMjXRG55HXasOxogSOGBLXQ+FZRkK5FM5g9jdcOJu/J68r5VWjdvrQ
tEnJaWroxZ6ij6uO0Q1r3jcyrxnMecEKrTzZ/IUGQXZj6XCnvQN00hgBgARZ4O0DlnKDmUT0zzc0
ZzZv3GfcdGD6MaFKRROBoQ5XGr9DH5hZ3I3RqHFMXryBVg/ksH8ps9z4XshMFMm5Hqmfz2VRMUWk
ObSeYMkdaKbn4Bz5AaIon/VeSd7whxliUMhI/2mreDPnTkQx7e6CkqXSIYasFakF0waLkTmi1O1R
VX8AmLCmlmkKtKQTa1cqkZ+XZ6UNZErgqiz9/8NkVPK58xuuucFM43d9GuzhcPYyfEXxzGpZbAB6
/JgO761YIsSXaCxGpZWn1ISP7K+BrdbbbNlXvehnoH7lKUrICMAk4cCoPAdj0rjPqhTnKJFH1Uqb
5Fqgq/1V5joY4nq1EezLFPTTkx8yuOeHPO5gWm3Gws4JapssGXjs8UhQOZjcd137tIifeS7LTd2Z
HNsW/4vWypGOttsWFmaDrW9OkAsQrNFhEGbOP1coa0/8cm3EJVSKjPxduRKX2TvJaONd0OIhasSy
fco/e4r3KCPhv2hctSUYxh+R7Tqse19uQSSS2VviGRNeF7gOJ3cc8Cc62Tpk0FkZ8qy7qBuvguua
WQrQT6Ugn34MoFu7ZYAbZxOOtLIZnP0Zqoz1egVkIG1kIAV5EbI/Ndt9pUtn0XAzap8yT4tLPY4T
h5mqDlZgUXThOCxBwePLzHYVc03RL3LH/FA/gk6ActrDvSB0CXTdWDqobJgenYaUSYnDzqq5IEux
FrVnOHHD7h1v67gg+hmnFaDFBxa7uVyzn/w+j76+BBGpTvZ2R0U6eQOeEGht53a4XM5hLinFCJSU
dvn533Qr0HXB3YtfHrcbeoZVh3zsJtgKWMJR5TEo5NxzBmgFOapPU65gD0ryLeeucmT37ESf4LX4
3Sgw/QF7UoZ7lsabZe/iLncGmuVIB3WU0V2ev8ReRZpz1i5dRCIK8QA0DBOVmrkgZqnRiAUc1HnM
vXTGSbEhvfnh5fGFBcFLJFRWsmFw4NgnDmHC6aEI32HfXsocbq2lk4vPhdwM9IXy23n8hzhuLzXi
vsOoHrOi2jM8ipaywEteCHjmzMHYjlob3P3APaQb2lxD08klVDygpvvmlTD3D+Shx0sJsrS4axLv
8kareV36c7KEhv3hEkdQhh8o9OLrwgbVdfAo5quOlT3hy4oGAQuY/l6yGFc7bR9wGq9HfUFuiciV
hObDm09hZhGqC496IQk+7lwDxqDSneSsDZl9mzO27bLH4w01Cc7bAEQ/EJmwaXpNPntpZI0TqJps
Q1Avm6+RexUYD6scEPxs4lXeKh+khpcwFVAjERoXS9ajDGgAblceceGVkHWBwgLW3GdmdZ/9cmeg
CGU0OAQ0hJQh98NbqWDkNsg4eC9hT8QVra61QiA5nDkVe5yvy0IVxHpJKFrY3psiHlwzLk9lzx7c
wBmhyDMsWS2FMTIl3inECu+8Rtr12hjTqVGpXjmxIOE+TrROt4RrvZsLwfvK040YuNWZ4GXVYZGh
nnJYN9LC46/Au7OU2p4CLpGUjaCnl8lWAn9NY4LkgLYktUUr4Of83jDp2Ioo8QAaBQVysjO3x0Um
geKYQkmqmueJybIjdSdCCHBfZbOCjmr7+3/Rklk3ZecJLmFhA6CrqIsUhiDOB1Gq87TOqSFYfJht
m0dMMY/9/ek7A+dzGKfqdTYiegTz/UvaEheTaYE1JrQde7vtWkZe0b4lzFn4BiTK9BtF6koICv7m
4oIybMmeXowZfSm1D0SdplevyqICMI8GKEYYbPfwM4O1C852Jz5BahCB8cyAPdyBdAp1SJqxjjoP
ah+D0qWoSiP5ckPtLjy3h8lvKUsSEy3PVJ5I54opS6igkKwrhoCXIb4gmEQ/OFX8HkxrmbhF0S4k
7CsUATcbqbU0vZqA23cWNoAZ/wduG3usStsONZpAQbAIZvcnhL2RCzqIsDBDEByudxiWb99ThYy5
U6NU/uJBxthZhXfUYJsQCat1nk4XGVLlW0pUNqSLGtuq/O3JmibvKsIu8gX+zMdekStwfe0QepoJ
mGzeeFEe4lr4r99R4f9uAENIIPf/iGbX0Kh2MH0ETjCoZVvKjHdwZzSMKUKVSEC2y3GJSGnBu7QT
buD//87S+5FHn3ju0pDZqQhDfLZYdX+uXO/vnjl3tjyo3Uv5op8Q6qZuUcKF42cevjcsKMM85tVj
fiFwGdqTA4wk1FeIMbihoa4UxH5ijpJ2G9JyOHCEyRGvmceKOjC8i84cPVDGYgwwd8Qog9WlMs+2
bwRVMS1vddAldEUfLL/isEIFofcvMrBmOzrlo3CJy1umWCiBkCdAx4H/kifw2T35c8l3cXGibf7e
Cg0u2YImEVq9IKQWUSZghiqL/iQXkgdGaPZS0XtpRPad4rqOqCdCx4+IeMrO4y3AAkAWWm44O93W
I68fDyvjiyM1BfgMCl5/PFGdcfpVNOg6op2VCVAsQuIM/FrkpMx89vcTwX/+NBaED7EBkCVWa5H+
Xy5CeYaMctRMs329FcEzNZ6DiZGrSj/+MDVW/TGYdj8CA79aJ84Q6ZcL1N/CITBsleTdlI0sQall
B6TQ9faaoib9RR+cHPCTIN+74k2fvxlncYp9NuuvB+zYIxvKE4TsrRdt+LSXvmRsyk9lLdK3wcFk
2BUqNUaNcC9ewISD0Q1xI2H3LhuimuKY6L3O1TmPT9lS8gHySfewuqIOqc42zwgyhZudByvZXwHL
9DzKVMtQ1v2jV/aTS6XTeA3IFbVwx+vDYspMNKJeLGq/C5qtB3OYx9juS3mGlpJn4LmjFGNEtUQ3
leVbkiSBhgmnXQnp1s0JIl1iomAkad+A10HaymkHk8ptGdmSydMHyXsd+JNMYfkxnXh1Ud/HQ2bO
AHZltYPEt7sI4mW9qRPypQZOdxus6Q+qYoL47e3bVBHATHP1thuqXBvmqU+ku8snNvT78i5Yt1be
CQQmVTqBZMdI5Nls8Ps7pA8A/dTm8x/TmXToBgND+W3MCBtSK9ZDrHq6bvx4TF7SQaMuesMYjVs0
YHcz25Y6aN0AJBDAtxkP4BRyS7PUrYuUudrG6JgNodEQ5R2Z4mB0nPs+sjwsY9OxREFcv7JjsLNV
W5ec3FiYHuc6s0HIwV2PZmJRIz9YqG6L+QwT6g2OPxnHaDLidxvoyjgBJfPSp+CqkbPTHlzFOrQL
shFV99tZr4/JV/odzVmKLo94njCNdJ1rYKQUwclKNcfJ5vs+OucmtF+EjQ0RApVydmmj9i6Ztra6
ptOFCbupSGbYDuumX1Xqmogk7M9dUupmPzjZuIerFnFxiZY5EY9HEj2jmwPm8eWlYATVYSlCEdf5
UmZrDxApPniIM4JNTyjK1wMyqxEr1fTQU2clxLx3Rv02WzAUJrbGEpL/77WgiNgQW+vUlddLWw01
xC7IN5Unz8U6n3RvTLXqAPGW4UDz37JFEQ8dYeFTUVxicWC3o3cVWTaLUbNmuPlGgKLo8iZeyARo
oBwEhJzKbUM6jrRGqPVyqmiRTtMfazIuGz9Cc8HmgaCbjvjGKhv0VU5T8onoKcbKeuataiNmF47W
ATgCqIziCRhPHBJkkocqlE1VKaROxu21I8bh8shq+1lphtS9vAskMWB/4GfP2wsea6zG4pMrgXXY
q9BfWR2LO3w5JcpuNkm8lwWZ1xth8YhFfssKtUAgZyVf3OaEihOW3YPGJhVG6n1MqDBbRbzL6t6L
wXIvc29hk/uN2VwLr1/gsy9BOTTFDx4b0g4G16F/tWsgsGnlqY1bVo+ppkZ8xKlvl4FmQkMjVFtp
vkTxn1gRCPJhijblghz03XZlVVFDwnpetymkDAu9LiWyc6Dxz9hE7rsGJz8OoeOlV0RmqLGwozU+
bE1CVGX/OHbto5l3tUwQ4EPDImJulfLzTttXPPkYH5Mo359jWWv/rMNMxve0mh4F/TxVFBSfRuNZ
2g7mQZFyMKs4GbpHs7VRFYqWP/0CApbzg18kLKHu+bUCOA1lanVPyi4y6gB2IWoO+LCkswks00Av
sf8mcQGrM5U4gjawW/W7xk+TW0czD0etLOlCNb+7bk4AInuhY9ZwYbMmRHMzTOynTj0hJeJPGNMv
LPcs+VVeUtQsx9H06in23rhd3yyV+CSDrZZzzmZ8NNg/yw5J7D19PKx54/GfGd/CglwXcLpRT1KD
eu6kMljnl8ZCz++n8rYAkpOPj33R5CdJxX+sbxv5HbmaTeWeLdGxv310Yj80tj5VOUDNP0xCv6nH
tQHu3GrcbD3Orc6h6tkyeOFKEpAVhoiNTtwjFku42SSPVCwZX9PWARactysX1DdIqO5wL81nVTQL
dxajG/5FRpT6Uay3OMlkBmiM5Ab9AVOg9F+EWSkgtHyVuZ9NIDVWHAyfGTgVG6O7ESx4L+6ojucM
a4bt5Fpv5rUp2FRKohJrSGr+Fev/u4TRuGjtBUMzwFBTJT4okRaB762+HaDGSRj6i7FvneNaCfPH
WrhN35wfW/PwMPIpK8/DKNzO5Grc5VzaItPBw6uCowSKOZhAZAxW6gx9SM9CACjjyEN9QveZ828x
ePp0NhgQy8T67M4m25HOZTeA7hvpfBC9Yw8DsVDsBtQ5kfuBht3CqkFNmAUUTY20RbNQBKa+Lcvd
dFKNnZVQxwOv9tJquu2q0eEy2mWDyiWnzvY8y2snBJwehTOWVm2VmAWgVHWeRtyKqTix/s+LO9By
Um1TCAnMIQKylNUsJVtrABx1mFS0OzrOLtyp9e44PAz+1S6B0noWEQ4JXXcgTa+3RxXMmenmeNCk
2S4nAsd/PpE0rQ8T89SStrc94B8oFmRqJ2eHVJx/K+Kx4qBVIYLVLfRpZohNyzwc0ogKQYHPRJ2t
rckYc7AnWpGvUcrjQCcE9cOAJA/jaX3abP4XMkHAhKwfNf3OoUexHVTLrV17CCZdVeT3RlchL5aG
vdvfB8O5IFL0bP9dJ9vZ4gHrgEHuagCDlQnp1cCdnu2P+Gwz4Bi+ukstujvWP8gMEXsaBaQGyOn8
HKEjCXBoTa/uhBbAMwpSN3qzZ4H1cRwsONueGsSiFip7pgpH+uuXsmVrRtwkyeNBg8oOYxx+TXpe
J4SmmzojFXJQFRn2LcE3IeLb3z5NUxeR+lDXWmjrX1rxx4YZmwvE2Rw5JwR+vVHFAi7lyoCUDe0P
nvhmrvGiT8qL5S4A1VVBPiqd+ucgidSDvB7L5NOgXdPfe+gbiAVJM9dU+X7ogfqgNHIkX9tMGoay
phf97AUAxc8tunwsyw/N+PYmg0X9RV3R3Z0R8DCDmSHDXg7qm1zKR3j6ArM4aUwAbuN1xvLpsm9C
JFRLhLvtnDzR3ItYTzHpkWXhtCOoJBRaTsVKfFsv15b716JU9OBT3RW9sJ5hNVK9V1Wimzu/ZE6h
EIPt9N6OR4NK0T/IYvVdy5cm52q09bPtKtbSjPolm/zKhERUfdzJpROjf+Cs1vY6cUh1uz2fmWrb
tt6UUwLxtwQ5ARR5E9x2E6tP74Dp+lDD+XTkKqZKzbAb1gRYvPEnQrjvOrMqxOryIS9RJ+IB3OWp
IwEtXQNoOGJPXDsmx+StTzWyzsDGqOvMRjPijvQdgd+s0gjeAA2fcwDXA4fN5GCmEKmzuih7rjss
Voi+i0gB6Il8t/is5e4cem8613EWYYt9YbYlBhRcmtpv5ZavOue243WeLrOH9HTcbEce/6ozy28W
aMcM+vxDEII5d7SyAhcLBUXq+svqgJYlz3jN15pX+sziADyWaOXGB6+swR/QeN8Sp4zkjTyI02tC
cMgzwdMLI5a2/ZkvAgLRhovFKOwYlTJavIsoI969n10XPJxQZuVTPAxv3dliAlAGSgnfB/LBL67U
BoiBCgHIa1hWGfAXmQy8lMvlH16smkcfLjXkDSYEh7L11neruaxCe8b7zphmJtT7ta6x8SwQQtTG
byVlv0zVvhBuwv5bKVzkR3MfbIBrs2F7TX/Ri4H0xyhZl8aYvMNt3+FZugaySkQCgchvFn2b7bzq
wgNfabKLbKNWYDmKewapd2VKahGx3VKKQpuDvEivCafPHjQmmTZsCQGFqMWCN1+uPwtXoCX7Z1Nh
YgKBKabHvt6wLNK4J4YnZF8EqlGp3AEtb+3t5joE/MlNHpGI6h8DGp5x4SthqZc573wGcS3Ny3OA
EkX2zG4ma8rXWGyzqYJ631EJ7FCuQQhUF5p5DiuiDo03FKmtT6StJoXxAS3wB4RfU7IlP6f2Vjt3
J1wcqZtlzOkqgTBqrSezTDl4KNrGsRGVuUuQc05wnmiohVYqoHJBh9Ejyv6XhuHWr1i9kIxWGhXz
yfMFAsqAd7Ud/yz7RgFv5ED6wUQISwn4Vk8AEdylLAy/lxWs1Rd/jV8W8i7G0y4vwaa1nxR4YFT3
H18JcZivqyMMCtWm0VnvOyUHGqlWWAILo+3EEhtjpvhnR5/RalBFiTGjU39CQjeIazzHDZpIdnyV
k6tltQVLkJnnlEiGe1TX588hzOO8iIcofW4bGDf+f8vXK/KIhdbd/urFwJNU9l4QI+sU6kQerOHj
jxx7B1IO9gRVkc1IwPIgwJPAoX/ie0tnRJd/b5aBbOW4X4cLzdsmEfWKPEPFkNTlrBMZPXXtSxN3
z8Ce96ERUWsD/533jeODni4oBYXsOVUUPqqP+IC50iSWibovYaNQJ38+RZlJf2E+PGSdSJ0FMQu0
bTGNvjyWySr+wYdeYB2I1ck1yi/4zOzlJKYyUDQCqk5DK1bxfHQfxRFkAhBvYyxrw8WFKEOCsXnk
hJ9OvPuiS89MY+vVj/hfELlh8HSdQ1yXNFsWHYprWOVvpGY6vceo2hN11ipLk/n7ocoOISW4ZPki
i/A3AESOcT7aML+GFxarsQ8EFo1OzGxwWMJ+xx8OVkvSq3vgXYgsoKGkyz/9TIbNB5/AB237X5TM
XQOz8AL404ooC5miRqawLbuRVeOb+warc6WuiW9nz4EKT0xrRCs+dA0H13Cp0q+FdkQxfgoTxANS
RYRd+ge3zUlKgTlMI7xh6bPIC5jsMdFWKp4H1ITRvviaW0IfAR5wHMqnbyXqPJxZTP7EFf96zJRt
ELeW42BZhFpQiIpXmp/WN0R8DXEvCmHSm+ueAjBGR1d6JHGsj6iHLBp2B09wVpP8kcvZ8JFhYKHf
R75874dtnPWxx4W3hmpZ85mOsLQv+kVdzarquAzdioCJr6s+i+brWz/AtB4HwXylw+8uh/NBlnRl
epxxcFXp5nBZzVKv85FoNgCQjrmdA6vMBpwUbOUnRPpEmvW4q0PBZpiM2X/QY1FiQhCdacv2m/nn
W03i0N76Wt6/6ol4hYpFjd7MUYK8YxEaUf4ToJ3Ipb/HEeK9xq4MjhzKXZut2l7omtJ3nj/3z+y6
F6RkM6obPEGtgcTYWPGSDZmZH8Dor0zykf4Qu2sJysM/kYltw4/F71vU/BRCiNV7X4uTJggl9Eg8
X2pDVNHvx6GXaoVFZwXDFG9JH2pkR5qoZVz7kOELdJgKLdMh/AqxdXVQ854QHfj7WbYFK/emjovA
iUNHFj8qSVw9IBoM0W1MJnS1zWrqaBCcCZ4W1mgWG+XIALyG/UqWvK0pXBq5T5AqhInthLVlAP23
zwhDlPrvlZ5G51GR5i5wJ1NVVb/Obv3KcBJeTNOjnAC8ZhinWNNfVZAzvnGhuNvpEZsPtM6cBGFT
09NhWbduFgv0x/swOrqPhGLn2/Wjn/njtBoOEHmMNM7eWG1UyRzcmEe35k5FkgdKU8x8bPtIShSc
VBFYUxx+ApjXAm4fViu/ndxbBG9c1rnMEThkw+nkM7aCPZfvjNi+uXNwcN0keS2nT9/c4VT/hq+p
P70vr1venQG4cQHyREOcwPFUvtoy/ae0sD1Mvzm3FMP8G+SMJzaPFsAXt9R3xK0ULf+Sk1iRQBES
6PdD5CyMO2QO4zwFEgPeA/2Cw6BTDuJO9jM4bGfJv7VLHbm/AG7CaB5T/ti7XjUZ3vDWfvo6h75I
x8vxkcxAMs8AeVBbBa0sPGC8cgVU/ygjAZxFWH4pGQ/MbYd4LenUMaec5i/DBT8xGVfGLIlWkDe3
dtxv/naMf+GeSJciM55mhdZ5blx+EGBGWhVAxJNrYnqSGW2ScQCF7nqih0j+T0jw5Z8TvbbUB+Fy
SZT4BeUPDdxEmtiyrJaJJcccMPeQlDPNJh3cmlejyk+k5+U/WpEe4dZ8fJiL8vPkdHZrEzySW2FG
tar9WWc+2L8DzcnfcgWp8XEwVtQQmZ3SL9s6deKYDgUegT9hA+F+9si59b5n+dJb1m+4TM0R6qD0
rnC205svYdevKGS4Eqz2Ofh8tuQ0a3TZOhqOGO9ovGQarigylYryYD+j+I+KBGmB0Jq2Ul037PkZ
NByxSHSYziqSOlLuwFWM3PFOePZsDLF4kSgqCNMQSbge0pC4tzAcfB8uxBQL+c4YlJ90TAYuMgLY
Wec2lgowaGh4LWNXgkeddvkYeTXG47j0CF9QnRN2FqeIZyCRDPNeIv2omLaUV5eiP77DNRt5sMRU
jTi2XCIEOb1R1osg/TeNyWuCoLmc4CIlexCrWxfmQUFk5v5e18lkTLVxxLhKZqY/hiaE9bCR4EVS
Ub5nGCasuiycLaGFsZg+QEql28j21t88p+kSqLq86WXfhEFp/wNt7gtEADJHIeGe0btx7ZqjZhcY
ovUImGfMDoQtxjlJoUdK+qclD8A2FsIEXMrdsVczSk3WPSNERqPm3+njUgjnGgK6EFOOuWZgCoOn
2MX+3VXaVkNBX95JxyebSxAkcKhfsrJETPpKt1q8aMAwRwsashnfB1XDsPkY4U41JmZhMPl7Kp8M
JYILjNwBVmj0OgJBC8jCsxOFtPjGLwHSx/0PWcGWcw4uyPYwmLUi/d1CxXDr/kHQF6rkYuvjOlZF
01aChbTAxIAI9NDf3ZEiBvhnoK/GYX5bX0ZDPh11r1xvQObcBIq+ERqAepdZf5YFmsq42vjEfoKs
qxyzLRVT8S85iNjs89zZp5wJFKnawWBCEnLmvyEPxlzBagXnRuJPcpuSD/VaHmlcCgJ6cjZfmpnD
La5qquUeHW9E0dT2fEFjOg/0oNbnH3Hf8yI0kepKoZb8b0oLoq0v34p0n202BeJeDg/vzfqiWQlh
GQj4+/qadjPTagzxpRWx35vRLVx+DaJUp8TGAEK1uZJ+3pcRBYcA/4A32VCdQGkjpq3lu/lpd/bl
LgZBQxwm8C0ndpn8sR1fae893SZP1D4/VtFtRtZkD8uvPmJ4hh2BLo6thKup+BVp/IvIp+HY5fkM
BuxScG6XeAM4V+PuRrd7di03MfW2oba62h1J695BORHmcnKOkJwT6dWEvEaZ9DYAzvUD1S5felZe
/2YXew+kFy4u2+ujvROCEUsNYjXbNRLqy7HPMFcdvjp1p0bU0Q3wmXo1ItI3e5K3VyDRiNlYJfuZ
fLB32bUUDQ9gjlsT8CBRiwwAEDlZzAZ5MomLvm52FiE0CRxbu3pgpQQKpbF4feI3Mb17Y0NRRXFz
JEdRCx00DcRMkEL52Cl74X2hoDHS8rqf9TGTW6YTYe8BAago5cNdU4U14J4B6zJ7j3xUaotGSUEO
KMaWPWJmIekucp+/T2RzP7XdzifA3u1m4EOatN1XKsJDqkqv3Lyzz7gy3P0TdMSQOtWJq13zLIls
rnGCb5PW2/VZu7njKpEx9sm/ADsIr3EkVVm44Gq0KGHlkY8HfDkd/1u7Ah22SFREwLDnNW+1Tmj1
nrtCv+M5EUYLJka3yh7ll9B7SpHN+Xz5Pd5XVu/d7wbzWItNOFR9bNs3iyJSwJ3lOd5FUYeY1GDg
FuljrHgaSYriMo4f/MTccEiRUy9X4jkZvXRaAkmjfbGjn4HKvQflIXhNAcQiNVlSbpXNzMLE6BKV
LF3zJK0QtUG0LW64clliXYvncXzXFM/9m/nTPSycck+d+lv5hV1afkUfD0C7kOjQe0qrDlm5KdWr
InbKWwyoiJgtpKnwVrHy85jc1h+OIFhxnSsEy2VNkYJCo+cMZjqFv8+Ywb2PbUYTntk6rkB4BZ/5
4IVNzwsyi4xLSEY0H5PZqFz91qTxjZSnGcfHdRNJYvOVlomKCzvMFdNZIlShxg+L/z5MmLJaFcTZ
kD/kZXhlRpB5dkZ46hMCqU0kMlCer6RH3D9D21djSJp4NPho8B49wVExolpviR7UxHFN2Fsg+llh
Qj2VBAfLvkl30vh7QfjM1pkeEkVZuCVMHkqz9MdP3lsOjDGkmFarbQa4cNojplNAu0jbK/AHZmAA
hnDW1mzd7FDVfhyZi6ugAHXpvmZNf5mbkk30GpALzl1uQVxe3jl4I51GqCku5jRBS2ri6HQSatRa
6l8F9DR94ixckPlXkdHmxgm+nPNricOijY+FTpAaYBmDLbQ9kdE9XhVq09vG5z3B8OFvvZzRPVmP
Ue7aGe8cn3UOo0fYXvWiFkVU9qOH559C4sSmTiqk+EQpYFfxtQiqYfqk3GJzeUYTb65JL5mQrueC
n2GjxDGutBzHlfjuy2s+x8LEj1FVwxqv0td8H0lKkPqMdwcbMiuGel/2nKVgPXGRSEuggL+Ns04S
8O6fnj3C5dx8x+81sT4b/z62ZkMaxERA1TL2yytQbvsuHnEDstLGj89pr8TKRpdp+3C4+ouRD4p9
ksXpstxiT1nIVrR0B/Ec4S0h2HEe+YGhW+4X2vs9tBjITrjghnmqdE/I0nIWvOT6La1efmev8VoK
IiTX+FtOHO+5t0mBDWG2kjGHmCiMoov2kaWHiZKllBsoiTxhzFSrjl3VVkznkJZCCHnnqLILRIPy
116g/VKPf6sXPkh0JLZ2573Hc5tmeLHmq47RH5Qnj8x/xwVfDgAoyNE0yCFubEb+6ZoueHoBEYto
U93TOQw77vkPw14qWX8lmMc2wSZbsCwfoqsNiCGmBIVOwK+uBudN6Oue+jQEpUegSyqpeZFggI42
FP7BnLsXcVnzCLFFcM7llzefbeVo28x3LMuGP+/bpBMK3lhTDecGDlw8lxL3ZdVgE6TGuVJn0f4S
eQcYwQqJHsb4MKaVKR75w3GjCkfVANZc6+2pw0ODiW9ulFg13OWmj8nJJ0W1/ZJQ7zb8NSNXepVg
OEd4t8RLBJrgsz0lDBa07kFzVIflyxJAlGL63gOman5T2FoDntAX02NrmrXRf4grZg/MGyDKLmCF
vxaF464/9fLhLHdKux2WmiehwDajOp0j37Tw2rqp6qs76uA30GjqL5IhPFmdy5tlKlrbgdO/5XZM
iI7TK2BMHZ2wPo1iHjbYs5w1D8/xrXhDJ9iTxsDDNh/vAFidOHZeM5acqfpslJtZngiA1BjTOtTp
jB0QegvL+3xgMj+V0QoYgbA99WQOP7KaclUwwNgbwRAJFgJiU9nIRrEcWm5S772An+pudgZR8ko0
bGmWsisczI2JklNo+n+BbnxZB1wQaNWLxyEQ0ZkQ+O0j7CCpfCdSKn94+hXQDH3CSPowF9tw11T4
61mjIMddfgEf0ppERxZBULVNy30JVZb6snew0vn/DTPMfdcjpnBeifVXhC7IZxo1qRLkaQ4+qbo6
MatxHExVAKJhyXfUMkx2WBYUIx+bit/x/IjUIaHMq4IlYvIu12mM3OL3hrxJ8I/V1/pcEWcnd67k
hsexJ/pFiOaMS+35fiK4FmdQ5MCW31aj9iEFQ/M8jK3IjyX0jvH0D3o00ulNfmN4zobRDJTA8U0d
0ULSu0hUSR5L/DQjRZcBBTeBqV7jPq4ngQMomY4hUqp51UD2ViktmPabhURadnduxxuq3FJRNQZs
AW5Y7ONDLB7hPMMUfcGB4eYNUKazcIcBnI/XFpl19tczr1JGh62yCz+1tAl5muvYaTzjlHcmjjz0
Z6qAFc9xylygZ6jM3/RsgQ3jfyPxU9DZNJY2z/9B7EjSJ0xFt26YKiyqKRVtBNC/7aDINWdJbt6b
TOmRxpV0amnqFMZKFeOdSRorrF8ElJe5n9YMmfOqUjjIOaJp7Xc0g7ORv17y3HRnaheo4CVSiz3o
Sg9AugXUEcS30mL0II5DLGbYfntaI/sxJqeBwfdlHBOcUQPLD+7NjbOX/YMdq5zmHWqK0kFaZ1wt
8mB88S9T/j1pPWYvDdbsmaVxHCim9WeVOwpgbPfHO7EDao5qzCBkTCazOnolGgpBUBmCfagU+eJD
+DgQDbUzblhYZc3L5yQD3nr3iSzt9ksNfQZCl3RF4T2RqrjUVfKwW9fAoL1BTmlm2yt91kqXvVQr
Li8AYZT65OAazMcH9a5AtLcFr3evMxvjaS9/Vu04dCDrlFv+mHo1BUbuh+l7fBocnDw8ZzpP+YoM
EsWIU/TPR411ogL/5Shx0xKiF2UAkNQVB80aQa1F/mqjyo4e4kfbptBR/6LVFKS2JGYrZBMGPnnq
JG1Mf4O64y2B70krc499ih7nMho0cC4P09+a81MO2GZV8AvQX12+bRzz8f4wXlscSQMjyuXdfv9l
hAOa9KzdCaxP+R3bXqkBFVRprfCfONgTZsCG58nHBkiudPpVCdjCGSz8A0v/r6TEZlWphUy/8Hls
giUNZbuOwXWEP3Y4sFlKOD4aQ7ftSN2YxfSitKnOmdkJNUF9i7yozoIOgUFPwwSOpaoWEAMqtq8S
IoM7b+l14afrjIBIxEi6D/5gaa3+baSVTkkHDP4odm3uTOe5wAC8cMvilzY8zQB/jHlJDdOp2aCm
B6nsriJCCg22oBy4KV8NXonZC4opSKsnE67QYW5tInYOjkPFICbE+eZr6yFeEIVueS365p5Q76S/
A/n6L2wvrEy5qnhG+x+XiYMZ9+dXnFpc0+mOt/Zhg2at1GQlr5xgg1WyLgnn7CjwOr7tRBW+lVa+
i9UDZQ3TK1r4ceipxKp8q/wyB69oqXlgoS4hgvD2Ed/POR6VZZonsdfjFdT2nJ2L0dxu1rG/obgX
mQGm/wK3Ko/IpNfTS7YO0Bsi0LlujhTuanNX1cpKwcp8xZHFrmrc2WvBjIPAq7eS/dw3rKyr0vE7
WQ5Kkv9ySdHjhZJa4A7bDWFJx9eptRyiCJgaEFun/HQ4ynMWRCv9XfuQZXezY5Bj50WvAK7khDck
RRkl0kN5ORw9uzz3cz4zwe9r4lF9D9EbisoFS9T34B8EJZ/XD3CvMw9ajhVu8eUq8j701E98sPp+
lmMTTmhTyP28qy6f73JJApAhBALWhbtga5XMwj3TAtoQejzGyfM+zyCsyS+vwHxpjPvCaPUm3Xeg
4/+FxtQCB4+SX9fVmOcOsBuAlwTyfgzw7ggl/5YI1w6azxYsC9Rb9kJz6bGE1SPZ/Y0angrES29x
a8DfrA6ezp9P848jxpBKg7ckxGCx+zRFzm+rMtwK3qMk7VRTpkP+N3X938HsrrFoESUAbRUJxVOQ
YYIPuf5/06N1JjurBxszXG+wLEVZpudaaRi6WjDyImxge/d7oMr43tTKxgpoJsxAy1RYnOJNQlkn
85J3ZT+JxMucJUC6zgzPRdt0ciRs9rFToNFX39vZQMF31r7gAgq2OYDfWoE9gc1WKGDFivJky8kC
VOddgR8g+FpxkzywLQEgKUsr4qIBAEmhBArDYKmIiFpgfuuuK4RtSYDNHhSuW3Ipuou8zs2B76Sb
4U9taDLCMHnzWXEh894hzMjmXTJ08m7hmWvdS8r9/eumvo6gZvut/VTrn4HmgL3jfqqgFpKcfa2l
OhwOkHp9F9JR3eDafmGddwIUxpIMFpVpIjkjoZbIwDsYqtYpPV+iYpDeGqYI+7BkceJGYw0dxazu
YFV7iXTTm56/P1p60yKWEtoowfFdyi0lKMsVuD48VV0RHj/2TMC5r0WNw1euhY4M66VsN6m72jGP
/4hS+il2x7JGG8W0iYeATxR6kAH8bwUJWIDmYn3yNalmnKZ5hHBA1U9jzPO7bKOdr9Tn0HOdZ19f
LVPec3fdGakazcKJw6bcuzsho0cxV70axW0/PqQnfs/P9O5HF2vQxpUAR/HbXuswRJVrXmQiH9lU
Hj7Q2xoHL53x7LjDl/oaSimtg+kZVMysdPEf6RBD0qWnWQ9DTX0gBwFBPuIOzC4IOTarc/LfSQtT
cyyLScBuy8PMYlnXvGvWuIpqZ1I1EIE70dY5NLzWW81nHhXzbqi3uasnzYR4fj7XkDtk6rX2s7X0
ZSUQKnVHbi1KXtgqz5DRMvpOsColnlJvOaJo5jx5HZ0xd+Wy2nIFa0w1a40MzsTLP+isYy4cOeOy
cX5+VivOULPpN6FJOePOZxdfv1gs30ypgKEK28QETlx65zsfR3OAs4s/hjN/grjzVvOwCPxi9nZt
t8IGyJlpMr8XmOfj+VJ6mg8DnzEWwX0NlfCLS+I7D1yB9HqD/KltfkrfO4CtJpP6ZbKqk+LswwFH
ELLuJkAR4vDTk4KsiUHOo+0NPMBXLoyDP25Bx6PUvkEFFt2DfqhxK8PEmfd4BVNl7UveC6dwZraD
KGiPUSgtDI66mivrZnqSSf/EVnXcNzGa9NNp2nF9OkgH1Glwg1Xv3z7vJHF0v0GqH/Gz8RfMFNyz
oevfhCivdW0WQf5HJCsYJNlG9BecDf95SPjt+Uht/Tm00aW9U2BEsMnFDAt5ndXaviq4wxJ9Hqb8
a9+a4wqzDKunqUAsokqcKrtEgEZUwHsng8U0YvrmvcoN3RtRgGbcOS6Z8mpR0hELJPcfQpXllP/K
6ScEcAhVQzUYeZA/rQ0QAoeAg16O1mqK2pjSvZBBzzc2SjTjbMaMGPyJ9Do2cO93YbRrElypLDhU
pM4iXn/M98HYNVlDWYmIKnxWLmzFslRxHk1kVdnzr5th5MQFcOQdGqQCiyOlDKCC71cIOFqZlxU8
XrVUkAvd6SNBy8ooH9q5z5zKLiBeLGNBS31E/stO+PKfskfbl8oHPjImInv0N+5+j29Ye+Y1+7c4
e8lrdPC9rhVKCwNil07K5g0YoXUxsScnt0IRdQ84be7CX5cOULMD3JliCVNHz5zi8p9ifCrADfrW
7qZeLePi6n3t4/QfhA8R7ivCRyhJLBcIrcbB7E0B+pR+B+5gTW2UpNqWOkqXV4nSz4NTwo1mlSO6
JyhBA8CCaeO+uXhrOARweZ+00VaP9zCCzdQZ3NLmyJdDUTnhEcgdVhx3X0yIX4zrWm9ZjfjnWCMP
yTln4V5xzVcQaZp8WgrSTSqriLb8yJXhZ9moFoN+xLB9BsAJ7f+W43BI5E6Nc3Y8xKMOORsolMdM
48VDYUxovjzVppErvahKOrp9KDSd4t9Qq3Ij0i/YZ2xFdh+gOTCss61XefBcDY8Qce6aLGT34pLp
d4A4qyGPisM+JC7YBXA1LOpyWX2I3S74DVlHIfSazaMDc3ojY2Asm/e1Sny4kmTKBSsqAoW1G+Hx
m3yeghKOVTKKIeoaaeksRe6ytK8obLQw3Q6Jvf35uxfxrStSpd0B9EUvoLASPHUtkU60tSzYMZMz
8VvPmCZ8eCuTvRsZltOS4PBNogDJal0d/zQ+WzGfOnUg4O4CoUKHy1b/atGhvooIVQSCk5Yevs0W
ofST4WMg7uLYQB/aiJm6A+IPZ/6nSKQcX1cEVcUkZwwDEgGb8GZERsxWYn8P4gFtqG0mwmyeO0sP
qvg1arhqPJvzFSR74IpwNQtA/vcFVaSLd1V+W/Dy1DIGOw5LK6BaRsZs4kfEf0nqMlwT6xUWO1Cu
pPWFAL2eQOzx6VeCU0EOZ0APqk5AmTYbx+NqVJxlMxNUhQu7n30Jpqf9YqupJA7muT2yTWb7d/Ck
DEMrkGKv0dmr/I8dr7BSK0+hh8g4ZhAktav2AQjyL1GBV3cm+xTyH2OlVKd7dU03Teudym5aliVq
oyehiovczWtOankZxmARViEDVNocTQ/4G3pOpmMbL0j634V9jCB9741sG9yaC2ZVFP8Knr/bPw63
piVtJbDa+SVE1SXmKY5Dy9d9WlZlGS0vy/ozk41+7j39ApzATmFGqYxGApG8wl6Mm4wPeDEWdFnw
xusU4zHjvhTXzO/kgQm8qwTUV2+/JSIIn0s1GyuWV4sGxjePWcEobRt6iMEQopEFigtVWqgbACgV
r29EKDAuSvazRORWt6viYFVQrIyB5NCpV+nhDE55+RUHoTL8mmEvxpuXkrLRXHHxloNp9IH0La1N
ybEUM2x9nnmZZFeR8jAWKpLyDv+pc5AxcrHdTtTL3S3W2+RioW+t30Mdx0WkeFXnkuflpffx7xrK
Ots7g+kYJzXNimCFyBzj6E+ZbV3fYdOArTwxr1PZAL9dteACmF5TS7pgdtP19Rsl2QXhplT2FKyk
eTFOtiK8IFn2T05p6tTT06k7RqvJ7Btz3jXND0E+eMVzhltWNs63Fuj8N0Vr1sovQfksrf0rH1/E
fTbEvjQBJdYX/pVjqA3N84IMPQa+UmX7YDMQPQ4d4+39Md0B4M4/h/wYE1jdghn8RGUrd02w4p0M
2GEk4Q2tKehDBeYp2OuuxCc2ygSQXLMbhHFUBGWLkQqmUZNxpXIM/5phbmIlTQ/cbmoalAQIJyK0
+E8UmsqMoH/rUTj5R/wN8+KoFl3ntu7m5ZiTCBBFZUYtPvQ7g43vL6hvJy2EiRqsQtNokeH+QadJ
p/R8GU8A7w8RPDH7L4mkyVw64F6RIYY2Za67O0cT/iczIAbFCC1cX9MjFtlBAwTo8qRd5MsuN4As
ZD0JgsW6ky6PGcbqvRgU1Ln/fszN+a7O3MGqZ0ijyhLczgsV0B6zkfIMvWlFE3wHFgw8B1tJmpqv
xVbdMa5ECd9L8Y6PkT/fg2+YJurQr1QRrG8OvDQWJEuLpxqvpZPnDI95IbMfmkivXQZe3aGXS8Kj
j1fFY+gCXCF+epnkxw0ZR4+xvAyMDZK2Z3RkZzxNyNaKfNtixyj0rZB0jM8OK42sEOy/hKngPLrT
s+bny1AW3PE5BqpBpslXUmiBoIlCxbYcWObW9B0LjUs9XMOC+ujUKW/PPyw380szqlx+kQ/qA32S
yYe6I2KOqJc3jYFCstl9MC4F83IW51CZItUuEIPD0xHL2OhGuIr5tVkLRD2eC4SKbR6QpnbLV+k5
sghL8x5qvkDJCxwtIVwWbMxWbTv70lQBiIyjp5RcM64Dx/57yJrrQfB8is+FjZeQkcPotv6w43KQ
qQE5cRuqNNqIW8Dne3T/pgdOLEwkmG1bMSLuAyZR3etiF/eFI/qn9r9WZPTg05guKQlDeOJ5bqX6
ix50rSuEZN6R2v3IChUobbTRfRQO5XJZLHdNvUSxIpPrTlea5OZa6OP907PUeqL1Lo1nvJhHdH1e
hrSwoxyjb5601+M7MDxkQi8hqvrxwQsH0rc2uN5KubhDl7NPmVG7kkvXWxBti+JQJKF8GXCELcBf
23IqPLbb20YzJapPd/bjJNNJ2ouc8+todJ4oiOmStq5pjKjCwCZzzZrL+dwrX+Y3KnsU8iagdhDr
uNPnfvgoxAQiLFwI4dhcu/NLJKHh/kCisQfyf0oUE/C7gcd0y7lc3JXfAArpPVcyU7cCCgC5+kKt
vwaQsAH3FLMCoFo0Gv2uqoSm6/zku09JoTAKOJC/WMLDXV12a2mlJqlJgYT3wdHHg+I6JNQISzXT
93WEaaUxXzAafPGjtRVelDyh1Tz0tmbpq/DV5QDDppxghzlzaf6+FKxV+wIFejWpFTNogXu1zokO
2b40TKTZc8k8XTcmF7dwKoQIefD1PYZKZU6bo7W6Q8Rsj58AEaLXLwoJ2bSDqgtrsxg+YzzwzIBv
9ygNihYAwnofcpZsM+bAP8q0St/+o4F/oJ5d087p4ULFI+Ql2LGaid6Z6Ogdh0aIulYIv+KAk7PR
zL5JJdx4KyGDx5FQUl5+4pJA8w8V94jDdtPadDv1n+YfKWyUE5EB/1vR071b3Wz+ZzkMmwVpw4p7
rLifcATUkauXLjkxXx6rxGMvRoXRe20lUrApzQP3DCJ5hda7mfvjmIPYo2zpXf/lzVfgItClEF63
7QqRNbx+Q6E0O9XRBv1AWQTBS+mhaozJnIFP615Rqz2uIkXOAPtVgqpptQnti+NrgPKAbdV50aLU
TR7P7hPIcMON5gDpgYTTOzLe6BOkXDHgoiBmC1i0FL5eE7GJyxNAJnMt/8boaV/AzOAUPfwpzlPk
Tgx+lmN5sfUcm2WCWSO7bsWkH1Y1Ux1ipYV1MN1Oyy2Z4lDTeg7ah8iSILfOCM5TP7WZdmOVYZlU
QaodxQP+obXK5wXlhyveZoHV+b4gI6a5hqQLG0CQmIgKfuS/ZKniyCKFn9oLQfqnAmc8kPQFOWTf
VbbokozMQ+CknV52iqMzghNQVnrIUu2ztjVe77DKwqytBEIBUw2OX8SrQiJIAbL5xAYIwh5LsJOx
OU5woNk1MWETB4f1DSFRebA84pN3vTRq/wokGcqt9py6HnpJlWiasg/B6HHiHdEPzqWI4WVBZmE1
1FqpcpImIMkTtirwQXNoj0q6o3HZbI0F4u3n7DrmlEB6TTcCYW4jqwABh3TXKrP3CLlzFSsa2eSN
tjakuxr0ikOgImX0k3iSk5Y80r/BNvfOtLV/yLMpddvUk+vqPBbixVD92vVoB8zfF+6eSafIXo7+
8IV2DpEUCN7sXCKrlcBAqe5p+2O9Vlp4iLE7ZJapYlHga99OkzCc4Gcl9GpU0cBLre3ztNLGm/my
Eqc3ogx1skJx0sqIdy/LN4Y1xSt+5CMVmFxAGmouO/f4w7qyNe9eUh58oF/Mnf10fcxMfOsAR0hR
G5bZKNE4yw/sciiqdLWL2Xi8qRSOPb6HTKwKJbOZcLMpsqfv29RNVCewWH1GN/xm+2y7IL/xlGkd
u/hYbDd+PaC1sTeFLcGrv/ZWeCUma8sfkMOO+mjasLEsDrAfSdbNn5S9nddSHoOrcDvItNkWSWm8
u4qWfCakZkzsPEGYbgqRYG591Vyn2GgI6Iv1qRJKHoNVH1MbrbQjJ0142aLq0XsjJZoqRYZjB7ms
lvsUI8sNwTffsAMSIY02qa7Vn6g7pPfmXNs6nRdoNwUtQDu22+UXbhVMFkxGuIMeEqrR45xv3sGb
0wL9YjNGvhL3RwX1eZRl+k3g+AL2JQ9eanT0r/oy6P9/PbgM760PBNQD+Dimi1YpcaglN8BT5BVj
161D7mgedkQHJIpzHoe7kxMSkTfRK2A0WOlV18uhXNsh3W1TNs9nBEUrD+LP30T+cIWeGlybOu78
2PFda1Lfy0TsQyJHfOqqS3iDxtRiuSm75FQzgDppGOLKvuZXEXSo5uGVNrjBYp3SQYk3fvhUoD6J
SIexJp69qY12wjWIYekKn072mFVkJBnZnHF5xDue9TI6TrOhw6+4Bkz4LiOmZC8y9yw6ziDY/m7M
kzU0HThcTvBSAJk22nVUsODOxRJpSUKFJUTXji1Z7mCEhR/6gf+p9J+vjtX4vk/MaojPfnK+pQqa
p6WPylslD1tTSKQcUeesp8jOMi2hzV/DJour/kTzJEl57mEXpK4GRb9GveLjkUKvQoAHf4+PSw+E
WvA+6C0VJkdDyGOclNo3Q8BjYqKHQYlFxcL+9UGxa3OuFr3Rcya02K4wcSQfgai6jkKHOYq5MkP4
sKN46JdUwBDFTnSsdIv1vns/BA/C5Tl3C+CpqWXLK5ryvJDATuvljk/JA3dd37+yRZJeTsyNqp5x
dHjffbp7Z9KD4ALxfns4cVJeegdcL4+FKG0lmOH2csFZ302v37cDMs5WevOdft1aIkBfa5zlV6p3
M5Ikb9X61f41EekS+0fElkPssjOI3uSha4pfZOr5J8UFEpUGgd3B1GDh8i315DW5mb5OrsW1M7/8
zoTMsAZQUbF9DShsp8v+ojRbQ931iZIxYEoB60KG/AErYi2STdpGjwDJRA/xD+0PClsq5BIvUoM+
DcyczNtRinO+qgyeLZBgMi4XxfFtR7bNTgZwvDVZCNmpVDshfmFivXzwOJ1p6Nvw4y+6HrJLdG0k
+d99Iz3O4kgbjDUzgIfomXnbkPGgyuUFg7AosGRUPTE2YpIc5Eain91CgoNbMlIV0w1UrGyVXYx0
RJXESWQB0dscdaMeK0RbtfKdRWNw10iO6HeIEkBBmp/r/AhFvutWYOEfDbWhnsG5GOldMv0x7vQE
ic5erp6SiX0O0TstYhujeUJAHeY670vKtAFp3GJCRbeKmM5Bwlle+etxA4RUZdp+7H8GcXT3PYM6
7akr4mwF+LPVtJO5FZ/3esw5vSH9JBGVuIujR0QE5tXlJhm3PthHFhFX44qN9SZYJqpiRCJHos4X
6yVssKbW+xzPUsbGICccbpp7S+tJYamd5091bhbE+wYOj+fdzojbW0FR7AHvu0N5pkV67Mbh4jGF
4mjAdDgs6Hl4JwcMse5DwSX86jqdx9rmO8+Sasp5ydqp6gSj9+hU34OdNhntwLv60ppdxBjSDhLl
KDEeMLWnxJK9yTmfjBAn93ZfoymZE2z9p019C0Bc7yyyf+3y6ToiYlDqiumL+qThS/knnCsfiXOX
WBrCq5pbV0xoX5kuFrfuMN/fv83GfOf2oGn6XsWDj3l/ezJFCind9TMwYPPyxt5IX2qE7kE1ATK4
O3GdcKkHhhB+G0E7av10BpCc9BEuizgTVVHk5saBBav9j/3dsnrynsHGwun0xWWEgX1+1cYTW1Nu
MSu5pmLODsZkvJopM3y7o+YzRJlQf7tiUFLWzRsXSY0VFyk6AIrXRQMPDiyp/H4dPKX1EmRTh361
Bb3QhehK1M487PsObkEWzShs8JKIAuNHk/tdDqmG3b6jX0iACo3A5iCYWCoGlrThYSOsbKRn3QLx
qRS6TVxPIsBH1UQ3EszQWcdnfvgFjmVYjsGyGAuFi10+FgjMocO86/FfZpW7WyzL6wfHmY42aPLr
cd6B/x7T43ky0Fa7sHqR063lPkI3WAmKnxl2vMoWgRO75aHapnMqed/tWpP+vUE9NZ0wHxhm+VRt
RfFDcKFdfdxMz6jxZDSV41zV62PcDepiiN6oOJkXoP6fZK3udNOMrpc/UXUWwwcztVnsKIziiin1
bKtsfcA8oUmrzDb/VOLqX69yD/eHJlF6auiLXfTMdxtXRsrXjqHkd23R90LfZ29o0cM5cC6iFhxV
Pz0B0RTaEjtipRZ1Mm4f6r2lZDfIEid3c/CTSyf4g26IUX2L//vc1mTqBGs+sEVEbWeNRlQ9Pgsn
EwZNRxaVZFFYeO6ZrQ2p6yrfq03hR7R5Ex5Wc/FmR21upflI2h+jefDVFJodZr74vNofRQOkdYYb
xJg/0doi39RRKTHE2NDImUFxm1Kinwvaqh8dpnamOsCqkfriVPwSItjsYQjspB7Wty3vFTaDPOax
Nyp+3zNObdxZ781Z3bDlIugjJs2brw1Roh1zeniHHwbh4V7/sM5TXcD8bUf28jvCm5bJsLnEHtLl
fa2HkHfVM03vloqkCuawD00EgeD9Caviyt5HiXjXn/WK2mWQo4bpn+n9y3rUN+exsjRIZ6B1C/HD
DUvcYhYUwgqxFtbtOiDB9LQDQEjp8SpHsqxmNCMXwbDf2yYi1KgUlQdUy42q2bOz2BjsMvEvMdSa
ei4KZhOwrMb37BG17j0KGdsH31DJNJvSFwRIox1JPkC6K6bIcKxWfaOwGRNabKDvubDFqvIRX59g
4pYOx1S5vFfqMrJ67BdCQWlW4s/j3j0kAsa4w8dUuOTMHu6sKf8EOXaLBzMVKXfVkfpe7rJ61rcR
dyeDWVHPwfL9VvdevSUq8djXFgCU8k2zTFKgoLZmQFgSgD1rPOZWIfrgMsZBOW0ymU3oa8JGBh7L
6qvHllSbFI+sWmAyE5Kr3Iw4QmKlmx3yg7fZi7VzE2V776i7mvrbSIXrZFcyL5ujpfc4lFtoE+Z7
9uRdj1qnewA8nxmw7m+KxAcsJi7SiZf2V9P4e6utXUraCCmJkTY3jrBZYXFS8BmWon75H7vutEyM
EDAp9y3vysUh8PSM1r7FZXw6eV749fyf9XE5sKIg506plRXXkqNd50BSJDitqts1aQ2lnSpLKMLb
SWw5mlQmAvygaN+XZEm8nwpL5JWDsnIdkJigR9TqEmd2O4TY2GUgCbNT40MxN79Ul/d2k4WLImF3
VsptG/iysKW2rCqxGLo0cFKjq3H8tJ45dhQDl76Adc819b1RUpr/s9wogSkcczRXdwlh03vaYavn
s1oBibfaLsRgmrPdgRwR4jPxm0WTYURAF4V8v3vW9ab62XjDNQUWxZhjqFayT03l17QbrJl6JABY
8Ky84iZvYcYyf4D0J51Y+1jCCkn6VmjKLNvpF+uADGWteV9wrGVCh8/2oPrU1XYObwz80ucxeCNE
POs48SLXk9BnVqZQYfZ6BqBUUfQZzKrhJCz+RImPS4mtiwycjTgB+bUZBnzXbVaUTKys/CNaFWG4
2LGZrL6vr4cllWwJgJvYGnnkOxwdcDUcCpeOmqBmAhWfC+KPoknno1RLmsvtmX3dGGN8wtvbN9vb
QrLplRHjt/03Vwqsjk/WM0mu09DPZmen/J8NiBW4WR+0XccZI8JMYypJ28emNX63cDyQO8y/RrJP
wUkJUC3zfvbSxd8OphZQU1PIcNzdL9IM3BBG/+vXYZnj00X1KrZ+y1WCEFuLfDTZOowbA+jcQF+Y
asSswUM7FE0XDMr+L2iu1X/T1JNxZ7BsUh2dCi4bqz2q0nTHYlX8SWLwH5+SJJm4YOLfmeC2xS0X
7HWGzxeXp9yT367/o9tCw+zs5svG8jrl5BNMAj+miU4Gb3NceVTeYphE5KoiPz/qWH4T0+Nqheb9
+p3krEz2f0I1yDUCOr9ANx0QrNsMpScOIjZ5g65VtwGZLstKcu25ck0w3JRnIchR5iRUCqnG+sv5
T8k7qUiI/i1NpZnjqasSFidZv4xcr8c1e+bCokFXK7CQnSe6TOyMcA0FwGbzvpa3VdxZM6Elq+gI
vPJV9S/2eXcT/SbMGbtjWHMUkLaCcTt74JL7nUU47d+74DyduPxyaqskko8ou5grv5ohvLxkp4C9
ZewsKP6W4tdFb/xUCtBhrqJaWrXpB6feCJpMIgtPR8+L+wZuOk5/WgGmgceo5dDEK16TUCSMl4in
9uNaekfLJX+xp8BzXozg5EStxBMfwNjutiCpr/WvPAF1s83CzTZ8+uZGQ4zmgSk0zUcG4Cw61XVj
efJ6nN2ZrNK2I+B45/PhDXcYlqKC5MR41SAWkMd+AfZX4Sqvi7Yd7dk6eMFVKS8duUiQl7S3FA1N
C1OzIkBheKUosWzZT4gIAdzSQseldiGkNfcX/87h6GSyGsrmMhnaaqvPCee9OTPN+aFnLFJ4pHl0
HTKybhqKh5b5ZRYJizL/P+MiuSFsNdevozYGY9OqDIJ3QVEhLXZBPwhZpe4q8cRBdxcj7euGCqPY
2UBxMcyRzFdH1+r4dOkMY7KM1Ci998ZytRvwiYsNQvOQiVpH9LBbUppnROjh8UV6R5ez24pLcG8z
rcves1lOhdgBU5SF1jRIeHAfZ3cjzYxXM2NgUiNjO1C4Deonjb8t613GgYDhDMrZgjQ6+fDRtdnw
TdPqt+UA5+dcYT5Y/RQqdR7eapKW2spX6Deku+m49ier6RdlZ5KnIi2/JsjUEX+r625djNNdhE4N
Gsv1sZvJVpuShsUcXbDjUoM4FS6M7c0vKi7IXHxJxtQnYpjUhGV7PUx2jcAeEbDJNpdZm7H7fGms
rKkm8zwMt0y2zSS5KmRbHLuwWTTaOS0789TSGey0187vX7G5B393quJUB4n+ZcZprMUv5BmkuubD
/MQtNU/iLDJcJi7+r+7qkOrp4QF/bTeIW+vaKYOraGz+xsU6sb5v/CajrvP6FJbVIN9D4VYA+pTk
SL61MCJ2LxuuZAdm8u/oUKBzTBPfPpRGGKds01tVoJkhEDIsse09GNERcF9Yu8qzulx5M+sHPV9L
GGv0HYfZXFHk2ygKTisaF7Y28eXFVJene2JnyoZYXZr7c2PcvIr+NeCb8Jny9JRPTz3cNBijLV/X
wzpKhO3sGbzeKYlrP9SQ9V8h7vzJMBrcfnpnFKSY0Vto95KA2Qmv1VG19UkosRycpOYpA3j0e91z
msrxSlbMECNHccMJAIS104pgH+vwEtuOGRnr3yKSz+7ZNfXclDz5VOqooT0WU5J6L+CmmpA13OaF
Zm6Onnt9d+bcNGYThID+uPZGR/eQvN6PeV6dU/I0PcAZsAMFt+FRKWevEpR8yKZDmWx0OjBH/Yeu
Cy2ZxhJbcrdJg9SsTJwmTPWbba6SMHDND1Mz6HqBV6SPA1DmmveROWRwNgcJo/hVzH1TT3P1ahhV
C59gY40e1yKbCerKgu9JH/8w37TDf7uBRoQEk5+xkHeg4iSVYB36TyTwdBTgEboqKyzLptKWAADT
QM88lbHo2r8zva4E0upYolIXTkyVqpbwUHaeQcgNb9wzHIHMkch6+w4DHxmSqAPAnVpS+eGF5ITn
+Fv+RpLBVPWdLhB9nMHEVefos124zzD2fMT2o9RPysmJxbu4mjrm58fSdKYq+Dej1uHMm1LxXjqp
UfNKMnj66eytEm9RXaKdyoKRnhWaspG7ra46Q+57e0MfpZAjlc4Sz6mNXK+8kGeQc9CokaJ4/pAV
uo9kyPZ9jpXW9vV8nUnsPG972UcQcvTHO3g+XeZDtX6Dto0SbnTvTeGoOcAy0kX108VVqB8L465u
kmoNehzX5LPY3sYf2gHSh/CAHPRDswx94oVn9elATnjFQ0UryUiewCFfjh6tKvR6GYGlleavKtJ1
FDirUCbtSMbUiBldUMpr2+ctBVv5TRQMqAwGWfvVRzLMuqyWDO8ab8earyFKVH7AGZ6TAaMo9c05
8UTOf6BnLWBgTcX5TSXpJTTCYIyYlz622/fFNLdM5z4WRjxfvhtf2KMZar/Ita8WQJQJat1WSrnc
taABfPo4CdEvND1ggTiV1wDudGMLkurnhjWKA+uPIDQhs9dqEapnVPaobLXiNbYnF3edmObzTOZt
7U+PiBeX+WlykctZdA4KqHjJMgZ5u9IfVVzhGl4T+06Crtr8Yeo48a44k4S0gq9Vre6xnf94a+Pe
RFRia6Ifm4BNI5rhqlipFJuM4uynIZJZmutB/y4LuJEeBM/fTW20asIR1zZEC5OugJwx3NkRQcBL
yuhMB66lzZp/Mo+A+SSr9p0Zz3ug1/1b1i68cSSudMfwqFa08xNdaoKb3f2hk1ZL5qMuE0OWheeL
RZes2IQT/eIlgWWb3kwo5sL+HcOI4hVoyLA3CEFihzH393VK4erJe7yMFfSoAgFUO6ibSLI9Ow8t
FP8VW/Ea1WwcEqB4/6D27YhnRogQZQoIEWH9qwNGT8WTAu/tgRljU4gfRkEvdcY8Mr7F/UHn+6ec
F3gb9uRA4zNTaNSvtkYhh2KY+4OoYs7QE1I7VxKOpjfkv0N6VlkNbxFpVYnuD3k2vnq2ghYr94IS
7dXiX6R3wL4Q72TDTWOs4rScGbH6zW8BRBefdN1NptGi8OYoGcwdz3XmUcwycXO7kxfjoOJeIWZN
CvN0I1PG9lvfTjC2T7kKhDRj2uaDtzbw+0O1eQLl+8FvshjqnTc/enjaoSleeS7oUqRRtpwlSIsJ
jUbNUVSwoRtdSkrL53dI8nhpLeGl10bRiufKXjk0YiJOGkdnAO0M7CwiRqJyeatLhatRQRc/BOuv
VXpgD9Zqw/wn2lg9zG9YVcht7UNbQxaw9H5UTuYWbrKgMhp2w/9bRX3gBilJzQigkGZJqDruS9lE
cl2YUUNlYFtYwRLAy1YZRNI+nCxO0K8SL0X2IdiRnYEa0BtH6ebl/Lm8EhaMDqVEta8RObUpU7lN
MEgtwN9Erp99W9lNU1jWKQCOJKDCnYTJNxlndfH9NfYx7XDJmxxInuUICYJThvyOpt2BUL+0HYqN
lHcwtvEoZ/XwiTCYBmtzNH9sgxFdUO6vK600jF3I/FwN9HP4PAySwb8CyozNtaqHOudqQZX8Z/Bm
JzqVr9bx7/xrRV3EaKd70jOwVGBJQ1R+WZPOdIOlcltd2DbRMB9DjyIi258BMYgga2Pn6Mm4vjV1
VDwA4ElR+0AOsu9jmgpM65d9fh8Lh2MIATPyzBsLgkiL9H71GpiPdyuK4DxGj6xGlq8hBNb+T6nB
3BCDiy6BBRfBloXRs9h4jM3dv0admIl+0gj+N//nTVapuJYZVWTwoeEilw5ypydqson54kEs0r5a
auVTQcDd3s/C/wCi5N5n+XQM2TNkT0RlD5frlsN9+DJwh8fezqxR58o0BEzWgBbB81u17hStN0g4
hH9B4QPXaWnukmu3ZLZK7vZlSFN1I7J/Yu18YVLzN4dgj8RtaEVp7nDuxdUJgCZNdJDGNNmw6D56
GaaIJdwAC3tupe886+CdVB3gRHV/47jv8w8tLmB5ltzhI+ofXEKPPrUp5V25ek48fSgYjbS5zi/l
Vr8k0/pbFRS1NQPjWOZJQ/yB4aIXLU2X0zQUPjyUj9LDn4haDMmIr+yG+8YqtsliZFUCFL+yBz9L
pEOiZ+gGhL/VTlrBZXosACqKEEW3UKibWoGFbJTrleJUim+lVpeqn5CIp+i3RjIJlRW7MA5LJ1BL
2UxRWhWSYgVtI29d8apXnqqqfKYgq377PtTlK4iPYZ+KxitIqGCbyqFJSExtrriEW/TAheEypzFL
MbSgj/rYvTSA/9yc2kZkIgdSD+vUarcWPFpZLluZGOvFkABW6jiq4gd5EAUcpUBFEMTq7DAgc7fd
zsH/j2jsfS7kseqxhHmGaoL0hQ0uC6sFNf5bkcave/+ML/gd4XBVXZG+Imn0LBUIepJ0ZzVJtXLY
wEsiMH4jlVAkBRk+mE9OzvN+oton+vTlWoymG7pXK+lLNQ6YTL3r6Fi/WO68guBvPj7CzLjp7kB7
Id/m8CZOMg9WfMaU9dMz9XfEVKGw9Vk/wTUwYpZapktguxJfVNQDhhj9ql7TA3ZaWPG8yqH1aVVq
PM8OzZL+VntsfNM4D0qGzG3n77DAgm5IxkjrdDpFifQxg4qA4ODr8wcKlrxX2FxwYMoeTSWao/q1
RoE6/uxu0kWA+1ElXZTdGiI8UJFdhDCYqr8lIrg8fqMIHXxe/nOPQ36WOdkLjNnYbpzJmCf+dtm0
Y713OiwTxl2LgPKRYPZzE4gAGOmadAWlenhKy6Frc0ieFBMkgb3xncOifk+BfyZw817t+ceVOvlH
SmIuoJEsvzqNY6uWl6IO1fPiG69RRmI+RipTJnSDJnlhm9RL1gz05r7e+Mrl/SyIPnm9cLrCHkLT
1vvqplPGl0SG+D+wVNkA9P4zSbwQ3sFKmqd3CgtkuV2VkJXT6fmFdscSghB++HRnXi8sZXOliWwf
Ulce7Uog6wAwIfdr4EIiBp6Gohr9ZuHFE3hYoR9IFZc2B08xnQkRgrlpsBp3dC+7Q7FbIrQQ9Hu3
UI/X2fLKuCgSnrUb1zpu0v7zu0eOLA/rf3bb8psNh/otUaFl6N3GRuxLqnqBxR39Gc/yKeWfhd/3
2DGEW9Y3n7hr1+NDeJe5apvKhicOvb6iTT1mo2q2DYsZOVoPP5N7yBZQsK29g+S0lhNJegafszZZ
xJx9v/+eJAgUlS/D05wVl72Iy8aNaVSSTuefAuLrvanLi0CBmp64r34cxjO8UAn9Rzj7/vsCggJ7
0EbuBJpaG/zFSQtd3mYMPNbQkxY2HGH3A3V0Y2pEBP/6X9IsDNf6TrEuqG/cW5xoFcJ0PSnODCMa
FFtM0mCHyj3HbUVnaq4L1QsWlePrLtBive1QbsYOH/cL7TLz5CvaY0NeKngu/qtiZb2jNtXCG46d
Y7isF6CSEYwjYqlQCPAQKpmlHTi1rWPcQDQkTyRMeOOzPhqZOJD6ywylKgl9mxe6fbCz0Fc/D61y
7dMy7a/iDkTleJY/HX2oQRhcj3iC7FcQQNy0PVT+rogEuZczS9MIGJrAFOHwy0k6DaM3Yf2egF93
QkqbEY5tGdbjd4Rd/zBKlZqC/Eb1VLgxhBH0YK+zc+VfbxZihMP/buXI2aIhjFX2zWF+jFy8euvh
f4eS/Kz3ILyx6tMc5P0JR4F3saawwP8hUd/tzIJoLzO0JoqeGh5gDl28Lu+J72fGIa80l1BOnWaH
gGc0JxouRj3F4y8M8GM9PgwsiVDHxpwtNvrYILCQsAMdf3MUrxRe5hiV4Px5bBQJzSMt2kcW6gx5
CH3xHrEmg7e8ig3rejrSjHYwdqpFO7nmGuojlHbAGKRdSqY8UuMSPOZzoEiG9jfrBQYtpqKtAPD3
pL8Nix+PscVK8YrY3rspCRw2Esc6ZvJkdHAv/KNShHxizQvGwC7iqgI9ISu6p09YSrkYzJMwybsU
t8ZESnaMPYl3DInUDP/OyXnghWDQkEsBdm3rpnDkfKLVyRz/fhqmMtQfWLUbdUQP0nX7ZwEcqTXC
Lrr+2IPfsuY4S59lcNrwuk6E42k19MyJ68vEUftMuwoOnt9UT0jMzd8R0ZjLGCt+Oi3RrF2F3pJC
zjfckrsfPX4f0e0c1J6Xj6dHw4snVUbwBIdUa62LdRvs5xO7gZaoF/mBotgH5QwX3tWZ4whxWoGj
PwFUHNuYGVmIA3bXPbdH6uSiqj8Pue4RnIHuYIdDi+hasLrr7DlDmogfoQ+1rBqduLsOwlxFHM3p
713X8s7yBGmX4CvwckAbzCphiGR1UeWx0gC3iQ5H0TwK+sRBv6iV15xCQVE3sRteUCuQ2qWtn/SU
sZvHQuyX6JgI6F67YTvo5rO1B3egMNAXvEIZdCypKY+HCXDYJ9GcaaTqnDj29+lP5122Ay0dcLFw
MtcRxP6NyvOcRzskJVhzfQJF1VG45i9xiplA6hxxYhI4Miqhs/Aihlyj7HI2dwygyTD4sT2MiqlX
xVzcAitBtekP/hAuslxXOMYad7lZ792Akrzna7Tcn57v46AgZrnhs5GgZbqKGVOwDysaVZMaFbwt
g/K2IVJezG0tNAMlu0/YNeoqL8CRNoW/6hMStYcuMSVM8WDIQ+ACWifcIc/4xEUa58JryV0qqmJx
OiD1a6Btfv97sbuzZSvWY8XaA4m/WNV1k9zI7mRzO4h9kO97z+dpYTJlZgrbAC6laTZ7kGrS5fmG
4cwCL8Gj9MjaWNdt+AhYq6Ab49kJ7L8lEES2P/YLLISrlO5oRc4B0QDucqdd/fZFnYJBr9/a038F
UTn5rSdjXVhxaNpw/CaW4UtbDWPXvD2NIExJB5p5OR+DKrHyBL2iAcS7nIWtEHhXffpd1WKgOKiO
Cym/aCrZJmNp021ZPKc9GCSIZZBqqbqjjdCUAh+Fa/l4zGbwv7CL1EarwtdtPVuKnIBwlYUg7br1
CtFWRIALL7iWIfx83FmuaVA6xwarKZfqquRl5RSrv0H/3IdGAVJFsF1RHNBOsppiHbfQJgfM+3RH
6//Iw1CX4B+B08CWC4XnNijcRad/1YIWMQE4RuCnfj0j4R6a8KAB8wDlDaIyQBuhxwAIZcW455AV
gp1RGCzCu8PPY6DyZzD+u9zmaynWz3wuCVs2IT6ia/aIr/H+HZ3FYwxaKoHOVQ5ipNIg4mVljPV7
ZwSOlqjxm1PMxGXtQTn8J5f2WNbDxRMZKNrQc4Zz5D4vEhoZ74yhMI+6ZvhOLFr/GxUnFO/6eone
QWhqJ5Nayn3BRLzq5ApizruOxVAyQyMQSn0OnJqktndFHtBz02i9Oaypz4Wi6tWpT153abie36fV
L7ecrWmdyJy73gHMURQQhgH/DXRuQTn8HwIHMUQ4vamyigrsnU+cxBWMlUKTfgPttZIBqc0EQO8U
KVC7gUImr//AZCBHm987ehzeTYHuJxKDut7ecD8O1YCd3DOLq/hVZdDVlJuAKoC2A6S0htO4QYIV
OxZS6cgbS5ZR2dhcJlZtrbYfAOsOipa4KWPlVRF6PEjp9ezZXldXY2p81xXkE3uJMnw9nBnR2QEu
AvZzNwPqdVQIZIdj54a+hoisiuGsa5OOEK1L0pZ3K113hgwMmql+gGjnDCUUPxtjJKQiu5onvFsh
ZoRsfAeZzNnoV9CR2U1L9VW7uRgOdPBKxfOxN7ELs55Uh7vl67THi7bIhoTk2ZlDMNgaIVielt9O
aTqRXAO0w6obiqARtJewrWXrVu0IUAEtPXfnzwFyOrILXwYY/9ahqrFskI3oEFIDj6AU8hkyM4Lu
tU0G1oOJgGETtSqSNmlBpxxylrDdUvd5769V8BZ84lj75++HGj+jTtm9XQINZhubksvJ9KiPTT09
hNqzXCMlgBRgOpY9QTvqY3jogN7eCtT5gt975CL1V5nF+MgfRM15Yhj98pJbqYvKV97uXhDTo/ss
BnjNMfsa1exGgP1ikCMLScBlSd3lUT3upMoJew4ApFyl+Oze//HcVVxXoorhiYgYdGC8UMxjKFk6
tkuPSOs/k2HwH8iE0Yn8brW33fZSiiqVq3mMD+pa3PYrskum+cFVt/uqyS4NQizo3gO1csy1Y5TZ
07sv9ajdfvkBoCLiXVR1OG3dRXcy6Ga2RjaylEV9EWqxW+kbCgVddWv369syzELE/EtiiWtUFEdj
3Oo6bqJtANgugp7/abGLooa1unXiP1hAGYt35jNAdaWrq3aOKnBu0qNUUp2/XvRLrYEOvXxf+zmw
2GfDCLMcwFAU0GBLOKOAcGt4tiCHBvnw+K5qVdZWk7zoCcjcVyxs3SaeZnYMts8PmLFlf9uGgz5G
cPnNFFmdDDu/rFNtKQkRO9iS2kXcNa5+yo104H6RD67fBq+gmAocsn+NlPr/dzfMaLnJ6aPH3cTr
WHzGLo7GIy21zkvxA303yDuTm5S/zC136jflOCiiMHhFNfXy3SOko7cmvFb6/0TjH62PF5QM7rUP
RHr3gEV1apbI/NCpWAh0hBIR10JhRubOz03yFvdDAYY2KKdLinFa3uJeTXcGLR32Py+Cg5faekgN
5m5RKUcwcF/bB0kTQ3AkdJo1VFxUnFNnrvYIeV3HjjINDoZSvxp59831zZUMDMZF204BK09EsYWG
5SaZwa5UnJ3OyRMBAqDdH0uS2cD/GOOzDXYJk5qmZ532qxN9kim0dpUCITyO5LoXja1x+iouUtWp
v+tFZ/JzJYqcSf6AN7lVv5QdA3+ww5fbz5vXUIRKmvVN3KgeqmvXe/WNvZjr9vgOHod65J+lw4PM
mveIP+tS72f7iSkfEkSl0AsMDOd1kr41zXLfT1UHCjw7TlClkkyiw9Cht1aI1PRGzGx3YCb2BI6X
2aq82icSdN3UpqI8y+YMy/UxZNwUKkIm3ze4Bc/QoZeyxnZ0qCdEt0t/7nuE+IFvs8+KcpsCo4Tu
RNOksafsLe55Xf9wVyDf5SydV/Mq7KtBDAeTr4JrKJUPP7oocqtELfYrXP/kDl3PPZ87lx7vHdRw
HMdLdzyRvuwt2ds90wgbxFbmoDBT8/C7lDyifhJ7qFRweYB1t9MzFWMB++pksaqL0ItAuPw4JCCp
XN6btZmbDMLCKitRgznp3jMECjRI5nYdPF7Q7k3PRa2tyTo3cXQWDXQedtyMW55SrVGqh9ZJlsKr
RMWdwo/WrFLk0yDF33I6IC+3fDlzgl7XzG4mwG4GQUWKbfuhAPhKWc2KfxKTv/3e4q8bDBV5gx3p
dSvMbJfcKDMp0xy8ptsagcPD6ym94A4dVnliKYbAQm6qbJVwEyocwKwqUcTS5k3Fs1QKbMlVKgFn
QKPxw5gY/PiLBsyQCI/DVEg7amos7nETgrQ2V11IAgDKhYBQ0zNt2C9eQbVzFcfyFqKwy/fH0tLw
XscmWwT2nVy3PyPtxaLgxzVrW2ivNPI1s+ZtaVxbisVe6/2YbRXINwpcbdVGZPKXV7kz0LnsSt3O
oHrTJLzW7EHSQOG4c38O3asOB31Zt+Les22sC7zC+FIoIs9XRrdM9uuJ+Hgoec+FxGYVdASRlOMi
Q6G3LEngmNtg/cUZhpeoqEwN3VTVE22lg9KLNo+4695Q5ODUsOfbt6II+Xn2Oiad20hmve1JhbvK
cBNpKCk7WwqHmqS2b7jxyvw4bOd31EO8uv7OaKlq5UHuklL4S7IOeZAEs3ivjMyxtwwtRtBC2VbW
P8mFboT4HUmfRtXSSVw6lwBLYOnxebqxgjoY++Ci6JIu62dyGP+EJysiWsCDbu6qkukLMHscBUfF
XeltYU7eRMB8RSciXLs218kVK09YAO65bOJJw0gz4qNtozO+FNcRDTNMIVJp+aW/7nkuz6TBKdHt
yvKaN/y2oPZGp3umejJ9XWpLe6bAkp+xV5Erpo7FWG6vnfMQeBqjpyYKfH1TH0encG+2VNCCFUeI
a9Bclql8azldXWzRJrdsd00wXM//z1xteAsd+P3KCVFaNsEhUXpITsInFQ7NwuJKR5Vka3hKUyu6
GCxSCLAw25U9TucnaTEjLMXVdG1sXI31DfynGpvOf9qIwetD6fB0yNXVlzM/a1Q62tMpXE8eRLnq
hvfdqKO9jsFbnTAHCvOxcaz2v7DXNDY502gGgJYnJjPCcYVIi2Ko4WJDOakmSpyHQW5HdolUdmV1
xBhX1C9A9SehzXZSqRp6Uivkfxvi4VEyR5LG8DoBlPgBoa6MaOcSG46KdyRys08u47FO8wSdGNGL
N+cfPHser+C7Of5qqEzBmAAW197ezF/IQjt2VcNVwevyn74SZ8jPDkeo/qo59hBCNIsuWzvJtW6s
VKbOzy8adlRvb9OSvM520Ep8JexLenSY9l1x5tURwAJ+4AFxJEe6U8hD8u0LDRS9lovFOeAwXiEZ
Tq/vffql1wqpAlawC3BKbRS9EeG1wgZTpBEFygfAxLy6eWHxOljPPMueLW2WFn9z5DlFA7qawu++
wd/4L+ROsya0Qzb3DDjthy85/tngAauEHsmH4Km7hwd93Joza1C2Z8LE74KQyqkpeqP1LwM/oD+m
ZHUPgiHpTD8WTm2FKLbx8oL2Tz5FIOGk8fHRjcYDyZeCW6b2BJ3xWBVOFjY+dQbbOJt1XBH8whPX
CkPgBAdK9fuBZI+5RFzEsAMfsDeqHFxblp+KJ6kR2yjngbKpVwQDm+Z09YyDCZ1QGJu45oUq5soe
2nXpsYVOfdvjULYGy8FlOv6AF3P/TiiDp+penbkeR4zNnQSyA5hExO4E/51sK/cHTLSPELcB/SbZ
dbYwmtHQLTIMtWML5NC6s5rlNfBIhHTys5mpuiFgvff+f1DFrpwRnAh93wydPWDzrK6lVZNiYXm7
l/Ebry5CdkcjcFzkqzGbWtgn3Jfa59I0nsLsnIU07DZSFRFQAixvrL4pGjL+5GPs5EQTZUvm28xA
EsERIkoaag08eIHvbeowxj6wmG6VktzQmH5zL4wgQbOTt0sawk8brn7lvwgb+Pc1Qrx37W7zjCJj
7fSrFPBFQfO0Luk6VhWz7KhX9y3Hyau8YQDZ9BK/U0jZRFyH9suwQIAAQS7ST45dTTWlau9ABAdc
D0BsNuH68imel25UJmuLe3U5iBKUJAxZ02/FW8LXAZJyRxn+I5NdUCFwiEOVwVykdIWhugb2Bjcv
SHc/YACtZv7KCNoevmKJWzu2hGnZ4vI544KxMFoETuRMqaj/990fUlTU3oBFeSCAMTNBpFrqMrWj
atUKGUYsRnpBHMLa8PhymTw1mhAZly4r7vAUPoE2G1q3EdG6u3roi6bwR+pJrzmfTAJXKPQ2Sz4L
eDfFB0VXbKy6BLcfHtfxkdG8GM9h8fMhQNGMVFN/c3mPTpcQC5Yn2XxDiao7F0JYDTibXDFD3zmv
xMfOfM3/OF8jyePjziysKdbwqUyGJZ5GsCdhl4E0ZYsnJOqSawZzEOIN+lGYNYVZCSYK/kHq3Oma
tmPbYfzneyTHs5NLDy2yy1EW9nYjCB9jFCjzMjbueMMAErw+uR8NitfzZBxU4TzScDVJbZdGk+Fi
IES5c2YTz5PAU3g8lQdo9IjmqN6LxM8zUt4oxkn+xjokGpsF/CNM4MKhXBBTGTr0xY2OO3L2b/pD
iLgTvbVA5IvHCGfRzfa+O/HXavOh7XzYfdYUc4fzUAKQ0POfgO4e2OZrhLPX7nEVepB5c6vD6ggU
56DrW2TSKYbbtxHejrvApVbQizgc2rzfgywaesPDPIhOzG3Domyx7LPMX2BwDyEjGyPDorgwAjyB
fASmX2BnAndxg+RVI7AcrsY5hFIu1AzuGSJyu42ckzE0qexGoPIy9e9khNy725xM5IxV7xRSkzRy
P9zQ3Rix6BpSOV9Ngc2fUte27PX7lgL3X1CIpA6IY/M9GyPaCHwAeTuJq/Yo2KdnoDBqHIT+/hxb
B8tNK3IowYUPjbqrr3WUGIYdGl4dq0P5sZTv0XeBdb5eqvWk4of999eXJRVUmCIfgJg9E4NKWVJ2
5PsXq0xgmz862Ptcw2izDO+qEjXPGXdbpEPU55tTS1TspVMbm0QfUG2If8/70A1xKsZfQnYXL5XI
Me2kTkH4DTQwix9RoUomQalnOSbrh+o8D2QIUD73Vd6+T5fkKn0KdqBESE5aBJ9Ln8Leows7upm9
QnOStJAaYO/Fmip+LXIw0DmKw0CcqLcxGt6EuL+GfZ3obXw45ALb/2ZJSQp9KcVYE/03JxvFjwF4
BSg3txBS/lFZjILFL++TUisLnwBckHhmuvrRicq6hNOzJuZLOySbwvxDgj/cdePUNVfKe4vEKv4c
3ryq2IkBVYqxg7foLdSmJuNUe8aQZYUTIJc3TzUUgo0O6hMYLMnEbB04ocA0qSCh99mvbrNNrpG+
ORDK+gaJw2hmK6aakH73jT7nGWuztvhjuwBPN5zvAadzDOyg1eIco4Lggy6wRQSlstbt1JX/wOA+
YguQgSDrKLFW5J+mqTsz+y56M/rba0BGyELjM+HGHcjJ3PorOToBDzdZ1wYh9MUbmBNdbQ6kXOtK
rO9Q/cleW5iZgRb6mFm/PZgRzH3fucsSAB/nV131bceYwDEMMHmnv4h/XeN21b5vwe+PMsR+4qxO
0vlwT3ZiL7ktGrulekLwjCfkk2l2V5ZgpN6Hfbaqey+cjM1AOofi8Fh8nziSW64alZcQldopL38l
XvdBpt+H2WvaM3A8IARSrJ21AjNDSH3MyuOLkooacX5Hhff+zfdTib7aQqFUqBXlpjEk1ZB/MQyj
dJKI5ImBazvyNYN10WGBXjVO5UnVlUKdNXXsYSm1Nog8btayY/+hklEgOC8ejYYQqW+tifhS7GxT
xVy6Fo1NAPsPSfQg9Ku8EEqjJdnIVIg/KQ6QgLqBS0udqKEnC7w1Uxx/8nj8vUE9QRqRvypcOlCz
E9dtj7/HeZMFIQIeX2aNpDcS9qdfaz3g5CdVwrNwAKuDUj9YxN6/gqdYQc2+y8uiUA8IZ22vVJ2c
w2Q/gE6Nzgw2RC9iK9mBXptJ0hpP9hsv0YCmSXW3U5RTFLpDMTEPtDVs7+KvKj8F16gTDzMuJjDy
hJnjzBaRdHoV5jpbighfnbUM3p81e5khoWdGk2DkKeIt+oYGR6qcywC//4IBigF7JVH+ICvfm98Y
nKnS/ltUpSqs91oa5GDn5sSWW0x7GLvyrxAi4DR8R4xEytFRp0jF4hBK2cR6C8ActFuv/Q0UGakZ
8kil+U39QDT0qN781JBWVtxnY/FcYI3lHZTgI4LrDUW7VVYB+zsEKD+vmOLxJ8TK25swtUad+Ze8
OvF3mGZUSf+YL4Ar7hk2o7VDCMZXK+/VWesdssr+7fTPYaN+DEmrecUc5iWHRkovX/7FoYpNDvsA
kir1lNydkeRuHZpFFeteAJgm/wadCTclvAvZOATc+YpyQ363p1rPbkKsIb6+Y2KA/1bwsQlJngfB
S189MQ2cswYor5OEWDIzFj6xor4mP4HAd7/MVc5CputTtBT/u2iUGRLZ1aT8La8BtUQX7YU+Zg7c
fEc+R3Qs2qlutaT45i88faxFnEI0f1wJxIH1GUCi1NVeWt9/wbG3ol9u9fyvrWoUoJ44SMhelrFi
kjGQR76d5yagPBC922EJAHM25p0EK4inFVrYEXsPnMxzLtBWSd3aCDzgpf5mYwNzk/ai9G2OrMZd
9X9ofsLIPEYBRp2+5BWPbBKoIUvr7oVzyOZRjf1aK01msKYDGQVI304WaddHoIRNbWzqiVRa8j2Y
faVPqxfdgh+9CBvJT4fn34SyNt4a+QTWIaxkj7KL1RwMnDK0j/HvCTHV2h3OrpotdMi/unzR0Or0
/ZA59EpZxCFGMvTwQMmSMjSqRAZYDVx8V8rglr9IJgZ+etdzHTV7rpePU3toTrg744YbMsFCUr/i
22M8NLaosDrgVpW6Ummb0foAySaxLge3xfelsbAjw+L7TW6XJGCveMOh79NCXOMwK2mGsem8zZAa
x+gCvrsL7ezCLbMLnS5OsFdsw4+Rs7poghjNFhhGwWxjSTH3XePPNSPv0GRfUZSoPidCeCeozFYl
29Pv3ko+dWvNswoZ+WaHm1LaC6vlvKRFDt4NqWL2E7cr1xk8VHC6o1hRsS32bKWqP3NafFaPYAZU
I2+RTg0gg3scAuyOtBJYW0717clOomWGudQMh5x4OS0MMNvs3Ld6olrNUoh4aBxQZn2MOztKmr4x
xRwzoxH7enr6C2rBwM9ZGvszTvcTZ2q2t1UeJj/2tCAGc2xQQQiGKWSKg0C9ZmI11IBrkMEwU3sI
mdMY6BFndeGHnr4YjAllxZxD9EMTha4JvLu8hQGKYf7l31KYZj4bKv8HoE+1hBawQqHK7bDReOMv
F39dPbPxtmBYsiC5Jrtem+aGIPsERnS//FixFjxUNo1a2mrIuKdh96uTRk5jnhFbzagENUP4aY46
4KAP1pS1k5E2LkT6QPnyzEFahrRAcWo1lRQB4YO3SE1SfV6RjwmmZY8ppv2mAIwLG9+eBCkcgF3e
5orciw22rP/Ic7FpDQnGB9qRc9TbToQNKmLnEL6UxWMfkg2YoC8VIgJGZnycxSx3wI36kQ8z45AW
qW9gvqFiC6nqbKW23m5WuLlYWK0vPYG1uKjD9X/kb3+ckVH3XrnjGchb1AeOF034mtFg5QLohS5W
T0ceoEFnQFtgj/4vyysfa2ZRra86tFNTBa8Ir9QQw1tsC2hvM1a5McyOmRRSHS2Ldkc15KKmx+i6
Hf9Nl+2aIp+9BKXHzjV9Kvgh0DTHo5qeo1aF/J5L1A8OnSSXmODKzPvZGSG7zrU3WPo3CJ5YW1p/
lBP896rL9idPQmFq8WqJ3/PawcAuywUpO6jv7DZXQDE3Na1/elkhpKHD0wkPiy/kyVXLzO9Z5LC+
fzhAvFicYm+QzA9833qRr2L02uxTqqaEcsKm8zbpjtQ/axX1/v+LeTFw1GfzQ1TNbe4jhq/VG2ba
VhkWRy0En37MxaG16p/872RaDyoo4uE9d9JFWl6+gB0sG7tz6iYBjmTKLeBrkrU4kZd+dUKv9r7k
cfURwp1aWF3GiMRKvJa/ZH09SVGCRBDw1uxxsJdsyoLunor6E4yID/OnamsnYjCfkmjM5j2IfK8+
nzpu1cePBrX+aqQEXcS15Xf3QCBEEDZMLEul9Wh0vrQC7EtJLsOpTJ0QgwlszxC9V0031HVUnLAi
mvRqphgRRaiCdsRmtfppJTY24zmsKhBX8F3a3W+c800V4t89q0Viw/MRa+rn3y2PlH1FEKCXAG30
/siWA3J2xI1ElNwJigPsx7gW2PmRvQiCPEsZf6gH4OvF/QNw/Px0qwdy5kG8nAQQG/xGegL3k5ro
uxdlOwhkyerxU/+O08Qv6uWFtjIg00Nv35QTrL6gESN2Fzp8oEElCncaIyG/QH1L54PSZ0JzSLOC
U2ugzgz/nnt5dan60zWPfxos436RFnj+b4kb63PyntH7MKu3/K/JihSXLbn9uPKj14WtRaQZNfrI
OmbDa4te1fbHjP6Ei9f8ed6ktFA3/3se7HPIuBSSmVeY99gB6IUvrfi7ygr9pjFmuRGNlXEgR2tx
Ily1O+8TYpgxkZqEiVy/OGjAjFweB538YGE2RbQZoBCAAYYtOzxk7m0uPC13MHSRxHm//vETS5Yv
4mlLY9OzZTrFgc4n+ZAGDrg59QEFTYoRYcKJYySxlO/LNDFMD+aSQDx6M+Qs6R4XgCG74EUD5HMz
Mt4i5tEGnN8O9eTBNZ3QdxBfjHNUT/h0Z+RfS65La/w+ehl/gYtw1YxGLIMiGZ8QlybaaBEO8Wog
f+b0Gkj4WNe23F8L21iHRvxtL0hNonWotaMFrqjF5SGlv7OllsMaQhUk+JPDeyqer1okGKJQ4ITh
DTOF0EsEhwRYMiT2ZIQuNWKaLKwUR7VEzVlq79wYNIa2CuuGINZs95i0S8L2HgYuPp8DuXdZVtYZ
5r0jcZQA1g+jbRGMO1pIm6I/aBBZg18FrS8nFzaGxP4CljobEWCt+K/eAAE41OCfwSo7mbaSwboP
wd2CH9kotCqynAUHjhukmNzjwBeU+01xQtJ96CwDQR3Ng7QU6tCBuxaPnqCvqkj8MqVa3H3BaGzQ
WcI/MKpDOuFVLvwMxfg2QYQmjzwJXr91nZwA22gLIz/HDVTQd3A+UQgMxJqtWeGvd6IuuQRCwAhe
XEy7gTQMnW+uNldzvxjpIEL9KzuT4tmN+3ghhIQZ7s0WEHv8PeYMphptMP2KhTZ4DPdqWc/R5WaL
glpLrFt1T2A3o4oKtF1+BEMWlmrJO1EWwp6Ixda8KdCCbkmK33n7xkIAxPPlBAStp9rRBR5GooUY
D1tntVR4h62KLeVnOt3zBKruA2ZkdAEI0U/cQbOunGCEp+MZcL2CjuRYkJAZTLS08fKkub3wRPOh
pzcDhrVrp4/Qturv9r6GxWrHuO39DBbemfptY4G1hRBhwHqsJrUERXHRMLuuWYAD2exqzIZhinOq
wveJpOtqTiaewI9rDmyO2sSBRyYpAHniKPtczHB4e4vG5nbLRfFYDjoQDoHYpc6eiSG73IMgdGSS
UHyg3Dn+P+f4epFe9aXBUH0eupRO1QdjLMA3ucdCrrwzfuvU2Q6zc/rvCQMWzoPbpL8RmU1vP1sz
4QN7fxz/QA7GTy4iz60nnSOncRDQijx9F4H67l2FX8yvyKkpWXtJ3BveIQcBaWCvNSBFZboWBFxA
MCzZl+gBOTD90VY7/VxX1m2TDG181M9SENhuwqVlNGAA2myaJN8z8TNqrvr4kvDtLKaCLqP3FoSJ
180zB0b2VD8bI84fX2Zt8O6AaltgFN9ffTlyzsH6O5gFijKjVvNt6Js6rTGjBY/pmGKYtTyptxI8
4xIOgo48gdEQ3Zbds4MM30fD20GiG35Fvm+I1l5SjQZvvt9hkpYC9KHDQEfCMCh4pmF045ZSNnOn
uw148YEukGpoSLN+iTwcmeFG1qA/AKirYFdy/obnhOBN1PrxoG7cB2xIE53so5kjWtim519247oo
LpMCHZe+//9MEFK7fWfTU1zpN744LG9bV09GOyvDfYE746U9JRz0bfVPmE95ZrIJ8o6f4oBTW1m6
Yb22s2BmZv1ub4C2MoVIqS1dhttoOm9kXFYNgKqF6ZWZBW6InT/+YsNez65ccNSR5yXJ+JBCX+kD
qpeSmC8O99h0hzWHQalaIbNWIncY5gtZCWnuEQpGl5sjJhKdF7AUlYP2LdjmOjxOn4X+dZ9YUuIk
pNxKCLY7S0wtaDIG0CXEBKshauLgDRMkD9dfCZ1SUSQEWIizLFXsYWQVOasRhhfCgh/TLwIilAcr
rZ599Wlll/hAWaKL1NngmWZKqqXeeTsZsj77L6gCTtwpwoHandLt7kICepKRsP6+R+gkKlq3iL/Z
dm0DkcI91W18JmdW6WlHbytZPN1LhcUW4hbHdFjHfCmgIa3QElNQDhdZCrTGbYaykBOBAmYzMWxl
VsjRSWQ1RXKOdMk9rSxprepw7uvQsYX1egq+9GELDXhu53/XqQ6jhSPqGwFlXI0/PQkTUXlmnnWV
zTMA4KJtmRiG8Atqy1oc6NyxAtXAElL0Tmx6xnz1xkOvXlDOLil2xpHS3oDKPnqFbMO+TqoyGcyu
na2JciOB13TqJqmxdiY3as/QlHJYvz5GIwqUvnbx7W93nILnZCREe/JbkQ7mcoPSnJi3XOo/By0Z
m9WSJ5CviwZAp5O24s6E/ZfzRjlWCWm5fMVbjCDXhKXkwxo3Tz8VISJ+frj+d0yhRdlS9TDalyN1
PhN8hbo1MT/W/OI8O+5GDf0D0VMsFVM3KIrwhKAl5jawrdQr1nIW1IaheM2sJ1kOKKAmD3qnS+i/
6XM7E4KeHvR+mEbsVMV3BR8OVf3fE5YhTJvx0z2zEvqJyBIB6JLfJDUKjkBO3sUuSgAxJCTO+vPU
VnQ5+uITgZdwmWeDiCkGjnUr0l/GOJxFjB0HNuSJy8LhvJLXLbmHaYnoO2Bm/Dl7gQh1fJbtImr+
qUydGs070OI2mcZiSYHlXdlPkfFUUMSsTKxRqwnXwZTcDDEEwEqojuqJpyERdecVEB4i3cNa9x3Q
O8nxpNJ48QPDXdmVPnRZTPY59T17MZICfg9WwVZoNMx2mQ8/S5SWRjYhOfv+vUmzd2ZvREgupM8y
tMzP0xIvSVULEsVAvx06YfrPneAIYPw/klbwUJJKouQDmCeenVWXnKCshIThsDs8uvgOJbvdpv6f
cDsMSFKOaCxXt8HCahioL6EBTRqudeHssoFxm7G5XXqPtqa12UsXlY1PRUPL5meGKFroB8oET2/L
1byBFywebnmP3Kz5O7s9zkuJUJ3rq9xojU2rok6Lu8fHNleV+dWyBxb3+q741W9y++bdiV6iZMgy
OCs4HKYC1mKcLTpsWjIesSulmpxXwRMZqLbSx0LVgJO9T3xp1thMVmhvIwCDDs8urym8usVR6g8F
os1z5P56nEHIe1JrKX2YeKRPH1G2DBSA36qVQl4TrMOSBqWDa56Q51aousflge3MRkVem5/+CWmz
tQQuN4lMJNBigFsfpeRzHkAHQqtzkj4QRECCbf5e3S1YOdgjVI6CWRbX9QR3+a9nAq6K9Q98Fs30
zJUnHXZWsq/6cB9nkvWPN3Zktgj5mmO3tMA+ELjk9Th/eSjvMG2BGBFfGgMYOmZK02WOpv+ki4+l
Blm5R4dxBvllmDCLnZJCcD/Ov9VTqR3kfTDoMFuVB2i6heZ7r51S5rlf59lynmlskjnsId8VS58h
vtsUx3BK0jNnDmrRZPX7cIiYNGhtGmMZcFhUJ6iT1qRjxBEj1WsfnY7T4TFaLkWevLnts1BkfuLQ
w7IFU2KFag2rSyDtlGxWucOIPCkgzgzTDzId4lejsq/fZnANiC5/+cCiAOpnwO/PT50c3hyDppZO
gpttjQNv/AN/UGXNsgkpyWDgxVMLeNZLsNDuBxEjyl28b2lY5Q76/so+4kFdFOJVymfnmQ1pTp5M
Qd1iv3Wms3VrChQ7j1bNPislLWVrJbFKcsz1/303aIr3dYhkt5z5BrRzN1U5HTLFsQc/Efpvbk9A
ZryNKoEruajKc8lYv9Dh/oxrfhvrmL/7jZmZ0Zb8pC1V88a/Sm+CiTU10k8Kq4oPr3k9UIU0o5KB
ThRWCXWvpVCn/YB9GPBis8/eXwRpm9fe61efMNlyqe2C7uqFnncQcBs89WuQEDMHhckYStVb9sSm
b/qoio1/Gof437g7eqR+v8MPfxKOoYL9TJA9GADXSGJbyP0G2TQybkZXKGDh4XCdySYLG7LBYhne
m9vG738dv5F7nUzr6VKBNQQ2IWo7uE+iA0c4phpNYueWiQEqNOn6Dd9jB274bO68zW/88UbJ2mZ7
OdUDXGNwm6A410tTaCcSvgv6JOTpKj9i7ZPSQ1SIdErLqbxXfz81F1SwoDgbetId6ps/g7xgG3Ka
4YRllrZXwWcQyLpAWpPyC2M+NlzjoLeMNb4joeVqOh3GHjhF2uJ1C/YqGILTho/X5t6bGRUP045k
Rw2Dnz72b11rbYgQQAY50/++7MMeuhBUPb3I5frSDlsbrnQVVvcu2/WK5uoRviKD/g5omyLAaRMK
pFHToRasCzBaWMAwcHu3jYaOLJ1SadBrTaLOSadZug+GzBChjUMU8SWoYVBiUH6HHuYWrZtscTIS
Go2XvwUV4+Yi7Tf+f0nraABfOKF1Qbj9qyXC/3fZbfokDdzh9xADcPzgKJ5PuC5jBcV+pYbNkM6K
/nuuxJUxY82RaAw9GFxFduBZ8IUF0QGWWYJ+ixyDa7NqMFkDtsOvygdFlB1EiXdvkO6NpOkdt/HV
Gh2qhtWFKuiKvYf1atcA6T+5UrXxUwgvhyx7LaxtE9lM44wsK7p2CXUiOV1gwSdt0XgxdR/81E5M
ZKFzexeo6LEcQQVgkQpJiNgs5Nv2TKEkS+cji175kIZF/seNeNAhMVrsVmfOpSycgN7IdazD57hL
ZiWMpZa3S4ZMho/uZZ+h/aCO6pexLgoULFkt/SEWxZA9yHQq9jJQt67OoYS767G3kF5CRSeLweJ1
WbFqQ0+z1aVYN1W+ykzwZ4gcNX4aQuJ+Q0NsUjmKMeYDG0zSxyi1ier3qo4fjfoc/BIYWeWa62nl
bLyLUV14Nt3Cl/N6NV2qOhoZ/lfi/oDK13WshUFUqfiyl2jVhveF71AZcaaKLaejH4etCbW/FNWD
OcwPpOtVX/YfteYWfstdxWPk2EeV4KQZg7/dpSjGB1w7pRotjbOjPv2A8TV3vEmyQbXhfw5PUTOT
4aEHCbvsOvhemBcRe+YJHtlx6HT/now8JSiz6F0XcQ2uBYlr64FKYl37Wagp5bAAajynAMuXFml6
ak6jfadCsrvYvd1SqdvbUEfd3nYUPkU9JIlSWmFSMTOJcpqg4S443grdezgH1l7u2ACPbrqMo9wN
RIBV9iDbDMoBP7Ujsk/6z1Z3nYBECBxGjmHYVp+ZrVRbj81Y54+tpXO8xfhAlUsL7LzA3rZ7YgM7
YYa88svNUtfrSYYVg0SzKMwf3Ii/mu9V4mbHPNYCvDLceOAsrTVHN6izbbmWOLIJepnzQk56K8PG
/nK/r/nfDJHqLDIO5t5lbgtbqFflvsymWyIyGfQh8CIHvXjHkyOFkK5boeZdmNIBpTczBYLomXx1
sSUwFKCymeQAcq7M6NtJJTjTVe96pmKPqo/cFgcCLbOhc4zd/P5sQJV4oxsDmdsJIEIcCVI0CLgI
TwMu+q74Tf75NJu+//xLTP6QOwgv/M1ES+3lfSN3piNxSp2SMErTnupAmUb7hyd++PhMgjH3F9IO
m7wborcy32V2bvoveKsiVieItLeg+F63rD9zyrLfIPHgYnBLo52jhypdl5kkJUzTArIqlPm1cvUX
tlI8Vu6t2mFQ8WVwBXVhHDcoqb6aU6r8STTtLTPsZeiIgdHPuBL5F7VRK57is8JzwjYsszQjM3vb
0uX4SIpl4cCGkiMadkvNU5hYMl35scywbolQ17yx10qPorCUZkmaq7+v6rV2tQnlDe+ZPBab3DLo
1E2O+0NpZpRtDdfYbhi/a3bH8Ku6UTE1F3s2wHekSo5u//CYOUzMaDHz4nd7/dA6kA/+/EENl4ji
GXs8+l2YzJHRA2JRV0zDSxBLBfhg+ICRgBASAcOIw8SLLSaBe7JATwsXhYPbP6Fr4MoIrn3XR3ad
5cprpKtJXl+a4Zb25iqQ1mu2Q4qNV/3mrzbQFigkgpxvo/4ILXsXeYZZgGoTL9XSlLHz98+qlinY
7GUrS4/KZU3KojSNidqcFVtnT762tgy2s0/eL226WAPtV3H+k2sKa8Cez4d/HxDAK3/GV53VI44Q
rkAaDuJH2ketT2otkfgoXCoA/tKyzaIWBzgQ1JFOI3ZdhWYU0N892YTNwrM2N+hTWgNXy7z/5hrL
AU+eHh+MZExOX3GK34zZ/X0eaby3YOwLNQzcv4tKdrohCknb1heoAsnC1k3zzHo+3kd09ACotl96
YGuHFIP0Br/xR0AU/C4Wp8MBIgl9EBBBlGaEpVDhP2tlB9HUgfQpGKb3H9VMo7G4XSz7keJ9w3F2
mYi9rmszZK7uJYMbYOlXRH5ZNlCWvU8uA7A9ZzpqCPWegxc5u43eql7Pp2l+MbfaVBcq606bNyIl
ZTqLUwdMrJpeIunf497RCb2kUT1E3s8NqoyYCk/4oZccLT06HeD62pp4hq71ZauZY8QCyagOl34r
TCuco9Inlof+512n4+6X+57kuo3+yZ6SbiO86lw+WFsxhAZln83xydi/Omz8zobhagl+Kv7On1gZ
M5qZHVY5hEaztezLQI3Bfe0TGjvngV7GlCSL8dct1YmfoleIIeocozR2s1pCBUDb55HwS4a1AGp+
nPk5d47nn7385ow4vj5QZfrW7/hNBRm3JxjbzHFOr2oXMtOiaUVzu2bMoPp2Na5fk08rdMFU+8D+
KM/IxDidOOTuMeZ5ZEJFodhNnxrZfn0FVJx7VKFsTzWSjzxtWdUK506QJGT5z5uErtgcTUVwdXFO
HR24bL2Xz665lys9E2MFTxgS+XJnCQbg3GeJTN247REluVwFWKtX9WTFzqMILwGv3reCTYPxSJpc
pEiJj4l+Q36dGBDC0LN04YRyNhV1wuMTK7z3Z9/yWP3G54K3n1WNEwh9lCcUG7hE6otB/n779tWL
dnvqwLB6DntJLQtg/dGCutq7Jo2P2bc2zG1viyGBIw+Gk1GvAe1NWrX6NhZTKPEk9hRF9zjwzS4D
ZMQWJlz0HxuBIwvycTgkSbZIQF+yTXN74w2fClFGQMQrH7AohHj4DLJMPJMZlAJcoA8OhvfYJ1xD
Hz/X3Sb1Cd/wvCUFx/5dOjwWa9vgrQaiRLpb+BfiuBB19o2/zp9vT1nwpL+q1ZrTa6CyJCWcdu8o
UaeDbMvMX50DChnxiJMfJuBfmqsQ7383rXkGd8+B52ePjrS8sAPof/cTcLmFJsWOc+zMJAF3y0eH
zf3qeWybzhfMpf/FrRlQW8FkUFew/M3lVswjkOy9NumQ8MiH7qSSaeKmiZALwdtNle5JuvioYVku
6ElpwepBlZPlmKsEuTN8s0t26NxJDVW4qjdGURw1nEvNMDh6jiR86Vj8ERV+ZxaTofYbTeefaKUV
bVbxomIN8mVnjsyRxh+EW/a/Hq2e9PCWYJRQM+GxlsWNfB0tcK70TogfffNlip96NTzK5oIaoIL9
r8ftnlSDad25QgXxeQ1YYpCV+Doek0i2Mg8L25SkFhwz3K+VH0foKD2LgGCHDUiDMCAmw1I+Xqve
0MsnMZj0gW4U1un6vp5tBqhkXqPuaNAc/WxJ9AVyYa4eXR3lxm2WkVd0Zg2cos29ldA3iX6R7r3l
R2DL9aKKvaje8KN/e1cEMcbqvdLwiUzkSGtVNhV4gkP8qqO1acasMlrNcNcySgAgY49DZ1yZJKUQ
mccLIZRPplUnqniV09abia4lTLlu/B1eGVC/RDN790Znwx+eZh0RdqZ072TpZQ1fJ8OYofIVcT2y
wgziGOJH9sFxqfjva+NseJSud2+XsH7Ps4VAvTv5fJ6KK95Mgd54+Mni3L0Pvw4wdBy8DScusoH2
tOZ/tWWYWbyoRNwkdtmOCuiFEDEb2/tIxBd8KEAwpg5RGrYHtzMU7KCnRyEdmUwybJunz0/uT4JH
dkzfiMp/MSc4ExukcDWpsXXRzPipWHySLz9S5CpL/ISTRAn3oV2sJN5LkD/sXfHIihtGeQg9+Eem
tPhp7SwD4mUmj3J55SfbqckQ23e3tjey+8Ji6XdY25uhtxn8xJxKnB+edYGdnBWHvQ5EbiH0NX9c
q1vEKIefj5AFmD9N3aXci38BPJDUmpHXbAX+1rQzNiWb2KITMsygRh73fOr4K2EADbR+aeYYmBc4
2kuXmnpUzvKU3KB573ZP8G+kAcd6jtJrdwifzYhvBC5KSf+xHjr6XfMxx0kmlRPVpHAQrUrZr4qY
g8U2jxH4rlOH8vtFnuUdeWNsg4/AH2ChI8L2d3V6HqcI64p1v1J04lQ1nWjn3dZBiK5cDiD5VjXd
JVZGwSc9kNdy17AMbWurNyGAhMQDURbXHRbm6nA9VbVDKmW9bYDbJWvuAiDAkDIhQ0skPbISRp29
wQfiCdEqZV1GzgpLpGU7N7Pm/Lhyds4Z6Xoik4/VGx5P9vON8kLEeK/2BheYWZpXCHuYbldoK2Hg
Ok5WiHSj0uSBc/ZEFjpNURmvnnRt0cpiVTZCKyrW+jNLp/D2IkpK3dDsHTFcs3HGkAFSXN4q89XB
7YnioGP+GT08KA2ErciSL0Kf2N0n/aLB2wMvLOlnKc0NuhjFukdu2yUkwSFUgaNWZ3eqiB7x/2ht
DtPPGYAX6EaGF58H5Mw5blUOoC0R1oBXEfMEsJllGD1Fi+D6tbH42b4EHaBaZ7qjMsSZAKk1IlYR
Xp4+OgJiWJtG6wtaZSiaw4Em7CXlaZA4wJcDt/bZnt3eGVKTLujndrsEajxuhmSdDIVafQxmqo0h
H5kibDW9EzuljzYZnd10XZwORH6na0tCDQjAwKvn6EBFp/LVIwuFi17RFqpdr1Izha/YeKoJtLw/
PH8wplekuUrf5xHNnx0QjQmiEJ59WueDYO302jRt2V7b0N1axaxcLG6JxZtNBCZx2pP27fNrzKng
WLwEnNpA3Tm7cTkGpdSb9HE3oWjJPjSwMJM3JTfJ+jN6uV3A/Nm8Lym2qetjzWJPmOzgqNtdZiQH
zBD7j9KcgwHj475EUEpFej9XmRXbuZ/9yrbTv8eKHwyJw5P9C7LdhJF9Z8kSqTTIEiCBflfSbyQ4
XTr3uztSqyZUv1tYWVQD+y2DvkM87Xv+WauBTvpeliiZQZF7iqHiXwtzBv9cTbn50vSrXq8Ni5nt
G+fVDHJUhlBKHCcHFNiUYXY6Jrak3dkHQdXGTF8zBHk3NOw+xqEGG4HeCKEjkdQprX6TE/xqnE5v
X/JWtxhQJ+RZRT1h0N3yZJSLpf2U0V2NSliAIc5vEd1TGzGkWz513G/XTOijaAUyRGqMEm+J6E6/
FnNy5fH/wFXsivJwJWHxW+oOYWZ1wA+YiwINw0dwKivo6DLSEGpGXA4AsoMwxU4Yf1K7BDN+NKgi
IoWYY5bf24I461ORR1vmkIZsiMjx3kqHdATcuM/i51F0D94+X6b+B8SNtx+UYUA4/tOE3q1oXxyj
O9eGY8H1LRvvX9DeSjtt7A2FWQ67GM9ODqH91gCyl1to3ceVpsDBELnyfuTuT+kvRlTHYr3PxIBu
mtzeYX2o8CJDeedts/AqbDnDLt5Ho8egVUy6HleBDgpRtU+zeTjNT8GC+G1/Q8uNit1qU5yPsitP
mayF2LRZcLnd4DcXnjWhlYjfq43fvbKiXW3jahEKpziAbCVte1tS4Cdn6of9saTaa5JyGq79I0py
goQA8AM8WmiSCpq7CPvtqdsWIi7eN8hXzvo6lJTTeHbDxnPY6NT+w/G5HoiCRog72vsYb0FQ5CTU
u1+uHSn1/Ee9uny2/5da0IiIByHLFxvPpBDVuq9A9pD7Vq8jHfnwpK1sIcOGlHlwNTuTcg8vmUpT
dEx7MHHclt4sChslSGMODQV+YhF68sR7Vr5sYlPXY4l64Qsny+PlumIk2P5YsCMMBhyCmAQVZNSm
17S/ByRS2O3xak5B8Wlc40ELgGeSPyyGcsIeQ/oPQJL49jIqA1IW3zQrSl7Rnhp7ocTVB9+lwY+o
UTRGnTAyyfBpWg7KvgfWFxWit0JxzuwcxFLjhMmTSwc+EZrbFc/ggzzje8PljLgW0uMJ2WAILg3u
quNT5bIo2l8En64EOzIvfjNS8FL1YYNc52GoUQ/67exFNgGR1mpxz6I5eehjXmVwpKcz2psLBIz1
2y6lkOAiX6m247H2wT3mdJZeHV7eUalE/3/XUgpslNi1rgcShrjBkFqewzJayTOol6PnUmw5PDLr
mZj3gBDXEIsVFb5m6Qi6VsUKprx3SQeSLlaH4TStWWQpdM+oVd9mt50TeK4jnZ294jtBHr2zH7B4
RZt7yJVL8wma5AWlsrSpOLuXGrW7sxH8Oq3TKi22XedRVK6F0YBye9Udcg4yQB7euWmeZFk2gCur
32/rZG0ff8HxMTFrntERbBvL6k73WyrJnk/FrP4WhYvJru0yml8Y1ZCmduZZ6Qm08JIqYGMPcsa2
yVmnaGcJRZ2GqBmsiqZNuI5/rrchfj88FSJiVYY6ur/mMhVQTuM0tUT5V/3MIpuuRaQGvbTxYJ2L
I7egNSvpgSA5dH0Z4K6GUOGQPiCgX2fjVtSiIXafMSMzn62p+7Agaz1aXwhRsMAXFlZHyM7XJUHa
F2syh6xYvqNXS3hbWXvp0XxBye0s2J9BfzrgjwF64jGoKcQshwp1FaxwOP7BuKmTPGKIPr36cXMD
JQwWZK7RdsYmQ3nsAQKR1sZR5IzaYXmbE8ARhjkyMJDoMpuzGxpWaa+fPOtz9me60GBYi9AMkRiA
3nOn07muX3P7JSj1wgkscP+79gOBBrC3PLmUJV6qViXQtkL7Jv5/FRJ0+YWLeYIkJY/lpzGmYmUd
ugntV1QoXJ6IwVtaheX7OhE2vFTLwU6JzoAqEHeRXKgtC0xVQf4LNPUvhB3N1l+92C+D/rLjJK59
uByEjUoQFO56RKKaQatJuhPPb9Xwx1mIcB9s5vauFBmUx6U/K8HuvzQAEA7Uu6K7oWRBJPEaSKeR
SeJCj8ZmyQTCbbFG7nX+ZBVYYSXaVscgT1AN2+bsWt4iIjNkxQi6ojt70Ll0fdkCJsVeLyd0HFyd
3Pq4Ats6DTiazVhqN1sNteqsT41/3shXHadwz+53UQHosyAIvziu7zV/+wmH6Rx2DW2F2NX0pgxw
ncOCgEAIIOdsH+eLUh3/tGi+Adt0Ld6k8czWjH6BSdQST4iF/Ki0ODCQZeu9EwVbio5sJZ8gSE6X
jy4hfWAFjCZlh3ImQoRRGoaOXOvvDoXlquoF7HUlEMMxJZCsBnMr7CoAGiVAENwEFouketOwnW/Z
s0zwrThoPvqxnKUV508IWWfcYHa/ZlzqY/+CEMcdBjHRV1NAi/QmQlIad0a8AxqgP9gIw67oS3Db
74LL7j7YeFSNdFcRYu/a9ZU7xEZVAqy7qfffe/J4mfdTr+bzCKxCASk2iqPQfkl8ZgQTlOVDufxj
mdGUXmlWlIoEdt+VoD74LDwW4i14649pc01qa2NJ9wT8HAhUosjqYWj0QXjMW+i2nEF9p9ymp9xu
07C6z3+xqMt1l21733z2GEBLQ5le+Sea8LhjxRlniKr2XoecC3Gqde94gvDIZNEQ5ET0octD22NI
DHek1lWuAVJWnjzNfLAF6EtnCWx9rnckNc+qHyBfStYu57vewqOJmpadiy7yDONWfJxuRBHNzA3K
HYi1vNbDDjY0PjmBw5ykurlzkVUkXO2fv3xyAxHG3yM1kVvyglPxEkgGr/6RMnF+K6EjUlXaiMQI
cYMA/CbZru5Vq0F9BQFxkmq9oPsd5qhVwajkp56XqNSaIv8Q4w/jycBA4w1ZWphEFhOqThVYnfKU
l6kriuiwAQamqz+b4DeVK8oBgZhLdJ/5YBepa4x52sBUB2BpdzcX+EKes9JMPfLHmYsL2wLLSIQx
fRApwjcaXXwxEWjc20wNh0RBvLBFCgCuGmUUQkkKZwbELwq+JiDR8DYFFsnokQh2Qbm9wqJX4nlC
ZDf/Ukas90QbICWgacGIG7aKAVpzlTRIHXXgAv/YLOQRex96popRs+r9o5vZVvm3nKo0prYY5Hu4
gnpqcIaRJzYn8nHq3WyQuGK4CgPuT4V5Gh+aWMAwhl3htSOzy9XK4zLuKFc227CkKxYm7+refa3T
hrxMAKqVMwiHGMbieAQ/9KnqC/4aWbAfkN00IwWIMgipBa9O9VPDRtdPmHzTZsIkV0QytjgzRH85
HOXKEW5zQuIVIW1d+K1x5NAB7yvahn8g588RP/YE9gWTptNs2qMF2l62n8HbNDbqUSQeHFiGMWZr
wXzna//iurDOQHjuY9eDS0nTV1zioVLL1OVprqcIT/J3HWDmvAV9G9p7gfeaR+81ahG49ErxpUeD
T/8be23c09WiRYKIY8WQNj9BDfxIXXN21fFGJED5+4kUsKqB0mldb3D328ZXkQujn5HKgCCIp/6f
woUwA/kt/gRWFLelAQaPvq8IousFaqxYXg3ypjmTlwJLBugtOfE8Um5ny/9X3VXRQ6vyeFcLz+yk
nG1a+rb2i4RpUOBN//2gB1cfY4YHQZ59Pyn0PAX4hEMuZEn4Jt2pAZoW1TCoby2+ZBCSh8PsH/cS
9GCEXmLZVo7c+J61m5N1hPEXBxKWJcOSvp0o4HF8xROmxrwxmP38PPX5hVXra1KIeX8RgquKLa1a
7ogWPWO259+fJtasU5LuIcpldTVBYaXcCOVjQaOFeIB7ir8YV9GGnrZnVwg2Z7gxzrVpLp8eqN2y
RVogurgemNZNy3YsOhFQ0GcCjLb8oDaa0TT6/78s7js9LiSLfSoFQLqSovntXJHOiUt2F7H8nPiC
MpsYIQ59w+tIRtZdJdCqWsVCx9R7SIgKdnWZM5m2wdBpNB//u+T5gfg8pqSSe6nlS9F9ZZszELz7
y2Tw90jpVnIrHY5C9vBVcYCAlkW0dqSVZfDxMC/ivKz7bXekK6fHBEphtsEKBk64Jm2pYoRUQy02
oBj6J0S60hOEGDw8KFRefJovexqXzyWSZYx18xjst41uxqPIwH/MECbyzgJYmi920w2qTvHyPUe3
3ofA6r8ohky4Gonc2p1jnj1FuJaZ9yBqkjdz5Rk8m+X/9AsKENBuDtfP6gNCLYPPGqipPwfMQf7M
hNwRe93+tc24t6SS++IbENCpjthSwA+EaMVK3FU0f4guLj4K5IIswlA+vhmN+YWWPKJVfl38pdjn
N79mu6kfCT9+7bJpmcFzIoc1hz3JT7Hd5mfq8Q7RyhvpDWCcGMBQue8OF8d1sJPy2VhA6WWQAB+h
LHTC3BjNfh5nFzsv5e9M9Pmk1Yqn1IqcAeUM6s0T2ho4BYJODGUcXwKnmu4XNRux07LQAxU0b7X8
DylSH2ObyPZh6jjcVzSk1iUkfrCZ5SPccxlgp2q/Bp2JflDi99q5f0UNiDCUB3gE/OBGX9/lypwg
Dq4dFjKefxQjpJlkcfC/VuM7Zintmw4BimaHv4MSnnjMpj2nelOgk75B1/fNhJm2Plu63/ENcmfC
RfdA3aC/BZUxerYMzTFhy1xLGs9eI8Ji8JirGKm7thIONUUV39Sg2+/LzG2TSkriVTSQH6qwo9iA
tdagBnlnKZj/lvP1QUMIYCIrbXmUXZliWUWOFF6uhIBmvngh7GMW5g/Yh++MgwsCZ9CY51gJMR26
KvMz+DLIZSJMTMM1LUMhOjASnqh5dG6MZpKC3XdUaA9HVs++dtFb4Z09jCT/Bs9p6id8Mzi3dpFB
JzcXI1rrUrqg+7e6IxQEFSRKHtWT0z0UFg2BMoCP8NBpL+E4PJdD/uv2A0VEfzm1pgFVLfPGo9OH
d47bxMvgwkw+hbK+UlgIZeU34FQBOEZMMh8ggrrcEvrDI9SfxyMTY+gNc2BbV/g0Fn4ghY9di42n
G0KChHmcp0fX7T2YIMRafFeyWio0mr06/KDzcWMXfVRdvsAx8apPa3L3UcK8VTAMjkKRY1mJVkP6
x+K0LhTxvGd18h2CME30OzZZ1OVna5+zB3TPRc5TbLMRKY8V4xTWLPqyaUys3oWOVJKaE0NZ2dCj
bGOqsZzRjKnZCTRqZDt0Krc3Ksnuf7Cy6bysC25otNN+fLNnk2z8QvvMUB5AOKvWkdMGtdv2ofG/
2O8NcKfV47amfllsE8MYQL+7Lc6rL1UZ0YXxMBryCorxH4fzNDlUlyJb+ZtK0kziEdP+dNj6OBXP
e48AnQf/xUULlFPG347vl7l7m0CAK9YmhF0kjmAM1HHcezJgHn7dosdjAwdPXwOlPjuKe+6QfGY5
aF0MFLKcVVC7Na2WVi0c62XKWmvqlubvMhZUkr0MkYzeCvKBXeSu7nLPGfjO4hGQZj/rwDRQdHhL
l88q1N1TNAkz3ObkFw9ThP6uGIP9f6yoHi/PUk8iTkQxJ1s/kMFeuGr3DzwxroNaE+Fif7pWMyOh
b0c+xBNnU5QIzBiu98sOdqjMJh1/YDCx7OIHkaNfJLJcUtrBRB+bGAIPxcwyrJLB3hzxynQlNPKt
0mudZNdvhWtI/F3Inyf84t2pBtI/jQAcIT8KlhljtZxS4bWwssKPHGOoJKjiNjL9PPjSo2zLHcVf
RZeO6lyKfPXygZ8ACVJ4TgcXyJzD3sh6g8uJTRi41AY2JMwRJIVJoeFzzWMlWVfR4wHjZGxKixgN
Zc5ZGrpwYccuBeJ8X7adfLC5lVekPwkd6vIOo7z/Q5jq3dzbQ4mnPiqt5GaOACEjaQG+7ExeDVwY
8SfhmHh4NhrGPbE0JpLIfKGdfVJQJFHKsdrr3hY4nqtgWXleUwGqptS3DoGTO9k9sSwbOXB2FNHO
EcJWNJOQSZaFJ1Y0i693k4CMs6zzQUOH/s/1Kldy2uDzFQtWWwDe6jpHSUpAK73PRZ/BvKrd1yJh
zA7RqouFusZC339uOGqXjR7mmpVuacVAH6BOSXSPUobrXcDGAUFNN+Zn65nOQ3oqnEqZC9SrndEV
rj+H9XFUoXaDEDuD9m2TWAYgB2p7g7O+QbnCv0VbO0ZQwC5aay6qOd3kj2GbLahFqEZIRXuTWkqL
CEr/wU2Re5ICVx53oVWNr05h06+IgGyJfXMIRHU/LU7EWP7peW5fzlC6lLnzuRY80SAM6m/k4eNy
JF5prRARH3Q85tblJBBIZA3fmVIr9VlSLIWL7haYbpjPb4odpiqoHnF0PRUvqMj2cqsbxv0v7l4E
1nC1QGxPbJ3FDCkN6qc12x2XpoyrpEm/OOvs3gYq0znPTujUWY8Quxqti9n4lKu3ujk/W3XrobHp
2JW8XZx3S01dOYfJxLKTuXfvThnjN4UYPb/cMtvYTvkZ8qDiWeaG0S7BWosA7sPXwcnY5OrcD/tP
FPGsHu8GNV+NXlQxaXZf0Bsm4FMUXwa4GPbKnr1w1+X2xTt9Vnlna/2aeB+6ROXpaCvTZsvbsZMm
ItXRGktVLkqTIWFjGfqX1Alt9V0Snq6MWQEZYI1x99ajzKJxgONKBt6Vk6xEkndCOA4NbplbT0rU
0c/aCXgkewACypggyXXNch1NDl+RcyaivepNk/YRdNlEB6DeMlojdW/zftGDQBxNiABzw8hHC41E
9hDYq/ePaAoPy1qP+cTt/ljUk5qlV7zkYUXNdo4zbE5J0SadMnKzrphuAAbA51CW6NU0edybHTUD
vYtFeYy9aFvIV7Fx5K6eDzqaJj0uJKf91bs1byxxuh3VimfZt/GBI5PQvcyJJIg9BzOKOjAXncu6
Wrj29hvnxAZM4fkNG6jHa3gJpWwtpVy7UVdQGLOvmIr7wOvuLqa5qUN+tVvx778Zr19tAKfzq8Uz
rwLuVfeCzh4J/pIowUVtQZJhbcUfWA8d0iP9CexSzGdJXt/qFfLjqgdR7YbaLgUk0lCFr/8gcwjb
Cqt2RytZAU0N4Os/361S+yyNpUnW236YNIuOrHnXM7xYPNqo/jOGucsxK8sQLbDukcSiwK294YU9
TBG5YSiFbpDxl09WBHCMENGLu4OxKALpFgSiyJiV1dYqxtE7pWE43k5MBj+y/cxt+uvLgr7fkx9W
FBy5shl7jxDbnEZe6d2tunnRTXJR0AyZZ1MU6aGTazUvu30u3pZHAr0N5FG9RVLbS5H1jwk/LkAN
PQ7Q29/WulIYwHPVQZQxefa4315sNuIyHnATaKpavVkyLRd/NoKtX2SGPnCD+WJaQKWnphrFN7FL
pFAWm/HUD/88xyvTqq9Bu7al+tO/XzYhbn6uMA7FCT34HXah9bHox3kMfPnWVQmaAtWlUBLtdUeM
wnMHRwF8+hBtAhb+DlDRKb3eRJ52yAJkRqtUq2aryWbxKwcHs7MY5DRdWqsLszW+V6kAc6KPAMH7
T03d8iM/39M/n/JPkYPCRD5wLiOkNoOGXbKSQIFcb1vCfzD/vib9sY1nftbx/XTVyzg4KfXXKkSo
oqVYF4IgEqA9ByU5CExLpZ7bcZTaRpXOfvPyGTTQ6dakXJPfkVZEz2QVaz9Iew1nLj8bYrtyRHYz
lgJRlH/nnOL2rbb8MKiOdOB/UJfJ/nymiK57D5ydP7zZ+MUXKbd+pJbTBTiPfTpIjgIleDm3DnZc
GV5ktEnitiGpVaX+BrLX2f9GRbQ3J+7FSlC76tcAvPdxuNv3dLlkh2RAhvSe/P7Adx23TBw+a/V4
Tm+ke9UVq9njCWHMoStwRCpMeQZTmpH1goKO71lvXKHBTymLVCqFoHyCV+nC0ZQn0CcgJbpQnatd
sfJdjQsVG5ZC97nJ/798BsE4vhOQN5vSpVX3o2nzVNozyFlAGfME3KZn5PcAu/qDc0w/zw65jyTE
S/UZlG15cSZYGZ7SIa9GKcbKA65WrBHrGchbcbcOR+lH/iPBdAgpYMtPpX7XZ9N4n4+BynhC6edh
cn9gJoOKNkzqY9W/MpaSMVSNdYB/moxMH3qTY1xBDkoriDP1Cw612C9ckyZnQyEiPyAyR+rfSY6u
yAr2gHibLmYqk7al6n1frl/X4yDoO3EIxntHKWhpdxslFj4GjU2SbUbtsFMTill/wff3/MHHabys
cBBVMybswuz9YZqrHqIr6BTIGkgQn/FKShHq+j85w6XN+9KdYCFbl8wG7vgAcQ1Y+EdRJGYBTOrV
8b4DCQgXrW+GMMSspTDwzotNGeg84lZ0pPZA3u6FFXMI4jQcmM2iJaHqNBk1nOABU3yu01ICt7qy
tzceVawa0PAw7SkIaHqeGiI9ZBTBD8D77mG054c1meyPCP/07otBA84X/Ve5W5zcSFxnZKQtuzpd
SpyDtajlRnyKkMHi9GSAICiecAqCwtfnFchI2rRinqE2VMgqPMV47ABEv/tTC2s1efqCKVLuB0wf
EK+72Y1Qmguexv68dEVD8G9ZulXxWFkOyn4ixoPFRA6b9FuR6iYTIdmv9r2TDzHlMsmQ38foqnh9
s+7e8HKwjKe+tDOUNP+tpKGhaeEKP1ZeWToem7wkoZ3uy3pqmB+8vg/NaR/5dJ5iTpYafY4poPAh
xbyGlampbdAda7kG9Rkjz1kxueXmW4pvkel1NRFPIkBjVhVmj0iGnwOlQx9HqX03MMSX/8TNrgGD
oRq+NVZlRMoDqCXwzVdVxrJl/JO5RYWW3N79z8P1ZgyuQmjpco5wZtuJ7UFPMxMg4P3fMZr5sCZo
5Z64GmFD4LQ/WI4p+fyKYCg2+3/AmXeChZn4laOAHTDfTlPqNUFVQmSpjEvmLJK7RFljj1opDcvj
yWSYnoV0XKb8Gfa/XDDzpTFbw+8OgjDcY9tLtv88k3DtgvJ+yoUSf4aeAq4yjsBSXgpKsSQy9dIO
62z5stUeU4/teXPGO2HrO2+MKc7j3JLlV+rIlNVZfmJuM7WDtYwiVkL4EKjOMeN4inMxH/riSiJF
pPGFK0znd+9aZ2dZS44rnLrDnr+72FjoXv5bjFY6gDUqbrjne0Gfe5y6r9VEftYIYpy7NiS8UUwp
mDWL5/TgJ9Ra1znL5I4ELvnCjlXHyxZXxKxSHRNGRz1ELIN5VRyXEIQu0NgXKAbEfB3vrOczWuDP
OaD9C2Ae0XGTfzb8aWTSPQovG4czlswpAjOwRlaijjG0EWrJIwmMKHZKiCnPmZXIkI29R+A0DYGl
xwsNoSSyMrIC9SRkgvP7aOqnxwbo3DgZCpCi0TJwU1w7RB6Kyj/lznZFGelZAYJSuwd+YafSqw2q
JfwmdczuFZ7GeFfbKkOX7e5XYexINhOdgqVQPUPJ6SDJPLLChCeCqPYvFl80gyvNqfSP2Zl8Je4R
YZiSpIUT1cGVT7Usf1P6+eYg1P7QDwdAABni+XWOUMqTAnYr+ImjoxWpz0Q6+p0ft6GrTfyZohXe
N3h617V67eZu2MPmF5vSPesq2YQ4J22JpI76RT3SrmJ/x7ZpOx3mUz5C0UPLPy48wpk+0nPjmBAq
DYHdZHV51sYlRDcMa32wlx+v5e4SOMePid/VPPmtqhB3s41j9TGK16/ncg4t/Pgogs2kv1gW2zBw
NJfMxEoFCo1ofG73kDFLlA6XICcP7gsAbXYKbk5I1crfZyhZ9k4WjGjp44oUOuBAYcQFSS/OZYi6
Y/nZdVFjQ7inz/8p3t5SLvBAz7Adlv2SUwDm8yLCgWtuak2EmT+SEJkfGJXcDHllzy8YtOnlWpEK
/QDsos4plxI21KmCrg/ZKvyxuDsb9Tl+CawCK2RlBE3QZpuwFZEV08/JFplT6Z/RPJR7WVZe28JE
VLTEtBnWN2VGuQGsDCS553003pa+UiuV45218edwluDxYGtPaUM6g/bILQKjSVwqp7GpnV9R8deJ
VLEtL+C0+3x2ifGUwoEWSBDY1EdyPkIdlY969B32aGuuOlgz9Gz/jUnFNEevtTS7luwql1RrL1RD
yGFygiXDWO/hdM85kIVFOhGt1X+RGUiBsUXuQJuN5UszHP/kabzmOIf5vUxjiP5druMsBguIUWyV
3dC/ZkwP6JqJz5nHn+489CV6OA768uxCuvcMKfCwu6HL5lJ9EAnEePbKaqzwZnONREon4Jum0Vd/
S0qyVaL5ToKnNy8cPg/f5qJ46VYuPBUoxyS3aQYbYYEjtHOn3q7UBPW37Qz81ZC6eKkTCDa0V9R9
ndFWGGmXhELvsXKrAX/I5ByI7j/cmvxAGX+t8hpXYT1Hr7g1MWK3a0Gy3W52wXcEU8xn2f2ZAT6Z
L6UjokMt/vlfQnnCbJSsnh/qD5yYMNd2Vcwn3jeCUSUefGDPASG88BNrMvr3rKjlXCwLj4DlVsfh
7eoP+Huq9qj9FQdet+Y8h/jbZ4VoL3TvRQqmtpKsAA4/QndO+SKSS8JsbI1sxMba/wKDaBAQiCLy
H4lp205BzdriBT70Z+2aEwoIx7FmSiQdYiTAqm9ft3VS89k8+3OsDapj3sCeYixEnlms97kYl2Li
+q3w5m3s0dS32025Ta6+7k5Qk+cjJqfGOjtGPOKl4EK8s+AowlFZuPhNyWmsa7uzBUmb+jpxl39P
N08MGd4WI1Zydp4HMPDc8+JUzsspIMCylU//yrMf+SVNSWYqQT14Qx4kYnEZZc6uhYa9g3C8lQlw
ZRtZzvKVzyMs9rcub17ERVTouGLmMh/fQm3c7C3kKTkHdlrczU/7W3N89DHfBblHKHVmPDWual1m
s91xa6LLMVXavmr6vTxuFEZzYLtLR+4Pe7avfHL/PM13ag1lQkgANbME5h9IjZ7f9MQzBQcqfXLM
pErfprYLsU/tuOnrFHydPLWwbmuSZAoqIHeK5sUxgb8B2AdHcl2wb0uXlp4392VdTiglrAQbWP9S
odJmCt8aDUDuRdXh649ESW4gGDiNWC3WZu6Z4U6T/Gzt8N1WVaoXgCz5GiJS522jvhvXSouZGWC5
qssbx87lfJqakmbN2Un4CcoQ1+9KORmMaMUsr4iAIuyQVG5dgYd1AOJJkLgTobJNSWw/xVXgEDZV
35Wc2oeqQp90OYgci8rFFFiU5k9h4wwnde6s15fE5CwC4/cmi1LyDstN+9VFFHP+DQktQkTDUsU9
/LUFYVidkuSnI7EPdTXK8E/lxDY8xN7KqOfVXu20KJykpcOwmIwjpWiixfTslwwU6D9bnSsxh9bN
9WXP3p9cXV86pSysy70bZbjvzCQ6K9CeVrgq/Qnm2sS1qP3xDmlmMnG4rMejE8fAG+RyZ57uh/NA
cEd2BWgE1mV3U1n+BHNEES4R/tWdg1nT58aRvVKwZP49PAxy5TUOSyY455UgvfNzAELKaFTBdT5P
+NxNZnCsFjdcQumwrC8T2IHSW7R4rsBr3F+CDrz7ARmO2fgUuRKCQ6ybdfJwCa0Q+H88CGMEbIYI
M44ucwxYO6FfkBxw/58JzoYgMqbrck0iUEUNa4yzknDDEWNQXvHb9uS/Zig+LDiVOg+ZA6HhkBkY
KctE4qSLWVTfWOqcUA1LeFq9PxA49QRYsb1TBKDTi6rAxS0q5kxErGA5n7Cv/esUe2Sp6FHbMVSF
RTxRC3nvWp7sWQ+oHu7HB9pq1ZUSnrhZNhXs15RVYYzS1+Bob8o9XpNDntRrWXfnp6ERcqWDRVmU
Y0Z9aBo26NRMoOF3h1NV1yj5+EPHeXDY8vIJ/pTNdLKsYirjyPAFqA585+4ROIuJMOUPRJq1cuV3
bJf5UfySC3K+FAWZdmRCYl3S0Iy07FZLUGrhiOxyxKmXIBaBUw4jeTyxdjppxU7JLTXVoZLT9nev
tBrn93tSuHU9lyCBvCK7TnxyNUM2GKqItgByVCAhjBmEuox0/o+UTzleAlJ2hwsy4HYbvW0Z9p5/
Ykrotz5XTZ8kKJRW4q5Lpo27DHPoATHglVmQYDd5Kmip0OyYPJxaun6JhOB6ag6+fn655ZxkQgSp
9f6kxtfyNccKEaKQABnxAhwR1qh0QzwdfZylaa4dOT55cQfeLr3U91uBosrgd3o4Nt+ZhbFmptRT
fMHmag1fbfmjdpsE5V1mLhIVg8wyMXAmLhePPluNegyZh3/xBlJB5OTQEPhUKsfMUH0+ES72SYz9
13O4ld5BZEYB3fiNic0T3dRos1dihDq9qUm2MWkRFggfNKxCvRW2SHB0A/Yujp8GilTyg4tEnvLB
Ne1b9snDwJ82cU0suwHzZsozxbTk0UR+5M7REW17E2yLs9qdvhLLKFx1ID3X1si9o9x8EgmiRxDT
pOlQytJCHT5DJXe8bNTBTC4Zb8bAnnUazQGA7MmU5GAotkz0SFeyI1hfW53Hq4V9SIzHy/yANkyt
limQftNVF0CHnMBRfKSJTfIz3Tkwg1rij8cYTMvIOTmOhxaIOyZ2KUHB6se/fDLoHtmU9IqfSDid
lB2WaKEiAmyfSqphJTVuYs2KLmFI829IHp8bDXfYrIoO5S/hzVNd7BHMWTuZNHRROVQcECePDuKA
7URLeP26ZgEsv3+bqbNZBLXBNQq4gMnL1r1bn3AEcBfja7kC8Lke4JcBuUx3lG/RmrinkCieDfTQ
I36Alo5Y5n19QurkWGwAjNuVRgyf/lXg6p8H6emv7igd/p/omr71jbpKhiACGrj81Ll9y+HW8Z7/
yrUtrx2OgyibELxIwrDD70oSyblT7KfIUduq7yCMR8RLGzGZgV1dQ2zBQ6tBw54URUpE0YMm/kup
MKx1D25qUPvkeCgQLtLHZ+1l0/4e3utO1NcYPJ+DW89mArFu/c6QczYuP5hQ8cX+K/thjOdi83Z4
wwIb1tkPtUUQmqeLo1vhRVlrSAhl58MBy/6epdXNrYbtmbogB1QgPPbLETOEje4x8JCq2KgDFvpL
rQY8UEM7Bmf7eZsXjt6SKAn2y1NHmHuQofgHV788yjXbIcqzm978IvJYWU7+2rnz540SGVbDimFC
+JqyVPOOho6zyn2UAv2kGtqoCDhzLcUTtOHVnrijHj5TFIZbfgcA81xQwzkhbdiT87eZ5mNFR1Fs
nWvvFtcWoeuaVEwyR8mewdUJZVqf5pgAoEGzZ3qif+W0gop1jyAcbptIosiNwarZhcF9X9XoFVVl
GEekL9FTsQbqX/1IaLJjyxK+ECnJiWay0gxKriRLxYk7QTkQezwVbhCNBrgGnnBWGZ1TqNi9OJHd
feKFNrqkUqMWzlW7eXDq6qaqqq2T6vaFwAGu05fn2rFEgA1sHt3/W2tt/Jm7cxPn678hov8oiadI
ZN263GrCjZjNibK5n0zjxbnEHrnS/UUO6inrop2ep7dzq7CeJBxfv5eWTv2LayadEFT5R4Us+hPx
2kCb8DmUmAMhRp5FcnscQaKltOebOnkVAJ8pcf0582aTOVN7G+VrM9OH8wphYAeGhZm5QqCOX4fN
jSKjFiTVMUf8cGbgFW6SOswVLmEBHzYhlzcFNlavVdf/NmQf3SRVE5u/MObPbir3EBFxPoz8FVHv
fIWcL9B131J8XM+7XRgQZT0s3mfi1FnOnuQW8MZG3yArMeuRslxbi+pAXoPMTM4ehFDKBGHxo+r6
tjB2a7TIE4DPGsee840RbrlhPuGnfRSCwekkQlPncIYtx48sBhpVybVkMgug0lzHSoFAcaxiBD4b
MJ+bdoO5cno4d7kp2thYPK51W9H9TMGOAyLT5ZhAkSen/tVEtvoWvmIDQ3eds63cu5grds+m4E3M
/EFs+Y1c52fyG+spXPzDzydJlzWUd269dLYNmVXyym259XX6LS8uZi/6YqbVqH33iNjeHqchAofO
TG1pOiKC1Wfntb3JSStTjNmtJiyr7wCBrqrhknSsd+hhml4PrHwIngwZsNE46QXw3kVInLN3nEu5
VirszDqYLzx3ax3uTly/OAVbhUtVfVkAtPq0JLl+fhPS+CI96X93CvfpSovPW2ElVzm0gacN0Mda
KZaEDPBslmCkkBOUIjeupX5a5BI4p4yadiWFLWJ+0UBm6nevYaZ5bBDwhmmBI9r93DTe2hugHG9x
wUGFXpnhlF8u05D9FHSWAMf1fbluFajzNezHu9v5zPYBAzDH4tr7VsPPjcSpKD+7OYXq4FDET4eD
xrx5u7znEoQhRgtcTKeZ7SDmQSioTvjNrpIdvqoJWaXjuV0EsXE44ATRCDO6nXhNPIU8UlpddHMX
KvY/agngu3V7fHhfAIJWQR3IbimqjVje8SMajHOOOzt3AtT/5Ht+jx8YpkjTE17zTl0UWHAPyKCY
je0YHjjqw+wRI94ESV/jaFOD8qGSFjKChPsPV/0KvRuJgDYhcE/xuNbSn03Q+qK5CTBvONgTMbUk
6WHa+yB2PkEOcdNd3fA+VypejHxhyMTX4eb7RuuWahFFig+dU7qOr5Acrau/fhC8eUrr219ZREbp
Y5mYEp1/2ZyR8hZkQa7rAEE93lwLT6H/vU2lp0MZNdGDTBI5TFXEPzQB01RC4xGXbrkiBUhEUhmX
WLvi1I5wXPtClJhkBXY3Amcuon7ZAqnrUymxjovqnMCdvnr8y9plxMtItKGxgYGoKt08g+r1iexg
kaGycg/dYp8dgxOHV9FAcqE09PiPcaB4ZBBj8t48T/yUsIUguSNKH4MzOqyBx8WrOgeNHQQl6Syv
nIQLMrfRADOtZx2CKkUC6T9bt1H8FOKVLRitlkvLomo17mbX1TBH3DDewuKu2+RmodO12chUyJMm
X9h81IAwfHZP1Im1dcOyHanVCcjB0yqG2rXt+XteaxvCIhwhQQZexkxybiDdWRgeVT2g5bX+rZxL
0AExj92Xiv7uE9w+4EHbg/n581V7qmpaAhL9qrBFYMPVZLkEXehs+cFOuuArwihw5/4aJOKdlEmu
kPBpnBhynNR8BUwWzdywrCqV4l5WJtMLRqhk9Dju3O1AliKPglFbDFFJgQekdn+VrktaQx1KZZoh
x591b4bt6ndVceCYWpbGQ2eTlaFJkIwoIJtPn8aRS3Z6jKVlR540Y5MvsZfFM3rqSmyd5VvqOY0P
SPSon+Udm+U10OfUyAwfvmIbNBYfpGwGNuKKjtyPTmKcpDpbcaoHS2Y3AZIEQzQFoBcx0xZsGcf/
zhdL5TMCxFJ4PWwZBbSBoQc8AmoV3efBXnaMidwq16NoZbfSqUY2pfmlHgb2h4N/3DJ11ApQwb89
7JfWv9xoqJufPJu/+q8DmLZZdekptwD170oda8xExATDsyAlXm4zXEZGASGgKzKkqNS0ts8c/KtT
gCmV5/ErZ301RhqqjXeWYOtmJ/Cp5JsdCwYfQaxKMPm1h18Xc5bFmoFaExcq3JWok/OiR/s5dzwP
hlfijzLUdMQ45iJYXj4c8p+rfOO1XASyxc8ro2771dCO6nPEBv5n2RTMQwIoQ4VObrwSGp+oiYhM
Bn+eSKIG8befjstdJxkG8XYN9b9pJfyRxCW9kUpz6y0b1sM9VICixbKhxc9b8dJYWFu46CTduAjF
aSwq4Wq0RxoLc3+7v1cWeNoTWI+qcxtqV6l6NMgrBhEJPEcUz5e1LgVEAoqdP1xRRA3ztNy4lwy3
L+1jZluk3XHUneGwN+kJ/qckCDp/kz3E+3w18+O3DdbIKurWRBjWLU2hZ7QESacV7pR1l74iEfKx
V4YOSoHiIS9c6WGkhI+ikgQT6Quu+wqi9Is2M2HuD2KjfvlO7KMxPXSR6kEwcOPR+1e/FWMjHNlj
xGRpzdk0aUN++cSkKGMnoh8OPhwOJjg0l0SPHdFWRKCSmmqKc5oRUp+PfNFd0T5+vNTbeE2xPZht
mQo0bbdf2ynL4PI8RKGulB9NiZLPkk+oKScYTvnut4mr72WQyHr3vth8EzwtdjunCLH2FVCW+H02
8TnevoPm9Uuu05FjJptDkH949nYbEfDimJmiNaSM/7pjtOWjc+OfMfcyKEzwpUUsCt0o7o6fzdwt
8n8q9XH/DpiPuRtackNkpCjmGBIjdz245StHS7rcF9rnzWv2iQfmKb3cRMVce8oIC+xXmgxQEIeF
oH0/U2bSq1U1QoMH8xXaq2DwUySMzwDFdqf15tvaNucmB4LnTdBawhYtgJr5oUnknBWkYaaqb/s1
GDV3Ldh69wRbbgGKe2dynG+Z8ILduFB/6PCR91I45Z5DWM0mmRKFYR5lnsR1OGonVsSCGOclg/IZ
oVxE3oT7pjO2oBJjyYc0IYIyf4KUYk9xqVfssdIPg3moFjRlIg5qj3OLZfXTVhd2yVKBWEsx8KAu
GoXM+8DWtWW36qvbD3MbWszRwzLThkxzu/Ij/s4nvqIW3M+jBGzFmyfgBGn7L49PEKDRsfNPdTjZ
YRGjMCxMo4kdem1ABPmfsYsKRlPxiWuG2rAM0gWEwqz2O4zNa6CHMM++y1UhT+eGhet2ti59UzL+
A1Db7djFGNH/KxTljN7rTkXc0ETvCiR0n6Te9RINTjz9+emI2m44sf8QxTZgxHJqsIhgn0XAoxrI
b+IoNHHV/TLk4XwNmfNhbiCVzmmGeTz7EBTgAHZ4nR1NKMPC+h12NFp5m3TmdOoWlnvb8ZO/HGw+
eTivYTxUpZuImnumqFmn5lpod/+Ij/og2iWwILCV2DfeG7u1Wa98R4MXtx7bSxhtXldvI9yaDLPg
PcoXv2EttXmkbroQBjiiDzdABHCG/CYwvwkwCHDwDYgb+X6YxVwy43cKwED+fcpyGokXkVyJCGM8
41Wrk1uEE/5uvUPqro8wJEMgwFQpRWSnDEEAAJVN2GVIyIER/CkuVrJPb0xIOAv+ruarMhIz3u/u
niS1OJwI225QsVUqUhZlGAQ0MTgXfmvMd0IcHJtCHdP/6xCcdv8/h3Xe/ckrraDcTYAYOIkocvnV
nGCXtgLH2WptuLSTcONXizF/+9abhxkN1wXSHzdUxDRUEhr040SJ+qtMnj/KU+fT96NQ0C3X8izz
ZMNo3ADjvL2nyKyFghD8shZ65CKC/IbMrlr6LdUJRs3ti59jp3fQrYXhTjekh9JX83dGxy9o5bLJ
l33SBf7jQmWEv4vDZ+LhEQMi1H1AczVuApRa36XpkopmmxYBTkQaFL6P5x5CRjmYd/tvufdhoQkP
Vs3dnHMaOV5Ax4jSVkPlbqwztzI87FKvSEhl+ld0ssnqwmOAfE6OnKDSViMMuixnnzYi4edl4dWV
imfSFqZESk07btcxH/9DtmKwKS6dgVGc4JYul1w8VHXK+VeO+giXe+ZYZha+fJCS7epLpNjcOhu0
R4Rn02f0j4InsifnnEP44H6iuezlUVRt5lrElpNgj31zBVPbbzR52RZlJFOUysCbY0GiE5xoo3QX
IeowzSC1mLbA5heLllgfKlX8M3HEkvchrFVFZ2+T0Gfhz14G32m/RV5EgFoXZZ3Q4Lye07Zr0PuR
rHuVCdT1hoFPqyYk/jKod44ad+glF0hV+If0LY4U3suEH42FGICfDYmmnNIvCHKHiO1mhFMnklR8
veMxkP/cHDYhVDifuUP4kdAHOL9ajSvWJ6Ps3aiv3jZ6wkdH46o+jp7Kt1gNNK7uIlKxygUcGU28
wQDTg6F3o7iNBBJU9SjLMFJm5J+tGouMvdpG+9H/G9qaREVVYbY8ZdGL3yvNc0O8UyfrrS9r44n2
SyN5mQOTzMH+kRAJRex2KdBY2oz25kehzL79xAl++3JqrvxlRBmiSBMjSocyAlferbK6QWsvw3n8
bXDd1I50hHB+Hz+Br519RsDv/E07QVRsPrXgNy8FYiEPwWXnjMzDEctAMj9vIUpu7hHNhljC5KH9
thtAqhXYEA7SvWBwkWBSPdLt2wbdxmrrlKraiiu5dtxuQLyYK2plseH6ZQdxvHycLlTzaxkm7nsX
Kf5U3muKopNOTrf9ierk7lz0HLWLCto/UD9MvnBWYMtwa4kRI9yQXJt0+L1f5Bc/XW+y6C5LFhAO
Sm+CtD9BMm4+q/RyN+Fl/nmDdYvPX4/Uw3yjcFQlKTn0k6ITylBWiBZ8LCK/WgLW+RW+Mk5acmPT
i4U7/9f3NhZ3W2EnyMj1VjXHGDwkh0i/eZ3Ckc8TfQirtFn4gMb/VDdQFkR+quAfMX5JK+WVfnfu
hT/AjNJcoyXftTbIIvpd+1EYHKTcNOq0j6XeFTarAxiKV0Iwfip4vwsnQiWElOUzstQytyq02CGz
Mab26bNFCR/k28dY+/QAeov/+npun36DFiOBrlYx1LntWqKXAWu1pDII3sdoVvTXMMZ+x4XLR0Zm
g5yjgKhCCdmUKgrMqFJZeG6euWBN+ik75Tfk3mTXb3ryPanIqwfNoRrzcv3gbxu93ui7lhhduV/T
ssAjESKk/XhZ4Kdacjzus8U+UH4asYA8aHq+kyNLw1+3U6ar80DFPnaMcpyXrigtr6fLATZSJVLi
FVMQIqNagyT8rUB2AB5adipDdVbpkJemGIXE91ZcqJ9Z5vM97op1Z1amKliYasdVxOBZnelmSN3a
QSiMykGJhAgck/FUqtKj7E9AWtArEIuZ8TUd6kJ3WtHoLN0BSbnT5qklpvwu2EpiAmmSMKsCiYE2
F6m4ko8YoLfrE2561h80jfNEQ5sqjy6+kNKmCzyOfcbd3nzDoC7opUhaQummUIEM49xdhQkf7Y6l
YX5iGUZn0Q7ui1rif+Iq5fgxkPhJ5wBf7SIBpv70rTmCbppOmkUT9ST0O4XyNYnIH/QC/vxqPVM5
PdrFCVrHBTSU+Uo4pKkjWwGBNYamLED2AqTNZG43nXIabDHX2bUqY3IxRcGrNeiyX8EXqgJdf029
efNBCAOku/gmmRt9s6WbU98GNiV7hFRKzVLWtrTFPYTum1WB+p4Tt3y/10+MtKh+0FFnuLkQFOV3
xCOpN2ZUfcRZcfmO6dvTfD9mTUQyG9ZUd9CcW9mzp461JFhA3r3aROHcMwnOBYBgjWAwTCNRGvvC
ui2sYwaoNHOou95cSGMeTGR8DFzbHws3ZTwXXOIJ7Rl4/aW1lQXLV4D0nxChBTG5YOZbz78nvr7G
ScT4nsOY2qcgNTCDV+oLOpXxJojT9coCQJko32P5o6zWVJ4N5i6bQnS7Y/S/T25N51BbkrFQ1B9W
5RM9BCX74Xo/BRb1tgphSEk/VD1puJg+xJNn3nQ8kSAE9+WS8C3MKcoZYylY92fx0KMpWmdfsNGy
TzCJtBpnRJn751viGMMPm/2fbOINkO5izshu9oj99SWOwQamGUUmpTbs/Dc0Q6lPqobKU+lZL873
4aO4S/ScslZOkmpeBUI+eyb10hZuTnjgnJu68dMg9Ig+pGHFdSidxTEjAnt21r5sPUgCkeZ94auv
ri7b0vMR5/ZXsLggk2p4B5P8oYvRmpl0BmpQSK2VUvzFpGYjc0UCQPj7WXkPohGeftERexyAD4DT
32ncVmt2eNvmCJ1miBTRGWUKeercIq/EXuTCCEh18CZGsrtmHMS86wvxB24wvImPtpH2+n52GLfb
A+lXj9hBr8HdqJI5Ou+TKwdNDvP6OxADRhCFbp/rBHk/5mB2yUkaTsNsw8KT25OWtUcAnXIIZq+w
LpduTfu+dbG7qPEGWwzlowkYWuU0fhFZChIQhmcdZrQ0gXt5IffC7xnFQF/6/InHAnixWkLxfc7a
ayb6xaQxozL6Aqw87oV/YadivFRZPQmRwjPh60ir9vjXg8J/2/wVzqYON3gGT3e2uzqmC4kcXbBg
jLwdkV7oN8D/pxZx8VwpI7XS1UexVc3EQbAvp7qzfFWMIzC1HaThod7pZCNbE013jzMimxNGJE8E
ZQTBuXP9mK9ffJLX0s8KO+8GIY+RYhxxw6VLa4a0FhdGYO8QNhgy2TSXjSouIUtqaavZGh68Y2gh
1Eef/eqVs4rPPIwhJB7QrFtC2wRlnGRClpmJz4AKurtS5BzdLtCgi+9qHABJVmdiPaAOvfJabBIN
ceGV6PpkMVrmyrfxVPpl7uUR0+pvzHyAMzy7jHUqR8dpmP7Er/Hp1CUiCKp2HBVPtgdkfwP7OAFZ
j6/Soi26Uo7fxjCC7/zQYDIYesyYVUuhc/3fab/YNAFp6pd7ub6P/UJ85D4+opSfSpyMZX1bfPv5
LoxczhGsLJhW1B9Z0gbhkqb34Mcp3k6suf+4D+16fPbiRYiKOWrzyAtGkmLgQcuBzO6ktZ+Bw5bL
vKCITCaL/PlD+pP9V2gWrkCO2DdCYG0sx8CmAQkAqkA8EbNDuEhIPU2kABVbbCNJDuj6ArDu5RB0
choU8pA6ac0GtNIg8xbauFYOtmAuAL/fRBAEf4bQe1GYddZMYWZLILSX6VIn/yqy/Tn6aYDkmWaL
axcJyZkuX5lKNFA6amNw8WtlRAquCKyjXq2MzZOFcjSXZZlyty+LApdXEoUP88Ny3OQbrjXbLb1O
FsElEy3UpqXBfUnu71ixqzq6B0cfxyYKZSamB5m9gIf7q3fdcua7uO7A40nTcU8pbEOmsZ/q+qb3
yOuHybVdbKlV/N+aJcF1ww997dYvj9Eetn4xcPjwZwL9XuScy+6eoCjcogc0HEJ9WflbLZuT9N9F
xTvOW8OlLZgMyJ6vl/XymGEaih7eJVDJME2FRow=
`protect end_protected

