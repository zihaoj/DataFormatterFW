

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
peElgUBnFYE95eKYTfZrpnIvdxmsESRHI8KsUslKl3wxGUHo4Q350QpQ5Daeisknn0jkGzHu55GX
rcWj5kY+nA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
foXL846WnMuQyS+KnySX+Um8/BzYDJh1L/Vkuxz872SKIxAGcCGxqYVxF57yWDQolsPqtbmbTxiD
2XI0fyevzAuClOgGeMP5ZM88Vm9zUmlH4Rixwqs38I9V1l2L8Gvg+NRN95ddYuuiy10Q/Pt4UEEs
qCjQhrRbXX1UTL3tnew=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S7LVSqsd7mNTg02/lZZbRNeWCeanJptVPdmW2TYWEaUfEG0f3QgDXN6cw/ZtDCxyH7QM4o1eCLDV
RxW6Rj+XGbob/LSYNDUSrRqgqf3cilsMzV16ouyMdQzKDi+/yGo5EbTxg3o3GyQMx7rclF1gU476
Kqle5cy0G5goKQaLHYAtAcuu5IyFw62vJJCwLKeyLk89phhJigrHhEAfHWqibymGa90qdDo172bZ
wzci461C/JZoOjYiTJSPfBMtWF+CQn60xf/t2CPjlSGdrCt+lEUMkQNtZUjOFas7Z2ND5N0JOffg
Oby33ERGSw64g78gh717FBsgC3DWgp1tEQ+Pcw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DE4yvRnHc7oO0HWP5V28l9C8UDq2AHTE+Xd/v7COjBqDFLp+G8yc4rfOTqjOcSMNsttRrOwsbcba
7YcOCAiaOLriUv1Gry3a7kcYiqvBODr6cEj4nGbLinNtjT5raCIA9alFqfNOgSGkheyTfqzDuGa0
z/F1Lzh+WG6J9HzTI58=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
reCKS58wk9DvCHzX2jTuq4IGql4vvQcZraOqLFE0gj+VqiVbOC7zHTOkYlRpG5HtC3W3yZbAF4YB
CbsiltQhm3AfPuNR3vYI2FGLfud7FKeiL++y6CbzGTaysnARY7/FTuNDhCX5jAVm3MFsFVB0Fn6h
m/iRfUJGvHOI4Maw+HD9o9rbNphlJF5aOxGMoI+JxKNMsk7o7W1F5Ce7gh/sReh39pbvT1zX2rjZ
sSrRI1kvWPBRd5pNUI0fINF9C/+wgu+qPRNx6NKuNsUKzV9LjYwEHd2rmNuPVZ2NADQdFTsgp0aa
4oOnxY0X3MMLNsSk5palQw8GZMQRc0Ls0J4dUg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103856)
`protect data_block
ET27/Ko5U6OnH2FTwkPrg+bz4jtw2MdR6r9qvQakK2dm2TrukFFTr1EqfWh8hYgS/OOdghNzW3yP
GbPVR5JKc2lIDmgBYLsUFU/XrDAzwRr7S4T5LQlQiFjLp4wHLUK69K36y9UDesZEshjwZcR8ELly
R2IAq/vf8x00o28J9KV1B31ALQevkwsEXhpUOfjunGCxULBz+AivHlofYUXaNXiQy4+rb0D9plQQ
fTVNwaumg5f6yPG15HaQsJQBowy+TFPXER8zEQeo7np0tT0tgtB1FYwbDpvppRDpAKsJkCkrd/xt
twhEgm4Ndx3ugiC0h1hGQzE3nVUCDEyDeLri2QmV2X1IjTSPqwKypVoey6xxVRYFaU3F/bCrEl2X
2A4FbFey5+Wo3wh0fS+rxJSqntHBvNMbQs0v/5KWBhfy7xFxOk8lmQSTmcymLAxaA+Hf0Nk1Jzze
+a2N+acsR1jdze6IEldoJMaNAu/1LDkA0LOY4eZ187L0a2WHzJDN6csLARRDzKqUfWBHvDUhl5sF
//uZEAvtE6ijRiHLdwDQCeHtx7Jz1W/wx8MqBjExpMSwJRn2XZU1ASeAWgsLYSrnsJS/sbbEfE8w
KjbX8LMxGX4Myz00RHfZGGLOdpODf9WyxrNYASRHEiE0/nHgiHQWRUsbIN8daFL5EfnxGEKxOxPX
G4TYFfIGl/9kcylvCsvloTnaxLN5Mt7PGwrTQic8NuXVpjJfOiolR/Bz3mRJqRIu+Cp99Ko9Vhme
H9tXg/Er3wFLQcg/gPKmbHwr/RoVdxg+w9jcHZnKg/pVt8boslgX6qBKdobKf6KDfRs/ayhg1wqc
HpT0fRFMaHFEX0U4OS/Gmvyp3sDSJlbMh57H/6sM5hoLnZ7acF+lWMtDIyk8VI8dDd3B/QuQfTlk
YaSEe2Qi6mCotupP2UbZWoIn+DKMbPPYmxDIwSqxHWBZI/eEleb3PGWHe/+170N+eKwPFbseq/xT
1nlFgxmCs/s+W/UOkVur267jiAgjOnDDbVnrKXZUZp4t4Ml4i+ay35GICA70yGztIrtbM0HB18Fn
L/jtUirpiPWVcRwKsxXOyEdX4bUVtjUfE20H7t26rpV3f1k74tuYhHC0S0h7PmNcZuQheiF2o3ON
hprvCX0De/leGbqzh+kn2eBtpSfh1gLZ3R9YxGBDjKLFZfkMZ6ZugentQp5VymDRj5A3wAEoeHTr
tvzHYEW3gU1xd2RiSwbtif0B5pjYHP/gWs6QwRDcusU+STsRieyhI6Sxd6M6zfzUSszhUBp8uYSJ
I5GCMe+ldnPuh8nM6W7O2z6sSlSdoZqP0H713LlJ9bsMdxyHrw0w3lk4oMGzI1VmVRS6Q2h/ofOr
WKKBLoqWzlCDS3rL3xex+tYJdtzuJpv5n8x9SJA4uisslHIIjJiXVML/T3WfvqH3VBXNS6GRZbq0
pLZXj2l4Cv2BVaPOQiBfe99eVbBBphvIFX0WNW42C++nE1rjxcyWJu71P4aFJR5lzVoqYV3K9b2P
xPN3Isbb78jzo4ovn/957MFMEIIRE+58pHg1peIoYTWtNaMHDPwOrAbuyNNlwcQjjZxTomuqF4Mw
TlYYxTQrt897QlmMfcGjIuW6p/GRz8GE73vz8D4zk1TfFFrmiIu60FEqZAPpSnNP78e3UBXXwX87
y3qRggHuONsDl7H7YaQA9WdpYzEZLCtUNDgs8Ap8epWMqqHF/GmwncKccRxkZTY8fVGR61kAj2J9
XAjpNAUmMr+J6bJNpsW6G5K/ZcRBGScATjHSRtscrsI6MVG9sLwl7m0i11APuB0OpePqYv39NtPG
V5VbJTPmrYBEznCWaJg4WxdkO6bggU830lBNUMXO8OXvkL/iWYXbjFj34BTF83+weVHREuV39NJr
3wq7VUqIOlZF/c2oi+wdjzss4oLrHqmLe4wZphCDx52X2WKw/XFMN47deG0H3Q0NjbiF1pfq3iPd
J432AlKkNQ35lLjmdKweVbmHPkXk6A4WFqIIw2K0aH7zJ2pL8wgCo9535LrqCfc/+jRo2qu+s0u0
B2eycmHsVJN5ytbB9dTGfcMqiMTyilNA5lztplaX1fOfOJqX21iQBGsYIK3pMO+km10+BO4HsZMC
7d3cUe2CTnFvwXv0tksf7Owe3MjiFgf05xtEVknsSSvCTpsUK6nK+ZPkPjagdZpROObrEcsZroo6
eTUwQboHHggTBJwDp3m5DRoOVH4/hmREdLADe81FzRa+D2G+/6HaMJD8Kfa4N89BV1kDqnSfJ83l
cCafj7isoxmMLpfk7VWPa9mNU+q1DIjO3dQjRewsE/dCSjfMkUJoD0AsWHNT96mB/nASgEpcntV3
DGmdH94b+TJvjfWCIVip441HIn8xV/n4uSZkio+H273HjAFSzBtvuUTRk8Ged1VxTr3b/Sc0cHwn
WlVhFnkeek7R7UjOAN8kzKBj+dfmOgj1EHDULdxUQMOdfkbTo2nonAvbhEjMkMACh0yAaeD466+z
BM0rD2KjjlC1emNgTR8RMlm9DWdzmayq5OSUOGOH3tv0PsL3EkCkQVRazknBNp557QnzgzNfz3u6
Tvgy83pdRlwr18BrqCBy4wm+KkYBmxQ4fl/pHDFIef38PuCROO3kOcjq1zGMO2WAnvisayfQN1S0
gq0KrTVvylYTxKTj0Cf1Juaz7FeAkDWLUOWj7wT3LdrpUhI5rQfaRI7mtbT+ye2GGrKZCUzDTWfp
BG3vQnl3MFvX4eRImoB5tDdJvJeDSdrq2+Xe5WKS5aLXmTcgFFV3GebcACxTuDYPV8Y/iucpD1rO
yy8msngAHMq0vN46fHj6mi3vlPS6YXksaNGKT1acukjhTB1dYG6e5k4O5JeVhW8p8hfNRSVZ7CCG
GiMITkiHjNcWYo4b8GqVEPlEai4jNHY90s2PPHM0awrY30W1xIbqdkXPLeb8LtO0EVxmKJtWnlFs
FcpFgMgbH3aiik7aRtieYNzZIe4ms8KqXkZK1J0iWHTwWVQ66pYYtezmEjixeUbAB9M4OVSp6w5H
gZ8GtJ3xwO8ART7wCmZ07B570GX9INQQGk/JcRe/Rz2ygOSmC+4TzZmlmgUh9itkvJjoFILtyR+q
JDx6c/wR5cgPvytcfCSZbe0iCTR1BS57OP0wjHUYf9i9k86S71YNmM/P0KEhfgy+QencXB1pnOP7
8/n5HR0zSXGkNrFqAotysWtiuRwVY3/BwxmmH4fyFA3lSpSSVxg6zEFcomplHxaC2ipNmsMJ+4Xd
8llu9DcxRXe53o3+bmjJF6I58XZ590SHPtjkykCvToOEMBuiETfBajWs61xnQoRNWlHAkW+uO2V0
hGRKHMW/3WEEdJ1nKChy29rQVCy8E2hWTF0wKi/w6FWX/btO5EGknSJwOpiwFgk1i8fp9GBu9i4J
DqA/TIVHdPYn+CY4ewd5W10j9sxWaLzXej2i8hB5nfGSFfRMhH+5WjxfAmghKTcsq6DqilLbxxWH
fGkEXhYBIPY9aSXRFhXEgOV0HhY5RMDI/NAd1axz+r3iiAmcf4oJEW0LrR+XRyirfdvM5fIlli3r
sCk9xfgB1+oWiCFK7SpdyM8AbqyEOHTkwAojscNZFMZbJ1n/gwaAe1yfsDkYHyHfZVi2Lz8uxSsR
/a7Rmx9KTCfyOtRb3MGwYBZEbhi88bKnuDepv+ZXgmmzLbjuZ9CS+QxJRHJRYO5nW78OJQtWyPyf
/Mfqzt/4EqzD2ov5KmqKyFPPW6zwRU+C6wEowb6SHtv/D9IlaT41dY9sWL6OmDHRgeyt1Zq9B/Hk
OIHm84vEJ/Mf/2vetz61jIknQr/pLmyfhBYp77ukqPYpB2cMbzCeY30XJEfWZrEE2MpjKCTdFiP5
XO8M4BkIEhsXvy3fuZcslVXaWiESJVzme0WPcrqdcyy83POQM1JQv1J/DjW1wAJAhVNmrTD63NKO
9kgZf4gXqrQy25smMZg4GAaTviNMuKmz9CzT0zEtjpUCwLUmT7W5khEEuON/C5pXdpImrfllvEQI
8bybO/eCgS6xWsoZyaxmNzuwrCq4XmZZ/StVaYf8zgAXWBSAYADNVz/H5HrCTaV5OEAuLljm8IxQ
nK32z6+5ArdkoS6+cBJ3mWIxmhF8CUvfiVykJyxedzEnuuVAqMGSfw9WB4n4pyThcI/skmSJEr/2
afxt+Si+lTbMPDJ+nu6aEVmo3Yjz9xsoczYhLRm4EBsChCSrZyFHlzCpAuV8KaJ4X7GtShJP+Dmr
ZcG4Wo6w8r0XtxQkFuaDRgYlR6kWFGG0ZQcCyKEvbLwxSUn5eGPzGk09hoozG+5bnXrNb5MJSTD9
JFup33lm0+pKi6XOOLw+w3buxUUgCbH4DO3Pt+tFq0f9jofxhcVYg403kT1ndowhH8TwYBhoMaQn
wfThSSCkadtCrBUPxuZmwJj97MzzSbbaoxSUCK/MM8r6IKUToarhWQXUsp46+dnpGTc+DTMawDrp
r4iaohw+qF955otj4JozOAiQ9jcf1KMmMWKCxo+4kZAkfFDTXrfvbMj5GZt+lAepS3i9vOZ8pk+H
fD2VGmRd46yYQAu4eBRi/LWfZ3mJciytMeQG/qvMZRQMQ5qgPt7IGCB8rwdG0Y3bvxbqSqiOUbmP
XfDY/zugPz320fkqhpsrgU1GgV5FVfi9gg+ZYaok+hI34OtOreSP1QGXTfR48A13XEyJu095p/mW
ysL7qoXOS2sS+vYi2akZcdaaZPgbEm90TSELr96m+DnkDQNuTTZKMETY/Cxhtyq4tvT/b73eD8As
AZ3AzVeNaWZZLmTT/G9fW2MvLnyPMEovl7IPokhqa+QaAub36gkBCexsLMD6I+IdynNrVUp+vmxQ
wEX2jRQmYeGI2M2aLWvFAtLHUpU4ZMqbvoK4QVQ33mQQ6hUWaUdrWeFbDWAbV2SlzQ/Phvufl6DP
Eg6ucfzok0e0W5DB89/GVPXBN2N9lO3Rn+C+wLvfac6SkKjaUocJrX0eN/nL7L9/3XEA/AKlznpE
crnD9+ZuHV5leTkz9mTLK5g9Nycwp1oDe6SxL9H2FgHffsO8I6OEX3nIPxxWC9NjAHmW0nnAq2oj
+kYPFTLWA7xUywMo1Ycw5YwMh51Y4HDqzl+LTMRKgO1/8j0YkILr9js8MzC1K9vOENNOqrzT06sm
FYrNzu5ZJSX3Jc3DtHQPlgPa65mvrKBWQ/SQAoLMV2lbyCbu4ZzG7K7/adxcKdtZ+2BTVDpYgQYF
ZeO6Fs+bnh3rEslNu2BtTt9LG4kvTS3Ljy9N3Xz/JqBngx8ts6bE3WyXvirlEuvcAD3mlUbvqP5r
DgNHeIHHPJsyMxQdwpMrMaqonQ3NfL6x3MPg12r/wVrUMlrSpbnsGu0rxFnPWL1Xy6qaWvtBOAaA
nFcYt8p2RnOwhOyhC6MHEMQvYE5qzD7INUfrYaFWaPHLXtYfAoIzhf/zrFF6FGztRNNclwVtEdET
qD3HCDk6T9pZSPiRcC6ZV19j094Yrrl3uUw2U2W2EYgd6+oYpj0ko57NRJVPOyLn0leVP3JOQLMH
5dis1INOo4HXLeCCpFidBLGpiKFq1IkF5MQk9/ygMmt0E+3iU0M6uooWjPaLi5XmetpxZZRPadRr
Z/k2FwSRKjNQIkKheOuNB/TjCfmk1BiiQymD0OKG1eKSWjj8OhZVBRbMI7l8ssZWAql7Cld98H52
8vZi02mv9ojwdKExfDBZa0ieVb0xpErwZYB9gG4R/hdOeWXqDFbVWy+lJGY5zgq/VixCSPbgzFHo
KUI97EPmtMmNG2hb38PpnPSmMaz6W0u1qnkhWYG/sr0GyEfoaiK3mvAItoiaeZEH41ew4vISmZhA
O0aJciPuZ68zNNGmtgnW+LRHTj+slAVmgOj7WiDAfi1Wi+eGKRiiTQG/WAdwBF7ScckrMFIYmyOG
+nHnAja+2NddjK/B2ACkhpZjr18Ke7g+MnhUnX2PE2HYnYKHUf+qmCdta6z3C14hlMkK/A0ajt7w
kJG5v/wpIk+JG/lIv2iYlXeA7MQqYN9PBqDXzASYMU2ei8+E1MRveqAIxusMzoIqQNw3GXhgzKZC
WXBqEWCRJBQZUYb6FK6Y0kY4wJ2dI/WYtqyzPT13k1Disdcs0oikelDMPdDWseM1Nn5KuYLAXVNE
vmob5N+53x7r7KFFu5omElnM4tbTdUkXsONNVqRz6bB5dOsopMQvzbwY35+rlhwa2xIS34nOYOcD
AyhCXUvAyb/173vXJVPOIl9wlERz9u2ocdJTldUOC9rbmoUKebKZEUCOvvctIajGmi5UcNgMQTUn
G1GNbSCPRsYHhe5Kdcny1t+2SE3He+9zH4tY+OBBF5NHIHCDXymJXPFuDEHl75I+5dx0/IYV7Bqj
p4gXKllFgRQSjKGFhXDIEgYYfW95yDX8ETqrSvNC5mtQgnPHF5z9o/CxAzaEh3WfRn9IczHARx85
I90eTmy90xb9XxKGIVxQqROsLAGk8gO1LuEQRIwVBIm4hU6JaFqmLPx5Tt8A7e4UU9ZUi/oLqChQ
eF3qpNZJiryqxeNOXEcbaHWCZGun/8IYsIarzw/7BUVvWfYZV1Ss/ZcIu48T9FdnrlxyEsy5hBvo
Na539Y6ccssRs5WqR95W0O2kPug7k21Hai0GNeVeceI0UoXH9V0iR0MeIXC/zeULLw82Mv5g4mIC
vz67A69wFCLL4lPGMHtHsKyUVAsU5Ru7LHq6gBIhtsQhNYsYX3DSTcJfrLLZT0OO8wpFDskUG8Dc
eXTTd30/YW5K6IhNDm4A5gWUOiEozQBpmcTQYXdkGznkkWmAPRf6Qdicf0fh96x8tFiMC1Zx2s/c
LV6TrRsrMhdADDc4zCj5BRHinGUCP5+Sk7eSNemlkMrDr1MKviMHjnt6srxJegSnTqe12cGNyoF1
Uj5VbaPnQ2zXJqoGiIVqLpfNxfLPW5v0hczkzWeRu98tdko+nmHtr1OKp+CJBaXEiJtp5Mg0kXnw
VwxOmh1dEB+XKyGnNAxrgYH3ZNvj1cUR99xw4DiYyQzy/yImMU5T4VBTKN4SqF98Pp4gqC/dAk/i
eBOBRHiPP+1uyVBlzKGe3xrVQ6hzekAjNs6tafXJA5mwoPsoCpN2/LDAeYGEXn2wCKM9WGAq1Lze
qHl9jd9MggAMZNvbPF0yxnHwaZV3mcOte4q7Qk64MYO3MxH1YLg2WNK8Vd+gbWCMZBdPbHLYW/DA
BxaNOhJrthxV95v5X8WrNhBJU7lwsaqdfILFx5knSbZYTifPXaN+4t8Kv1e8uSwUWL30wVBFO75K
bXUrI3dF9GUkINzpsTt2xjt/kUuoR27RW3LKinGbu8q0qGh8/ybuGaGg4T5knjJqem3UDzKmnwx7
zpK2/U3tuw4nWg4Ot+/obvq36riD+0xQnbqpHrHF1wJbkx7uvqd43P4Nxz/V93XFsYRSpk5QOnYW
Y8WQ1ZKsS4wJe3TIJtu4ncPe52AeEfrEQ7YPEHefrCibPTMJTboignlRbMzr6GvHJSD+ggxyeCmj
oxCs2MaIUJw3fXDh+oawclvscTwDoQduSSf6GoB9ylKO245MezEhCl7qULPhNQcDKX0MLp4tQME+
6SEUGtL1Pzxmpgl0h9v8fjFd2xE3n7e4MbBFq4oR0+5bUb8l/FIkSpQ2r6sb2mUqyOSjhBcapTHD
VcGzKTrQiL1ItckXtaGzdlyC9r51ISIAS/tfmgEsqwyIGpsqN1PRrLfusUiUORjadOkyznWVpDE1
m2LM8tjGNFox8djRmU7LxXjDQVxk8LHvSrXeG2wOIICRYwRrv6RFPFueoqrhKmNGdrFUN/6ypVLt
awxxGYw3ZPUav32ppUGgsQA/BkXLzBFMuFBvDZUyJ8XGYfoJqzdW80HZR0umPvy8o52teQAyy/ET
mR+UF7dZRka+KFz6ClxiH6wmhpB4FF9H4nlo5Obt/+6Q4YJMWfA1q+SOMweKWxQEPCvotSK7m8G5
dXxTs8GNGdHS2Uj/Rua/Gzq5j0HDRyW2T67bDCb6OQRDn5uqi2JjW9f5qR5AaNTPlA/x5sqgC6Oh
05Q7d0XEDpOoULhRYaERD6oZMpp6u08HDiS8pgyTyDmep7RRtoNE4/P14OjlPhdoPtaoQ7mzMH1C
4eTD8BiSK+nwTVAARb0AnWFNw0i00az/NzgNHDWiaB/5+GrQ35couoSpZUXZlAfxbzpdbcJ4F1cO
tlhBs0IqBjRku8LIw2nsvrZBZP6cPJeKCy4kUdon3pOAxrjUInwHAiQOV7+vBrQOFANsMFfZrzX6
jle2cSRodRAulzmbdLdcjx9T6TLiVCJpENYNfPk/uNUV8/54hruBkgxkdBcd1/ZCwl8j/KbtfznO
EAK8LrG5ziIPr8NX4jxxutBTOG/o4iMQwEUdISR889N+gp2MSfx+UnhF4SvjzfU0GJ/FntXM/Gdj
3+vZdRJGGixLKglPnTYNcoUrrQ7ndW5yeX/gL3zug3IDeJ9RxdEnFHOF1GQbn92aPOivyuioI721
uMB9Rh4xzgsuA0bGb00FhugHWv6k9l1u1b/G4OZKcPn09Qev8LFSO7BYr0DLrnomRS27ON3UgMkF
vPnDbQmHYwD5JgrXShDxmrNKT5Va+4gGBFG3vNqCUtE1B8EkGHKeAjv9baVVVUOLlelZfVB1MA2E
wxrxwHmoWf1Xbjj1iqEdOD81WLmpkWOh1iao5r4OHOaR4k1LYEc7zqNuCxIMmvKyxd8TPaSh7X7g
S024/aRUor1g/p0WeSfzuHvkTdpVDUtg90G+hZaeTPIcHcrpG9NhpO/t/NVESEtdXGvFRvK6jfTX
LzZXw92ly43wrqAkdnZ1Mrl+g/NOx22xRv+VF7Q1DCPFPh9tnjK0KHBqprnRB17UzdCe+q9RWsWg
Jo9YLVWwnRstqv4Bo03/+HqHELgPaoCLriVjzLrhrnc36CdFCPYaVNnoozl4CkW9taeqA2sKnCjw
OJzuwjlcNAMxdHXfr4kZKK3CnmCrRzPLe5tBr7ROtPwYACoEarHdtruAQFkjEiKGS76UwNEoGK/a
jeF1maIdYJdNw82Xmvah/OppPbgs9xL4LbteeodfN1zCBtUhjvxz7NKfLKCnI9HJv0q180j4a6+h
BntvSfpUc4CsJwAnV7eYvy1AzUdXn5n4rXLZF7Ftb6m3H9oJCiEiDIwvCcSGTGWEJqq1dbafTQ+y
7HNvGCWzmqMLVP9m4a8nzCHGO3YncN8dYFFJ40iLKZAcXMNC6TkzwmPaTVql+MMRN0rZ0+rtrReo
B2QjTKvnqg7FU1mcTHDk9dg0SgVBBEGetr9B08S3w8cPls9kb/ZHGXihAzNZaZdL2zAVPn7dshpk
aIhnNCBNfuMeSY7YMzIeX1XXU5LmdpqPTpyqSh9Y/HewLBPa+ZQYUxl6QqW6cCffoL/lllg/Rjpb
7gkpDNRINFueqX2auY6W6F+EsVLE0JdA5yNHMxDJnyZPyTkiX+9GV4OCAuqeVdkwAOxnG1AEdKNa
Tb2sN0bqzRFQHKj+hov1bIA6qgId3wKCLEh8xPTnczlelM+JA2KiEdLEwWVBlYOTARapQ08qLpej
9LTBUixwLAil5pFrur1gfYcN2ANQ2uqdHKMb3BlRhQTRQQ/Tz0zY5UUgk6YJ7FmmH9VQUBkBSGBI
6hWY9rZfMRvNqkX0GqCoSr7Gl9tiISXo+NychZq/vG2dKTMFkj7g06L81gmKlAV766OEJq7Tb7M1
8ACt7ypQKqv3J7hmsfPpow3hR7Or8h+H+VHZe8GkVAhfkl+5KdBBCiOqaCGLPpmVnxkjBORG1tm2
90BqP/NLWl/4lANHNcC7bRghHvXxgXXONyWtOE9cX9S+Kvma0UaskKSp/Vo4mU8phNmi4vZnmPOB
karPmpEb3qD3t5WsD1Ajsa0w1mrYhO97ki/mqE9l/6qOqh+mbxEjKwKf/O6oGzy/LWSAObxCfBBx
dQpu1oOj0UgpTu+BVkO0Hcx/xR9jRwncHOncCbS+O1fh1aBbCJITqNBbTZeRSujU7Mu+JE/NCrUl
R6sfoaz+5v7kQa2dcPDXhQSMA9Eqg1uG48aSmvOUy86azNBCeHT+K7qhccE9ylSEAFdAr+knKvbx
4W7+rmcTJ8XOvtuzD+kfh0h434a2vjBS3lNIpsYPLWKxL8qf0kR/ss0VnW26wVoOsIef6gQSaFfD
n6IFHbaYdw2J0i2b3rLAStXSQxS11kGGKljh+yJ9JztOpITueVrqE9vVEQ85SiejhuFkIPtMf4h4
fIWnhO/kCZQ3+dYNKJCZwRwb/8Lu2CKmNaelmex0HitcYaNO1ZUSJ4c7aVIvbhjrapEDV0RZbwHe
mg9ffFiL7nCVv7dq0oC/5Bwr3Ci0/ILsEM9DbHGk9VetdXwXczUqaQEmr144qSZEmiWp4Ssprwo4
tYNQRsMq2lEw83I+vAcIK2MVRX6C165yiMocw4WDJ8lqI1TlNxLodkKcmRQeECxyjA8ky+7S/aiv
2uTnnw1vuaeoz7rAJBkwyKMl+moSldluuxy/TaDXSy6ndirXzKRAUdOFxHGmtzhnoGlrwXsVyjjS
uWje4ORv/VGwavKaVYOKEwVDB3aBjOL/SAVSXUL9KfuajjrvOGDLLW+MISKyhAJEaxB8YgKpw89l
kp4ICcdAvKxZJZmoMiMCJOu+zuUwpOTokAGMFEBtMHT7wznIjG8+Z27MVEYlEYHT3Wac2hK4t0kk
Dh13TC/i4QvS4ozmtqMpV86MiibSJ4bC7hgxDSoM7XZ1IKDUkiEkeNwN8fW9EU3DYLh5Q+R/Dkvn
4sX2ZMpxcPLvXC/fg0eyRko7cw5es9RjFCkegDtqw7xrhsQ23La47DrkQx2CIjRvYEKYrvHYh5o4
BtjWpVVywWz2ZOKCs9hoBhJX80PN+xeVuPaOWUTXR502nj/vSWki25/qEO0KXa0tsfkLfOV9mfjg
rqVbHgeossqKZii/JO5OiwtVMjczFwifaTgiwaYLv8xwaN/HHy5fiINkZKfIkCU/1PZ3UH0w5e2m
AsrFXGGoUAwCDpo+xv/CoUIC+7reNBnubd2vrNQmT3douogU0Kbwcs+BHOhdu0AWPlmkD1dIDkXt
SLVs8OJaOHNIgu3O90kNU3Qd9yP1MV3gZB69aarc9/CtDLwl2bg5AdIMbu0zpcmm9EuogBJPsK+B
Qs4DMpJyzQ0vS5R9EP+uD4P0W7p+k48+8ajL17oF/+oieOHXHFQDRcEN1EXNAOFsan43eWdrhOX+
gLkaribgaMR1WyQIUAqQuregWjO2SjM70QQ/BALXr9ibdwG9F8FuKdzncq7gIbQZMtmocjqcBq1H
1P/BDa9xdZtJqZqbztxCPLtpwmYxyk4RBVkAb3bhjZQD7XJ9wMBYgB/RiJz2TEtCqamcM6Zs5Apt
TL8n4q7na09+hlhRFaAl12gMxeUUxTzA/MRq5eZyuRs2OHR3wWEixWQW6jqnerlFjSrpzeDIARv/
rWkrAOBNSr6qsU2iVxysioG/h7cHXXNFVYHtiGKNsYi9VcVvjwJzDJhUuVT5F66JtSYqBYu+ehFQ
shHHPhAbYH2WJFmuv1TSW9O22V6WncIJjMlSPu8nq8c3WffvO/Mgw2uBAx+CF+tBPRRtgZUGxXXq
qR9d2mg+s4E8gpgH+Kj4WZlugiQdXkbZGw/3gpC5mc3dasAuw+aP6uMdrzwnUEHvh8zRQ1j+nxPj
15nV28zCwCnAE8mqGuKEfQXIPo+xv27Xe/PbyRKUmqrxyWlZB4zVih1h+76l1mG3sQPgO0ZYWAOv
UEHM+KcxubjcPsGEfQdlJ28vEPy/ykOJ6zHX3EjiYcQg/OhhjnUUDVl/8W0skQB6roOCLdwpurzr
G0HzJp8wcJEPg8DeOx157C5cgv6uwSalBX5BQBVJ291rSjkD01581mS3jWRg0yv6tUSvoz3yG4zF
2CL/74wOoTbqwBWk5/zXZ/dl2hj/1m7jhFf6q9+eoN8ldbxedSIaTXHFFwqz5Td/4awlU1a4XiH1
X2B5VNv6G0mdQh4qPUzPMFV6tv0uxRoAZZvkrU7B1E0j0JDuXze2dNeSSR5MBBPHqFXdWBG7JnHt
hDcsxYPaXpnwVej09fUf3X5hQs2pxur7egvC0PpOpONz9INaTod+AMLr5tN8d7tgHj+blY1q3df/
xfBelUhxLkRGBrqE2B4d5HxAqOdBvbVLgEy1uoQzIqnvo0zd2eS/851lmptIHft3zou5Sv2cCXwP
5S8PTxJcBK4AYtpi5p0AgmSV2+Aa/3FZAdh3FVdpNkc0dWQk5dAeCqzf2v99Ksz5cjnH7mbTk13j
sxQ1Lz6JtRwKVnMiTrT0hvvbd//Jp5B344wdaxW4IO2O/gjDpbPnffrrp4MFv3C/VunopDso7p5n
K+NBjJ1N/GY8lqbm5EpXrohSpIj/uemDYIu5B8IIFK3r4uypDQhkYNzr9+WQQIeQwPPMeM2UEkLd
hCHVt7gqPf9O+EXbOtJbZtnV6NrP8kPP0/7pPNAf3HXB6WloYAiOUhtuqKKF8KgN78xBjOjFPrmw
YT7eQ3lHjWELxDuPEmK5aa6ggdG0vXbMmjXXlENX+isXBkFz4MF06x/komQPFaAq6O/bBTHwoef8
Pm/sjfQVvNSA+9G37pI3yoFN8DhqT8VQsuGFArW7Y95i+3oLuVw8v5cjglui2X001ApBHY8xJzeK
pqXHKUQsS9p3/weRza9mUvWqHQyEC+cOo/m5iwMnNN3uGggtOguCLyYNiolbJ4QNuqlwqctRgBt+
EAT6orkHNF2eZjCcwNxbJacIRlBqWXLGPgbQEepgcrh6WqGmodjjMXDFYQsw/zYfyhsA3DN3oSok
hv/bkQ5ukGcAqJq8EZ7LFd6i5lxrk1SshcVu3wTmkKeNLTR1nspvn3wituRvtMmLRALz2MDTZbtM
n1R8Ir3Ksjd3tyrN0zadL4FBeEEq8Aq2/AG1zwq0RCIFfUCjiG9azjJXXOOUnQ2R8oR+QhOA1Vc9
r6j65Kx/4oYzQNvazIwatom5+xZlj8g4fik3btYSjKFHhtUqlfwImOiWM5fuiO/pG/bPgAVp4Ms1
MFngwTnpECsz66B9j79i5JeNjwlNx1VMHwcZDYOOzeamJ7eaiyKnvJ7mwwVhg16fqNEehnGZuD13
tZe7teFcLi12kOut95uFy36QOwoMQDlYbN+bLHXLmYuQxId9qxoDcPm8CxWzzaWJGB7d3a2CSvK4
QLhIWxpE5K76OCQKP0uTWWszm1EowAungw5GPCMt/UHp4t+CG9Osrc5IIVF2E5RTbQg1367bq9RH
w2YX5KPYq8p9o5V0j/sDLRs+Xd8lCr7RGAQDL+rJ1OBIhStvoy2MsWgY9wd4TLfm7A0UnwqSvmiy
9+8EjgOEyI3jxCOItyD7YRWD2CVFyopOgOwfNqo6dqtU1jHwzS+nnB+0MDCnZsX3simlbpVvKAQb
aruboL8B6aEEmmqeixiZUfHNPOJHf4xDSoIBMIcHudnz7m4R5QPrdIudMxijtUq3K0kJo4PqCnqR
ThAMUsFu0dLM290iPimd1MaAgl/RRNX+d8htgG3/3ngGcHP31p04KFw9FpMEt6Z7npecAUCOZc2O
2+92/t7e0hpvcTCrfpbMOfBadxf00c2Ck5x6yiZOLc28QQccePs7ivhPea3qPfSeOYJBygMpd8Zd
eZOrNVfOFzgA2PkTHKGYe74fvKnvshn/nfBBFLksGzastP1FAtDyTUYJPbC/CHLXvCO1gHMrcQkt
p+6As4iOsB5OfF9PncdFxS2KmasWIjq7OY/xTK4ZM0fIJicQPzhceMWFfZkrDYNDOhmKKk186YY1
pWqZS+ZPvKKWEzXUCwSo9VpMbYtwEZwa1SqXQNCnbXOrqg6UgoTzD+36O/JHwmS6UXa5IfhvJt3r
/ixOFjSPDg7f8aPiZjEHIDZhX1KqvVLG5s+F2eeKWh6YR3qr17phgqVxaHvoN5LM3P5l70Ez5EpP
oa12HapQaGZZFbeRzV2k6LcV3TPrkBC6Ok1Jwdk6jV8PsTojJcCKvfkK294RUrygBw8DzN4/M9xM
e64PLoKAfU4azIH9/Y+v8F1OHl8FDXEcjqYPG5AJQXoHunVCwzOtnEvsFiWsA7oTCd+4s2icfq1i
XEPTDZoJGZ3N5knOXMNYxaipCJ/orlHakqwas9NPmdFSlPCIXNDL3+GaIC/b0ARwhNsEi2G2s/M+
2Qt7+LBtOBMPLx7ktuY/inPom76qMho5AvrCJgOny4OqQJDusfDLTycIbqcFC0fBp/TePJermrQq
A53slhWBR5pIs0GAQip8HqT91rn8iO6jD9MfSXXapvAZ+qL7+bkhlr/rTNkYEsTHiozsg9tRp8wB
PPHagOqVLT5761j91TaXtXYno3voUYrAmj7CSupxm6eWFWlU882JHIaW6cKMTvsmpnROYZzwa8Fp
m2apibquUy186xichpXE5RzSCdYkZ54kbG0/c+yU0JG7Ka+YzaDblYLKkvwGbbt+AbdVgTmyGUsT
PQ1tY4nURlK6ajusd0+uAwpjlEomHhnf+w+WbFmC6vACBT7umpN7c9jUblEfikUknFFqb8BYaTAf
eaDOiHw3RxOE91ddeE0wWJcwSlao9HVt//vxepVcW8ouPlPffrkKz1vG/5BMDgG0O+H7pYHkXLZg
CQVglVvvbbW1kb7531E65Fg9e3RFaTxab1UUj5hgKZ8xNcS2fIeuHu7AxUJCzBQoRwtRUa9nh4+0
+IFntN5oPyWV1kO1PawpWZxypiiRThBLtwZmgrEhlFvAWwmapgOMRqCdhEr0+JfeDXz4gPYEv+bz
/+mRpn9gq/zCZpG4ShudSuH9DyEVqSzcUZnTH5Xr6pjlRXoyNB0qqePTLBpbcj7pegeRwLs4cfzz
H5YSChWqGcqPk0+kkMJOT/rKkmL9LfmKy3zcSmuk6hWZycQSOicyIa15B2soXp889g+TPWSW6+kM
Fh8Oo4QANNMK+Uq1ntQ/VU819ZyFMkqxq0QvX0n56zvYlRoMnKfx2ENpG+OSRhWtjlzzKYRHMd1u
HJGxns1iVPSqY0L7Y43uLPewAtMIpwPWJQ+mgkIpWjL4ER4Pgaaw9K64r/89Rfwp+7bifD7NRB34
Tgaz3r+MvlxkAXCESXKij6x9fq95s8ItPx4Pu+EnOt8iWRUMic5/Sdx92h2KC0gpYtvinC8OUPjK
5ZVy0JWDT/IBLw195Byr2q1QO74ZiwcQcWNihhfEGYlYWuUfm0bDgeAWYiRdvwwqm4TNStFUyIRk
RCqCzu3Adbfdi4aRHkid7MYcipq8GR05ixA7I+iI98+u+SCSks6weVxG3fheB4stRVGNA5EJVKI7
cDvPXJRx/mSw6Mc+Q7FZLIZaR4WPgbIPDC5roPFQn7BPys1BtVAaZb2j05lojAiFckG/QhmZJiJr
vYMqssfh20iswRWzt8UgQat5LIw67QVu99BVU71o7zP9tp3YE03mQ0VIVzq41ChyXb6DczNx2gUa
EFjhs9GtO+H2jQzGsWtH/YyCfcdIg37YRCKA3b3ZggbCKV6y8qcPOermWEZLoKv4Plz/Sekib64P
vzZ1OrZ6OPRkA/GGKgERIN9kdP7dSRP5rD+YyeZH4zSKM6K837m/wHcW5gGVn/frOxK96ZZR5D3G
78mG7ObcEwf1dp/9BIA8vRgfIEdN4ypU1KyenvA+naBCFfbPCPFTuYtNBXq3p1FnU45oZ2q4BUGn
xLS0/k2qYh1UsZjXHvfqEKvWFxXwX8clVI2oVSVNowWf0KvgSMq42EKTH4sk1ypHCFbVyU3XQCLy
kjKezqq4nW1t336zDQUl690FUQGZTpD4YnSjXBA/qsm14keb2gWGOEeYkcGAqMd7sHWI972vgkG7
fcvlvuRNlJI6g9Hg5PMRoH6AOhyQELKfZNwgqBmPGgryN01h25RvbqD2/6DKrn2qsjLnEy1GfyvJ
LAoL5ZeQLh2IqAJvvXtlnnkjuA6vMye4XfWHjxG0IIn7G7T/CIte8RrBoI64ReCNrEOPJO87NI96
X2A4fULMHOy86997/B6/5lKMLS6RhwtfExpqS4J5DfGjU4AO2YLoghstHafGxr1Gb6QZQH9oEpnp
TCSO4Mfvw0sLRu9iuvuvZvF96u/qK6BGn1wDIZjI5wmxCFna4BwOasTWQNl2OugKeEd7/qO9Ag2Z
aYQqwKiDjp5p9CPFj2IpGew0pp4hiVHeChGFKRXTFu9fOsLf91I0o7dOIe5yY3+Y44i5aXZ/zr8x
GIkd1sM4LZD8tjQqXDpyxCRI82NAazmH1Pe/rGCRpTO1wq7Rhyhb2KIP8TKDOVl9IfIOSOHWh2bp
muAixVFlUDoHgigfVgQH1VkOaVlZZOQunmfpzkpdSF06cgFZ8PRjO79O/PaFrLqBEBTJObZrFR8f
bpKf8t1oq2nP3AUQX2SEsaXYS00fbiFoj2RhA4nOREQ9LxUJ0oZQvdBJtI2U1iylF22ML8DAn1CA
2EZWT4nZOMjDuNKIkOAPJECrPbp8e6znjj5TLIMuBFHp5CF6QfVcO22ZJon3Ktlbq7piG6GsGh4V
d+tau0p0gW7imk+FAmAJQ53wyqexv7OOAZYCppZmvR6sZX1vJdnk0Ww0tbmRu2v7uJTU/Wvh1L4L
B2TdGrkafoO4Yqwmse5DCWzyRAY+3Kbeq125grIKqQ14tC4E7ITKCP7HZstsbFByef/LGtN5+zIk
NihOSCaEDH00cZtqZZ935srAlow+uk+8CkomvxQvNoi25QddYN78fBhQmQgGVhp+9Pjvoktw5i28
5RCGf5R4F8AoxEVFDwc9oij2AGTOWbxbZK4akgCzJ5kNhqYnEAXltwgziBxzgXBAnabBOHe1Iggn
uRV/n5xlaxYNsHyfOqdQdsWsNuyivlETm9huhwkUXj9+Fv4UJpgh3ZcgpYU+1+r1tti8ZlPnsa0N
6skeaUtE9JDwWFZVYeSijTVOZyD9ndDorG3GNVnqhPadvEyhLl6wbfKGsBL2tlmMeLc2kNsVfwzs
QTtHBuNzmLYlVy3FRvdZunrgL4kUYwbub7hIvD6L+t8hqeuD5wZz1ELivvlvzPCPALauf/rGhYXB
lXJs0gc+kfUzBH06t/GQpxKVfvfgRTuuxerEG2Wtn0JmZQegddwmZqkvguLlLLm7qPVlVFdY1MkY
s+0xWYu8IAPn49z+BGBAICKxzyXIrZTKfOMnIDV6sP+6xmbi3jvakRPyOlj+qGVTqRuGOG0qOzEl
Xbx5yLyBJLwA+mmKb5UZOhHICNxaGPHrTT1apTEks0hUVgnuZTfggbIruzU+q+NuZZjqs8pw1wnj
sSbb2N0v5E3eDnSVyQaluH9/tQxyeoLuUO0m/FDuK68fLomr3OI3WF6wivRNciTVAxlwcMknBXnQ
cdSWkKGdQqXgWR046HSAFqz00vJXjKNw/QT0wed3y6QgJ/HobgJuOIo1qWxk/6uIWlc9YG8H/5/t
J/jUxel1QGNXRWYQ3d9HVwCsjSk2RtcwOfSTHqwyNsJbe7vE93tVjG2MGMtP9ndhKBNVhVCg5a7X
gVek95Hyg1BTFKt0yDZme9TZX5NTe5Ln+TSD4qjGSla2hdSyxu4GPlSjHO9ldqRlcai/334g0Afb
Erxf/eBfNMK8+gnPHFPZ/+tAQzS/ODH97rlGCpwvyKVEmNsydDqhO9+0v7bhW+LP+HWTyxiLSRDt
r5V0K4B+WGHK9ZuraLh511FsNOqSXQElYDnbga+Ckc5J2D5ZbFngAij5rmsyC8l8K23hBOcNiKUw
RTv/0S0kBter2H1aDK/W9FEb926TnPbTaxFtNchgqU2HMnfsHkPcdCVxJz7AKNJ3I4raXLVU5D6h
FK2du1owNd9jjEu/r429HdPczulKb0NJ7ED7TgM/3BgfGqoBd/syG3Evf9Q6JPDHpomwk7VVse+r
p+qLfLVkiwgj0hOCa5TeMczLdMy8R306fSvDAHkV1m7wecnVHa6/JrOCBEJEtNBg4oCgof9bPYwl
Nv64U+j6aBI/YJFuD9mrG9V+EY5g5dfMIJ/dkzUpaBa8Re1xt2BY/hgxr6c1kaIL9i4pe2ZkyrCx
+EBVUp8E3X8WhTI8g0sr0GpmWH8+wLIoK96jFQtlj6d2M539DklAYDuOfH9GwsG7MI/bZrkA/qPJ
EfPJ+Q6R+bNao4c/g1hjTzqxU+udR+gPubvoVxFuZ8aoPL5yOOZflhkv82MIAI1RcsZIwBg4KYun
d/K9xwT2uQDGI2lOrVOwZz7tIB39197tR3QwhQ1lw2z7xsqEyvU6YROhNtXpW7xrJc/gMDEiuaCy
RBoUeW3RkzhQLtQH1caKRjf7rPCTbbnLuMdxVy/mfChRQDCv69wriK3Vf5QbnrAovLDCWrul129m
7ZGhUUSmBjr7wZoKbpZCm1vLz5ZLWWwLgtsZwhloQ5vsZoIjeXXDWTgxKnXYCO4a5NhCNNup7LjF
Qdcrw5bBo7wnhVkeaeEi8sMfJcwtEp1yiTDO2o8Sn37rV75QYNLMg7viQFPJOovLh8TUkHmlzoBU
gKzzFhjdnDWkTQNtQuyTRT+FaZJGYsV/601ON/3KOv+Ag7zvGwsGUJtoCncHTsv73kEKXGROjTrG
B6S/q8uz+RYiaNfvw85sibpMw1jpRU5gIA29Tuc9KXhrKbzxnoyxq1tevE/ZAN9o72wXN9uGFt8d
QmysS7eS4SzWxxYWUm71yydskIk/1XbQ5k36ZDrKLJOf5YYZa4S2e0N4V6ipqlw+XGCzfUzmRNlS
ojk/uAtb8MDDqfB+Br/jFbnCoQ8MyLiZrzYTOAG9LM6NYcTWzntCQYT4/Elr13nF+Hnm6K1jN/hO
idWhuCM000Cxh1r6ZFaNcY03P8ZX8xeM8Uez+KKAHRgnuc+jGSXXqS1R/67AM96y7ZgkE2RHlSB3
6WFqcObJkrzO34GJxs/+EUgg/1wXHNH5rLdeSyGUkBbTazy/knHjo532dJ5Wqgx93H5PRRGQYllU
IkUpXAJhTUQ6al3dweOo8gtbCYMY+anSAi9IB/xUOml3DSw75KaSp45wZcX1KGwNq+LjGf/qn4Qc
YqDELgE+lj5aqoRjnvZiUbKuJejLQFjAlo9XC+/1XgPQnH8Ov3OwV8U9yngt8xe6ijcFtDsLdLDR
A0fB5r2SE7T3xV+aSRdKDivIPbkujvDD2EY2rmGy+HVv9xT5PQx94/6VFpxxZMCfU4Cec58ze4l2
S5Rk9FZaG+oiBgDZsXG5M0GN8wW0DxQQ/QZNUKfOU+NZRPF/4tDwJ6qhN0T9Ls+HaRXza2agdNj8
miIbXbFS4ePrYVfg2BwsxEzaLJzG25LBLf6+zZhvxO7M8rP3O6y3ETzpMEmVEKqUD3b+0Q3Rkk4G
gzeLKPh+zEkvdLp1hPEOO2eV7C7f+24d54Y/n9ZQ019eRkBu9EbmisgwM5xr40SUcFALW1WZSq73
A5VuOLDZX2LbmSeh5BSLfRkg0NazMfIKFxbI8CbovZmLoaoYpZ1TU8EqLFNsJPCu1X+q/S1uLw4S
RuZB3K36neaHdzz6q5ft2U1Tmyb9s9WfIIQpmoW5fgJfKNdvdaYUg01+xPA/utYJ99Ad9IFQetzc
9kCcenX4lPhg6qdq6nJrqujK2dIMEAKiyBbEO+J83BPJe/acOR193jOe0zBdDq4OBcZB7V1AV4M6
BXbJrwqW3tXgZF0/v9jIZdGeF64akQkLfn5p2g95lbkLw3/VZfyIwuizeyMqPoqYHJco7G/Yw2A2
XThd89RNPYbffLy/lFrVMX8WSQ+l/cX1r6BQ0le0E0XecOYabJ9Q5tr1FNitdULwaOVm15TXEEQe
qc/6gJoTmiF6jPYZr0wE+TxH1KyKl5LHtRMN0T16KRYUIzBPpI2XzAL4iZzRRbhuTd9CVXk+DwWR
R0wHZrmdvPGW8rH8E2U4zzprL75N6xUHy3W0o5Ymwp5S42qIvLqLgMUAzmnm6j49LDlw5tMiKdj5
0H4fk9Yd8Ok2ItbyulHja0UNv9UEDljTpML4VcLM2TIyDEY1AV9j8UOosOvXgL3WV49vA82u4GZD
vuC9Wb2XmH6zB50CBshmmwPA7LW3eog+v464oVTsxdg6RtcFu411sKzWVN/WISa1FuXtMzNjZ0tb
kQqI8Qa1Ol+njieiNrDeqVa2gpg9e0M2Mar/7IN0zT69bARdXgc7UAw/fRZtVYxIKBe0Uaaxne+g
NVacsu/NYNYhN+sUjDD+APPxQ6AK95oKHgINOYUrnzSGnszSfHboqzJ/IBihUZfFWdXZo/KMBRkj
V/MU5OLqpgQ9LbYHluF03HXx3dYRKXThYL+Xnf8AKBIJqEnrsVBb6zwD211tgkPAQiNm8q9SAdRd
HI9xj7o+i0qiUpubUzClNLtqonaG0IeHpzRJBboXN0oBn3zGtJyhyxptjf6huAahC3GKmTlz0vJk
xSkUOC8/nyw3n/CC56AwVGRj0/z8OVog5k9xEiCciC1pXgbq75qQqFDCWELVjM8R+JcNXEPSQdjJ
YpaqdpSqJKKp870qDpu424csTEAR0Q1w0/ujq03ZIcpE3aQAIAZ2vzt7lF1aI74DGr3oNUXkh073
faTsoKO8D9Not6QSLBxaZP20lzL+606oqMUoLNKxJflgYyUxzVjJ0TAIyaNidgIBnFuGlLN4LtLe
Jx5W0sBE3yNWm487JzTCNibBs72YK7vkA1MVRfcARQU/Wgl0CvdcDpSgVSzwDJGgabnj1OG0rYxk
jXgJT7NORI2+ttiSapNIIVsqOicKebe/TX/N/JnkSdAh5boke9LIDRZRiOeF4MV2Kt+QYuUVCw/E
02CRx+FoBbwkempN9yK46kUqwXBbvkv+XytPw8A10LnGEYCWvT0oWyYVw4w5o9oDqboi5Ez9/2qu
sxj25f569C2C6Bm5RdPAKta4th3hMQqk8mmb0rsfrRg7d2yADPhgPrFjNUf8rL6da1yyKEzgAGuv
oTzoKLdqhzYMxPiE+FGs5wAiXcrPoTg9x8CkJVjOMXAA2FnN0V0O5X2QDHXesXkv0sfoVv4JrpoG
aCh8R5FcqvpgyHN78F7v4KOuHhSJQPBhjHzeLK1bDRLmhsj9GQIXitS9UOz5fI3o/uLSoVvfkOWx
dJqe9sCfw54qKiGJZ8JSd3r+9SeTJxMbO6Ig7rO7WM6ZWh0ceURJKBM1n4pSrukhKK/u68D1d230
e/blGBb+tJ7TdnYnbmhrXsAKJv/LBY+KzMJAkf/Z2SZqy/kcLs2Qk9uriT8iTcCprb1HM9cULV6C
0SZZFPiGhULaSGqvSt5kp9+cXtQqv/tKYUtbMc8NOCwf+qqKKGpxyVbNl+8dmGgauYVqz5d5yE/r
ouEsA+JBaI1CETfjFfwMkA1MDO/dSXVazsckMRFF4f+A1MRGf27BbQ2n/0SR+q6+sOBzkjN8NeKG
ux683vVjeWQgTlEjAVIeCH5WNorS0oBUFxKz/DsWzWJ/Yhr8Od2hhZaHc9ASfW7LWtmJ1aoEexS1
Aka8L/T1m6QyXje9K/xwNy1rbSypjZlrQSu5q4bDWn0YSQeuY81u5QzbfmE7TCWgLDcX1TkUGCDx
TDZdqC+3qy+Bv+n3ZhmYUqYDyjQkVUu7nD0eVZJ2qx6dYWFYzsd0pIxs+I9+J2+fJS+3zDGeF3hM
HE3Voh3TSDUxm+ssT6dMFSBaeEEsWXKhsUKX8Q86dzYAHWaZzdUfWRIEVAhkKcqkymEVy6nY3vL6
2tdKz9wUj31ur0H5jhsY71t66nWFjjeTjzMiVHK7+FUgSx+MTfXDgtCwn1sDpsi2uuEfVzt9su50
XuAC+Ubfv4a+nwtBzakV8I81wsS0XGlz0FjllkFh6j58AC5sIa7ZC03ypLqHagfZnOpOE/t5U2ei
mBEg5Zgd9dSjSu0qfImREUAfsOaPAstXaFKb4VWGFCAXkZETwP02Z1tC4Rmfw8p4EKOLns9qACMe
t+sW5BTOeHBqse7PDXEubptWqfO8ievJz4uvjUGZQmZU9nqjxrK0UFXi5BAyXwgQ9Kbt4M8WyvKj
86C9o33gJMp3LVw1BvDiSSsk0Ic63QMYAOSQjLln59hS8zgsX40tbPOcfhujChJx44mLpcbfY4+u
oKVyWdU+JquRpXtlRBLiv6k2kQwooo47GiEi0HzP9XKUpXSEoljuYhGj+Vd9GJigj3f8q7QsnrxS
4DNTessmgDb4pfZ/PFWu+ANxCOiw7b4pMGo77SDPW8kNI2LqeXr7IUWY5Jjq7jz5IHKSGdsIOWec
XnpZ7zIq6ByAPjiB8hZHvK2iSygo+ie3PxGQFSUtTc5dkGq+EHMOZRtHR7AXo6SUKpvKJsWBvoh+
qY7DzAiIq1hFcRAAPzYkgjGIBlR5rOrV7+18BniLUFvZMiKAsZxzQGGntTb1mCXXwgx9OwnHy+cQ
AJXKGcS1dTXWuV2A3PbhLyJNZaiMI4Z9zEycE+ATo1FieCG+qZpbFm7tcI6tybwMVYXlrYMCkXAo
mQRUDO7kv/UTIf7CYDLv9Tv3IZrjz1Tya0nw7Q622y/9gQ7dJZgD5Ilc9q4QqmrdjBRQASHLZUhj
v/fVET5lzsh6kGjRSZjHcgUzRhwmGBahRgoxynkrrW3k90XuEoDgdbWrLDmnCqB2lvcJhINOIyT1
5S13G6aRyJRoyv97tPTQRphBVLCAy26FyZDw/HiyF6J7o7daxFNlCDq23H71uKt0VMskebZGWUSW
Bu84v6KZ3CbRkahwX3hq2Rx69Uk1x+WaJ9LkGXs4hOOfvs3FRth1uIZHdYNVI9mCehTZ/LkgkKBL
ZiF2Rk8ff2nFC0g4/pbScF5mQTrBechLN24g56Y1e8YnSoWSwNsOmUhrHzXOiiGGyEBdRwtA7PwI
egLWtJJy+fJae8fbXKQy0wXj+vbA7dG8iYKjrdwxUownG03qf8QxdJ02szdmB32/4EDP9qW4RdCT
YxMS7I5B+srTS5r7ZrBhYAPURaCkneMauvEE0SyCulLCoGRYXFOgbVSQEbKcrAm1dKpw7lDOkueE
Ov67fmGn/TdWLC8qZzBsskPwqiTTXydFvoT/39RsmRJQmXhF4SAo8XWcMfqil2uyHw0lqPPXB3yA
+EkF0jg7uRxXE+mKdzIzjwHehOPCkfzkdeLV3MSI1Y2M60KgEshZ9tbuWFU8iNCcsUfwNQ3f/YGc
X9JpOf3pn5UNg9edY/yeXZywKwozV8an9yn+5g16/5uB/h27VMaCwBxjEMJs5OndCfpr5He7jIAP
FzxMJ4PNTPhSwT4xsbAh0aLgKETDMcJ10SdbhbMKyKHMuRhGjMM4If+5NvmTV3PbT/ita2I8hqYw
1A+BNPIbDmHp3Pt7spUnIHjchDbj25ShmTsg+/EI9TNv3MO/R8e6dTy5U+6T+TlPhQuLQr0UewIm
BBNavG2GyMvQfhxMWhX9ef3wxqpAVwlmgc6kqnldElOIllmj19TH5xrRX0lbLz72kaN6kwUr89Yu
4oqezfRfXaroX23Oz7KLgpMAcxHv/3d+x+jKj735Z9zewziJhH9HsYkIF/hW3uJEjFyhYCDVD9Jp
PLRCC/W8p8R3VVofsV/Idy9a9na7jvcX7MFsrOK7YJf5XQJ9QZpVu4ajmGMtXOPiORm5DamVf8u4
XrPg7i0GfGpCSIY9J9r9wgmFfBFmLUZ7Ln7LGOMQbWy7rBQXXoeGMWSLb5fCU76j9oEuqJx+sCHm
cj7RhwDKpt0vkcvMwhJ/w5rZGqDSMOn1KwuumOxCox5BGmznoJCmk/xVGwIx1wmpOs0ZDepEpCNf
09yXKSupzo/ZS/J9maTJKHlofnum/2ru4kxvjOWzveulFJX7a9zthoGnyKnHBU6zas+eU9xKwNNu
ApPpNVt+Vux/uwV8uip9zOznYMVzbUf9XKz9nGJCdpOPaJQou/ZIBNpg6jV3slTDrdB5htiODXE/
YAx1Wi1f6BgXdvqQc1x4HoqfLhpSPIEFO/vZA9eHMouvJOlELgo5Mr2AuYdEf6xcCkfb9NHzI3i8
i8GXXtOiQN1Y6SBE82GpZPknQBMCsbhEs8NwdE48sl8V9HAmYHX3Klkj/Rqp69AWTmwwnxEExNX0
g6GZo7nF7rZjKITmxbmfGgDJEJJQzkQZqb+SAgb52zEGnx5glu6rq82f/mFotFHESu2KumBFTwQi
0DoZAcNS40cUQNmlFsf/qukWw3qaX6yjyfoHhnfuovdQLNaIr8Tj1YOkMFD2ekhXCJrY4Jzno0l4
T0zSwr5SFoPp4L3sou3ScJYmvNmQdUYXDgA3E7yLxtDpiZWmBbM5aUD+vbThz6D8G14gjd6hNqi6
jSE7zOrFeoJhx+Woa0Ftn4DWtVU4/Az8ZSxBEfEtlJxtY6h9jfMa+dIcmeCobBEdrwvB2c3ddjTP
8fVZ0RkLckcz7ZWJ69p4im5SLJvRXSnm09sz3qx1mrnHiy2FO5HCdE4FNXcvAWSSVUEoHQ5UQmwe
NNGasqUyLPkMvC3LSJpIkSckES4dJSX+5/8G1dOJ0JIRiiscMKUzWSQZ62qyMfOl7+A1a6cu2idp
NqVK2FMiFxA44etNrvlRfG+n9CLaGLfH1gAaGdtEkNAtrmZCiQn0URPg0JVgxVCXV9MQkwqcnwZu
7dGZ4JYrfZiz44DNZIdpuvf+Pn97VuwjGBhsU7CZlH9WBzJkS1kXEmrbbtIunqVBaYa51j09X3Tc
XUN0mFKz2hcmU2/rSy3UdkJsBC0GXrzAWoWtcBfyl/Gk0dpev5es+f/mrHta26UM85XInBX0USrO
AHJ3iwHg4x3ib5t+uzCPIe+iw1psXJokwMNp2p5zaOuvuIesTqsCBdqjTH9XBU8FwrDUpjlzfMpt
bor+uyTEt0dErijCco3oxI2XoeZWO492BaNhHXqgzV8l+PoSaX3c11jB/PUER9kqCBp8w3NInFpT
dyjiq11itzqaLaCmUDEfEdB/HoB3OCNYboJAp+o8UtFQWo/8HfHh5CxKTWJ0pY+en+s/inT9pnqg
teHB8mEcG+gQXM6v+p67p6Hxr8aDYevwHnHY848RjsydKXx2Q5BtK7FqlDq6UjjwvAtM86EXg/2Z
iRDOwB/TlcNSaaXf8cCH5hufCqWY7hyESVe3YoDBfCV+cn4mLPbp2nem3Wnc3rk5f5Grc5xeQ4EV
xLqcLBvMbdRC2f4jx8ZnEWotZhUyygGjzqpQvDzQ64RHgzp2qIbeoKpg6UKy1qHsHfaN1aJJzXsd
dsrQb/bpkYAqkcE7qLLYEr8yfNR4+Yl4ymwBYOA1P4kFAoTqFqBq4SMeOhE92NdXJ305eCAzkmin
0VyW+De6XPNG0tYQ9SVTRQ6Vh9jp/YMQ6++9e24RjVMmlhekKyD8YESE4GUT4qWxPcHRSWxju1n6
D08FegaTMwUfnKuKX80j8XX+1sio6E2MWstXlZAeEWHrChY9Ed2H4LWpHrJc057gx6wixrBFbgA+
hf5JowP2thOJzoMunz4vKWap/9FfHfQYFN7HE3+wy1wOrrRllSyslCFbnt9KIsm8gvFeiOxkT1wY
tufhFd2w+SloMdvVzcIKGIW29suCFGroz97pJrzuVHghgahUG+Oy0w6L5khRBtbdzLrfeN1xigxU
JmyWRL7yRM4qO4rjorlYlXkPWEwtmuYwU1MwYl2to2Vi7+1FArUSN0au1WEvtsCfB5obnScXraxO
JmbPONoKUmStV5yKmYDxbGawRLcv5Xjqwr4/sNKFOy5oBB6QRsMnNddulsE1QQzNncPKSAaylR2D
tFwyq+Sv45Eh/WDDCaU4XfPu1cYGBQ167BDWI5bgA/Vi05yGzdUSkoDYeBsgoskNE4u+RUt3Fczr
3z97JgkuR0lFS9d2LfOyWnheaiKqzdo+1zWvZBTtocHAVBN/VG4almTXJaAzpt5Phk9tesXwg0Mi
FaVsKci6lhV84sQxDZzCOc++kLBnPpEtVnwdRCrtv1IPKp19t+qvx3bSIDnmYbY9qsptQDDQOhod
schLZInK5N7sCkxtP1OnxayXTkX59l79ICvWO4n9f/cCGyUw4nFY1RbsWTn5oTVO63Gp/GLVRJmn
u2Y7QYBSAdLQxwHLPQuKla7j2zL9Rwa1rKtBg51EGaAwBEhKFimUK1d68LiW2cMhzJAvOxYXnahj
KPtfSGVdTA7KosexLUzYvU94JIj7o7DqIN1AAI1HyKlhvh2ynQaaBQ+nMJDTDTnkP+WZs4VNJHBB
CQdcRP2VL4FBXRquUWgNm8KlVFSUVQjAp7pZzye0V/cKTtn7wcY96fwkuHm0I1++uYSFI3dHLiMN
e3Sz5w+mKDFS0PjZmu1EOk29uk2Vktv9t8P+gyVoVRKHG80JeeOrAi5hPRXtSNQE+eTPd7Y3NjHd
hxZCS8+3y7swhbtiqO+iF/xBm8M9j7NfA3b71SOHAOGRsmZ1M77osVGJoNM03oG5eNUoQOl4bhw3
XCEstAJmJH3+DprMlg6EhnQhquCGvyEGqEOvx6u5eyntQmm/4cd6jo18lkymfb6J7k7IBAXU8n51
qoxK5Qtasxf0+d7k2uUKK4AAaI8gYPGczyUB97rhXf5hi4Q7jU12nJvjxO+/RiVlfwSNkFQ8NW/w
UFkSUoUuyct4iv9hYPZDXxJd/nAiUn8BnWA8gqaZ9lhvobMZdqdK2Vc1j9pY8shFV0bTMnpbr7jT
QnZMQwtKLQdk7v+PvCFxU7msqWddbln/dw8XeC8NBH2AtsM/paMk8ZVS3tU4SdeY4bZBKT4i0leO
BjsrQGJcNVClIPcJ6srPij20EBdxnypFl3J2+4ZXPc7deE9CycEivM4sJi4OvC0ZLS5GC+/xJNyS
IRcCUx7c4HMFdNvgI8cP6ABXS2ar+yWxWMa0zvG2QuYkoyiuzV1/sfR8L7BkjmUa8RjKR+eb+2kt
wNlMAlGbTJutXZIPGCo8xRGxx5+pemhUE/ZX/597F7yZQP7zqopJZZTPnrtrQedTtP28XPIDXriB
CPx2GmKioZBb8tjMPml/nW5OpE80w7wLAYbj/d/RSiGSV9qsjRQlqCXUxwj2YqAVP+4514+NXq8Y
QXLn5pyjrvKZ7wg9+JwHVvBlHUNY2SumnlYi5l9BHJdWamBMtYcvsrIqx126SKjOatdSCi3R8QMJ
H+ShN1POf7FSy+kiGKO4YhV9iNZ0FWomV1GUCx5wKhnwnSqs4zqWbhqkRWK/NTX4+ywxC9C7R55Y
LHpq6aEc7bQYAqZrKLc58c3BwgyfpErepIZysxG9AnoaSSc2aBBt3nAo+Tlu8qv4J/zUXP79WCPo
zH0G3MHHogV1tvNJxtxBCO+799QJtI4K3JvkG9d4tB27kw6vpnvKsf/YWEaW+EI5LCE/OE2PsHQK
43lCI8+wzM+wR8yHBPDtWkBhek92s/MkkyMbgOVC0EJs+ANHsM350LXpHjLBJdXTAuwoum/pJH2g
HnVrtaTYgKgOnwRqvhECjtYVwYVR+VtdqGR+JSwvCESfRCvhwnghNDhY9K+7QyJhw9SUu8V2tNpY
TkvVZKCvHBY4KVKMjZ4iEGrMYpJMlwxmD/FSVrn4PEzW3OtNM+Ze2cobFRwaSPtgpJ9yU8tlQFkE
1lVv7IlY7OpK8U9iHw+Y1p6nIUB7GgK+4fuWt6Iy2TVXlMr4ML0FcgsjeCj56g/Xx0B1edWmNwy6
Nv4bdbgem8ph0kH7LBQWOXDv/EdnNHe/iSk99m9/4R+TG9nnsYT3BUHTPNEHNktwTX+SXxJcuIjX
xjilUcN+y/Gixz2xs4NzY3n+Ou8c4ulMhaMTc/Uhbjsj8mLf1cWCE4KpJV6/jlJwjt2cl7cDl2Ya
Bttt2yuxTeqRhbiBXlKAwyQPGtEC8QMTezrPLLT7FeJ2P1x6RbBllVXIhwEGz1Z72c1OwCtugBtI
kBWLFL6/Oyz/fknw7e02Ii4hxAe5nwJHQ//wBC1JTs1R+62p+vV2RLeisNol4xN7PrlqWNYin2u6
llrhG2rctVlMAy6uDf5kNE7uAowlWOwIJilZrG9MRNWqQmwWBcWqMgmTQ+dAqShMtEPCPaXQvqbL
N4JcAv9OpLk0/NlLpxvh7AQHX8Gh3Zk3SYQtPIBth8GI9+43qdfgt7FgZo/+ENXCPksBvRy6Lx/W
zG1rE2Us1BfOjdDTM41LcTU1y/+la/I4l+LDzNIdjU9Crs0Ao/jLK90BWdkNy6d7cHbFij1zcPQ3
a6U3rU5iqo3orUtdEtHWTSMTvre5AfI9fUMczM1qBDLHioBWLgZ2fPBgWRCi2vev2Qfm9pHU8Tdu
ljOnlMj9UBCCybi0URy2+WFnGG19tymmCF7hpwkw51G+ki5KapU5PzTCdiPrYbMErao5ZnaBlSsV
q+hK6fhCKRtMwxvULJmRWDJeIMuuWt5Xmk5By4mvG+f54QldNaWDUoKbcIB8p9afB64xwNvh2GwN
jI2zWdBerwG0VFSl09jLuNEcles2LcYAHHhxox7KXdhFZoDsydWF2g96MGkHaW5mmu6Gn97gxgIW
O7QB58v9ZorHQx9HJO3ziuqTbjJ48Ox1JnnI/7/OhIN6t64b3Y5m6L3J0gpLysHiqBpMjRmogOgb
Ez+0ounACh6F5zvesPlOO8x58RX1xzpglOIrpBNOaKW4rn81JxTP/Ov1n9NGxfdbzG2sWcBf/Mal
lj5xVmSPv4Er+VVtMlB4p9a4+LY3kmorKPCo+dA2cvG64avvlOCRru5mu5LXp39ANboD797c2/wO
hrAZsdasPOGl8VqPfodo8AjZPIhqLaYsd80eu+uBsN2anWDTpVD4yjzbQ42Kq03prvaT/PQcBIbQ
sM2m10zsRLpwqMlR+DaRPD4ylz18dyxEy/KmPoK3a0Yj14cgeOrzgcdA9M27OeJMiEsHPRZa2UVJ
mtWp0CkJvuxNnEasxMqWyXkKSWmBRI6vsqVPMaOFFz0rj5/aAlOjKcIMh/1/9bXVqBVa/CHlN8w9
OZn2JmjRv/wqNPMVmiGGRhL4ExzqWQZ2/2Js3YHNCZDldDh2Xi4uZmNRy5igQd4j010mcZD2eZQ5
jBIpb6fOPS6pkywiTUTGR8LMifhpiYUJbsr/ZNl2kx1QEh0zqTwHe4v2/KbyEuB2sXYDga/AMEwc
An76a3PwbVsTksFBUo5SIYpkRZZUPgh+f51Zpj9bGJyqVdmQIX/oXQFwE37zbMwJEm46kR/VAMCe
klw9LBhSuYoql+JPPgMET8SK4dWDfDLMUMDWKgGIsWz8BKjA6cTfpbI5B0NOAre2KEZIO2dMB9B0
2BCd/i11rz/eS04uonAQyEm6dJZ8oOZchb0oJv+L9cNcsJvHBhsIrByQlgHM/gQM67vFab4FtyDu
u1aBIgMQmEoE7riXuyqUgEDUcmqc0wRYX/6adXQ9Np7XWVhfuASDl8tECvJtYqdmQ+/raEWTrWSH
ii21uPqxzKnzqXQNfjhzXpIx6eWJuzSztCeTQ9niEjwm/x1sdjVrpvdmVu7OYHr8FcRQ4fKSOid0
IZOfsrMQyZ6lViE138HQ4gIxT5imhCj3c8lE/lUvjUdiB+rfp46R7ACN5zWjDmdRAv3XwmRLT4yY
J26s9PScVODQJWSMQt+8B0aX9/7/YNMFNdt4By8kLxezbEM+wSuR3vHY3zwFSd37RUwujQAYsF1e
XisZGETmxcXgwR6ppqI7l2OafvjRxILACmxitxwNJblb3/98y5ejRV8MPkKcDHnWvMtx+4qXUemU
oS2y3fblDHodNwzc3ftRn/zVjAVgh1k+OS9U62pFatTw8VN6JvyKuWNNc8hjHfIOC5W3PigAjig8
jrWt3bbsVKSUmav2MD2Sg9ILbliHJXCLOkzbrWqI3GCfP5lfIkUAzV1tRXSV+/7u0lJDKKL5WicN
zfkNj7AfmFTBatQ2jgl4bYHOVt9bRkFUm+bCeduyQDmCTAY7TqoytdopWjqKXjwvDMDLuJUT1o6A
awSkAQ+dcTbpAQ2KGQwLffyDVONhf9vr9S8as9KxJEFFG8XgvCxzQ5QgS3BoD3X9gUySaMYysTg3
+/SGGoC7rmXZO8enrpAX2FRIzBP+0SgUT+U/OUf73kM8uxVj6/VKT85CqWxCbu2G0ShtbuWMZ1C9
46HvDQs5XHy2U0dIx7kcv2VBcqwBmCaqFbOwOFgVT9CizdRm6jx/yvhKWZQo/DrNrNz77t36DBwN
QCCAV6Ut5ufn7rsbDBzvPuQppT0EHoIZE8EXkrW+dUK9VzOrQz/eDT2wRumEx8T8Fav52o6U7U5V
J1P1J5oMR3aA3KoYHPuci/rgGOzQVo2rhJHC8XF0NMiXA6uZF1nK/6ZMCAHYErScUG/c2ng9z//n
fkU3mxgVJhVOaaKd6+I9y3EQsFiABbDb+fI/6Y9XlkydW6AyyJD3DtEiOwbEoN+kSLVNGurrh1yf
55Ff4PNau9Of7BcobbCs0VSbrmTzLn/0yz8h3L/qVjw+mamrjGOrm1e33R8u78yFLaPiU2t01Duy
d7CHrN3z9CMCmFl/xbjbrVY4pYiD2U7pVuP27f4eCV3p6sjGovHBMBpKmoODTTM87WcKrKGIAtxK
TKQHycXHEfmlKR/4tGN/I4JUfVJwtn299W+hRpunC9ozaIwNADZ12TxbxtG6EfISPPF80E6xi4xm
p17iOn3W/HRjXnCwdtnqbKtWKXYyUMvygGk0XEKRT1vPgjEtkAgO2FGs1qhx8Dgrnak+jugA3mHc
YTmYOfFc0S/XjIpUzBJoLoU0pj+6UK3svo5kVadPwm55gn2StcQYr/Fa6ugKv13YdJHVZ9qp5g70
a2aHPqpxbFtp8QWnmg+ChsslehtqqCTS24XTFxCXmjxGAJUjE1OonDPRRYqBdvs3CEI2gSbRMLXM
n0U4bovgiiC+tzShDvZtXSNCEhH3BAUt/c4ZAUt+vbBdqzYtnqToS931MAZorJNA/xrswSKbAiKW
2ST5RVY09HdH5EwrtpfGNF8yUGatfSP7T18zBPbgnilXZ0S60icz5h8Pyk7OOTZJwrFUIX4hE4gS
sAN98BNOxEllTHKLTdXIoraRBTgQENLwzNS3WAAAlAX6zEXTHdpCRf+A7pJOmIuDuVa1zYHjsGWB
niG4OSLDucwpKxoT3XAEfhDvqdKqgKzV7iLKMUwsuIijcQyG/e6nuBvCA6ZO2lkcfqQ5ahyQ8rqm
QC1gXs0hYRf8vw9sr3HSNoZ3x6bzpyySm8WZOmfGL+EUBLIP7txhCoczeRyuJwl3YqM/luvuz8++
2iqD1AZUAfS60pJcMVBDrfU9mFWjf8US5WgdOTWq9wXkcK9CmG8wjznimv0q58Ok2smOyRcPF5R0
GNOyvdK9gYZuH8u4Wpm7z2YarKTLxzOTYP/fbUsFFczzWVD8kHfh253pRLKFGU5lTB9RjGOB/Xvw
Pca+xz2lzIJy5pfe+PEe9ksJD7jdkXr+yh6RFeg6ebRXExdLkFTrg6swzFx1afNX6bvG0OjhREsf
Dagrm+KwoIurOiH8F3zzfo8OdBjl5ymr+4UEwSZ2+IHpN2ebvDxA2LFSHZZppZ2c/ITI9o4iJhYR
dVIy4IQXT+B44SYQOSsApFKT25Oj48Lv3uWvsJgN+zcg/JmyQu+PeY4rn359gb0BJ13BHXr6HLF+
jt89E4A0tvRtONes7isywaWIkV4gPYM79EkNzOpWWWFwjn/tkHnVLvnIT/xkDZ3X4IP57aXNxfOa
x7GAug3r/dMopoAIm2+tcjr0qv+niLe2aKk4vBc25wx+OzXVt3caxO+NRf7RBxTJmtF/zb9MdaSR
9MiFzcU5SlOoGwSMfa5+xgqnYyitquHXUzXYvhoYC4igpznw/vJ6IxMxlkJ9RVZR/USBZxK5/qHD
G8URrYZS5IPh/rUxXc7SbMv//4Fqvnqc8oxGGIbmkQ8ZRoe3XhvQfvkOXjd+pE9VRDa9qFY3dPXm
EexrFFLZJUH8Z5YPS9P/V2Wh96dKl+5C316pqcttDj1AvPRu4DRHE/5jMcGLzF+XYFaCfv6aUfBE
xwQ4mis2J0ZwHvjue+R+CJfc7b6rGsi5Mr8CUKNjA9aHONpVRSTy54Qi9A2cZkxZF3cYIzPCvHkb
eag+voVKg2H5egCEMs6jKuwbXEGxAQ3zSB/3kvcU/ghLtIK40YHlzA4KQz7TklFST4R6zDXVsuZX
oYLU6nnxmAOR0ANpqQTLENwLjc4aPzixHgpl1ucAg1q301gZ4jfiYqz9mKLiqDBix03F2jjflU0F
BBnasNGGWBW7Nuk19p7TAFTv1Vuk0iClEsb3j7heBb80jnlrhn8vjv/gt/HgcfvagYOktJcJR9IR
LX09kPzFIyyn1BJcp2PsDlcMUjHi+9+6y2QtwqeXwYnatZJXgOYJjd+xH4pkWeJ7Qos0n2mCUryg
mHztBS+vzny0IfWoxxJMGoevIxoZYA9Hc5UbVYg/m3me+1C7+xxfovM01UK3ZNQh2H4hlQ4vOMsO
b4caL80Soq4E1Us8bOiUvz80VQOkaz4LqST/Js70VorD+jp6ENjBK/FuW8fN71+3DTjiaXf7pZ/F
N9vQrhMt61R0JGvGaTT0UYgFAdgTWZ+uPgI9Tr8FrLxCvfoHo88G/WgKkUmggWsUEVLlBuD7JblD
doKjgH4vv6bFZghLdJsEPbAwWhX5m+fvlKnQyKNpNLM52SfPBnW9dpYDBqXMpAxooFwAyNTDhHKk
/s/cvnIGXldaf/KkAsEgj595wlkgj6kagqa3jjzTupbTe8q4GvWW/780xd/mZZs5tylkVwAfHHTl
3hCJFTZ7fP7WKX8xm/E6ERaXmHjnxDWp/UuZgJVNyZFjXk+jhADJ0wJJbJ5vyFey2BeU+/+ZYOBk
O5yGscRFJiGjyBsZwQovXTYupwxz6Wl5PwtTQ11fGJWgo79zDkKLW6QEmkGJy19puQPIOIGszCX2
UALYBk2uqD1nYfEstTKseS0cDJ6tp3I5pG+73bvE6qfdVSOg8xqcrJcT8gFMzyQZgROWHyKlj8SB
7UgWLBoNKKihwi5eQ3IiM2G7+/vfLwmPV1M8z+SpM525nzR3xEqqV470pYZDG9e5oW8CK2H649/j
yOjI8kS1wgTFVh9l7slJ6ys7N4vkMcasVXrhvhw5r5XdGRVEmMFTiPpRHTqycyANKfyu6/amVljF
gKEQoneIuOrK++ZzapJvOnaFsdxlgFNGRv3NJPNvQLTWSKE0Cr2MfUomjR98tGDGizv/4gav9GCu
EAiOjpj2TP9TAD2G60r6hriRsZiuetwUKQiYZgRtLvhnDjXhXSAr60cUCOJqh2C5gbtBO7Hz+au9
FQdyhItiUVVfrYXfxXL4MIbb5QAzAWyPxaUNXCu5/xLFFDpN/HqxEQSKrkN2cfsWhqsbyUKwbwpy
GYGUkUyqHKbJEKg3RY2PE6ebaJMMF/+Frn5cN3G9mYU2COKx7C3Oduj5Gr7VViywsXz/+7YVtD3y
WzOItkJUAZuAua/k+te1BY083iV8RWtIrpi2IOiIFx3mze4Xed8fAbiiIWmT3ZYjyPne2CppbdE+
yk810L+K95pmQOoKCSKxuk1qpJZQgyFLauBpaT7WOYzOvJ4aFF8Bg6BQCaLbutaB6NTVww0Tm0TK
Jjcp8jFTbykNgWw73xBfIEKe6bzRsDY1pLtFnhMfEPpnqB/qII6DyRCc8rr5JcTnE6bPMMFqanc4
Drh/vTY421fiAxsp3BM7Tb+7jG83xlf9Ts3VSZb62IkYsX3toQ1eRpWSoHnEVEE9UyrzzkD0TXfd
dVGJYlpAXDEvPQIxBfjxcljZi3iQLm3VwU9qj5zicgJs5Ehai0rKOydpM2e1TMUcDe9P0fib0wyY
I6RVd1yL0aDamIbwYDUD7kXXBA42kcC7q+qnTeaQyC606OZ99rI6xUC4ub1cCAhoUFrikpHNod6Z
CC+diIllpiAmwuzkGgBkeLvqa8n9CLEMWFYlogRVwCSp6LD570ks4dD3a8cU5YZUXYhnadnNnPi8
eqi9eJNt5ZCoeTOiyvF8ZxphL07keBtcLL/SPUPLGlh9ig7BGeXN2kxXuRyyPhGLzPK0qLLDeeot
6Nrm8rEXM8sXxBTNyJtK4maEQuJH3Sh2RRuOeqASZRvYs5KVoCN+blb5TL33k3QyA3ZYtrzFx0CM
ToA1QZ6tDsbCAcZ1bwfWQ2qpEc/lhkhTDEqhbSHglGdXGp89tNY0eM7ddPG7WMbfrdtQTFkzrohr
7IEqCHgqV40ccCT6xGUpMXj4DyjwugnQ13ckLdyvWhFyRoGuXlsnOyH0Oca5BlGZH2HQ9cF9s7N+
IEXeHybrh0tUsaxFJmEX9FGJrbVvFucwI4Ad9EDL01F97RScvAtXHIc4kCUmZvicFtvFM09IngN3
Ov/2W8tIS5IOz7aJgcgM2mq1chqkdramUKZav88H5efuwMCiSL6u2J1yVy9wB9n+Wt+Z/OuSi/bM
4zL+VO88rh8W+Ap9fcw8vtSOfl5v/3fqKquruJ9vyxtwxq9lE1jJ5jq2Be338aVix5MHO5LK7X+G
kqo6Ls1nEUE4KeMY7JMmFuTCH61OeqOsphmZsvfhAvl3FWSFf4yCG/IXHt1Roeeby/UZJO6Apv4U
KfrcZFcjIx77HWnQDEHJbWn+aEHNAxzfX/zmjZAwC5yfwhKIghAh8J6IOsWeCa6g1Cbs0ALFtX0n
ivrHR2xFNZr3R7LcmE+0KuL6My+hR3g4pB4YGSONhvp+dEatPbtuOoWKp9yk9tRfXqtDw1iESK3n
s7qQUMSNerxrgFHKV6+zWvBGyk25Vo92NrV4xmV5HZqfYlivwZ7RXe10H8GmvD5bRNl9ifNKj9Ne
E00DgVxpmUP7P1R3nDK2akw9PDkHiWihkva2jx92Km1z5JTdd128Qu3it3IvDpRdmYDrVO9cr+4h
b0pQDZLfzYw0OoiyRpayfOHRF1vookjJ6Y/qTCL0JkMmt2bfSB8Mkcl9g+suw03YMUZ0rGhlFxlD
N1qgi7/o47cKtVwa/MfNtY8LQ2WDSYFjJ+symjdONw+Hvkrunpg0domQTJlCVIr2STM2eDypU4t/
5diKjVM3aWBBPu0GKpXYeB14IFpqNItnwWluplygT/l549Q+oel7eVooqcl/DMye5S14wX7RiJBd
l9eQ13aDa7OLPwXngwuO4J/C2759XKGGAwnemXaJdpCTRaxCNZ0pxVbHYimfr/Nx1+KoLMIhl52e
wr0WyYYqVFEl0ASz0j0H5/BYbs8zpfqxTCvBXl1E67yaivF+yFuJy2gzw0vW24GSvvVDP6Rhz1ef
RVxAJ+eSxCOQYVo0p0jUnghrvSuvtqTTDGNGfI97Dj0ty1jGRQ+DbZpKZsp6pLMNUFLZnBPoXw+J
qdA2GeT3LBjTYsUouUvq5gDZ2AQcq8EpPzNWUojP3IipViTZqrShvxsjngOgGC7j9X2l2CyCEwin
hLEkWPCTadvBY3TJh2yDLc6HQ3dnrYaI1bOMNgW4fLxlsMA3hj0UQC0etRCRHD5YJbY2HxpxqefV
zCQP1Ad1bqIr0kSjGJabO7zSXifywdxmQfHq0SMHmlBlZOB0TTfrIwWgDJ4FZ/udqPPWMeOFiCEt
+0b2OrXmkJF3h4vlioAKJtVCYckK2IOhoUKB6uDQc7R+DVfj40zOxKjYtdQvzqdjLyyYGtY8lltG
yfVK/dcNNSwbfNCrHmVcfKFe60CxVnnPN7uI4GpJhxWZOUUsS+b6iymiIB3lwVzpGHsNnRzQ/RkH
y9jobYXHSQUbO+c5Vj3bbv5ssg8O3VbnqQS3LmQ/hAdSCG8R56fVkxVFfq+zLgASGysbQiqKOjcf
/g2Pd10TclGbKHeQY141amdkmkqJ1OCnAgP0OvEH6qVmWDrzhdbdQbMc/SQd6FOirT5xV6jktbDS
nVUIxDETg/EMdbvWCDm/8wIBoaNAjEhioD7iqeNe7MCEDn3Vd17M4HzKJwW69eeTIF+M1OjqDIi8
jqSmTGH5z/XvVnH7tCjAQ/x+v448Ony4qFibjrmk9yUWXBcw09Kz9mav5/yEGy1oowIdRQiT9r2m
PUmZNgTN1Z7PF+jb9L86wcTALueswiMf9CIgwKJakSdpwaPLrKdCbE8CVicsGidw09cQIgf2BC9R
RMnrRhPJS3o8sA1TrmQnNlUtjiOOXTTNg4qvxnkGJkaTvxMXVmHjtb8sHDlOrExVRy6rzso1XMbP
C7RwdIZKsrDctQTPj3gChU7iiJmEeXztDZbsihaBauOeqblUA+6G0w/VNoaeKlD0KPZnh0+fKo4S
STtfcx1fDfuCZ4/cd7XyY6ddjIW9Ij8AldPG4tAjm+fiC3M9zR406X57zQJqcQ4p0QcNiZkhTghi
LhfAHGdnPHiRzAC0behYnUCULaPS8nv8VFPDKX0Y5qL7avNR7o1JVxytNaWMA2X8Bi3RNZBPmeZ8
4OP6O95jEm1JiWwNhkA0Ro0vTAxl8sBcEujXkutDu6QL6Ovwx7YfP3Dj7O1r4DjkWlvmDBX+inlF
3tfmTPGd+arPwTxBf+fh8M0BDwDYTNOfnpyi8/Jikih/aWqy5wuHuxTyCnKUlQ60GqLcfmu0OZVS
N3O9oyL61HL+1fHipbVUPdCF/PXiYTzKLHbyo33PDhbBCkUhUbPxB2wrwdLiTlSYjKgYnviqXfAP
w7yQwpkEuvJQ0emgS9KzEEGz9pPPIfw/08UiEoB1Fvj6Fs02/y8/x6rh/3hv5z2/WDAKzKdagS1y
Vh3C5M13VaJOfuIF4Wmi43jJhVb/ksl68yng56p69+8ZGP8zCIGK3a7S1OQNlegnIvsxME0QHWc+
p4L/tzrUMqBnTG6uXuKz53dZeAbel1hmrbcHPhyz7KKfSvUrFbTP510s/RPnCoxiC2j89TW9yDWV
QJ/S+f4f0OWtIB0jLkPfxIR/pkUvBfyctLweQQVXmnuGK0Wxcz0SB6s+LAYpu7+AP8ibQdjjQ3es
yJUotu6WOg96jXUVFWYt4YkptMw/0T8ZeqGvtQcLBV2mOGv9E/MbwsRGKA4QPKwgnHmqXLce3chw
d9a39zpeWz1pjnh0njLZhKYRDVXC2epXMAy9NXdHdVdTUYep5ZQFOZJ8g2xLCMSB/5fI8+1jtIZi
+yOX5a1yB4jeT/Fb29g+JyDnbJeVrp+Xo3fNwdJMNceJZkLUM/DU9Bg0Hy/Dajbr3khMnjLzD70r
izZ0cpWC5WJgngY8D6s+CjNB3HBOkYyIO5w6+THcCHMoCbkBQmvwOOOX2GkPCs9/ThTU1S9hH2bW
CyhZcQY2+DfrEVSZ3noxT8311+idyutNQtN0s3nOulrRDWGg7OX3Xxw1h8/7xJMqn/H0ityw57NP
dclAwNHSN6RvJcvRgIDf76vMDn5k+de9O6U49L6O/sgYUvAiIWAXqhVQ/Ij1ZpHyW421QHaWpHen
oLbRYKP/43Pc7G9I3tq9+de0dUehqReV06Km4u7h1InwZF0MywHACbFC+naX6s5x2WHjgn3CAUuV
GP2RvUTu2HAbIy7le/Omo06Ee85mTrVRl9kT7xaZogGbboiE9UYGAKVIbpJw2mVEArMP59qjnJD9
lonNEoUEuV944NmGO0PyAqlFYDPj7Lx9w9FAklfJYgZHyBpKV7v9811fGOTgyuxso67l0ySMUylX
3aLUjGbxAiNn4cSLp4dQ18allDS/DlP4hsS/7cb2IGW8AvDgja5ZQo1bfYUcuk66snblQHqFoYgg
mDZBfQ7L0vLoqCWDdp2qkHSUVZgmd2E3ttOfVbV1QQCVgDQlJ18+vLRGTrjJWOwLCwPyFNYCZAQY
DEgo+EHEjSFY5YhV+dgBQWUOf3bwL0VXU8zILowPt2fy6CXCne/oECM+1vIrr3FTrG9RV1sehibW
maVgkOpqu3R0b/G92EvHqO+K7Os085xu9dcNZcCv4ghF+mgoWRmZFhhivDRRtKNctB2d6htVpJDL
tccx/eJDj7aHZkzToP3QRknEgXrs+SCTLm8Ryci9CE3LVWMKaxDHwSRP61c0HO+kxqXXTuQpgTcT
a6WCiBajrNyeT0ejXnapzEdDIvUYfQkLoIu+EK2xL51D4qBwwd74nsymR0rdLepUJTqzNzEdMLJU
80hICR/F49qbfyd3S6VdjGfamUXeYtXiqzlyia47BZoK3x2fdeBmLZoR6y0Dc94PKrfFnDXHADyu
iFQ3ECdnxC5YzJ0Xki4/KcbWmlaqTZhsxl3cu2TtITGXiENdwacH82274GBDIdVKE0jocLUPTYDP
GuLrRu0pAmiMClxyjz7fQ0Y+rpq8VjMj4o6gFBR0SHflJVLaWke8Ppb9kDw9Ioj4pYQRV7q9bX/j
CmE3XvtS1ZAOeJD1JOmYgw0cPxEorTPZEDTVQ2XSt6klW4/Uh9/Xb+i0AatH3RckeThhUXhSYabq
kDvmS8ZWhHbQGIWxcBfv4yfyHwg9q/TS0ijWrhKvhO1YkUFLggDOE2VzcbSZIG4i0ho1IC5S0IKg
kEUvZP1aRR5gaq/lp/DPR3+7gk7pJ7KLhyrh/s54CfUaoLlXkiSQx23WOXVVop+FpD/9x5NxhdLG
onTAcwhYBGuzuGDEaPnDQxFZMe+5K2R7EDpa45gGb4HFraIazN0rmnaTaQQACuMeSbWV9AOHy8sp
mMSEeawzNTHssBZuPmbrgRa3yGHuAWKfMURyXxPtbJfOt8m9aeeiVviqk4Lv2lYtWAzGJA3NNTg+
Nw0/ySsfE5wz4bCgTrgswp4uFu26fQK1TvliaIgLYQjqsjNVcZlWoSagyKH1QsaX9lZ2kWuXdjDQ
EgTCBwamENmc1/TgwjM48EVoulh6nM8hM5jKU4bXmfPMJtBFEcg5Sreg29asO5syTu5Hy5VkiRH+
eStnzDU0NKgtqo0ksf4LNSEvjMeDAbFN/dl4PLjsqrrTfzfhtx0qRGbo/Rxkz4yINC28P0LLDszi
jalJ2TQgvjZRRqPXhJZuqMS1uhxTx5nJcZKTOUq7c9D1wq2gJYm8UkWjpf7Z/ZRgqAIIWDvbN2bY
pUtcBB7fLhjCW9SrmO1fRa2Jkpo4JerciTouaqQ/XrZA6yz3bq1X+fhW3YnvCQ8964un11R3DZ6d
s2TRhBL2aLul/a+dk3+je47ZjctVWFxDtN+bkCg0lWePKgRO/E4ylVn/ZCRoSWdpe0zVWm6aDoLx
4yiL0AdZu/27qPSps7WLpUNH3rwPjkobGaQrP3+I6JSHxg9PV8wStGVK4qyQPkpIT5TXKTboCjvU
AinsIWWIfbs1SsKzocz3xfum/zpWNQ47/pP+5f3ZQutorHsZwNiIfBaAVGHIBV/QX1VPaZKs/Kme
ciYEROlaZRRrpyM9pR/f95U6xActd9jEMetu6r8cpluQNFG0jQK8VpScUjFMeGIRdAWW4+PF3FBX
TJ+gKNoaQa+GlH1UQWDrMKrKGgQKWzCullwu7hyAZgsu6b0hUPVMvFJ8gi7Tu+oHVY0fB5luW8j1
hi2zgQt/fti9Dp3+4wRjx30SdYM7Zgv92ooKmOc5VfgK9SctAQXax7IFHEiRq6lHPa+S5bnowLU6
fVLJBq2a+Mw4AXcPY6i+FQGgXh+2N+HINgoYMBWscZfhr7P1E9p1MNQdnvAILQwetdMQaCGL1IaW
Hb+n8y3oE+adhRgXqfxZ9mznHAXraf6e4WLVeIA+3t+yrMf36n8+rrDSZ8ZvXyAaSBCiaMW1rQS0
pqd0XxU1BWoMv1R/Yud2Km/+xm2zIlI5+DRxChS15VsswSoZMCs8Rc6RjK3d/BfZDGd7sIf0T0BT
UwykCCPCfYrND3Kj0ttLPjI2vAICYVPz7VaqtiuF+djtUpzlbQUtmxI30AdWeC57AWFn1+lGuo1Y
chLsfW4vF1fRf0W0ry6XujSc4m+SgQmq+N/NkTIbWeckrNWH/FcOfOkfVar5ZnZgxZxV+5vufqjC
7+EowD0oIxFJH+vx5zupBYUyyfGJl3RwXHhaxBmv+7tBlABugPZfhJeZ+9DrLRm/IG9wH1ggopEo
rEryZpCPdAKITlz/yTQmnaToYg6kTl6P8sKRvoeJH8XcA93ISeqnEQd5h20ChLEWfwWiuw4HnA8M
6z7RWQ7+eDrBLJ3HvWXJMuactF9MEWP1xWrciGQeJmoHPR6hJiO4p79oKI474SxalQ369CKNKssB
FEmya3Fo/gpeY0B872tEpFQ3c75Ec104Ho0zv9Nm4muDdPytgKlcN0UCoATPYacRO+/HKq+MHSmQ
9Krsmq0X6mzThZemiLW3slRAK5xUkLxkleBwbDNWvZ9RDgIkyLmXRl914so5zEs2C+5Zjpv90jMC
IytVYsobx9zictTjibPb9ZTsxuc/ZDnni8jkvcC9YpnpIMLEgVAVR1cmjtxuBTyKq94+ymp1oVip
IFrtZTyZ+aafA4ubmEEht6n7v2685FXnsVZ7hc1WvCCqC45MhutDaVDW9gOQ8qmJp0Stbt3gx48E
4Y+jZEFb43Nmo+ec26TZDEEY5nRZGJsCFpGci+pvnEdjzbE3repr4wNNv7evRHKsgned81Jhn6wa
F8tqefiN79VjdpVWDZu3LTOSOnFTxKVeebHsoYfh4cr3GOaSURCoMNWpnCbA+LcwGdPkbduYj9Ue
XHvNuM5c0vtTAeLDB5n0xoYxdOspZMwgDQH6hOJ5VuC1LXYd21cNFYYH1rJKUrz4oeuamRtw9zz2
Mdx+xmTei3Nrn9xl0lEQseAMtGbK7/2wOJEL8ETz40lbDFRYohs5yIjpTP+vAbwAsuGX+7dkut8K
Cgg3kMwRWItSLU2+7jWKHKhmRfteyRYy26GYPj5M79SK8/+bXw1AloKBVRUNw3KPA3TgETbVxCYh
BfPIGbeC788ZICch2pcVVz/dmUxUOkKu1NYiDLcM5kGrAJAe2mmwAUriESjLvqCePT03BzYkTGyP
MnIKz+ZCPBDXDCciSg1QodPlsLo52kIP4nNwvwTVDEOUcV41tPfdYe+2Byx/fctmdSaPQ3cSAf0g
JQ8mEHzy6R6629XmwG0W6nRx5fGtX8sXFSYz5pQTMt9G6EcgruReKmIhiEBaqhS0/JVUjVCBrv/r
RdVCorcUK+iaoFEHfQQtmtIonHb1am163XiizMkFqM9WPdUV1/IJU+CqjESnrBlUqup6L6AVAFN+
UJ7hl/Eo70OrRkJwMJ75zBqDI2f7Kh7KPTmv8FtDwHIK9zcLboWA/L6JExfZnpCORAHCzcRdVj2Z
IktdkqlKe8Dq99XAophhYOmhn1aoVE6E3YkDA83cgt8ZOUVP+zX7NuzYsQaPtk7tjtZU8faqkQ5P
5vbDpPg2K6T9h2J2aY0OTfL3tlRMA5+PA02kg0GlDlj2eWp+L0Is+L1BJ0b2N4GLkMvgXoQNhEWx
cDqnArZA6UVx//8YL16CNpS3SNpEAtKX62P34lBdsSRs/2XyYQhYDxsGYNBIer7Hg+6qe0Yk0OXG
iQuw2JOIo47jUEsoJeAsrdWZ109pt2jYKr3MSH0RUDM2PQzfxBSxOy4B7KMGxeGv3xWS7sj6k8Nv
c+gxdsWD+DyAerv61rrfzjAMgGvlEN1jGDSWoKo8ZtcHYwtvmfZeJickudnth4DME58QVwOXsgmg
KdYMS8pffjtTQ8r8wj8FQsJ0mzRDp6KSw9NdZTa9gIQUmBG/RBJBpLiVNKrQHmgUXW1N/6jtNNqK
uybhuJKqIuQysDv8tcQSlP4ll3r9WV/DRZynySzMdO8k4itExm54QNhHU+lRGqulxJP3GYN9mr2T
utIi6qa5FMIZoAjvnlSxRk3PhOqsPj4fx7DBluqz/KJI7TjfUPH9+st4Sh4gQYa+LferuxiQ4c9N
r4QF5cL9sNW2IS9hz5GJ0W0feyxRkVrHf+WsNXJ1eIjHwVOQCJwKH3riNC2zSAPgO5oENS3QVLsz
fsCmbpJuGh2VLEKnIRTV+k4HVf7qpJ2dszWjNmZUMJq0bIqjHDaKBUK/OCJI5YhL0WhRjYW3CwSm
Mh8BIGu0D2xtNXAIsnCZOEtmmkqQHBX02cHrDpqRXbJbVJPnaPndJlGx2uZnYRAN/nlChSppvsER
aw5jkQzXnkKz1IEDshhT1Oo6rHKfQG7OOB4dXd2cUNb3E7x/iiBSuxjesztIvRmtC6bocusaDAGz
/aQMGCrXz0kjPIIEPpYNeWJxSRqxoFQjBv4szMCWGHNFVLLrMpUwzbf39gZ6UdUTBd5H5kqoslHt
s0KX3d4xnfoC1facTe/iPSvSiKT+iwRYg2wfA1gIFH74DfZlzjNwPXGVm4gLehOQkwCd+H6ZYKL7
MNYcOPw4JdYrfkttqdj9rTa/8Na16wJ7cUNrXxwaZw5tDhNfSB/87sijxUjyrzAZGWh0WsuN081K
KgpOetwxxrHVrj5SjOHIsyvuxYJ1AHdCPfAXr0ol6n3EcOJqDYy1er7T/kkLaYe4uv0zGsaFLni3
tUwJnO7XrUnzCODhMhl9ANg4kwa6cKRhfcvreScYmTFarKh7ggJzg5IO5kVCCUOODIIFQRuedAbx
mtE5/8OFR0NWaMYtzBZSCDOX1m92h2zjq42c2oLda9DYmThctsg/GqR0gBxalgWQOhw1ELPEOf/J
gzbdgSFdsFpPzrYEcpQQyta/hi+wrYmfzLrpm5HinyaZdBhLGoBtJyRhLGJbBqI1EMbWP6OeVVuF
KyvLabFqgLOwgsfRN7mG87jOYvmhKkV/j+vzP8mLrKMJ4+CZ7/uCp/+MhtdZSo+e9T8OIYXCQ8sK
MvUp1O099SixHaDzlLkwGHMyHzEJwtxQubCZOpoFwK+xq7EM5Nume+KU8pJ+jLLNqC6e4ZXhGjG4
lpwZ3TmpM/Juln++ShHyFxcDBWBTqUVJBDjffvODKHJJOpAz1iTSsVYhuJnJ6Gj50oFSC1U8B63p
tDp5yiPxYrkPvS4LRgZ/+7dsIx1cyQj51F+R3cnMATWHrOPEdj283vWtqTK0o7wmXUCWdd235k2+
0QZUMA0QRfvYvlHmkKq4IUjdmYVQxg97spmz9nbHEcyHimPa/nvfJ3J+3MUlS9b9uW4RnvIYQj/2
3reo1iZ5Ty2/5pQZTNjdcdFz3ial+15y60s6WDpqRlMLpQ6m4cfQlvsBhCGhztiu8dq6gnNjDiQT
FzC54xh62JGuUPXajdf8ArFlUX00tsUJ8qi2M4UgIVlVs3lSmWf370oG2DQ4NHBa2w0pPZdycCrT
Ic4gUlBHiQuOt9vRz/X+dgckQSCfOy8L8NqN494J2YNZoMM6+h0+uoRkb0bC0Mp/Q141rd56geKk
jhz2FzlfvDNax23YUPntHdVEWp6/pPDVcr+ecmp67PR9Wyz1ijjwJrSwYG8hwon06aBcbqWePZFW
fwtWdLRGFkdbhj0TnTm7rZ4hwO8RAu//3jYC3tJJR5JTs3J5ytkwSLCqu7zP6odDz4Cr9vSL4PAj
bLNAi/cnv7e+MmSk8fRKZq8RDU/T2MG10p8aL9Qb0ZvXMsLk76I0KuJsy4jslwz16jgtUsXi8mL3
qsWOgB/ocpcN1vMDD1p+kC4jiDp7D2eLKG/EOVkY+s8U886F0Si3ebozXuqg05xOCPDzoFxUUp+g
Ab0TGBfui+fPGbkaiJVRMUjV7PyRjwelCK55EdxC/x0stLk21jV68IiWKxgMVDQfjNmszKDMgfFK
aytQRsOOXLOBMq56L3SwZRdIdPQAMSAUcxCR9YJQHPxVvvOTBwbUmp+jFSp+LKJjJsC+OYWuKSDg
PSIXW2NkTnxLFhM+yHLwLlsmM7X6/Gon2hdiqFIgyIpOIfTHiw75HUaOZluJ4kpJjwMVb3vCUG/I
Sl2pNvvlvJAAqBngtG35eqHQAD0eosmAzKuNK9w9DkKsnM39YUC+US4omSuma4TRlWwtEVnFg9uG
ZtgePuXgXVmZ8QJSKEXbU885gFH+xgJkeajZcJRWBlw3z+jPX9B/cM4zhInzEdgAHNUEcPJc4+DZ
snlAPZc9/6kn5Ljj9n58yrkjs5Ts9QeqfaM3uJXfztI0iHeHSxDY1iQP3Sp5eBFRPpVUySsNKSMF
vgJf/ApDRNB2efOUtiNbrUoMuTSXh+2UuAK1KEJOsirOwwbLRMtwYQDG1HKUFMR91TBfLGrTcegE
ZBeBnyfeR5TbG9azTQX+9VuCeLIgGIJp/UsV5wKc1Svh7X80bIypPDtZdZ7vlrAPfFmPX3f9pOBM
neyjZ21BEWZHjAUKuLJ4/7P0emaIpOXw4aZHvmjui4TsakSkMFZKjpcuJyj5tGliVu6EQ24QhZzs
sN3aDFeczPZz0Cmu2tyePru17dk7lNcV5fFwn0YsyXnqhx3CsM5GyDCwLYv9nQINpAf4ntCgTjGy
8yoEacua1x6BeIhHydXkERiG/yI9uGcZZgmApcpbi6cAeoED7OSyv5r7FFNz8iPFaGPvRrrhH8iH
CYAOZHNoudNBTJKKlCX2e5bASQZxw+wbPo2+vzzG+F1MKSaPiDwMNIgh6KJOtO3I9QzWS0rW1TjK
WuRz1nAkpcx69ZPajxfWpEBEQmoBAXFBTAFKhyMuR+VM2o8lBNQaFXawyFWUFnj5Sv7v13UsihfP
kMxCod1W884t1lSswI0ZdktrI0We6S+8AZpQ85L3nKL26Bp7LwD+HWYzo23AZgt2msw2D7pzq64a
pzAfKSDnqDyLwiTyMfpU/GUV2mnXIqkOa8lXy35fbBMitd4b/qZHmPvGgEY3iAKVksV6H5dLWDON
DJMZCJyhNBXzaVpxh8iYznbSQwF0aIVFfwgMuuTRNhOAHQfxwkCagleASFjrNR69hiyG6GADLzcd
Fy6cPTwfPS+yu5f/ZBxyJTecOlsMul4FqPoEudiFiBLvw9IFkX9tum7Ffdj/9Z3tIcFaLeNfHe29
BG/BMzuD+iESF9tkhoI1vw3UjuEYlnMmh8DAdM7MBbBy3BqAtI3XdQpQeMYcsdW7oS2ED1FqWIuS
iRhikV8IEwgrfnWlewY1CCFhd2JwzclD9gfTDf9QXgSHXjTEqSDHd0IBUpslwa2gCyFlUkJumbHW
ESj/bIMyPKiC3rGSQexw7ntCpXJQrXbOQX45i3XGrhQdsAlUa8hG9A+1kko0Mv264f5f70Kciq6i
A1aRh53KSQ/BSv+WOasWas6+k6TCsrtjRjBqD6CPORKKMtC7zEfdKu+2abc8rPCZJ7y3sUb7uoBi
RJkb0y0CRZu67DIPRcMXnEog3ZjQ0eeDiHt7vwPVC+56yOSc7Ut0FeMkREvyjlNNvfGOfHuWUUYc
mXDKrEH0G4Eo6LrH6eYLWpyZmX1xT9PexwH1Z4xz0Q5XezzybdYjyyVBjeZCKqyGwz+gFovLMORj
IBpQcVOlvgaehbpVZEzpTddRjXhV6HwpC+wotzd3lgofbuNfkHjDULYlcJ/hBQEGzNFYy2OfWVSo
2MD+rWaeH6vyYtqSO6/mWsVC/+w6fn8RY8/FT0j7RAeGUt6OIXKs619YEr0bhXHQyPyz205GLL5u
tSn6NcPR9QE4Sd2iBuv3uugSmJm6KOALRBC9sMOlN5cYg80ScCUFQkz7WU/l32gZvIDyONzb1qpa
9H69NEHYrGwsOP44zMh9Z+AaYCJVhP8uYS42FaQv0+w3VY3KOxcb2nYWztUX8HweGTTEM9CaCF+3
wkiqg5KP7mttsKni55/77I40XCCm49AQumofFqgVCqoXXz9U2qtT+FMZCsKRd6JZ5KEGJnbc4Qnh
ufL/OSqoZwNcr9WMe4fcUgKaKKWi3K2baGO2Q+ogBQQiETbAMT4CBoyqUnL3uNyvCoSVD9d6dvOI
dstAPpd9vSQyL0BwqCDVnwHSC3QV3Htz4EXwJFMztykUY3rmb0w6b/6XbRVq+66gGscfZmp7FSp/
aVohbXmEJfDtCLdE7cLY81jOYYq6RXGqhvQyTpD0x+vGiq8/6QZ1oiBhBDT1Hf4sFfsoNanpvIe4
xchZ+MLe5XBxGlhIdVStkRWMLwukowsGlmDSAYEJQKH1AO67KIh0rEO+IdIdU9Kygm/rAAsNjEkr
CJZCR2crE/A8tvhoO7wN1zTm6OI4ygZ+U8NbySVYXKSUnrMEez0F8SMXbFtIP3O2BBJzg4TKqeft
HOEU888NDsT89qqSWh2unlbga3gKm32FEX4Udw7OFWVj2KBoF/S9R74rMpmAKU/bnHZilvvaPK9Z
MvrLyQuoO8IapQ/x3WD8NpfPr7B7hxmRl7/GJjWK1ZiRJI4UWh04YhgOtEHS/GHz6gnG1lQDNqrw
E5ELFaRpsRz8t+6DDbrEJpdnLA91ILrIFfy/eAUJ1JV3YleCzAKCzVoe+7uSLGL1gR+54UT+Gleq
uAx3JpDVZKkXR6EkkYzAr4iOziteDRC6YcrN4nQ8xXSmEhuuIJfFJmnh+2IKQMRrkLBs8RxmhicO
+74tKVrOPKqa/GywDiy399L7gSfXHffTOlXexAyMPmXPS7Htkf/ZGDYR1mJ5wKYk5dN+AnL/R55d
lx0NTrXsWSyuUMQ7LNdhkCNlZew6loNe+8FKQ91bKOsCXwKhEqjCsvA3kB5oIid/jvC7OFHZGSTC
SQhh2ZnougCqF9Cpbs2tPHpboKTqo1FbNiFxnUYRx6lTMPbYCcatAb6t0q03h5C8wzkC+F2z23zq
Szi+ClnSRJ+64qBVMCZYiWP401ep1pTS2+5IszhV7XFt6YdVR9ZRnKl3yrdu2azQY+I+m/R4UsEm
F8pR+fYBXmDZbwqtTA19k8H1FiOLnb6LfaKk2HdnjKc4+zAjEkewVGnaFJGC1SM/t/TrzEVapu/U
oSFBNPtSxSnZu3sV5K4G1bnnkSN9L5+1sqZ1YWaWthu2kBLldMW8UG08ijls1p7aszVOsFgpUJ5w
7HibPCMgUxHyD/w4IppV9cBreIVMn6RJ6tFgawOs0sL7vl0herjeKUJS9LOWgKnfWuUYr0M+fLVz
+NDFiPjeRxyuyUV/iUdwu6IO/Ro456tydQMeI5Dyt1xc0cqItAqIdIhOwtiIvYmZMnPrUuu3Yj+f
Oejc0DHHZhiidYZd9cS17upEkmxVqjX8fkJ5OnHpw4Nzs2m7dyW9KnPSpurpiJFhMDFQ31Nz95iM
slG5RCZDqQmuQfW1tQkkAdvBpjpDdPsqz5nTQQnygu2xJ+brsP735JfLpL7gAJn/aQN6pUOWymKC
EsMvJsBdKDSLqblRRnpGhXENeyzMh3C9/P4gYsRVt2OmbHmFH4CWUnA9m6aZt3SgGATtsgG6D5+V
cZRG24HIhOv8MTFmU2knZh6QN9bGlC0ldoCRtXah0j1A5kThxSykcytegEgltuEtn+kYoQk9Kztm
7WXeBMlKAZQp8C5Wc+xEdjaDG2OcBu3UfRmZqsrlL8K5H5iGyw4vF3etqXRJHLMpctOsAb/qYAhK
dYmN0IqssBDnd71EvdPqUT0r5Q0l12RK3lHbczrL7ecAnbcA57MvH/auoLGSY5FzAG9bbVpdKsL2
9z/mDd7E2hi/RhLE8ybIeoMK7cjbUXOqpGgOy8CBTl8YJiqVO+yQBUlpPRWX9l661K/TGDBvtscr
fx4gud4WelrQ8Cv57iOkvCwApifpnngAqM6iSq8ChejMQiW8V8inhGNNJ3rKpHvp+2RI5s/lzJpt
yueX2xP0RMt2KaYzR8klTqNxsrCw17VZxd+iSnpsqu/Lpyu6SBLlBbfzi/xx8J7mQICD6KIM16NV
GyaaT9DcuQMDyNhrHNYjcUT+HgOuUnqHbMzo0y2XdPOYrVHkL7Ui79GxdJ93wx8Zr2f5ZUvnX6F9
XFwWFvFnwMPgWGkTiRz+jwh0r6gVsZLHPE4udP0eR0wZq+yWLPo9kU17V3Qi1ScUskSDHk5RqmA9
fX0g2YERyjxKkRgUu7kzDL5cyibWvz1TE/RMfS19U2/JOKnqu7Xa5I3N28m+3Uvhj6zIQ6K34RIm
bRnXiv3maGY4EQ04uYfB6m5QdkRB5IVbfo9US/iB7ekcN4bHW6TbQW2IPVoB1xpgt5JLVLVDU1K5
w8huynI6CdcoDKQbCaFc6z0vkyjeIoBJFXN786A5/bmSGOn3p8gNjPlqC5r5L4l8P7fr/DJRylFG
kpa+o/6Aqqmd8iFkg3GEn+ZzOttCX1luhISCqN5g3mOG8VFnPMmYV3KPjQtbc8l+KtdKT/b08PJS
lCZVczeN7i0XA5BuwMfR+193M7hfn+EIilQDDb9nsqyN2A///Lmt5KEyQar5YU1pMQ4VEqFZ5XaN
W2O3SmsW6StTgAn+NymX6yt/oEFI/YX0tSQJiOjnr3M2FT7XEi1QEB5XDMk2SE08VrD1084vo4Rk
xlz0RdM7TAu+ANysZxCT8+GyBMeZf6O+C9RIGmwpU8W0wHwNbgZmy2Qrg6nv5HrhrFTC/xhNrZXs
ecQ9fsYfbOcuIhkjmn6aBBZ+9vGEYP0r7t/GEEXBlUBk9hYLCWFVze4ifLbVvZqCpJNPiWzIEcA/
jmuR8EOWrkHN7DNrlWGQ62tSvrPcJPpL+PBkEkrf2YqZdgzNBioSIg+YayZVtUF8/VMcgmkqSw3s
Zj0x9shv0/JMyyQGey667wB82HKFB73WMkR+wDQdKXW9whRaalp1CBXFHjghcVISs02IerC0WsVF
UUf2pAqii4km967fv4IIeQ/iReCE9g/0Lls/nUlo55oKxECD2yDFCvn7APedIef3zqIQBRkOlLLb
VnhbdA+7opEZPheh8Rpou2OaiOkXd35c0h7GDrxBXaQuyYV/9PayQyRFm40s0+QjYGjKGNHamKqR
9An93NDMEHEYHhXKjtDgIRXNYzyM8Zrish2Y8PioauJ1CK9KhMc29td60IGK4RmIQaKg9/prwGTj
OcrvrN70N4RRB8n9tYoAo0mitlZ6CmGKsj+YlVrdYrjfx0L9266o4lSD3SCxp8FMicsc3eRqgbD5
Lb7Sjdq9g4gRs6kXzCIqtKfI2VurRVGvguIC1QoZb2io4huZmAd3WPVkX1w02UVLL7+1vFCIglVn
720regsPH9RLrjMTiXGu2WhyU0kxrtlKiKaGTDELrBs/ZVKg0qK7ghd560SblGHUQbC/OBG89vne
/Bw6qqhyMWoSs3d0tK8kVC3RGMJxPlZuK6sc1nYE5Tji/bdl86Rqo7WDu7rO6j5W1++L3oPp75ts
lVtcPI3Gj0faJywsaSrv/wA3Kw4q2iKruy6TzRVE+H8DHZmEtWCZnmJRqGEz5gMByUKI697R+KTn
MlOTCI6ZKMn9CpvNEKoFtdCz2YfZkV/OINTNGzPjzKgml0QFtIVOLrDOvWSxRlfeURYRjZzWa8rN
y16XDrdD5RiqSrp7Lyq+klomzvT8ap1OJDrdFqss8lZ1zJev7qjBSoK75iRC6fEqxH4G6iaf9jX7
M/ZjTej7D+uRXqCm341Sv41I0K7+HZDTs+w0YLksIvTpwoeUgC23zgr7MJp1VKt68fZhA43h8Ujv
fo7ski3DFGmaypKDFU6ACoiZq+IvWWEIH3gJdRM8VWzP0Dx4ymWLaqARw/JWNq42e3UCY8Np8Lju
0fCxQj8MVmlExNQGqkdVv1Xm2bbOn2tqkNxfXiqj63vG2b3pFWTFuM/3Sm5jKIgBXYJv1FX7Vjpi
2Ah3P4E6VuBdQBuWHR7u3kzXqHvJoWk364pvPVS5hL/CvJ6lURoPGuNJpSfgNtafxXDUukBliTGk
wHCkftrYVNzcacvaQA2j2dm/YRqnwr7c1kzRyASEx7o1HU8nUWslb7wAmifVjtynCGwWK1otzLTu
usC6LlTbSQ+zJdnnPqphXid7/euwNng8f1GSL23jyJhtNRkgbeNg610UXKr7Bzqdjy5hAJTwurHL
u3Y4DhXQ3dLziLn1yZMfu59H74l9am/3zei7S/Jl1Uk2D3JcThg6170ZasMNSsO4/My9OgBENm3z
mftE1bWQEBlO7yE3IYCOEtZxcUMny/LTU4RvCaAwkAvqQOBQge6uUYOoSAWqyLWxJBlXd8QlXZXY
W3r0kz372Lx0X3gUfbNxJ1ZVlj/58gIQzx/ykPqdapo7nwlTktA2rdp/pMNbVh2IskwG4Frmgj45
v0MlAzDix/2z3P/RWbDHrbZy3nP/O2ocQ2XtvgGlAi0y/kyNZA0/LCeIk0bEVTL6ZS7nY6znWbVq
+qjZSUxDfujlAtqHHZm0QCnPHKcTBnFrWIGkWt9SXUX4m6cSIDbKtyJLDicMBJRyUByfCyMN1+4q
SurF+Xk3VnKB4tgQYvh84kb5+5lX7yTtaAgJ5PFMRyi/pdgvVUZKjtYpOSTtl/pM0+gQYa0b6/MV
hnSH9R4Zgvou8KL32nY6tp8EJy4/F4aRUp7vKHXyomwksodhm8uI2ilrbM5yOUkmSaY4qoNtV0mb
gNNefRwyf1tgknv8BtfIL9AzMtg3bbcVAgaPI/sbavzn0zpNM0tAIJbzVEVxhuPiQDqCEEcKcVxg
08e0dnqgTEze9Yq/SLbdLEj/RQz3eD93Mrng69TxAjIqeFuEFCcUL0eFsxtGdfF1dWW0x6GBFaJp
QyXxPq6+V2wddvQjugHDb0uCdOOoFCozt4C6gibjD6meH0Tqs+BnF6DvNQr0v5E79/i9mL9ixJKO
wK1dQEpAdU2vO/6ncKE0Nw0YnNLQCc9fjqOojymI/iaYvjkB0bEcAtJjcrwgz0eeXs7C7t+s+gg+
1zpgY5xVZwyADSLAwZHazGcYGMFBg422GQCTiCt7IORdBsS2RHeiGiSg7L+rk5iPm7Fz6fHWX69g
fvh4T0NwUaq9ERhVuAIc6s3jmvEFV0ThCwhIzvkwkVYHJD7Ld81gke3XVxrgKIJ6LdM9y1JUalvj
gxxqDlf6M9qGPYEZ4xfaLz2/HDzDh57LbOp+u6rSbHxehfCXyYOsOlpfycs7oAb6wPsdyOUzszDP
ortEQYKvtUNvqh51CLVeEXZGeTIaV0+Woo0YEEMkVNzIrTZnlensygFWJ8jsriBSLMH3s2EacNKO
UzbYScz6Q6Zwzpjg+RJuroM59Mpth011xRxyGEwBOLWZpHSzRm0Ovna7vrI7jef0FPVjpwMXiOf7
OWLg59lqvC73XZHbTtBZfrzY2942BUWuQckysFGdzjYZgUq33teIXbUwDNAhyt4OywTCQ68leCsi
fyuY5YbVqJkiD2yjCWPt32DF6h15zucdLkMFecmpK/r74dBva2QVsYuu/yQUBddvKnVk+VfxPCYv
ogxLtl/DpqWH9fG/YcXmk3Z2/7QdnfzSQbIYxk3epqZ1fF2OleQpV1Y7PZlvWWcqly1Bx8RAvDTH
TCEz0IDMrJ8wtwszEqtlDqPsF/3NWNrkOfxJv0CypJ29QV9zWV+DH9MTiwM8UdcjozM/N/vTLJ6d
wlgp7fr7+ntIf6gePZWKNyi4ydfzGhq4ShEboQiTJ55i7WcyCVfhlvmYpcr0CA2LbdY6q1kGXeSt
PZPoEcn3E3k3QmQH0bHfN4ePbi1X2w1EeIa7Pe32W73pyIEEhyw6wgtYTRvQfmYm7Zpycm8MeL/l
IYe3SsAy5kU6JUm8kYQaxKVzolGKKvVXXzch6C0/PD0n9NwSfJd+cRBPHKKvLeSpcmLcmap3RbyN
VqBK92pKkC6YeZoi/nvbJFDKHJppar++INb8s/l72cf1ibITWJCnS7wzgoxdqVCZH5IhAow5C+o5
HsVBKXCEuxiOtuuKv7TFgXWqxNA3XsdKWpmrO897e8IdgyuG9JBpJlhjPOrksDDfbV9Mz7ZAOub1
fgqdByKBt0/5J9SzO/GVjF6LE0XgSKr1wYolSoid6FFMszWfM360b7xk/wij5x44un/iSGYx+aW7
ZsRZmyW6N7oIEHjnSkZHiqArG//2hCvWef62LxBkj5EVZ8ZuhaMZ3rwR6RsyJ97zA2qDZyEmub+X
2656EOU8Np6zo3qe8IhZu0rz7UWw7JOXdJrnPGl1e6jlPda9adsTB88juq7/dHEv2uodIhRJBK3T
Ryf7Rjxy9aOOqipLclKdy+MtuW18Z+djIWMo9qx0GXIUpnEHVxubgODlvGEJzC1Vxmx9J4QC5xGc
EKp8AXMaNLX2NWJ1SOaHM6wH4mzsyFK5xygvYWyoPiYhYtNLuf6CEYpjSlKmW8j3qvlyWYU2Ofg1
irgo6qZuASOVpYCakwRujHzAYAtMImR1080ltuBvmaNuVJ5wsRE+8hBHgQ5VN4AdzMsyouqf8kRK
Td3U8jgCWTccT4ANiAsWg5qyCc48bSdh2leWwO+bnPo4l55KBFEVZ8JqNKjkN3ql+yTlO+tSzWLl
mHTGdWJX4q/nJjN9/aaJVPTjd3I7lbvA1PCkz33oJWJp9N11bjNxYvnxyFlEwBcI6BuZ8vNEI6jE
LeSxAeng96XHwY0CS5AuPEnPMg1FJQkHqHuoe7ceMkOn3RngOIV1pKD/CBuZnkubUiBQ7rB3eHW0
BMfbm6D0AdWQcws7MR5cox71BI/e+saML86o+ArO8Wvp81SwbkMWAp74rIzRdDbxpuNmX89CSkL8
lye6w4U8MAwYVkMXxVe3sfXlfgwMzajJ/ArvJcUl/OlxpCMCcKY3paeVVInxhUhUd9BPiU2p/PQ7
DL7wuo//6/dolBhHhT7qNOVeud8D1blLC1FPpfvifkv4mWd4oN+Wla5mL5/0swGFy5nRhEdu7sfF
MOgcNIF2fzY5HSeZotasSLEtnq+pNrMZN+X9ssY/rO/kuyZ4M4m1MtAFzIztGhxupxETWeQIGSKj
hwIj+bxvMj6++KW5MoyR6Ij+M1eNVAglfDkIKrO98sEXEWNSQwOHODeGzCdGgtQfS+P21kzFsAuw
VL1DIkbbQkEJIOemDB50S8I9PSsPtYO5bcovKcmQp3PEgQS3EkmtKhDXvxoVqor9SRBhyYEhi5SO
vkozULxcip0rQd/8EVuhNunkUSo9hDjsWvln9ik03x6yuqWn2E8fku9E9l5a7LHa63t2clIEXc9X
7Rw39zi87eEihajiJsQ8HbkSecziG5R/jFaK465aeOLwZQKcKoqgH0wxFB/eBM63HgE0G0gThwYj
DfDdoWfuEaaJCSvp+o1EniK8xcypYqJdGokPNn5IUFUeedIz32n9rVbTIUJbQpjhgqJPRQGwP4Ue
X+VAyPAVEUpGC0p+LVtCVFtzIlnoZHAo8OBdaXEUSJi00Mdb3D8vh45VJRvPwmfyDxRHh3IAKLe4
vKP3m2qFnDf9pUaNH9yxsrtJNYxTkDDRKtuS14jUWEQ1yE7kWDXS1ksQ+k2bBubEeNsbIlvIVKtd
HAOzNyoMuG+Pj42rkopB/7FqRNnyzcWBh4dtYE6TL6/VrU1+xl1umVuG/Zp7u/iI/0UNrIKtQnD6
SgdfGPi2KVYfeY8m3PHAjWezFCockRDquoGKUTpM/cR8lycBguF0Hqx2KOlxb8KSF+qW6V7qI5H/
X5PvejuRChbQ7yb9iTSX25loon8/WINhrHOUoagLcGO5+tvSeYa6WVONRjYTsKb9v/cA5UpAWJmz
y4EMlqcXf0oUamnTfqM34QaqV0WHHrAUNNF7qmL+iOEw+NkejLFJCqYPh3X7vPdKWd/ByOBKtYFB
yBUF4vGtifbp3esvJgY5Y+yjgnIgcS5YU5WXHWQMa2LnZvdbA4Erigu2zloEJfqzzMI0X7+2CBQ3
KRro4mLAopeEEb8qMWyi3VVIb8+6NFHVM6HzkersIYpw+i+1+F6oiRyL/v49DVvGiwZHhtA3itge
O4EOjkD5E1Uos5BxRK/wY5uX/sGiAAcPGJVX5mvysjWSZ/uN1NQ4k0CRAWIAsk5ZhVMFhvmMakUx
bIbs8Gs4fosjJBzMrzl1m7pNYNTmYSvb8QAlYAoF5pFopPM2MW24xDm1X6yxGCwLxM754Iy+Eoso
iWUhriEzzUWXwqnfFxFohHtypyEOdwRgRgfrjcWXNB7UVNqEbYWWV14D25B6e09muPqrBOdbN+fD
vj+h4FxPmLPPLk3mI+4fjclpgr1/nhw4sUa2itw97JzbfNcWqBDV9PY0NwIykusUg4jAyPm8VfxG
cYQ5xFVCPBEYMyQDpGmwKypXnf6fxKuwpTJ/YpbQTo4NTqVZNZor6mYFsE1eToJVijQxlHUc6Wb7
QY/Mt2ib3IlPf2R3O8o3U+r4xq442aHq0b4pDgo2wZRJFG+fmhIqe6K1Jdy79n8GVm4IWIwJp8VG
Gj9wUkvRocPcGyZ1WFTQ1IVCf3p6+RkCzzGCPJdL923Cq+NyoVdYaVMksNOBriUNy1G1PpELVEsb
q1FimGpOv6ugTYNQtVAP/BsuGLo750WIVAijcf68QXgpIvyS6qoWdX09C6b2Yvo/Lzx1OzpCW3uO
c5ygCY2pXXakNLHK1Ij1SYULhef0iZ5NyE8CphWWTYNiId/pF7jkgHXR4O3D1+6nDsXnI7CXfohB
di4VCsikhBt3Vv55KPBJD/7R+eRrr0m+ZrsmozOq5uYbHCqK1GZ+1j1Fe5ZqTKOEAePQdEOFoasT
9XA+y73Tx9QS3x5svgafInl7F5bFhr/KQCehr8Wq4YMMyPETjMoDbF2VNYV1Afn47KymYA9bnaqV
PaWBOAKjJDQSO2vrzNB9niJi72bDBccoUIhrbkLB+q2r/UcTTex/8uv8Dr80fpqPUx2bRoTKX0H3
RAlKAcs+9Vu39yFEn3Q/Yc0SjkgmmnCWgpafnRhvSAHpIZMD7OtdRiknL7tkcVQGv9ZWDyA6vE0A
djy4uUNst/v6f/TZ04RDTJkxq2Rlaz+fccnywjBctzZZ59xE71A5X39SZWdOj7imUwfXjnqvmuVg
ItLTepBKGZ3E/wW2QAKWMlR6lbUlNHjcSjir+eozfY3Q/35D4CT2ppdullUtgwSd9MnyB0B/UDXj
vcojvq6rkJOR9+lYJUgfP1p5Pz5MTKMHBny/S16us0vXBHHYYQ1esD2I83eIx8mAz5hoskEF7DMj
izqlBmHY9OunBeJ68N5HNGS2frPfbYgfxeyLta0y4BE1M5FnI4LL6HmkgshStXTiEwg6d4PJSFFt
4d5+Ox5Qvh1IfZr5kAw20UiesH2ZHOU+VFAQKSktNRNzinF6HID0aW9pnlOnxiK/K3Wk+Gy4oJB7
dkkC94x6Butt7fYkvJlrtXOgA+EgXZNq8CK3h7nJ3Fvm4Xm2L59P9hKamV9taiZiUtPr9lY3C53N
C3Bh7wbJ4VKBRRau4kgW/t6JBF4UQ/nBCkpivbTDhXstUUfBwwaYVTDhi5FUfB4GStfD27Le4Zir
lBtyxzEv+E5HZl90HzStMJfrWk81fhzJ2jijHuN7AiUC20dmT3cYnzFtLOulc6NPqZv/zKQtwOwA
QLLLRGEFoheeAg61pXYlYDLlU5Q27jI3mOxHLQecv6CLTn2E67ArT7yQp8wX8mKG0CU6B+eEkkRj
jNtY/DaUd52TYhH72hXmedpM1V7NleeZSIXXxq7zDu2p8zp4194+dr9fgQSmQwGTp2Rvyc8SUf71
Acr0XF7FKUmnbAmmCFpVbznm9WNO7n67J5m+DfJa9kUKtyPGEwvd/vIJDb/NCElJ3SnIbacq3BSb
BQFGMq1V9SrcWutqhevx526BDoEu5uHehzy7whQrHuiDnlZd0A8Rs6j+7mwrvFF49odViCgXLZQ2
DJJwFSXFDYvE19kGxoT+ISKO3fiVKuF2xAEG4W27DMxnZZEwRIr4HbxDG9sIxv+uSj5gnHRHcRQE
ihEzl8XncK56PEiv+HcYSbUndvT5r/+vun9vIyynywVspm+uO82vdHRlbuGEeQB5BSj7HXueibNP
ACjGU6qpeE8yB1GfTEjtODZ8j6+icSL2lc0hJ0l2nZfwjNGSbOVkmnPGsB8YT36XMiKAhVXMApD2
U1I2ac0He2wA0/Lp8ztooFtkaw1gDAVm0qId2tVo7u+SLYsnwh4+xtbhmsgL/uILFlpsDmxnItjF
EIiYtFx5p1L+Q5fthaw4O765GyXA3yeyvhslO/gP94xPZ+WNVv5BadJdICenKDt9/xbRRdIoygpR
wBHcJEhYOGe0pwICFih0TEfTzC9KvWGOZaP+hv4wpIxVm0fFdA1fbBwsMNBHmrUa0w3p/YRnpeEu
tWe5ztqfUtorlFXjY45Pf7hobBSHlHqrzd0b8QJcM/1AuY35lTPehPmN02vivz24lKWhdV1426Bb
xiDq27QeC19gvabfu4C2UcakrO1n45VoWHDA/SHR6kouXzmqpOqvPBIZBkQXhBzqBnCAdOhHg70f
A6nKwF376IXUDF6tKWNZnqQtOkFmh7j5ZIfFVgXPcfJKJRCYcJZJKxMl+A9eMtEL8mAOSuOcpyL/
QvIbC0An5mVEngnxpblfPALIWr5PIJ/JPl0Hr95QuqGcX3LplPbDW2yrCPcwMcXY99zPBaqipmvN
6HZAE3y4+ByYW1Lxd75ZqdBPQhyV/ZxwujZlZL3cx2EyMoGypLlPh4efWHqb/0E4ZAxTCgIQ1mQq
TSzWdvTzGaQjtb0DZtgd3VCQt8YBOGkf8zwjSHGBrMDteVBefAr00kOal4QvbgiytqZnyG2Ka+S/
Pe7ENlIwnbe52BQqx3h5m8MUax/kJIY1Y7PWLWgaBqqhiAcAtQOwI3sepF3OGGRNkEg6PCi6jQHe
uLhYktfXzrn17S7BFtTVty1Nc/iquIRIjjFyUVBwSSQNBD1gQ/89rJDKU3pobvUBmpbQ78TJsgq6
PzzvdqTtExAM1LobCFaGwVDaVeKz4vY+yTHudej5cfPyAHkURge6cNgSmvAUSH2qNEsVfxTcY9ON
Y5Ol3PLm7LGPO08ULkQolux0iHVhtLp0qNi7o2+A+pKNKc8t/onT6cvSN+EA4igQIb/0iZcsCxiL
EwqL42fEritqSDV3rnaagwyvEu5jTn1gn/1tOInlXJm1cBcX9IVF+CtkwXowXqZSrGZTKL9KP3fd
DZVCrlv0I4ObXaw4adOx5bTbZqLZWgkzxnDXRWIzo3Ya3IlJZ/AbBfTY/3N/Jzv/pBfcAF5Za9A7
nNN498P0bNdAmZNgd2P8UVZkNYVlTTeYRfrI6Gp2vwAA+queAevEJt8eeJTjbzCBOr+cWC67joh2
Vp6gLBvDwQnWgMcxo6nQGd6XGiRE5JDtluAkXWohyJ1uUrKTXx9HVOZd560mIt2AH3pxubj2YW18
LTz9tJBFOK8XBmuva7QCh4FwhJJPZKLxIR4VFKK+TavKzRRuuf4ziDqPd0ZHGpX4WbyiiO8fjMCF
r07YRv/YY7gs51x/ri8WDQEVIZ+/scKrdTRX/43/zQZudDYAUyTD10EKkKg1RcrZqir6p+UiL+Ln
hZ8B3jqNv1rjjt8gSRUM6fPrvWm2TfDkPFYUhxZpvdN71z/zfBmnQ/WiL7PWyXkpm9hGJKzUjJ6B
QyrVYsqtu8cAgBuMTg9aLbUZdtmKW7Vq2teC5Ae0cxpMDEWZ8qYUN6Bz2tb0vma1KFJOpzVIOER5
9pR0X517SVptEEXffMTxjO1DPBR/0egRxxlq7hbP7JN8rsrc2MFJLQts6iyZ6QxoYsr5pDN9WRrz
ILA5svyD7shIi+YIo1He8QG3cIWFpim6hWFhHiafsvTFhL78KuIVKyGiQ3yt8ldYNUVEVda0onuE
E4ytwmnAm4wh/TXdtq4RvfdNpYYJwkh5YO7bp9In+i7An8kEWH3rkATY/6v1yHs/aOKbwsNrhS7U
p+M8CigfRLVmkzrPCPWeseo9GoecBSOHG5yqWnR9Kf+VI50cKy4ubSWQilBuA5+YFo/MsCkD1hBG
t0Lgg9ZLsZ/4pwU4X5EI3ZwJ5JVrubYmxJdnoJ0GFQGSKOi6yOvh0YYz4uoXxYo5RZ4Amq6fLNA7
JJolTTb0JvnGsAson+m21vb1E+GT1j8XwH0AS7bJ1xMUmdjXxZA4dz/2gsN+D1LSxrliUhyBZDHk
2H1u3MiYDGhF5FifLWjdZrdlbhTojCt+CXMUoBFWEzPdMtbmC5uwtmOSGW/rKmxNVhFgwrMXL9Jg
jo7pyQhs0GDk/O2M7RFVF1tZAewduceHGEzdyaIzyTx2L32etqbHv3pt4laijWX8l5C6xQ3g+57f
iVKSiy3KG6sHERuzG6vPFLDqjDofTtaJeiNv/5UiFJvqt4+sMarsqVLfuKPLSF/i+2eKDY0FjUfh
a7BCEcgPHYLU2Ibfs4yQKCbKppnqU5xUwu0EJl6Nf9gjCO4FYnsX+kvIMw0yInfSJPj/e1I0gAco
RAdq8JNlSTQ34EZoROTOvpRD37B3PhXjBo23ouyyYZxo40YFcOAoTzkvbeR+ws9IJlIGwGcqP+aW
LL+M3RY7wfMNk+JeaLXRutdevx1WyCZai5xsJ7QKF1GeK6tLmZTXcn+jT8A/3NxRbxBo5PW86OB9
cV9bJOEvtIdhV2qDrpkVESTozmwqZzM9WNb5u5QNJQwjmeuuSm+jON3FLGEwmSC7EqFWCBXte7AF
+HPp9YTXYluw0QXZeUfGK5CgU+fgR1pT6ewCTPQMVI7yoa5/leUh55pQ333II1uxc+y1JygO4DUR
J8ofQCK9s3GmPVrrL5Jhi51zU8EFO2C8O+wgO0dQmHlllX96880b4EXxoBbouWKsyRsacerWG15o
U3p0iewqnKcfajiT/iAzKJFVffVSNSpUjX+/ewDMUFOMEgEJfvuah8l5uN3aEg5xoSyUO/UIS0Lm
Y/6eNP1++zN5T8uGV3YuTKheTLplnmHnyXP8D/0/jf3LnA6VdZHG1VMdktNDU3IBo4ozh+YJkcjA
r2+9Ol/dDREZKXK7VfRyy40zyzDuRIzbBeqIvH3XsiWpMv/QTXDH9g46f6ejfuiy82fwgYmsCsdH
hT7qdpZYpnWghNjoN2jdCNmXsHy6H3JtmCnS29vdZTLBvImyi8T1KRDfrqDG2FEBwe3XpKreu8D0
XnTdE8N38zHJu8u//nWw1LZa53sT6cgfH9BGVyJdl9eUYP5GOlANmBrBvgQ7vdAY2kDbWGKYg1nL
IUykli1FEhjFliM7dJP/k89IenfhyKwWykEkAWS/9sT3Z8Yh3T6ANxNGn9p5HivONLTd+5NPI3U4
Cu8rStw0Gn+T81nn9+s1aRfg1PwnxpFRf7LBGdnUbGv1wsn7lP7PJpF+E/8uvgkR+wuIkllE/mhA
Wbp6KGSgz7SKKkxOiDDwGszIrrHXXkWVqdZ+8d6AAy1awyj+kfOltD/DfgB68Vz7zUlTBWZOP6p0
dJSnRwj4C/xFJ4uqrflSMpq0xztlRkOsxwvKfaCwTYXscvJOYkdAXuRDtpu7zJ7gQQZu2A5+8TYO
btb6SRgwYwHq79d52vTqw3Td0iRCx5ZtoaHnyouappwykfvEeFz2JNjAzmbgtvfx45wftzDUIsan
mMwJZHfixg8FpQg7eCkkzVDLzq1WJX3wi41ZpsbfHOo6DRqC4HldbmiZ35enuq6tALg7cWk0xLzc
q3qk/ySIP6mt/3algeV2ttlKHyvh0mXG0+EGvq0/XWySH1NGJeHJPWzZh7TywehO3JFnAU+zh1qk
W5kOJqlFjBRHxNGo4MjJz5ukqB1asyd1axVdFrl6DeWyye2OMtlL3Vf3boLsvkYrGoSMjBaJhu53
cAEGmdyKCrbjnD9TEqSlg29TwcuhPQr8HY/mBj1J0SVX8Uwa97HFI1Uh+3yRGaaZgBmEK5TWc8PU
42PvSYJKyT6XMgXjJcz1U+rJthqMgSStRM0Pwdtbydy/8WyOLNyEnl78KA0wMq5F8w0gjN1XM/A1
OhW/619uQhfjMF0y/uB6TSYcMXEohsdZB7SHWacQ2JTl/lM69fP2WgzlUW7i0xe15nEJ0b9Y9cZd
sZHF8bnybYR3viLEgkgwsKYMB+wE1g2SNgZaBt9aWmRUeMYYjLtamaiT9Eo+h2biy5yMWXzfomeB
q13Kei+/+NGECTNs8JKQSmp/XAMUYwxELsFiFmrmINqGx7OuxqQbTYpO1WA1qTreee4OZQhj3AOR
M+JHrahFdhTIs/rSnMS7icNCRpsKLVStq1Uv7aJGKKF4sk3x4w/IF6fYypXknMiMPZ2kSB3pl3ES
1ouwazt1tN2digQgYwWm/bOKVJStFndOAOs9SEz78yNahJMuHXg6OTFjZe1/XjrJ4tcaYPOyJ9Bb
pyM5VEI6xlv/nmyA8skyuX5uOiI+SF/LnhUMyKv2XoXf03Zj+4RwuuwMmUWdN9Pl8L3uZQfc17Q0
cOwfwZkDikL4Z2nDXlu2FLJCr+t3p5pVM2CB+rUp7mZwVNlk+mBuntZgrZP826cN0/K9LDYaOgLT
HEi1KoQw0wAdoLSfCmcsiV5gacdk1/KxKoP3ZTXsdr0hQPFRVgLod+E/Yzh47R3D9CMl1cwNcuNX
ru0ZF+FtHMSc4u7SpFB/rZYI0VQhl5/5ig2cwXO9vxFR37UddxLh9H/olixUIgMFjes7HiMHYx0V
4S5BKfTuuyrBo49COtaxLFYhC97rtfoA+lVRSqiKkNtGbtBmZxbTSG47uXOhB6wB1oboweiedPoP
zp4oWr+Kop2qPBTN/1m58v3ZfoMiTkKZRFuMCS0fVbVZqAG8+/Xei8opyyZoEiWOMsaHV+EJ1Aeh
dP8GwrkkWgZ+nLJrxDUdYqbryAVRK0W5xrsD4afUvoyRlmJtKuhfAPn/NG263HhMokJRQwVYHS0B
vTEQHvmpO2MeOVjn4HwwHv4jk8mSmw5K1oEthVWrngyQRtKaSJwbNmAVaNgDTtfdgTKcL87WcEHC
kFA1Y7VVD5z6m9JdOJA/vHsxoUn8gA+JaMu+w7ANUiFL56ilYIaW+fdIX2QdRCrT7wnjZyYy2uyS
cRCCOQXxK2d/C8QfkspjInwCpvDrCZb0ZkefiD3+t+vgnFCHVdlgpg8ZXU3T4BWx3jZogbhU94i8
+kPmiKuBa2VgT9JyG+v2UyVhRS/DMcEIE05UcnfFlTYDrEn6IKR3KxsYbeWl6+Eom2zC+b4qi8Lh
OQ0I69xApNSw5Pti99ikKHI/Je/K7au5tEZtSn4z9ESoxoe6xi3Qd/P9Pxwz9L5orF0oiF2+iM2A
8SXlFRkEfFBtni+HBvypqql3NIeEsGRu0vegApAU3CkbPqXP14OiNxpSyxv9j9sPkkWxw1T4PVBi
tUUbCCrsSaIARplW50sgQ0oLJzStCLvzFL1MvSxusswnqDK0CJmFWFw2/tAZhW9vqxo94MQGH/2S
HNX9uxW49NDO0ppy1yfBneEvQqnryeZmBj5p/uuDPN25dHM33lTKS060jY8it4M7mg9fZno0sB0H
Oq7iy5mqnVjoyypy8cMOKnM0YJt2kEd3wImaLIvQWRIl2Xx3UYsEAqOPio8Cxs+Z/OBHxZmEjUsn
4o05eYuPBLqk8xTR3dPYpQ+Z8hpNaF0Ynk0JGhxhHqhzhHcd3XcQAj20U8VVGNc9q1Oaf33UVMXi
XPAz6DmDgQdSIZ5hIeHSbfAb9rr2G0u/YVCobX0LNnuxbt75AGaIa4x1/mr187gw63vCIxxL35zp
0OgVgzFccMqNtQ7q66w1+AVPWdoJ3cj+xRPBEt5seKdQLKmbDCWm6Ib08gPtQrWuIrEy3R8+DMHL
RnBbPK0rbf6geeaZEv4XHN5CtfGKCo9KcQPF7pT/WbZtaJc657M/X22mIXSjoP1G0S5mq/LdIUuh
1VFd/NhMJTzflH+QwYhh3dLy7G2yxd0V+fKwr9YlLx2RORDU8FSzLGl3FjADB7hplmqSlwQQJqIc
QEsTuSSpBvVmvizXZeERNTxybJ6VFKJVO2SYf+ELhtCNHcCWFWI/KMkLHb9Q2a/rA+IosiqG30OJ
9FD7ED0Fj+/v5l878HxADmbVnMqWS2o3yziZ3cVw5EIIIS7sdFwGeJ38xQcoUaB9Yu0vXlC+3m0e
MCZjDpecs+wYYg5IQWe8VZj6I/aNA6lFjguWUoeUjO+HDMTny+Bv5rHU+ziwwUuYCirAFWUEE8mF
iSF/JVyUZhc9Vdnatf8D1zicTE1nXgbWV22jxa3pfbQlywpaWfs4p85q1mrSwh/+ojZlLMzwfAk7
dWJ0hhaGX0ndYjUINSffn4d9+fSO4dLtF3K/cAybW22Qq+1pjPrlshVnj8yxtGI9z9u+TTYwiBtA
TurgrJnjPkr3q3X5zZsknT/bsWRnEtjZ1mJ9FUz1BBS5qhxKa0QU9+V/G/eleNEvtjl9esn++Cl7
g3dhHuDqmQn94C6YWcocbP7Kq5QqMvObwgZpme6TqQMzZjw1i+Zq60Um9OrDCdr24cUvu+/kk22A
foXWzPTp+SGD3GuaEE/tCZGrsqDKZiHVzY7hvrzm3ZpCgMIPdpInsCZR3+A6xg/B2rS02I7ae59O
Zj+0OBW6XORUhrKDsyH5oLLpI3iU2cquu2vJ4d3Pm5XDzYW9Z0O3/1WPRg52Z3Ovtc1jDgdoLW2h
RoCLuHpdVWuy6ifIWtHd8JnRrxwlu4tN5B3pCHsnUuc6RiwIAfsqmGnz3Mc+qo4m4r1uDu48jEu1
L1kje1ku3/98ZoErSjZxMbdNVRLt/+onQv72/LL+qk/DT8lkL/r7A7SnEqLTueFIyveFQHWnecRJ
oNEzCivF4PzyepBbO+/ZcyURQ/2yQXhv8ZmrTdEAtBwJw/9gXXQo+V+8U3UV82o/Zr2CF+iF0ki4
ZTKiAhPFBmbwI3DfaZUOhMK/KHl2J4yALfXe0x9sAfKKz6WK9cFH9K2jN3i353QDkIFn9htrJd2q
dRdgfrAkbSKDmwJlmBjCr7dOQNLhWVnNJ4vPBF8njmxFRbragy2WEb68EJzeXx5zfDm+TmHG7bPu
5NlClNABqtP9nNcFbRuBLg7ZwetK6HjiHJw+s0U+gQy3BUwPZOVKJVkyKS/iqTkDI7BRqXW/j1gz
Q/eeHtMz22il9GQkxIgEOTWRL5CFcZHV6/tptkW5OfQTLMYhT9Zit7+d8x528nmZIEXNNw6elVGW
pYAnviTLgunHn9EmUMREJsP6Bu2/+A3qrIjj1FPxDZ5KylaoWFmVevLC0lnpsydFio6OxZH9BYEE
XvJVoKcUN8DvNtkYRh8gfosuqBcSoyKq27MfaePEvz6hR6b4iWhOLJCnzVzfJ/On9d19gbf4gn4s
np2WvEmNaxewrq3SWCUxzbSQqgjaAgtQC190MxW0x6KZ3t37thseBvbUtQIu1hwFxVMuEksIcY85
YazkHWOC9qVFdOAZxDTQzM38RyY8IDJLH4S0s5+rUOj5JxaoJZWICm3DdgR7C0oJoSHIYCrjVPzp
OCxY6sP8RIc4ryfBCqe/r7x8J1zFweye3VSXDjVsq5uoPavIAZZLQk8ppLg8BBXflKEpSDreXDeY
x9tP00Hvlg6TMazVbDDlcMXf3u0PmBmPsU2c87wc5yiaXnWNCnWSMoopEB77NVU+yrKzX7WY454w
ChriKoRfTvGgM5xB59eJoeX9BecVhmZqUw+my6SVSNzshHcyUWFdlXOOjVrAN3Az+sEQpSFa5v3J
IBbAg0wlcuoc8P3uoQky5mplz3ZLUPS35kQvtA1bjaxq9BVpHiXQF4F10AEcjc3Wce53QXR0U5cc
h0SMbnXdGdP3HcO6GzL78Q8meUqLXA5ugFSFDL6HKBSG+zk55t/jYO4plQz806P+bhrydJ7O1p99
LD/2Mo+oWT5mdtoZyh0Z2wmN5CwWGOLAUY4Pcexv0HpIm1joDthm8x5CDeFRrs9DSwnoFDKP9Scb
r6IuB1umCPRTyd81206b7o4LpgO4tKI6d0QfJIr8cUhSkDt9Y8/gmcahdP2k9L8SoyfiubOn/lJZ
vj/r17b8oRBl3VgDiZk27CCl5Y+n74pfHGy0xZAI0MVlHbtNVZCutF3arUQ7p/pOC2peUk+ooATf
0vOVhLhzzBKIWNBmgpk4JNYvb/25mLsp30YUZXIXzFIps0M+sPoKb2PFMKgNynt4wEzgpH+4OaNL
t1I5e9Nr4bhWA2O8a8Rpbwc9GxxZA2vPwFPJln5pIm+EYunZ79gJQZpYfY2sWX881BezlMWNrRj3
UY4xPxuNT47Xnm5uCOCAVmM8YLHsNX8xtwFJJY/RR3ylH/NjQV+GFB6j86dnUpW5rIII4h8pGTAj
E7QmtHuarQ5qqoCGWj3S3tPCQyxgVKwbYTDH9ZLGW3yIUANbtIYCCMy/hd1xn+KqMNj8f+Y3sOlo
JwXN8R9nISvqEZKTpXo2mDgERbFe2qgtGJVuObJ89yJU/3WVBCzsikSK1JUeL8ODrTSB1/s6jCDw
PbPu+EPKPQGU1DKKai9XGYKnT2zWTe4moO7g0sCGG88b6BCgDE/e6ws8FsOUgiDa26S3apsNpG7Q
iNRm2d8sqqd4HA7SMxqkYjXX2QM30v26LWjBYJXhZN/YLO0YyHnuYREoPXgl/TWgI0xWI+p8crwR
ALd9B1jWF/uXO5Locji8/7sJRuv+FpZaOETjiDssWtud3b9QMVQW3rGN91iLeRhyLDgHsq90YA4S
q6UNuC7wQ074WRmFGa3OeQaohqr3Ejhlu3b5oe9YcCWbDoN2lnBo5Oz0XEUWAZC8RbbwKj4e/cPW
9czna1NRQw/ZxIIgy14QL2em3JVbgJejdNUucmKnvThgxGv6utEBJ+7imwTkTLpzN/rEHgzaq0jR
8/AOITc7sqYKUCf7fAzi3ETOVRCzB8ke+zDD5wGMLKz4hIa1RYuAFwki2Z6h+XDJ6AF2DdG32ges
RROw3KmnDwX/70JSYiR9p96ggTyxAwLs8P/fjjk2oVsDWcuQ57BVF3QXSSYsvi90DU8qe3Nt88nf
No1k2yHJIkDhLXy2iYESkRWtDVwRF2cOT3lfYh7KcrhFJN4oL6alMvnR9By8cAMNQFKTgpY2IL07
gWOZg9QlDG7T1z8T+p8vDMmBsebykaLrDBwxGfoKxJ9fsvjOW2eU0fvp1XfZP+geTcV5OBiB/YhH
YnxiEQ9qFdkeu4xNw8FTBIN8tuELOTypHhyZ84U010CvixTUUnCuG2+aAnGPaMnO8xPGXXJZdaqS
MSSodsLbeqIL4yU2nvTJ/jNp3VzQXEQR0PaLLNTrxahtGCYPGhURYhrdlogg3vrpTaxsTGAPK4Wq
/cgz/QK7uTlFh0WNWwHRDmQe4ZKlkIRJnegrTsXmDdgX8jR0Dnf8DQ9PfUfRdzphMNq3LB316//0
qALGgpUHViyUWessj/ocvxO/cTZEmiFpJBQ7HJ0evgvBWgTG1jTntEaH0+nKfQmFVfUIsux0b/SJ
DDziH0k0sAlUXRX//YKp86iCkFsF/TLIWzkKEFrjvaCQD2Ux7vc6UnUSA+xDw8MMGYOTuHCkiowW
3U8wNv87KxN0fiEHg3NcrDBwdee6KfouOUNNe97GXbVcndV2V4ZNT1kLIOuidR7DDqf+qR1oESue
Nl3UGkD9NFEsP2ftWoY09gwiAvCVYYgwZOjWKy0aIbVMLj6SFQDrSjWLd+2PlDcJp4GENOBxx6VK
t4ENPjrhjrZ+rnFiOxWqF8uJX7eOZdN2pnq/1FWVZOd9g8R9WEZFZUqXjspc+nYXgQMhtzkB+s1p
qEy3LSy4O8CZLULgBWnNh8FSJSL+g7kbmMPDAe9vkT7AY9uK7oO89qCHeGSySGbb7SdvtTBqPE5X
9aSdJP6pYuoe5j8s4HvjIOxS+OVPPaURgULeQeFOBzcHiWGnui61myzR19KKLwYKI8spYZh8dxvh
Jp8Z++UOM2uH9gkDtFci3r/JunqLra4vvx2I3HzOdKhQDreqhOg9VOzSJmREnl5d3CqVx4mIUPi+
M88O8jemS/nSDrfhPiLgll79cOy3xQP6Z/iz+z/rE0IyheKRjLq+5rusd4i7Xe1rZEGAwxmGHJ4V
aYXCrulvRa+MX330fxaO7Bcd91aiLzhzxV3kpVyGOZ/yUqTGfsBkG4xWsxCNSwMpPfZ/fCkAP4dG
+Ff0tnffeNm3yQZFIe099nDQRyqwvU9F+55AzQJQ9j4Zl8dYAf9KiH4wwz6X1B9TaN8BJ65AMyqK
/jCqAfv9k68lljSUgMs9HMtd+cHM9E3CzKlbgkvzc/Wy5aDqNWIyGXV6ihIcf0xte0CpsS7cGFba
j3l4waPvJtueu946Iqrs2Lc6wfpYzHC6KakoPDbpvL2bkrawk8BsUDRUB8Og/S4Rji1oPyRJrH80
mPwZ6ZETuu3CKkPPFpN3dyMpSXB9XUQTPaU7tPURpYeWAtasfbljAc47xODoNWTr7RZDU8x+JAKj
okzcsD3Ovad/vz7KPbYNj8Zt6HlOtfYdmHVFDHKu+vMIx5VgLiNyJ8kpGReGkDTjXdkphIioAcjG
IbUz/4jTPc/d/CkxuKVxZUnir8ZmR3vtH8A63FLp46tR5bh1OpP6bpCYmNw3KGKh0lAQzHD1py4k
q0ts1/1HGrvZLbD881kgizFCOhmm2D+c5xbQj+r8NqPbvpLU/sYGYUN7duwj2mQOXYfvfkOMLe8A
dPQzBT+ryhw1IbqO3sSSGWeJ1+Zu/VjnmEQHBkIqAdx+mTXT12X4XJutWccPVa7PCH3FVUc4tHWU
AO0ekX22ytSK7+bfpxgyxBi/KNCTboaxsw27JZc80wwXsJcs+7Nz5bKRPDCOVLFXfmGnTSaavtWC
4THynRimawV1WHnJxRZcnuXxyapPoe+w5dYwmsqqFdCqouZKXXQP74lGl/nhWV4oWH5e4K2fcbAA
7E9PeR5HSCwcGC4/+5LDgsVXgwB3SNkFtLBa8laivKXQU6DPYckYeiQugr0Hd4zbafyOKVVdPCRk
PZVbPtb6iZEzW1PjvesYCqV6GJV6L0zQ7FA3ctL2SYXT5avk4sfIj4+bwx1bs1EV4+afTZhjevEs
5lROro/x8PADv7zCfi22nIsz5bd8F3ArOoX7UYrhdee7QqRrxg2CJSdRw9yPPR484Zboy0Qlt/jI
itIHm2bOE8ivvujxgDChcLejTkNUaZd84HE3szhiRD6XFf1uqw6eim5ysQEGMSfQlU1bG1YtDYlF
7kZRBi/CneeG0th2KzMZwTb7sjVWijDU/3+EPlHRko1vpiaUGDD39HGa9yeuHvaOuPDzo3PfTF6Z
OiFpnvusosZOQqooPHF3GRInaduvbNAJziJzk7Vu+1K1nXoroJ9EmW3AeFK0djiZVYzbNepwoNFN
ydmmE0y2y/oj4SSlkfRPVM95ifDZtouJRwQl1JIuhonsOPIQIsDArm9QVMt+6bMUiTbBEmiyH5TS
WpyO2hQYdv20goSKLhdLdv1TCMCDaRbYfs+3mtbj2Mn5fwruxgfZwqufWPwRsn7WSXZE/T0cR+nS
hMl4iiiXVuQlvNay3um//4nGQJ/ltTB+A2+RN1jxM1edpUfbiHEuTDcLERu7d8H8HPtvcmDST7fL
Bd/bfDIdfiDdtHfOP42vsknp1N90jT8FWfZl0+2aE8nFDHF21o4KYCHmqsbjLyfUF6O5heQ5NG9c
Ynecw2YwgALSNucwuAd4fuaJCg71pZIzi6WBnG8QFVVGpdItPc8Gu7DgVyrWc0Qb/oOKMmDMpioL
iqSGsgwVMIvMN9SvKVb2/40Nr6qv3w6/2s97Lo6CX3N6gVXe/RMpL6KkgGuTpp697tU3SSU20K6b
DW0NyRpZyPkXQSVkLG6KMQZmk1VepxWWgM6sWp7ZxdfNuz+K4cyKYKMAQioeU8msteiRfd/kz1S+
CveXDsu9m70DrQ0aoJu40P34fvMXBJFCK47nDL45svL4G7LpgYpRXJbaY3f6lrA7OVyrM3rXCOA1
B/3bZKG48ATq1AQrVqbV40sfdhgnBWI2+Vx4QpNEVE75ZOHEMEAh1VN6GRFvqVo2tqFy7bEUGd82
z0Op5qlwLI85KjKNjvoqIiUCXuU9bjxWZ3Ogjl0zc4/pQFoSkyS8Wu8+gUx3SxyIzTvTqIAirOa1
oFjOIE2cjqIWu8/weMd1pZRkI3pMssfIOqmdb9fwWPhtIPsxl3VuUher82NgYGme12yUZmFAt1jy
NYSeAsK+lfQW0+iTvnLjCInoWtMhAG4yOqJ++BB/gwMlfkx9Em6zsRkPM3e9ZkocygUUbURmtIaC
pkgCDx40xFiSDIkU21C9s0iooO3P+cjy3j6gn5f6ywCAxW8U515wJiQv2l3fpp9SK5u6WS+5LGW7
JKCj31LGBkjy1SSgHN4Fjj/5LzkMisa7xE9Bzsp64pf3OwyjaQhQfSABkCty9cUIE8XXbjD743Of
OOwl/itU5BARxox8IqvPZWtwcgCtPCTnL380SsYy/RiPT5feRuJdJWs0SrRGMd9Pm537E0EfFzTe
zu8hpaKtIaqS0csXWGerI3GrrEsnhthWJT4g9PzH/8ra7a+x/n4NcI0rYnMt2jrusWDJHZMBR9dW
FGbjc7XLygwsnGibNE4mKSFi70jXu00t7Q8rUwWB6RA+cGRLKpF5G8z5rjGr5TVb8IYF9K/G5qah
O7Fj+FaLRRgR3z0ehVobx0cDj/6TqS1UUhzxtylYZ88TOMTeBnbUPJBU32EEarGU7YvMlvyTmCld
oAee9F5JOCxPqFQOTaI7jiCy8b+L5RRGVv1jV1XtOoVfacd72mgVAXYCyjW+o0B0xYlK7pCceXXn
Ws8+vTJtJtc8R3l7wJ9mCuvEbb3DtAILqahGHgZExzEjvv2aCzdok0hKs/72hFaFOEaPUYQP6iOs
1mWv8J8DyDfunvNfm1ui+5Fc7JX/QKnHpshTI970uzdd8Tu/H3LqgfyVkzR5uIm7BbFNl2Wmzcs9
NXcMextYoSAdaZJOccFRw80dd986BZMqckuKFqAQADIyTpqhOcV0HlShoAyGNosHBEKlxyRS4LV6
suARw65YriV3pWs6JvWSDELSenTxP4Th4uQgtj0+Aku6G1tOXV8oPHtHj8l9J6th4CSazBoNx6OE
5j1yT/niJMGKsO+9g19tlPMGmnUFn0KRjUjCTV2CSHZiv1nNeL6ygkvPysLo5U/M3pep7ZOKT2jp
o68o6Mh2faoTXyRSuQeoviirZmNq/rFoaQkLpxUfp0SNfhketHdhcCrcJcywB03AfWh4hWyHWDfw
MxrX7JoxyDWiK2D7SF1C3GHAH5gf9iGn4k/UNt9sy1uDbTyg3B512VPKuz1HoBAM2Nd8QqqKR+FD
Kozfmz/X+S6mzrmEvveEah2a4yvXUZPPULFwRvMK2t1QxMGdz8NdoTf3hhvuip60kDQn1aZa/6sd
dF36XBGLILb2+xPgujiUsdAgGE99NusZiVaP2jF530P9zWUdddBKk2aB8lqPnn3KHZZZ34vz4OpS
JJpgvP4R6VKBiurXUHoqjAjpTXNCJMoADNZrS0xIeGIKQgcRoiQUeHk8y0otWd+YzVPHmqOYNuTX
36b1SyHy7fmeuAsyOJJRfj2EOYIUa5qm6mHUKwEOLOgv9wzY0SmEd2L+ElfWFvAz/qLydabY2Wh9
yJMQVYyCZv1X5EPnScCbSuPXhTkwo0qfEPygG7IthwEyMVQQZopd/mxG+hS0ToY16EEYp3SbY+aL
26AkfOYNl9qxey0Q/kEyFymgJunMiA1+tz1v7fonSi5vv/dv7vF3OV5MHIXvn9oqi3TKoR+utNAs
zxTBsdvvx/dsB+46egF1R4x7N+nn9DykH/ickeY3fORgsBSzYtr3gvq2mR5+mLLWojHLFRzpfczQ
U+XNXUOY+gftPx3hFbsbdMx0HyJcQz8IrUgPdfpdP1a88nLpiHNVz4fc2HO+oBqedmvCzI6Blxry
4SkviJE+SDIOkWKLOgT1kBvGGVAibYhMFBDak4diuYKlgO026dte1vxA8dHVO5H8jhn1vJBpNZb/
BYg022ffKMVYPeBY8gLwc+AiM5xhyW+tKx2vIbjcSWGYI0rDh6SjXHKtGHJgcgHjBKdduxze1Y4Z
bIlaRy/LvbzL81P4cU1A0i6s5XeIaauC6klfKuzou2tbR16W7ulBmQ6tOhnQMrk9jTbkrhPaYNfx
N08ENH8DqHGsF6056CK4+VyptpwjaUahoKUrWwKBi+Z8SY5dG4Mz6at7vn9TlSy8f5DTgb/KgI+b
FIWQcWliv+EYen4wxT5a+B08hUMWDnlCGU+tnwFhOhjp9BDCAG8+lD3cfH99o662jjKTeiptVt9D
Ampsef5m7goejVKQTbzViigSGrLOAMWUcFMBT+L+pxIiZHUpaBy1BTukAQaSkDN68HC2rBh+17gj
J6WT2vywOoNpFHFNQWYoNq8rR+gVbwZ2epYm0FbSQ5YecbeSO3spXIqvHLhWgHFY3IuPW7txlQL/
R0CPZ6836F24qUiF/b2r9tR3/TFk4MEDBbDfpJ3cCzcwHMoDh5/Jw4xNq2h7PkxhgEv4aSQo6y9w
M4bm9/Ve7xqammBRT6zYOcpr9a2C9oemyqpbFb/hHqIk2saeDeI4MT+nlDfxiWrblG7N30O3EhwC
aEPk5gb2XNfu8qfdsyaMk4y+RHCCiYo6aTs/MCgWWlTvLaoloCRhMytrA0aMAlw2VIJrhvfswBYE
HFPfy1QJPqEp7NJUXjHdyWIiyhGdjXzUAoq4+aiWDVIxusx+r5Eh3Ku5jJjpwe1bHwc+I1lueATJ
jtWB2b/8smqP1fvBtJmKBWIc2+uyIcx4MoT35C1XyB6rCmcWPqhZ9jEuyM199sKGlqf+T1jLvwu+
4KhGpIEGJqK2tGk4xqWieveKFFdG5Rgj2znIEhskzx9yu6O1FfHh5Q/QJeGPnIpKYOXI0YBBFEcZ
wOZ7JkwPAdnfGeI//DbrnMiKRzJKS19p8fZJQ4GhsS2nyNS6fe/vtrgKJJzEslmpEWlUBwUrkV1U
t7XsOTKW/4Wj3/kP/YMfm7zK2MUyriX8PjF0Gws7OPmNpqJPvNjA5ON3FWXLT7UPxe5gRnnqfZtw
0NPmuGFTuWOd1j5ncQ4/UKyhL0eGUjYwz2CwBVFUYQK30dBVQ5GyMXFeoxHBN9NOkg0Irgo3HzM6
shwd5WJ1h1AS8cnsmnm736X7LKeFtqmvha77M2RcuAviWacwsQ4JZVyIWr72kSU2hAlwE+rUVaVF
rwssgSIGEY3dnd5F1LJqYHsVXexUq71qLZvzxnusMUQpKZodBN80c23qITnVvGqQG/69huPjT8wv
zNC110D5QGm1JbV7t1V3BE6q4fsXSiAaakQK9mupZDUylUY4T+9kjslXKkG/a2ASR0DGcxiIDrHs
KFaGcG9bijSitgxth8dFBZNMxRcyp1qaXaYBBwzgE9bjqwaeuJo1BLPx2ghrtV00yqmwCesd4y5g
sipTVTtiHSt0viAWmO8tMfuty6mNtWd+6IwDDyibmSGv5+EhAyKeKLBDSWm89u09w1V8y30nUtP/
EHn0AeQXpWHIwsJ4m2PsIVk/qCpv/rGEjgpL59gEB/5Gzz5U4Tz/GLkMmPNYQ73fHAsNNWXqZjEN
whcSnn31dKX6M79iQgeLwjLhgaCD6Zu5KFZtcK0wXh3UZ0SJbz/ZZLBfOXKMzIy5caA7Kj2r3PhT
YiCrFXloO9U3A2uzXdzYD7V9OyhtXMPCNjiur6MsKrqbZCWFreF4qLB2gMYKNeUDhxBV9vks/kLl
MKt4Jnw4FlZAiKYoDhcHx5qDQNabmrBm/xIzBR3WILFx3UxywcSOUOYwphpIJkByan01l9ZQpG5q
zbQc21dWiIVGp5j+HqZ13saWb7aRP9nclkqHqpBONBTPMUk9WAtAjvt9beHZXnLLZklCKrwNtFoZ
Vf+NDUyglAkct0aZWqDBH1p8TaueFI8OZ8/eVOlk+BO+qBvjX7di5zXuJljJMFunhvOBK5kEaX7/
ZlZKLkrHbWtFvb6NajbMKQ3zkvuE6GlxMlA7bE5df6iRpRZnxWsUnESagHE8oRbUYho0oezXa2AN
ce9fs1jGAQnx+NggANbPf7xNnjNdx+puOWje0CisNLIs0IRaUlZ4i+ciCN4LksUaKknsiPsXcAeD
XyP09lV7rlmHFnZJA0tCg+aHPJnOBDIl8VoKpJsT2QfSjrZOE44kxyzaZuYPsBJLaVsRvBATlkTY
n7X9gxZi4puKd9M5rZXhcSgf2opilQRloV7BO10Jy4PuyjxWNzq7gA+NTOAa3PVC3e7KRYCCz40j
4L7s1lNN+dPgFkAFWBdV5ieE64/giiZ6M80PzjZP/z2ZdH/7KHVqZxO/1JB16ZOPVJIb5IdkFeX7
h3oZDD2uBIyLUTmlOQmHUfdI6WzudkMmOcc9QqSQiJ2YnGDCGnWF1ItL105FYIac3vyNtXlaEa5l
xLyQcmNWxHjzus6bFzCeuerkBRA7kvO4EAR/StUiXR03SD9+gpi4ry+drb0tF0Y5dK0IusYyFRgv
LuV/D4z9VfiCq3z1FVYuE8y3XKHS06JVRuFH5PpTqn0MszErk3eY4rzfdW8YH6Qu5JWyvavnqO0S
A+Zh+fIL48R8OHRh2602pTLw5ZbDVBe+rSGV/UfLeKMwD8ileMnsz/RvFQpS6zdeVF/MDP+pd6RJ
0AcuYT9IJfqeAsdfccKKfcu/xvLmVdcL6azohWia2p+WpRpqLnFQ4PXsVuHBXD60MbhdD+QE37KM
s/PuRFu1lnrfgxM9s085vS7GUBiGJE/v/CZE8IzuewWEw50zcUmdee93LxF3MkRGr0v364gjcC5W
0IvCnSne0ybegz1VyODBnXfi/hTMzNB7TBgJgs04/6v1WtKWFL5OrcNIA6ndVn2jHSMo7CthidoC
6fVF1zL75HmXc60pAeIDJZxAVPJwZiqGP1thOR4ZC22oSOvdzdBAPWQlMSIsEZF2WAAPWpoUYs8b
ocUQRU1CmF+O8pJJL+4KvPbzJxwfViaytQGqyBcaOQsUz5ss7n2liDmv7V1wfnik+g5NSOLth6SG
e5Yhwl6ht41wKtn9F4GISeHkXdgeewNvYnxSgl8OU15omlA7pkhKb5BjRLL0FgYtpttw5cQp8Ot+
hWIUSFxMaHXRR0trEyBpCrwHQbQwIAFfWX7O/+fnbDyOklazDHGrAHRVJX8uUTXD0o3gFBJiRDFZ
iJA9npy5NOEuQAOTiVyTzeF3Stp8UkTD+0K/x7wVDhyNZjujNNDazFtW31qvj7O88mcWa9fOxlSY
CCdjZPEdyMnb8wGphiCgzpbQlexDZmKHLNWe0Rmu3fgYIGbyH6fyvO2cprAAsmbqCKPsiIj/1E8t
66hIl7nY9Rr5daCo6uu2quwHqCcduCWx6ziGuoVRwIYWg0Adt8Gqdw5zXPzxpatZhNhRYhdB/Err
lnQmHIBnTWrQQxjRZL7NyRnwto+Pu2+K/Tlv0KFmYAFtmo0FEtq38ZNX42Af3t6CGRaLv/GpAiib
H7KTnie3NASaPv0QtN7hI/ggBPdxdY7zMQBpIHfXv9TtNyGNfXcmChXo0xIzxkMJlWSoh4DQygDb
I6CHzCOrEvdg0Vd53oMejLOxsuJpE0122q8OQS1XsSIaSgohL5lFdLyzhDvXV+ExF4R4wFPZXNku
0TNUUf4tROftb8wtIss8VNvacMgIe5NUIPYHg6fvBYBter6am0zq87dbgYzzmUaplYVrRbKamdOT
eTdlBZPIHx5IHlJqP1iXhG3hwwNjK42TtFtu/UpnqohXok+vc0Rh4Ik2i7og5W2X9sNUM18S5ApC
k1Um5rLz1f4GyiNfLWMQWb24qbDgW+fM+dePya2WAOm7W/3/9IsM6Kh+mxbWvQRjJGyS6teUu7N0
wBawboFJ21nhIfn0OoHn9awQh+zjXz1yCF3RKU+zyxEJBDZaY2Zv3L6UldgvMHLwQgIw3fIG7oTv
WHiu29mwosY8e5D0ky0Wy86uxRz7HuqIi6BPlkreBjhkbFWe4Kd0yYwk6XeHlwYHm9m02497HfsU
TtvA+WAomwBsQDK42uZIbkk8K682E5+yxqmMjRXqFLpOGvChulOk48Li1ZCLcSx5u8/THaOHyNWl
Fz19iu2/g8poM0/8pqFV6nolAvYa7+9M30MlTz9IdMQt5DKtK06vuuE4xHbl3MfQbCgz1AjuqcxX
trJc3Md7leHZ6QanOXriCPnQinazQDyUYWxwmh5zLyHdm0g7kPbEy8LG6zmQBmkqDQz3D8HXm/5v
0DaCn4rPeRv3L0EZp4mupmquBIkDotbUUMJyCX6WDhBhYTtFmB6Zki129bg2C9GzXqnzJdoWSVjs
jY316ArDPjiApQU5n0j5DHo51Gt5k2uUvwmlRaVQC0TI9+aQOC2jSc6zytLnBIlaKFDDwjhQ+kNg
aH4B3x6oA03lnNAJmM48UEbHAwRvR2zrU/RWARYZHjjyEsZNUBT/N3FC0/XcFJtSBL5zRnWLRORz
VhAXkhwNCDTxf9WAN7ioszEGCc9qGiJEtLRcOYjS9nyn5Jeq5s6E8/b1qbJpzaa4e72pK/nWG1Ae
ErMsaiT6NwWIJa04NwEWMKHfzIP199gp3h8mHRIhfh667FCekCZW3UJRiMG9flpIxpDbu0Jyryuv
BQoawbPbS/MK2LIK7v+xYXXXL3tC2QcvB6woxAnBdpWKs4RTXDxs7/ndqVabOevr7NBVNCVp26F5
1DUcuc3fVqOxqwt2an95/6j6RuDOvhf/Rl5jMxmNE30lcuFjkpyx8HLF2Z2ZW4J6duxY4ZAcKd0f
WkIXKgFQCve9JHe+F8U7d9JDaSPIRjuIgn8aLJ8YkbdRwQxUj7i4pCuGZHmLqP2Oun7HimsUN+/T
Hs05lkalIUePCX8XL/d4qoHw0znuDHfwoO8nrz8J+lD58d0PyIIA5oP4+f09O3F1PuStcXOs8/M1
+7uwRLY8pifuVHQjJDaso2ZtkoRKCDwDkZu9HmpCsswT8/YQyrj/fFmAS+mrEUj6YWu9X2x2gLFY
Dlm1uRE52kV67KXS/QhbzWflobfagPe9R5ZB6aY9LJUpbnLfL2D0xLULF3M3tqJx0BEx47mlneRi
7xUOo1kwcUuFWYSojkmfiSloKF3V3eSC60sdIUD+j9Q7yHtT2VgAbB8iV9HaVGqVkZfpzk3F9NNs
FE9OqOWVH6CJfZuyTkp+l249tuJc0K3WQFiduvnDGSOlXn/KZW01nrDbrestRmnpfFi/A0oYFtHI
g+KrX1kYZ8ngQMi/HPeBIKkCbGbzZ1+PeSrbjpXu8vhEB27aR7++g2PF81Yv7+96paeOVjrWSh9K
XRi65h+fe63fgx+rFJ03Z+GQV4Ivyk7oMecW1kUVzdFgnuA3MWc27jbpRw+uFY1RzaEY9UKUm4Uo
REl1+k4Tk3RhYEcFGfJFHT1bIE4mf5pqLxPdvqPCcXs8BU1zOkqbmpaZFR7VMwl0QtcAnrCRdLAh
Cysf4PlAexN3dSZ4ZAZJ6CBWxU3b6vFbK5okRmjGjdt7/O5VmXkmFLLF1H+yD1N9SjpgeujqJc+/
tORkRpgkCgxp8bRdHF+I/ZKEmPUKQgD6kqDnez4gdTY5XRQLWUA2PnAZYArXCh6xbWsZwDUTrFXM
4vQVtdjvLWI/oZ6EOGPs+nYqfQrm71kgScXfpiJg1vD4zKnBn58jCpFluw0du3/aJGDptn5UOKdi
H5fcc6dBWE28S2v7z/Kst5ttZYQhxg6GacIaoUMvb1BNfb6s8Nlmxqu89+7SxB2iTFhTAuO6vmbl
K1wPjZzcnTdFnB4qmME5a+YqtglAENpU7tWf0qRERAn+vUxTimnr7Gpgz9COuqnYxYCTdN4zO/Ws
8hRpc/ItMp5tm+rz0uQCQa7kH+7xgKFo2tyCiHV3o+FEJ+6lq7tz/LubK/f2GIXNs3AanodvzBBJ
A8qqD5AdYSBeqd+LErLjlg/pp0TpH2baH8GONoA8B3WXwsB3Zr/WC38UP/viUXt+bytWbv7ETJQd
jx1THDVACVNFgCDzWDphTfAOd82ICja9oj8do9SJ2mZ00kWCpf9bxYwVU42ojQMozM+t0ydJuV27
dCD1Y/D7W7XhEilbED6QpmbYvlCet/ULcIoAqNqN82trNsSBTJvjaGBkLjiA5GmE3tTDS10xUnf2
7ZCPcwzvBSNQJT5wQ8eNQH0MQPJnnBkXl20L/2YB71dpl6yLUcnruNGCMqBF3Yw3VRbGXcV4hcLf
McMxuSFra55wh/OITFR7ma1DPRoepKmlzigF1jtA5636veaL78MzhAIZR4qDrMYYIxXaodLUv41s
a0kvi54Yq1Lhi36RaMJeOx5kVpH+Ysr1wMK0kElqwlt3E8yctNTiFY4y5we9CWKv65ePn/rAT0l9
i1TYCz+VMCZ5Fi894VXtTFGZpNFrCrTLWy5Q7s4oWCuW7VTeNe6tR2PFmOU9sTtj48MBgpF/Zhra
04nvL+0EPMtb+mbr08sHbZPfnhUEjlt07kcbsDnAbGhJSkABmyaVk9ujtmqVyCiiL60qtqJPEywD
D3E1QoE78kaJK1c4Phv6J5lAbcnkK8iemuHf+DWyC5mFQhy9GoSf1eF9/ipXxijNwVpsonUxa+B2
Y7/KrrKervhLIHslZYXJRlYP2Jd5IVzrumB/8cdilFP2qt5xfw9pMWsKsPmVpJG1YepblW/BOel2
m6jvKacBXXHWOrhfC6Zj7XpjmwY0zcCeyMHPsK1QKo8IJcE9Y1bTeD5OhYlgbjy2f8nWFTFU9478
GKLjL80TDhQ4jLeii5Cgvo3Vi/qC18F3bRerKvS1PsGvPzFsjy8CnVfKRR3qYR0cQt5zlqrcnHil
YzEvkN9wAzzgDm2P3vuAH4adHTJEvMvGtSPnS8HEEU0VPiIiCYIEtqDDd9L24idTPiHIC2/hJEQz
SYVCZ5w1eyHogNf3E+HgksbLD0Te2E9P08tPbhwZsC8lba1yNHZzebhuM46f3V9HjDCtbkWU4f7A
BYvqj7BHEMj6zrEljxcxczuJhHwcvJ1c6DdEpmQ2/OFRIqdO6MEr5HBLRfGOe8mZt45rsYVLbpjP
JM7MbOTxWGnAtdoOyNi1jb6yNXbwi+taQJ+MW5yi4Z4TOVvn4VEh0QRTlXuc9L0JXX0Of4QMosf0
yexjplvNFxoeCkvxyFfjMWyywKDc1BZ5DpEZ4yCUsUlUXIlOux7QqW802A/dJ3+7vdDQQOPNhxhs
Hmq3i3c2uSxoiWQ7VsHfM7/sNavi8XK8Fxw362zmKy6FY7w1RotnSn/Fq/U+m3+jxA+M1nZ6LWqS
z0jcOhxB/IcU9UZcJhOCGZ0NEqWnYz/8vtLz881rFDWRu5/zigrR8rpOhB0wOzbTx5hSGdO2fPvZ
w29QDSZ7hbPrmA4BJXD9lgfp7rVPhq+5lhXUFztGMu7Ytxj1rNvLkQwW5JDiuurESqgm5TAy4QP1
kprvc2qhIng30yT40JxNqrxKYSIMOPXj/awbVySCc2xy2N/8RU8G5hU8pyAi8MNiYD5nPSSkH9t8
JVjdLW++0agJkOr2ysJ2OgFTGy7Vx8nul6Bsg+oYiJ+cOjH3oBYtnGquIQNt5RQqBynNSyRBTRgK
O3HGodNm4FC72IaYbsqUN++IC0ONU4dU5Lu8zIWfMf/TwhtFsFsu1meLlJ9un1ajmkjBvS95lhkS
8l/Q5rGQkv/TRhOLuiwrdJmHRzl1mnyLLlrkZfZpn0FKLraSlYw01vkKAVOghWaEj5QgLJu74Wt8
dfGv6JXjAYnAcYocqgGsnnMm3vK+94FkDqRWzFxFpu7Ka57MjBCmEQ1CJ2LGc4VzD/R3ShRiBVrC
xxw6gNU2oy9cf9LpEcaYMVb7ZPwN1Lzf7djeYmyeftCvfArAScvFv0+lWAAPA0tJpQsWLa37dZHT
r0WX7DpjFDhjBIIfE8scb/KV3sHAB87JWR0HnNe2pgWE7J7X5BskfECS0OXdmODL1Ux8c1Ek2b3A
LDxXVJxA9uUVHiqfXgujSzSe/kGLcxwtJDHJIJ4DGA0X4cq+ltTf275LSmfdl6N9G59oVhJ5Nnrg
uW3upzF2fNCbZYczCmqpX7jE1BXYK9puH0uFJuPgPuSmf4uXLcFaUJGzQ2BRqfirkTg88huMv/Qt
Cu268G+44fVxHsrRzlqu2nuVsS8EbN/B4+d+qkcfTgufq3o0H8ub+ONnAFi3awfGdOKw6f7ozVg7
4dRttSktI4wo2WlxWsvODftaYl6uj9i8bd15ndBgT+nilBYZE5/epcicbjGTqBKtWRE6h8Robm4t
y5V9Z0N49FfQgxdD/dmyAXRJcxyzGrcTcC7oC7to+mX9sDnhAYLffHVSRad3PIJnV3NNdvQGZCu/
9iL7JeoHlTEZSi5upj8yyrdCM5aURJhVcWtPDpdv4DPuL7AEBaweAPzQ8p10L7qR9DxMzygkDyyy
cXBJJLkn2PCpso/VGyl5qyX14W3IzUHRybilBn85Th8NN/EK4GO0PWu7JEvnw90oIoDsEnzwfjtX
YRlVTiFuWKGzFsbRhW+/YNgdfvJmckowB3FZiSRVU1jhFilLicSKjAjcx7FRqqh7NHTBVNdrl61K
t4QL8pR7O3ZlrWa1PsmucccwM0kab2qX8WSvX7Tnqky4n+oKWyGALaZrDF3KmUECusJ3pOgI3MZa
LTWKIYdTE75helUiBn0C7fyZlC9aPF+V1JFs7SzvX7GzaydYbgSZroCw4XyrHt5UDPyfMca/RgWD
sT6lmQpLkPNwUtpjqtSQX4CjmrbwO2u5/BJFhALuJNt710LNs4CBfSCuHqkV+65NVBrCTfRkE2bX
1hLVdhsVnLi4cBCO4TxOUg0XSFYANFxbZhf5qxSyC/vMg9lhxUAqN6fq/C9wG87W4bnDoY1y/RQ2
6LkmpcIm5yF1pBYpHNSbc8Zz4Z88AhJPbdW4VxIr7BWGcucVN0yBc+C0ChWdDTr9d93QCtHWaOs7
YbvUyEGGDEHvaN86ry4GHcehZWMPZ5N3FFgmfZgWs2zj2tuJXyB39fmQVnp1bUXyiaNkFUutlDxD
RPczO7TZxRMSzv9ciEEruhGPuGJ5rBwz2e771h1dusFAKfRAlGrAIid0Na9o8OJeb4UVsZGeaKxU
xSUGrjrKbKfuIOhtn5Qv2XBucusphlckUfiJ5njAMG+kRbqlhFyl+vVzZnNzAewfE9Gguin2MvJ8
OP4L7S0eQeJwYZptuOeaSE9ALiOQRqHvFlCivBPO2YJu8pJ/tOqZ46nSE0LpSgsMAc4r5fZz2d6z
v5LSooXWynZniSP1cQS3wuhXqFFEmosvjmdjyPSrq47yuDS4bBuGJYcp/jxbPiBYyrFriGeQhO5i
eQzFAHhhOACyRODFiMX5LcrKvsWbU9bjDm0FyRMzi3eiVNyqbUwctSOvZNeixwNNeSSF+x5apIHM
/Q8s8cj34ogtk5OtsHxt58naKl3tzwnxprmMhEiSBJJw8n1EZ54xW/e2p7Dp7FCyIX33zQOOtznt
9gD0pNCuH++7kPiK9Thaj3GmIulTPHMslWT0kZPuWosqmYS3yNJiPhiqg9ryin43DLgggY2wzjPT
XhTx81trAj7zXwUFaSS8ak5cJ+2FmkLG4MT3qI7+zoc38ZWL7mxfoNYPFzZh82auFK8Pfe1CrOx8
I+W0YmKE4GuF0C85EnBYGNTLw7bliX25SjjXVgSgHKKhEsr8fKdpWeQQmFNqPV/xTm/FMxGIa8R5
N28195PEEYhbyFV35R3DeK/J0aT3LNtjulB1PIXhKy2IgACv3i0yJBalaKTuFT2Ew1t6eYgAcEyC
XjSnAGrSDN7QNbAa3d2T9CuASVogSRG1QBA1tC1ZfRNsXPldZ30GSbpEpIllWxGGsv/FVvYs0Gsh
GGdca+EHIQdp29amBJVQgMYhJdIeGqYNdJzfR9LRUCUqJggHC+FYkC07+DhGR+6kUEQAoX7ugO/K
pQfDHX63ZrcME9lqasJNJk28a/mdbiLa9F7BilZQqkSZGx2TwKjOFXWN0+ALV0ZoeWb5033Qsp0x
Kwer6V3RHEwHwtoYRRywc4Y9jMkBOueEPLlXWyQ0fEukRgb8gXIdxQ1QJRO5KsHfViQz5HAHx1TE
q/d2gDnKPzh2hHiJAADxXR9przV2KrS/Vwz2VC81NRkPySFd2HCFJAVo8sGBoHat+TumCxNW1cHB
cACJLP2wqXgXES7e7d1bqDB5+cOEdwYacSuC5QJEg2JcORvJfsgDO5o3pVMLycoVu9dutDwGXUHx
EUN4eE1g5X4A9omZVm5QH9HWohI+Gmp5C/g6EOpLCbFwujZUABtTcSn2W0yF2G2lS91zL0VvD4VD
lrQ4wZ3fd6bcHSfTlMRHVyviebMnISb95wJAkyns7EXDGX1wTD/WwdKDhHvPvN/w26vYz9TZlleW
G0MZlQwTIbMAipEsPZIIkebK+g5kydNyht4/nGu9QoYEsAYl014AxS3gbPUH0nSlXfKseuAc9GUy
VdfwWZMfBqq4W8xVCbvHUSqrHH5iAXWO58Kv2fqw4mXCi4umnB7HOgZBjyA+zpCSmFmOv+Mt1TtG
NGmdDJClDe+UC9YEhCUVHNigMJakynFduG7ZWWl4VH5hNYRdk6liwgJIPkfJ4TcHMOm5LLKSVgBU
3VXR5vtKgRddKhr4v0ACpQ3nk4wMxu28jXYD/PyTcS3RTFHZEK9auKc5x/yGKIFlO8AZCUZyBsBg
fzBqf0/AZetwOjUsTkJpwh+ca4swXBvxQOuSPBk8zK/7M7YJXFfvgKHOkqGhRqSmk+VoBZcTq/7G
bDUJMFK6b5gqLaBrS2fIWVV0aUVd3lALJ77B8O4QSrmsKMT8vUtqMIAuNjMWaN1KXteNz3SPwe1E
ecuK9ADR0zUeasrT4nVTsuDxMPNxwFfjCvdNXTGRng7AcUXaTwX2RngwjmzPfirzX2opjSXMeTQ4
XcgPtpJpt2FwOjfeYxIUJLJZUkeOdKANLR6LclaiIWrOytFN6On0nu483C9g6mjzxOAQkJvu9TQS
ZiD3NUVpKwNdVv/DHtNj27SniFmRiSk5U7Y8inewsr69z2S25JzQ7WN9oREdMEiKxRJ7RmuzS3Zu
vTB2kl3m0xWxns5IOtxxiAvQs+RTWT8b2oSDpv7yraaXE06FC1T3Ta+u+3EytLyqEYDayOToGzVT
PNGJIsnvhl5pq/UK+NJz5G/3zOoULdKliROrhPKGG5obQuJ4D7Pglsd4lK2Sv0IsdpxCjF4GCyDK
lK1YzKVz1S41WTm6sKmRBNGAL9euYope/n9KnQe/VK0LykAlOVH3s7mWarneB6A+BXzTNCqSs2Xh
30RJIm8vpkdzGF18IEyRa1j4fnrtbLqmvO8npSjNL3/pnsIe3bVOJqF+upmvYGKrE/zgsLJh9M/X
SWf8+YOUqP24nHNAyTSwe3F5R4EEcns52Y6cnkE5io79WcyuHmeUkXe11lIOggYnkT3+amBinNLU
dcgFIPZmJoRfsF/AxmLhynCYJIkYSxasW1xpfcdgJsagkIIhkVilzVvOX4a2GRpIZ4kMObRJZPR+
g5s/Yp+ueymomkWza1BviwjF68/s/4VxKGlY43j78G1Mv9bBnVZw3wg+CaNLOXQPj4su66HzD/hK
nbL+/e/Z847I80QqqoN+TW4GGXgoyEca+HiPuT0QWaZIWig/Olm6y1OF5m3L6L91fWIuoIG47GGq
/SciZW96nNDeyKedu3BWfhMJGz43/G+dEfAl4GEVT+CZUUy7pTquQGf4cDx0ZdFgmjdDqHeTW8I4
D0wYRcLluvfRUIRLTlYLshHQba/8z+6hsc+qHUcIYLEABhQ8CFancPW8z1Y7BBiLESEUYPU7BTvY
0gtWtYyVjunMqsekrSggHzVmAfiZoSpMh0BkREt4YX6OhR/H8QUsH5zWyp8T/b8ztYUqG3q5yHJO
3Xolq0/7kXwlQVRpfeI41/ExqlPGiPvDCHpp8KKZStu7/ibtyNm2zc0DjvOms2ZyJEkn7U+s0YHH
kpuy2bjrH8UOPvPeL9pd9MdeD0+Lhhg7VFmFiD+dKiTUL3bf5IiIx5ULYTiIzuKhLZkwsV7YDGIf
sXnzRVFZQ9W3Y+oYZUhb/b4g+EDfX6287NWqv++18z/gwhxXZrKrqZGOGhic4yulER/GKBEGcx5X
/mvsp5qAFEDgMhZS3oiFHS9HyiCzlh2pg2xE/kyziNH19ZzA39OxOhH72IjVK0C5YQAsiDioxTB6
tKBqKpkeEy+vOMWqnwlc7l4L506SNFK01j5TCXnywTdSfFACPFCQq/NGXokx8sLaNjy/UKp+m8mm
ab1qHwbBFM6nggFPzwZxhNQFlFpglvwRDyswNsSpvwfLPCkxdZRPt4lTWesWd8Kk9UqsOaPNQdxC
LM3Bw8QlaySsV67sVGfrhLF2fRxS78uB+DXzBRC9/AXo4vuzQ2INC2wnF9bb7yTIY1ALujb7x+Bm
H2SMw/XQPc/AW3DPVIdA9TVp3fJj6Xm0mqh9kG2ChYinfD+3qAqwsHfaxAH+gwbGIXFT2VB3X/qN
TYMOhQeHTspzpvusn6PKC/qnEYt1gqFxCU9SJZQnigQ9T8Ul2W/WY+ee6XbvrtgCv9LokEqLrcCv
iAAWioc3BNR16EkztfFZvdMEPrAJ3XrpnTYwPa+OFAwMCG60v5eZlkHn7I8UtadiXDorT96474Lw
NFRhKYl3tOpmjGW/Zn2DY5P85QtSsj2R6HKL/MbJFf1fYuicgnkvh0KURWLEtLrE+zb3TgKBN7RX
Z1opKewbwLlkfvRdEh4TyoUZCLzGgZ6lZ9R81CoNPNUMBjfHjmdXHBi8qs+xO7PjL73asBzDh+S3
eFfx8R4yRyvXQOyOAG3lUQhED6pOsZc5OaofBJZonTZGntEvhJK+lbKwal7XYy2L7DnwqxMdXMxV
jyXM+NP4kOERqQNhDFmPumSdPbVPeO3QpMUvYHc4eO1CgRZYRBm0hu/EzBW2FMVMV1/Crhyp9Nmd
JUTKd4B82NmtjlJUvyuLH/AT+tXSfEmTm3+rW3tJP0MX/zoP2niM+X8owFzaX6aXeV2nMMUUXyCQ
XMt29O7LZ96Azw0fKLvG5+pE62WnwYprMjz4QT359U/wsXMgtkIoum28NWStDf4SciCbcnHaJZ3h
HikpVMyQ6ATkIFrYWSYbLl7iwkuQ0n4wbJZrX7JZv55SvgUb4JvC+OVj3PE7D1PYqdsxPncWnbDS
xomUq8lTCeg5mZIaZn2TrFGtEO2QmejKR9C6Jjh7Q3+Fhx+F+oarptRxwgAgqoATsdaySqV/rPzS
FfbNc6/6HmlCSaAWQMvlL0GTq6R4SIAKllal/G4sPcgvtyOegjdJzjLtxCYq4C1ExvxJ7dSVSXYl
4x6KefKUm80zBjGvHPfWW48lKDlZhJopxg9WISrbn0rkBcDj2NmlBpb3Tfw4zHY0kG840AQEfzCe
tO5kLIXNfykR3YnWiVU/CBEgmPZP1nUnRVN8XzyT4opPt/YJxwRGSgMhPh3Fhx4bkYPwiXv40SDD
DwTIQkDIyazU8dNcKbYWZQfOwF3xpLoHhGwpHREuyxXAiqHg5jA/yFEwIgQ8m3emCNTlum5ehxHJ
FvyAoqC2coC52ua2UxdsbB1/SCJIe3P60K0TuQNAj2lxWa4MzgDgRVDvax3e2PXCAInzhSGvqTHQ
iF2u0RZ19T7d9GihnRPipyiBADTq/HaT1gd4JQTZev7Zsoxm+Ir9KFdNXrFDEZs1WAqttjS5mcbw
di43iryzh331NVrhaeddpx3P7dZjmfm8mVGSSo04xMjj+4x6kO0jgwOxiITVvYWfFc3CtJ+amSa6
r3ry6coNjCIg4pndHakgq0+nX8Q/m0clsycumHq9dcuv4I3AK/d1To1QtschE7qOAPFgd5eCAMmB
4f8iP3k657tkeNxBQQDkRfcB0jvs82+Ioxm4SPW9/s9B5p1N4VKk9zsc3XsCiUcUBKHEH6aCntKg
lvho4LA2aSe7Z4dB660P7QU9SAu/XLzy1QqahcI8G2q08tVfhmexyAtjof94o1vEIA2GkaNmJcZa
begwcBe/T5La82OTygBAA67YMNkHme9JemavQieZs5QIGA0tpy94v0zL5Q8J8VNJ9c5WmDlsTOQ4
OSWedGmoL4tHwvctFOSNBa0zt2UDrSSWEqhWz2GxiL6sEB3NvCfLKWVRk9TJ48ueNhDgWSttszl8
MVl6daSzvb+5LvP8rdxza+jR4K/Dak+0hr0M9KjIxVWU0HmJUGFjq1P+x2oQCWaGvbzoqkXib+pN
0UHRCkGF58WS3U3AghjpCpN7UT4Ha+GyqYQFfRS2zOuRgNHRnXKKqRhA/AKKXB8jhMjOsePY8Jsx
Bg7ZNWm7E32QawLsS4sTiy+6ofKx1vCXdnGr+bzaUThC+y6aDiLKPjzDJxI4e1yzeY2j22ryigSi
0m9B3BUwD+suYTBA8DF81mMz759NHlWVCnpTaivpYdFB8VFt2e1t4MobhO261ohl8hywtz4+CoT1
bpZAtDENqdzqHd6MgJ0QzPW5V1x1dH5q0IIe8seRkaC4W45zS7mYLsg+M6qZZiuFs60Lojk1WFqi
f5TfOEgdNzDHqUCYHVPA6mPkKmxyTUI40I36Kkt6lHG74Uzzz0plrs0cClQjODR8ngUG94OJXYM9
UrPgc+CC5ro2txSj3ZnAbSvQ5dpONKOZvSNfuDKsOYWrOJPik+/TgS1SWxqkh+fSsBAGTqV/8ggV
dvgLymO2gJbKPi7DyDOHy8Kvtw2h/0KFXFmPzT1Hdx9ZybEbCTGLji9OJACfiP60llINu9LLhRSB
cO+RaCuZpjNE8lcoJ8K772NlTDOfjfDtFeVsP04aLLikY0nfJ+NG8f/RSJGh9iD0l4lig8AqFmqL
dia3vq+OpgA2MmqZ4kkBHlTpRjPB10OKTD36us7rINqwsnUc8lVXWk7WOSeGR9IJxVlTQb75zDiu
BNMy0074Wag7d2yQnnO+eVS13Otz7Z0vlFcgTO0A4usxzjsVNgZ520gYL+6rx1ozfksmUtzmQsrX
OuO7ZJ+LQgXN9aTGXYcbD9IIXrnzi82Dez/ct+BA3kei+UKOWRfQq/K/YLGnfISqtNrVhNhc/yOK
ADfr82N7O506bPS/MyeWaZi/VNFTLo/FP7D3ezMitSypQAxmn9ZKf0PEoE06sDupFDOHI3mP4Aze
JVKUA4DTBxfbEOHAF8ZEpURNA/RzJ+jYPViyZlIYdoouVDsWIJYIDxxN62J02conwn15zxeGzjr7
wdcoHaWVR3oOvmW+2CmmGI9PJKxlzDowWk3u0HMLLfgrHyT3KrFb6erTOoYBwmsQx7sjfmomkccw
PbOICkrMYy9QUpgZBew753Vw3NZI5vlWNgaktJ4WRyeUItJFubXoDvNW7dmXEzHkiSJJeGwqIF6Q
1KejGumcVpoDIi3rJGOnp3ghzOb1EOSTzpbA/nPPYlAW/lUXHeQNeaonBgRmc4sxYJdfDppIpWcd
1jU+ZQNpvzemb4wVW+VfANXO0dqial7DntkJ+MikWAyp8ORLc1VeFHkpZ98VGQ5WVgWK7k50xEp/
QT9xmTXjuLQB8UWntaJJBUQXm7ia23s1t3ajIQsyAqWuqbHDmOyJRpo87+Ob4ZhZVDoyDiA5/nlC
Flb0HmIELGoGhf3bo/+qxTGlDceda6bZFzB3XAtSh9aANcD6MXxF524wrdDrWYNn5eLJO8LwOgoV
I91kVX5SV/R/UyeiCbCRW3JzwRCBA2fnp481qENab1cTvPANxW89xkUs95i9BIQXo0YsWD9QLr1G
QwQJK9d5U29aWLAD2BINhN/80ynHO8MH5zY9n57GXW2E932cWaYLcKP0vH0hEcrKIRcF3rQhCD3l
NVeANvBcMJWwLlJ2XSp7OkLex6N8FdCpDoZhRpnA2eyavdCmPKRGK/dm7Mb+R55yRdzW/8ybOdm7
TOEqCVqHo5Or4TqaKaJJOEidOFImXxar4MjTjSedl0SV6AeWzR4VbTui8vi+VkSxUSOOSPrjNl3n
PBre2aP+Ja9NLmvpVDomgKK6iskDEUWMFAVqFm1k91dzXik+8m9cNmFZpxye1423eINHBqsVFZPq
2jFrXzxJx9Tn1dbVm93eQSQQ2hOMNIhES9E7owwO3bZyaXAh4QqZQ7ND7axNYiQAWROL3SnSzyA1
E1/3LtBQ67ntV3Eh1UHP2XiBAx2fyoHCKoxdFkLfsIk32OrB2dCnk1LIOQz4pWzA4txtSL60/hof
mjZRXrAqud7OHTrCUiUelpTMHmDvCgKE/5y1xLuqryWX13BhbpPyhCY3PdEhMDZUlW462tJvduDD
M3SfYQSP+nZCKmsbHtZKZ91jmWsmTrTAlDQXjwALOTAFHRVZO4uHcf+KSHwgekhxXfQb+WNTG6QX
Ve1PG5mYMkEGi+FdoNVHWStjMH8+azlc6r6yVAl8RmIPUCHXyGLUPGqlhvbxEUxYUtzaYGbfUkKH
MI4O0LoBMSDjSN4KR92VFRW1yzdiFoFHCEjwj9odsNIO3D32PehHVzmWZnILHhzcIipRhVmYUzVi
99j0u/FchJA5PP8aOlWxMBhHw6w4FY7/JnCMeCMyVPbyrhqMDRaQglAoRrT5M4EdRTuavtYMHAX/
9m3FG/auCqi03CNF3v1mpZx6dJet7sD6TE5P2CIUHZs9wi7zQKBlOHPtvIVz9AGZqKH14E1rJfj/
Lz0er1OHfTvJEXU/JOtIqKH0DZgFK5HjQGt9Oj43pq3jIaemFtFDU5NbsQdVh+1HVFFQQh4szk0x
L77hwbDTTSGYwYWSw0g5IawR1rYgGhuI2rFwO/Y/Nd2ErjvGgJ7b5wHHnfSjLsDsYFJM4rYlplUS
Lx29pURglPSpD9+ExK2/CxwRxpHBr9mhwZUEGDdmyfmBfC3WHEkRFIN+d67WNxWv+0AtEXsqFaqR
FvDvbJ2O36JGmPCU3BFJOap80TE8DAtFRJqbTU/fhRoc7ai9QkbZkfauMokTYVk7dMq8Rz0X4L58
himMg/7p7sc+OLoXOrWEAmpA0K17iA+xQIRk3tHpJPyka+y5CyN4WGZqMzE3en25J8DyaV/l6EwS
bMUAyyPnHDHFvU0+fuowrGVAllXgnF3ILM9QPdirGZPlLE0MAiWJiYD96su5xKMXcfB1Yt27i5bz
afHRo1EPG64N3/mfiurvKlrVSc3T2QQ88UreMjLFl5teH88/W76WKoNz3DbDHd0C+rb9n44GdDC1
l/eI3QOn+mULWah9tE0tGUMdOJLOjKWzvYZ+75UHDgc+5JubWIjb6jttAQNUrmQaS02jFECNye7P
XLctlJBa4hFvD24W/7h8zfy/OmortgKurbKojsg1n9vkuTu/Bmuvk+9jEMwA9GrZkoLglOqGHYuN
vrsPKAJ2rcuYPEx/0Fd4tm+ZKMp7FyHmW6XO9FH8+rL2oOErdrOWTcx8fyCLVGl4ek+QMUjbeez+
n0fzoPh3lQ5q+sSWLzYQzKpXY9j0o4Ue8CCdQVvPFL/H9OicEu/XyYpMciR6lSJlQvpAeVmTqgr6
9GFhdtIhrRty/OMBMCnSBkP2zeo+RqJ2F0YwACDggHfRrops7t5FhSb+g4Tzm5qXmimkdtizelmH
m79v8BOWwVssniEo3O8+Tq/8AbT1uocMMyesEC7xpVtY/h4B/QtiTSxEuipt+d4oqx7DHJOcDO5g
j7972vQvchYLQmkWMvtIpV+IhfsdSbjl54Yx6lBcfpgReN1A5uo8QmxNwt8J0SO3b/+VCjgjbYxY
NJjItbgnE53nWWAcz+uUbhKiP+vANq4GUa2kQEPBIyTF9DtpXkTpHqYkvx4B4CibdeakKoCLuNqe
+vmy6CBZbzncA8h/uZpV4k1hHYMB8/gN4wkPIFbrgq3oKH+6rtBM4LA2BFkWTQ1dn/eoBufZnem7
MQ0OKd9RyYgJ1K4Gi/pDVVD3NmhUwnrw1gxUEEZO/cCsW6kAnEhPx1Hd0jJ/5MXdpqsr9yTM5/K3
oLSKyWTgTvhB//A/2YNvBs1YGZX0VBDducv2I41SPFXjOPtN/TUXPgHZZDqITK6vzlUYAIyZvAIe
N+7ySXF5ZOxixCzSDuXih2N4rni/3jPdalrUxV9+Zw1E3oLJV5jcO9hLdL/1qPx1Xra4IhSUm8Ly
J+iZqstAbfChqSkWRG1uyNKXLPBzFagTD7eFz8xUGA59omGLFY8TDeStq3R1rFKJYwW9OPdmHnGI
I1Lve4madlF79qKW4O0DZHLlP33Bdv25ZN2jc6vsiX7lHNpMrOxyykbjpq7wlMvkr9Azp+uu2HSr
YFxKzm5Vifk9sQmA0SnK/GLwTTqrfOFQTnTvYZM4pFQO06/xuXNs0oZULmdBDUmHZwPr0jCXkSiz
cmAg+mzktyWRl4Wt7NKgBd4ZsVJcqEQhRhdGy1y4FzVPS81A/GUADDSIMW3zB2rzb0pyGAN75EZy
S8Iw25VhYDz1lYqjQD005dVFtnMn3ov7wQXR3Diwabm+LdZFDJmBQJhlbGqpuwmqh2Kd17nYHo3X
pRbR9UryNLQvHbuVpfRB62JGNb8RdmrIYUaNzGBEd3ljwoeJsRU1GjDFrfOZ9+vT5wzI9VEOi9Rr
Y8UUOyG8PGIvLAAf4mosoNgmDjjhoFi90/IOMO6SoH5UYZJhP53Ue1P1Fnf4lHc+OdIeFze0dKwA
HkHZBsE9A3f4LcD2n7Tm9zcq3L8tjvh/qJhff3B0rYR+8AiYryHo0cGCIU4UQCxv0XwbtCPgVk4g
ynnGQf6G+/aHZYKW7eG1EAMuPCf75Hc8u/tv9fVH6aQuyMhzjjakG4a6TtGQgGY8iKQedjNh41aj
bFJS2s2yx9XF4/MtZpdevbucpr0/AY5pAbqUzQ9UEUf97uNhtXmGHcj6aUQzsTZiAaElXo47ORZI
kZj6+GRkpNsRbud49axxzcudS27dnqyqF8xxT0OXvD/o90pkU7WbzTxfZa5AN3HIfaBmxxW2JJ6j
Q+9+3+eLsuq3ZRKOvVO9Bs5SW67TD/ZhezqQsQEsWMv9ZLsnNFnfiuggTOWINgnt4cw8EeFZctXC
fiBJDij4w7/Qu0olK+YnNlo2MdulyUXIQznTXu3KFRtsL+23kEEIYyjML0CwuPs7IhYpsju5Bemg
V3H/T1jayw9IJqPbpgCiZxsE0fPbHFKVQGjJDMve9MbhgoDR5UOL21ybRRSrnsshaT420sO+q4B6
ieclu4K1UmD57szzMFjsKp9uyFCDhyigQyNaqZF3B4bFHhPwzd4Eaix6RV969gDwhdYMfOegJAVq
SkeVCoysM3t4+r2HTNW4MwbZ5OXmRKctyUPtYdhJG0M5tzm5GTvV0okhThmN3B0FDZSL0HVZWdME
/dWb/fl6uG067ZZOSlhkMghgEc2b2ytFstGQpvzT/JQR39Ig/HhxcRlPsb2RfHLTvaHNQfRESQhK
hvz6y7c94lFMqTWmjw/C26oTSE+y0+zqnslVBmaYm68NcpgPU5KpNdcHbZgUFglf5beypLfTLIbG
KC0YClu7IDcBHnGex4UdFAwWHEx9yvUgyxVwpnwPuP5cXdkEYBcWQ7NXXKUk6sFXWNAlmlb0zJL8
23bI+OdKaUvuaF2hXDZowCagLyltO7nwWtcWHkwonttKLvWC6FPRIZfPttZxyKxG2obiyg9AnfYg
OrrRx5CgX+FQJmfrTy744Q4BN52Ju4fmbLKp3ve4aU45eaEpzCaYRjnCI6wedygXEshL1Duo7Wdb
7SX4X/JIA+5YUW1DZnD/k0W4EyAiKLuC5tVFDmHI+IclVyVuGk0Xb7BED1ApNguazI+4eXKTE1jB
pi9gRN0jrYSTN0cZUSkO8hX6fxKuhzuqTe687RAO08RUyzG3fFgUyYiEa7zs3lesvXoSMgO5JmR0
nDlt4iTeX1HJ5BDBw3XJcOLbicsA98gTDs0BQw76Q1P2iFNmK8TQqXbvUHAfJDWbHI7YGNdV7n/Q
M+hiXCN9o0o+HQQ1LYEQg3QsGv+lgGWlgC+oU+QXpjcm8wNjZK766t9tvhx9oQPgyqzryWA2vn6a
MHulBGHVliJHtl3svATo9KO4IurnCn2IKOIycDCyI20O9aJJ6TJJmbXAv+v7wqy1hFwnryhBYjcJ
ZvFlLOPFC9ak0G7N2xQELpUIveOhz+Z5a2R+VSq425D1sQO2ZaEM27+alnROJMcJU9fUEFCsQ+BF
PoowFX48Ab0n1Yi2vkbsQlM020PPYP9+WGjLsTcALngusUo+HiD1Od5qdpwh+mSu5HrDocafHPeA
dIsez3Xy3jeFwiN/go4YPRjx/qVRC1dIbFsU+wpxrUqDP7lJ1uz7gAzIgomC++zxDw9skpL6GbMv
NCKa/r7aZBd4sREm53juaMUb+qFtTWp+hJmQgzVGQkVMimtcJrwdcqYfxd87TblqlJgUWBXK0qkj
AiDbjSzLIuaRuwLVTX6oH/Qix+yTVixwB8+P5qOF57LHWphhqKNcqW4Q3Vly58W/yryM1CiLg+JE
L/NBs7pl8kSxp2nRuYmNlIKAJeMMIXWBv9Ipk/HXf04yccpb6mkva9vxy6rCFvEvhORXPfrtIEFs
cVfUx+Z1O4/CmdHdlpTwdxHRNClgb6h6S/Yvt0j70CXIz5gQ0G5qpF+WsdTxIVWcNjsmJqecV9+2
u7jexiapMgQPbQdJt9bwYhPfyzMs2KpPXdh6lECyYw3BX4biOTO0Zt8431OavN+x+8Pi5HIEFixI
ub/NFmaRbH4eXhNwjPVZn789BaRUVvgwSz6fDPKdqPHuoZzM7N+KUcx9y4M7F5ejrtUVwcBlePDY
4r3RSSr1hUqWUK2WvRxAP/tFKoY1DfRE+ElKv6zSPA7ncSkV7RvElU3LfrXv9bt66RWT8GMSC1d6
IuZuQzS0NDWk2IhnsFzdo+plty97QDZFSsh9+4tobHB5jQKZC42vjL+n+qFbBjvbw17uBDLn+Lr7
0R+B30FAfrKSvY2ZhqoulDQ2CiAPG/rh2aGV3mAArCY7fS7EsIaD3RbGbcRbrsi2ZtsIuFT4/hjI
vzIoZJ+M/WdUZB+uAt3meh4uGY1kG9QpcChMfps5SVFK0s0flFUD4xUReSlLiDIoUAAFrU1oGMbB
/znlRYOJq3Ag5nq+jq2ftviFq9H1eQ3J39Dq98DOY61aWEHL6ElJy8umPDfV3M95xZRUnMQOKzCZ
5pisdTxZQDi7VRsA2ZaLAC8poz/J7U8oPGTuo43QngmKEzNxOFxF5Ux024JfIsdFt5Hvpve19ypb
ASplR1f++ox7hsF+A42dxsMeCy4lCWm0KZPMio5mrSpQiUChau5YtmDlMnm/KHJsZsFV9P521af6
1wuqZDabZpRiM3oHVnDUfRTkt2QbG2LUY5iNJht24GHtzJgx2DXAU3kiPF2oEQUrSvuNsV8Xum3o
RPJ4e7QDY4UJXxreTq/UoZxYyW2Xju1msp1msaiSDYskP9PkQmxzWNU+biQdASt3Lkrc9DJETp5G
xA2TeB79tkM25rjuuyKH7D9hGwnUMn1Oirse8ufAvUhINz6A0vn25VVWFMM9sjtX173tW+P1lRNy
5M3n3hf05T+nRp/aVhsPkYv6MZpQ0D6UULWupn+RXacQC31Orurzvi12huAR386JPMvSB/4AhW7/
FLl4Rab5IFYrgFqF5DuAOurz1nwIVxIUPIzEBBEEYrrgvZCp1hlNex9A5J2Hrvr4K18I5Ssj1JtG
z75CJWNNwpZWoycdC3yek0SWKX71R3IHUPUDVFOAgJPnly+/WbEmnZLyt8ra+WKSjclfwKOpJbyM
DqjJWtvzEondP8YkxxJR2h8PTJmEUEPEs0tAsjvkUbfXv8FsQbqlL/M1PSXTz6pTqwqkELAuFof7
s6K1/MMGVJafB71cCqo2YENzV7K/JtvGbiuEAk9zZbQdY2R+SpqDnCpI6MYZ33bkZROoiJLcn3Fm
KcnB70pjU6GC2CMDhxyIYWcrryRwbufoW+JHQasZBjvZ/Nt8lIg8ckG4p1Ru2q0GQ2P+cwxvwEvw
MVN5vXCnX2v0GHSfgXbkPOHB4Vnc2Y8go1cjmowpvkSG2ONgWIrQmnQWGTFK4+NIAs+YwmTtzpx/
y/ixV77VTpdW9Qi8HSziS0hCnmJFOHt9+ytgWb/N33v+iuGuVwT37i2khCtIJyl9mqlfQvLCcvgj
duwGp7L/SEq5IgU0sBwf948mKf+z+t7V2JGjG8kEnWHmd1J2HHVzwhkge7nqZ9BlYmSUlT5kVx6X
6/pPb6u5rax943fMqpFf9PY61OecdYXQEanOERKJjdqkINl2VksZgoNl2pNf70ehvYIaDmZ30cmJ
QiDblh2/mSWJo+v7tISTNdLKO5Dqw/QUYAuCthxxxT0+IgwmytuBqQ0wn30Xra16Q2hDRzCkyM/H
IWWCz0fNvBAYU4koRFQ2jzyEzJrbi6Qr3Pd/yJqStykIQoPu4Z/hJUviXobN6zvR7YeMw4wpGGb5
c7NVxcE5zqXMGvBjb4oEbGwID9YaTt5o3FepzyMPPCNbDvgTUMfKu+2NB/CaN3HYyS+4GK8cCB8g
WcuLKLE442VgYBj5slkbya5QKev1Y/GxbTeYYDNE+++tBEDwoXXQAsd1J6tZVtXlDK5GheIsyrRs
yn1Ng3TbtTlZt7SLGAsc8e2w7fLnL3Jc7EZ3hO4vCImCHUqG6yqLqSzvb8qGKhl+XQjfjclYx/s2
HdDjTh9ehlwC5hXfRrQLBSSMBTBmk8jqHnVmqN7WeRKGUyx1tSUHEBL+2sYs8UD14eEoFwzP+1Kr
pH7d43ukvoxUIxX3C2byBbezpjDRsRdmbIFViVG7epHLarOAF6ptp+w/CsdkHYQ8QVgEkYhz7GNe
BYzU8q5nmL1VEGoBDHHf1CoGKIWrOX3CpaZzsE0mF0pTDSQNmiLlmCC2QfmAjR4e9ZrbSmUjdVvG
7gGf3Qnn3V5ve+zmLzXqlJINylo6u7dPFK4207syBNfWwh20/8MUg1wkkgrXruBG6NnwvYsXComR
u6cpMFCXHghC7dhqLQSmv/0LrvtUan8sSZK6OtlftD8PHibr+YIl9F2OBKcEpSqYYphueP2LEzhG
JE5T+CKCPVCTWavpNoGrpEdTrZYUYeNWRIfBlPl1tyI5XFIllVhwZ1AW1KgjBrbIncstZuvRQRaE
Ct55Vf6ezXQns434kyeWKtRHml/dOFhhKd7RdOCmaqlaZLHn6GgPu33lPh5mD4sJThxlC51ZDS4A
7ozxX10Krf37YIZKEhNHfyNglPP5tSQLWAkUvTBpkMOEy2a4ovOoxT1Qr3Bv6LdWn/ZaLupttfk2
fFkKcU3dkg+GnkC1z0YSjRzgfHTaEK3vyMn97/ZPUfm0tSj0vV9eruWmx1KRMwiJvAMFjcWMN5pl
ilkHreFc0L09VBgSszi5BoFhnPIicahUp4lYIknbGNBLKFzeFosF0c0Mz/Hw29VEko12takjm25t
moauvCQfME3VFy2rCZtSEvRzaUlUcT6SRmzfSGP6+S7kdOz8vYEYXG7Oul66exSAsiE9SWqTR0Id
gNgElQEYxNUv8AywxpEzWptooKZPuitw71MyOtK88hQYUjvy4/HETM5tCOP1UNowsrdKnXVQAn5s
tw8Mla3nle9IawszNpUCtQAI8g6PmWogHXNUjfePtS6sqn9gm1Ly5hYoMBn76sYIHByvNxAufo7n
Ky9hc6tBF5Rdwbn3xZ6OUsUEZsXVdC9D044yYwGmYHL/B47cQOMLtgIUz5XwnMxef58ACgXME9g3
3MuDxKys5gDp0E9O252QxXk7wPydg1FfXtNZxwLcjtXf729UdIOjqREdxSfb4F+gMx6RFdtTA2z3
sKJLtNqOFh2spZQ76QQtgTkineZSHhWKWMlWDhZn7blwZuy6yDYlQRciOyzeXFAHsFGUoA0DG3yQ
oMUTGNiM64yf5oD+h2vwX4GyBNSJXj7ngtkjK7sBxCOE0nd+4msyq4SsjjloQ/dnUgCytLJQQ8Z5
yf2pzbB08BGinxLmZQKANu9jBwdSB+mPm01e6eGHvRTuqoHSu/xV90YO+/5WMnKkfwnFKSuHpBVs
+Eb3k3aC1dgJpz83w46whVxXflYT6s4wWJZvL+kF24u6uLDMXAzAp9TZKKfBXxOmQvQXiZCPhapO
HMuowArtOp4Pi85do/wZd0/49MWvWePvmkzPGTgtuDybCRLHwkxsuWHRUYgWy3sdKE5o3UmW88ro
wo/g0BD/iSI8jCFpwDBK/vJ4A1m7dRh09/5lW6ynA5spWhj22dvTNHF1kqOH0SetefuM7+pmhA6K
6XyrGnueAel0u9e4gxHJ/K4oOtVnRVRTih9g8kp7HZhPBuxLYKfQ/ItjOLDhJgWBuIcTqsfoG3Ec
xhxR9NMHUjq8PqXPMK9KAkDtxNtO5OSb95RCKQdJ1aoH9puue+ytDa8V8Z8Ru6E9IHcO3d3AXIMH
HhL1RmVNBVWRFaetIH2Jv49BaYtu82BU8+W46EeVL8qJltVKuX9PF09qOqipXfwYJUrZnck6MQqZ
jvfSjH1vwMnecnSue1X3hPKgq/+FXdDjn0ngEaXees0ki6FUbjVlMXNm2YMMsVGjI1rGgLC4lM63
KhOAzvrbPUOiqxpLAzx6GkQ5ubw5NnPw70tCEtjQw5uOIIyfrEG2JNAm6jbTN4Cqum9LDb/64hZh
T9ojZdPv30nhheUKaamxkHYv9zGwr2Kq8JBLeTZeFJ1OD613nGux/4z5/YZzP2BO673qXxZ+EZC7
c+E59si8L/C7BU4DSmbIXBhttZUloGmuyoqPlq+3QKu1of35xKsYd3HSqXxXU3pCHEqQAwRrDlPm
C+lDnjJtq3HAfngOjFubunXPi4GKqEuQcLFDfdqpjDaG1dX6rhGGs+vGiVQUxJCmhbWZpblyfedd
0Ch70gC5kXGiHD7muDNfu/C4Qx9sLY3LJd90MUDjQF8LbeJ/EwZ6rP8botqBJ7jS0kvKu1fiBPz2
TL2DKfkolUksxaft22N2phg/SMLVpq5cIPozlqMYFaVekRWd7mmvadeSScsSh9eWEU6RmS9Lmeo0
OtJw/D7IOkcQoeNwrhHwgBaEjEvPZ4CV2TQytlJlbH46QxIZkUEuUUHESVF0/n4107bHkEcMugsV
uUZAeulQXlA3YGJlZLwB6aKA1VbWJHGPJv9nicxYSuIEM7UwwKi7FchWn2bQoB7LYoVQ8SVre4Ih
yY/F3EcxtlleqlikCpomGOUz8BbSNA1PDjBiBsQj3dUtM8MfzAnE92sOCWEJc6dbvE6eIy9o3uK4
ZHND/W1WcU8EJiG+7bwwYHutEs/KxJyaiMgy6xQ/44Y7OwKlDy7VHVXMg54W2qquhKLHb5OON8QU
7m+iJajB5QkCExOV+IMnY69j9QGb80OJOVnxd/mbeFBM06vXjT5KypIkA7Y9mokWxqsdcfmB826r
j7TPiYM7sRysGfHSGWkEbhf2HlAdqa9g14OIjup8KwOU2LS8er8EreqQt4CcwDv3ybMWLk8jgPR3
Nq0Cq9B1Z1wlOVcg38ZK0nZRQpj0GJwulM/l3e8vNPbrx9x5lV5CHiiUlBtH+RlIb2KxcMhKDkih
Vi4alfd9bSOEYNUmE/3GTQgRMGf+xxM+mgK9NcgEMK8ygAPJ+n9eLL4GOdvQ96m46YmuZ8kl7etD
z2BhWaAi/yUDDJ2p19t9nIgjMgDV7ljqSnSB2a/x0oLndEUwv0wcM1nhu4FMLd7JIaRkGnYVCmIP
jRiTzaMnPiOLGw7/kMzbpCI0rsiDFlk7nIa8F8Uit3Ks9qfrNBeiRmP/rgJh+Nee2LVUpzQzJa1J
XmKPmmkbuQ9jwpS/qqzDlDGa5txlM0OBAQnFp8NHC106MgceI8An3sWWWPOzSk849Vd60EUSWJ0S
b3q0XmsW7r+IJBE19r+6tlrT5yBFGLJVIfJ5kzJ6t5cvD3WzHyQKGYuq7I+CI114+jmInisprljR
jbE0d6cL8a+oIFJZaWnbIiMSvPDrxxLusKRvyFYiOttxdta2DARSDcj3UkejwHYjFhk4uQyA7Pwa
muQAST58QhaDBzMuPWYZIqso0YCKAbyZdaWonM7OHxNcXmwPHNzmzM8oIolQE5IYGFgMLgaD4+G+
oOOadnENg4VPw7RkKgNfzlI3sxAVr0MvrRkl20kHIaYrGbgVJQ+cY1UFSKoqLMJEy9VNhTnUjcZ6
qEhZ+kAVfHuDhNz8zsxbVw0KJV5hAler1g0QdM5V0hQrsd9r2/4hXHN7FQ9FN54rsVmSvcCZpiam
1U4VH24u7NA2SUzVKnMcLge/p7EvLsY095/kD96KLPXxqT8+FwAtXVn6CamPhb8oqPlDlsgbYroZ
bGcd8iNgXz1jioU+LHtnOng0uurYU3BXQOyaCswkcAOJjKVba0wYiNYmvASAu7UwGNmAtGWz5lCI
717D2NyDLptOBvcnhGCxUfVexj+Tpz0LhDxDyBDAl3eZYyiCF7j7Xt1IXD63Eb3ve7+RREaEAB/h
9j8opvaHPfxCa7jKhG/lbT0wiQUKzjb+TPThLUzYr82OWYp20HClXrOD8DW5KPGDFckEj5gaT80q
g22FLd6eDkzejTakvCU4Fp1ILkNhL1wLtGrCGjgkUIWvPPPpBJRW66Yv1ugxzySuLR7FYlcbHUk/
6TE6FNE122iGzlP37w3EakT+ujBKmKa2gW+PlmVaRhJqAr1wXObRqnXJ3g4vUBayZXNt1XaVGs7c
I9Pque2UpdfpQeb+mzA42Nzr2soZv1ByMarx9EQhsssJ0L7c38LSzIbz8zP0Z5SQlBIupxybBTkp
JoEkbX0RjF6icT2WH0KAgP1kKrr7TIqn9yJIWYWtgpX4lwMZmm10mLIW/SIuPNXTASjQOLebKaLC
J30qt1JLvPlUGUsxOW5a4C677hQcMiwE9B8QfWJgIzVRc///wWmogQTpZvY+wtpjl1ZrtnQK5fFZ
47xU7Ahxr3OWW8roFAD8Gb7RSjBP63gLdbGDwQ6E/aDcpTpmo7CxmixbWQrDgKkPjp/wwPuE4T8z
qH7Am1CEPJpE3/05CMwIyFLqbHrLXbW/dtEMoopGd+sNPBAp20J+qtZV2JDDesAB6cSBOHiXrgUy
Bof2zHIgsKa9ssdNZ8JJtTtOTLgKQUFOZzWIGXcJu1E0aiauXyNF0NMEzBX9OYVc8tfo/XDlRy2K
UxEXHD5OOQ0fztWa3nQ3vkUFqG2bedPduJmaVdMTe7VGvWx5xRbWEUd8rTkUIZQgAE2qdfgYGKGS
IzC0MZD5aBqEWduYSosQnPL5a83so5W34IzmBCDhpu3JBZrt4QU1U2PjjbKehi/BhcEts8KKiCZL
onwvhwEcbLRqKCH6n7EQjunsxqpqXaKvMoX4Qrsld6Qu61Y1dlMjIglWhBHFr1UFgEXjf3+qfH2C
92j6IyC7+PhDsvlUYJtaN9rbYpbxC7WroaDVkzQzQgDW5gMFEEOB4xKd/qBragsdDZ5ScarHGdmQ
C0bRoX9o41pguFdV+Wc6oPFzJtNBW2Ep7Jv2AmVmOAa7EcH8cbjkwV0L8+WHeoldopSns5+D2Fv2
8OCFekApc1Sn4GN3v1I8vbfSkfKRJ3bHemNPz8uYjLN7tbpdB/b5ATRo3VWTXKZ4KFde7YmxqJqd
I63n/+8KEOSQMOuUoT8NVb4tJs+nFIasa13hP/pfE+0FE01P0BFyqKKZOZH4sLISK1adi8bxAg0E
RNbYROofS/L7a//InhEqUs5bCx8KBXfJl1jJQkjBan8DWmBv69o2X/xBY/oes5yjnKAxDGgaop6G
CSM3mj5NnV1nJ+5sDBbRZYKcKdAonemhol4WYgcgbHeC9Rl5Lrd/nnYr7tPrd8PtTbKoRbX1tcBi
4+0ddxiHT7sg2KhVCV0RfaGRdoDRy9Mvar1CFW1pn/KuG9blQ2q6Kmzy2r/ooYLfDf6qMGNo+NTq
GEQLcZBY3DQztPQHi+d9sZ+bLTogJzzQAJ6mgOSQCe39UD9M7+/n+WlEY+7bD2h2Rpo6y8BK3ekZ
b80fIayBhWaDjeIgifjsB+8Hi/slHDnfMo4ZsuEKJj/KNoNl9szebr+E1o7942XabauWhD5m4kkk
tYRzaUX2dIzWO/lLboyUzpmnYcpQrDm6E1P0LIJU+qOzL8EeR70h2Tvo/yy+LsybI3P7hEwQuYPh
Y+cflequQGKzIK8F1VkMepaNDY7KWXeiXqVQv9pFB9CtEZTYbfd7UKvuKFGq4OlNCT0V9kU3iQYk
RQzUg+39eQIWxXZNN92yJl+qqYk5JOOL9Bc5elupyHVUyj4mMz4j0u+4oQO7BJyJBQl+4+hTVs+s
VQCOB0zUsVopEi62eFa+v4A+4Ru3bRXUtHzrdC8idTVubrJfX/rQF8hqP8OPCW0c3VmINR1tbG7p
ckcpaqYnv8OUd6KxQrL25ycyMGEVi5FBYzhYH34pPzPpR2oaJLLDILh8kQhOWYzgDeXD/afXSh5Y
sfipeBOAnGtkulfR5XxLLTSTYTdZ5F35672xzNz0lNB2tSWZB9dersLmVU0stgAvkXi6ot4u3qAH
03GWHVC+0U6VAdzkp1CrHZYFDqhao0Rkz/iCuPGTHVGMwRmqnzbiS1FXguvsUso30ziEsf6oYiVT
MDrOtMDUkHHklwtddbHoM3hj26ZGWGf4o6ucKAh+ulqGE4Ajve/lLTjYiDeAf2Jcv7b560WHuvlh
KiVsfwiAThFsWC8g6gcIk8/lvodzEalS2pFZfTnOEOhqkFMvfUk5p9k3HpQmVCrkOKhZSMqxZsES
yaw71bnlcQ62UG1ou0GR2hFeJt0Z+WNcI3e0vYFmRWJNaKyHB5zGCV8gctNkYyz4oBAV0yKPN68A
Iil/NpkCd3KRlrCX6HbWTIsL6oIJS+ViaLbIqNAGm+P/Ok4U4OflvAa5Ouzmav8OguZrvfT/nO+U
OoesLJY/9G2xRx84+H1YzuKT8hGiwpOQVEH65CP+RMrVdqcszplnKbujG17Gy5elINkKkW1xK5Ij
3Rp/F1MhRidKyFTiEuN3xX+lW6Jf8MIkZdxKStgpoUamPqXWCsAdro5rWTdDLF/Sd+QKCorvZPnA
KnQTABOdm4+BvlDmdvs2s0rr4WBMohKu55PXekF64XKTqoyyzboXd6hqjevjxRU7DiZQ1M84YGQ9
nW7fTDbKnypqYCtHH6uOG8GTIsdWeBR4uwhR5IAF8mWbY1UUm22zSmSqEi8rqYvOSuw3jGDV4axl
dqXVQ3ybhvs1u1J3D6ypr7ioLXZrhE/pHgJL/9scWRcph9KR/19wwpT2bNOGhDxWgYZtqtHlBme4
Uk58Vii++FkiX4VctxfJxxq92QU5qRP6C8ggNfGwLXZJnkMj0k40MVzbdzIKGbYRyFmX6D+FFim1
vnLt5UrH2CkPcqSEq2Pfwc4eZ5TUaXOqPiyXkXCCIlDVu8G/cTn9zVroA8GYbSxH9NJc4FRiLCHG
gw4TEKO0HTq5R9Vwm9EdFrfPnycFD1ZpepvPz3/cAfmuqMK8pObbEa2GO0zGjjJ7QTBAiuor3Yyg
lgbYiZq4kULV+MS4vSombMZB7RgTHjFxNNGpBJYe9zhXTHqwp9qHDHotAWKfuPpJOrx5WvYZPrrQ
8yne0irivsZow648kPJ3FuS+lTf+Oj2BI620ezo2x3ky9txO2VN+4xGg/HSoxQGDGKX2xH53Ooy5
ctjwviAQ+xG+l274ks3VF5DczLHihtT7gurveRhgPRzubjGqFC5GuLRbV4NfeVkqpkMfWkVkCGwX
E0co8vC4zaA1DJk98+Vrk0WsOutvu0yKkXERhFvQ7XeeOj309+xmWtFVKc0WSvPcjUTYTsdUnQ8N
gCECBIFtTk0PMsNnKyvbMr158UNyDWj6KpeXN4SQwS7bC4gOdGm+ASavGX0KECY6gGZz3RDJ90XF
j+ppsEl14Jv6IR3Jwa79U3xDlprz/5wN8gVJKHqkSO7DsrPDAePo53DpmhZCLWj0gBGULMP5NWSJ
UE50IIg3q0M1ygSNl1nbW0okpc4O8vWF5Ac1+alZ0l9f66ElZLmwKl0eyQzifsnSzzraMsyzvGT3
OXcBTcLgFIjLKaZghtU+JKLIOrSJhd6TSKui7ycl4H/zNrhYZzKqtXrXgLEJ7r8YoltRuJHg7Lhb
MxBxf/CD58RB6IMUkug+qBdSuOJaYbHx1IK20bgm3ELwLdbSTPNkynWqD1iK6H2/57SQjOqJ7PgE
pJ51h6ljROeiTeNuK1v5Shwq73Hruwf3GcvsjkLKtcAu6PuKOxIKPrasAvamZMUdPT+RAScbLe2C
BmVMFbEqWVZX8bJit8NPoZ0biMzsU5MNZILPH/xwHfKexUHh/lFVjE88ENkV2zY/Fj4WmSPetN5Y
mArsRbv8JkVDZGZynToYCgljIQOrRb7cw/NbsyFMEp2BaBS2W6BYfAnSi+JvaRqn1bRzPOrw943g
B/+oPgB9+/O+u4vWrD7riYrr3iC2UHTrh7T5d55BxldkjTE544zXByZviwDMp7OICXXnZg13hPRU
qtiFifjxdGoC88G+ii6cb4s1aJ2/kWjbDD+w1ZC6ZU2c8BAslBE6JKvh3plL+/oDW9I4X1hyT39m
+CncBwBLv4TFxqDln5z8MxOy+LKtLedJfHXGQFD2GRmti0aNMxqywWBKC0oH1g3Cz7OY/pFhaUb5
zKzkwOfsoiYwmDEkQqIUgBx3Zl35/XIpMzYOM7uyaRgJn2EYZZPsjNYqnr9Gui/kvbSDJymVZ08a
+uZkjTBngTRC2jpK8itQbp00qGTowZyPYc0n0jdvYCi9SBRjf8p5qNy9HVYq6vAszyhn9lzBuTjR
kaIl816cSj1lcoqaHYAUZY6CtPgvElS3AA3pg70gIl6uemtpXznVHqJdmAClUln4v6WM68bJgzBf
4TB1WY+ZGrh2wxXd+I0kghN+m7Pyw1CI5iBAvMPLQfxt9m1k2BBSxYt0D2b74iAfHNmugkh+ffKp
yNAbw1raycJbnOyNfBei/Hseh6wtNAK+JrLEbD/579XSPzLUzma+w0LH80aYdW/1GIRKahEhBQBi
9oFBE7K71cfkA0UDOqafjfgpdIDx1GL8M+n9dZaRBmIKwcwqApBTQTMlx4c1kYweekpqubzz/wVk
hiC95X6TsfGS9nQ1hYH1LTPhWgfbGWXLkRV9BZGW6XMjNRmIyKBHLb7mcGAcZ92W0q3txBaHHlI4
N6R0UxZpfpxNvojxJiZukhInaTlFbjyL6dCZT3XvCYB87ImWYrYSb7lnYKkoHwqq8SDEihZDKqcl
6tEtr0XdoN/D4QUf/DgROe5b8DasvmaGKC3GW91HHw6nOm7p6yNagIbnDxHXwSGMfBTkSBn7pvTJ
Mc57hCQKW4fTHBdby3t3CArizniHutSgdFxRHjNGo9SYPiaK967tW2+3QUtiq+nA9kubEP+dkSQy
V7cJvPtmfoejtDX9ekBpVOyJkPzBoAtVqF0iU2mZLxufhkUm9IrQlEdZrMGALVQVRPk/qpiHlmkL
t7EY87DXcZcg+vEJiIJbcfuKwzV05QVTguMFkCezMiycisCxFBvnl0gIdiDzJHwBYDoDRLbuKRMY
zCuWNd87bwB7MJsq9DDz3ExtAXztrATwolW9lDSeTFv06TkjpYkj+TemKRFSK/Kjfkfnh2ug87Uu
tOyN3jM0/wPc0ZPt2m60T1v9vq7poxOjmC4H8FfSOjrwAVp86zGV49Y1zU9pOr295UpZp7QsYTgJ
XnXlgwKmFUriZ0+CmMI47aitlahkJeyT4G3zhwOL+H4zeBm7zA/ew4SF17LmwTDYtWlZ789H07f6
tCO4di8nNKq1gc+zKbMfwuUaLAeLQ1flIpFN0ILF4hD77C2brG7QrPz1LsY1SvdFUroYXyF6DizO
Qt2gkJMfEGMwBHNKxDHAuuL6pztKe5Q7WR2c3DRB55rIWJI645YFQf1Kde5OTXCUlwaXkZl+SskF
Rb8Apk0YK2gT4EEc/mSN/v48ZPz2tW/rhdZf52+hruhKPPtU60YgsmqXdT185+vOuLBaR8DRIhCD
ER5rNSvGZFim3ZvFburZ2F/nbXu8eSuDKgnvDNhCwT0FkQ0/aPlGSxdzkNNjV5UFKRmqXnPhIUXZ
5ZbjYfDF2B7IVokrxY62cz5R2AqNqjmrg/wCBs2s7fd9Iq6l1kewwcDJjZmkpUTarPrQyptP8d6H
Uv1SDNH8PrbQir7WMJZlUtwboMQWNaGgmIQDE76cTuuZJ2Uazq7VhprnRf7mUFndK9w/Zmga5Pbk
q95LaW27mwJA6eVNY0pjSfxFm18wBoMEnUWY/0Bf72VI+Zb8rgmPSj7NulPQGwkZmL6yka+nXmWD
XyxqLYvmxOIqI93Tj3gk11VCHO0v2oztXPi4PhDYfuNJRkV9heeTKGkTpuAQEu0XkRXpeo5YjFbJ
LVUs7GKKjOOWS4hE79Apxh8YmBThoXLcc1s+FfdB+7izm18EXSZYopVTE8ugw5bnC3kbRSI6UY1A
OVHjVt+H7e0UAiV3SpPUDDI8A8l94TmowUwRB56ZcqTwjxfdQSB/Ss0ggNxxBzH+lBFZ9RfAZm4B
sRbbMPKzQFDj5rQwxfhw2sjJIN5N0qfni/q7V4xD+kHnHVJe2FWpIuArrt2807AxD+a0mFiq6Dyd
Qy+MSOBRTEyS9Oq4QXuhLO82NChKjBaJ32oObmlFZT1vWMh3/F+womKiKr2iuIXsxEHuxql9h9Ga
Fu9wbDd9YQjYESbNllCceqFyGPCqzBQpcSo2tNwQZjUA5whZYo9hq6UBXsegojkAw2udhjwkxcmF
spqahIHlHBsZys67YOm7JHs9vaeEONQC+820WUkEXpwDPE36yq4Cm/TTRRPTMtS60FYXCbcbC6rk
ncha0+E/K+UV5xs3ymHXn81u6V44ed8TXTXAHxqv5fFfhc5iCAaLDBc0JL5GJYCyr6lpn0FfJHnZ
t3SdF7YU5q8xetcC5gdwP/DYHPz0vRicYAgHmhhN9H0ZW5oPdVzrUPy943dzKkkdXKkShdMXRLQO
7gTQKI3Kde5WCEvSWcAGkSbxExJzyltel0pwCQYnTP866gPuQW6PJ7PpfEwha+8Jme8Am340P9SO
usgVnlv5s8hqOc8FcOglOPKD5LzG4hA2HzsSxJxWi0dEC5gAWJDFvo7QhrxqXnIbYVMPDmhWj4C+
juj7uTqNBOCpqSBH1oh+j+o/PZ/wzc3RXBp3U7OvK5yvY/vaHfm500CKA/BPT6YyNLkIAKRzflTE
fldNd/kM2OC0iK4SRYQixLNSWVj+/UBXiO5bcDuXP8vCZNVWMFc8XHD/XZA60ghRc0TmJ5ectUCP
kVDQ9zPsO6W/90r1Mn3CcImIaZxzeJal/nXl3chtgeoedHWbsOAVpysrf3P/pQ8ldlrXDjfv+9oA
H4V4qbyC9UCZhbi4dytCZiCKW5BfPGWLlhhSeKQTqlpcMaAzCOdqwN/N5ieDti/dg87r9ff9/C9E
EWp26kCGKQ1AcM2Cv1hVTZ0mp6+gPa2fOkEWru1Gb2zq12ceRWvUTZmsDNUfe/VBpWTrc/NwTtLX
wUgTfXgsrAhjZShSRPCBQw/uGO+/Duwxi5/sgdCS6pbi6T0Hc+d8JjpFfNAcZUWMoe4eaZIody4c
XK1GBLcli8PJVHtnCXPv5e1ajccOznmle8fZYIRczrAYyTL0mdtj4Q3HeQRnSf0EdVFpMorijQWp
1GWu17VhFPZLrUWVJTOgDVI4VBCZIYPg2/IZCbgCGZWhpUDKCefw//awtxUt4XKkq/AAkqGTfyc+
lhNc3cHl6RmiBbbX0VlcH52wKYYMrEI+UlLgeEY9uGHCndcLQH+mxViYRW0atTYZ2bX3wlifrYHc
9aE8emk/5HTS++4Mwe5tmA9n3O93WTap1vOc1sASfaE0kWCQdP1N0pNfDOhg1itDTsvjSq+V7DQp
ZIKd2ZxFE3VnTRz8VH3DsaoKRYCR8ITNFBN1Rs7PgoSnVCfSW3oPpBQZudymo8Px9lKEF0mpUKM0
3dFarSgW0s5fjnLXhs7QWjw2FalFAgusctGBwC0YnxjRikvXIBSU/RjdfU56vsqKyzqEWIhRNnS7
+STJv77ow+CsHhW9DMwaOGV/3bFmuyC90nxMFonQRWxaNLXGhDrjll+aR4KOO0fJS5w1rOCv2/uH
qFb1izqrD62qv8M2LklZrJj3K2MAuUonzidk0PkaRNTXUDzBjzrg5Hskh1mGpm6jWIBF4z3ntflq
FyIUc7uMkojNla2gNbRXvHvsBzcmCUjbCaLaiuOkOiQIo2jRVgwHu/gekVYGLTDwdboHGYyUH0IF
gmJZlzHErXJKyZVagsZF9mw9eogi688FjL8LkzbiXcWix0YTdIVYO6f0jmqbdXJdmodg9VpzyBFq
6FX+8nEFw0AjGxC39CiudjRAJ2V93gZqgBcB6kUvqFvA8/koyNZlttSU/zJe/JmBhK9y5Qdrh9gA
17NyjpObDNuDpRK+bn+GrbyLKQWTvSBSvTjQU4pxq3FiDrdnO0+aa64OPyKJ7V1bBt87YgL4DtdS
mZeSASCLNGCKB3wGBriIub6WOc80qhHcLdjPUi2sRCLtcK5SM+pIIO1aaqywMrQQ9t/EvnaB+J1X
eDi4V9M6UZZahsYiRn1Q1B/h+b7A0vW4mM083DJmNSyFQD9HV5c319kxDpGDQgOkAUydilHtVdIS
mHTAHPB43vr3DpKp9ESlkJP35IAe2r5ioZ18yKjqEqTb58v9khta5cpk2YLk67slZ1hFR9Om9EE4
cmf5H+0/4qiffuTFfLES7tb3+CqCSCd/IrtoCx/ljNnixWvFs85xn31kvm8nUNkvxUW1RZvPMEe/
Pr0fcdpoGM4YH1c6SVCcgiE2DlQUPQnYqDi68TSL5eoZk7qQAhwUVUtqea7tLRDUsvfdwsQcuuZr
QtA0oPdMmG0lSFJfV0swDPceKZp97oFPJOuYk1n+9gdqVJe6yVO21fedoS79TJJb6bSEt44lM5G4
mfUY8Mcgy2NWuwhsn1vebfheqe9GKijDg99oft3vZ337RkjqapM8g7xQucUgdrQ2glQIrot5hwWj
AshiHr2nHYNtoPnxnm6uBNDTdJ+tT9Cbe8Mrt4zWxGE8jsBIOL69ykYOH96Artk/p8ZdkD1r/SvA
uSlupZ/TaymtZbW6w7m17DhQWAiHw9af/p+7pd+BVzfw1x3XOqVFAuiIugvA3RnbvZiv/K5bU1fy
Af0Yv0WFRQb5hlm//kUmj5uz3kOQZ0JJvXeNeUVKwI4P0GH+SrHdOisSETODwsQRLZYZalGkl/3o
R4zEL+APWXXSiRDzhoM86S/B9x+dPSFEW7Bd4eHHPoQOzTCbzyS+WquMUKU61sTge/LaKqzbVyZd
yudiFZDYHUBrAMSrw4KA2CcdhAPfcLzG7+CUOly2EXLCeWW9i9KpjVhdSI+IKFeW7/UqjnC8sBot
BxXCSJ54J1CGocox0xWKg1KZ6A3MUA0ygKEniUGLSD27UIQOYkfIP57HJr9sRl1yuH8vn+G1XCBs
z+VgdafoIHqcQ+YsBWPy/IXjnqbY/QxgmKu1175rzT2HChU+5WJvDXVsrKM/xtxFhO+aIlqoCA7x
AIYcoIAcig8bU3vrRgz9fADtregMQLDRUJ7BzOZ00KWBfou1L8vwlSi4JajJnVyaqJ7JDK2cJ4bM
qpL9SDIwcvJCGPy3sHrfBtIjmx/UbIzIYbLiGCPsL11Q0Ydt4taw4Ifq44TmKba9PXUngKU9H0z6
ZWhgmsG5hTf59HKN9aIooU0k/Jqo38cqflA3ih1rdzRKlxee7vN70kavaN49jioP7BI37rT9p84h
kgCCMstqjCDsaDxhi6Srvhjs9dT4kcfouV42s1saJmlG4zmUnawCRC95/AhUHCCGQfVIGCEGJCoR
jIgWJ7C0PIJG3iJUEQX27gw/we3PAkA6Z5PysIUgtvbmqLGrCpslaCWZraP9m98e7G/Khi6Qt6KE
oxu5t6hyRBUZ4AAnAsZPCdRI3QinAVZoT+ttUQb3UQwpOKIQWKymK2e/98Ec8K6K/UofzfqhvBls
GKczZE3fenx8XQKmEZW9PCIHNeQwUva8GcX2PnWh1JWXjXpaJMfTDBB1+aIq90ndW5UvFc+BcjKD
4lye4WT1aZKdIo8y1VR9Kb8AuoyhJHy5X4qAmJfSBN0rS8yGrQP7ywVtwCn9cgHbzqBdZReJ8ULR
y9WgT9mJjwHRaDCdO75zNIfWeM7nJYLDBzHYwa7Y0n6vODJeCHYrNgND2uBsd8ovgBE8VjkOCXim
lTZdy2n9tpat/+aoM49O4zqgodqg14FF6J8aMrWtUBUAb8JjHkWtU+b5AZj0AjeSXU1aPX6wQQGf
v6PaJXDP0CX94PMnMOGguX18P7LCVkTXlVAwFkfoUUj2l5u4OA16pnqXdayjSWXtj8ltnkqoSVZN
+VKck3PyK9D8CsU4iCjg6NfrMqIb7GdY7F4mhIc1T4lzIg+R7QFEvYFh+9ZuNeu/ycDnt3Tbwl3u
QuOaA3JTGS4M7ofIi2u8JCKaXRkxJxsOf0Jc2qRl6bvfdlffdvJTrkr3ve8on1AQjGLZQzi/F0Fb
Z7rT6HKUIHUTk6TcuO+6Y/DJGvlAWC9YK7srqIFIc51RiXilzJBteXlOaPFpHmb26A+jSodZXl3d
FTp92s2xBUcv0Ke/42T/Eye/4u+SvfOGvLFYyNHvzYRZMfRJly6eRdiALTjrV7CXZD9VlwZuIeos
MGVFfLKgpnLXAlE0ngNBilffrwKamIBbjlxZEYFzS066bq8kYTEtavX+GyaTmwgfE0tDLsQxd10v
lLydV9K+mKeC0/7GKSBDITgi7GiJNVHIyyDzkLuB2cN+yPYw5D60Vxl3fmHutBurPwJyisKKPgo5
R9pN7TG9lOJ1aZLbI9n7VW8TAqtRxIh8Wds8ls8Naf4GP5+0lVPWplQUJmVPh/fHVnfpwX8lJHDr
TaiPHySulDdBiXfcxPoB9ZWThnqwyjcoG82u/G9PdbtQAVhPWZzaA5fOrVald09v52G+NPM8oAh6
8kgLV+Rg6MIxnMLnmhkvR5nUSLSwiAMV5U5K6ANk/8UOumZLqIB7JB1QlnZQL4i0LFa59aWEEJEV
9jqrJvwS2YoYXGezL1fYwHakLoeey1ykrdWG9wx/5KhBqg5B52Dm+MDyJYVRYQtzYDIgetiiaxxo
WXnc3kH+7KRUVOEofD3lUbbWC47lY/0YzRncJI9qs06w6Ze5G1Wl+zPpDgf5sTy6nJEgjpnL7Jxn
NTUZd4jif9siBs2lojxADfcnstJzq0ReRHjkfoSJdsrhHRlWFYikRTuxe64Wa2jlc3VGw0CYoAf2
UTH5oKFDFa7iACI1nG52ej0359knEMAxbSQI7DLqqYXdF/AhRnoNk9jy1WAvlWbCwocTke9lN1kG
HL5kDAsrO5oPalyYu+ZhLHKqHdKczNT6r9TNSUnjaEg2NuCTu+UL1ywqZ5d7e8QbuD73wPJL6G19
o4cwZBCT5j0ftT5LXq8ssU+aKP/lFlAvW7U+OCJ4AJUea+iogiyPa20jiotkdQwTCOQS/2KpHaes
IkhkfqzJgVtYvyVX7IhUdYF4el2V8R3bFS6EuclnqKaOPm+QlqOQvululpFPz/aGuxSzEUVsfrse
BrIjVqSAJvEzmcbZjCT0iduDrhEu/x85jZmb92Xk50nf2jycejWZrtJ9UCdadzVUhksp7R+TJkba
EAvEmvWCH2QZaaWOV6wefS6EKPpMh6hJcZrqLGP5jscGms3CKQhazQeRGWfvKmRxi+LyWpmeiDlg
G7SqksVlWYaR+XP91FiRBCLYPqIdeP6lNd8Y0B8vXraRW3Hj+4pQTYsrmaQMHjozK8zyaDP0tHdU
QqbbD1WbwHA4ZfLy/UZ9+VxSH2bEC2lK1vGhFCRR/NvcYwpOqVot2gSVRTbSxdbiYfLCg3SZCXi3
bbwzGAx7poatdTkKp5TwrCNqQnOwp+n6CWP5W9e7efNARgp8b/cXAZFqmYQNo4Z5IsujjYVqwWky
rgYQQ0PxCURiQZEl/ILcKYITwLeAPEsquLLnKaAV6NDD57Ovfu3iwhp5B/jp5EevTiABf2I1CtYv
ag/3cCSlGhwV+W/1aUf8yyXBpGc31456L0d7eK86Q4TjAwkIW+C65WxzhFnRIHj0tgFEup8N9FDT
+Q/c6bBN3cMsBSBFZkLxz6r5MXPN8FW5PaMNpPpn+eR5ZEo0s1w8cPlN4+0J9l0Cc47PLKX/LdDk
WnQD2pg2UcaU4s7BDNR2JHNcoSVPxAz7WTV2HZhFsnIVWbC+05eO/kqkLmiD4PL5ADe68zaXPAYc
ntSUGMfqmXeu5UdijaPUFWaPZzxvDP6+Gl1Qxoz6NaIlF0mGzBx91KYlFO83meE1m2lumKbpF8/d
ip5vcVeAvxS7Ol6iu42gnWxz+esyi5sCZgqbrkZzDEG2lLh83N2PsMzfYDFISaklsxiHtJpRkx/u
eAQGgwOLxx5wdF0UA16+F8EDdKZube8mwJxblCWVWQEO+nECSRmsygwuBwFxAUMcpXlKQwIoeW+b
CPLxNRvKRUMQnDGFhOK0DwL2oqzzIUsSg76BVqfOxFoFlgp5ToUp7u5AvyWnkBc5fthxbMFwv2oY
4L5ttJb/i53qvKRp2axrup6+46nttDWsJiGSzVXzxxl31Kj/w3sWHur1p7aNZB6B1bV0+zlUvM3O
l2+200NcH9Y3cRAriXbx9nvZXVv1h19euF2SuKQT/fZxbWwohzD/vbVkgus+EnSlR/pY+z3gvo8v
OkoD0Q56iyJOSAvBbutwaZCexWmGPfXb6Yz8u0e0Y7JvGxwwcuUC8i8CJFmLA/UjxZeXK45dkYB5
Tvs5DrqBSkKR2U6vZiwO5CHwDvz/HNmXDI6WybWNt1tEvMaMF+M0Lhu6fThO/dy0IeHeiV4LjvMd
IQmDTkI3QaIGvM/9R7ZY9u3MScXotEktIfQZU0EhDzbY1oipy9KuucVkzl8+lFr0LznJLQSMYim0
3tqYM05n1ty4qKpDpNhfC4QW6DtRzJOJwqSQJY0GCT4w0cKj36rJvKT94Z7AwUuBX9bIIhvBcOM+
dS/MXWmvGECE4Pk13TkjEr1wtzbvrig6j75KLFbKCLsUg5hG4opzHoMhNsUqHemY3Q9EWDpHOeJq
48Vbk+HGp9IX5jC0da8ERN2zQFoPW+cR+aKU3ituKMXANm37cLxZlEKOFTCIh/HmtKgY9nTgftFa
LyQQpuQUrbGM/wv5S97oGwJGZFH7GwaqiBeuhITwgat1XM5aNAaF+NL4icap6xwc/mpVklavKQkG
oYrd0hF3C7I0zRweAa00pikOVe4YPdEuCRnb+8y7mgdicOS4JNuR3/4ar0+GBDsC9LDrcQpEMLrH
/BNeqP6MuI+MZejx3Mjho+PsRYRrQi91cYx/p8EedqM/zCP49jSzFB7JYvIS/v31ds2NjtZYFPG3
R5pbMHFjqzJ0dncMXqXLbeWQn6v48YWT2lvKYb2iFJbjGOuozwCzi9F8DiP06bzAwIAuBHnUlLvm
Se+SR3aWqShFTiSRlhnkhw8osCDjEL+S3kqcFiDQG8H/Ba9IT76r1IaDzfZFSTy91mMpiYRTcm/e
oMZQF6UxbR8gl35TBjjO+q0v4Oy+Wl7F3uu9mkYLcoSmL4Hl6XX9TbwFx8OTvE/q9nxsjfvzUX3e
5CO+2XFFAfvnDF7ImoKGnWZuy1szPaoy7c8J8yG8+LO/N8E58rpMQewxzoVujTgBASEDBAByVhS7
iGD7dD91kEsTHKIeoR8O8USJutMjk9U42+OBnKUYeB2iFVbVQuSGNiAaohJZZzD+MFxZP/oYBISx
G79udU1ksSq+k6Eml3q3A3H5tAb4kp/pBRoktj5UemoL24MVH2ukPRPxopcttLoDS8ajFr32bU0V
944dH+2AZcPP6/ZxEo47MrNGW6fD+c9LIJ7nug1n4Jwlei15jn88nsEa/5MMCmggz3U/2vTaU+H8
lSsGXHQaR9zUIzPuhLAtGmQGyNJ9gJYfcUDJGKukqUE1Loki0m1iMX3TkgqsrfkhqlycbPOyaexg
qWG8idfn0WyFuV9T0Rw65aTrWc7iGXMznPuGnIb6F59noaYAqp7iNRWXldMyyLWZCtrOrKdzexRR
UOj3namqi9Lo9GZrrqGyfKmaePsue8rqEphozs1bJxnceDXDwQ/YYQg0bbLSCOdqeA5LDlK7nedc
0yY6wpXUyWPYJMOsszrDH9wgqQc7Z+epsTUXC3apsL2SI9QDlIE+ccMiJcVa4pjb5vsfh5at+d6E
rRFGl1qM0/UhPhNHN8ADHcO1rZ212+gJQC3hbLtyxk/M2mV92VExm3DAbGpmXDF1aTpHka7BHJ6n
WYsromRqhILXuQObY6aLMBoUAf5ydYZG1jDQr42zvWQiANwdaq4a7844HwZaHxrp9v2h+vnIqLww
mIYXXDUTRyTVN6FQNOyuS6heHjq2lH2K/V1lRrWkEFuMgJtZgiF4rWEDKtoFTdCIbDzEHuwQYWJO
/wXOlw6qgjeYddfBSLZ03j1GCqxntCQqkmKpaNiBsYP6M29anL/kg22AB27oDTiOH7C5YG65+Ind
FSx9Z46TanCWFeVBcB7u9r2TEot9rptOvT1T4BC0x4QOyswgGkcypLovUdrxvv6I9dDMkGaFG0fg
0RPOoFGaL/BBoajZ+SIEjIUdjPDPaAXxI07mu/ZKlJ4DZ1hg8in8PXWvGYAS4EjHcrVdWdSwTmCB
5ErK60jvrlEamdSO7ikXEHJynVgxCWf7gyj9QEUd+wsXD7/Vye3/MzM1WQNppX31CySj1Fk3s1y4
+fDitDv0TgYWS8p9ARaax0wWXU1l3ARA20EvTML8u9RwOKPjbbIgwN/GnNaJ69OmBJnBt+Ml30y9
eEmzjUaeXROxEiVCFY/jgILGysXJcIiQONT4bslyOUv9hMaHvt+dgEnlrF9leDzMqHhVMvEgKzgb
eLzdaHIAeqlib7M+bltggVXNkzcxRFrIQSfCJ+5wrqU7eRwsbiPQsip78aZ2wTotzOH3tC9DqZAQ
qtOOoOfSxVWyMd4AcpsddXv5zjmvTm9s8tN8xab0fs1Kyfyub6gdRmWDLsSV/SUlA3l2X2glFjJR
Kmn2pUmdKKMLuArQ6GobI9E96m6OQpMlKp0HNXf98xEC45mBXP1YvcrPRt29PJQk8IXlZebC2H5J
ioKCsOv0HWEfyNzgcsein432zpyPDGfBua4LGqRARoJfEc5zKyaQ0ZDwZp+MiKHxoDNw/g3NrE10
oRds2dh2DqIvPbMnLvlJRqescCNWLncLznFK4PFdoVXkMqCjuBHJxQ0zy/p6Lifh8DN8PAAUwn4b
NXDSeCz04vSRaH85sp165XfpqAoY9MvnodkjIrMhrS9etEbRkEJo8Dzkv+E+Ht5NfdjQeszOALXh
GfJN8d4l5S0eLNwzn9wgR/w9BMy40I03xc0pR28ssxmshaMItGt+4/O4UBsADsu/H8nxpst8dupt
+vuFN/4IA4Q6wf2rKxrCKV99lVmgYyRPI5MupThrATtUy3mCcO6Lw3S72GFDlfVdm9QDMboJeRSg
2lA1CrMkJ3hKN0Lt2RoVOB4HyruLWcMoiN4K340hXKPv0m1hUq/gJmOrSLCCm/suM/zx2ycAA3jY
ElFxxQqH3Fvqwi5OxpmqjkNQqBFm4mvinnuliKPex+m43UfMrU3s/nj59tbh/zqm+ECbD691C0Fe
enpfTaMuZ6Gne8BglLDF2EHq5X1vDZKaFJAcg0rSW7PKggEju7/gJe0DUM/zWoKrkrwxVu0b/WUI
E4/6GXNvyddFcDrGebcfOyyMGWtkh/R1BYwbluIaMrG/+0ZuHiHiIMwED7CTAh/rA/5PoE0eNZrZ
9fo2hMBwd/AG8tyWYqq1Vu/eYbVTMQk5kwQakmDmrtrnYnkX0OolBRlY+EMGad75sFjdTYMlXxhQ
IGuxGpp7s/zH2jEEFFe/Vg/6GzBCGFdliLqVgYjQwO2ZSuIsmZsBUL/0n403VsQnlzD+Sz+VwpXM
UXFf6gYTpfIPR712DLHxVcsbIQeG9DfU9MNPZL9UwLI9R8k+caQFYeLem28k9qXlnnHpDULa9o99
HCJt8zlbGZ8u9Muul9uiSBnUtLGDCvpONMwBYz7gzJDnOcNxOSuPqk3VdCMZ805x8YrQNy/GQ/hE
RMqf4rykoBiQyYOLvoHUYYKJr5xEeXIQ9BKPhyM5mz1LiN4FqSRVhUgO/yTwWBHvtd0exbTk8Bx+
FhKcy4DJgos6hlXe74ni4JEpky5ZOFKOEgREyFaMmKCHud9yfX0jTORX81YSBI5DstLD1/AiBmxz
Yhjp+LMPI0gibkjctUKN6WS9cZ55aw5vcBBNDljzdaMmntBTvTSK5o3NSzUwCyQtW+C+fXJgFVhr
nynUyztHD7HF9kR8caT6tdMal5CU7JBpfQflmk1i0z1K10LMkXxVjNbxllIz3VT5Tf3weC827Uls
kve56jKtuIxxrqaQs3ULvIgIsHMv67RNovkbC5HjH1FCIG0SzrCcrl6Kg2xpO1ZyWZSqTHRVjGB4
rPNxWDYOjIp7vJM1kJUjGckjrKpVtLjWZb83yaju48mZkyeL+gUtnae6J5KFpv4Bn99XJwi78dOl
QRda8OPqhxOMfzQ3t3Vp114syBCATEGwwWhBcq1q4J3ObZ/zmUAMTna6c5Zcj5EJzT5Ct75fAsJn
TvYDfedBQjjEtkVKYznI8HoVMuo/LlHUG98hHfvLuj4/Y0RqxdDebOjRgqdWvzWOWqxAaE9hHhU/
lEDzo8b54IUKP5DvjzUBjGl0gwzsjI/yNywl8Oa9UCTQzwjlkUmkif5/9arhySOLCv8SbHbj5xmI
OaTOGe+zfdyvDRWKVlwnksIXuA6Vor6zee4cMPBB7wgp8R9b+AGQugyVumZKEtM0iZ2bEQL0ydTb
YMgh36STvrXPtmc6AhA14Qpydlx0HT05YrziNveBaxzqj8YTMaMFYLdKQhX5W84dlDwNAUREJnev
j4l5+mo8e4Zhx4sYF8EdTflsIG3XUnndEzdByuVw20Z+xhlOSiq7DzYPIh8VPevTnKYY5FU32NLE
hYBfbzBRckCxtNDZgeVfLuso4qzI2fYnIkpfm6uhAa8nrA984+Q/dcKRUrNxYcezdAUqpwXXDeAB
QzmdFH2LJF6j+XpLdho48Fkg7LNV7bM8Jn5lldaAr47h6+an6aK3g4taKo0RTxmahD2ezsgSxUBF
u9K/yYiU/el5OdRd3bv1txFZ4hLr8QclrAcOKtXDLdHjdjaEMiNLxSNOfrj/lr/R/rGUmTkw/YgS
roFObz2Btg5LWHVB2uyXvVXR5eHsuupD26zx+zNvrqmLyl5zWCxEY95gJ2ihdXg8vkOJHzGmF47o
aWYrZQbAgdxF6rQ+NXkQ3NZN2NVeTlZ+hKWfse4X8eyV8XOkjEG70GFgoLhaCRbjohZ+t7i17HRY
hVT5Go07J9hl5tXSuDWZqFrGPM4GzxRf/N/gw1rUFtX7oaJtBk8sqzcf/sDmSql6iFFq324OPzrX
hcCASjKTanb0Htedf+kAAvD44epTo8IzZMujLjXM7FmF7aLzGZITkbaY8zGWkb7LRM1+SaAC/+nJ
doleNFGdEt4g1PfckeZ2JI0AcqSbCgEAs9aD//0aHLETQTiLbd8odSZiJsaUuHx37ERye+HKN7kC
YogJtRWx33g5udJJTMHKvrG5r15+u0KR5kvtynxmjZp8VxtYYgS2Msz9KW5IYEYV1MV6pxYFg/Ya
8jym/W2Kg1hC2XwlXQrdkL+OIus7X9VuO1LmM7nstV6VkGHXeMgfoGILxUuFGcUaxbblwdc3Y8wL
lSv7kkCmURsUiMpHrRw3iiaYaKW62dc4a2IdWK3igyMjPc4xsudmLXxr+8OBFN8uTzdUIyuEyI77
R/iSJjHK1qBKZD88wZwWGEIhZJ/ugB3BuZqnKHePtkVIGXuO3Wo43fwlSisaWBF9fus23jXbcpuw
2sjYYyHZbY9uz+bYVKpHSDFOq0CLf7IswCyEsJvUAd7J8ALxN1KAb018o17LrdjZRQGW9zwBrhfB
S37mif9Qz2nxEcXVAQypIf6/j7Hwulu/9jt5Ct7peDXeKQ/kPSFBLTIUe7UHF923JgsjxeGOUvUa
X7yZfeGSgW2L4o3q03dGbYBtR+ozxNNGcSMY8oDyXh9/NAN6p9m0GLvmqSh5E8G9yQuUAGUEL0QA
9CwRD7nzKmdqmeu9pC50GL4RSf6JtP/AZfgfdDSTFCy/WPxVPdkXqYXShyVi1qKnIkWN2hUMAA5a
eYArvlQXhHc9fnbanPz+6dN7L+WzJiN3hjJOq6MQGOeJR67kE0qk0cIIbby5ESMKad+N0mq16Vs3
uD1LUnkEMyX+4K3SyEUx030SB8jGI+ZFMSI+oykMtykGhwZrGtgi51O5kwJdRxTumTIRRMBnbgTO
43pVIYHXXz8L8oeZLkQ/wTbsP/lGmfcTK2qFV+7ImZvmx2yjvtVgyOSepdMvtdswp3rqh2vOvdkx
bU+Pgp/lXhoYmvLc2yhq6XvVHVEWArNnCOoVZu5+OlM7OjiOFCle4BhlpldF94y697troOwVzY0k
Wx/k7Ew4sZp2cll6Ed2zcyr990lpl84jjttSIR0ZotTiVUw35fAHp/pIz21WcFj57Er0VRMNcnKW
5/JICKg8p7xXQUnAzYwrakfnATHwu1V6IflT/ylCi4CAxDu8IOkU6P7QLSGR0RRYKeOeqjGzFKMx
EKPNIrRAf7UTQTee332mGkMsmV5Xtdda+0N8cddiiV1o6L1JPpUF/RIGI64tMoek7m3h6bEZi/B1
Y4qXJdj9nWCIPVIQa25r79n2pfL/Qr3g+r52SCgirLP99T3TIo3ocYBdzuQLmEC76j5kYfhlplds
UnRKDtYU/W5UA2ViXT4g85DXazOXda5Km2oU+lnxPRkDQovpcdkA0HBWbF3Thwudx7htSxv7gVhf
BIAI3Mps2dJEFbANxVhCHB1Lamm9XTHWLDCdROjcpApS3THqzxENJb9iiIvJepiyQn7feDbNJKFV
yqWL9OOdHxU2+/9pj2H7lR/xtBQaib5+VcPEHkP+5edqI9V6iXbWxxs/gz1JaFX2kWhiW7O0gl47
LxWyxe26M/BzIgL/nm75PM+vntCEOUBMbi1484UO5BPE2V37Oora9wTERI3vzBQCc5NMZpXIcC+G
KhYWR0g/2Xof/ByvIK63vqlp3DwLms7uP/jMpDv0D3pL+7ZpUlmDF4Y2V8Pd3RZQ8328mlWP/OKw
u/VGbTVHoQwK80+e0JuuUfFRVGCbrbZiEzeCvLeygfK459u6iasf3dSDi9LGFte4eKQ+wa1lHD7h
0VQSvFomw5kRjfVPiKZVDB2wolZK0GL1DZ/GNPiEtQIq4hKak4HCWXY2ZV5EDYsTECuSTMmUMskj
kQHUs0/l567u8hlEbtIv1QSxG/AtCe9q/PyRu4iDFOHa5HkoWlZZZprBKrOVzL9Yo4eiAiBwIMzl
huh6N5OUwJFPlMmUw9qkaE+SiZZtblBA0CScbvAbQHgM7dua6oEXWC+vNyPhNcCtaH2V1e/GVwE6
vFQnYqrd2HYyTwrnJ34Gx/RoGNbUFAGcEkwsmGm0OJKW3vh74J138QFBMAn0yLhhgcq07zihv0Ka
+uvNyWZH1JBdgGeFIJp+K3By+HXEuUnCB/CLNMxk2kRVMf4mhbVLBaQHYvn1+VBZSFOTdQlI1KNk
3Ivzj62bRW3L4yLB7qAYPUpNXHXn8RfndNteFJSZFkQJB9wO8pJC88jjlR2mIhmZzWVV2C0DhIvj
zjf3V8DiYZW0BZrkxBtilRH7LvBQCJG4Vf3tfg1roNRSJoPeth8rI3whyMQZn4GNwKyA9FxOeEHK
dHtEy6UgFLrFQDtP2alsflOqpoVgfU/1PM4azVf3Ms6PT5O466dohBnMDuceoi7Qd7Q13dfR3n9Z
fck+Y8wfJfrHcnxam0igSbVmGqeFppMH6JVOLIPZcyrgJP4hYwmoI+zM3JsuW+UUbCiN4bDMftwN
jSiM+gB+07TMGqmoGyEw9kUHcWPFyg78cvPNLVKgLrtUaDIBlxacdiAr3LGl8lnp04fjafVwg+GU
LWo79faAjSWeXUAlS8SwQ8hwlSQrVS8np2WvQai6ylTFhk4nhgfJl76M87rOjfvu30Q9m78/DkB7
oxkwbs0KlfMiZ3RomUBn9NwA09GnXK6wY9SRU0N8cOvj9rKYAUdrLYZLXnZs90qEuRsM5XhWbmt7
68PLhHxediCQioBh3Naheilz/AQX9h6MZW/lc1g/sCGW4uJU8rCQPDZqc/6v2vzs249ifiFmcrD/
slsk1cVL5XYTJbiwoVN4yVKFQyhF3ws8JDx/YQZ+Yr/AyeONxN0w81qr6oMvw0k4diHdNWRyaS19
7KE8sWH+nA/X9Q+tyf81okHwOB7gW/6Yfi1xfWn7MXlJpaMZZ58vyuL+pwyvrQ18i8gJpAXJ8XXp
60kHKLSbaspt/+d68Lgp1jtoE4FPwRc7jERqHEa95/MhF9KESOivmGuKsldQxZFa4eyX8uj/c/av
6uXOKmf8U89n61u1n2KNW6vOpgSUoIaBtZGuXLtNQwbawy5M7Q+iMLrv/5zbhPTEjM9ODkvaQLbQ
07KsEF2bW3ovc8iWZ155JOruHUaiTn1U7pe3gkHxcwlHT8ME1lRZa8sv5JCYzYSCnK1dT/GLVA/h
kavxvr8Dm98ba6VOxlPyaF9sIP16/9FOwBRNygDN5ldAMseXx8DtS9QXwmhfCFyNpvwu/x2A8Apw
nb0JuNowyZPd4l06V3IUWUsGcNjRxYWq7myIyV/dhsEaLF0Z2jRMJKTOJyrAC/x7Eex+QNr99dyq
3Qb+cCNY4ZjxBhUNsNA35TnlR8SaWIelYIm7SrC0y3ivHn/8V+GK2K20JAX4Vg4DZ4DQ9vXS2c8+
mx70kmc1WxSgVy7pO8UPeqOOTVrn0mhxC9xQ+qzwtsp6iAWIkaMTkCM6w+OBKOQCGTy1WweyAkN7
kUiPYPQtDZu6SgbGYAf2f4KmUOQQxnFG3HPl49Oq/bNH3ovTUu3mPgME0DsVyVIEGFA08kCRFI36
JgMWEz46J/wboeMZY5XcQQTlPluB+FPM+39dmJu/eS/9ri1prMkPP2iigMSFo/5aqVqz1AdMHZK+
9ZWJmxTq/RJm0nKDnDRu6bAJQoULdayyo/cx1CnNRWs4UW+r0VOtba8PD3H5NSfZ5zosNWCZE+Ah
YCgsLUgSvC4KuvPFI7cLPMOYAxIgPI3GIFACRByT6x6OskIL8MWZ4QKbXjhNOtYI3UCKyuPECKqx
WkCnkmk0LPPf+MfRX8keQLbUYpQpXuWkABHJDUnmN6CQ5l7/Zd0ktkb0k4mpCszWNsAcYhOdpaQY
XSwMbYF3/xlBrpbsAegvyMfZaElFBI61MFp1xVooy8hCGdaMPUVicNBxrzDMPG4pyTskmKfFo93l
Wy7vrV/gYO2hrJgC6FyGoffU/ajlQur1VRQrNyxr4+i/NkVpMfIggH80IEZ9spqLk9g7QLSYIMfQ
JET4Ooa7s0n95jcZfStWLts6cIraYrhzC7TScZ8jhJgSjkue3/cgId1SKlu+2eqU7tIXm1+BkPRV
n5q2mviiV0hhJ8AxWRYi7R71MxRLK+w9GRhQO29N8kGoiCSh8NwSVK2fDEZBZ+JI/IWzEdx4HzH7
qffBRwwBF3Sbw0ERuQ6GnxXEhO1kjgLwEY42EcH4KmjDkma49Q2P4gn0DGCdb13Rintg+A85Zrc9
GIURHVlRvGal1AowqY3h9S1q2VwLUvYIiGTd+lv1yLvwevK0i1UoHzoE4sWApdY4gWJlJr7uq59C
AJX+IrFaHWtgSXXEuzHRBx8r3vQODlJ1RSGocxTwnIyhisy8E2vCr0U1chg7+SY2faBCcZQ8FnNs
Y4Hxgd+FvHhY/+wfB6OYPZv8GYuUI3NY/sqpBeIzTtEtsJO3PbqX6zF5wzUnd1w8yJoptxPD6VZa
/sywiZWtzpguo92/2we8uyCIbZPBdYYdenGPmxjOalsypLme7jXyg2SZuQyPRKhF0tSUPACSnyUv
C/TyDeHLm+VuASL6ne7Xxzc7RylwFVq2eAv5cWCUr0gdQ0b6ZvIJQcB1P8GjIuDVMTPFYtYcSEag
2uF10d82GtOslI+BcKisZ1Q4ffDKAml0ONiA1jIcjnDZzXYVotCBOERi4FROOkRn2q8EU9++FvTC
Ak5C6CGNBCEQdsOBVP/IzW/GgFkFPU6e179aW3FNoFgkadZAo44Zlz0AlgfSuiMlfRAo/sep2bCu
ENaE8jpD/jS0njnfkSFynlLmb1iLv4iXcTx0pCihqs1hdq+f34PvvC7MBoLljP1isEevfDaZx0MM
sqQRWLn55XtMew3qddHZNRIchMlEPWkwH16QDly+LTsvFB5+Qfcoz7QljY5eP8+KpjKGp6BV83NE
Fr/aLxRViIIcCF1xRFCnVnXzLlqA3cepY2+wtzw96sR1oqPX6AotUyXc7HaCKJyekB8Zc7V/91Fn
vCYLMP3AG6Jc1FE4CnY4rGJzZNqa6+WMaOgsy9+mwF99C1sGAJ2P0J+x6sVrd6avprewI5Ie8nXz
P+j+U+F6+ZYwJ1OTGyaNE/ZwdlQx/c6ni8G+wg/g9lZ+R/oevvoxlDE6nMk+mm92nn7lkSHdXkqA
IoBR8voNLrH2agr4RrqrQYcXaR3NIssaiqF3iEKSJpD7gG8C9hg6JYtHElMnb2pkAS2/WsQcgDBD
UtYd7Vmjiq/MrNg4W4Znons/QDQHIid8d32VBkypd/ClovMT6KG3UfH7r0lQ4afw8eTNGuYP8oQh
daeO1LNV7PwIxr4j2k2df1/yD8cNbJCKEqTWLO+3f/Epd7QdHb8pQKj4AqCFb0AYaSck72UWbMs9
LUG381t+KDcqcCYY+641IgJ/3w5qdLyt0dwUj1uMxPgxgSbe5o0Qt0Pm6JpudgWxbVguURKs/qG0
lcYWy2JaQlDY9+7uE2KjhsRLgWar8BQBB/1hSzwJmzuNWd1P3o1tSVytgxPb8q+H0dRmcqROoz/f
HmRDDSlMMiuN1VtDY0jkgcNhzdRY6W5PA0oER6YOcEA4Drw6nP3EYhLmIa5oFQ+Ux9B+vhDdtAGP
iZ9dt8xcxh0m81iWujrSdXM4B8l3p36BkWqSAODaqXVE4y97uDLKx/tf+wenDAr36fJmSTWc2Mh9
lLPGBv3Qi5Hi8osFFjg4E8godDccYHGU5wpkDvGUrSpwwXlhZDITKXrV5peL5ftLIMmfs0mS8fyU
dEt8nwO6+MS/431PM8vmpgu2/o1/gpD3+u9pX5owX+YwZrxS2J0bRRFoeOQ4feJmhN25e0eVhHHp
ApYR/qxnl9oxS/xxz3R34QLzzepL+/bOvD8EbtkLGWyhmRPliDWFLcBDKEZixHsHF0F9OoTdRFOi
XpjNurJfWpG1LKGHL97bB4QfzuL+EJpcC5f4oHxoD9FAR2DjPe2XCgAF0Xiv9q9cgnYLNl+W3JjI
t86vxpr8YL/VIH2AO8cwfGTDmxxONcPGYbCN7cmwC9RnPXCe0aWzbWWg5zfwRGsperujljQlV2s+
XkxT2/c0xyMae6ynK9mH8E7FP0u3RauxuC96zpogCcsJung/yiLX7UijFrHRe+ZbOi9hXBhfo3Yz
XiDOggOrHB5OOhekbgEOTfAg4IcMpelmwk+8oWAPhGfY9oB991VH+IJh1kO6gHC0gKcq6rYhHqyw
8sIlKP0UQsKy32BQMgjWuoJY/tpgUoPeMLbnyHqzCiOZmZnQ9O5JFdJH2TGPw4J3GBVzt36CFr1t
w/zNxq1kgeE7eQvRxvTDeRHoV1HHjBK5FIRaIgjVfjERTcl2krb+y7OYlUDQjKHHLrzqHTAL/pDQ
1xhfqdxvCBVxnW9hpCuP+3gSsQc7d6hF29wOOdl6wu27vTnRfkfFCm/6qq/F24OEMbbtnSRSITsV
+/dAQC9TFTGFs5T33FRdgvXnls8JXME/9bB5o4bx6UtyDx9NurMi+D0EY0L+7lfo880hmDrsnSbk
17UiamyV8x+wXKjBnSe9D4/kcEJGtrLEt3J4wixHFdZHbJZA4SifeyaLTi32cmSbIDE//zxJlTRF
7DzX965OLcHVLFhNzpCgPakWOdxz0Ai7f9FYTm6LtWMZjeUrz31lIiq4vizv87zMWn632RS1Xs7o
UiCfXsCwGmMJgiOq/A5kv1ZftENypaaS6mD+lSCnbaDT9QCpuv2s2VSkrHBCNLzcesEeRoEg7aF8
IjuHDoz2hh6Kkr272NLChfcuer9u3EtYn1t1QMvysgv8XfoUo8Jl93NzUYA5f7v2iJOqvnsubCVM
Y9ofFck2Cl+G0aZUKJrm9tRcsao3iJAMok3s5TYxFfF2eEeV0gcIRHHzyl0iiEMzpmiQnAywBAP/
YUHa+pdv/VZUgZceArhtj724tP3JPKFjf4iQagiQ5ucSKc+TobOL7RLy5R8vAfOY0w/QPlYaDlMu
WAik9+706b74l37Khi4o59uwXbs3vwOnFlwwAaknbUthH2KB3dU9D6hUZBKr2KaLoc7OULwFVe0p
fZSoUo9QRqLxZe8fCzBC/XJzPrYzG95EL8hoqaYmq9x1mtSuIQxyOerLC9+2/7hRWlqa1KJu1qIB
eH6X4px++7mqAbwUh0zYc5bodFPHmmBrM7jWMfcle6VZRF44HrKmlRX0TvlkhHSj1UfwyatKyZcO
+C6BkCjXd/9pvhHPz/WwQ9/tlW5v4dF1FxvsAgIRKhBdNV60aE1al0DT3Y1LPg/vBLG/kpXhFM6e
mQ/LsdsXoR1GkPy1JLE7dRlXOT4r3GBf3Km0UDW4J4RlcuVdQivs5SBpWeq0TL9MWsFIiKdtvwGz
QxN+QRCU1rByg4XJmr3M0QbpDZWktKyz24ZjjgdQRtH+w2Y4yFvBRDID0eXUAsn/1gvSgGdPU+FA
gq4+vXlilJT4okzCM/uy9QKv5M/B12QbaIAOOydrJFol7tVQqY8nAVEv7BoTaO9DR+pKTQJ3YFnb
/9jrsIf1W1A+6rWby6EMBz122/U6aHtOd49bGh+Up8S/Q9AR98VHwka6aApK+hR1YnEqQ435/WCy
lbRf8k649h4dfXAg5op1MgMC46ByrCGGv7RefNlwH5isBlP2V0ZNpel2NIYYrjp5B7kmdAbcJ2Rb
Wz+ANl+or3jl5K0ehkpLC+IbiPgBfqiIUXMxitQpi82qvMpnzUtX+Ef6MEji/pYJEnrND8j1fuYA
S59oW8plcdFIP9eq/geKJdWwCj2rA16Ms1VTqfs2arVNkfv+by5UhF5wex7kJ2MIpohmK0lNBZES
MXF09FUraBJiH5s2uI+9mGInObPBlM5ajpDvMs9XJV2pmoQkUr7aN4gWkm5vYuOvrruKO9Uveqvz
2WEw1DDVP4/oStq/45YRwxGiBJUKIzC4rMoRI81KqRci/CLa/QLJk+0K43SKlwQ3d2S7D1DkbLPK
GPxuwJnoO5JvrlrYJBBmzu15GpadXS/Jj5d7fPT9FnY0ZP3ruXve2GFWNcTLK44cbKvohE3NB4PD
5ivshQFgGKayTq4kem4z4WoE0WW4RTIutZyNUu60IYw3rhIuZVirtB8HZLRmzE7Wmca5W10Nv/AO
pI4P11XPup3XPXQv+EmeRz89NmkOxwEXRA96BVw28RVs4KLDx0f6HuhSRv74zSKYJPMXf3RRWmCz
/nYx78WEUVPMC+UB79WSzMtDWRJK2OVOm6pwF39kxTfhr10ZSz913iINrwwFoieZ3y7QyDZ+kypG
V3EAxRMtN/+k+VbCthXK8Mf5/42DuZTF7MJBXMACnAQll0ppgnoxBm3rLh4DhMnx+u/7+fim0Z9k
/M8yN07Z4eDTadizTAhayKBdYwDu0BMZg5Yi3sl/uQXWYDApfreVF3BVpPu1jiR1qQexIuxLScIR
oBWHSjd+UAfZyLsu2pQJjRvAQYqLZtluwUBRcM/uRC1sAqgO6uBORWUGfuTS0Ly75Q1oYD5LXwhf
n8/a6Ai/6lAZRJTcmJ63cpHjgThk+i8/l1oY/Y4liDT1Gm8IIs1y199+cwx5mo8fTFfRrXMEgl8E
qVS7nwF+GoZo5mVeABTqSeQXW/liJ+uTpyGNhycwTGULLE4wCsF0MyIHxFaalFfAXFV36sDWx409
96zDotxDcKmWI1hDZ0XESXWLlB8FzGJktlfgMjl9MPgA2yMQzg4j2yHbDoEUba38AeLPRxymBAys
d8DBvZb0PPOuZ96TQlEosWm6tTKI/al/LpQOqWHLqTu8nvRlq/yvxwi7MvGMHzbkxlhsLQkKSenV
wSA4r2yTLVk1GOD4K1pkpm8RqYHvnxkqTRRFtkInn+xGdLxNJpA+t1AdLi2Ja457mJz2CtfCBLnq
SpHyVSiXKREkubmKMaUVyibLNjXj7cX1tmAerkiAxAWFk3uqVg5w3s4SxHr7gTQOZmppbPPzeWrK
PM4qJvdhMrkeIU9/g6O1fYDiS1CnVnrB+/x7MQ/D5rTcbg1Uk3gPTp0FqNAtq0jVsApO2CRya3uw
QK9ZqxITDbltg8WAZo1mFyHRlGD/I3TrVuwuQG9gX4b3oew5AysEW8HWjvliQNyHjGZ1ov5esx3n
teFcdEeBMYRKOb6sh2enE6zGUEF0MUSS2yrHwVOgoTMkUmuhhwu9aIYt74anXDgA6+t5fVP7omQN
kEjyDqLgb2nsiHFBF0s7rw6ki2UzWUfjpagWMCoju8Q8aCqBnw4xUnBq3AVCNbsQ6bnBIo/vsKeN
izvUL/JLsivVUe2WmBa2mBNIigO18RK7UppTmZBsgoVRjrmwYzUGcftKKcdVJiGYzNMGFTKtzYfd
LK3whmgznfMM2m9HkZ2KBTFv43RwWylCGaUUSksw7mJQ4KFrCW1sMhB5DnM76HaGZmiKB927y9NG
qOWXCrGJGWJ5YQdFOG/7n2eVJjyaM2BcSq2wuHgX5tlbW8PWcmoJIdC3A1dOmb2NZLbi+fM0aulh
Tuy9wV4ZGD56SVu0A0M90IVvsFeRmztWnt2A56bWsMFo5ViXWvaTdYC9PuvHe8NwLHBdR/702XJL
lT1IwhlvpU5S9xTVTdbKiIEIxpqXkQZ8MTFFTUMn+tB016ub7DavmIZCPopf+8DvGdvzXkeKMTZg
5FoHJdyzwRRF1uTJLfD4zb9nUQKfhE3UEEFb4FCKHDSi/S5pn8w7fPSeFme9D/qhjR9mf0UUQnmb
P/vozv0lQlKinB7oxU0T561Z14biozVC7waV/83ScrkvX1ogjj1xfpT9plTAmj+RUC/gJeTBUCGB
86UJqFy7hmZ0wUMk1f8GJ4/U/EYeifaA//J0tNA6QBh56signAR++mbQZ6Wu+8ELwBPL7MoObOPt
JBtd15jbqLDIui92McIGECODPuAk4n5Qy8kOGWXsoyhsEPkKZoXjIp1FNVjT1cgBKDEA/0Ttdolp
VXuloPElM4fUxlXrFm0MJCr1q8CIwPbCdeMIr0noZc6eVEqkivZDTLHriR+FUUlE74M+2pcE3mUH
h76CmCbkibOH+mUYyRDCz9LgIn99juba6GqbCC9suP6cZaeZSPQoCVhCEPlcEsE6GdLCOpUfSQ3C
WpzITl63hSjDVTcw4Hp9VLzB4/Ea0SwrgW+LeL283Fmho9vysQr+RcS2jhlfSabzhQppFXs2aXbG
ntt6MWG0lXwk5O/sltogzO732KyCI4U50GfKSoaHYzCpxGynkMHZtNmJg33vJUfpeKCn+oMdw1fL
oCFQY/D/MArVCRBN+zVZ/zo7h2qMWfhJ1beGZpcsffFnPnEnuh/mQCCgW9Xn38FQxHD4dyi1rKei
bNqdJ9n78oukJgE56PZOpfYAY6DpOeGy2dxL0ajjYdb4zSA9rEEr122bMr85PO27HL3pfTDYDd4W
nk+BA0CxBxWxZDNQ4wvW6PHdunChtxVvZhkBL7KumHIvjwUJiFAAarSHRDaUSrr8e5x1EjMT576e
pzleqhixfnV5/AFYMRPcQjvexXE1ANc3Lrpw/BuO42a7F/hVjGAGpCmPnTASwx4qfISnSDVgsG4W
xK46Yv/VUzyUCAN7fR7M44hAHt3vW3Qg8YD1NjhQNtLkPA1fLtTrQZ/u5SSdgx5UPNe1ZaKOfRaZ
AynDXRqju+Zs0kW/SpjNucRqDi4KrS9DR+oEF23o5xKNVE3X99Teh22mOq5ZrFWgde/LCYD8gvJK
kpWItV6X+ApuD050rUlS9p/n6UcZc7OPvrszSk+KqwQaxVohzNjf9jqJ7zXTCjIK/ErUwIYthjxP
Wi328KPL2+divJqL2zcX9BxsE+Tx2bgzP1+WKIL4A+b/TSvPcG4EFTb2ctIs5t8+oeFL5V2R9u0t
OW0pKM5k1L5ntE+qwfW/fclQpWbgUdX7yOdg80MIX/zzYJAmjfO6porP40w7i4YUagB/yIO7Q3jC
OwZl8IhpdHb69JY+Ah4GV3g9rir4BduScFFXyNDgLAMS5dTPMQf/VVwS5RnbYPy0h2fJKLqNjFky
S8xlTfjmBubPsR5VjTm81LI1G0TO8EWMjX2/dsrO1dFlPuTCTWllHg5d37ytMs4otZdxer46pOlm
ptEOlJAmoJqwyZCx+Cge27LI9Kh1DdcNhGQCVJkeWRXTCNjUmJKF45kNgxVY2ip9KSNouDaPbP+k
R1FJHAP2KI4ZAIKRtPNVXSXDZKw2yYpHXrC362Kaxb/MC/shTY3/vBKICGuAappdmPyf8PKRTDjO
moTupYRG/iNxteNey6RkthasXM2zK5apfPY1Oa4pV7+dRRIT6WHi2Gu1Q+zxmlXfDWuwyGyT6Ior
AWC7/k4kS6OxSKnCfKEOnhJx1lSw1lpFbkdG8u14EHJ0Eo4acShnFMx2zxyb9L7Vc5k7ustKp2Al
FcW0LOs2RkoDPfw9QALYHydhx8HUF3Ak8TrW9c8OYs8MrWZF0fDuw0nwUVHiRTSOJUfJ3DU2IpgD
uKAN/HuoVlBqkEbfx2CGzUO/7DW3Bb1srA41w/gbH9TdPtY/7HO0Ncw5F9jff7E3KORlrSATnNCb
aOHIqwwT7lAiOSVQ259JvRDNaPH/XTLUT2CpmXEzQ4dhTUDybXsrWcnLBIzNmay1hJ6bEVq1+1iO
Ql/ADWKu4FV057rJOikqCEAjtBtcoLOICPhDh3OScQWQuTcobYL7I9IyvvuxDmSYoFs1jJ8X2coH
xK4iC77FLq2iMuToMg7kcdY2VK1DLLM9ekhkFkLU9Q72dPw9tzZi50lvDkTXkGdgN+n2kDnyRRtO
/S6I4n89Fvf7Atua7dcx0RpJTdRijkhKOH50HUqHj+cAaAw11KXN9Fshs4IQyoayISyVlF3At9KB
bRBZXWRYxK7enrbAyTs3oceGYliIepaISsJuf/aWQceiQ0wA/xMqiwj87KI6unMjWfNJsK/MZfl+
t1i/fcK5SIn0w3WtKQZwEiVUMHel9bJ0sMYJkdT8OPV0CyOxihchI0hBJBN84KDUxv/LFYbPO8EY
Pq6BE4cnuXg/qgHeEtQeubLrObODaPGhJx+8RdEG4BaxpwdqYMt8CoVgy0+46YsCpq7KtsMhVf4M
Qgw+kKFvIm2n+DPzXsq8yD7Y678JqfDWuTQR4al8zTb+B1zwXfUhysmnkYTYzIYLj3FuljPwdhh2
3KiXdrOPHjwuQob9EuPk9RdU44qwJtXg/T0E1G9Vq0r4BCrs4SMQalgxIjHbteCe8ZuuqirxVkK6
If7Ez6MXN4ICviKP+vk1NWvVDlogHEkpQmFRxq5wSg0ec9onwwPiFL0AhCZRyMofigqbpBlJ5Fj+
gcZh2qPLfUiM0VwCFW4Inil25sCbDOhPcgtyzcYvXohq97gtNEo8VAcFpcbcUYgTEEUkpkgbM52g
CXR4zoCB/1qEr+hHx6w07O6kQ8sC8P7W4h78xvJ0qs739pBu8BThrpxU7H5PRuHdtvfdGp0um6CB
Jmmrrg6O4iMGEMvlRcT3eQsSasIwPF8/K5F+EuVMROXA6x8NNNeuUpqxFXwWwckoAqDNZRFH2jNH
kysjacKR5Acbj8fFGGrUyn4v7O3DGjwJUaHAPbzihxti99xMS8GlOLit+DZO+2+321yNhgdOS7a2
zeQ8NeGOg1MqfWSRXiIMI/x3GH8jMd5u3FkD89AbR7l033YCRSHEZ3VxcHIoPxdlPeVmTdV6/q29
/RlUKULD71WRXJpPk0zLZlbvkQfQFifwqyKtMm4aH2VeeggLzGmgJKatJW5oUcXo4asJ8eiLpfnV
X+iA/wc32adtXPQtKv5WwLrqP3b6rFtuwvi7fHbeu7R/iEz4NwH99xTrkzMXC9Y/DpnLWcd/R/Zz
9QJ7bcOl7DEWjm9MYjTFhZmXSl/fVnr6goEpPxYqyv2O3mrMJE+iL7i5ywEb6nX1jFRdOhN3cMsy
lZFQGDJhXwgRp/rhuXNvERWCBXaWjt55J9ZLsn9g3/jaNjUv4K7SMJLcBdE/tAZWCNa3s+nvmyPH
iWfx2nsQx3XLCKj3N9KvXzaZlePn1YinWDYHTA1ZHnvcY5zt6kyE7I5lBam8ZoWmisgQxybrAP54
1nbllInrPlS8E16EfIkx+K67ZRCSip2lQqhNBEErie5LPythjei8VjtftL4AEtV5Fx+GytmqpV8R
mfhQcBZEOhKXrhCTjaUSPgSsEFw3dFyYVhu6Daci8A6Q86RblRv2iYThFhgeJCc10bNPKeZGzeHN
csfVFndaw2fgqLvK4VT3rOl2I8jQZy7uC0Hv/HXYplnBuov22BQgmalpZd7QmX1hkTnneDkvO9zv
f1293cXe24cJyQZNn5z19rWOlepmWvJmUoyJTbTDdb1SS6zEKv+JCboeCkkAT93yOycjgV9Jnd9e
sV4JgrII/ZL2Gk7vKSfiQrz3RRMey/YdV7c02Srrjb+r4He4F1KYMKiCRxxrRM/GK8w5aVkvpzHY
ZrpOYWe4A+LFIYSwbA7DREGmMKuknebYZj3dH1FqubRjeeo5N+0g2hFcg0jGA3xm4Q5E7X41Xmmi
Aj3qRbAwxuVe9DiczPGNzg4ushQOu0n2NXVp6LqdEIM4EZ9YeyHt/ndFANmJK/+sZV6aLuiaRHKt
iqTEY4wEEuL3z2mAkYQ26pV+RbJNQDfYw3NHVzz1+r+3kNnOaqEAkg4AXEgIjHiXYSQnhnTV02Ip
3ZUvH/eY0wXbmd6J/td7mM/X7hi0Fs626fFtlaZ6p42LEXWAGqI8XGA1j+PmCQwzfD6IZJC4Eo76
RNAcYWlK/4Iei8w4wuyBTC9+8HnHG2T3pqGN1A1ywwHmTLfHFyZa+7vY9idU7y5BpSJXc3XcCtX+
RFOss8NkTCYYGbgX2UWNPun1QCgI4MHxJl4oV0uwcpRK5JZxZTqURibbUOWb+LVymvX0xx63SjOp
kK1jdo7xpsC/7BGTjkdcQ4JGLZD+sdY8qXTt+clpocsmeXQo8Qw0r+dGyJzj3t67JBN/v9xBpgj2
VyMaYjUW/hGYluZ4P66E8pasngw/q0YKw83mDKMDzpVgnNo352P3gkNBwriNuY8K+/3xclOpOcO6
ZjnEJvECAZuYnrXRH38yTB59bEWVMrPm3qnjMVAMvT+eNIcR13RGshlxm32OFSe2vFar5EvVVvOP
N8+wKg2dvTLfJvd/TW3aAk30MUqCzWkMPy9pV2zDe0mfv28aPoTbP8seFewJB0aSXMvePEPqo9q/
DQfhqB8dj45Jw03rz6TzUdOMwX83mMpJpsx/MVqr3b3h2MYXFu3d0bFZ3LjqnU3Q8P3tLDhvltVk
4ePUCDBPD1pLBLkhajt/JvWnfwJNfXkMlfYqRC7Fr3/3WyWaoqcSAAhOiJfalaputZzkOJjZMMS3
DNUF4b4XRAs7hnooR7flV2oLzSIobjJeXHXwjES1KoVs50vupWrYDmDXRGQn6uDrOzUb3QPXML5m
Hcm6pmizPedtSoL+OCwprdWnJ9B2XSDXubTXFrdOgVyDZ0lKatylgOVj1Y+x085xQt1fecDH6GzP
9pve2F2bh43/PToNQGmcOZRAEYOtyc7HRYqb37as6gFx/Neg6DQPCT7V8SJjiwibPMa4/aC1yPYY
+udkMqCHStd0AZCrZuUMMnFwIK1zh6M3O1EyvXgpaZBeOzkO7rYlwbSlJ2JQx8FVG8oDyUWmCNuu
xSd2lBXjo2Kl1RPMUDhCdYw6WBbSOXPxVY3ok9mVGtl5QkpMCbuXT7MGaL73ppKJSmjX/UyeBY0i
sao2rG5CGc4EOGXZzrov2p+wG3VRvtnN3tePnUxzYFcdHpmr3ttHm0VydBpRh1BnKwN4xS58g0BC
3QZDSNLZaOI4/zXQdjOWuoh+QtbFmoTHQLoy9khAcHKINToOwSkVSVMs47O+7dxn+1bIilWrukDi
UbcpatvIZVHYpuLYAqVZYYKqLMPGPa8tonHO/79MHOe76uJPNjjKA0vH5CUU+NrDdcXI8O5f5gGn
VcQvzOmL6uix5scEWVexw4kkhGRQE3fVJD6HoS4nvTetPEqcvNEc1KcPkIYr7XNfFlGBx2Vukurn
OaXFhb2SlokV5VWL2hcMKCijD/w0dZ9BhgpqlGJ2v4pIw62Y/dBbXnZNmusZSeoQhwmXeSekE5sw
EiKrWFAUGbW3l4vcl25G392uYjslJ9/Th/xcIhF4By0wrg8y1EkPwWk1kQnxVzZGeXEkfWM2oYlF
oq1Gm9JweCHG49pXJM0ACi3GLmTIng4VL0KBAFFHi+QuOplM/gZ3cGkcOyjuVgfJeG0QiJjmQmIn
c1PIi9CFMQfF/xAdxq2pY1o3Dy63n11/joJJAW5QXgDgWDKUAgXozSZtaNfRjhxbrf7GZLVbmkqV
VN1vK/BxrnyZyiZVy9La57J8bTtCHVGZohZ4u+Mx/myF1/lSRbI1fjzoMKQSxFLmmUiSXYUnTjMo
B8sjOTaRjW6FErNx7yKAYx5bmqxulRqX8FBKDv3mXDN3tIbJ6dtK/9aiubeeViBTh9lYzPfT5aPt
Ge0th3a+OzdokPxLYIK7mNGgo06oO57lakO4FK9gHO2hEoytI6EDsspzU9HCoxBimDUocR9RqWhS
Sf1buNDPQwO7l5a4W1xHhyE30n4iBhvfiKnvHwHAp5Azh+qTWYD0g8wOUMM1OhOXdFJHVhHUkTFU
pEsPyKzqmsBLw/tcIm22dEknxV74JYcKms+tlgMDhjzzBsBbhCSnuHja1utEISlLt/WzDSeahqrC
L4MSkSXa+r+5VCbDNRNaLYNot/CoxgviAseU2uO+ulZjNIYSKGdHkBNySviDFtYb+5esslWmFxAf
23qXjlzj3mYjlZ3+uIqbwWExkRT9bD/ZmAmRAzAlImfSnO7/i7lQahCWKeb43DOudp6XRrWUkw2D
DsAKrJ/T4sy9oNEiyL2ZeSMuKCVgxkUtjRZ6+k0Znn6tKehydY6GYHwwT0Lw18ppFx7x269ecwOG
3FpoU3P/o0tAcVCR/kEeXFWDd71s5I2rjtjNHqKitEZy7uykPi0yjmcoPXPycUzJ3SgAJMyrckvO
vmX3kVmvkty+uoFx+02zBcX1/M7Z8Ka28dp0m4NPyqE8YplI7UZkumruJqr6yl7h3UWZESMG6dNj
FM/MHzupQKsEPnxRdzN8zR4VRyCRc24FnliS/oppmo/+thwATVD51aEmGMoTxvwmYlQUJ2PJe0Nj
lJwiIBLi1KRkXby0SIRdF5Az+b3my5kXyfsNxPkpRANleosji6sx1rYHIfSnV3cOJufYhhd9c9Ky
hixvWs50wVzus247nPjrz8laSWG2nyR+8CjHLt7zEj229rYyw2ZXsYf0ARvpnqGgT+CDtDDptCX/
Vs0hhibkmwaUil2CRjomzBu6SMIkSewm6S/1rw7/mvNbtXUg/rQurfvFvP8yhhqOxDcnWB2Yz92n
BeaPaYwVKnJylAfN3j+V8ydVEp95EK8LBgg1CDWmP/2AKnDgpE5c/RPNieUoGKlqbkE3hDfO9wp1
82tM+M6bE0kpISAufOTUAfRPKgpZRCNeRiDKm8qNoI+MOttocWiJ8HA/mBk4e3s+oAofpzByWKLL
hSBxwibuGyvKHZISkZCUTAVtBZU6+YOvIySeIxmCTApHyAPI+z2rvhI4cr5Ma/iYpdIbu77wUhKr
ON6lcRaiBFj4nZOZxWerML2MMD54UjiloMJvHFXKPqH5oarv6cfde1vc6oOVv1yYfsJ/X3Js9a+G
YmyHKijtpfiCqZgAwr4sq73QcVa5ITLgIL2/QDsPmKLuLl99HUD829I5slGuarWBnQjYDIXscd3v
Mz6bIIXfO3ChjGpaLy/obSw3UUqW/Oh60T60ZcpzatIDbQReS51Y53SgvatgnmQ/97PfpE14KZbs
O+SF6Eak1nuDPBDFapPja8sc4TwKN1bwpl8funD90QCv/jJRpTJ4/jsWd18pDg8kvF9+5505FmK3
BW+ddkTm9MJZXoH1FL0cZ0y1OgbkIEdQQgu6/Jpbs5l9ZSvIBPcbOFF46x3y7JKnH9qAEoXP0NpG
vVQqfUWanwy/TT/hhE3LPvkUUvAqj8ST1jJpNIdhlQnZ3PHrX6/dPi/FVIZWC0RMBNIHvIoc3bS0
p+lrJ+RxcHZboQHRvmUBV9TbzD8p6H64LPFhtvk4of1sjvjoDB/35wnRXPSrko91UfSHZNQpgJbC
7kpQ0IV7RFP9zssXO4DMbVcM+yxrV3nvdAc2ksknmKycWF8+ziLqo9DjMzeBLf/sVxeY2YfckVOp
iJ3YE74ziJAoQIXBq63jAPUnzlwMY/AuGYWS9HJR7x3G/dtkSztvWb1Ynl92SGwMub/3g40XcH7k
O3O5JOLMEXE7vK3DsCIDwGKoWjMfUeRdorOSVB7JR1/QBtLz0825rtFoXEL0ugmAAqWjOi8VQft0
T9Ca9WMLsLeELnisFr23VWDG5JU+BOjqCIOD2WJE3CBCCXk7Ozw1Efb9viPEUYriS2Twr2WpOYHS
qbc/tydUi64yld0gJ6TPtth6lseSIZ7Qz4BD7sK7XxsPReqyfKtWEo6mJ9uc9TRU01FOwzHSxccn
QpU4KaKYR0Pe34Kw6P1m57+yBiqQMrxw+Vwrv8NbQRrIPQbM+oRcG+n9Up8dS8SSshg4UZ983oy9
JemXLqu5grv2ZBszxqVT1GEu3JlYkdmhuKI+1YYji95HzhKGuv0dm7OQUBNDHrXzQ/58ez/3dhrO
Cf7kcqAC97BMGiKpAv3alzU/oJazYNWHZQEXGnGVN06AnAUzyS2e029+IZj0zQOce50vE5rbLd0B
mDhBsNWgJNv9uTk0vAfuauHcZiwkCoKJN/Pm8whMFWuNqDfzBqZwFFQcbtlroBx9JBOezn1nJ5VL
3QsQ46x4yd6KjuAJJ41Bozi89FgA8F76kpGE4rhFSHmlEz7bKkU/J684P5fdqP11fiNqUpadKqSQ
aMSFMbBdCzqmycbyPC5bGFXwNZZp89KivI/qrlyMpNp9JsrNujXQqmnd6m1ZPRh/zIWgSr54YT1q
VhfsV0xhx2rot03KoDUYXixrmWLbrjIWqvhhoSR5WTkqiMcqEe9HKp9TotXekPa+amHbusvPXUF1
muqzB/4TBlhFimlGgcjZYM/n+4Z/cns3sUvElIK8ahGgmVEl8xSgLQuxPEu3CrgsJqZwSKCCsVWc
egShqcDgJaB3YKZp5CBtrrnJ/SLaj5C9wrqWG2RkFQTjYZAUNpLnR98uNpp8uPOHoaddo48WeQDl
mh8mXZvYjTi83xT23ILqboLFUJnTmi4n0mwLxwHRmWFN1JVIeOhBN0kgWpgknZJ7pVEQS6QbSdix
tyrrctngBr02lHC6opsvRIUozjh165rfcmOsIGQkXDM4URhaEaE+M5A60dOUvK32z/qv2YrJmZT8
aWvngTNhO3tdXj015l0fp3WupsGKYAorkNUTstEwFwAUSKb5y2u8PulkaVGR0/i3e2l6G5fosxG0
rjPq/oaJq/DhaR+XZUon4dIB3nHUKJJYXPa8RYMgBvPLuw16U9wdWFA3dtTjT3a4OOVLmNrE31cd
WhhW5Yg8Mf18Q67nSB4ujZHJRTJCnhWecbCGxBmPLhI8dmsRa77H7Uez1zHLHoxFgiPoOvaEnpXx
ZK2ZX9ikiFKHJu49AHE37zXEMUu9fVGVBvZtlfPOnSWdGs1TZRevsSlT5bBV/JJwjs5gxe71vBIU
MYKX6ElCF7ir8DJdWCRRVTXs6rjTN2fio6tD4iT9uHwQa+ASF/bFj9UMmUJjBUBXC8A4i2+QlT40
BcLcsIfe2lQn2da0XvbPKlhgT5z/SV+SS6EfdKANg8MBY2m4XMRomcRvH8qavVWj86N0sfkfhJOP
p2NxpYQkvSASjN2ZIRVD1/bNDt+GM/78N0ZipGowN/Xkz/4G5NiLAL4JmTzcQ4JfsmmjYSpu2Hwq
+C7pRi76l3VXdIEY5DYhc6cR5A2/duBxnwUToQws8fbQgBPQILMtKmmLgFNpxAskrYuireYtde4G
6H27Y8/qQuDX8MnCH50lS05h9LICvbciTZzIBYVCsbL3X0G6kdlqgSh5EjNrnInYSmraarehsZQZ
M5nwbPD/qO1d6wjzTZER656WXPljnj9hVGByS38mhOwpOYGAq0XzgkTTMw90mbff1ODlapAe0mKr
yJVaVV4Cw7HO+JqtlSpUoq3Jqbp5oRFUaRAp9zgewCKmzHwYB4olITnFV47ztJRTCOS2pMEKUORR
fP6TaCrEh3JaaMBF4s4NxioRXRs6LvPvQIgiPYsmZ2EeckB5AUUyxBTaYVEwrk8qQ69cwzQJYzhA
XIRjCrtsAOQ58eqV6Vb8oAT4zNK6zycs4sQQOGKH1iGaDQR6C0rjy8r06TkbkavQNZK4eQupasMH
hPhjgiSpP4qfjpC9APqIZEF9Q2hxLrkrq9rIm4/5dzSsH6Z1RVxCtMXNYAxvxM2Kwfz3gfvF9Wxc
jffWCSf+9+/fswuEMLZJ0s+1Gm5dPV1a8VBS6hpHWGt0EbPxRMA0gdrkaw8vZIuQoB2KvNlokfRr
btV9eoCAWRYn2fQGOuk6kYrxsOjfmNU+aTrvzvojXml4Ljrq/LERaCNLtycnh6eP9Ktteo/P8luk
gSRSZmItOG3jI65t8K6CFRtsMw89HP0YKW7dK1FxFDmFIk0MhaqAKJLBpBI1xgSOm+DK9ckcAGaS
bi55KebZRe89cN1e1VVVgcW5ogudZsI+D0WejshvC+Gqii9hLRX4L+RyEnrETCAGL0LortM3Tobi
1hIorY+fiF3FbHx5MTEqhYp0lO31Hq92+3a/IYUtwA1GSIyBC65nalVrxen2LG5FiVNseevV+Nrp
ndyQdUNlXaMGSFg4AuMAgXBJnbrCjLiRAlJIe3GOIUnBu7Fn28vokxm8PiqMOEzB2VY9A/VDe/FL
kKXoFUmVx2peT78HMgq333nIWgzqeUEmsyUdexYqqjta7Iik1pFaLEWvjKVcUHz0FNV4DkghJktr
QlYKeFfquMoTyECWJsUwAUwGJfOaqoTS9ESEuZt2e4yuMSyDl/xRAm8msK6ugVxjvoXB03pIkZoy
7597snk2Xqth4ZCBfLKsjPrz5UGRfAJZpWDA+5NBewH9aG1PQBtzFejPVUqWjY9piSCwsblRKliz
kEGzs6WDQG8+goZ2yAm23/3HTR51cd+/iUaBhf7BvpdNVVzJPxocU6NJp2wUc63d23VbBGYepjPw
wmpGg/u7DP+qH9SHHGFf84Cjs3UEpl+ZHNFhvmA0PimZRVkOpOqWnZMRgG2XW6UiP/9wEEM+m9mH
ipwb65w0U9GmkaBNI+S759GADkCI3JStuUPSYsXBh8NGKUSQ/pA471dsfxqYTxKuKsazebaJN8iz
/f31+qNZIM+1wRZSNSVcUIe0EGZ6V+Q/fH8iEDjbIxg3+qBDrR25Cpb3HETYE5GLzNwzGpnrqigT
1iZ75fLGjFkXWUjfUUERVHv379aOEtcwoOwVLYtRI1ZiI9mSqrvD269hel3I4FUUGf9jvs154lmI
n2ZzLhSDvYxdECDgdhkef0gUfKsAt6IS7OdkhFRUPgEActPLu1GPIZlQ2ZUsGVPFkMOyxmQLRKQZ
Jsb+W8CKdDrclh66NmDQK5dD+Lv4d8ba3brSUV9FX9xdkOTzF6mWaVCt4gj/qHZN982ibM54Pdkn
dtZDaelt8i8HZyQEzTDUzmOb5i5YU6NsonoH6srh1ot18NiFlm1v0FIvXtfOKmCcB40qhoEzRK71
lb9xgZ6avC8qTDRdcco5o/jOqwCqg4W32TMLoFaGjKwbVVsG5nXTl1DsOXo2h/iQspca4J3rgJrg
i95mqn1JTESsFZzfSrgVeRW34j0GtVSW5Jnq5Otm8dk1WqyGw14IpJHlGkf+6xR/L3JOHJsmK2VZ
mx7o9zHYC+d9A/04WnwYdzKlMNDJAKicBLgt8ilB68UpIY0PjSYFhwXAjz4ToCDdHWS1MvcrVfDO
VOpL0nfu/9UTJTSczVuMXCcew07sOoYnJ4DZSksGn6IDs2BeLwrvwMp6ME0Mm+/C4IzewnpIr/Lj
sCVYkuBoYIBK1m0GKCcwEDykymK7js0Cl/P3fOUaRHYBWJ7mt8Jcnqkvv/93gk7hLkU2++gJevFx
ezwSHz9tNjdLuPA+jIelHLYJOmK8r3XPKJ+DE3TdaaBK+RDwZ9yKebnvJL1BHWthWrwIQk1I2Drc
eTBSEhX/+nwcIW3TWCiqwJTvL8p0kSS6JQOdC/489dztw6Y+nDP0bZMEumg9Uj4DrfAurOuO29fw
0/ft5oSzLfSV4DDFZOQyvD/aXKQ7TtYHfATRwMtKPrjkZExQw5Ol+qZyKlv+VPNn0s3Vr8v+VuXh
PXtKkZs/FObBM5589BsbiagkPg0WRT06D68gm5XHlilpoKpWyvUi2bMH67qsfxUcyB1O8bOPaYa2
CeQsOnfZFVhQpm12NGewwh7LNfemOtFaB5afDEnj+BDUSbr3D5BCIk1gbYZBEBeuYJlTiMzbIpIN
W8Ka5sslw4Fy2NWOIo62Jd2TdUwsmoDL2cuW535PZ4s1TiY02idcA999AulZZNR5lfR+xujh3vXd
HvPnzbr0/thmwYM7lXu3sAF33Q1Sh6PPLZrU6kqOJ4/LaXJy+FEiDzbuJZm+mxIGhj02xoA58x/j
vEa5/9pL/krz9g5pUsVVke4mlk3924/8D6a2WEx93oKuG/YJ00miSiJOQQvaOfP7Ge5MLeL6tSt3
FKlrIQXc3DBOYhZAGCBvR/NvAA5ic45ZSjpSJqif5znCoCaWxKOcftkE134pismP7R+jiLtQGe2M
/i8XJu7T/nrZo14v8y55CrzefrCvETl94n+uamMY6hPbhPefSGK4j/hXoxmvmywOEMhMIjlN1v3B
nPQlvaBJhx57E6ip/GCMzPMw80ZbDpMvkgvirGfEcBl5O1U3DkblMwMaq06T6R4uJW2Ruo1bp9E0
F6BuXNZnkaaJGMWrhkAl2uFeVuYciltLVWY3MFchxejLl8p4qVgM4uVkH5B011rWfU2Fwq/VQnhA
ec7iU19gjJRjtnDxSp6izENLUBokq+PE5mr0t54slIkTdqGI37I3KQNcMhnYiJmr8Ee5O/jHDlFx
5upjyMVy9FhsnowOIWFGFxXsbrJjplklFJP3wazWupNmYsu96Y36W+mg9t6Z2QfFXxKsENOqlNmF
UYe98TrvQCZzrYjKBJtben9cN4Sl/5dv/ErdGM4s4bpI+SoflYo/0hWqs3WCKnEXkz81hXlPhdcm
fXmGxldG2RKJRoxxAdmPaTZHmng8ANtR+cNBQpm6m0EH7Tw8teLG/lwDjDG51uOh3JndQJlOTtkn
u/qVG6US3V07Ohs2rfel+DhwTqzEG/J1Mlcym5/bF9Q6JVl3Xj0H5wdUWHjlYrX6tQmF58ILNpcu
bjWZmokVRmfD26jCDP5V4o/w/VUw6ypDDCSeXs6hqjq2ybYUJLCe5n88dxtK0ztw0/a27xj3pKvS
ocBzWKkmJCJUrCSFwisnurJgVSOHeOvRQjJfXQnTEITzD6ENpIyztzJCHWQemHbhO/nbq2fyEu2S
6o0Y9R+nx7s5Uv4goRDbVVWi1xTxGR4Og1+m685U2taTrVZ5CO/PhK3UhCcj2VNeHrNvy1/dclfp
a9v2UR2XAZl0BTe/liOFsaTG2kz193a7pcsDZ7dti5Cy9d5FSijxocc14U7JtHHQp+Evi8cUcI3H
pbkAMkM+4HL5cgavyrHCq54UXVhU2AirO/ne2yAjwAmSbUDOP8G/7eHi0aUl5l9D5MHnVruCsGKT
OJTLB9i0bH7pybtF9u5mxheIKvV6i2qSpO5em3naFHOuJGyqBWYPe8KrzZXeY+F4cwSR+Gp6WhZh
UAEE2sEugI8dCBDyDfB7cElJSXcNsdZRDARc3H8x7hj9IP0J32aQocdgAro/SHLUkFVDtkehJict
RCsIM9ZHnowMsNweRsUMSYylRuiWIQSovKVgfYBFa3ssFos5IX4pXjvUQnmdYDT/hUB+a+IgQeQ6
F5ioD7Rvm9XoI+pGMxMQr457Km0Uz7PyMe3nFWmQiZh+g5sxJsCDYe/e2frwYODjeKCd7zw6NMRJ
UgPVFHE2MVoFgxMCFs4JP02fQjS86Puadp+IwcI2z0wVpdhiuKZNDWMBsDrPz58XJpNq9nN0HOP0
zpTGswgfnWwK69mdb2fIU9z4iiZOc2Yd8SXdRdPK5mtxwmYvDTY48OyWthYH1iKjDajS/wOGnmBI
dNhLY3lrn9jF/TbhiwIfynrd70eGMjD1ImnS+F0GmD95jiWxmHesT0VFmordwe63W9ocsyTxi9V9
IGZ+fpQ1otwh/YvAQdgyuIUG9XQQVmGu86jPbfLQ2NtaL8GM45Ho95em40kPylxhhuOCv7YdzOHk
nZkFXJEiwmeA2tOXbgiMf3691cIfG8ZCpPU9NaV5oQjhBPNbVS9YgCGFkiULqkUVocD2TiVYrJfw
bJfSQY1FSNV3O6jli0kQHK6T6n3vuSq/M9FRT5hneadHJZ5WRgFLLZY/2APq78Kj9Xz2Ox0HRNMV
RepVS5OBDKQs6r3ViTE1JDt5gx574V/sL2r6M/l1ni8i7F/ADe4eWdJpHnUvFsDKqRhH9MAlNenO
+1FWbDdVOFCYRq/OU/IWO+3EFROUNA2Q1t6cQAJvYoUPk0S52U1nlOarvjJNMyxnr4cd/8ltS1ZQ
8+IIQXvSGP0vDIG6mmWBxBw5d4CsCkqH7iq7ytnAb0V9Z3g1h8Hx9cy590TF+JAgmkdz/a094VGn
m1ksngvYPiXp0P30adnlnQFQV8/SfJo1t6ThdOX1Zvp9/XREgETf4etdB2JTJZPxwydzjHXALdFa
S5WHB/g71mKDAG7et9FkHLm4hSELud16lh1ungtTPpydmUezApTKo+Mz7PT8aGoRMcrJcrE/8t4D
8NDNIF6Q3SCzTcFo8XIMj9kChIe2xl0c8aTzQoWea8IoDwa60kE6sapfTaIaBxPsZOQ/5a+MBImo
HmY+90iLEGD3XtRKHRTetXEi15TQzLPfohmIBm1wcaZJRoa+ACHHyAdOiollJJl/7esGMBp9aW2g
eayUuyuVKWSNp0wI6mRvxe2LG9Va0z1k285IoHThZEnkbyTcvNKvv9uv7irXIrr3dScMwP6p8SIm
QeBsnBIw40hYFhT1qqzKIyNguyXpx+zOOUKE5llV/Rax/XOnVCYhBIL7WUFdGfKPwdLI/8rrB47h
+jDJqcZTp4wJzMozbvoBd76VZKHZxD4cREQXfjSpCHFUPY1utLhaRIqmKfk03kYFJAkcDcAZJFcj
nDw1a/oPV3X54Xbm6SI6LrqJkKl3+XoECiwa2wnJwM3QFhX0ujUlFYBRoMBxwD9fNxGSAIMiwrpN
KFlJx0wwyyy7uBjxCivoM5vUH3NzXfrwdJnGQf9El8PCuHN1aasCYL2mlFFiinEPrwfKt+z3QrhD
w+iMcDcZCHGWkQF4rWfcn88AmQZGmRBkRK3ShjYIIP0rgGd0uiKqGwMvHz3NgRScgH36N89U58et
hYuGS3XtrSpZLBRQanqtegdQtKhOw7UPE5dAl6Z+5PPsEHIY4YWqkzBbJXEn3ZDKHuPKkD16/yE6
+YuNpgwVnaW1xtxnDqi1d5kBTJ6GA0hyTn720iKQYm3C7N9ZFwHZU1VvRln7Vr61lZhg/PZ/ZcFo
vusWDuN9sEU9DYmlS49Msl1XOjahutLDfe85XsaEH0XYorfql2Jv6rSwSvFw2zwMpV9CzxOY0+dr
C3YUKkoHwRc3nHadn9OygkFQc7Xd3gN/laYiZEnWtqB/uMKn0C8qXrVnEgy9w8mgdb1dl7e6DL8h
NI0sB/4OxoptpIAJrRGXu8dG92nktkmEEMVFbBjyQBH3txZYtbx4rDspE5aIZaV+fltY2ntDNLTd
6xt2Q2MpDFnuqGQQAOojT+C2+gAiqBM+ebW04OAo5yPH9tE2IZaJQvQtsCqA2quRUnnEafHQFXpp
L2A2jmNmHO00QLPdFfwIJsMFeF3eWXk6a1u6Jj7htPgIUxohyPnF3Dq2QsMFQdQ6TeAZGC38T/hq
RuW+5be0Qtq3Uhf5FKOMDCJ5haICAHqcTKBbQ1KpBP0aok5UBip0PKcK2P9vZ8Y4nbpr/MCfhEjv
eTQ=
`protect end_protected

