

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
aCDLXtVrULWJvV+ER7T5zOiyyIpooXEDGQ31qY2Gso7MygDjVHK1QZMmLZ2ktJwbwa+ZwfV8CEox
1N2CBFa/uw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZHaI03S6AJ5DAkcQ8Qa5VLNoTA73wS5g+J+D4nyvJh66O+vaV9OmiHTbJMZCKN26yj30r7urlL+O
o7Ne3QEdHhR6EVtEZhL9fX06u1GwvUeYLPmTw/BJdHyKgDmd+9C4+DxNXSxnv1FW6XBREzTyHRif
D8Dh5qWHw6ZRpCZoQLQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Hz0NvGkQAzZh8jguIKoDqgUfWtUuXP9xr3NKkeIoOA4Y5NTp4KNH1olKBiZZh7DkBTNhKiX1J++r
OYmUo4nfRKfU8fGiMGkBx5TFNnlCwgxSAcfZw3KvE38bCseRSBw8AjjY7htrZPRaIppOfcmLU2pH
UIhN6Y8n0QUDiZpTaArLhTZtihGwO4cK+ZUUAPN63xhYEoc8FWLz1LcLQtUT+72HxnT8C5l7nvyL
qbhvUrc9WgaMOxVIHNIt8ah/LvHEQFjc2DVoeMo5ZF+V7JGYiyLSKWboEByyGPXcBI0V9MuMKeFe
CFbNZ91ovnfO/L0GOw9BVpzYS+jnTGLx9iA/Zg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Dqd1vX03WX72jg8g21dMBfn37fglj9IcNuGCtS/BkF+fVt2DC67gTDXpb5UvWRHGxYhjhAyFngv4
f+/cUqiFehoWkynFGfbw9HsLRSVwsSFST7+YShYHL4gSqXQc4T+9w8USxr3YxXzjpCbADPhP8F20
bitJur5ELvsZC7EWlfw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BkipnOWyv43QAd3KdHQpXHtHFLb3FIa8QngJvXphENRJl73YeC3wDgRiCndqpXatmfMYIL6/fo5n
6WIvbkJKl/doLyJEo8If1jB2qbpz5mGEHOh+uJwibPVN5CSP7LtYj4BsT3IyCaCsb/DUk5si8ays
jAXr+m6ka+gVz8P2lmx6BYKpTDV68Obl0j1Vadi89hYJJ893Tuq2EN4DigIzFUE7GB6Ta0pow3V6
jQ+ZiK4tHjkMrJyXG8fdIqo1Sr8nBWCnLygUJb/t2P61L7aUReGH2YBSQlw7/n52QQMH9c0SaHHE
Nj+KGtPFq9CWw229xQZsFzGM3FBamycIpVPXnQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VCYGICqcGstADU8xhghKf0/3vDYSjwwJngUAuvhKrcJl67mSfB9uJAW1UOqoWcHqUMwRW100Dqkh
Sv2H30f2aHqb0v05G7EABv+VlUdaN5oSi3+XWfEueT+RN2mCVNEfd2w7rc4VwtBqe63LVcVwpCmo
5nAU7LFH9ECIewkiC+/XB5BRTlI5qXAYREoMiVT+2L6accCgRTiRc1vzp1sx4F/uqeYfwUwd4rTK
Q0Yjg97+as+IU7Xyb9QXlZtka7M1hfOZT8KelsEfdTTs8kKWyfo8R/o7HeXhy3mh3xlD6H2QT5nD
98uuFaFZJLpfmHq8XK8qdO1HqdSCgHqm1a1lpw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 112432)
`protect data_block
5PQZjeOwY7ePjBAw/FuL58wEUkRb6GAFRV5J6agVwLb92l4kKJflKZ5DdYeBIU0eEF068JY5kCnO
UWcYBuv6PS7H/2WxEg0UwQeGyRmpFQMA+zWAefz1KCKDn6kywbrLiqFWPcSVEcU9mvoWJjf55yQB
qkWATuzPZL6FfHPKpslIwx7B632qSiMNkP8nK8hrW2iSx4Z1pWq9UIOu5m52WqZsCX0VQGmY9Omu
+w1nATsAbbS3ITeGc+l7GZfmu6dPeUl3M5OH82R9BF3+2rr/R0zKP/g2MLaHETTlTV15nV4GRRKx
FB7q6mIE4YP+uUQJzpTbo3Q2TsZNm6/u90Covp5a+VI8AKz+4XXVlRNq5L2B0GRIxGrh1YuSAfEs
XX79/q/SM8+5+OhQ2AxORbnNvJs6ZDw6TruZzaYHqzH37isCua8bvsOLXu5yOC831uZgV5y28TtJ
YY0zpKpQQ9nyoe3AxolRGP+3Z2AzbgwEAb6RPBXtd0/xYO8Lsdr+MjZOP/9rzqg2172x+qxGqy6u
WHsdS9ELkBG0YNmBqoIZ+Ua7ftq9Ec0AYUwaOW60YXGtgHkPVvoUHE+DK3ZGPwf5utSXQ6zXG7I4
eHXOgX208k2ufVkYE/fVVzj+RdwijH7qOGlKZNXiV6L7j3U4ehCJShqMXQRiOYm35VKm9jgQ6nce
pN0M8L7WEeMzwBx0O/GfApc12uULctSqEVkUfpD9Y8CWZebyHOSHbUXqi/eaDnlOd5kExK1kwqZT
lXaZo1iCKg0y0pX0Yy43m8GicnEHDEXH75fVldqPZ8HBMhhY94RWnCVRGyBaAcrJCeqfyK5+HxXx
BO/JjjIHSNuOn8gAoz1bdnTwYTJEiBSsnUrcz8bYb6EdpTSGnGrLpgAG22mOK7pU/OAzPFBI2ILB
WJ0+ok/w+QQOe+dy+XDagS1KJLAQ6mg8KoGSephI46hbTCljDOpEsEbUfjPC0UKM9yh4370eKJE2
yiuMtf8EaFjNruH42E2rXs4INjcdzs09tPYCKHxIsXmhZ3B2p1S35KnjSVsn4cG70ufMY9/cRh0N
U0xc66drJlQ2kgbXcxJVhuzaGuQKRXXo3q7iAykuhLAV2i92rdHg7Dax7aSdPrPhudoxdDfdEh2/
ABPYyJlBTwoOSE6LPJb3olCWzLtaXajahAKrhlWKzFozgPbg5JP3W3KXIjoSnRcz0r/w9g/74Rip
HD5l4/GARJSiwIdVJWr28oMAH9ifuQuTkBAItbr3sO1b4KiUVIGE3FNa3WjLP2DG+fw3ECrr/fnr
DhBFnyQNyosu2EH1OkITy3M07lS+tz48VmDPs3+Yew+oi2vyPYf0A+yR8rO9vOioS8Qb7KXvv/fJ
lRB0fJCHiRzkHl3G9F6576H/AO4XkyNV8+1uDI9+Wo16H/UU9ikBWTuc6YgeIaGBJeA3aqiBPjfY
leeYpRjt/PlhiFxaK6DmJHWiVljfjXJj4otje38RtwStVfDc13MLH+u5BWOfaZJuSzSgSe3RhJd5
h7aFkd/NDK9EdcN4oUDNXkf1gFA8Wu2wCOHVx7hp9dIabZjCGeI2ylA7KRLehDg0oA0hv9g3hrG5
YGx5Vr6UwWsK4APXzOPHl7s/JsBjAmSluFGX1XsGU+KxAa3/1SM8cVZH12Pn1IbN4fEWzWBFkSML
YiP0bdEPTLvlr08uChDFvo4zWjs84Mx/DrbkQbUhLry2IeM06gu93aPhSS82CQPZybr/Me8zm5Kn
DZXbzxvGIbaloR1OQh0LpZ27CC5HAHHqXcb6ebec+6x2EpKhjbwOpzVTjmfesJ3Epo8Z1CcpRJBf
26xq0xC5+jMC/QQIDLsaPgqHI18jfBYOfbE7uae+4JjUa0hiEJAK3m6kBhwWr1X7BsP0iZKCA3Ai
PiK78DXBJGsRL+ok6egOS2o4zRDsU0ZmN0br8EduHetBlPoUG8bQyin66cM6RYlqM1nH56uWc5/p
Uv7E9Ycg5zOOnt+F1l8BoY9ZQCRQ83nOVXlpeXOO2dW07Hh7+d4QtBGvM+cBTA0oor/BJxbW/0Ks
LFOm5dZlRNwqz4ftHJ9PvcTdiR00vFIwSQvykX9NU38KRaiIwpV7UX5OjHNcuy8iRWRTPlt8NPDw
lrkQGKMaHwUhkFLPRmkJfNxOEKzU5l41rqnH66Uj92IV/YoOeyEhR+gWpqJT1GocUwH2bynxBGy1
Txqf6EAN5OqqO0AarehqRZ0yFZw1B1CKsWGQ9Rp7Sb1FMFCVNKut1M+rgViL5QsyrbzpRUQ37Pf2
j/xyDwVHD769plFNHe8TY0vIbLREa+qVm6DNCRDGRAL4Qrxt+JLlFyJaw2F6DuDADl/jTaOwUqRL
SU5g+dR4x4oEeP0h+slSIH3uhgG/EjM1p1CvRVGffgc0uo1X67+K1kyCthQi7lu1VeokevJt49FL
dP4e2/DC6zS8ScQqVYrOIGN4k/lKTrFqTk9x1btT9BVKdclpt1kLrE780yZbNMHJDLkkUVDn+pDr
oAvdgeVK9fnzRPijPdFgcmBvAAs2il4Ts/LsWjFE6CYsMVJuPIvnsEwPTDoaCg0+LaUyCoEYoqnZ
gRBGLMnvQcbxihjrYrvqJS2WqCeCpz0iNnWQBrz4d1xShP1KD3W50M70RG9Y7ipv8AxHW09pcdah
Y+6OPi2kHYYL/p53mzO/+0Et0yKrxdptqoVqRM+6I33jy2UtdQf83c3e6i6M634rYW4FsB5C/jb4
fIo/XEOioW2vV0lhfe3oGQbBQ2FlcELzMDzUYZ2nzMOTLVORso3vcTm18tit2jfJbWxTyCKfYP8i
gQDSqKutdagvfMuHFFj9KzF73oZ+93ZhPV9X5E65/DM/xBl2mwydDzmAMFrlbs0kKBrI53e8nWd8
jSr4sDp3Wl/wqePuoTSSAgrQM8b4eSV+yUvX993iFgP/02qY1knEep6kjB9hHiiBEtQFiLt5y2dl
UJAAOjBeXKCSBoVMqwqUBj8mf2TY4/vYbtBCbOeMbTUwEqp0LkS6F6juzwPoZ1dPnUNIkMVq/ueB
02IZIRb4XPYYIG2H4wF2tuDbojuIGZPL+mmUsZcSOEXKx2LO/C0Fl3tThgwaLY2gWlckzUHRavid
1vpG4QJQDX+n94LX+paet+O95c0Fl0dLKMDpPuGG19clmmESbx6ohG1NVOaHZ0FTFSHVdbc3aBK9
u1m8UopfMtObe9ntbmgTh/ilEpyb1JO7UXiOP9h3kMWx0/NOrFAMU2++SrIcRi6wDL6EA2w+H/8c
yCrp7w3D6sGl6nFet22GjKmxzCWZ4EyoaA1gZ6gHbLNVVIlW91JrHpsIC09ISdIr5J8gj27FFKEA
zBZDs6rohgxldGHreo3fZiCOcCS2g4gXvzCLouKmaXZz2Ui/1Tz/Xr29dJQLApjR1frdP4Bd6pz0
gYARh73qYw6wseR8nuuUKry5W55r2szGwGDxh6s1L+cTt28n2n0Wz/u7M85nbwho7JFbaWzXXmDq
ZMIjeoaf8fIrqqIc/LClv2myLkquS5bPKtEwBTi3zNL0KNFelu5DdnvszjHFCf2U7Nn9bmj0n+An
WAaf7y27vDDVDWZITZIRmAxcrUwo5GQaM8HB+jWeOwiWTxQ8fR/lQGRrXgTYkow5lYG1aWqkkWM2
nMyWBg2MKJYcVRoYBOz9PfuYzFl3OE+jCTNVXrJ2x28MqDNJoSfbh5QX5T4kQI8t8HdOKoQ3pMzp
i1IU1l4qsbMKRY6T0kmiDJz1XVi91UCxa61HK0lSxrNrO22XzpR77XMpnjms9zIIVYtSQdPtpRk4
vfgJH9akx+lBxf959Q26813uabaleY2WchrVT39f0d5CH6aHNFoy7vb6uSFDA1IPFSRuRYdxpOZX
jfRTaDuyBrkdjpowWQXMFEZ22W4N4EqwSebIQdlDZSjjmqR0NBOlItblfcuBV7RniD9gwSueUaZW
+tDcTan5c0gdNONRqivVfhcsntd6SsgbQhi2kA4Un6874bUrFawqX/Is1lWroFGWAdoCxqUuZUaR
jmw6KYMax97PgAsSQC3a/VEc6cTra1Ov+Kp+5JvXEJSMD6brXY5Y3GEXhe1jZt4qFYjD6tdvjgQL
5bMgzZYPbyxz08MZF/+eaK3eW0M1P4HsKT0KQvbCbZgLSsFYUU8162BRWoCj6gj3svi8yuCFoD5x
QBZOJCQvB81e5Z1UUpC3z2N4Cy2CdUgQHCCEgS+Q7CKZEB4b1koGLKYfZlWWf84G5or4Jz9ooEo1
P8am5CMJMMJBWG16yaeRw+NxEfKMxKxJKOp2Px/dFaf5QW6nm79Jl5CiSr8PvSh8X90DhRk2RiVU
Oqe0ts2q2ZQEB78dSyShUn06zzcWHGLieMvelOnzCmcbekzodp2V1JkaFanFcmiSiubs/P+6f1ay
IYJ//wutZ97SDbXYvwzWEN7+p1qSoR6SmCYYw8sSVBnBVIM9rtE+v2cUgwQGqv220h7YATUzFXZr
EPlQZvtyDiJvtR0qMTZRhfX67XKWWCoseV8/70oOt0OchvO9yQYaq1LblRpPnYwkEgwKt2f6BrRP
qBquknNdjlCSKx8QPbEAWYBj5cgGI8r5ZcSLk6/O05rgiRLu8CStQ1V3mT4v4wtTYm+umzZXUdAh
2reFcfkyck6f0+4IFQMCXmG3L3OO9B6ckrOYN2186axhfJ1GoqNdZ9VPvNNKBFVhdTaqTbiRXwRf
tN72UAYe9vH5kLCDuH1BKE+mR1y7WeTU1xeF4fC2qwO+3sferG2gs63wlQrhxrgh/bGT7ujaTXJL
WOSyHCBQcLl3z6XjizeQkpTKMH8JkIKfCfqDVMToClZuJbYWgIiI4ibJhbARKiaOYLkMV73jmcO9
Pjr17ZFlyS+R8YqlVwDw11wNaJknqq3t02opsDM4ZCs+ymoYeFVYLI4ljr59mtCsgPmtC+98/zA8
LOCZVZh02Pbx/7MIEoYqWSyDooUPyu0XyXfevpFu/6cLXwyQr2QBTCVO6wKE6x2oIe4Pu4Wf5331
Spp7Ru6CdbgzVR8YZ2ciHnb7NPh+yVjNBGIGy0bjXqLDakE8t5Iozxapq/jt5E3sUqBwiOadWUYj
GN25fZqnlQ+Lt58hA+bpE+yLDe0g41oFdTdWXA7KyMmMyntscxU+Ma+Kk2noUnI94iSF+w7VEI/i
C2GAZeYPPSl+MJ+hTkVFFhxtTTTa+HsjLU1BVo/hfcafGNw++F8613Xl2bQ1OZXcsPLmwstXtBVW
vfmI+xHPQDUG1D/pWQ/d0AAnYefidO71AbZ6ABUV3F27vXmqKYMSHvDz/JzvQumlJco5NC3yWopV
sf6s1ezMfViQrM8bvZ5vwhHX90F6alFTz4SIEv7ljZeuq7YMR/xARwvaHXP68QZ0ez8QS0rqwIgT
sRjGtASXyy6CcAzNfXaXOiNOuEK4Z+IttJ+7jWl5QaYoSls1m5HMdq+d+87Ss3QVnUD/qQixVlSQ
g3RezSVaLQZJ9KCe+Zk1czah1/u1JHiP7OMhXcVt3OIHzvdnUZt7xeIb/eZ5o3FCahT1T9fi9SsE
yswYTFSRCHtn0NPcN9GRKnFue9LUBJ2KPwKErVrUpoC805YBiwP8iqpjShMDgaHK70ldxICAqjtt
Htt6GjCCDH4ADErvss2cN2S9kpsyYc1CWLnTrbMp3Pe121qKKeRyA7/5+hSoDVStQ1+qyCkSpRrV
eToQGntIK2QJ8uCEEQtNIyLHUjuaLnZKPEuje+y8cvjJ7H0DuRgKOzcvRES7aMVr+NB2S+eh3Q4k
5lIT9uRn6Wjt5bcXb32bZm7OrayDM2k70oQFP5jJmz1LgmQiK17NXDu9RjjvoMEAImcktj74Aq/i
rQ8JshMb3alABofLlrBBzH7aCRfCQ4gOu5Cv+07kL2RAcpHlS3xDc1DJYOGVjyC9gWBNVgP3N6bU
OwJjuNDFQIUlewryKy4s9I/WzoiTPZVlOJf6yoscCNFQX9+mk4/XTNV+3jr+c0JUT9y11XZKqsvV
YXYa6FYjs7pSM4EpAmqcHucVV348ba3RitZCBFZORrFcvgklsUiNK0EwMx4EZSmCwFD+2WRdjg6/
YPVJ71Gm7+OQTeTyoQJnAvNlkYd2svplPVL6eczFoRROtzCT5Qs71JD45WIj2VZaVsHJjoH/4gaF
FVO0PCryAODjDACeuK12lVHyQlr5yZdYW1BAa3QQ1+gc9+Zvbxvh4BLcHBgE/MgNcYRq2jwPEHFs
vJKtScAse6O+xz2KDtaSgqB3dN4+GpP0RY358O4MXGq4Pmyewp3A3W71QuorqA+Ay+H8X0wP4Qbd
T6ATemxZoaxWHSmpbG3xEiPrTtGb5ZpS6bu+XEVLOpCgj6XCQYGZiMBvnDBZ1tMBuzq2rACq41EC
X4yg0M7RLj+83JfppQPdz5BvPo/huS3+CwcGfItlE78fyWF5FNuaTF3As9JGCEimtwvUkML0/pQV
GePeoMX2BsE5YmfVe1FH8CD46MclYQjkfcskQKeoZ14g6fGW28vTVZp+jV2qVDLlR6E1dHdqzGcZ
bJf+HTxnXjebm2nD4lQLF/SD0qwQvfoYJLeADcrSH3L4j9ccDl3cryX9WDzN4KcM3394v6OBwOlf
9bhEpQKQQ1hC8XVOX92+q7f+BBlBviFM/g0v0u8icb/Bz+H+NygzJOKHrfB3jZYuko/l5ZW1QBLY
rK6uxDw88SyQP4FwryxStcPdReIUvIviE7Omi7nbLdzP4d6wfK3cLb/mgUNqTxeWiJdgwaYKC6KW
OXdgeM4NiZrsZg5j8tQ3cmDOpouCwuOU94Mpxb4Wr8Wh1xfg0hF8UJgpAGGsPg2bsEPRqz945i4c
6AdV5LzeKH7YWnA7b+wtrKxSCdAMl5I21ccxTLzh1tzalcavUQGGfUBflucLiG2w59ULGqzdUvv5
dKfDRa2GmGkFcfQVijnSyfaWpEXVrGfrytc0i9luUmCQ1ljIcEMUwNTrr+4HtidmfATBrqdC4V8r
dgXjV1ui/yAEffOnUnZdoJkc5EhKbOTaEBODSV/3rHgsU34Q3AQz4D5hKV8mp/XzBp+ORgUTytXc
2MndsPxoyuTh0I0hDRsuUrVwrnuB5evINEAV2WjsjkvunQ4DoCq+Ner3JyqHtWG+PwBOpjK0NgvS
q0EIIM1v6S+PRoyLdyUKbjaXeAfONOOXNOgLWDjwW1Up0I3otHyq7fwaCT8uEqKRXc3fcRhWaAT2
0CrDgyUBB632ejjeVSfhzwNXnF8XFsia/q/UJUvDgi7CXoF7R4qw9SG1sXofd3pHo3WXRoPZc6rB
TLPKM4jG9znuVXvy0MMKryhU4gy1d3gMDiX8q0h7gD0IsSrAj80oDqWi5Kji8vQU4CQmQgRoNvcW
LjQlAj8Xkdu+LDrIDhxLyWmSqyYlPMO9fRIJ503kJCykU5imIRiMx/1r3mcNGVQnzR6V6Iyh3BCM
t9zYriwzFlmNJYyMcgFVdTT5m5Ehe9eNdPJlqNfT16BSo4ojdBFqsFw/B531akzU+RtQGU0lE/aA
qCpPpi8jnhlLjX0kDLtfI5b5BigN1pZvllg1Wwi79e5AgRjMCys6jcoxhcAzIqX17s7qwPX/KCFZ
rOLQ9SAreceH7fOPQuJ5umYEhWK8VWOILr78Bw2N5ojoLUVjp9DS7TOdNQ17cYOSXXSLJkINcPJO
/xC3ZDxuAhxjg9d4prt9xf9T78vj3XKEFqQF5rA7D/rUvMn5R2AzMW87xwfrevzVISw2L9HGu77Y
tTWhPmkO5mDO0U3HzbzzkiAMvuk7tXC4+GvfCJLmiWOYzlqq5vy+1vS8Ls4W2PwqMPHj2nOvGB7J
AuXvKz+bntShZppdS3PV0pznsQ43vKaH1Xn30xDHhoND5sTH8LDZBvMu096Va+IGfxYTvTifs06T
562HDF8UrYJ8OyXKbwclNp+NTyM0DlXRUunZqwxBKcVRmbgoC8tg+ka2sbf7nKwYR5Baiw91FL4A
eSNOahDIP7pw54yt1oaIgetfaYKVZpoDZrNRVGxzOkPXwvMTvvRhO+e2xS9BJfx3HMhVvZWYRo9z
4OGtkcRP3T7MoKOHVGERvLaCiqAjP++Dt8THYW6IRFy7OhsYkUF2CJ8PFS5gZz1AsC4Q3JDzveEj
EjusHihvJp87KtaksO2seHaeaBQU5RRlPNQH8/ktxqDKM8dfiISpsOJCgPbt/DJUYTJoMqJbplI1
A33QpQ/C2vUTK4DQHVx4XsfzqbDoinCKmlR9lEaLrTZZ1ARI1dv6720fTZ7jXg1Sfu83QCf4t63S
b7IBBHZ4e48hW6HDX5MKIJe+ufkwjlXtxVBKHQraJkxSVZbvCDq514KNWv/W1houpp7N36kAoe2f
R2Y8B2eNNChOUGOHEIUE3/9PVJ5MJbZ/vONKx2kH9IrDC8YaUSkurXwg7bfgWAXriCumu21CemFY
yEHrZFLdyjGCXGUIP8CWx73T34Wc9Y5YuChMfDGgvTLJK151+Dd1Oh04GVt+PLPge23MPl/mx8l5
GDMqtOiWHomgjdeACUWLh7LRuCCQWVZgCb3fSSvMhkZ5nFTgW5wWeKmvgvsvlp6tQA1DspUsLNZp
cGNy/XrxD/bNTOOaWkW81ZsRCzVDj/pzYkYa8u4yrQJKr1OK7osdjXnNV182Ue6k4CGi8iPic7Nf
MI+njRZS5hf99TTvHeKE25cM3d86FrHmQ3T3O8NAL35hRsNuPnMaFX2QwgBfnqH+yHFAIz5nKcQt
z4j//mKKCfXYu2fGaX5zA2JQn7iMSruw+VGmtoZRpLuPvzLY6wHD/s2v69JcwcedUHHB6aAKg/zQ
NqBiOGwW4KfCZ+YjSV9ChdiUK8ypxwbchbGfif11OSklGu6PJExr18fcKAvO/AfRacBJ0p+QnwDd
vOIi+geRfHVjzaz9bTgV2ze8h6KNqRGyGZgVWV84gHeUe6dOWnOqBqgaDj97W+FCYSBpZJItAlMU
npMuWGjSIr1whsGm7Ygfi7B0owtPJjc5rH9uTj70w6n4qtGLsLaKFbZKB8TP97qDCtntiOzi+KAS
NJj+Fkp5fdlEMxNBTIFPweOI7h9eAMLpDAD3hr821G4oHjYS9XJUG+B353ibaiEkdbDbhdNTygiG
D0Iq+2i4TGg5X9UaUlCqcBJ9sjoQZNawmFJLF9yVlaLq7YsakVnOie2dPvt5MkagUiY0jMO8YwEc
cn1ECoSv8pFemkBenzZd1h6DK+HCYO+Symun3rLQzBOaW2Yk6BYO19AKMBZIJRbc/EcQqh758xhl
3unFXelWHHBYze2MaZzgt6NmL9FanrPuYQoKdOYaj2xHIgJbpmMeHXjBFDYPljYzueVgN3JF9NO7
x9C3vWIAV9MwkS5lWYZ22OGeSgRBVnDD+VDXgEycb21B4JFioSOyn/fgX+C0+nkDL2b9FLOPJYjR
imtBDlWzeq9+U6DtvkuLL09EFaKF2KKpLLW6M6yVZi0qgGEewBpoKDh5/lbpCOwmKeo36KCpIScM
MNvhoMr7B56klSoTM/X45WQf7G/7ULsjO/UzU307uOQn3g3Fc1IjqWPYm7ag1I2C6KBGlIqgvrKP
wnIfh8U32GT/I8KPwVPDYF5P1t1DaK/fNWGJhiC6JfCXm+7UYd2pop7tuV/RciodNJjW1oBufEKt
d0QWFiHeRuZVZtRNoQmDa8YKS6fECL+2MT7ZmF6xSokYhVAb+XqcCOCAtE5EC9IgTe31nm+WePx5
i5RyGcLqGZru2iidCMrAlavxbt3K+iRDPbrAB4NHQp4X8bvQek+ExAVXeDd/LSRJcuUAQnXV6f5i
MaAjFU5tkX+btyhUQmDmI/WVlIcY+SDw1mqnBfQJPHlHECPhDR/hcZMahaBjgqPzKqmgPvmGKLZz
emCp5vmQOfPU2sveTAaJyhGqSNIMW8RkuUiSlhCHEoFXxcQi/+WXkg/yxEbN0QpsEG5GApxkB46w
KgprUXY9GvCA3iYqrguPwhUwHFRTysrl1KZNNN4+nhNMsywi9mNZ6KQMXdHSq+dqupy2JzHzvvsI
z4MypMGUjoXEGRHhfH9HIud6s7Dz2o9ZfjtiYQ48tL/pLJnIR39j7I1VggDDXLQDEBfLKQTSrIKD
m7EwE+7FlVLRmzFxoKsIau+TiGDep/8+TyIW5ADTw4pCCJC2k4loGzp8HgjOOSQciaxKWd8fTsuS
DVTLDG4o4k5/MKk1FxVNJD1v5QhOvTCtwf5tr0nHQbq/XHD+1WA/zRAa4ArL0sLiG0xzAKP6YRZw
/wLOtATIPMCN3x+6oAfpvNGT5EZRfA2Id0s4lQVpbghgAIdqn+ue+Jrn42aHXETt/1jdMhNttb6I
kA3q3HZ5iiopN3Dcp792oAvUGUtHWZGXS4T9ruEDRQv1sYZcYTMw9M+Cz1HJvN7pRMzq+GQ3rsiP
ZNey6cDgREWu6wjXdS+9v9nvIdtP0elBY3adSVfJLKM1QxyP+4/QmiZeDxvO31yoHfgghv1rqu7J
gyTcr1L/0W0SR3FaIJKsyZIwgDxvKgzrH70Rmj2TiR0mgfUrt6ZyeLGcx0tdRNd5bsLKnqVucACy
/SydiOli+nvuW326MeR7JdVbkKfAXE9fitgSELQ0N7dQIqfnwH25lMrLqXlDUdDRuolEmVN3eIx8
USY7+xs7y2S6kUn/G7tY/4VtlW9MOVkqp9DYbnUkhkIrFvgmTmm4lNJYiI7KQke3Cajtp5AMgL5Z
X8+Xc/decAXT+Cco2APYTk4uWXfjwFis2S+yd+PXkbR0JaBOGDiL3kANR2TbpGOGKoN8T8Pcy0kf
yPhuKmNpx2NPTC6p5Y/4H81zNFqsiChg3EwECv0bfoBUYPEg6ILvZvDd2H5Fl7VBjSC9b5cTyK1b
KEp07RLDY1gZCTt3cOPG//QOrjdmYKkpe6dCeulknRnbifuhgeODupLtbBM7yzqkvln+rvOW6ePW
YHcFFN5gkMSMfnSRyLD0nuHYmFHd3vjmpPhELHbBp68MY2M3TT4E1goehUoo2+suBaRk3x8LjsQU
UFNVKOUhkVkYarAjLxUp8iFfAMOrBwYk+g+r73eR032LtPgp8D7bQHkoiWUXZyB9b+9qTov9o3+A
qSvRdlRiFOylYEkOXokXarXP3MPVKQuvImfn8AVueKkzj0AUYKW4DNf2t9fLfwYZN86BVtJD4Qzt
NAMxw0vgKwnwutAPPkN3P86f5CU0shpdA8Rlt+NIP3z+mnk18+vzaGziC24M0vODSLMvElS4ZzPw
fSq28qwNhQ/+yQbUkrgqWNbX7hZ+zDn+7qnf6z/Qbcx8XBbvbg5OwSJQgdzOq7gCFem8y7CW4yhN
hSco38/AgD1XuqlkuCACuVeoQUKeta8jc8LFPwMFzh20HwfAI3jbqPv0tJ/DVBjw/gZ466MOhDNt
zm/lAb/TjBsYYFKk6nlxzPBuylbZKxsLj9/OdcXAtATuoBGtuzWiUQnHJccdyTnGXWqXzK0jYKGf
9wIQyr6vyjStjfMvp5etzNGVyWMCDhr7MrB8XmhWbr+nIS06s8bmFaNuqJY+52o9QQecpMAod3nR
wPQ4wPxeMmz04dTXnblecsgaiiSuJPtW2D+pK6LDalRDOanf2aazxHtujrVbhGL8R/ObjZvxq3R7
KnjB2S3/VLwYR3YFPVEGRx2ayZdR4AYUsqicHl1LybJaXaMI0CHxAMZIfzoO9N2GdvbzyRJpBDX0
3VUVeh9ZHXdz3HQLoIvFhTgzJ3xdZ4NU48qASpk/P8+kgWUW53t09UdtEbiOI3Jgm641xNaDnxbS
bSZKt99HSaBLPxtxgUE00METvn0noQZE5TQl+NZpa9ZpM42uIteg57/ArN+mVEfHE7gWAzbNrhPi
jnFfr1gvuV+u/PI7MegsDDByHT3iuNF+m/rEJfUW3hHzwHq2EYDbAjDHQVZUeyPkwfwusqQW3fVq
HE5JR0zT9836MXK4Tn1McSP2vyKOT1VJnZv1ZWzIB8Kq/EjTVMQsReolfbLPutdxXMbZPWKMOVnQ
TQ4cYnAX5niXF91DlXDulip9lQ66LCbB+gjeZzEVPlSoKPaGg5Xuqp36A4Ul7pJPyc04Y5xacwu6
LZn691vkeKZ8JoS5mnE7CSSALL3zbYTvFmNAcGGmwDMhIE+qHCdTAIRZefSlASRUu3c42n5uVMXd
tlEtCgDbyMXgoWJnOcd+keBchMYxPdKrJ0fGkVWpVs92NsYaGvk6+B0IsbKgABx2/p1VqyAsAoa4
Urc1ozFFCmLi7Ll7DxHjsJ8G22Qd+eapO2XyGGehVbGbBWTm0UuT0yM0ZICptG/HSDGi/sUC35UJ
Rdx8k6OUiJvExDlpnmLRperY6Ce/pQdIXohw34cuTqD3vN0gsGMs0jc5UQMtO01aPK+qnFQwHmz+
cFSwoa+qy00NY2Qoh+YOfo3QrSn9uhGafspvkfdIHrvXZLY5z/fr4SFp2dp8OKCcxL0R6oeJI0op
PMOWNu8uwxWqgh6lYSs5C0UnmXKj9IqttwHhmAnBO0X5zG65jpZLmu1TZBT8CHF1S3iuE8jVuY5C
s2Q0S/4HnU1ZIwXnXPD4RxrnRQzTZdZRuqW6mjSjnj1HzGYCSt0KgvM9dre4mVFd7iHdD96o4Xg6
4E8qSFTrXhcwC3Zf3YaNLHHT6aAbS6sb3Oq6EzbKWkgiACVIbYc8WjDBElXSdiz4L4ewfa7dyQ13
Uhml2Cjd/4Wo4dGTIorg6SSISD4c6a/hMhefaWJXT9FPyCwDPa4S6DEVSy5NMDReIlgTiS85rGV0
lr4Hmqv5ozRNDtS5sHkVSDWnxRTwAp+GmqbJ58KVSupb5xOuPvRCUjKgmbwcjbuZEf3Ooij27/T+
ggWi3bq/lI9g+3lX5QxtkKkG6hJr6cN8KGy4jsh93x4UXdL95lQl+kf1R7LIQUZs22hkLsPpGJSN
C3RLkBp+1Dhjx/qd5ipnd+f3JwPATRr+/wS7Hxw5ocXLsEdoLo+0UxRGFIVWMd/qiSPpTLGWN8C+
LqaHbqLG+3ldXmFXCeZfL+t0cOB+axyUx+H4w5A5JFl6vNauEG+MEM81VWcxYtUy+6I3FjO8J6iw
xI6nbbj7e7Ap2Kd4XLcg2XSmuNZLK2XeT2HGB4TccrRQ/ep8u1OFsZhc7gc1EptTM079w4N0v6dC
5ctf9c1Qc8XwxVuZz93F03mQbNZBiIby49IUV2/qZnh0w8uz73UkX2IrHK9iW/xxfDXv9geupy0a
pktiHTBB3ARYIf+irzmyaKAdsnQtmBMI5m/qx1GGUpKapxYr3K9I3mj4RI5ZkzxCllrxLzEXnhoq
SpQsWNf6HlUAIksJm1ohxbnexk1WBVny644EVAuL1g8C6rDIdejtoR1rI2CuSi8PK4B5Q9OKHko4
hB+ELGXeJzpWG4bxmdBRBCGwerWLifUbRYJwfEMUt0OmCjek6clF9gXCKgrmXRpaVAive9iYjEwn
isd8JDEJYbxzAAjI1hLEHhIzRUxm6gKXLptyS5twBEm21rikNZUWf+FvV8qmYyIA7WcxDtF3ftzE
hi6RmwGmxWonkMto2Y51v+JDfpv+pAcv5a1YY8b4uZrA0Kg7rpIJjMmFtiC8JepxBZR+esmcHL4V
k6OWEU0DMWkUcbS/5GrGkf1AYKAsradg1SnKnybKCiocKTUVkxRv4TwuHPtaJHma2BaolJMyCd7c
biNPfhlPXU9L5Co6l+1M5w7kFldP1/ATsTTDhgiomw1cbCV5AgN6tBewQVDsbKl7Cg8INNUGJaFZ
fg/+ChPjo6S3dBtjnwJaT/GYjS97BMKbVPiMxhPQl7Zu6+anY26Z24dBj5rXQekkdALPY88dA3J/
JFG7nFR9ZKFIbxER+qPZyJK09MwoYMXoQjNf/f/LXScz1VW6GPssV2FMKs5pSnrGBn4aL+T/yuXG
oIWzJFMBANmVP9XNBDL56dG6Dnjli/ID4HswPE9ekTiCYRqaIHFJWNvFKnexm2hQqAziyWunv/4n
isMlnj+UDjjOAGyB/of5mOrt9kpuFU07UcJAQvtGiylGeqWsIGhEM4zCDSWp1gyuajSPA2CLsDCd
WRQrt+Mbo12CfamIC7uHCAXlHdTr4UIlyJBlrVJ3nHgKZHjQoYHxD2UyX67P489NR2MopMuLRRsl
nTOqk8CebSTdUg9+UdB2IY57WXR4flZsCWIjgXbnnvRhu8nWdW9bSvYldvEz16GRZ/aPMUTxhr5J
6tGEcxijwiBhmQKiaH3xe7hhZy174T8A9UvHveSttRWuRm9SYrp3VptJKRaSTkkgSrDbtjFNqR/F
gYxSF+nJfXTN9rNzHHdthgnD3dz0wCcJk/QRQQ1dHvdYD2mOQsiZx6o7jULBPejpHgNlV/aOy+Yp
t1GWYDUoi9yta6kQj5S1uMhhtAMUBkpB9JlFxBfsegIt9w37qZIY+TpO1mhQBo0/JiLck/m63ldO
YhluXk+AlxZKcc5wHuNoDX+SQDF6OiRJ8hrhs4rZ/ahNHU6UHQiQZryOcAp8KpDjxJMEmWyaMXgL
WgqZ7ecGyqGXOSBskKNL6L7MH4tS/nX2Nzd9uRuGTJsDgAFk+RfH5uVnG/JGItg/WFchPPv6YgvV
d9vr1+Qz4cGddjhwBw4XeM0FMsUu9wXbhJIoNwWY4+IOUPuEZ9YW3T899V6WEMdE7jTDTCz8ygQe
WQE/jNpepHBWneIBK9Lhfr4r4GyFclTjR6x/QWTnL6Ny2eMprtTJGc9UV/jIEYTvCgoN2x6V5Ojc
GGUnDwbZKehQaguxsLqbcMJcTsNSM9xY9Pv9GV25vPU1t382GQ60q9TMqt7rpBG0lI1aHzsIgS39
5YL8szhABdYq/AF0rUhWIS8tyclEO1Y8LJiVkWpmTkoMqESvAauWO86dBJ1bpsECPmcPuXuBrF2v
VoO3MbSTJZolSVehdca0d8/qes6ar5UPYb+KEQLSq3X13/p/mvln6pK0SNkRAbVjnKYWZMVZYvjj
rXYYaYkAxFOnQc4RH++52aUJ4PpmEQUNHybofe98X2/vQYOehpQ/5m56M4IFBIlyZspOkfLB733B
v445t32gCtutCFNEFSE4McOhlm/OXcxMka+lElTnHyvvmm/z95Q2tDLdGZ35cNQbOrEoBFYZLSOB
GvaEzEqrN9c1+Iz97/TM0vBRSGTQf7VIV54ByLV7I+OAQ3AeBUcRtA5p0CGbN79BHUtXyhEB7qJ9
KuxGT97krjOqaCLEz5fxFAi8npKhpsnnC0oCfjKP8jEAJThaQkT8x7l9MPQKCc+KSNb0DaK0U6/b
u7kBazVRjBB8i4FXozjCVUS6GyF1rtIUYkrDaBUJC83bGAtUmLrAfdI0M7zp2/qsvsf8HYq7g066
4j4876o0ruKmxAhIxWZwg9cgttt9GKejdG9ApJUjesUwSQ+Zyy5vPUCBMDxd9AhcLhIXmZine+Xd
qmvLELXTW1jWLY7+X8/dotrYjJM9LwZFs7dYxa2D488gaEr/VXAF4ts8A6gvwzMzZ3vUL4Fv5GZc
q6KZHhgUnaTp9hNK8tZxy/7LmpDZ/DlGarwHt7UQLO2KYUmJTK3vXtFLghX5hNKYh9wVAxWiO5za
BmzGAqNpM6LVU6oXhAGdnYyQbQuay4+1nkH/7bw97c/nyVuvidTpgzHP+uammvl4mGf0kJz6UM/n
dHkY993k6RPNaLRhM+mo67xwZW0o+M7uAcE8CXLhC7ck2Y9Ke9Edz9d1yQJ0MsNQbNPcwE5B+zhW
WL9t3nyElf48qoEISTV8UNL61hkQI2c+TyR8JdBrIx2o49P7Dhcv0l+5MJfTnXqiYLUBExSTz3Mi
T5vDemCOkMr6n3sZuNXqss6+90D9Chr+y3P2oL7bFQtVAPw7yXzQKRcT8Y7FGfADpRT3T1J/EMHf
H1hUjUqnQXENtr2bPghVi/U7QM2y4LFze8M6Tc3lFZnH+JXkdMQisZfwVzxVBT8Z+q5953ZhHIk1
jfZlWMSc0Aj7ghtu9t3L9cyjQoWZkwfutPAoFBVT5gjDhkwa4GGAottjrVBusZ28ArFniUahHlyz
DvuD3AtJG94YNSuuS9n7KnXILYUqoPvU8Dp3K4IpsPDf4GoJomZMOx67jHwnPy6Ey8Mip1srHF/Q
p8pI+KFlsYqCASmAGTFlrUGK2Buk4/f88DVC6DNErw9D+MJ367mnKtJWgbMXi27Sut93JBDECWk0
tnQwn4dDm9xk+Zgn3qf47dUtg3pDNHCAMXv4eCBBzXYBZK2Fvsm4FGryduMpnTKhtRuYBcw2vgy7
tHJ09/TcCxDFwKcvGh07Jy0daO4WWgtnfcgIrG2nqQJCLjcW5QZUUiiMHu6H57iWt4BfNER3Gi6a
td0zPvpTmkMdRhU3PLet2AoLFN7NIqwI5psE2GZMzYiU6fcj5G0fBsVJFYhYk+b+8LRzcqAjy3Wj
JSiCpdEhT9uYSdRuvQDBFbNKOIU7Q5WWhknZlmX0Y4F2VBZbN7jir0B4d1m2y//GCpHMxG+dof2w
woadqnlLQSuyES8CQu9L6m8V36VLPPTAYycHj00dTGjJ3Ohsj+p7z/MMmOZ+H2TyCYOXBWnnDl23
zHlvD0MrS0lfeu2Vt41VJLUKmsFdmZCtUNgb9yEtrJgK8Nq6NdFE9Tj6ihNCBTgFI+soMMCKQm2E
M96poSxFtKNGQxLiYnATxbfP/xfLNQCmR1tFxUegSK7CgLx60jdd4Pt+mafHHPh8AMw3velYhyNb
a1OSlPKOyLFd0/h/1PCvqkoXoOaMKsS5lxxenDxQPeakuYvyrGThxUuKPcPgrYslBBLpfoCwbcGw
pE+sHipENPCUUFjtkc83rW85SXoE4llOyuCO26yW85TntTZ3Zw0fZL+99FRp3qosaETgp3ePlRw8
CVO+9Es+MPpqLAqbG9n2ncAmWdCdt07AgbCkWdLsuRzeI1WeX8mm3dSuLqM4+kHUqd3ocXwKoJVt
DjgWbYOGo9uzEUfDisfPsjX68SfLBBZ2Qs63W41RPRj9a9XjSvoI/fmRgylo15jZbi/6vs9gwzRW
AjNeT1U5oiXHDxmvvU2KSh7H4NS6F/dqpgmq3vZLAMTQZ9E/vKciki6AVVSWa7TraygohpvMx4s0
Q8cZwb1l2/3gEP5/ZdAZPM3XZYJcUgp2SJpPQ4kPNB18itRu3AP/INGSHs76shReyg0IvFXqsvov
9EhLwRi2RcRLeejvegx+OUPdCHFS4th0yeENit43oVTFNqRAds4lYpugMBoMOjCjXLRKrbVqzm8t
6RY4uCg7scRgDPuaDjs/687VoxIm/H4lbARvyvMxr/wz7U4+W5coE8BD3pN9eXqxun7+kt+W0pNt
/hdsasJkhGamHukz0t5DRUa5C5ftMUSmt/eQxwI0pnfosVRN0N8p1Q2WoW1/9UaB5SDx4KU5/Zwl
dU+xA8VKorx+EX5HhN8xrjLEOuwPslyPa+7+MEiAzcVZV97p7NYWGs4CudPf6cJQUTeQ6hFX3NgJ
fKAY2GSivUJSeEcSzlKr77/PogtknV4rlUUpVOD0TUlfbcTKp/6IJqLf4QG1bCsJ1gmVGTeNcA5c
5JT3qVpXTogwrXQ7bKWBNywP+1fE+/mYCuS+3GMPEBkZl99K3q4ZGa56mx/4pffcUr+co6H5C9GD
WwH5HZBzKcCvXNP1uuX7gUBoZ/SlCkmgC2QYsfpMng99gwu/6uKTcTu5FYC67sEpUQMR6m+5GmJ8
TGP2zM+At6YcxHZFfBfE6bdtg9WVgkd3WmtaIeK1FFOhyVtzDkzbVY3YNGooBa9qkX9p7w4XCrYX
zfRHjvSWkudrPdPczV2GoWKzlwTYhKyh2zk+vA3P6LvwPl8n48qzwxr/ZCDgPtt5DC9CnWIwWyyF
05XihrL0dyepWVgCadLSU1xn634ngvy/K1nDXQjV5ayRRGGdLPXbdfpBI7Vd7MSsQTc36FyONcva
7k+4t6hDyya05boLcQbKdaO/FQDOLhTT5SFHyWhAUZ9pV+QWzngprXQdVFR29g7N2i067dcukm2k
55yKWt85vaInA9PO2SXPc5y6UAFXN3vhizegiht7JZeH5LngS4Jc+gRxSPYCahGEsNfNdYJHsAcV
t0iPWwjhBpekIJQQwCJ1jsmoN5k/sIBcZaAVlJQO90DJbG11B+LrV2fnyiRh2LUvLmHhFlFsynjy
QxKUsf717t3MbYO2rwNFSCpCu93ZUxYWw4qTOVB7jjzGnja4/Evtl8o38BmqexB2hBfPxzc3h8kJ
NHkiuMmd1NQquGXEK29MlMwbruXKbQz8oZtbd/7BcxSi4HKfP4Gp19QfoUp9+j1gTQcHSbG164vm
MwADauq/vxMBgi2yCIkrCYiqmfpdlgO9M+2mHFOv/b6HbnPwjQvj7vu7apo/WSmmpI6bqfPUanzt
Gk4X0ixpVRdTVsWEY2VPdqdcWGgiwcf0UamKrIMSFflj/d5f2SLfkitc/dB2vnOOt4hNsaB6EJHT
47YOyNw3UXxxt4mmlCkxfjT7CCPLedHDnpQ7XsBTiPkXY3IEaRh5WTaSJ+SceZvI+K6NxLcgt/bo
N0zzBy0SqF54NbMg9xiqjUzvR9mlHD1afeDc1uRhmuFsBAKaeq7NsoEO4QPLmo+uZt6mWne51FNb
0BCGLG5MqCmDrnoYSkwtKD0uvEE+Nf7Ou9avByyiMTl7EsZjiYmJTCbpqST1qj/0m/AXt3Y+YXiK
4wGJw3bCLbMzkrCqMR0doTTjIP4D7bl6zWMJM9KLEnjQn7dTzunL8X/iZRkLvnSuqEISoNzFOcpp
lpCuZVNEdJyCfrifpm+NmsLMBs0dz2Znf67Jm6aNADyFEjFbEAjbBnWm7qJBizQtGjzx1XfeQP1V
pBXJvLwIboSn2+cpbvG4x9HTRn7W6+ulEbnQct7P2+RlyjOJ4d++TIzwdnWPzdO1nHI5yWVmQ4ic
PFzkVBoWn6zU4n9hAVoIf6VFOf0aIZyY3Ml7tQc2V8k94zhFHKOMelCJa6/gk9DmCwcQg/4Mm4GN
BENnEYoc0J/H3PbZxmaSPanbtawC1fL/aaHmv9Gg25cZlKrFAt6FXMOoX0HkhMq+9Y+LQUmtKsIA
Y/HnuPxhr/gUBFKA8H0ypB+OPHenrz6W+hBJ5+yjsHnW8bKMxaWh8yOwDKl288YH1NtMJ041QOKR
tILAdjxqjZX0nyyBXfjoUoyl0QScq2YXXQJZOeoFJORJ45iBnDOy0tANsJrk7SJxzUGhl+iYfoKm
vpsh16nrwfiI1wr7q2u0JYqjAHIyrgRsslLc/pJNGSm5hScDWz/TPqr/Ik6sTg52Hxtx3ujLTsGT
0ElwN94d5Rx8Zs/qgjGg8PIi2VYu0VP6lTHLMxiQ/L2swqFLjyDfqE1EQAOQN0jzteAkSzfCLis8
0FjVHc1KHRtKnF6YLmLTYAS+59zPcv/g3MwsP/OUC0ip9Kzg7BEHCYKiawwhniBKBBuExMZajXmV
AGAkAeJMivdkgdi9QzKIZPvu6poKx1Kb5xFgHhUp9Ko3b7TSo3DPdmuKRYi0rOpfW7zHFSRYyjVc
UAmrcfzFKUo1rWQYT1ev9V8/XR26tF2TD0N28C20DjVd1EAAIApnBds9BFFiBDTIrFooAxEYWOKN
DSTaoP/OA5Ckt8dL/zDq5pynJMqii45qhN+5v17e/Bf7Ln9e0Gfsav+lsDDGd9DX652RjzLKnb8+
+dARZUSIMNlMaU2Nuw7il4RKXabk3hix1fGXnHVKVqqvelEYcFhaezLGI01mpzykrUCSTaBKKCOf
oc1z8zjTAA9DMXxzVJCbSGlhLeS5z6BF3p89AmIzlWDRaPfIW9roXO71kCIAEZmIR48w7mRzsgIw
ZzupeT2BKZZXn8NoG1ZWdnkQ49UI1PmFjacsQcAvGB6dHGF+bW11QynTDSJsdlkyJ8PfkkVE5zR3
Dr1OAy8t1FEfqMcLzmKgB6eurRdC9WnL+QPydPVd6onn0fK0Bjey21FhR0w1wMjHTiQesA+00x9h
L5kZd34nyGAG1PiAHtdmmqNDKYHxUH0iE9DVCMkutet/wa/skRvqhzK/agauhPRWhHh62xNrHSbo
0nG39PSYL3D8MlitnG3B1L4zNCyKFJDk9D1k5AkwGjpl+A03R+VlC4mPQ7ALCSc/sQ0yY12HbOHx
XUDIgC06Ob7gxuF8tnGXFSimkvtal5cswK/7Vx/a467Ijv907l0JSgtSdbAcaYRfHFuj7Sqg3tTc
op8xDnfpR1yD4CzHZirrwN5FQjhEaCLNt+Zju+WzRtjV+0NpDJEsdkjMIPWZYbaqtiXEhXhR3wrX
G7ULdnB/esxqJhOQmwz4pyoMjcHDzhnT2Qn/sQWRGm6pv1JZgh+qeMdXvht7BTCBo4reVX6i544X
8BauJoD5DCcezpWeAzC3/zP9qATRy0sI+F+ihvo+0t1cmjo00PLya8UXGbxYW3nTcHLZxv0mGGx+
t+99uWKtHerLoEg/oYgqSF7KiJlpIA6PoRexsF376NZ4Wh+r6BCE+WkpcZVYL6UXkThT/po4CAh5
SCGPjfcXFd1kJm173/F/QE32Vga9w4xJRcNEpVLLun92ux5LJ9YVKOAuay+9M0ZQa0aWI+cL302N
0DYPWQJ5ZDAXKx5fADum0yb8vnizkkaikWVMKwVizZA97pBkEfd9DeuNiQdIPZ2RnX/yzBwKnh4E
UabyPf5PKlZUDmyjFdTXi42vL31CYfnueDzsJMa7WzYhID+TUOiZUuuklpB6PzNUVYT1Jho90wp0
fy5EIGOGI16UaOYLYgYxZ78cFshcQcjx+JGjb8lg9YMJYrkMY1XapasVAxcK7NrKGb2+FJaR2y9b
AcqE9ZqVzVGwcfQZU8YRKmn/5hU5kTFTS/RlTUQsAKLuYjPcco4nukrrP8FARqaH95XWQD53gBYQ
hUz4Gfp0m2lvF+m+YO3R8cmCkg0CreQI2SMdYtp5Up18n5+52R7WsgRAr/4pdl3pCLncTSKlFgOi
cycwq7HUqae1rpes6vHXjs8P86b85JjseTbo3ne2bn+ftWqNzjFS5VccnS1UslcIXYJy/dPRbnYp
SvelT3E4mzOVv1K1uQDi+aI8dSBzRejbPKoNxi04bVJ4yTWfjo5lYcNT7Ix5EQ8IHlN/dL1eRDu0
n4CJxDho7p/gQvyEPUWBE5ONm5eiDHJTR3UngYT8T0lK3ox6g21hYpQT8R3rRW3K5o18B1mW0BO+
y7aUWC9Jc5XtPLOD4HLykWajslH8SQ2l62vkgFl9hD88K1dQst+SlcueSZ0nGM3mvDWM13OctWXa
ydZsxOl8Synu9sh04HZKtTLm+vhcnxQRW2Nmqhsv+OkGZ4Yjt/1wAvrbGy0wMIz8RAkgWvs5v9tQ
AEWNrYGsYkOq4Fo96n8ffc7WD7XqGbLS9mo6HCd665gZHya56jHgxsMIryde/VzlYhmLpWu4hy9G
UxYhG6mop4cUaLRtJeT9W760YABeh5nX0jGVC0H/rdEuAv4/1t9KyQE5w9xSJ+45HQmG7u2DM75O
dJxDuWPaFxV2IZ3oo4WsBnuo/vwHaV5snbCGFwlxt2aIF3FGJpHY2Og0zusRjnBnSa61i1ChtHhx
fc8O8ARGieeNAB1+WeTwKS2sCKxjyQrLwfkm0WOBNvOBy0GGI3zgIm7c7oZyHcjwdtZwTb/Nc8px
JJ1wOmbLXHg3lX43rBCXUD+wo41gujx+yBhlFXqRaqqBl6rLevTk0SWrexVdTHI/jWhqpMGKrBn7
cV9Z6HOnzVrJCoL/u7SPjY9z5bM3ZoDrIum1UhEW/BGW39o3zfCGFFZINL5IXWL1wu2QMlAqRkU2
HRoUGRRNDPYhba3byBmZNQBWyvSa4zxFx9oeck+IvJTwN7fVuUf+KHQioXTfPQx9rxsK00aWMKwU
HtM7t6K+tyJ6vQ5Nae3n2Xn4SnCMP7MbW47D121f3JrpdcC5+m+3/5wp3bdeOvkvzzQHVGaoWC8x
PofAL81bWSo3Oq3uueaahNkfl0oGFeJlKaO4uWn6ioTGKYhGgBskV+akvSr3/t016hjxWGksE9Qy
GyiS9Dx1wLl4c7nrboMM9COHkx3Na+U+x/C4ZloQMtPBcG5C+t9U8Kn4I0paTYKS9numhdIX3AbY
caDZGJ5pbD9H0R6x66RHCmyrTA+NFzC4R2L4KxEv5BC1MmphgCIinUY9KPo9zOfGJ+ZIpXfDtTpz
ZfJBHtgtgxHpKGqm6txQrzdVKlNSwJmtbpRjoq4LWlciNbh3O6CYSy8aidJ4vKoktdmmWndNlsu/
LROd1WD54wpYsMeIoA06wRn9LijFLrXNwSmzFCRJ+F49uObpI+bXq5qwiEA9s6z9Si7Dv5D4Egkx
yS6pCXW/ym/XmYvt+urQStOTNXVIYS43Zt+kxt2suGAYiRMAToGLJK9jSFnCW1mU3xTTmyF2c2Jc
ZUP4kUFIP2s7ftATgZDa74UPQOy7QAzOCrwvDy/YF+rSvz6DtH9tGPazVxQvMmJVH+B8qnpd+Z2r
RAplBFvg28Z9eWwfjmY0O0FlKhck9RrepSzfQI0Fkkxwc+1/Ue4lC0ztxZD1uRULSSQXm2y8gGq7
V8y2RtGOtWtG+koYLcsyxj1mKeNHskwAVXmVYZv0zCLJeNp4/V71RrWPJRhK1dTdLjtk+7MRy6ho
EJE1RgNYC99nPi+WRFBA+PpfnGmoEudRxzHEsTG2PhPw7X+1w6ll+RisA/ZJ5tUYMunQyXGER3YY
CD2VkJG4vktf7dGE3ypoBUGKP5L+vQvweJVndw68to84MPg63y8PfrOa6fOmOk3n1JPE7Qglzxnw
uAuHj7eJVZJ4u28IPJdKx5WYyK+TXIuWaciajXHSS5Xk+yNBzeUhTeKI6rW+X13ME5X8glEoKg4C
p3xPHtBFtKpeVSoLpzL4qHu7i0PyQLppmuVjuSudBYPSIBSIqzBBHHdGCaqKFXAvS2/KrTqW3DUB
/QqxqwwwM7LhSJuZy9i+0cx9uf4pKuVaCNJzxtZ7zOWnLuZCBVaaG93/SlZ8NZtW+k3vZEk1cd/n
cHH5dQQN5ZiUBBgpPIzBtHXmRUqqG8LBctYYm4QoOK6sqi6u1c4aYR6VL3fICaFTa5ESKWgcgsgR
TtD2UNFbMB72jxd/FUlfI//L4pEbkqH9ytn8ZiJL/Ka5QQVjvChJ3+/BUoHNQk1IYiONwyA2M/kM
vnlpNye1dFUdK4/6871fqkqvqC1FkZZQABVKfWbvDxdnSdrzbAQNLSATihBBSshGhXXZfH4+dWfI
C/oKWT7HAXmFr33Mp8JHcoxs6ElRes8Vuosq6zfDXoHO3AZjpDhehLtWTS+DynVaBrmV6SMFVBq1
XxYFGIFGptGnfUBbUSsLbJxud4y+wTcLM22hcjZUg16GlMR3Ql62DFOO+rurSPnOLrFzg7Tr97WL
Zu/yGWUCAlbO0Pz+nPnzZCidwdKJ+cFkhKdttR1+KSO8nyfGqPcTP2jt5RAETzmp8UoFE1KkbOuG
Dd0YR+IO2o2QDRPbvDUiw4EBqFhqYUC8gmW4bTwbR+aq2cSyj9/yfVHfdMm7x6ZhQwuJ+2dpNi+L
6WZsfvdpubhxussiOGemkMjW4eN9jolLPZE36m/0jt+2lXLBOgsZoVmPlDo6hGzRVwTAiqtibnTl
ji3LhRCpOifeObtQ4idkO3IY35zTePidKi4/n5iKVQkRMY10dJEE8HIRle4u56CEV46Mw6p7nY+l
LotLdqZJdgQ7AqKvcHhuidQwGyuI/zFaJffMIBoveMb0oE/wZhCK6DlVH1MUNe5GGgkTPymL6VPl
1kyPA7Hb/gZxrpxqBkO+mFhJXIEyjCoYAEElL5+AYlYEFyBsdHUQtl8S/XzHZVJuZ86VOu60f2CV
sIWGdwlm72Z+flfkdpFl/uyjxavSFgdaJjRXAy0+BfvNUbpkIJPszO+yTnOzS6Cc4vdDJDH9iNGK
Ssbtk/R4woua4yoAHvM0tPi6Q3QZH1CtmWyMyxTZz5H3gyeakj7N2MluEmMbaBVEOSEbsTX9+Yrl
T8NwqoHzOPtdIURLiNAgCpBygjs64b9ceGJUZAReroytr0CW0kmMT8t/8whrFBPno5ref1Px4YWb
GXSNG4Xk8zDr6FRgb4Sy8uhM7MZKQoNOC9zp56tBYEBvSkOgbMKfm4ptHgNICx9ocbjG1Y6PLRDK
4TPZbl7nvcPKuE6wJxB2RUlK6TE92lvZ6n8bxazJh5ojl4HcRXP6uii6HCnne57Czt37FwzVrSd+
uqyQLjIdrxc0waQdFBPtI8IAnz5KHKsqf6n4xnJn4+h5AIqdRra3yrrj8zHpJjeF6mRyYPS5VL32
wb4B7IOmFteqpuJXn6bO9rHCIn+Wqcw5OeXsE9AgRgPgXAWm5wh8CHSNCzW4kJEArhYxNcbRhS3z
m+U9gaZqUxxz3Kof/8jt/30OjGgzXesETG4y22SdnF4wbz+OIITCnvKRAdc7zt/kF8Cog0O3Mmtd
oODYublkS3dzvzCt3+c+ZqKO363GBMxCC+1elVh5UoaMk41nBBqEllGWNx0Ikl9SLdKg5M+H1QLD
yOAd0Au/4q7Bp8Awa1hPfsIWXpCw/lE2Jf0RSknzsNOaTkE3psRVUc66gbB/rM2vC+z8Kl+9gd2t
y/avOEa9cq6sBgN1uoDOqK9hupI/xewoQuitPti+RFAx/og4OkTEMPZuynfgBW/Kmro9h9VXi65E
SXPZmvApyQTATIVMaCpAj2H+nLTBOUQEwNGtuTh/4C6CuCOJZHvAYxSQ1O0UFpvidFYhZfh1fXX5
D/xmHvu3PhpiZI4xhdALQwtMglV9KTzzFMYvnzLlc3k+p+880V8VECOk8DLix78vJyWfO2KTUvtc
o+H8BEppoBF3gg1MuSXXsLkkGGCVeq2kUyo7C/ol4XZV+jLugdqe0/R8G1N+HL2mAerFAwl9leKe
NGfiFd+i8AxLyhqPwsFcStPouoLwk2s0d9peyy9sBwW5+BCdezOf3/FQ2X4uFYxZhJ1exgFCRhFT
CzH7VQEWkhWNW1jyyLJ3qqLKOzNYDyxfpb4g0lK5+EMCaaCVbhhAC23FRA5vZ8VgEYqA+dOyuIxa
Xe4hzc//f2b3EH0bEwMd5b3LSFeG+jqy+9LSvo+6Ag1sMkrBrn2mlEOtzBV+yvQt4+/XFOefG01k
D3cFvRCQPwXzP0V8fziJyE5+rTI9GVI8w/GArW9/OUJOZrOZqGL2qiXc1G1rKTifWUhf6zsx4XlX
JESSEJD6Ymr+wDCmJ/9oLileM8GYHmDDtlEBnFo9diuZaPr0G7zH6IlB0ckkGeozT1ybwk9r3Mwk
jItrQn/Ftvf8gmY+l2YOQW06Exql/+ESlgVIGEAi0QPq6iwtJo+0uGqqIXfNXxsVVVlO8I2JRYkr
vJzBHtJpr2WTYsrchTFjTbYHrG9C060jXOnkL40j2vrK1Qnfk8FoyDi9RL4OmqBMyX7cQitJ4Sop
Nf1JeTeJQwsLFHIuSjFpMQ2IQAQfwnrNKBvmIJrlUoo+05i5ULXcO5tHYKNNE3XZ5UYyu235gpVT
SDeRe/BEzIPL8cCLqVKXwmtYMXG5qqyk1RrjcNapU+6b+n+JTZS+BcBcUUZL5L2wX8oXTK01oFXR
xBCr7oTz0aMsHdgat+QRk81B+rWsOPxkaSimlSxFIvXLH89VxODfYEm87jpwtUgYnPpRl2cFdfj3
h4CtxAbmQDKiQl7ojkj+RSqMBXDdOZrq8+gTomto11umA5jgMPZPU/i7E2aVUFl2MueOXPrwdzAE
vaMgZYNxKg2PePsrLonN4KbWOZ49Wx6ADRtmp1+19PjlSOSTIha6+8uckizUvCdCGoHJO3ta0vpr
CTycHkB66PMtWMd/PqtdjMKZ6nVpoow9ExY9n3KnIjfCK+SdMRUIHpl+X1n54/ylPzyZWOte33ju
DjSEeFwsE17En8CpwviVuRKilV5yY2K95b/yUry9ZRpoMvd/htW2++4HPfER2k3+zUBzlwOSuH82
wBkMXkn1kBxEZgmxkTBkfZbiRxW+jDJX0XDAK8Aq65ie1hEDpqE97o9wXPatWsegSCh39F7nZvB0
oRKt+5vzl5/GJ93a3DJWxQ+EhRoGBouHmMxfS2h/1Qzl8gsmgBAHGek0vkoJgEiOo80vAtO313WI
8ahTySmjUrogUC4J2TbpVFGR+oyw4INFHIxxbEo7FqmB7VKI0EmI3mUqqWJqKHWS2yGbNAcs3/xC
xmnVCwfWVnGVryI2AqgyXId1YbE0JOnoDlbfOlpj1jJE1cUnHfeSb1B6eR7OJ8ChDgp3heKuBNYw
2t+Mly9VZG3FVXGTj4YOxsuT20J8jCzhdeHClliM5Bzya42ArEVpxm7JaQ0E/IOE219K2lqDAj30
R4BWheuCPqgF8fWzWq61NLoaKOXGgrhv5Qr+GJrFSDGVPEIXyGeIu3U1SuLyQWSIKeS5MMsBGnDF
zI0gGYpROVaLtAFQPI9JXno5pIRBErjnQdYK5W4xdWDuLn0h8M9bM7YliVohjWPPWQ4n1o/rHDLc
8xTv8zF1iO2r7OViSV/T2nl70tBBsywA1xaFft45p96eWkN3AzXmwAwc0JTed0CivaRCb74twXEg
DqTGiU2YW12WH3wjc/v3Q0QECAaqOc7IK+SZowj0/9+Xw6rCAh7L9gNO9qq9cVDDpU7b/FTxDZyN
tuwW1yU6yw43AEB+3qoP8Q5yHTGcNwiVVWgSowW3xxrW+4O95BSyuaLiuRPfrbXMxpIZsD3zAHfT
1M7v+aH60qk+sD2Sv1alyb5zPA75bqIyrOIdBdMFJjWpd7/YMb1DQd9K/hzJoGDFuIsJ5CKM8xSF
rmUzpMidyWUNDK3Hyuj3/GYak3zo5VmVjUvRY/CNooQlvmU/onJPUoCu2zekLwLWP13cPUYrpqbg
nsK5KWR/Unt2stW02qtjdqCinAAfnV/d6cjtvEOt00bmu7bEa5SHwMxkXi1FZ+nXmGELRyDLEYbh
tDocPgls4LPe0ONIqJmdWru0x5TrovErZxXttDAwqV3TE7sMTzFaSMv4QBbNetbN7rONcmRguVUj
1BaLpUH1cKpln4SwW/IBGrMNafyCA+wGSHfVfRqbfQ22etniABuPvWguwZkG+wZa+Qa7FmkeRfUT
UNoYgGo7i387VPxPJa7avkGA6Ci3DSCKt4u9ObnIanBrBnfc+xzkpzlExDucNDnHsLfHt000n30E
5P1l8RWO9pzmq0YCqm1v3FLeaEV1nZ1uXw+ybCmvA7mkyOurJbxpdFY1vjqy8aGVANI4qzPzlAdi
Fc2WXm5ogF0BjrSvE+QbhN6f5hyqPWXc6H4iFrKNbePkrF/UxprjDgionHeu0jOgK+JPmkR+3ZPO
Bb1PwUzttfYoirAinK1GJ3iUliyCeH68MrT7DMcHooJngNife4GkqkEGcFjedE0NvUbHTWjlOkno
Ob5swqZgaAe0KNnnK1WBPEMstwX8zMyg4XZ4KCVqTVMUku9D1TgWy2zt/S53xCxLVCt4rAkBm6WW
+V5Qxi6dNPlQe0jdK9MCUYmmtIToAlvkPwDyq7KqqgHfs7OOcV/tyU3gN+wT6212aa1Mdu1C9Q5Q
MqHkkk/GUIkRRztMm+Linn+E7Xd8+39d3J4dw6v15r0U9Fr1MxsdFJnd4n0uiNvanwpNkz6VXWOy
CYaI4hBUKo4yiyxQ7hcmVAhl2ENBP0ToJvAMshKGQn7XO1IaAisxIpsFwBDBtTJRB9FiCF9YT0Z6
mAfwLrNpeahSCbUMDdet+iXi9RRk4OuS0S37wAdOCS70VbJvmHK8SMUnHebTp8aiLTS7Jkfi9cO2
ShYgw0ObSD52gw4bSGrnSVaCNPbm6ubLLcWhAMsu9uihZsp2mZKHFen0ldxEK6mh6OCfhK4g94/4
JIZMhoAcztj11mNTW4XjmN+bBDscuj2MOkcBJc3CONQ5PGYqRQjOgQhu37sCdQwD8pEEM8cueQ5U
wExGbbgN2AMLC9L3qRYSfMqh8NzVLEalGMsXe1zg2p+Xb5k+kJCT6tLJSJ2rgRTygp1y97eKYJGM
T6MEKQQyp3mgiplqexTkNmGGTWta4gSP3dTACViOe/aXwhFyjZC5819+0GN8s9NOcJXNNGmQa8ir
mCcUzgyQvYQgeBE/noo3r5UalCOB4T7l5C2sPJNixycSJpUaWYC2lU7aYPNr+Kjvu+QK7tT1aYgg
48HO0UMWVARNievb2nR758NKcTSO/38eFhpO6fRk+M/90ZkBXPyZRbHU4gzYRV27NRdgKrNt52Sg
pdIAP6X1Gi8W+sNYMJidojyZhZ3hxGQFVoRtc+nREO503jIHmoFciX2fvIX4le8nAi5O6IxrXtZ5
MObLWcnNT8LwGY30wsKq6Lff5L8vKJCu5UqrVveBFvin9sUHKuwlH68q0ABSdcGLAuz+Ykj1m7U9
dZPlgqFJYUhtYt8mr5taM5pt7BOamDtluLwy4m3wP08CfkSXh3otUctYP57cAxBe3wrhZYbIBitl
0y+/k4U49ajI6v3E5VHLCoGem555yRsAvB5rOLEdc76JKwQrfowv6rrHqkq3KY2e1YPO8Afzs43n
AX2DyJ/0Skd4UylWe4Rhzq9tViUSZWxudqJZiNiT7trGL45maG/5EwEakat0kOS9Iu3VYNUjHUdb
M84oCi6pbNX+qPyPiVc3EMmXvF3jR6DZUI0FwhyxQxecvN2UWAh6JtgyeWQG55Htz1bcHBwAmyN1
iGTSf3gSMkDbIgFMQ3QREDDGe/fOqAOt+zPBledbd6H9ZXcVA2mcIhmXdiWi/ZNBsxvxq/3piBp4
+myTF3kNa2RXxj9WPJc2LsXUCKJt7YL6LW0tcLmkEZ67oP5QmvZXr63nWOn4YEroM43s9bLOLZn6
ez/AvFmd0y9jcbX5Wq6ujGke+6pqTGek0Z+3W7rJbsLjQyfjoAWLc6Q1ek9rNqZ68WdMZ0t+xy6C
y9jd6/pAQG/8A5lvDHzqH0XQZQoaX/4ksuUlARlT1pk1Bop9fK8AUJr588NaXpArbESGkTZESuLT
JJn3JGWZ15jT34LVwhQiZ4qCIhbkFd/y9c0LkfrOsoAmW26qWlgOPHwJ4qlc5STGUa7gk/Ko/fAW
Y5uQx7rxQsjWCn/FFvZnOH7H1GEE/Uydz8LH2wzyyU1xCw9zDCWUWrMfhym64BSZKkoKqK+qTTau
yN/jnP2peqKGfHV0UFBpBpqsGZlfmmuBywmo2EQw/p4hePfjeFl5SCKvWf6kvARVDMx6Fi56qDC9
9pxx3oAWu7/JPspC30z0XRXqebyLmLL7rcpF/19OK2HUouccP9WUgWOmU1XTR6EIWWZnUdwG5IKq
2YsR5yOwCMAmGtaIz2qmZtAngXtZhPLqMRwLQb5lfUYHRgAYG9WO+aT/sERvu14O1Yi4wceDz4jZ
USnxBWpbQ7x9dhWvpHsRHpPaN7ax+ntfqrR9Xq+fDroNM9H2Slhl5EKDm3LkNnwnQlPQf0rgBUzk
3yBM71FRqp7BQVcwTekQx2c0OBFshTU4paqUw8GBRYGdIJCACue5CB/AmchnkFPctLvERJO90pCQ
UnBFXcm9Z+n3FVFHWZUOC9IvkpmzSF+jmWTHZTgSWHhatvwtCEdBPADfQDeLzzmhucTPDhSZrRfh
MXcqeN7vhpe62H4Ebmk6mOajs5Kpyw/fmiE6oxPHBscyAHo5hDVkR5T9+pxhc+ind1exz6mojqYD
hxmc55qPcH7u0CzUni+udxD9vKBjzJ5icNCrdgQo//3bFtg346GmY1537tldXPPCvtSsF8pDKuIQ
SQV/PeB88To18z7sGtDAoVvf8WCTBORTzPmQG+gGo8xj9ED7dFYhb/8MSS7NGaNO2hAkf8dJA6TJ
PtzLEO+S74o8bqQkQmXFVed0CBhuHjMdp5gyaAoKU4nLc7bxd3544ANIMybmBtqrZ5dJ4KsWmaHw
BrIkCLrdS1jYRPUikhB5ZMfuKOER3hGaTWRkvjzgLoPmaZppyGdFl6ekEQ3KBjlNSykUwTj3cShf
2087WwSxbifNDT3o9bJvYZpEpiULufMuN0qzFYblQ98hbmPvaQabnYo8aUhciVVVGwDUavPjjjUV
GMh56u9c1211xOk0KWpFRfdMm50pqidp8vBwfQjCxsKuzCpbvGpKkFRKLl4m/ETouL7E2d8kl1zl
AtMib/XT1Gj79otgfNRDxyETeRaewpNuJ25et0Qmb8oBYH6V/bV6BjexRmaGCjuqYlEMcT4/PWA6
6iJefCjw0HY0HRs4DtxC4Jn18eUjswvRKceOokV4F8dy49szr7a6VZFv6z6LMiCkH/wUS72SnxeU
/w4CLK09DadAO8tAYFetJM0XIbu0bvCHKgh5Bx/ltrMTuB/Wv3UI/gBcKYYYR2y291Ez1BXmU0d9
Ms7O5U9IIHzC2awLAytOaeosHoA6DYQopac/HcBtlIDcUU2zB0cTnnkD7+wjt6fo7zRk998EpTKg
cCDw2Iy8HLKnS7K4Ts/wBulB8s6BDo3I3KxwobU9bS+4UGPYzN9JVaKE+YE3cvs/xuNi7HNx6SC4
9BIoypajXxl7Yp6nhJ3atQXUP9i7EodcBKUIZ9g9ctVUTQjrmuvd5FQKqOBb79vsx18DVH5pduik
9ReqDnS1JhA1hodKgPL/z9r+I2sQHfVmQ/q0hkPpJ5wFTfSBiXqRccA/TOE33K8UPhSxhrk8dfdm
8eKBzRBTpeQlqI6nWwufF1kpa7F/FBDZBPsxiRdlGvHegy+21b6/XN5RUCZPogyJPKeCUow6RAcg
YQD4BErR5jIuwjmZhzhlzU8/sHBwTrCc9DBNGfoqJNtxHFN7HaBZ8NcvLMLAs6RqXRnlMMd8DYnf
vlNn9g84nvAAeqWoXYiVbYXOV7EDsx66KtAP4WlOjWlun+fVtpWoNZsa1lQprFRMZcuZBQogqhhD
u2ilIlrCnbxhJGvhfh5tze7StiZXBz/K/QyhkNzNNHzDFI7zAqLX/5i6GOmVkzh2cXLWZRYHRsuQ
hFyxD85kq5TyjwnGs/zDh3WrIANy7VFAgO8rckspuovMVnwXdOFHMRRwR+ItbvyvWvgnfYrK+yqB
YcBXZZRXG+zeFwX31e3fryKW3gxY+oDyTADc6gBUhLFh/jI1LV0UV5xNUI8tMM0U7/X/lr93d4s7
jK/zqcROEiVItCz3GMNq876TCF5Lz1P2BaGDG4ThDQ0UyLdMrIu6GgNIjCAF7QdZE5wQ1fHN2TYl
KYLve8GywcW5Gqe83xjm070jBdcPBmF2EWXFFo5ZeWzRv3wwj2KmG9W7MZchbCyccTqqKURdT8AW
d8rHX0VOW4uD7CWwtwSM7DrXwWHix49AF10/AOmIRr38xg2hRprP47DSZ87PlJn69TKsowkE931n
sPGeweJJC0O8QE3GMPKAqfwGRhrCtpY0XAhoT/bakTKE7ZDZSEmkRDI5dKzgFTKzne74/iYe76f/
YB0XZK70FAHRLXsFDhewqErWajjtCAch/rf/ymT8mki4RpspPTKsAszz/qPOSwzvI/53ROrKaR7S
dp2vLMp+zBigA57MVO20sT9OSHVi3yzo3D9VLSgM9tZCNOLDXVW4TSS0+Y/Oyai3qrnT/jASTFhX
nAvgFHM9hupbUwOJNBYGLIPl+DINZdh/FIhjSQ0PA4r0WAd3WI17HYKgDDKCdH0cvBSa/47VwM44
PgWrJSgaPhLWGZLy/lp6vLFiSRJfYX1Tl33Wg998BJf0YctYnf88fGhFX5y+hAF/DyX8aSeqZUoA
w3nrMV5GZ8zeEEYhKqPh42v4S758FDEUmDE5KAQ9d+/ktgvmV+4Gq1bNVaMeXdkRPj8ppfdz29yi
MvMVMW8eYLjKGyoEAmgBrtZCctrDGFCBr4aK9sOxwpOuKKu2xKS9nm1v6nNK1yOvP04YqQXr+2Oy
AgDO8gS0bWK7lskdzL82aq4KhtVL6lmVP5cjISTRg6onQSRforFSJ3LpzJ2xI30brhOauoPs5jA+
PzDTEp+lP05A5E8axxZaGUIalIL0YD6lW31VER19jyqBAb79m8TcT8IIZrAeIyl4eD5bRZpINrKJ
htnoHaxTfmly4erLZagRuv9SOpr+wQ7IrmTwBfo6+t3SxUJ+CtnUv5y5B72tSw5h4LmmTgTC3PSv
KF/qRSNTJnfah+cmI+fbiXzMhJGy9UCrCnB60YQGKJkMPkEnh4k7+sK7O/nPsG3lwGLE/VXYwTZF
qaVNbCNp7iym9Dar2tM2F8HpORF39Ba+hO4zCbjVS95etn+f+WZKXROguEolnHiP3fT8IHgNxhqs
xLaOfs1Nnrn4BN7eXNhdzE0DQY4DHAZObGmI8FmG+n8AkBGGgnREF8FYMTBDaAMtoSl5nAHCrh7+
x6Cx9kxphYfZvHw8uGR3ysXLTvMCWP4SkSezdGyWw3OZOdDoEu9ViF8Q2ah+YXDQwXTIyGwv+lag
s6mNuqjWgz2DUnaWhYL4WPkXBf7cidWS94iWyH8T0XStGrO/ay3QWqw8/VijDhVR4c6lGGPY3ibo
wLNng+C8iRwIgUmxRLXhJgiE5wxj7pFrgoyzKzMtLzTwc5DvQgztqpZiAD9IzxNfVmbAR1ZdKQ1R
9uapNrBuATpXLsIUvXzqGkDQely662SYMEXWFZEblF4rxDU3Krmt7RbDBCC+32+TgXO9XpXs69dG
3K53Wn0oeXybKp+NVZdMv1eJEJ8xVZVJ5bmKk/VhxJ7tUV4eu1dSxzEOu+xHl+QqaVQZRrGky3q1
r17gpKe9VBD2lNkah4ep0GefySDUOShbWalClPqw8U/W6i2/HIhWGgnjR/9rS31VD4LbAN2akeg7
kZnoWGtVApPF1hCy+vSG1sXe45inmxpThcubKBx5OLg/X9wiG6O1YP9Mm21j7znrsf3Fe9KiOSjF
Qe5mq8YUVO2G+xMSJ6cxnUh3AjVFaAGLrhX3OsuMSE7FgIOKbRedj0SyHvQ+i/w8lPuV6KiqphHI
ruz2K0y3v89JBM14l32sBwwg1oXnlMC0FSkocScql8HyXbty1L8eDDMlJupQWnLpQh+Fs4iEhSPx
njhDHqafUAaBDYXN/nTltAE94mqs8bxevlfzJfDvLCn3rgZdPviV16e5A5EdLWHWyrZwyUt/+CoT
fj+BBhtV+NLBbldT4slpoMB172dlN2x+hqG+lnK+9J89mZve3cWuTaNZB9WcEdNlpQvm72wg4Mgh
a6oaBi229WXVgK3jvx3WAUM/UCnVblSlmR/6ZfeJ1jLEPlv+SInV2QQHAD0Li8woNxUk4dJi4fV0
u1GGIMAER5U2dxv2OQ8OoVBTEL90xPxSOrY2iX5cvGfyJiteS5dnS1IbS0QyGPnEYqrMqqdOOSbQ
JFGbGUor2nXz6LsIIfwlUzk0mLSiqqOolyUhC8gZ9NjJRNI6Xw+Uu2trCsg8Y/hN4QfvGRYQZpHl
6G52ZlwhkUfp4iSsN28Un2VIqF7kyrUviAl2U9KmEQjUvc1CUdL2LJxGdmA9dS2O8V5mZyH5Dnrf
3x4+iHB5ETVldo1dRI4gqSyzmLhvF0J5ByAa5imd+8RlcEzBa7qWVfruAFeNvvuGihOwMOPoI+ec
ausaUe7cQHT5iLUZvM5jW9VX+yVxID8eyDHckllUpJp66gTQThZmeYj+7fYO4WnSNWTU7uj3UcH/
pP6hsbed38VgdICw5wHHBF8IKPPzmKK+UWGNnueaIQIBYlP1x3lpMwQpfJuQlKED1geDzZTG5yyy
Zrn1wh6vx65px9Sz4c5uKcfPcx2g7Cdu/4DP4Rav+M5X5yp4hEI/aqAkhSjSnmpNIAaciW4eXmcb
Rhg4c8gBfA1AJI4ACx3rVFPWxeBZXbVetvWmMdfqnRdN/faynm0TOW4QcHy5fCfFvD+MIejkYza7
aVGq60/ETBOWOic2YI/el6BSz7cOptWRQ0pQAt3GbeAyR14RezQCYvB91DJGRgoafTt3lJnbB5iz
nGoOSpbfO3OPmO9WWHlQBHsbF7IQ0AuoPS6fVtu+5f2Mk+/EANrTHyuQ3NoqcCtkgQLxUHkoF7gI
ivljWecJuF7MCn8+B6S3LpILmd2z1eLUgYo6YAphFWXKU3xCEgqI7m3EKpy8mVdoFWajJripD+Oc
f455j+uIyD6vwq9X9kr4ogXHnn+8R3lrslMTGlshnnYPMKUBe1s37fBv0LK0r0SWkjH5jSLmAAeX
rUa4lH5qYAmfitJWmGoK7BfWBiLq8xkIqc9V4WepfnX7zlaZE7n93K8zDGfn9qWif3RirNcUXWlH
BkVryqvttD5XkRn9zV11/c9HauF9DJZhEtlMR49IxojOq9+au8pwOJ4dbHCt5CfN5spPHb/udKho
uCIiit59RXCvXOAPD4xC8RfykvH2SgG31NkiX3v/TbFspVKmxDx9G/K2CLPSc0uiQz/NSp59gyrC
Xomig/5KRwecjykXFutmBPsk9w8S1V3jX/iU/Ee1oH0nbMqXc0LH+ka9AQTHlrFfflh/C/pK23sc
SM/bVt2nLZugcezZxV7AEuER+3NfvoL7IDSk9uCVFCiEXjXY4FmBHADmSTjR8dnN5un4A0bNqbd3
4MWRES8IaAvlTO9a1r42buT3eqvSRpiNVH3/qEUPzrO/H4HL9O41NPWA6kO/GZHVA9QCN3MTxHZF
DMaxn/3ZRdhf0Mz+oEnEP+ouNMyVu7YoQO3Iy02dBNHZaqR0mBjc20WtPXWc1EVcKdwS3N1oGYr2
ZKBWaspr39sBE/z47JCaj2FtxFqloM5frP4gVoXcf59EXTThWKCXnHbEZn2qSIMOPU99c10X3XnI
K20kMEo6eMGuEdVsLKpL48Uhs+I9+Pk3ExfxjytLLwnWYU5t+LJnsDcrlA8cguaIR4DohTYqS3j0
pa6mJs1N9PKDAVtkew5OxLHxhwTYm6mDDb4b9CfRvutdsuV/1obxk9wyY0pPxG4sOzixobVuFW7U
TvsWxqKU2eslaCB9mxWnkQsYO1UZXJ9K21bV0B0pUin9e+C6d9lGJUHTTmjdO/xrnXB9tzyXMpHy
N7pitjKHrRyFsxtTU43j8eCf70rSL7KOu8BkPODoTx+j4LoWyE/Fe9N6VH0uFQCf3quetsl20TT4
oluvQTlZdqO6Y3dbIuod8M9zRmuUFvkIa3MnA82Cdi7wiq+qE/LYHW6FEsfI+dplGU9s56Lww/1M
Z1Li1avZC697TVytvu6MZHHqeZkDhcTWuIsqAdeXOrHuQ2w1f/lMRj9jipOlQZa4eimPmYaG0CP2
Ne7JaE9l4XblJokKo6+gAr6acZWukwkyFuNZ+0bYRaQ3FAmBUfOHsQzbCSGBVzV52MTxOuiTc2Aq
tdNKRRre1qOqcJD1XKmFVBK7Wvjp48trJo+K9KMUPS6bv37ZskYdrGIZLkuc7CxKAsU7rayC3SC4
oAw9zmzOngBe9PcFU1uJEMUuV/nnWYu8XiT3jrmo/cc5p8xb9ulUNzXomwxCIHREUbmIX+CxG4UJ
FxMpkBvm3bOrk8F80rjwfULh5mY91+q2RYZn23403AaMUGhMrkSjIXMaaLpX4xnW4FW3nY0PDvSy
3faR8vAgEFRIEYv11LktZljnzaey39RGWtCYwmN0LroDbocIO5oqMvTpg0xMggL91txU9ZLavHJz
soY2xVlqVx3P2sSO4D9ydERoqLFpH/9ZsWFZEDaz9zg8tHq2f8EY+bwUfFyMuxZYtSrpp1Q0tYFD
x2lalv0yjK3we3+S1f9eaUwsWhWQRyQ6D1bVBpoaPpdDWQD1JLAdAfZlqMONHNcXXGvecT5dZesu
vclumozWSwbS3EP11QX7ExyUaoplI/xgXpTdm+IitcFIJCtduOFBFh1omnJxwAYZcJjy4VWfV2tj
2hH6o6FdaGiAuZFOlpkaYfjj5N7kCKSSKVT2mDuMmYZ3NsBMFRyckOiK1hbTphTBv5GKSRCzkbg0
wZVECVVWQ8a7OEmHhbaqjGjbHGV7FkS0RJyS3nDd0Y6EDCJJNlyf04tEK+hP8IDzD0+buE9zKxLX
yhdv/dlHEnHMVpO9R7EoRMWMwn2UEG/wHJ9lrr6ioevYktnVpfeFzl+jt7bC9hOb6R0dmSHiXD0B
52d2+I21PNaFhcVm8vZLoIr2AU0Sy1dZvP54sr4uzF88HZvQQ5yT06Fy4HhAJGF4acOV5jZ2MAPX
pnNSkjgWfDJijfkjygQlDkBQ5Rfzo9y22lSOPaxfnZb2K5xBNeHapdrikFpuCw9CLwu+PWo6Jsel
dCW3B83MWQ1q89QmK3iGr8ZPV+LcpqKq4Ti1tfvORHsDq/rBBrx8ws4FmMY89mQB8wGDG8oPBnf6
Sho0GeMjjkJXQUSPXozLnqPHaVgG5iWg/9viYq7PfnXDiHndAXuYtoBfgzui12Rj9No6fmcAT4Bs
23NwVkqb50xIgDWOkUVbv7h26KraFOo1wnRpz0JjNQbo515o6+SHI2twt/OUJG4SZ/bvAveJ+KBq
g9qKR1GQh8qNKHcS1N0F4Rh0o0aoIy5rBJGF0lzmPMD4PCSY/e3n9GPfVKN1SyMBr4zzCPaflvdt
txm7+rer89BskkQ8Cs1JkZkNtyaeHwybKvNzKnXMRa6RSq+GNErSHrk+h+Wcx+vf6zXt/ZD0xbPK
cgGPLJjggQV9mcfC/hvjZsxtqrcM15PzptaGG+LKmM692uSXvW2KPoCXVmIN2VvrtKNLcrC3ncAj
kUPBudim60xx1WIgqmkU9buhB9AFhsrP/TYN3OxXG5uEQS/V8krvs+Mp3/A8HFR7PHUtyVaFDEP2
4RNR1AFRoIAmC6VGrQRhOHmGYnOKdHIvaqjOCxe7zRjue+Si3UoWni6HrReS1g57jLzH1wXReWjc
x706mmK08vPw9aQ4kkrkwn27kCkiCA76KVF3YDMJiH6lpQ7XAJ+QWWlMqCVohLie8kgPbwphK/DM
jFjPJ5BawTD9Qddf30atzSzFV5gt6MuQvuGgM11Qi89jRzTmgRhfJJxWzNZHPRRJArVtg9Og0cCn
Yv3/QAMAk1CNWSePSaDLTRXzaueH/DQCziKKkosMMViP5oTs4Wh9LFOTB3RFehHFWmYNpqqVBlCo
UCnmsI9qjQvquu6v+2+nuem+h2NUnPsjza59mN+U48Wxh0AYVUPSmbHwKknPMANarfbZs3vJWegX
S75po4qX6LgGOqLX+4+lbiBOO/upX8O4TeI1bXUn7gZ839nNft06yZRfwgUzKJq8oQ+jLjxIB+iO
RZrkL+fpXSVFtaVOC+RgzC6dMEXDfUU5NYt8Hf6GyKjjWb8MhLuIdGFMzTdVUZE8YSccn8k4ecbO
q/AaTLAr2zA79o7lEpEAIwuQjeD/zf3CiwCyJJmOafxxHv8Wf4RrLZvTeco6EFse86KGQSzd3QR7
XTNV8Iftco9HVBTLvLyVzXzcfmLsDOXorfgaWUImQ7XSCl08oI4QGLRTR9Jm/Vcs81x5Mt3/HbbR
OQXnsGz9CvLOj+JxK60kfRjOB29mmvxe9F7xU2HVJ844cQ+Spa2wgB43DamAm4khwc6s77xMUi74
d5fFRbjGE9AzhAkGv1DPHNh4OrVZsJ/0lpcsNf6y/tfDNQ+SLKnbFR1cTwxoczAIfTiseBxDO8Eh
2lnGRxU1bRZK37SOA76kM9ACR/v7RfKna8NagCWWA9oErr+De2QYopn3GhSyqMz4OdKXRGQWfGGT
3TFnvAVxOQNgzPU0TV+d5tuYdv+xsyR3Db6/7sY6Pt1tECJT/S1qth7hUAoVi05w4dnLbw5s2jBe
XM+ICyOcRKt8R1L40mdneaG2BXYcpORvEe88J7D49gOWNOl9UFAnTOawwsHYpUSBvHGED0tHH035
5Bz9RcRgsyVxhr/KrafA/3NxySbcUAT32a80HewEYzlT2h9rFzKslLb/7RwxgewKTwqTuRmnFf0R
p3XaMASa2gR6rI0DmfiV7xIbJ+3cFdBLJtWOSiTpRXyghTW22Y8sIjWgJAB6uw59+fxAe2jsjBHz
gHCZxlGyBD6lCVvo0kQVrWWOBjvvxuk4wemzFYV+Gq8vNMka2SxSCh5dEcM1LN1gHtcT+Rb4Qqie
HVZ+HKOYij+s1Lp9ES8cozuiSOU0XposmDtRIWrDf88wQs4QmLQn/likr9B+JQQL4ls++g9ORy4L
rdaKlYggwwLAzC3xvr0IdTlvs9huxsGr6yh35AryaLi5ETLa+w5ApF2qA9N33mENTTbiE9Mqv60W
biFg0h4xNRvKY7f80X0KSkZg6seqADTU3bloBcsZuoZtQs8qI8uDQFGmpSE8VtwE6Z4h09tKCtAD
+ghEVUuwNUoOrAYLcL0OGbeuK+VAoOp25GbS4+wtjjAqbCVUa2IEzELw3Net8qgfN5lx1PwMIowU
ukvpuyDKQreOkVohaUKxlx42x6kr9wRTxPBrFTkYVCBKhDCxDUf4NN7sUaVjg2f96p0pPd2ej03d
VaYxsTdww6P+2fHCcoDq6QHloXmqsDv9FUzGHzDOqycOrikvPnURv6wGuhUYT07xBlrdu2ww0cCH
4iO5ZuZiD6AT/JW26f62YpP3z3J9QL1vTB33jtbuNBfxbzwoBGgr2ON60UdOe+xPiQgw4Lyo5b77
Kk+HO+iQ1wOKdOTQ505of+w4HFSzljPvJYiL0ty2MoAqcPuB1az8+lbhWITGY2g4l6WsqqwOnED/
7UduRW/Z3tJUmctR0vYsqHBONn3Xaoxup10jC1Gz5xmnwOMip9yuETwc1/H703FzyEElc7fYiPva
5rPP5PYdtLkqJeojR30blnsPYcsJNLW8n2hct5Dehafy9QuV8cABgyZp6O1xPI0k/Iw+izO45U0V
09DCr07KuDQgf/mR7Si+XNtNFaLMo2v8YiqIU8UHNOG/haNvXrDpfOuMgqPF8yKtpJ7tN/gryLR5
+uvJnz6fPkL1sYSKn1/oqnftQelN7qj5/XO+r0+QAsZAQhIwRB7TV1I75Mi2zK/tuGib7/Lj81rV
UT4uH2LytnSY5uTFqgQ2CXzgUhh5AiT8oma4r/S7zpvj3A6CVkc3IcnNNLTag5KES7L0zweOMGCF
puRK4GNzdauYj3Cb4dH0tzAxpqgH973Lv0sdkBCDRkFMi4naIuQvrMvsOKdaj4LtLhkCsnnDKCXJ
yI6IPWJ+fpV5hQejQnRRdYh0iA6+ERthcqAbriHZFqvYkekalmax3+Xg4fXULmzwDMuYbrLEJEHu
oa4NxLGr8XxiV606GDUnOGO4+d/BknVL8oYPgOcxvWfQYzySxV5vnt6ZlbjWXqE/FhL1/LfIjr3k
unL+8xgbYzXiPMOFu/cFB8BEp1dmcG3XsfYRNFvuY1nvSMDYa4Lxpj+ajfjW4anYkCPKZitBzpCR
uid82Ja6lv4CXLUJmrOaiQf066+ggiLeBqTSp8PKtFF52RaGLtOfgK2EtW0cTK+QC0if4OfoeSiy
TDSeuX+n3FTbFJ6yh8Ov7sq2zFnQqxr/GYJI1afw8nSsvCSzoOCu9TO6m8AX7Y9BOplPvg+iW1Ur
5WbgZEU8qAAoezQ2cAYlYXn9SgbIqHNXU6P3o83mI0PgS7iPEqrWW0UKlB2ZjbUKWCCIsb8D9aYk
um34ErIGJVn6kbp2u7hfCFjQhKTwMBL7O89feukmSrjr36BrREg50C3dZbLOgaqJeVW3OFh9EVIR
5Jujx/EVftUbupC96mIzs+OnElqLAlJE9CfUpU59L+aAuCgAJCi/fja0qvoPNZ7ShUApLdPd2leO
h+omzhcgz/OTVKilzadXQXOVAacR48cn3Xsp/FX9aBmok6ngCeRBI/aSaFWGpqSKCrb1V/LH7RpU
KmAbEvPnHpCTGamiXXurqvWKytbYzVEkWwAZFcFFcDPfF9VmaSSmQWv79+5UR7jqh1cekTiWKq4s
6IZJm35bsBi6s14mjr+ShMnlsicMD7hJNSXGU2IvqYE4xDdptZ4UMQeIx1u+HvrTKb0KIkpZPcFp
O0LxqSxe7u3kYXwV6xHx0q/GJQcyeWAxMunaGDPXsvunQwQVdqskYl36o9G4HF73RLDUf4C7Z/m6
f+5iym1hwFb3z4ETrH94TjCrPNRpDnXciYKCaTTYAXfEMisCDtQDf0U8YwEXA2WNXEXV2C5dwrr7
xnR1hVrnh8mYWh+AfGebxFj4Ib1xXMQt1EPBIpzFpSB0EStZufszvdl/a9YhlVGd+Hoy+F5C7YRv
n6Uv2r4SmxfoJ4eZRZqCuNvluqwPCCpb+R3SXxJ+HX085NEoEHnpH6VHj2efN6h8bz0jMuCkNIYX
CCFan1b0axGu7823SY/5ljuJB5nSEBXmCJ1JgBkP7Lqvs+dFbMrvpJWkY321/fpJyEkBFwvxEB7y
7EFo3dJ06F/GQs/CF7LEejNHAQ4WbQX8StRHBqLNE4FzqPbnFnHDDAOM5TxNumwGH3S3bApsbBtb
NOxZU9nylr39zB3kfMjsmBBeK0e+Pp9kLPcGprq+hzK0mdKv1iEW5w8EK2bJVfyaBZN3w0lghooF
uMeVORIZoc33pb90NKeNj7jhcefsaJ4mUOpW10A+NDzgWWSsvMUhYGzknLN+r5kJ/cMUSvXJHBln
/wQ3dlcE6m46edYg4u+7rnXAIDYwlpHzPPNUE8u/51Hew9Ro9HU4OfgizpDQo46JP+uTqemZ4gbR
rN/0Dk02JwRoWHzeB3/Y5My9/ZzbCI6/oRtuJDpbCnPtzICVgKQgIlHboY/Zbtm1T98LhH+kzThi
N02HZSbYfSChPM+Euwn25+CmUlXsEWXC6roc6BX7JJcK/nyKnFhuQH4B71XAdpNFrj+bHDu8YDel
euyihdbQC4iC2XzZ85qphyVNx8dKCP+gF7Q4v1/wN0t4nzy29SnKG3gQnZWkcNllueHXMsBVP+Cq
BBA9SosbNkLgiZjkv3FINK3W5lUzDHY2YIBzWq9SpX47/HkLDXSBR7qwY3P4PQbMCgQ8twZgxJiK
oiur+O2XfLROxDMEsIjhKgq3inLmfwkIZRTwmRb3dix/bRRNvZ/QEh3CJtt0fEzqg0jHn/Bw35Zc
AajlZce3KJPvz8UJdfOkQ/jwHB/xFz33UGZHDAcQNgMRwQAGtdJkUkY8bkmhyw05SRtHD6Z8qECl
nttka7JLs7RYYxnPSC8zcrPcgDSeQyx0+2kcCnmzz22bqGOERWzncnenc4koY5iN7qJvObo61iF7
etgGiDqua+1STrE/alQvHpFiojCPvEyAYXqFWiLw9Cr+l3KbkX0lkdoTMJ/suDOT/Ef8CaOJogJt
2KDUkEvhHh+4OHZ3UG0Bea9DWSBY/e0VjcMbi++KMKDA/3as+6KXuJ2GNWQlRVW+z2N44OFeE7xw
2dvS9DnjVo5MZzx10FZ61oItk7XBBQpUE2naMX+WMN6YN8UupxTaXvY81e6zUmr5lfGKIxuH+osw
NuGTR8bqc8y9K7d3HcRnajtxPQRa7h8uOmXBksOH9shwF5sprCRYn5689odnRO9Q2tJE7kX3D8Ad
PxkAU3WmrYLjv39hWlvOD5kN7VA3QwCaml1J64jmNJMvY8h/EIlZogLLJfqiwheyc5WcrJuw4c6g
jPta5TkGGaYNlRPjOKFBwmR83UD6hzJ4IbmIZoxFZtE8mj747MByNQMWbNc4A2n2gtW275nSYjAp
mXSomZOitRxuFbaSThGWMBGO8CMEL0yC0o7FcqgTOTYVdHgREyD2KnDvQ3a0A5e/CDTrX2Wa8Dhi
E6wA7eKx7uIec8O2pqBNt56jbDAMa7Qxs9+bbKdQvfySH+LQNVeDRW12/8WC263G4Iri4jZjzmy/
B+7ckbm/yuyKKQ4z/o87jUwRalIwxd/JT14qxw7rS2rScoV6KXGnBNAmV/HX6gKlnGp0onVg5ydc
pnmU03wBR6PXxdZWJINMgY2v4bdyrCNlbxyKZHbrZvkJCZXhK/qviu32HVxhePhgbaCitimFbpvN
KnIqPzUO0rUi0NKX4gQocXsSIZE6blgdYBNje5me8ebuO06+e8zglGog4ouByB7TFD1JgMp3jkUY
NqCOBOZiCJ5pt3pxVbQtCJm7/mhhd6nYGZyHQfO8QpR/OKyYJSYZVSFF3Ii4g5ZkmyIV4PwlVlzV
ruzs2OOdcec0NZzEKtS6wHncGWWjWYh6Em10+VP/yVYOEZMHhFYfJoV3MaEzl0g15p3WpgVpDNQp
XyxedOLVz1CyltSUWqPTtpmXZQS9Zy8uSxH04pRKX/nsoI/YOPV/4lnnDF7nqasmqEDy2tDfxC7d
nUZTDJIjwZtKI+cyfNxjMb6pyXkc8ZXum8aC74O3ZJTtAkv3JudYSR7HS4vLyTQjyBeC0o4z6W4r
iLPNviq6UpUdwXOgBVoKokaQuYQBEZVswj4KBAw6gWw7iqHF1KPlRep3abdL+CXqtiQx20srJlXv
bzSc2JyUcahYh4QniytnqlCwlWmwwNE8uiZxz/ZSYKc/eA0goi71HI+t+Pe4JSANzGhkQEjcq+/H
RVKbyFqHmwZOKudKYoGCMAxO63xICBK8RXpIn4Cw8ADVg1Ci29PGnF3EQb+bk855vm8dxotXSUpu
NNgeasOshtPxiif5tDehCf5fLWLQsTou6liyUokN1UzN66SD1s53qhsV8JLPN1RFDJvd21wZpSqr
4THuvTDSP5EmjT6VORwfdKBhMTcF2Fd9LNmyAzUcQGTpk1vuYWjdV4pqqjQ6D3jQjjT0gvlQaNBY
3cVUvBoZ2OOo9U0bfOQCbYYbedlEzMkSxyqBuTWI5LkRxUb7/qRVHr0+fCo+6PG/XI2tLwSH98KE
LdFyk1c4WBTBWQ8Z4Jpb+ssXI1yC9omA/pc3BDe8W2393RL1Br+coLwNt7gvskNdUY/l0iAA6fXc
KD1TPF9Pd5ye0dQtsErWg0b1B+WexW7CeorziN/ql6p6x8muYeu+nPZH5uT//lNQNJi+vu5XzFIx
siUvIi8U/f5MH7N2ipwYxQIpQgA4bNwJohg1aY/jo11DM0lCWsAtH+9u9u9F1w8J3bRExu7+3/Cw
+91CDvM5OOjx2aMYEwGwfGLKGzFCTF0zMcjKG1abfZMjvPExjYKzJ5nPT/j68Cw7UyexxEpl1cBM
YE7gDU5WRIMcD8xqlRai0vkAkyOM/WR4JXDZguXWlWarnTcR+hmiN800a1dFJv3qeyCm6mpOtz/z
0OYfY4KjQ0dYyf/hDi9sicgOt+sloQ4sVlKN9T+G+JpGb+lMdyKIwj6P4LXriU5/s4jsnHVhSAsW
YBTyDKc9kZ3dTQkXA1HzKG8D6N8vZC6+rO6BIepWcW4NKoioWJuxiY1LEAG4yckosB4PfxwxYSmM
b30xjJKtg1OIl77jaHrsrUeeD7z7gx5h9x42KGgDgWLccM+wB6FS0qWe+XvZ5k2QZRX0RJmrtu15
ceHgRgw5SQxONFUQwydYfqHvyXelXA/mfaLtvsxRVYcCbhBobk9fjH5n0suTub8b6XtBLdyXID5Y
qyduVM7dKA67r+1HzNR7NJeqBFVMJprddGl6mLkqjot0h/ES6ZKauKP5wHcETejXocpea2wkTsGw
AwnXxPsJjG91xV4hMz6UPi+hW83zKz9zx5NvY+T+dtLVJ7yZFyMY8Q7K67lYwzRMH6nM/8DvSH8j
kQ+sTCuEYItgl1aZRj5T8nF7S51Xpti6V6/Rsj0DX0+8UT8bJ7Kk6GH9E7XTqXCxKkZMZ/IE5EIg
eS9YbN4gcUT/odugyqkCv+1HmJ3DbgsLr1oEqmbNiZYCkT1BINXyCDENGLkpaH8yjB90fepFfuFO
FxlkGf3BJ4ejh/j5WC2MjqfnKkaVy5BVuYULRaVixgQAti/KkFQBDRRpXt+/mCae9jiEJEoE9+fi
oZ4xS05yBcPFwYQOa4P22EWvF9RE1g7cSCqN+dG58PTkUOeTT8Lh63cASMQmYFfs+5sWxHZdYrUM
ARw0zLBAavScU3TrPHEACCt15O4CRGNs1wHe+tXIwe4GdL84fFbAGVCphejXWG4XZwpaUOescp+I
VUv3Dx5WHcCtgjoQ4NSqQ++1rAm0CK3GSLTjmL7MizFB9bAX/EAdUf9C4igXRbglczMKyOar5GtG
SBFvNBmsf+2BDv+mlN2dUKCN0/OAaeS/4zZG37NlSWLE7Gb0lWvFtdRFnPiLTJbMlK3NW9RISYC+
QjHDziC66wGmqyvdwyl4WFZmTiMHnKoNJX8WRN9dQZcX1WUPUaoLPYpZn3/Vhbe0nZ+Zh7fFlfmE
VYYOkIkt/sICRC9ZjzPhsqBgd/IqLASqfD7LfNrXgcDJwcuq82BDZiPALA1T8I0dLZosHSEOAReC
e79t/M5p0DYCo66u/uU71NIucfSU4E0NNsVGJuZRT1RSkk+8+wDPbDppLZQ8P7WGmOp+rUqnLgdD
BVBMZ3oiuA/kXHjzHZ8lRSIvEzMWzXLPNQ9mF1o7USqjor4XSZVkFj0d8VjbArxaoUEDuEg0xtMG
7FUgXINVF32GJ4Y4bLI7ywfhdxovL6KQ4FNnmiW4uqSMamU5qlgArbyvxqjPZzkPtqX+M28HCJhg
X85O8HjgHmhY/wdLwhWHdLNo1cXzn0x1aVz61TmnKv3KQWQ4iIjKHtyZL1balRhqY2MWeF2ujc1+
zLMoXAXpj+GZC3Ib/2TnVuHO9RDOyZP0W8YdaZDMLoDdWTyh65qJLoI4WgHBwHbYuTPeADJx02/W
Bk037NyP60ECga15qkkfgmCu6nkmlUEniizrXKF3dfuwBb2wt2nqv/+/N/JAhsRm1NBfy8/jP6ha
utZxqqZ9nrJZH/KDJJRlFYdDzvn8R2KXBX2peIxf1Em9UBbkk0AJINBM0A6hCnBYCWtmfKD//cAm
sdAfaRcKxDRXs2ZedDeo9mawbAP+X2BS5LC6Xhi3VJCi+XE+FxbQCiLpZavqUTV/U3zzyrTPfiML
kFfV+jDAwi2nOZ5al/N6nF7lIKKXg1uq/Lvz3i9IsTo2o0zcVALcraDz5U6yA8JT71Sb6apjOjVL
DoLgdaIJMEOAiEPNjUKc/4MSzjRjcEDrmx59UahWMGsZlxOmdLiqgs+v7SRWH4QdsOnvsg+C6xT+
qmVK6i2P2tL7Y6Yroq1jdsUGJiHlhaUb64sC8FFaen0hi4s58ap+8mwRCdq64Ww2juhCFDxmHb/c
c5oES+vDXawyMFQIlH99AQLvOxCex2yv1YGPi74KCbNG8d1DkSHjeQ2ckMQ24wMVDoEGkB/N+Ns4
FIKukuFh21lEO4+dsVZ8o+C29vwKDDak4TCG7i4YhmhpKygN0CM+9ob8zVm/HpjAFTz+J1QGatrt
gHVQZpQTer5ceip2Urb/LH2CbVWEPcmO5PK9Lup2JRcqXxIZfzc1OsvhbAHgpcWymW5yvANe5gpH
OYHVclqhcSzfFe2Qh8icls6h9aQLGeA5jijErdK1U/iq12brpPiNu6Tc4rHpd5hKbQUH01PLSMPb
uNH1dj4XNHWHj6X82QUyqcFkHh+QyPxlUA7rznsGuHT4KT2Gu55/xArPBHO6V5v9KxAOErvWoyEr
NSjTW54pT0REKW8UziRrccSQa6+cFylQiwNo3/AGKNKEpJ+IUN6mZ9yWfVjTm/u69NBvyO7Xkzsa
5q2ePn5kMSNFkIpIQawavKRxXVuVfNLFe+cY9prItOqDlKYVvF63pbaBofj2e0fJxnauOjVOYm+c
cRn8MsV098XO6JoqJJ73kNPgRSSPd5C1hvOKAjwAuOCk2csFSTWzYoJdyqdy2qR0X7YcUzGyb6sn
GSOTLQC05dUgP/gQo1rGChaHaSPYPnBC+ZVTNpxcwq5O9M9PjOiB641gkMVbsGuMyqbaoswYAZU5
ksYBHnMwe4MQe4q7WmWXxYdV90LwMfoUlvEGjOw/ab1VDKyYQU0os0aX1COcKjIaA+5B/ygDbUYI
PvFpdhDeZpRrOAASME9SXRMaeEV7GpHkmRMUyWa5t1e+3DW+e5AbxMWwcyJwN+ej5NcxHqOUHBpS
XkpxcwYyZsFGFu/rfHugzwM5/X3/VjxwxrKRkYvPZdxafWphT3kwgNkl3kL/c4WooZaiMFA1ca6C
KNYp1Naml+XGvZKiwjNcZ8IWG8nsfEYkL9U6bv4rGFT8Lwt79gElg0AwcewN0NWm+FjfHxtLLsXK
Ce93jYS66YgwSJ6w6OBkauQrTpUXsH8dnipcLwfiPhb97v21p6rhf2MORXKE33MdKJvYpu3pyC19
3sEJ6HwpIMI1n15JJGL8V2Yl/J3fD3sIbpzDBCOGAONPSlkrW/xFDprpJLZ80E8saluuSInD1cHt
8FF/SfkVJL1XaZpRWjwvsSoCEJLmYf50YbNzBwGCnbxVTbrsl3ISDjKi1I7/9QW7ocRCA6ciMIcX
4olUqnzA/F2Crf3AwRQpTFT23NC661Q8RSSOmp9lW3xpjXo/6Hy6x2SMB450+1PbbPgqBR8nLe4+
EGoWMxSbEKkgreJ++XGsIdFa31EoMLYyLnBkczoVNfjFXfJPJnJEXexh85rmyDq2is1YP9D3gSUF
gwI+KVK+Jy6UhoUDHMuBHyJkUy8AhDHHiaZOVqUMynGOPfzUrpy/lrMIEoX7uFZkpgfOdjGXJKpe
toIZgm8lCej8yG2J/4PUi+QbhMVOwdyBZ+MBhqL76ACR1dX+jM8OA3lUixhaIpCecn41Cw/9Uxak
tSxy5rtUYvhVMzmQy9HFgtxXzZ986eg272XnG0Vx4Zv58pfBYOEilDTlR0oKMbbxAhngkjKneakE
n7opXQoetVtGMDfIVadRMQzAuuF5MPyw3nnxmaqtiev7uQu28B8lF0bokqSN6Mkongu/udS9rGqo
qvgbe4Rc5c88Q5mrFOwYiiah9sp0aLeaVf9B/1BVoHJi3a8ARqyfDOci+owrdVS0UlCylqHB4eQR
khrD7wOgJmZGbkLNX0Ef99ziZmAy6H+Qf5GR+cYTlVlG7QlmpFzkQpYyhfV8RuIabvNMGBDG4tAe
voCGeFiVW0ptofchA09NNu3ts7iaD9pAjlmvJ797ycfgdeT6wkrpGH3iiNhqzmSIR4aBmgnFTihS
swMXnyQq6W9JHSgaLOOoe748g0evuI8rjr+nRRQlkqKSb/WQ2eNwbazs510SquEKT82T3EBtpyPp
fyTGvg0x7VhLpdfasg4TqEj723Uzrs/tc7BVqLIO1shgNIn8YiuwkWqE9LsQ2oGlR3WFIp7C3G1T
1qrE6Lbu44OQWEFb6pKC2CsSZiv5qyJpal85GNxOSzFpoemLa3ynRGSM+OSfYFWNXkCPCcqhh7CD
NjOsK5jGxfOQKA/9ybOgkmr6WzfQ7WXB/wJMA7v5NPJgWGaqrgUDXDfmeo93h+XWfznIq55vQddx
lG/aO8JG8RdkyUd5l9jg0rDhJn+R7kH++wr7ChYC6SsGcH4kI1KYDfHkFgkF+FEbmVc7b/GaxfMQ
J9TziQwbZVM2MSZ7Ka6LyfPC9m2OdFCPXcxD/26AgF2rZ3vWN6aFCW9GhPlOayuqdOx6KoCgyZQd
VjalLPoEBvvppzltjvE3BgY7goENYO6xw3YlN8CkI6UO+tm9hFG1yMDcxW7VvFm4j66JX7WBWWJ7
S9wC1MuQa0o6WRwzxzCMWvn64nIQV6sCGex7CNeoJmK1+veuZnLQspsBpkR66hW60crbSiFnVjrd
zpIec5uFk4Qu6ejwmyjDTJSI21+r70V4TKv/Rm9UwGFm2c+hpTb2pb9ZJUb9931yyHjt3h7yhsOx
Q72PQz5rCmKc4NRj9FXZL912Y1Zm91q9CyBiV75F37Ga5oue0IuWc1uswK4ZmGgzV/2XrNpXZZnQ
R9YQRBqZHpCW8LMJQjcK1kEq5SBdhZvih9+f2xkBzPkaDKYu1GvLRLzCX2n1tzXVljmyXlzA1H98
t/55JYyiK8ikqdYEb1rzgHDLxpFmIhiRcZKUJHXvpcOABi5aSFbRr42tQSzWJ614xsr7cGXQnmsr
hjrooMs6vssQkyPseIgE1hIYy4m7HAEsv6GCs2YmaLeftzs71k4Y9cxVnX8a030ToYsVQ4uKWnki
9NHUXXpoE0z6b3y0PbtqagNm7f2RGk3moFH0HWS8/vifgkAkdxzjAcX7bOlI2ZaSc5GcamFwz/C9
s2EUR0TH9ei5RWTuhzP2NyGDbMQyFwOd+QJUD6oLXkjB6AF9yxiiBoC3aBizukGn/5cJBI9n/e87
q7Ip+JKU+gEk3MwL6IsIt2+ZPpHSFqV4iXcM/OT7rNB10W7ynyMA/7uWwMJcbyoEjdtHlRIPBLtp
ganjUiZLaXx+/ZkScDMoBqISHRJuLlbMZI3q9I0c9TvoXiisSZrxsaQl9thDfUR7xoYLPnyBgyX9
I6bTsDvo/xNA6dCaoCHGVNDXVlClyAHqLZpA5EAmP7jYGJ3kkMhULmth55REUn5FXKIsPU9gaX2T
EF9osJPcBOmLsZNmEfk9G1ZG2WA7mdE+AsA3LanF4lWhsr67hj/gs79pHAUhkc/ORp5mqz30SGRM
bIKzFcd38FAqRIZMjkWrGs+ErBs94ffz+nC78YIL/he1MasB7luzMeVnv3pcUfgjZyGHUCNRUSsp
NiLURjOkBCPDeBej4h5jJxWsdHuPYYzJ4j5ngt22ln0TB3yYQcbNGxX0jh7+/12Voit5rHDiZGOb
M8FEM0Luda7tgCqo0gUfQ0Kw0QWRqB9Creq4zFqIeIPmFOBKWTe+417xCNkMV2b38r3Tk+ilvUGe
fRdenUjizn4bxYRZIIOVgUQrLE2AyBVJJ6lLggiqzSlm2CrBcnhDrwGSaidK9HHUvnDm0PuMojfT
/rNrVF5QcUahda3i8h22PwveaDyHsxoXW/TEiqlMxWPtVesJoEUL+fjUZULlanpA8L2NUlEdXaKW
Pf6NIcXiRLBUSgZsis4ElVsZhs10DkVLiLUwBBMKUs/SzFT3zCbkb1dHRbUhust78FVytTdQmM+0
kpiMYg4qmgEEb+IVGwuP/78sDdJB0M/5vWUu8N80w6wFnFSR8j/0QMQQ/Vq8WAr6GlyRjwV91tEt
gsMWq0mwgW/8wXTmx1eKbblUmGu1QNPBuN79KjkurWmDZhdKicKTSIMAv8jWebouT7vGOE597EC3
iCoVno7H+PDHb9rKk8yKGU+IQXSwlzvSirI2tT3z/vtKmKyXWeyoW9OvnkZ+iUZh+qR3UUCDZzJ/
B+MjQewCIR+Y/XpMGZaZDl8+yRkMBk1/ysJtKErdCqE3/3y+i4HOi5YG5ObgKLoxArgCO+2ZCoEk
aC49nQQOuPxYwcgOtnI5+VtqQZU+P7awutZIC3SVelLODQqtyhlYtKL3NQNZykxJuYQOuF8cf6TO
iNNJcC4wH1Ag+ihCG1fCEkZXIwS9vp0KRHcPg8igqe9UJMJR5Glh8CqPzt5JIHgdxV120nWIwRtD
JNGn61VZHfL5czvtXxPnmXrgBRDzzPW8QgwfQ2rz/TfxQJtNT2hdTXBVV/6GXtFkUuFj3ln84I6Z
emFPtklVAdj7naCjJ1pZtC4l5mtUbDSbNvX1lFImYnFpr7HsLWrDS5qdfQOeb90k06gF2J4O5WEl
7NqGX6AUYmHrw+CJ4Wl5whBRvcdQcg9v3DXw191D+Lzd42LJKfJ0dn6Rk4UWQaOvOLhvisQ509JQ
u+wNNeW5kOg0h8wLsk5GtKRfXrqFFSc8jdsENqAxjVR20IKkhzznxfOltWwnGLKAWxIOZ33Sqgfz
7qV7NMbcWK8u9fU0zpOOXuBv5wUu2nG8qXxLe6rHxEuFyJlurkMtFnSUGQ9BfEXE168SpILUPxhq
cJ7JZIc/KGiUzqXMpg9OuYahxSaWGp+5Vm+83y5QF5hpdxxNfaw5Gq1RXLWpkg1Z8k7+8EMtF/NW
obnh3C3NicQISsZLw/7RsiHjRK6QRIHtNEJd2yVL5Q4S422B+3npsdG3MWdqODykmWEx5ythbp3o
ui2oSEgesNHFLV3LwBKBzHyJ7lNrAvWTt/HYFkfHe+zpx1FcjTafB8VGr4LknMpCoABb7A8ubD7V
ZAm2+EcMxf75DNKCTFhFyzFYgf4AnVXdJRJrR/K3qmcLwLss7EUR74h8jlWWd3xdn2QkTx7kyByr
D1pj4nIl+bedT//V4T+ZvHTS1B2Vp9MJbBwr2MD4y938v63we5NwcTetrOt5FCjdAD/Nppu6/ULg
OaAUAh0BnGAme2MFqSePJc+gtKkaj3/Axp+wrL6SNYdFUdjMd5sFLEb54gaD3fy+fThpnmuUDAUJ
N0T3MDO4ipQEXhb4OQBtvqf4HYM7dM0L2Tjb0LiNIkwEZmbH6kSSCtTWCuFJx1fu3yPrRYT5aXyd
iGUcKULeYTI2ussjP/V7V+xxSjVODPIAbMmq4akaxcTmL3hXUFIaLhfSMSQX6XU57x5OIUJ1YXSy
hiUgSD6EW1QzEhFTvtEruAcaQ7kU6pBTXArFW2eOtEOLtl5F69I8VwgIgl7aqVyi8sZDukU/kH6U
hGzUx90vDrarx1TNGjl/hGX8/BDHcDMmOzR2ng6zxO7KESjIy52c5fIGo5dpnLydBhr6g1nhwZmP
QChYdkaF8j9iV6f3mUAu9PiFlYnk1zkpFUeYV10VP/3OfTTdqxoyTRnFoc50oUV6NToalmm3pK1L
oiBc55K69Whvofe436SDi1ViPH4cWiUJWOijfvUF24ZGE0ZtJhAB9uO1sH+Z4hc3WLON1STcREEh
2GX+Z+6qOBy0bu0OT3Urp+6/QvXQeuPjs6WIXLO2X/sJZ84McG61X7wnB2zFqzavTmtrb+sZ0FSe
e5t2gGoMkAoopyC0YmIPzDgo3bG2pZEDGUwBXTZIN+b1GuIquwwzIbvoaBltFZzbkE7gbx08vuCf
8BGi4jNyNogHkMi4tVOMSVqHQIyZUmj4yvcChPGtklfQv6s4bHt48BGm8a3B7HkbgXg7eXQsMenc
IN17Gpq7qu9Bh1GSDaMS6ORdmYkc6GOX1yRsQSfhL2VYsXn6foZAVS6eEaTI2aC/g+9CDFNIn2cd
GMICLFSdyoP/KWxi47IEc1Y7kpMiC7fYqKlK3sz5sT1MYrgP3zk82v4fuRioKfjqiDYxJTmcrA30
EuNyuYoJWfsGAmwtkX8so47dM92G1ooAYTVQc/r77/ccPZg6AUTB4gG6cKLzeJhlo4B8uqs2kyQi
6wHcD9hux/8iPUmjYybSchlKMbIHo3bRYpwxeGDsqYzgvrrUvi7bm65uhxRfwjHF3psC6IqJbdKr
j1pOobmL5MWl2iBSLaWVYJXylcpbvByCZnb0/N5PEOjivwSVihK+T6OpvI1xw2K/xri0Ron3gjZa
PVMTV0tAmQbMrMTomX4lK7WXE6TeeLnTydmXCUy0U2vSA3Bfct84bdt3qYcwjR/jVmi+k2TQsOR/
a1uJOoCsPPVc5FBpzAqunXjscku0cpJPdsA7xmnhyHxSXIuNO6L/icrudTYhxZN24BuLTJRubbhk
iUAMLNOoGvFSVyap1sg/aaExU9QmW/rB99tOAN9gZZS29Us6WbNbml6cnw1lhRbG1gPeLkO3FFDk
/CJ9rSwt0X87plrWwZ3aWCL1NJzrL1nqg0QhIiNMogXGLeLuNu5ibC0V4EStAiv8EVD6wNWG4csA
R16tYI4AoDa9n68l2iCTavxzaaLdl9M3De7feYZawqSvF3/lyE4cY5W4c9fFDTOu3oy8FLfLJSTQ
yANk/7GMp8JFy1gWuF/A9GnFiNgW9ASzgZ+bWsQj2KD7OBBjiL/6a3DoU4Si7cUi+qnzTDKTiVL9
sV1RnzMwA2VGtt+tu6i8en84A+l9a1pI3gzTdRyuPzm2VZonuAtgCMHBJondGRQ17zZRg1q5/RwK
xKztfFagAQjMpJ408EHKTSqeDEVyR8yFTwDcOJSmmSMTDWTFLNAQAkOvetL8cZ3+EFmS8hbU3Bk6
A73JfhbX5n7sfTVpq5f23mSkCcJibRV0nSwtKHHA8vzritJ+jUBVjraLwX0ekTSwzLbwAbQbmE9+
EmCxKmKgbMU3zupQmkK0H92/cO2H1pbD2yJ1NmYXB/qERpGobwefgUWM/zGYR1XwtLJxk4WSrlTK
tei0fo8fxmKCLVyL3H15AfGz1ZCFFBAGABl+4J/F+TC7dM2pQimxIHFpBuatfS9Td38vGSHIObdT
jmAQ4LhpUxWO/m3Em/BTHJUPSf8dLD/WC825+cUnpJbEFxqCJU1x36+dnSZEobjHwWLDmoyBQtSz
SO5BrhNev7S/8lz6PR/0eJLrOPSUcQf9m2EmkGtVSv8HpsuRSUldrWC5A/+0dKhEzPmw2EGyUlfO
6Q8AQ3J2zW5FyuA+nAcR+AVJ6HXqtomEkQK+829aMf9+4vNzoxWKYDJvjdIwZFS5J6/+TnaMZzGq
/a2g36v6ULC5UA42DJVQIQ+996wdcM29Hvw1V6efVO817YTryZF1j517lVBhn/E1ykmT4u526XK1
gsBcPRfBhSvHRdqzA2vV0suxgJlFBuG5zzs4jZnSNkOpZTcYxRJ93YND2oyDOJoFKgIei0hC302f
48xXfW+Wt2xEWMF/QbMAY31oJX7+8tu8jcBUH4opjiIpfDgQAPjd6uR8ONm9TtLaXff0vnx2+PeE
UtCkGY/GtQE/aygMOSW4rhygxOmiRlxObjsZzmTaR5QaaOK5ZNhyf5wGYpRzOsTjNlS+dXc/50x0
agpcm9PmD22QpjxBu60uQzlHrDz1q0gSTebHaRbgyCQRyb7YHe1DEfuiOP3JGE2Plj/FLu0jxYhL
HL+i/NcxiKXx3GoIcmMKthqCeBTd70l/w8ImlNXX+EWg3gJgXMbNJhKbywDiguToEgvsvZcbfa5L
IDGDhL7Ab2Qch6cxdDp42VMQmUOM7tFCLASyeAu1WSxoU9NiQOUNxO9Eau7ReLntROlwW2flHwYb
ZWK2Gxgtr1/mu75sL8Lkb3K7qrirZQ91WpL8Qia6xlLAkHfx1zw4ZPBeNNWY7XCIEg8tsDz00mAd
jRAdeCsf8fjI/taAhq+ax9+BNV1UGj2LSKHBYXDLC1+78OEY6zjodIJiE9/sXSmQH23kKmKXkQWr
I8U2qCVzWhvVSxGwVdX1ItmofBmR/jNTx87xEFATG3GAwjVUvOUusmfxYwoyO4RPcRE8K+YILg1b
LAhgUfFDkwHmOR/R3f9EXUTjYx6M7f+Kn0aiGPYTzCb7zqtA2KTje4xBI+HEbOCc7ZJ33zGBX54W
/QnkM12rZsRdkdcWOO2hOYmUZCNVs+q8Hm8FthShtofAEdbxWe3VtB61irghYu4NGbCBLr1ebBPq
OjJin5BMbBpaydVS/3F7W8wzO7GTPMPNgGN3Vs75dWn1zodwSD9pgKFmwWvbVBRPvaaEjtz841aw
k8FL6ED/rsxWIT4EFqVsG4k8yd60Y0vQPjoX7LuHunx+Qa+7x03W7WyObMcG47H4vZhhdonHLQrj
fvwIyVIaNyxnI/jMw0CmZL/DIKHV9TyWWnUYnRDi0bKaymW2iLHEircps0PSzW1TNXB48HsPDcfC
+SEGmYHO90HSEuA3jYhAvw90mIDZCeElw+kicya+CMMrCoXNJQVUv4YRIuEnWH/5KbrGt00uug/5
uZubUUC74rma5yNi0UnMyC3YrfKSS1/swBqICidmuo56Qy0PmG3PsVuuaHZPkRBKLuPzr8/3J3TZ
TO0jgjJJuBm1GrlhiVHnn8ZtYkSPwia2XziFTPd5afS1QtJvLpWR7j/mi6jPZK3f1adsKFaF+R16
TH65KcpOSL+6j10wrg8iP4bkw6Xb/uHg1AVWGx6Zr8nooU350B1/mIdjrz2IhfqsaWqzeMp4+Ha6
ukuOTQAyiZ9C8OBWTIscUmmVIaRYinJ+bCci0dZ1a3WMmvc5Nc3CtMPrNEAIyrWwpwXXsww45/QQ
qNyyliB4sDiCPo1j+qR2ITOpwNVqF4ivyAOWqZcV4z5VaT0eSh1SwStEVUbpvAmQ+K9XnmkV9q84
DmdBHdIzLs+ixMJozLJPLSTzo7NXacLvbC9OSJcrwo6nwm2UhgDk+QPyNhaYFyNo41JK0bdiIQQD
e+0PMOHdIHRGZ8XKwgyY5OlqMx8iUEWKhiDPFujo8izFpVdbAXJPUYMnWGrfzrbjnpVo6Ia3ULqF
I8sVAN3hkJYXps8D8IZgQIxzPRz3O7iFBVnapCuA5k5A4FLpfvFXwtI/p2ExY8kaRyyxQbxd+56D
mze251zNSFJ7kyn8L6yyLHXr9fxjlOcdfJm4mIfO5YWVrSUSNuh57XNB2xbnpgxR1jCQb9wtMEaC
KIHJU2o7SvJewuR745jogceTIKCrAFpIc0QK2cfbufJWg391+BkpFXlpHew+WXft72WaQNmVI5qy
LJrdyPWcpSYBFFbKhMO8KtqgdTzfeow/q+K2G5Pq9BTotEr4grRZsFJxbehiHYtsbud7aPdzIB3d
8HnQ4iF6J1Gv+0Jd3WoCEiZMNbv/cTLjXS+mD7y5srZipyiyF8jzcVltNexTIPYYEL+NwozLTkdX
IPTrXYmIbCW/7BfiOjt26hshpUP1hdDAIxUETYyI25ep0hqbpl4U5TdgZ2riNga8NnxUMK00KbHv
ponbsZMZ7CPbA/6nG8y4p1PhED8wGftjiuT3Dcpb7t/nRt0sEIhvJahloaM9OZnh6SanG0pmGVJd
KdhfQXsspwzffPNcANeJzSELUZDjOMTFqpteT8rSehnb/Hs60fGsKgjrtCzAq0MoxkKVzUT0CG+w
MhICUm0N9yxozJ5U818TRThFABAhNQccjEu08J/1XZJarv5q50VJf1y8rh5wSnGKDwyANu9zAJmS
XqDmO8ywamf1B0QsC6L5FUJ5M74T0MjtI4NtBAfMP/IuttPRi5se01XPY32MA47xFi688BonNgTF
xR3eyemChvbo3XEhxZHM/kMNeVjwwAdKda136X1239UHaRtjFZ3R4W1h2Wznxhoz2weLgwRk8ocd
8KfwEe37oMpIwHWI9qHvR2wvUL2aoh5QnPwNuCYdv57AlpDeAWxtDjLHOoJGGI24pLUnWQHn8Mo8
BDlSisJn/l3fjcoNQQDRqiCjjP2xLkvv9eU2/RC7aCIwnnkmkslZOrnvLcLLATDTpHEHH9gB4Tg/
+O2dk3o3sFGD0b9fKTol+rvDbUdeUgXshVuOMHt8qrb9XLwxozTVnIQs+jNObQV1Ww3TxqYyFzmB
KaTC5mRxcq+DNpXMfTVCD9ZqFpakK/IhIslVfgxx4raGwJ6C8XLarB57yaXxPWhhxodXDcBaE6/H
78zVLTQQLv+4utj4ACz3Pi6nKqxL6UIg5tWs4XzZKfsvBlgKbMfR7yZyiW7kTzyIc9qMup5b5bU0
tnwJHEGjkHzh2fbIuTcVLQuN9ZVCs+LeHoyO50PR6ie9I/M45DzRGmMRAIlsgnu3vIdewSsbw7oq
n5HBaCAsWcKl+/o7Zf6WS8kxHcszQ0IayCiA0wGGx4gmVYJ/9GvH4mY2uKv3wWuSc/yZLVGnquNy
pxt1qo29GNN1F4HPpDpoFAjQZQYDACWv85TPSGrkro7Cgbi0ZiY+3QPLdHjYOJUMl7kcOv7jRLfp
hSISTDnzdCQJJ/AQ66wPiWpuBxfEoOTSXv7mMeG71NL+QIhQkBLiHzU+WzKF2m0yxlKCJKgJu5g9
9QV3k7sWI1PqbFJRLNi0J9XODc28CTb2Gd4gwaSYQnmappTlnLSp2N0Xj+dxX7JHxhWm/GluSc/c
Ihb88kp+WjDcrqaTAfIT0dOPvMji3AcfZkHIdRqNj7w0rCDhHXyAubXZOH2c7eUfddLZU6jB/pHf
Fj0FFIlJ78BW0SG4LXS2AZY3eR35wtCAh6X/f010duV20++H88gvRlO351C9GdFDGsfxR29j/kQQ
KOq1+IkUre/FAPT/cLJtLW3r3wDrldqagrgC6OhK8yn+Wt2AgfhgESip9pmNdP32tpvf1KgeR3ZQ
5WLWtFW5c+dNezOB0AVzUVjYukcaZOWeMGDxclsjvZFK9oYHweAkOZ8hkfSlR2mTGi1ybG0q7kX+
tII23Ec7Ocp2wihiEVMGH++9qx+ItTDrPJAMJmIqUP7IiA0CAJ+CG4Sav8pt0HYTaykircm9M6UD
VjAwt9pYX+Rt4QBgXy7q3Nz2lFADr0kIOr0VG8kFL6k+xVBIBnUFoGzfTZzNxKZ/e40VXw+fI/Qk
yM4X2f7zQ3smlBwoRfTA4QeNaMMMy0TzNsvU4smQ+orvUZr2P+6kMLKOaK6fmeSc0m3tYZVnIwIs
DtdrfH3EBS/TcWmM6KSz/q+9Q4LgIDqOyziGUYnH9yGnjPBzEbxl+WhD/486AW+Xpdfs/GCr+vTS
ZcthbTgnJSosOJYOigxbtJZtgPWStZGv8CO2WAQhTXoibuH1VxUmA+vFdhibubvJSiPAVi8KAcWU
4Zd2pxvoNPzHWH7WikmrqfllOrMq2nVMdP0IvnUBZZWxYfAD6lw5UuEOSvTfgZwA968hJSAHGWtM
hmrzYYWlC2V5M95DhBaLxY0umL0hwz86F521F14Js8m+FzXOPc3D1TarvmkNqWIoZZvHqaT2Ym/o
8e1vlaPAr7mUCTaXcJJmH5lZVXwOULmnDsqLTcAephYmjm4f9Scm4DbjD1EyDUBWLeCpzoem9aZE
zVX+pDLa5m3omhYI8T9+xXBzNNVxf57hZ/1aR/xrmg1UNaITT6287FbPdnhnPo0LaYRMf0ebjioI
G3VrddsY2pTSgde0aemwYLVrsOISmZGPFW12n0PFMAYtLMNxVzqzuVfot1apNGvjetzyr0LSk51e
b3q2L4f/ndKEZ07JWbZ1KJD7PPy7ht8Mk5SZFldrABTSYJYbXTeYrUOKqe+lq+3BzdBHHyO73AGv
MGEzLJFDPvV47NH7fRDEfM6/vDNHvXxrY/kw0IuJp8611GqHCjo1X/Y1qqChk91L9b7g4AN9Jl1V
3PG8wdNvsufXXwOws0xy7yM3rm6jHQtxr79sWMVMxFKw480gGdwKVnGDtEsQnuL7jrDxWp4Y1F4p
pF4reVrt1TNra8KwMn3+BRpYKU3+LQ/NiX/2r5ofe+Mcei9xpF7SVfVFrPD080hXDZRgT46HZXYl
gNNeu/fV+OIlmgC+RpoHRp7On5uyMrdrxZ1+r3Bf0tpluCMwXZYxdWCPVZPVWRgaAtAstk3a/9dP
36Dah1Vft4GGUYfvoWL2rLUvD/lw51x3grazi2xT66/8quxXygBkl76CatR+Td6/MwiPcniHroSa
ZKxP2WixRn359zq0rNWkLm7aT1m5DNvkNEEEipN9OuT8kpI/7lXK4IFCiM09CByfSqeu/pgrQbw8
w01I66LiChsrPYYegw7SGmCrAJYJviW+TGX/r/aR2OPrAbQImFlpkySIcz1l48wSyk76lFk087kx
yycUEEYrTIpgavjnDRXUV/rLWGuE6e45VAp/RV5yjr2FnuP0Bo1aI4fgMXyob7rLMmuoZO93SBeY
ATLcDpGqtRiiflb0QXXnz0ZU/uZuvbfItLfg6fcjQgM57xJ+hqhf0GG1hOYUJ/p8F2G/ZgBJzRwE
tRCbdlskzhIXS91csMlWZk3cqNAhfPtta5hn/+abuU13DZTO3XMGc1CQXtKv+VoYkt+Xjixk4MAJ
+m5A0sDJ4Szrcg5auPUrwkWgOA8S3/ZdZgSxEddvAD5eL9CT5cLjRzqv8NilbCRynCHEXiuuXG0N
o+voGGUzITkDqY6WHLi9LCqinNo2VjJosHW6b0p7KMryjtjM1zwmPuhUS+T6NH5jtKwK6hy1GXPi
a8blBBNcVxAilxZxvGAm+fnejOLdCzTSm695Iy90g1p5AVqPgfx3PXI3+4Uk6lJbg45h8q/3B5uH
9q9PPv7BNd3mpXP3a/C0gJa5j/1Z37pSqWFNd67OZcCijnZFcpavTRFHv9u9migBsJ//h+bAnmfr
QirjoqZcXpKK97UJ5PadiNrx9Si50Ee58YEEqJa6C7slQORhhjqGCp7ojNmpYsyPHhhaESNal5aM
WzXyXhD3oWFMJCOXLyZM9msGVbhpkeos9RLl0uBYcxi2Xu8HN5NFhaEwTVxDkwc1VchliDWlgqyz
B8FPTnIgpsM1YI2sxDRiBEsJ/nTLJ9p/RKNg6Yg1MUN7YfLBKJQ+5shaQTn4REBFiGFoRdBp8aGK
T5XMXQRkf+tsHq3hBN3uuKnMVrqGJ6T88MoawIFlKKhkTF3nRNpTXHljoBNBb/H1PzRgxd5m3ngK
aNix5O3q++iIPBcXqn0DCnKWYcYSRmmAJ6jPyjetS/0UnM8ATQU1VYeinpNrpOxPuMvKjFf8z8cR
KDS8uwzsaLiXgEeVJpLKpwkp8b1O3hiriW2zbpl+dCH9wRfIER2BwjR4Ng1agrBI9ThjDUpcIY1R
pjEA1KtAG6RqYsLm692ApQvDlsMQMBaySsHMRdtvfqwZ88jqo8gkN2MQtImHk/6mEqSQoQG6K+aT
BOw3aAhwH/byGL7S4MGUxqBdzQN6YGL3S9eYPZn7xaczPZOVF8UWupyJ5/OO2i+bp7X/u7sMs+5L
a8iI3Tsg7d+VMCmriM48ZgvAOxtNT7wBPYS49SmU1vJX4DWGAW9PVhuCmZiWeOI2kZJ4CkaksXZz
BgAFyDGdRE64mRZOTBXwBDr0cBK32sGVRwnZxdOp+UBxg3MZOou05d+ANzQE7AEAxTEDyXiNe9nY
JnzluSogInwDcfwnJlF10Swvlk9JwsiE2eiahO01d88W4Q6/znk4d14eRzpYZIHFJzavlNGDk4lC
EXpCX+4vkZKm67rDRYVKHqfa/u5Gz/Es36K0K+O2TfNQKBCOAeMMBcf+MDOAlb8lE2I0mK50wAu+
ZiJlhII5anE2E7hRh//EY/Auj2tRaGNKlKppCENkVkjqsDGfYQOHKgSrQxIrab6okHqHe32qEQ0b
2PFk36uMEIpeSZj73OMLVrp80B8qfxonHYHyD93w6bK+DZHbP4k0nqPMMxQDKuJjclFtIbznhSuZ
xWknvLYLvG8dUR6gFTe3GT46Lre2f4UEkABnkXkA1nt4TTU4HTtVrhZ574cKxIX1geZTX0tAhy7m
BUr7QLjm9UoChB1+T1R6jy13J2TexP0SZjoOymc2NpllGb0+Jv9YBP+I7zVQaeJOyiaqM3F89Cad
LIkwuNr8qipODW8GnL+VocOILcFVH3HMtFceny/DS3tAmhtEloseKLeb4EivgJtEZ1tNxbHcMCrk
d9KkjnyIwHWChg7Ghs7uuohmdv6KoliYkWOCWVQGYfwbYftan51yKKtgYWypC5VfCeh6Gm4yB0Pv
gDXfUYM8m20Az088BjpcuZe7d6HZgp2KN148E85GoVGIVQWuWJHzjOXumDSz666dWB7dRJ9cIBl+
S86qvcmKkC8zqXQxIMaqK6NzFGXSL5u1z/QwU4SV8US1FEhBONxWGgJqfkUix3SJ+5IjsJWcEm9q
wcbWNoh45PKWqcrLuqjJNblGejVqiF48wklJEzZ4sJkKt5N1eSplvlYTNSZzAMCN8lvyWznpQaAq
gblCTvoowjQMvvLyPDf0PqQzPAWGhvzaAwu1Vd+82G0Zj1aZUctpqhAhQVb3z+ydS+8vBvI+j/++
YP2hspts1AcLWiWFtOdTTTw7XSP0Z9yaF4FGH8v17ulwrLM5i17RYJvBwZZa7fSTRmwnYky9ayCC
MxSPGOdVxt9l2JtOPesVP0qYVAQ5imDpLc7oIUIL1v6gLqwNy+tBSxn+aYi0ysKSzbMWLwi32nE2
rlZWwkLPtuIpNlpLOosgtY9oiINVp//5mJZPbOa0xeImF0RE3arRl/giHO1ukMUIE/UMQkEzmlVG
OKuvfLEyLYMZjTB94IAtB3IP4mSLP5V7y5ecwU+4KNaZbO9qQMoK8POE98+q76A02QaLXvFa4eRe
EsngCdtLf7CrrSzGX4WZWfbX7XpyQ6aLx/1ThknrvskReVUxy4UbTm3ix71KHMMwHKsYZP/jXK5Y
hhVGuDsHUChlWV2gVPHq06kWax4fIezxiJSShmLYOBEqkhUnyL3KV5M4DEoOOpSq7nlc6CvKY4k8
jeGnYj4UOkidsC5NYa2aU3G3/+4qgrS6bk5WZaDoIeoJQyfpU4p65+AKNWKPyUkJ1JekiY4kUnHI
HeMneKI0OVesFbia3ilqtlA5l4pxDVz5zlT0bQILfA10Rwrd74e4V85MJGuQ5Z5jmyoswZEOh6XZ
cD9PKhD43yLpt5mmYW1ILE7+D77HwmfyptN159aUF426PYXdCoxxVxpVSbzpc0eATiIVM9CJFS4M
dcxZvzLlvDOMsnUj3zqbKQSJjnpe1eeVqQs1FAX1kqw1WsNTFAg5nrDaKvRDaKB0Lj2dV036z1WI
dGC4I7iMDe6clooVAomMWXxBEHMeGxPk7GzDbjn3ir16SHBFtK3QB2ZlLq+m6398cKtzEPBHFyid
7nfFNJyzYqhatpBDl5mXs6E5WF9fK2b8T8bpITw/9B8x5leciG/3hfnzXgqQcnjMEpsWIlLHECgS
umY7KeY/J/nclt43jxUcaRwqBNO2cEq3q9W6v+e69aZMMZvRnDnHP4Fes+TWuO6DXtc6dWQbK1vN
S5qHPLUeXo+dWmtrkeUQI2rL0HLjex7jDYxwTtDS/hksEsJge38GFIcel5mIAgT5lkZZ2HvvhUOM
V2k8qXBoLEx6x5n7JvdZZhKbq8XmYO8N+bjQOVyBySCANImYio9f8YSJHC9Xg3vykcInuRWpnnjH
lu5Z9UUsTOERaB9bnQOT9HTtl1jyaWRNq8CPrbp8bKTqnUhq6H70eTXaFnjvzaiFF2mWmELXbEk7
8G8U9junyVAW2FNhX3bOOWG4UdBFvVy5HXcALfcX+czrKmkKNuI/ZPAinn2rSsJZN/Vw2e5IHARS
qQ9eIQDR+EeG0wuizHHJpxeSDDoAVt99sHem++phi5T7jZLvyZ/e9WL/lUzsE0dwOdYAY4gVt1Fx
SHp/mMAS8SAULjPk8X4P+mc6mM0B4QC5ZFRoXV6VMsD6WlUDSJiO5k54PhdNWJjlGkrOHAjq2Cu5
m0Dq+fNI0x5iIkb5x7frW5Dg63oERghFmKuvM8tx06m+b9sMQFFowF7x7WJ9EPgKzpbu0MWz0JRG
d7znrl9n0wRIGrAA4LuHVMVmvCOkkytYGtpdnvigscr1OqbMDzkC/qk4i05+rQFBD/e6LErNUhgN
CmYdhBLt35qnZPgAf6VOyjFH6Y+UdQZgvi2lHnnWwPMBhgH2IZJyXQuuUV8wAWJoO5ep63B5M+z9
farnb+aIf/3hx+dkjLV1QXW8h3QSTMtswvz9xr8ify7riXFNe09oPpBtfAI4at1BocXxZ/60++Dc
fk/RzjkJM3UIS5BuPs9ToUmtiayvuAu1EzIGUpGgYHtC66afXLcB4hO3yiKUV2hShijp60d5kcbx
j3M/qsnO/fXMQif7YC4L5MDzoxPkWWdd+bZtnbSv6NGGsrJf2xGTY8M/a79NUgF74RoW8zhrwTYB
3prRchfCB8Ooa/brsexDAuUquXSP4Pq/u57k7By/YjVMCokA227/kozVGrRLlDKMfOCAZ74PzjZb
gV+PFv6blPwbSMxWayEKck/o5LAECaTxvmE8czgRpIEtVOno+ddPzpx8bx9SCWuN5zT+rieTRFib
dTCJwPiii7OjoLy2MwvoMUEVERnm0ObgXjcpEP5CeTtXfz+UfBxUgbAOpnHVJAFijJoZm19c0XoE
8FahTdftxziaS+Bws8o+t9MvGHecPQ/tsmr2ZUZ8TMZjvfh0IanYCZHKGmavHmSfsPPHBWazcN95
ZitzcWLJsknHzz7HPdNUw5ONnN5ZOttmURuC/9pCN9wCKSx9xsi7zXD6/UJPBpgd0HoO+2aqkkNI
z2B5IqTjowC5tJ2awHuj5qWYJJI+K1cnYPc40wogSpb6HS2sAexlkOsD2xqVrc6Wj0F3MGnBifRC
2cUwsiEnMwwxWtgq5zzy1345CcnodsxN2sVjF9C9jGw2tL5LNn7NP3qzenZUd4uFAIPhPtrR0PoY
n0chEiG2le6pvTu95B2G92FFT8DIonhQIwYMedca6RCkLEYKtyNJNjo8oycC3oWqG1op5GVvga4h
iEpDPT06SNRv8UjEFIkQ7bGsCuzU/mj12KKjRWoC2sr8x+6HdZ9xeTCqN7TlqdRwX9IQ25atBP03
T0GG52HoX70cEMc64ou2wrCUMT0URrnah4QULtzC5qmpnuun6SgWiYywDVJEo6OowymsnMksjATP
hjSIu6eZuxlQ95kwoLpAcjGklT5YZTmQOa7lfbsco0fSWXkGSihv5YuB0M6SbFQD7yMwRU9b+KID
iFcLm9qojU0qlcsO+AoZfxjKY0BfWvjLgdan0PFXox5fr0K39w+n2AY55aZZ68+q34UCHKd9ryqS
Fe04twOP+MwDgAEhHEWTZJwD/xJVrwEvveP/LkoA2j+uizLa1+mNQdF0+qpB9WctgXDCVBbUtORA
66cmIT9fx+BefOZQzkwpTe7aC+Pi3sh/gTZyMTU4QiEfmH1NRZAUOg3fSz9QfA+lIoqU/MB3EGMO
XvmV0iNTQcU73Az9jg148MjIUPoMXFJIoI36a+H6DkbJNXRQ8eS8KJ/+VcsIlOgJzkUKZWHstYPA
sZdDnIhG59dCb3tNEWoNLKI1XHps0VXZRnUWxp4/lWLpYgr3Xhji0d78kPJVbDUZpaFSliC4p+5l
w1M2VWUvwo0c+IH68+De2i54IEMJjNf9OUhdGtlUc40sPenjVmgxOWgthGy2goKSIAt1USiwNkCa
wSK/F5Ku8ql+U94A2/+3g+XZy7PBN7NAhSgUU5MpThjpWklsEnFNYPBzbkWjWj8TLFDT1mGwQhIS
gtIB5wf7aUC5A6CxiePALFXppWoniZ3zYjVMbRlIyBCYVqclYnJXy96CKv2Z8Q95R+dMyBzbX27l
66aZMyEC/Fu2G+IzeM6qofRYt3zqZjPynq4NegLURGMnFhAyl9mssaK3g06s8YVh/nLCEl+dJNif
aS7nGQyfKWEUc5oT6EkX7VVl3G8DwePwnlsPlql26gjdivBmVTCDwBjc/DGNUJy2lEy0PpswJLMx
UnE7bEo1kUn5jkMppGM2lhCZrqWcxa/DKaghatcVzS8dscYMZJ1900y+fmS7v/SPm3VuRcsFiaEG
4N3lQgDoh5kUYSm5KCi2sA2AFRq3zTIx8u8eFi2TYeS+cKOai4DGI4hx98mdYzf0G6FvloHJRb4u
q4RPkZgwaqZFREnuxNeSIhXPxdwhnenN+FgEZe6RWzvwuSLUTf9xxT+zAqBG3O5w8mAxq0M3a7vf
31sRFa8eKqH6MO5SfpGlHjdwHbJ9fX58i+97ue/6f2IyAyCbiM3d2iE5wL/5RxnnZC5syjqb9GQJ
cWfg/q6nb9l2sDFLYjD05OkHrRiWTYlgrUYIHHwZNqJ1SdzgcS53a9Opsa1MOqQd1Ml9sXBhqQs+
2kj42qnPq8QqiFSk7M2OxOevr18KIxegZr8thhA76Px1YaElitQGCqk1SytTaCCHCcNUBYwGcGKo
Dliuv5R5ixCPwENossH9CAJGeUN5YQzeTaRtfXdXB9BeX/ooBmt0666L5If9LUP9h87/xqBP0EJB
vS93LWVhYMS+aRGnscqP7Hl4mOPRb8bI2BtgJpjZYyiM8rhxmXnxXeCMToeyARhzg1O9jRamY4ZP
4K538lt0aFjGCi0kcCIc29HCjkeMzTM4afik6VE0Hq56ghk8Z0U3ib6StKaqLsP7Dl4aq1LWv3rB
ctbNByHpu7VgB/DfThdg/j8d+F/WDOHawVzv9E9QRt4U1jwBhYICbmDaxfYD20m+2NAYM9MDOEZw
N7cgZ2Z8KIQRWmaaxGHKLKJNoQJXNcbxTT1t0juzFTNbjnEy9gWsk4xewMs3D94NkLzSkCK+LW3W
iSqLjmXcmxNE8BRK13X5dcL8oVc35AMYefC77XhWHf8clC7HloCo1TFfEw3k3H7RrpNVOK7jvgwQ
XO6gbUM0Ofqy1tGx3dH+Q6+yeHeebrISzqe5+98wZabt3ypAXzO5wLGDLzH7ft25sKySfaJ9iql0
twT+QmzNwROtu5rBLS52Or4gOpXULpKTq3zFaL+tAT+OgfkjC11nOxdR+mArwabVERL1A6ZouQWX
xMp2/e5wkMNLFo+Uj0W10NA6ePhrZjP8NwozmfrlinugHHCQedYsTTfIFwpb1Lw477wDihMry49D
3ohHI2tM//QUQg5cIDvIYEb02cAIzRnTSucYL89pxaI5aGoCto7H9bJWcmjGE96L4s7R29Aj3AHz
wVSR/AXMgYHmNTrctM2NScRBkvrJaMIrvYumj/EN/CfUIFTerYrTR5xqc+zZHKzQs/NMrhkK17K7
kx+FIbDQw8cAwHRXM4K8tJYv3yoaelvMH9E+T1xBPutzLd+No6h77EYa7NnDgpUFFEy/Me26pnqe
TjepFvw8DkU/2LmVRP9UY7jHhoui66MobvDyn23epnBC1gFc8L9iVseCcgXaJzYyhmmpX9HjidvM
GxEjWgxwj328NZxY0ic5VPzMtvNN1qGtFy1E9lB4J04OeQ0EyF6IqgnJ6+gtWpjU0XuVh0D7y3PB
3AxmzZ9CNPklzCJYeVZbArCLmWnculkIYydrk7DwrcrW7zYteceEIK6VfHQL6tQs4wEfGav+lern
uWR76ZSg7RMI8WyjW/A/K25ChKt/7g5rM28v1DWdbE+y7J/dLvcXN/cBoc/ms1N7HzXuP24Iuiki
lGjz02suwnLcBEL3/QZkVMwDxVoW0x98luarXC2TtGfFc/hb1kWgb1aDEnRVAUIpDOkeQdyuUAlm
wh3bUc7kSCrGa76KXH1lqihLU+KDBl7oVHIkcCYarIfPeKsHKFrD16WEE+s21HW3zJjjsYEvsiCc
D0A5IwtUX38v8SKTzsNUN+N2R9F88Q7ecGHPx3agDWS2kmiIuy2uhtCmbr1gtQb5yYxR1gRLZsrC
fAiYW4uLwLqjoFZGGq/rhcbYjQuI/cKGtFuUlMNaSb3uKDUpAyBFhoATKs40x4OHJKRWVN90YLbr
yPyrjkxMZkKLYg53LeKjOzCBcHC94NQhWmDZKhQEALWV24PozFZSIqcK1gaZ9BL5fkmo+o6bRGf9
/Hc1PXoZ87GMH8UECywfFvHYe19R3pNSu4i9HoujxEVaW+9hEvTQatV51uokamq339axDPSYR+o8
zbPcYDqdeqFzZOFGC3SGfp8XObdNO5u/M/3VMxhi3skxIZo7xvhkTMfK9bzhBynxSRZln2Ka+JE7
YiK7Kt7SHGpBTLKKG8pW6TCkH+2oZSNrXmVxG3JHR24m3OXa/Egzz0EmoMJQcTLTKvdrgx2jv9oG
4JoV/avgc4r7mZ7R8aN082Gf3PLm5Qxml8Zco6ckbDvz3/dMtHcQsSeoefDtFP3TPPSTAUayK6Qj
MokyYGmqNp2e8aKfcLWlP0ZKI6INDPKhT8I97Hx9nH7g/vKFmn6nqBwkCACQB8rEBojcZ7ZXUllS
ntFwhdXQ2DB3AiQ/4WUmhruxRTwR/wGNZZjFluHRF0wVZGXgC/wvVunEq8X5jpk+FRJBtBwlzZNT
2LU+D+t5N65dIVvr8CHTys6r3mhD170VjGITup3yaCcRPh+krGe+5UY2JCiUzeztqg8Aj2yD6ULG
LTWdjLzckg+S2kHEbl5eEbyGtk+b3GHON5cWurtFMWzjDiK1nUp6U3apneH0/PSeRxSl+9qkMVPF
IEmhSJxPed6U6U8J06ZJVxULKnr+K1G680wKleKmDbnmDEff4BUv/E/eCURpNE/XqaNbBwAajgHM
bcip6sWVRbvpKQ/vAqkIOCG+VpsoX5Fs33Uw114CiHMjF5aySEBgBxt3sVs2WkBHhuC9oUmoaTh/
4gDPVh02ZYhhWOmS2j0XPBhlZpuJ3Q7d8dP3w2XX6blc5/j+4eIWbiXzdWyOeKuNz3oU8xuJxDL+
yrMEmui55GjmPAawkNPqt9yCMdEp3pVPH3iW/zbba/PzRsECwtvq7WRtpGROs5Q4/NSHpy2azMSm
qhWRX5q+wKU1+fEh6fEbknxFP+WfH3NgvaRMAx3QGg1UdxTz+k2VuUFNcfKV3Xq6d/ybT2Ruv8yz
xOqqTUpR1BiZWJc5hIw2MmDN/qWNsYNjhtJGaWOjzoRJ7SKV9rWzS+Boi8/NEPtCgFReX2XbGRAR
PYOlcWu0KOfBk2bK5HS2bXTM7rxU4vrX5u21whwI5oycDY0n7Ws8o1IvvMfAHatTHTqdxIFVCTNU
5Mr3KS5Xf3vNFDcqT8sm+t5A2UuDq5sySe05CtWVAV0gGcUVqhfDyj49XxcIl5mWfVdTJ/ItVft4
Ex0s7dJN7yOMlBjGwpw07Nvh/aZECHcBqs8jhe8knG4PmtW2Z5GUYI0QRM1F2gqivHY9dkgSILzp
+AMO+a9uvPM95POxroVL9lnGymVHUP69Ir/vgi+gBNEH7ofR7cFJlYj+5o1EV3056rFcb7xVua7k
TZA/mtKcqZux4v33Qa308CnHTaVfS00KUCOsSNEoI+0ueXThmeDablM6jfo67QiGJEz5OwQpGZ7U
lpT6XN2Xa3Lhy43ShHan1sRsHgaNhQ8AZWGC/MU5YwMiludv+M+3Bxiw2au5WWs7JF0mel52F2fm
8lO9H8I3B++jBGTVUmBvxdDDJbWCreEY5mTJgGnDbpJG26pEvtC4sEVPeSMlzNUAo29WqnCgDeKh
YOljouxEc9/gZHD3llEdvoiqlwcR4XNrh/p4m7l0XdgyqoY+Y2o12x7RaOzVgKin3+W4BuvJvF0e
bj0J4xPOwKyNkA8x17JBrhtaqA4wa9mRDYeW0ouA+LbC9ac8NrYISnyKogKpII5hntQwm7Ub5nSC
MeWDFslZt/VhGOGevOxcMcYS26y3g4I6Yn7ysDXJ4HlMcp3iXuWMJafvljI6EjGkj3kWuUxP2k84
N0qxSB4AeGiz7gO85MOk2O7Jt/rjSFfIeWs8oC1B9RpnJChf3bgj0Zh5tIb+wMBcWQ5DgSUMbOjH
S9jUmhmT80wAMhy7BqC7MIPBtNfzdOzot5RuxqQVi/MkVts+fK2AC+VhCxIscR9iBnWgVFp7SP4r
TcZVDmExBcUHaadqy8EeHNJvMxv8fsbjldQSnEFqM/RB8HYwC7vqwZVpzZLGfn8GsNQdh4mBw8wj
k3DN73k5AM2s5hqmsh8Ldk/85PTb4o5GCctFIurrfao9KwU50eG2J3/wcSe+/CnpWKuThyqt5uaL
XedhsIzpSr0FT5SIsgTQBCRtZWF9ydecj9X4JG2SsHWgCi/9/lJQZyZu54LMefUBdZQ0rgkX9Gja
p5P4Al/+ylYAl53j5C/NBAFIEUx/7yeSNF62IEgir2KbsZXgfadYitGDy0HL/rtsIky1xUZCXzuL
kWllvSJrXOoQcwjB1CedIdN8XZz+6EUvMNdVqByAelldDDSyMYR8/BNIAfgQBh+j3+DUBU5iEaWx
IzRC8FO3Fzm85vx8GyjgJ3g0hqRomf6cXB2WpItOU7+p7vSjHX5914vPk1RrfPbPzkiBgw8UpEdh
NEzDhqDPa5o96V3q5L1caJiWKqR9BsysuoHC2F2nnC8wNrOw5spr9HYhfUDxSId338H1819uAA1X
Qo+DWvrGkRGkWztM/FkaHwk2smXARVvAC+1VOe43zgAQzwjnDQ5Lbq6yZ3CFz4jw0hS55AwrDBWs
+VTfzgH63eMwwddppsa2In/Xdg26oYsWaCjypPdFJ2XR6A/WQvAwU2RNM50Lc02vSAPBJ6lJmxGi
6CUHffm8rwGiVbV97WwuuTrJDWdruZVHB8BT8iH9qqUJjMoCevDRBSMs9LszTsU3CWxZHzVhenK2
Kx4J2MGe0EPG4g0+vumx09cPMdMOsqI1su9zhHr84nQR3DkU0RN17iaFcPV3ZLzEKtl1nycwHJAw
MMbAHzcwVPGICJLcyvhQAJgIspfJhu7z5GA+yaYeI6aNbF2FzW+96XZo4wV/nTrn06uHidIqMTno
SPDsIAb3+Dyxnwq/gDgQ+DEELOEZBCSmT/2R+rrsPDv9wZH1LpC5yhGvWnQIj3OYmgnJ7rroxcGA
GQNJ2dwPnuHo4J8cwJ0SXYOl0k9jG45BK9iyjol0Q60xKwru0XEj23DcftXgpB1r9qbB2xJsQih7
GNORAp8L/UrvfVhQ/qV46WvPio3hAQ+BEjQqL+eZWl5W+BzS8pUO4Un9lh2GvdEIWPyEOItI/R/f
LZoTzLA9TiF/ihviGrl4x99fZKRxg5h/fqHP4Z9+KLeOjFVtZdNEHxta9w6HSmwBhZVZ+WD2MXaz
PeVecOzE0eVWEylAH18g2o2HbSFtiekuWdQ9FTwPl/GBaf4KfumRPx766IQQkib1r48evYFGABwm
BlvroOc+mX9iFX2xk8YaG23BFk34eQipLsc7U9tsjdubMC/UXunXq3wAFJahfSxokcSD5eY7ogEe
O+RH/B+VHGJPVo7FpeBOyp1MNRKif+J5puqLsb2ok8aHb0NceJrlMzyX/Bd9Bp07S0O9nE9ekUnq
wSwAghBtYQ7W8T5O412sitjrp2iPbrFGc/ubjeuX5BVJgGjj5tuJ5IcmN1y6CZDbUeR8olEaghMY
eWIZzOLLT22eTYB89rcz+qOGKpkv61WvzlosZ5GEW35JXu0rktwSQVb/5+6fcsjRXDR/JwHAn0FO
A9T0zwVrqlCcbOPNHWnR0LOD9EHgWe5J1T4Bm1PUYFhN/+LaRAvTQACLV/Actm21TAOACTUnh3aY
bbxdskWFmDTrbL7G5Y5zRauWUzHByS/HKYZZX0hCUQ6CqfgTFTOEPY5F1YwCti2nbPt4dpt4KjPp
Cc/0h3GtQz3257GZ/rLdzodAqIQl+JqoK3aUPUUgvzONuxJqI1/mJ2rC+d4KMauk7HL+iQIdOIJf
2YuFjYI9nYdqEhT/EKqLsPWT9zBLGL0ES6i6B/LAoDluYC5v4tQLPWuGuZU8pRnUvuhux+cS4Uef
nzaIBNxyHzCD55DeZ/DU6Gb7+bXa4rkt1ejKtdY4wcV4FeQaylr8XJroKJRN+6NRl/ww5O1Td97j
gVM0owzh3ataUtWmhid+xaxbPjTBbhKJ5jzQ+QVBw4OBJ623BB9YeQ4UoSJejwEwk7sRDykr1Su7
+TRPN/j3omatGGoVDcodOhEEYKOe+6563Dgr0ENI1C1gpbWJNiFpV5AZhCVQrSU8QIJMsXHeRL7U
dYFRJTzvu59VbX6OrTkxO9uajM54H+NEbZM2GLkq6iS6whKagK8sImbnFegw9XYLOfQzhH/v/iV5
kJ6dFaGPktqwYyLBuA4J7rNw4PifaWtJOM7jBpZHJ4/gELe3vOtVlMRrQNLraaVwSYQ/He2looYm
RTnTdo35Lq8IN/8MXtxRDvf73LsoyqBas9gavaQLTLITwDNMTvgDsYzqeTMMMolyNc3lk4xu1seE
QeHBL4ocDQBozVmGmj0TYceOS9PMY0sseaQG6yCtQQDOHY6whHW/Mo4F5MpfQSfX3TdWOL2sYfOq
mffbsXLvYuckK2v2NzGk2ghEvXru5NjJiZWM488wc7YpNkEEIlmNljv741aqUKpUm17tfRhiz9Qj
gMqLumLkXoDOREKZQRQASjvEAJYEkpslQ5nIyzu2yxCP8Xj/syjiSNfW3bF/5w8xW+pmgKlaYw6k
vO2JdPRT/a3lAZc4gPodtNxjv8MnAKzBo/gWrG9yiWLIVl79b7KmupPER1T6T/XbTsdSRCw0+C7+
YsKLa0/J8upBHAdvbpEXuhNk+v34ABNtkYW74gKpY8X/0OO5a+e3Jgv7Z//gjHRG2rYWx7kD/K/e
TFwHcTf2oAjrbb5DFYB2z3sE+wMAtrqfNLgqLjBfsQ6i0fg6MAKIPyCwwGSct4BLNElZZIFJVowY
YrjJ08pYl0CpEXpcNgjBmxIyP6Yv8+9UlILL9+1h+nUJ2Cd2ssh5JxE8yV5UjKDrsv582XzLwKmx
UjTJfzYK44VFhA6TJILTn/4rxEOJo8dLsHD66FqQImQhg3aHFWkErSoj41fIL73TSwXrwLga4Tba
a/lypBiBE1cYQlMKwHsojoj0TlrZYK8IrtnmSpm0QnDsFKJKoOHoMYh7XyINMlUUy4p/s3oPrqLZ
5mlk4u0sAUDC2v51lSGCNRWscPpLESPSUeO1KdMwOutdG+wlOe8hUoJNJgXy7gmKcFDtoeJWoayw
JA+PL9xrWoFEYwHtiTDujL0QR3FvHX+JwBYbhtqnX7ownCW32AbkSaZGMtmsOcfeVznm3qyMpxjR
XGTkIK9OYvwbWi0bIo03NgPU2avNthv2Xfxktrc37yQJnG/jTlaVVTzj+lseTjJvPb2SiJufa1bN
jhqekllgmqus0oK4jz7ynoEE3mVFTXH1Q1ky4yD6GmbcdUDLcSiPEXftvNqQXOFmUxVZ6rY8f1JP
uIHeZRKfakazEeGTv3PFsrHMq8qU02bSVIilEe2ntX2EvMbK6Y112xN4v9Qs+EzthcCu4IEu+bQg
pOnBmtN21E2RN6Ow4QXYY3Dt1oRI6B9Z569FfI0V0u5SUMgnd9HEYpSaatSaBNdjcGc6FE3pxEKt
WPzMSBrdESjidvQpM+E0L5O5joIJrx8Q/nP0f0vBPCRsNNn9hCsoaSUwNzehYM3Hb6KBQ/qXH3+A
UZ7WeoibTg1WdLETe6vLv7v4ERaZ34v1PFRBn5XOz+voFa5XFQxvn1RKlvIy9U/gXBsxPOV1OX/+
lBaDc4dYGo3LdBexRlx+HtTbzX5ynT0R38F3/q8/qbvwa3si/FN22/5Q8MOMz4V/7Z8L6R+Dj6Gx
PoVwZu9UVanortr1kAooPWZoQkvfd/xJsyZS8kbKqON6yf8ak2eiWGD1YYoPtXFDyIu3rp0QqjXo
CZLNSVBs9DOKqpza9cvWw+rQVjdWoWzFZJyfNBlgPYcwe/pI6D+ZRU5DzjLXVkrEXXzQUhxMIerA
8SDWo7t8HdxDcKR4xRJdFnjEMiO3NSdgPubkxLK641Zqga6JeXEItGcHzjgF6Hu+9LhCrlsxaw5o
Pl5jgEEMG/6LHF4/EQf2KI6naz1pbXF9EjjdmEhETm+PiIEtupMloPq7RE1i4mQYMn74JElwZ/uL
OENbQ0okt1P04stlm4OgHqO8z8dIEOk3Seu+AZ56JBABMO0p/N4sVpB6nTZ39Ory5nWWqgVgadjx
FFRF5mq8SboAUTlfQj/Zps2SeDvN8ZrkuZMn5kh2TswTXrGJ/LoPkIvJPYOcI9tc15apkxGXQUjz
wKf+Onn25ghL+46ybCtm67+9Lxjk0qURjADlsjGBkRknnXxpnrOxKg0M71Po1JF5+WIvWgTq0WDR
bzvLbQaUdTpn0d/ODZXWdGOdWbvkZUcBaokHz+ly2fa2DpDCbi6dr6YPIjJHoOvjE+Y9zRgBsMKE
eMk1d80nkf3TMs6/ocjiBsUe385X+eZ80dOZ0VoO5DIyoih9UP4wjKjDw/Jm3YPqH3rTV3mo91tU
uRTlE5sXbZEDTRAf1kdoDQzYfQMjk6ahC0Nt3qfoZcDy7qLdyxTwaDRVaDMq5wGYCSYeCrm7w42e
lp/HA6tOmuFMBIxxuUin/Ei15du7p8Li/fGUGHZrcXFBvwTkWtTVUoIJmQC+HZ6zvs5EENqXAJ2Q
FsHVni3N+jOwaEKxPaa6252151qoaYWlsHqHCL6RK9eDO6tTjCdkct/46xXoOHqAEiyFbiR3eGs9
BjG4iO2iDazwdk7FP6c9INWqvkbSUmyEz+SbZMcUl5DjkJrfmYhWi/yEoTFeZoONVCx9rSlT746J
XZBVOOkC2yG+Jg0M9WIS8uATP1FZikaqqoDX8/EY5f+tg09k1SAzVGkrs+4zN2F98PV13K6A2eSG
4G9x+j9T9LJBoes1I1Hgx/Rkt5NmeLyQpkY59pyUTIReHgTfmDAQescS6VsNpJe5Q1Ie9tjv0lQ1
fdY/01Wmy5z3WYcoFjIxPJ5+kl7Gf6epIFTCBtl8s/Ow2LVCh6V1t4jIsTzglaiH9xgRBStbUGtA
surkzfSRSWugpaXNBpD/zjOFwtb//rgxQHl8qHNXjtJk6ei2/LSyY6Ft15fm0/ZPke52KCO4Leqr
xgq0WEpUIsmuwJwmEllqFy8GhE49jKY6cr8se6Yd/H5SljL5mVrU6O0ypJ3SrTJWwqKTpym0dRFz
Z8TxM6Apxj3q0b9qJsDW+mhxr59qw8+qU01S+7X2Waj6veQVxjFgt9QZGOgZssgVgGubsjeGAh1N
YdWk3uLUrnwU8dh3yipwmzeaINIEJ7lWdLN6Dha2txW2JuxQoFHS6gzab6BpK6O6MGq2c7x6RfDQ
WaOEF91YWayOZAasnsJMhQgiEje3Ir9SMNneK3OxjmIoY2P8bxe91AFYpzqxG3XqPj4Bx0B6Ykcy
lX2oj7MBr2HcNzh7eCaSd0RPI3Z9+BVF/KnCqjqljFBFaqW6H5BEhLL+6KGeDQZYw+QxE8NGSFdE
cdsPAEDKCYaL7ynFhrlaO5H+nvR0HqHMvm9RLKYeVV4JG2g7/Ou7sgcrlY6glCjsk1nLPwNAFW6v
49IHM2b4aiTfXq53YKxSk5zm1hT775blCMWumyZrOvIqa/qxCrvVRU4ej56gn9Wm1QP1/RIuTDEJ
O+/9bsNv0JIZf++8AEFwAz07UntzRzCaR4kDAyzTKXjPrOnjJwzhC4p2x1AzNW9N4t4YEE1kbm3U
j4ea9xmTz7ouIMWD7HeA8pwnH/xfc373rCGedyG5PPR6omUHyIsGKapvyJ6Vthc7vdyI/SuZHEnG
1jQz3t7ZLAVOzAiaLJIVSTsBidONhhumbw32vmLnnh3HSLwAsODfTP3HgqXcXuCzQMCtiAAzSV2o
glid/QdE4M9FOkrrTYIVW4lO6nKnjOyF18fykI/FjNm3r8c7+wISW5oP0Blbv9OfCwuDOF/quNss
GezaxwQBZ4mfLL/V/uZ27emfq+LR6dkyajzIj8MWK75cG31Rt1eFoecxMIGc+VSAnjmKabv/abAw
IGJPYU0MW5ARkkR78/5zDPxOehVOsLW7CITOfgxmHcq8kLMob6ye3TOqMFnmgCFc0qivk1nuM27Z
0vlQVT4OGbA5DigiAXFjKuGcwENpjarExy3DmTcFHDsi0B+DpP9RzT8DFDjONksLVgdt7TqyyiQ4
GsPmmhX/SDw3A2DBY3yi1HWVLR5xSuSyzIPYcLK2o+zNu2aW417oS0EjS6+C9EYnYueIkagv3hQs
lX/E2gSWho158grKzJT3olsKXhKwR4M8aIhMAT3d8cR0KKl+nyrrQffu4lm/Pqakn1gP1HJVC+IT
GiX6H6A3nZeEEn6Y163K3Bh6NH0qmkcxFubYdjBVQb9/JPgh58z0on8jCFXG6J2D4e1FzDledInd
JlvXkyHPioLA8uQ8TWySrVairtZdTXhfYHoJKFOMOM9mPflIm2aWi5Qnp4MMZRPUfwCkOOti38fo
T3stOWqIIws72UeoBGCOljp5M2jNjBqJfabH3WZgTyBCy1xv3n7xeVg/o+s2boEuXGfu7cu85CAE
Z8t8ATnWrGIh9ZO4od3VM7FgSlgijuC1EhZCBjlcGKsYY1toxB8dB6/T/Dga4BiH4bPKAQ9lfO04
hXA4YeSUQC/X2iZjSm8ySk2yTW1YR30hdRXb/EQoV6zI0XRPZa6SQvNZf2cwlQYqeLJuStMaRVlK
e/VNCboAK+A7EyCcFnRAdlkbKGnqYxaKgaJM/hPlMb8YkRhFV7AoTPtTK2KwIr8POPRkbE8+PLuQ
ZLBZ4rg4VXwN+1qQ2Zz8gzYwi8RNdRic+HwdDkEeVkKhxcEAONzANbFkQIiTeAk8BXO/bPnfJQ9y
NUtpX6mf52N/gsoabD0Ji8MFUgKtVOpilZKvcSGnlwQvWZwzGnSVt9NtIkXJKPKNmPz3kvFjGCXK
nAe1zf4KRUXb09v/NM8TyZsacXWWB05OvVYp0KUnhehlEnCDfljXrCVT4x6NOE0INZmKBURC3lL1
90hClTjiUErMWDKgrdFH3F6/L+1uHd+H9Y/bJOky6EFMoNIACtl1rr81BGA2//K30RI6AaFev4rX
g5YEA3Xsfci2sSq2+kixgAwedix23J570F53pAJXBOzrvtVjYFioyNeU4ZEluaKpW/mCmx1f3Ksq
c3F47XaZBRDPYwOPL5Lyb9qNtge1o1x9KSrExlSeSG8mBw4VM8zP++5c91e+Ta0w2uYWTgcTAzFH
jnlfkfNNOjIU49ysN7huEi53sHhRqySWB/XGf+U63mLabaL3XMqGah+crb/G9B39KKF0dS1/SvxE
m9Ot+dDHk2HnEKqgpaafuZ9Jyn/6TnNo2Y9YdSd/eWwIxGGkJZpoThhxWEUWSeBKIhLNvTUb3NGL
xu1Rxt7EERLr2P3I856U+7+DGH8n7ANdARROtzmOdkCKKFlXCIlgvzV0BTGfq8YUh94YUcbc/sKY
3+ZXT9jxT/6d9lwgnR203T3Idc2Bthxw0W+OKopYxZmwODmOHL0QN9BHl45bWHcMtusfcHzz1QB+
T+MwnoTMKqRWz8XMePfrG/Oxosx81WjXKRItgP/APmAr0O2CUr+iHVt8B7wPsTAMysoVDT5XF5Pe
5IHPCe66emJMyasKxBD+JFAHHQWiWxeRq7fRVnk0MYG/cLp3PxXm3cvGsgqvY811oix60QX6R2we
caq6OHfudGsu55iwQe8D0mbvtFnf8AdYYootPCo7Cvwez4Mg/dl/QzK7gS5tDL4FJ8+w9r04cr+C
u+d7UoTYz7CD2lueDV4k82OD+dX9asDLhZ3D6NIxKy60G5yi9qrMHwWHXOI6qaXfxHUPQbUcTH92
7iQfLARPCYMv7hhmzcmjVolWXz3LBSkqnAMTbeoKpx7cCbl89ZwmXXRKMTqGZX2HkglaNAokUfaa
rmTrFZ+A+Rp3m8fH25EGGZzfaWvYMMXvLRD6QQmAoGhBjfq7oTGiQrgf9DNwmFqHjynrITnKBADT
4qO2xW1pp0vSCvsPlIluSL194E/vxOJzEyJcH3INPABzMG3bJ0RS879Z/TAZfyH+Aci5qoca4f57
gSuSzNjiRMzCG/AEWi/9LJgKJ68GIVjSnpgk1o/HlhCssSCqnqy3X9fFZlp46LdXcoG+AJUk9Mur
VeKqv/3cYOLNI6AVvbl1+h5HKc5EXrNBVmL6Vamf2Bj6FP15cLxafsmBNcxFvgoXUX6BtDQJCQVg
r/gKHMgFgTzyAeZPj+WwHbqCq3zXeu9FMaA4BdscyWNDvuGhWQideA3TAaeOdRvBir5KsTLHNUTX
fZ2C4nP/SIgCvFDeLS3bas018IuON0giSyUQoZbJ7pSrU1ngrz1R9UJ3QrCJA8rhNWeS+rBzbt0N
q/YxXQ92TNbO1Ro5ovU/kC/qbX8GLhvET/BFbk08rkHkj4Mo5hF7NdNz1JDwrYESqZ6Wf5sJqJyb
0Ntg7XrNakO9/RsWNJ9itQdKyKHw2dvRka3/7CcJTPhqkXhI5cj4TcBE9x8m+So0pTrdQ6glglul
WTb/NIhTAiUqa101qY5iaYRrcxj3tkihEMaHOT82pf5UI8yqe08XH5VBQuLMD5os3k1B0z5p2odJ
ka29vGJLoSyua9cHhzT2Ba4weqUy9BRBgwU2H0eZx3pJVq4k+m3M1PrDUpU3i+O1xciX2ndu4Lbh
qEjKEWFGhtbIlfhz1fJX0ZBIux8C/MjyZTFd8RZGyuVSYKnOnaUy6B1RwR28VxbtGfO3BZ57Ona4
QemoMJeYASc0F5yrPo3E8ejlMtfVpe8xe5fTqxe68l11NegIcnVQPoePq6hRI9YbU/CnsadkWqnD
jKeeZL62tEiA7FInu3Dg7juy+6F330VqHU6flGUiEL1TvuaJBpOMabPPNoEwmXr8T5/Ef7naLPWA
LpmnahkDuovMqO9yimi8YFINPa1z0if8ufLx2l4Nkr7OnlrMAxJUSns107vsc5jeWYsLZiqgObR2
z7TdNktdFas6VeHTjQOF8h3I1s0tJuv0f70W5R3IcQNVDdh+wMCh2r0goagOiGQbqUk2Ux1veA/9
opSepW/DWti6XsgQaO6g33TYpEIqGuMrS6Wmq1z4Ddf/9oD/xfswuYx9yC+VWHUW7kBMPj1rPEel
uiEatUznm2fZsPMkuoj5t4MBimuldMzoLWN+K9kBkUZFwOnwRFkI6qibYcjqf7YHrO7vfJ6M8Hmd
2m2+fNKRlopciCXEaCsNQOqP9PbsbpCIprK0zdL38ZIqsCcIB6iQxgRfl+Rz7s5gWk6K0k/yW7dK
kWDjWTpUHpgeN3c+GUfDMdP2X5Cz8gFy3gqoJJmlQPyhRHd7QOpahmrwB2t4IhNnDVlhxcnTfoIy
E/GNf0PuBJoWV8p2wumqGxmrJ0khzImET/wluMGRUje0bMpiUBO4qFS9GAZ2fjpg3tTEQ6xIKQcr
Mt6fAWNQclhG49iZUvwqi67HiHXThjZJGlLRTXUDEILpGcsKyYCA1j32M80LaezxjZWvuSY9MW3t
EQXyt45hsQP+sT0NGYs6t9/SN0py95TRZtDFETZqmM4rZA/f7JtW7lVSOQh2N/k8rJDRLjgUCbKP
sY7WosfDa/8aReviFXrIyCuWKP1NKnf6FmtLPkKhGdOTZs0m9v0OIv7gC9ucJ1mO8qDfgnGiKfVm
FopCXnLjJTIePoBx3w4WLcf6BBzg++m1S2fvd7f/UVimn0J56nZTMqWlhAHmufEH+gWE9oXjRTbZ
pEHIIb792E64s8wWzoII7SUt+Sdiq/BnO+aP7HXpgsEORHIo/kja1Q99MTa54KMuvBDVrBRXZ3Fw
la9Qtcr8qI/sqqgoXVH5HS1Vb4d/k5xONWOYsCCHo0MO+qjCx0QfcSDsNCdXgN+tCAO6wesm+WiP
6MiHmdQwTsJmSIUAhjEdQ53CWLptrgduuFwZfz4huW8yFr0KSZJrgLptdt4olnGpzu8Lz33qjSdl
N8L1m/HldwMJtnKhdu4vjjscTZYzVfjau7tHgvmgl1PrYi8+yM/zloJPCVBCRIcPR8JHz6TfXQOF
Y+4bhHknJTALIhOJVDazqv8x2FochrcZY/seaSewqdAz3+D1AeqUBj4/Fh8GpUF4DUQmOlkcIc7h
JUGoJCmtnURbvPDpdWlmYSy+FA/HuIRdKUyiNAgGl1lBY2mq0lx115IF+OZC/ynAs5YUj5HRgrai
bGLaLC+e2OUJkF7+99neR/Dq4CQdIVFqa7mlQF8eYFo8Pyq9tfUXQdz+yU0KppsNRXHrYXvWCUt9
d8MyylRvcoUMgxeIk8xUCBpxDammSCcIfqMY/NN/XM/7Jo6M9LLC1MA1UfPUWOh4nYjd+gSJkeFt
DzLxfnZZuce3H+JnH2B9QnH2AbVcDbLNuCu94MeB4nzg8GVlMMHIIPfg7vI/PETr85icGTCZU2oB
efMOZjbg5grAobXMJ/XquLeMi6IPzzedohpuIWe+gpofPyrLskGgfasvCxMbEo9HUUAfrantlHAo
w4LrK2nGvkVpfQcXPUcofnhXXpxdYipow9VFuJu4AWSoplv5fUkn7spkTLT778kyZ/OJU3ZEL3nV
D316ToZdxFf4WAjlGJs92bNEcgWsUCfuXG1rwxXN9GRWhW4FMtCW1ZgoeD672VoXCUugwlrw9V6s
nKRCP6YAhDW5/JEWf5aOtmLcJWe3F+OFJSDpZyg3EXp4Gqoht545mp1U1jHi4nepFQeIEzaCibLa
fJvcwrwBNVlCMeeUOSxE32AS9c+Jpk3UXZ3HTK/0HTU332hzLzxcuVUCqP0xmP2+558+XoBp1AB2
u7hv4dGIjLNlBRrC97fazEbGTJN+GlFeww/Qsa8jsOmIFpQf4OwZtWQur1UYJMlhHbi6eO7LCH7/
c4zFLbNYDLq+yaoVEx2srhUkNXrLY75w32A6w7vrXA3ls3AuuZBSnsyOi1OeTcGgyvOgijtM3RLo
4rOqel5Ht979qSEa4Y4d5jzYtvtICsPolWhVOQpVyhzKAz0OHOrtd1x2p3OMu14CHSEFgagO3/k2
sI0GevA+wYFA0efnK5cZWgIVeaTRUvkrSihlNaYhfIun2mYlcIzxQjgN8EbSWza08gbAyYYbRXeb
wBE6rBbnx+WkRVGahg8nxWe0ebxqrk+6bn1ZZgw4XYoljS67n7XNOM4KDhSrkvJSGi1oWZYO+9Ok
V/g7/PyLK/lSoy6T2neA5+HerSuffDsArSf3VHoEUVaivTBQWCEt4NHrFsbSdkc6WUjVJhZvfoqW
6HwEaf/vdZuVWD0UESzkuhuGtQAnfpWxqqz80HDQ9NrwJieEiZujsAPmY6TC8oX2uaE8H3oECqWG
WVoGufQUotP00tkEOIqTNN3oIIin56LLwwpqDIy72kHCamB0dbMTXlA7iJX8ZjhhlSWDolJX+dzl
FyT4xTCjmmYoe8qMq1OiSVWKGqhV7mWt0aNs2LX1IYzX1zIWVBhrWpJb955vMksK0RehgQMqU6Rv
R1RexpbIwZQE6RVKcIsPVKCqRYK9UMAViBB87ucsQBjPPFERIHQSHwbGCR9ePS1cX6+OEA/o3as0
F0UAdvpYHQe9X7Xd4E++QRsLO6vq4On6sQgjlcNSR28Owjl8Av4Lxetp1co1ODetNkZWCzeVDQEq
HkBPe3FLZ6SQxAzfnUi2lNCOT1JzlUMpgo4Abz0a5tFJ7F1n5NHuWeWyRu2NUo67BrV/ZMa+MdCd
SQ7COmRYPzKStUSrTSlvZYvIhIH5bOkdzBOhR130yNOgXnyU5VVG4nFcILpLzbSdKEeT66vxnazo
jzz4i462EMl6nZBrE5pLivS9L8fFlj4De/i4PkTG/WqWxKcly4neMfmeQWi7myjjRxK1DuuDQD8I
sHM8C3lzu8aaJyGc7cXdE9RgH8JI5tqUARIgmLW7022AkelQc+fNaqCy/gMxW+jFwMfIEoYcbjLh
LL6kPVmW70hWG4FXJV0o9K09DPNURPRBU7YvtHr3HYTHRlnuM00+xgOBZJP+C9x0/rSC7hXFhnLC
VHDux9ro0M5hZ9fBc21KM7/Hqd6kbIBjr51cGhbtOcYLmXHYk0AmAmqbc2IDJDWzOvLXTczj1VEz
c0ij1UtlVI9PvKFO2hh2Sx7ElSLONJsTn/oIMmo//Wtb/zI6WPxKmXppMLBnKo1UhrS2Ly528m9i
HdqQNsSSFn4oDbhQZH/BP89oBLBTvLqLopJ+fn86M8g4/USLp64GETmrtoUKLIrWQU7VP2dUhqd2
GoIjB/nF2Bm1+P+tyMmRkehmuYJOlUuJYK6BSoVCSWY1/ugF1pSm17VZ/O+wU/cYb9xMvu6SGeH/
Ixnduv1u3vHJfkSWJzhspDVl5klPkqCtRGsDoixBGr+Qe434EVdiJNTpJeqU9CKdGWn/j4Ympd7s
kub2dfOKQ2glX6RspPXWF7xo2AAd9CZpMASKZW/ArflAVMUohM+KPaDNdBvmS/iBmK+M7i9Cfoj9
GHt54+4wbj4/c/+nLlM4Bi/gIZUm/NhWqrFPlLFZWEHeeqcy3A8NtOAJ7TB4L/vjyVAVcOTWM9V9
+qMSUU2B/FQvtZziqJ6WbRwE78bIoj0O265qFa2t2c73CS1xAyqk5E8qRslGbFlid36cKSwB7zpp
MhRQTCiQB3I9/CctfJLW61qIU/vg0naVSGGi1KsiTQG900tmRZ6IwEvivse6baiK6PvkSZr5ycCO
BTGoyOaNHOLPRAXfsLm/xf9Ra1X1j/d9XM80mrB4aQUoH7hQl3p0Tuose3Tc+1JDJkxXfMghIAP+
qlJsZmKtTrEBYMcJ083Q2tThrwQeKXDtuRr/UlPZ25IuYRTJp2tShc68KS9dVC2I+9m1XFGbp2vv
WO5BvpqJTuEt9cSz/97xbvnpHXP+MxX+iESaFSSMmL2/eVnIwqDC3PiVA1LoHMqCCSSuWi+rGbcg
mwyF5Ru+Z5SYwLP5jdrxeSAAatQfvwvaeD6SV61/GjTMUzL3DGrZMhx+xtcWv+QCEOmFYivK28sa
V4uDlOA6D+B/wrlJgdLwczjCFvzbsZe1w1PwcAcZl0cXiH8S6I6redf0eUe9V9EP2MwjWJhVM/CK
1YCqeQfKuk3vzfcuKqFwB/W+x1goofCXm8ioeiJpVTrLcqOrC+ZtJCEgtMpdpjO9VylTFRevZz7N
BwMnTJfz1LZG8KxIrZuAcRDb8KmJBDks9Dv4wUnmuxNxRaX7mq0dhgWnNqk7pyA0Eh0Wip0DMTim
kClhul5YWFKP4O5H0eL/T7hA/UDl9OXZNaerKRu/bLbgyK+foVxMZ/++WID1R6fXpLnvIyxfpCYD
1FTt7hu6nptdvArnQ2i7LKZ8MkKKnTRv0xGBoQkNzI74hhH7kgaSXSkoUpRdDD7q884zAFNWlFLU
7+VY6Qh6yKtuIexVobOE609eeo9SOGwGvACJsYjmS/vtfiq0yuLp1Up4695/2Oe8+ks6QXNTiosN
3wtcesmBCw3y1jW40/U/Mn+K6GR9CAHIkfTUYBS0e+hWT+vX/F4D8CCgnfDbVmlNXGPz2EVD4e1R
PcUS7ypSd8Y1N+SWSLPSmqBqW19dSoUo4GBdRe88NF32ORwS+yYDCnR8FRrmb7D4mwxUCPD/+YlV
efZtshGDA/ceYGl0ZLTyptbJLxoHAWMyJku/oeTua0aoUXfvxY+sRsQGIyDinzIl27FVLSwT4HKa
pdsE+cCO7Xn9QiUiheGE1gSLp80kwvQG5qrqaALFUTRHkoZ4d/wUXywaaV7X+ScspBrmy+KqbVOV
wfpAysqzB9M+ujf0OYU/bn1xVn34VK3De8DGGEC7ONrlffiyljbttwV2b79cTgN45Ysn5nibjGf/
1wL3QJyx5nC5TOxR7Zcy2R7yitJR7qJcqcH+kk1JCqNi+2RO+dRAU6VWW0C4phHqF8GvaNE2cdhF
bDZ6220mecZ+4iXe1bS1MTerypaCvhXXkrKSNzNuIJPU47XlmNJSkrtDm5BOUGqTAYfuMzFkd+5H
1fL+LIjGqGu55Dw+Zhk7BJ0OToEqot7545bdCL9vYI7qnm5vWxdmrUy3dMl+ZbpU5lA7nHI+3GrK
tVByhlaK7xPEkk78+bPgP3sMlL8VSL6isfIJZAB7lIaZdRGrh0m4fpuGPbMbv3ZH3mULbM6Zkqi0
3qy0a0Jx2kfUyyeVjCSjjgcvOlkUGRADe0RbTAX5PALsRNKptY3fRWtWX2q8+1Tj5jbwTMPi5EpO
L322h2Ck/JJMCxeH3WP0JSIAhQl+uextrNuZ7WVr+AYPkS7M0BjgGZoQHoqzSA2YEitw5qjG14ZK
sG1baOqF7UH8CXvR59ZMFA80vGqMUHI2/yOYqX2fRYMwfIgIQa7L0uUUcUBh1G/MZpI7vIsMxgcO
yuGetJcJE43Li8A5/WqCKF+Jx5fwGaVDuOMv3437wV3esUfpeeEmWIyFzaF5ndoxoHw0j0wvGDP5
bi2fVw8bex+gq2b17lLIvYP4rXmibHuvpWd9yUWLz3ThQpyw1lmY0BMHwuzObxmMKkselTHs1+gf
z/8OmxME7equfUKUal/FclkRHzz6H4V6QaPSBRUphzJK3B+jh1b7sEn+L05j18R44Ssq2CQKZeD+
LJOB32rbgZN0k+hQG4sWOCpMZEVC8I61FVreRIcdYm13SVZJ1HsuOIWMl27PQe5ENwcgbUc8Kiht
rEp++rDwROa+eHlXyZ0t7tzXZp8Zd80NDBZCEoy7kt/51h4fxAxU9jBL8AJI7OP8iOpmiWcgfU27
qlLmsusRW/bo0jELMuNEqNZAktDZr6MbXtmXhl1D/lTZ455gGIobbDPgasGk9hpo95wOiAOg9cs0
lJBqFHDB/87aCib50Om6E/0h8YgVQC5PM3QnG8x0TR/dc0ycZKanHMkChoUFjjAhp02gxOur1egm
T1Wn4AixnoFAXem4Z8s/ulkIi+ryB3TRL13+t9xGA/j4cUAPEZlr6p4+CldXb71eHV4Uf1RxCDWj
CfD63aJNXHTfqjce+LjaVzww5cS/LcONHR6qGA2k6qaz5vSYgIDUmCLgMPcff+qeTirHujLnIvdS
ZSKzHikoIXuVMk4k577uFpONKtm7pZbzzWxujMOlweXiADkglTdkJykrpRLIyzCGii9eg0rJWzL2
09wcGSncqOWO1BERo5zgNqqEfbpih9c7XRNmImEE3n+i+4wESznltEtm7e+Kcc8F7ldCaj1f2Vv4
RcJ9zwr8p68xd7KcPK0456kIQ3ocqi4AW9LGZ7p9PJROUiZbR4jAVhbnRW6IENuOIyt5PWbLBfKE
DIsGcBbO9UN/M3pSS5717h9NZ1EnM1OMEXwJBCcgvehwtF0vNX1lR1gVHS0lJ9/C9aP+rttUdgkV
GG3QCgedXxQQg70tnwXFGXuh7zqlkMy8OvldwIiAirY/zRVEs82aYSg3Rbi/2xpD79rq5qZvsyZb
TKftt5Egu/ZwmAsaKd/ppPsSqR3PnSD8IMuoydIROXfjeBXwrDqEVTBhdAnJ4wRJiywkp64l6o42
c4zMYcbcxHGQ41EGYrixcAdBLA6Ya8bWeETPUw490hQ2usZ9h3L5g2P/DzNKuwYoLJPJdbTMPASR
pKADaMU7MkuCqN/BIlqvetz/7QrNpuyCWwfo3soaXScLt0RQyYV6jBh134Nu3UFxhgtbhNfRFI8F
xvyugC9dCXfKjh040jDlVBp0M/9SGaCqVvd9Tt2nC0Cahduc1l9Q6NoarZG9nkIfeK5p4cvo8R9g
L9waOKWk1QNNpY6BbFbwyH/AJZoor7tjrSZm2IR0893US5H8Pc8AqnazWj4q4jljLYkfYJwwVkJm
8HX+SESHtJ2PK4pWoJuS2c1OAN0auseC2DzX6OvGA8DY+YYfRwLW8EEMfDh0wmZ6p6R/jTvAXrKS
KpblbFyD0zrU7nEMAZUOmuT8aLZnEbB+ThyU0QEtNBtGs8nH+ZPUr9YaP0fz3JFzl7SMbFgyr8TW
WSnrgnDaAst8zTXjAi4EdZAoK+TRym85bPdywp628CMryOPQFkiaXM93XgKCoi6vAoYOrudKdyia
JWbWyrlZNxTeAULSaK5R52838WKF2uwA8eI9s5IyOB0pbigsv/EU2juHr+OaiIhUtemHTQQ9Ae3a
JfQm6fsh64sAvGU1+UOx0chc2wmtox0QL2/LnbOtGamnxEWma7Ch7/CBQMrKWcgs5Q10hw8Pq8Hr
0vIxxKEpL5lWwz/w4AjH9Vr+hZZmJxuWobIGPzau+Yc0HXWrxix0MkdUE6Rbprjlzl2X4GboaqE5
DiVt4c22E0w2FJq9XCQCExgDOvBqji5MB8T1rlQyaZ3DPzgsCyGjHB3FyOkxO0scYU6uiiHNh2A4
0iMQCprtK5P4D5OxG4p47m4liLjGP9oRNjhdUnBG5OjKTVIaQ3qrURJrDarqwoDQQ/39azvfVpH1
kHcV2Tm1owD35hhD8s16VyIWWszV7P0oxeLHQGyJhqX1Ll+fJ/AzS/mYCl2r3RQcwjy54hFSkHYe
+uwKdd40TG8Sh76wYWx5yn/f0X6akF8aX47hwH3Ec8vcKBH32SHUWPCTg2q2dTncxsYga8hveOI3
7f/8G+H3wb+RfwbRtPqm8GQQSkrl2WVXpE7AvUfqVkCg9hYOcE8ZzVUxNK2e7aPbDPl9gthUx3wL
hw2YjcsLqMwlygJ1t6t+iRxzzKvxoqJ1QEPgImV4dmbbTjv+EnUmBk/Wef4rUR5cSzuWyTrawj7w
wJBC7CWCryPJ8hKxsxnSREKBdGyHuaXdh0HbqqvWe+mPouWtorXvEQDqOwQUN57G5KkoMaxd1aQw
Grfkvim20QJYKBImBlStDEekwqyFWfAJNQLhP3ut7udHeYCPCMEMf+twrgLf6QylgDnBwmPwDBnP
hEhGbD7mZlxNDhedLGPSqjHEj93HA4B6I+uTC62szHyP9KHos8zSC+o+n1pcOWAPFGQ50ky6vPAp
hXKHnyBFNFq/EBzCTKzNVgbBrEdi4rAfQ0Jb7pJLGcg6vGbgEDmmUD4mHaepkWU3r+cxCZ37e7Sm
fetAK4BTOSHd334CWaltglvzdple1m+DbzgrhXFumesHGbUv1b9OaJzywN1AR1JaMI1kYQ6tm+5P
mqAmk4/Gu6cdZm7fki/QL0brcFU1vaIXpKH+AZWcO8Go7Blcki8pXOaq8vDe1HedO9XC60F2AifZ
GVL1kMm3Wody3RB9mwiqMqutEZM3Rb0/dhzWfBCY4043s5jEy9nnfV0+Z3TbVvGp58YfjNFiIhlE
fBXyG7Zyw7XB8rOIcn+KzVOd+KkjZrhun96CX3TYf4Y12k9wFA+0j1hTDSb0gOoAO96VlCdu38TC
1bFG1TpI2CRbdPcmLhdxnGL1VPOE34xyQhLcfAEWbb4Ky2h74oA39skLplIggCkZQo9p4eHDlMDU
rvdZOTfZcIe5ZHetm91TMeVs6+57XgTml3BO+ekfPCRY6kX9HDvtRfV8uohaG4OmbjLEdQy3cU0+
MAuXSDXm23H09xbaqWWGxgDfr9iza1MZokbeQXtiY49iyTVzYTCuG52FhpT9dMKXhzDrO4+qUiR9
9Ew9fof4E/CCRBXGGIOH0mvGx+5h20jfiFwfKFANv1KamHMDXeRhEltO3ztkusotxoYgPFo9tXPJ
yVBEoDbvq5jLid9J5XSYTPzgWn4RjEU4xQSOhLrO2jGBpQgNvHvfKpc9mI9lpLxkbJiqc97NDZld
476DERG7oLvff0HFMLrpA71YjOKKcU9S5NfUzRxj63AyjOS6SYWsCGeRzQNWsULcXcbk++LbVym9
lzGARL7wYgmQUxgiDDK87arceTn6UeFF5g71c5AHt0c14ATwVh2NTrWorY6KRh1eZs9yACH5c0CX
HxbMfPjWUa0kVuHRwRmqScyisQw2Is5c5+rXHZYFF6NlmsVDCyIb9pjltjE/38IuycuUPfqfsWnZ
UOk2N+9ANQvHwqKaqvrO7BrhRSSrT+7ySImPyAPy/2wKgRHp4VVe1PSvAi8dP1h4WMArccMAZv9a
2c+U+HRODzfJyHibWyf163SEwUNFoAOyMiwGhzhclbtd/quHJAXhMduIerz4bTRReE+Oy4djLK3L
OPYeG7sqxZioOZ7yAb+h24aDkk7cPahdfYZ+I31dPvPJKrKpNBMGUqm+VjO6hjN2CvJOZBBiE8H7
Nwx+L+3tAbRGRXfgcHQ/wbQzGDWGDz+DIg6jaa+cWiOkGnv/T//jB4uSqL0HwTE5qBjyjKXU9Ir8
QpEYz9F0T2eElTsnpi+/RSYVvmZTqNDtyodCXb2H3RFPFc9FPElpJdjMqJDSkYgC6mGXdEVVRNs+
USrY8E4wfZbTtPFwtVL/e754oiMugjXQdZCz0SDCkI+ah/yKFht9p73OfVa2dbUFpwzhPht89ZsI
DCche/jGdEyosdtuy94k4+gPy+vWZNugyjwpQDO9OwmaGKOleshddF2t/FBpy+2ocdMYLhvA64ib
t3eUVT0QlrTn1s1Yrf+Mp/b+Duhuhv4gNG4VtQwiUOt5OGMrBVCO+wM2jhsB4TA+z8RVIVAjlQXu
fgjnvToXKmstike88XGOrtuNCm7CJPlpH831QDpXnXsmJCFT6Tpv9RhbzlsYd6fXx99+GWA3UJSs
OQVSfVVv35gSicT2f6ivsXsSkRzn8xCPfiy5k+b1hDEwlv6gNibeVMWXu3lpGEFDQBwWOko0NOm4
mNZdvUUM5friMFFcayp0pIdMKsvAtJa7yti+twaB0zNsIzJdYlrzTmyy/UTn95qne+u8GQFNaHHm
uAFPp4wHTQ8v5Mle8OEp7D7oXCG2ZlveKR9Y/NqWaxCh+AvYBKWNuaWRgCGQKQrNIjYKK/cNiEok
9EQ+i5J2b6Y4sxoLNCv2APDatS2xIYaQVRK35zY4HhV24wxO+BPYZeVGKI/FPppxSLW59UQLT6Dv
6Wzxk6QhORAsZR5jN8PzT8g1+Bys3cC6T+cljQuBtSpIYOVlmzrG8DMLETVMVxMEkdr6vs3jy/yw
EByotsoVkoF+KN01JpT8eafyWlf77wgeCvV04S6/eR3NhHjADG3rq3W9ktY1J7uR/ZUNzSfDWzee
lHZVBZUTBYSdbk8fmGxkvXxVGFaks/qBTPLg4pvlnrnaDzeoWcP388093yOFsjgFADTwDmIRsxjP
rSbHys/wCsW94xEF9mOuAaR2tQAsW4oGPY6BTvE9EUy/kdtSdhPM1ikwxQlkt/9ru2vYj0oLoXco
LHPoRd1W+UE6AA/gDBTQq/l//68cM7U1sAHo7bJsOTh8aDsjZSE/PpuOgpALsESCugn3oj2HQFoa
hxZM1sRHFK5C89X4VdjiJcU7jZwjaaxaHWzy7KkRq8WVOeEiYEBUCoezcXXvhKhxprKyPkSGDWKr
bIpXzTbJzxnrsMTyHjPOtzTD3uO3j05iygk55rOEuRsoGotBGBnC83qPTJwO8Tq8lYAhQOnWr8tq
O/JzC3hxsP0SDmSWpEkaYATpuxY0jDcWlpaGHnulhbwExMFQmS7eC6zc+iLLXSKCx2/tvmbfsdDu
u5/8u4bphdvm0/uELKacYRFKtK9DzoJV4gw7AsyuccHLHKGmrG9QwKTfUlT2PCxTNfsdMGWccSxg
nDRKyVh3xmX1HasAP6Awvlk6+o8XuGNCxMQZVWSa7RvtW3q8mjHh6UZ4ZWCU2bC5nqS5pBXbNHeJ
slaEx9OtfSkhZD+G5CxLz9R07NjYDi8MrUo+NHleqoX5tAyWt80qINSv2t1V5/yEvt29hR3/k1z1
oJfoF+IZsS7shsO0TqHLDrFl96jOuH92cyTh/R2/kxjlYdUB78JCtaeacWhctZKkiX0KDwHawE1I
eDXpA6BSxk8qUxu3JcG8muNONqvdgznriZjKCjCKq0LTFodyB3fAQKhVXZW9r0T3la6PQ9+xQQiY
QS7Sh6OMDTTIHwR52F49V8AEC4ivQqm2fpM+GXuBSr9uwMKOZwEIfnlH9YD8IEgbEMkKzSOfs311
6bqA1yIAkL7m3Xy4iG/hNnwoNJ7lUkpE/ufL2dNv1No+ixq4Y4qHxy2NtInnm2NQcXnMHUfeUy0u
2vAWXkYhvLyesCNfNJOstOW9yJQpVNeZiLthRl5QODaOcXPWGd3mmW+/+AqU4/YToJqRAkjtUvFC
V8lF7fZq6Cp49gYRKYp9317Kpq3fhVOiUoKQOQ0WqYFjqP7xHFRJzfBDQa6DPB1CGgW+HvV/xyjD
rOwHjJSPcZ5O2GGxBv5coCB+5HaTe23ARSiLdJCemOQV35davVzd72f/mGWx5j2IQdt7bBRZq67G
pDh4TPryWEHpQsIn8kABNXTjYva5GU2tq8Z+WtlMzsqJ+s7wAuKH2td/AWSEMnv5MBzUU/E0Irla
ScA3DIbwulrz7/NEgDmxfft2K+cgpB9urDOMOEKnOTTeqb+IuvASUJnfBB/a/FzvJ+Z9BExGaXmG
wl8W4vw8hLqLHb4OUxeczkQ1aFyP+amMwSQ5qL3t5egCFFn9PsGQSFO3wiLUuPHbWXZrHq7RP9oU
vWVIJqGdLiO/TxWexsg9b2ZTqlFz+kbdzfq3/CuVu4rDjsQfBDaP+/qErOi5eefyYt80AbuNCcD3
tjLRX47pYuzk8yufaJTzC+EsuCjmkeR/fpQVZUCoX+PRxY5w3UQl4/aaafw1+cOp+O1lrkGSH2kP
AI9YSfZR/cpLOF9jyz3rQrQV66YgpbaY1u2umJluA4CC8nPbRlaO7uhF6zIMZCoCdLptabKep+Ax
Z6Qw0qZJ66yQNoLXrEt9zBsbEPoeqoDIb2QtG4UksYY4z+l4rsIDF9nA9Lh9sTSDYA5ACqe/uarn
z7W/b6AuPDUGgkodW81HztkNd3KaCPQvmMHLLLzXw+huue9maUcpvhXAAH2EcQ1PECmIIuffeYvc
vXxKAK+KPmUuAEV7qS9EfYram/fWARKgpdrrIwHRl5j/aVSUCZAKcvSXDV9jKHmBktjwXtjL1Wq3
kxhbuAF5hJHdK6gA6UZ4csfQM6MgqI+Ylw5M5Zdr/pQxzb8rJpDEaNtTkbMa7Q8nKTwgCb49+BDC
92pD1x2LqAtY4UKKiOtTK8SJ3AKcTlyxqrzUbprlvJ3C4NPgNqwGKQDK+aTLwXDlYhsxqDO3Sax2
9nmsysLUt0ldkzYZ3Xu+KWg/5c+4GWz5ZJj8TK6fPmykZumHebL8k3eYPBMYA92VG/WNauYqdmIo
xSzbKIvcOjsZ4dnyB+LEdTU2Le54ofnM5dO+WkKKMarVRwVwdOX1wraQOOQhdMy/va4q1pNUmC1H
DOHspkuUgWLyFhvWKrOEW0YTVr/Coh2hRu+uXq8OxOdORl4S17jY95lkRL87kE9rFhaRayATBml0
7L+rXXryEA+6Vqn23PclRNPIvi3tr3cUbsiTI5lqCXE5DAhQ4wvCqduAeywGX/+imBX+QV8pAgAX
XH5ekW275DH1uKeKEBZpXbrzQWwX6+N09Ras8iu4p4AllfOZElRKVqyHOEHQFC356m6PDIFtkNmA
mx1OCUJVLm5gjHMFOp4T0IvWifD4F7xAHzPe/aCVob93wpwX4B+nVltafWhWhqiUIMDoz5paH2/A
jRdD+LQETEGUhqqbkJ80EWwIZBQou+CBH54j8Y9KMurB1eNSlG39Bhas80qr7702ZtOLN2aBJ/Lc
3n/bswAAtQLM6uZqW8/+imte4rAivIn5DgMkxfPxPsqVYi0lnrhKsIcm8hLIXvNZvsd0+ro4ftU8
Y2lZuBXWOOHz6aOx0Jrq/KvuwrGymWvBix+7UN7KokUz3dzO06ZSYBvdTM7q+k+CUJgFzuaFQCL/
FyVKwNlhPM6QdtCs7qLpENpj+3N8dmLCj7tlfjvZhzQmIw7HgzW7IRNkvvD/SWe6H4oagvgWdbck
RbBIJXtCw5Nd7ce+LZ1WqHfN6QxcShXClj56idsHszLA4KkIbCTJecnUzcRyMrjlu9SJ5w9Llyr2
waBd2Tf6NjZKlzwJRKS1JupGhl3Yba9wf0Rmv7QljTemWNunmOOVEyfv8h+2LnJWZv8mGPw575wv
LTKFvS69rcP/q0KY/KmBPzuY7JGyEONentJEXOEsfSzi7qSmTHg42+slZHdY1H876CegU7O1tYQf
rKrenjyjSwpsMZ32J57yHzhXScpvLZ5evUP8P+N4VK+m6iVUNyfDpxspk3qm9VXG8tKetupsu9ta
e5q4yLkO16tB8ZtYlzR8K2c4V6FnbO6/eaI0QDiWckrDq70ufgOmgoSfuKDUzv6TkR0I0pn8o4Sd
l2wBXami+1fQ0PvQgkIRkMHIyAFW70KX7lq+4Ak5TJ+BCRqqf5K0xnqpqWLmrRfirIda7Gb1NWqJ
flaiHaEjBGyYFglzdXAh15KxeEgJMqNxtpUelMK3Kb+ohKb60cFI+dlu73pGGRwbaRO6oEMkp8z6
M/GnS0lZFcWXCywJTeShlvTDLyiCiu2NckXEjEcHd+yTm8VBufJ8aI4LdIoarphUgFcvDsBZ7bOU
AVoOFo+MG9pvK0iIFpogV32iytF68NF33Q4BCwkpWG+omDpndjxF2llfYnGMaPiPEEbkWh8s9ukD
yA54RuYlP8KuSAUVxuFO1T//lmXaLwKQC6Tv4bTzOaLKbTeymTRw6TEtRNapA/md+Wyc1on/9Eh3
7HwBnKcedbjZOC57AOdFppAnANse2SW1WdWCd67aWak0cqWundZW4Tw2piK2zNbHQE9ywqXuUQX+
iUZ58CapaW8uxHV8iSWaXHyqzRTH1lflsFfJxDPtJay6f20Xs/mYevB2peUNrm/MWlrgjfR7WQVm
fV5U4bGdBogRWtp+PXt44y74zzZgMxr3yqvY7zFc5xl4z2iGK/GR6HatSIDzN4u1IZwhPGXIoBwr
EES7qdcMm+CtoadC6ieoBRulLVQ//A5ys/N/P6A9LFcvgEb75oa/wMymPkpAGCqnQeBy2nOlTzS4
lxVPyI4paiRV0Ej9PBqqHMMzKXsqOYg4t34jKzS/Xr4mzKOTmgWsIAh7cx/JNV9UDYJRXXyFYmxD
+hfAkgMNOathV0sztqCmr7EOhx33B7hArCMdYimOyw8YA2oR51FUSvQkrGjlGyy5v2M+2ksT01au
HYCW+kzkF+DkK8vPgwi6lvdgHVy/xgcanG1Zj21H+PaiwLdHm31mRMvyk0cWC9obO0T1vEnSuDCO
uf682GoQATUdxYag4vvsel+l5i3juaQlbxnYOnRaMAbdTCHh0vDts+TxlkS7ampHdJEEb7o+8gbV
7o8bt8Id6Li1iZ5sHvLZYJ6M457P+u0mUNA87qbeC6KqYdYQAUgrEzOw59FOr0Cghz9/E08wWWeg
DiKXPK3SshzL4cgOS6VhMXZT4dY89Y8Q+nmgSFUAxVpzgBlqLatlJ8Ii9rV93l3gmV/T3goxwiwU
zjjOCVsB9wMdukAieE9V0E1I6Ru8b6LOKxjL1TgRQEjT+Q9FsUpPJg6FUNfdCbeODjIkqjjDUDSa
ZRq8rz4Yi4FKTvwQ7fvdYkObeS529QSjZivtF3kFuL8WR0EYCWkLAf5qzmvEUcvrVzOCXwI9b1Hs
llkj+mEW21NZwVxH8V8KSWG6xrMXbvJmcf6CvqmMIlPjX70kLKA4zgFd+OL0NZFvcYyDhxHoBnmy
OdXcX09bEc2rsavoHDzqf1RAVT/OdEfsTqD979vng+8Xej3FC8IwfHHpaRbswiUesHAVbGwhymat
yXKIwudFOiHNAmT/T2D8lxaJTI4lv9IYe9yH0Un0SY7DuTHBrBg+iyIkQFfm73fhh+oM3qg2xKLy
4gwBSOGxK3aJY5ZA+rOHQJiZt2Hu1LkxJ/Cp1mnAZ23+PiahY5wQHlqTDWs9SvQPNQiG8Wkbt9y9
NhWTLVMVGAH3vte2/eWzlQ4tFqASGFbTiDnFUXrt13k219rTNTuT20OGxnov+aK27M6EsN/+LKtV
yKmPTpqdPutwq2xCdakldiMi/E4YKv0nb8foqM4KMgvbszwRj4JLzQ4Ax4g/U0JXPmE+kt3QoeUW
c4yel02/OOBrBkqaV8S2fjsTp6OYqeRdXa8x3wgqdcTfKjTTLTyjc1jvtFjSk2qUJLhWDY/hJ5Y9
zbOLBvxXgYZKceiBA2NgT6qWvMDX+uJrm19G+Up6348A6k0Pxrk3SKty8Rb1mPInqOsdGb12l6lz
Xeq7MUPqRG+Og0KeJvky0gsB3haG7Q7uMgaXW2jz4ae3e9LCK3Ju2zjBhkMI1tyyyKTSxqHYT1GV
2cxCzy2ENaf6VZTqZSvEUxLp23zdc4q/P4PHgTfZbFd+0HYiEhOmdWWo7OtShL/hbyr29Yi1DYx8
+B3lqTxjoeKg53yf6fFrgoa0LXtK4qSF0fB1zclgVYdOO7krWybZTd8FJLH7z99gVkKWSS36RESl
rL/f4LGbkMaLAIPArmA+MGAZptF17wXkNdKIO3QJuKoUqFI4XwWmZw90KyVFSFFEitroV2hz46np
UfWjIalU2urEwRjfF4VATFILheC60ty5vYzcdXyYM792AnhL87IJSP9gnpGltrUliUf1W4RjrSlP
ZcMem+NLM4Xf/XFmgQCH663QKjg9Uo9V36AMUwUCWzKbsYwVykuFnF4CYPFxn4Jwws7y/YTs7pO2
S3tHKqRqr0hhtvl6Vu4akV6kIVDwimGBKZtNAYWS1/kup9eiSrJ/WkPs0971DVnqIEDMBfCeBcp3
SekefJ5ik7pcPvITU3qXnN6kR1eTGi+ukw14l5efxzz5JSVzPJ1RW0jN3Pq2Djne/v5afoHzRvwB
05IhUvSkcenD2tG3nmYF+OH2gfQnQBiv4OZ7jISGG8QuW2Hdbg2tHooNh4FEEPDJ+LPLgy4C3kE5
qYp5OKmWqMN81/FxE/mWq8cybDJD1SS/PnOty8KpxHa377E9pr4ie99CKmML93sfprdS7rXFV8+4
YLJFQoKKjp7wZ1UJ2R8ZNKZoLjuUmNTXaKKOC6/2LNW1KZdRhbSyua7ccK/BqUJOgH8ElZIvfUey
KAN+TTwWe2pQlm1cTGT7KmJI492+B7uz2UVt0EDZnxExZMt+Szu1L68zmyOEv000N1ZQ/ajswVD5
W2jVvfO7j96bM8jnbSxF7+pV7uVgG6Gqk0r6RIgw5i+zaxrbLSgQWvaKvYJT9rQ4Gq6DUekpNTex
BIXYE+N3F4QpQaIdzqXQYHaHEsD9Xq6ALzgrpYqsTyJCfYNHiID9EsuWA1P0pmf9p4JQ4oJKtToR
9lHjeDPvqdWBZkACrr/dqyhRZusflIMgqlszYyonRKRmPk6t0aY/PNsebisBhwfN0J2iyevTns1R
8MVJviGipRB+O/RY/OO4REqIiG2HjBbar+desX+UMQT/2ExraOMnSiRwHg1BPCkFAUDtswLxJGTx
Cw4FS3c8I2U+S5ldUCtrmfTmRizurrbIr7GiwCvwMXKvrf1nyYNViBpqTxdjsoNJAFNd+NPO/GNw
/uuGCVQt9/l+fsbejl3s6SRoCfruEpZDEVkh8mbkcyn9IN4U75ZKZ+XR77eg0hCeh5k0CJiT/7Ew
yzTWHrKKtUYYcGXXtU/PBaBFUTKa7UdqF8VJfsXTNxgAWChN7zrge1VsiVwPJ/zzsHzdceUOqpNt
ITW2H/DUp0YNjTNsaHLSi733lR22Dgrr6aDBC3471gPqwS9B/SV4obp0XlojPwWEUHlcCKFCEq/w
lDlWex1vhKZuqGUh81lZJ3lX1FopCemdZBS/rZbydPv3NgOIPkstbX4bV3oE5Norkq1alR9sY7Sn
EcUbxD4VX6mviuf9BxqVYnkcDqLhs7szzsp8lwvrUsZVxfVZjPAtJBePxBU72druNYrCyf6i0HK6
RFJskleDnhXLlJV1RycRSGhGfsmmQpjaGjtjMBe4HtWz5sHxdfRIYRw4cR80koS4MoK8izsbY2OI
ZekHag+F6BaOuK/zsvXfnpy9qB1pJ11lPhbdMd2VVQKkLLZ/3oFLmD39YBYe4SHLiDcls6oDZqb6
DrMnn8s1g4BKfyvaYPq4I41VTgiyX3nfW6sFxIP3M+E8vmdC8um21aeJW0Y0WddAber383fRBihO
k/U/cw5yCrRXvZwLQy582BXrod6h4yp0B4cLgpA+JQGGiQfpIy9C3NfjAeS79D9nbKpamOYHVj4h
7HdeztML20JRG7JemABD1fliwCFVqf7+GpdvzS6FnaYp4IeMgmOi8BQlZLcegOyQXzdoz7P1FgzB
izR8MlEfq2qRjWvOYLwI+yTS1JXks57Bn+/2ZcXOsUHPmCgJ8PMtZvV9cBwzkmpcbnquPx2IRjZY
n/IrydgrFQRa/yzjBRhhC+IMm1igea/mLzm3Fpmla0Y4mkjtPucfwQy4UZPrACxYBEr4fhpbhimj
Sy2T1vyc7wdl7yAlHRdRxKAifIotD67e2d8bte7bKihyb5b3sBon9EX61UXyPuyC/zFxWQdPrCJA
P6V/2FxlpELbaD51ydue3MAr4041jT75MRmaGanqnDhSmxFppc7C+cTk0qcz83n19/ef3Nj0Wroe
uY9FKZWRnze53MYbTezlExxx30s7wFd0yGkAU9/N11XwL1cmMw1lF3kILKJv+MXC9BM24ggeC+3U
xq+mfj2KGN4tA9vz4sSi0Lb+wo1RZ6Nk67TGykUdEW+YZ7wG9W1wHd/5b4dHlvrlcS+06+i6onI0
LcCEmC94yzBx4ojrDSFJ9E1zJIZJkSxBPvno9CNLd+MRM8yo2Nf73snEvnpFYwUAFd8ANPwZmiEE
liw/Q5xtGROenX7bbahC8aIRRz1oGvHpJLxlXsj6JZxc7fvIqCaA1otqcsaWI/O4ib+gCN5hCU/M
8KiGyWSI/nHXalpqeiIv7aRUmHleaoRA57XAJ/tV2I3POd3/diFB9M6wgImiCJ5OIg9gNjdhSbIB
+WFNZUygtd1mwpARpaGAuhNJfstfkaLZ0xkQlWSEcuQTlrGcgwzs9gNbsGzQ8xG7YHMhdWvunGBI
xR+TzGEbk7gNNJI+s87IAt2SZrjWYv+Og2s1/8jkrb322d1Vnn9xZn1piQw4a+rfqFIvkmZfwzXo
im7nsZDuFnL8EmkJa+CheiWeV5mS4BkdSpxy1H+KtKH/lJqEGQ02j29T7f8Z8IZLjxEoVZJmA5l6
XvlTV5j3n8ufa5j38jri8H/GxFcjb39AqY6Pab6uxLrjRhB6tdpKlPnIX1eU+a39dmKroiX/CNEf
a0UoNZnh0YjLShec2SJ/6Bhn0bGZx7IPXM/fVa2EdTYJDUcCARVvepP3aTF3+tqqDgf6vnStTnKw
MjeUvui0Dw35MDUm+fD9g0fPcQRpvxxxZ1ihxVtmorZzT18aGk4BHecK44fjHQY2od4EKgQVRt9s
9yBzPdVyUSFXjV8GtugbSaV3Pw63hjhG4GrM8kvrn5vBIYZN5GJEcVIVOWxvtx5lFsMU3HFS7OFs
4hQmn4cO/KniySdOAfTQwvTnZEoyphmsmtD7pg1n4bhJEpnrxidcVzLJVaHuld7urlEofOIYUD4j
F0jsRR9CbrGF9Z7o7lGPsbpQ65V5U+V8pxNnMAXa8YCP4sDqphUIMCOL2Yu7yEjnpnD6ROMEGzfZ
Gzsr/y2qWdXxFldaPv8bz4TnRlmXf3jx/9F01yn/eQZyU8vTpetObqeu6nP4NDUA/wC3wze/Rozf
Gk/OF0c8oIB7vUfcP6NYyHL8DLvGFHNIGLK6aEkjghVMooYPl10r/iBESiRyPIiROlF9xXG3L25x
HGoW7lntqecXjJPUNyvfHfStSegHu7bkKWYsspmHuYkR16BADpZQt6gY+KBf1DM4CAL+0tTEsmRq
1byYohYN2SdyJZsOeBhiH4aMpfYgGikvyxMIQsCTXR9yIPenC5Epvkcv7Wkn3IDGibn8OfZbSgl1
PrIoI7qm2r1b+SBcUzc0vjP18MsjG64JDwWareAwK+OWjoxj+fkqJyW6k4nVC7wxxwQbikx9FCX8
d5C/w6TsFOAUtQCRFYGnMB9qiGzxtaaiy4beB97sibMvnbndpxHJKytkJLQOmk9L6sfb7+JjvFCh
xZ+lx3x6EfzoDWiMQMUQiij52EsimA1P1R9FZE18ul3cgYy2gRaw80uSyS6i9FxlcCmCBhIBSHqD
xjmkBNmTFzs5l/WANpzjhBfpFUNlNIffj+kBJ+UJf3eL2Q6SzUq7KDFugRUNOgFXhASClOB4P0Pe
J7jCD/+L4AlCpxAuHjo+mRzX/tdSqXfq9M8EKCRZ4MWWwafqruZpqvcCbxsxKUi+Oa+DJvtSDrG6
NDmfBQmzh4iUp6ZdeVLcMYK+Jp52Ap8S6Ca8slHhSsEtc6NYhG5C6dBgNCmrg45UcY0ZQgLkqZ8M
T8RTJafF1hjHHA0HoqpXNRCgD6nDyhdlzl5I3aDJfqVhhvxDaOTHGSfVMeMPeB3p9mKgX1HY6cR6
MG21Hhpa63RxtoI6qq9wMCYAqoa5Lsi/j0BQBP5pm0q7ICtQSlGcf4PloJljDKQIOsHw9Tj/PheQ
IhvpQHCN9bxE0PPrvNU1cRhGMene3rT3z45iloL4u+hDK47Kl3uvJef8KUPcurt7u1EVxYwaClTa
Wv8kaf4lWjj2kV5q1n/71h9ZCF945P6u/g6plFN3C9Yctnurxx/AAJ3NipfqjEU/cQE765X5QgqA
kPEz2WHP7jumKAm9YCQljTbprCotinSAhhvzaR+nwtwHpxnNEjGVK9T7Y8rqZ0uWPxwBNhK8M9lb
AxQlfBU4urT+BcTDmJhbxXoShumMMSQWQn6BdZkiicsMfahI5mazjMW/ThMk32hToH53uHqo6Ewa
wAVZPg9SgiCTmmB0ODYC1GMnc+3aYo3qLZQQ7U/R+FQRhGYVLiyZnq6Y09qf5S+dXArVB7hMNu34
xT9DPUu8TIYNltrBN21y7LGi6Tpfz+LsydIq7r27AYSYd38Z39vZHexlgVNUW08KLszRNmu83c91
rGgk9Xw0wYisnx9CnfHMaG6Sxr/GQ4DcX3Seb9rlBC7Z7mqTsm/fMLL1SO59p+J6C0+yiYMuzB4c
Vyda43Mj/ldJNfzi9BLbYIrz0WBNbzRlx3FOgcXx4HyPpVL+RJHX02EZZK88JYtOqmiv6dGufwkY
vmirbl4kv2jHi4bYM8OQ9fhUQJjYAz5nGfGTkWy5QV5JHRRQs4YA7PJ9r1V2lF9rvy7XTQxzpIu+
Yju8guKGcQIn8WFY4Il05zTQxKXHXC7cMDMU2ejLlWzbHyU4dWAk8VggHn/c9h0i8M/IXVcG3B9+
xO0w6aiLT95szG8wLOXncRofUDkU6Bv9flUERTLX5aACUkstLVkQRZVhJCNSVtDFECAoO8IPW2Yg
4KEf3NgylgYm32un1lV/ERZpDAXwkr8AF4EBu5zCtf2RVq8yJgkEz5Nb9dEYACRk2hW6Ec2CGPQh
dLFqw/vfAd8vM2AJsucXR54ymMLOPfkfTqTfD7jwb5TIJrj9kogJOffibN88UV8JKdYhbVwFCeTM
GdrrWNyEJgDVP0lrqroJSmaex7lDB/v0CcUOyV1Xxj2z0WjwWENT9BCX78B7HIzdWlCzWy5ZhPq6
h95z5wEfzajuf2qOh14espieCejt3rOb8J9erj7936pnNzFlAyjOvtQnkFyd0t1o8gRj0H2eoGat
iFp4wXlzGiAuOUmbVXfu0mtLUemueW8fuUDRnoXzOWPKOlJ9XPO7siz8EZloMQeV++vl6HYsaX5n
qU4BePgXPJGE4yLmSyJI2oCiBTB4w0xawNnYJrysrAcu4KR02QJ7BUM8foZpfVoL2wsPHnMSgfMV
DQS8NoPs0JPL2JdrW8p/FyBSf9aEoU+G9eg8najItGYq2zCF8KmqCZ8x0qtL5CxK0pbUBPy85tLj
vQD5Emz7x3qc3zEBhyk8D198NC++q5a2O2VpudDuopE+dLCo8avBdKzD05pJ+12VJh3hPjbUs3g2
zB7nyrvGOBVlhog2ANZUaIoOfT2jk/prC2XM0zryPZsuOY3SdTGg1k3J1m0gZ0MqmVyEYmuuGsbI
x7A2crUwEzUUK1h5hXsWNo9v9XbyInFZ/6K8J3BXQ+syq3sZ/r1TXiIcc5N8unjSo8pdz5WMRs6r
hE7bBzUn0JZBF8/DBBtckKBy9dAqPe5fmIXBENU9R+ZIHZJN8wfczWJSvIVsQ2C1tuzhSGbgJcQ3
XwloUFYQRwSfFhFQpDrvTmOHDwta+VQ+y5spmCBGVMtVYv/byUyEUEX6JlSRxMA2t7nIAsjH/b0J
RN0AHp4nV6EsTag3+ew4dWNiMMv3QvlboQt5uVEF/8IMLia1MP3PTQGXyi/pcyogILzB1DZYEbjY
k52ql77wEw8z8RET2X4i3Gvv7P5tr0ffDydttjTFfRRilHwaR/KSppQFQOELBvL6ItbS1Wu4QgCc
d6/O+1CI+jN5y1NOlWkv+hc7lFIku+i9v9GHbH4+QdY4iS/X0NgRkjin72aQQzU+VVrtEGG21rHU
mWKpa5moqv8EMzvFRZztcXoe9RhiTyWTP+EnTAg04p057LW+BG8Ldy2A0TlUwL9lxOQ7DkNJpSWZ
tJcs9jZGs4AIY4TsrnTa1cLcPkYKu0mhWX7PmaM4wPsZV8vpA6sW/45KkcJnKT5lXxFyy/kr65jD
iSA8w34zqkeZ0C7WOKv8l5uAPOIFr35jWyCyDhlOY5WMNoX1/z8ZMM1d6FwnQzYJ81imBRX4zf+r
nWO+HbJNaHKCGjVKDl58YyVOFm+OIk4KWk/gihqQCYKzhNApp5FltKJpVNdWDHzw15pZoaiPkNbt
Cwufn2jyHX0rq+HW827okmL5qcyFpnFvAuoWO7IH4EgJonVPrlJHposjEWoE0iMH3XFt6aQ4i/Yb
93DteBwsLsjiPbn5iL7GSwhGt58eFUhL+881SgCh2fomO0VwW4CZ3hG4UyCpOQ7olaMkoEkjigJj
FqblTNJo7ARzXXr6lXz5To7DzAzwZ+0/8co/QYJingK0gGdQyZwyYdqtjN83iAhGax+7ZKFPpe8W
rFaqTyXnbgr7pg8lJ79oNpo1jZbbM33dkaqmm7YbSvZqh9OHGFTp9PRGwa/DjcnvpobQ7TI4dH1M
+c63uPUN19mL3SZCaCe/7j3L1Dr1s/VxOl8bNc1UUV2iPEnOz05dGg1/cKrNo1OrvN4T/SsHbI7U
7s4DqGnFBcdQRIRDZuOSIHjXZq5r+XrxVtbAL2VNR1VSToFX7eaIs9E8Vkmm7w3Hvdo9OCdLUSFl
MlTVLN8e2VgSnUdE1RC4WWaKKWTItD8uVhL0GqyBAZ9dVSLZ4zNyD8ttGnO3TteBevzj3ruHeJdt
w6cSMl3zncCZ1BWVD62nvsQYh4kGZU8L//5X8x3joZNZ/K0t+fSnbS2VhNiMr9jz0XQYvgmnuyp3
LD5OJkED9dprWHY9pHw3FYXyeuvRS2WAkPaQEshQUeYeZj6n93PZdg9/i/8eHlx5nCfNgEL1YpYL
2cBPlhehv9CDfWhI2ggpqVbn0Z5PFbCAy0lvsnohcKeHiTemB4Vx+0m9Gr6UmXoaSEQWgbl4KitD
8kXMU5FlBogAaXVH35oOneLGt6h2atT78NoMJMp6Y+V67ro/j4HdLvFGqdqDYpP7YJN/g6dXRTeV
eTRvZnQB0jI8tMskKCudc3edbOW8AOzjT3t3kKNnnvFVS6V/wWkVd4wyyxLgf82FIyujJJLHt8DJ
qD/gBSL/XcTadkz8MvckB4LhEkdx0pbTjFOw2yf0VAc1ga28FGu7EUeFyzLPMJ28fo9WneRFbTE9
BPaMmXrwVs0N8S/NDCTo86tx7UUBUknjGYpz+qTBLWG9HByK3dE7k+YmiOPfwYtkmlyS+xHF9bdd
nK6Gunn7LD0MKEnYGNMfst1iS/EFuFEhVRF9ubo2h36baRWoE+86jMiledy9rZwyh5nSfCvNZkdj
pcmnhPkboAX/22xxETBj6mSl1EYEUxIsCKCsvQfOqoBavsfwRdrmC8DTb62HXlJ8SHVkVdA1KS3b
NBZLXhIkjYSJH3/+eG0vd5dmLr4Nc4l/3Es6wtDewp5A1n1b/omzN4wM3Sx2Mq0mse50QMY55YGR
LayJ24zNsDLDTAKx4LZ/IDO0vtXl3evTV0/EZEF6WMbzHBPuROQxNJh167az01MF24TEriFYtBm6
Gq8p5mg2Bd8NgNQvHj83KmdwRtZ5sLAnPe3Z8XgOP6C/SHGgbAaj/9y03OdeX9sHefG+Z2Zjujva
RFbomf8CI03xhz4LtAHuEBY+NM3Rqs7MOz19Ib0o4sEAQWd2lE7gDBjeKhMZKtB1cmH4sUrvIXju
NHsvZ59o0tOmu7KAvjPMPG72Wa8QomN/5C+emxtyUW4ssqVTq3uFOdiyGsooBoOWzY1Gfh9UyXzw
QNtvq62zjp9c3Dsw009o2yEXDAmY/Gu+vciGD1MBx7xckwDagNl/LAeyrkTQHl4VOKs7hEDhQFIa
QXh/y6WmxvdHDkrJjE94GfUQlENXanFAlFGM+JOw0gCkLc1ZsjPIXQvdl2tWN2H6stoDFDEke57s
hgJ2faCzi80llJB8mTsqnjMXHfhm4klGK6AHD4emH1MFakJP4KjWik9WknWYqYKAzEsXFykl4PJY
RdkszYSQTBdTPS6FEPsoV7YxNi/igsH8PVWVdF1Uz1WYgngAxKoZtto/ceyJiCjoPjMQp+JPAEzb
Um3IoNz5gzh5XGtwhrHF0xM10XCGERUDth17dFBr3ggDtb9pBasiQhapSFAk/I27H3x4Et7LQYF8
oOZmKWKjPMjP1/CqWZ7f1syLkOFy962OjcxfuJCZ8SFjdYXiCv62baDrXv3pc7WO05VHu7SvFuuv
fTl/BoQ2ho6mYu33Gso3pwH7Q6wQTQ3tsIHvnHDK8Q9zWf8RTkO4YR5dEFtpH/seZvjbGRsdB41j
XibagJBQUATjoI9ydNyuJFxA6tWxy7Xe4s90glU6tbz9TOWT+R6kC9MWqnTMRPwNUJYUW8vj1FX9
I3NKS+rFaaGl8eEX/X9vsLNVBWbMGQPzo1CDM/rS6DKrNhA8+B+ratxGWwG6arh2krmwD4hPT8ur
I5gkiN3z92WQOXortEP6i4sKeSyTeqLQhJVQ8PQPUtZf4uFtxy7qVU75XdS9KpMXEH+ZAXQXwIh3
zrGF5sedisVORw2COlnoE//52kovuE0glAkJJeZuEEXNsM81ARl4GxtSljf/uM8GVzYWg3XKm8Qj
CLNgoleOBb734OVUiT3OUBFdxdAxP5WFvo+Vfnhc9Xfzwm9cshTjDwfQpWUNu4CA6kLcF9mt6PTX
TqsdBZz7hzy6cfjoEG5ekrhLCdoi7TPS3A8m/7m3Tc5fXd63stkuI8DssVGSgI7nOL1oSC8OK1y2
kFTTnZc1BN+fjjkxXYF+lcYgBfXwCtsQ3NZErhH9sbLdqYEwDDGQe0LLB1mqBmuyx66Uc2ORhMRl
VjvjzwAgxI0KqR9QB0JQA/v29HGZwN+pgQcKmhaiU2aOoXUPZzIjylarJ44Q6Zb/QIP9VXzPetjU
GLu8AGjISvh9+YxpcUxdih62PAvbwN6yjk/1ZM5F7B+t7AL6tfHbxs3Tywllakslxpvokcb62Yfs
dRL/NyEjQqcPqh81VRsFTPR4UnTjD4hUv5X5O8V1xwSvy1YhjWyJS2maGPcIsLO6Ds5vE7/T6hrq
uht1ZV28+cbrO1tYmtz00COUmubMjUbS8iMICVmvHARb5+N9/BiZ9TQ+bwJNUWjTRjMNjZcTyGQa
Oda+6qubDcpH71yF+uwFjQ2Qf0I7sGKLBJvC92uySPHMqA2Lb9v3t4c6Qnk/Hw9Kf5KiumIcwLhQ
pu26XuYv9iXm3l49X8k7j0HeckUZpvSywJka7Ups/DQSI1c2B09DYGXVED/AdDA9ufm6qPJJquBi
YhedI8uezDl0UKx3M/xbPa/I/Uec3oB8Yzzpef9SvsxuiV8E3chvcj/EwImLE18s+5VMEK24UXp5
8fvmV/cFXs11tZVXFLviZRjfC3hcyoEavQ3D1nj1ak/+fHn+YqNoB8l7R/2oAjiht7nTrubZtyW8
MsN4SOqutFg1FITp10hz9cDIOCxjnmikCjqP6QwtjjPxKRuWfBRDEMbCANu8T/iE5jJbu0ulhv9R
ULPSbnHtO/p1DcxriCAvy80N77fmEodwiktgYzQm1r0pxwb5FAFYnWjgQYcriVmgN1mFscdIqgEY
ML5euVyIzpkIPa0Cu77zKYqW5ZXsaAhq744n/gd2tekohn8opXfNfW7qw6xBSlvKCRzAgj08OqVq
PGtUT+P+KOR6Hsni4O+1mxTxsgsd+e4Ens+0MDXagCqCl3AoScyZEHjMjtSGkjBA/0qQTaWG74DE
QYf0NJyHvdPWNqlSOEDoPmJcMHh40jsMPVBGHas4yMbJMBS4SHk1iD11Tz6Pqe/GM3rl5JzSZFSd
Xmnodq6WYW+rknGOkJruxL1p/pej8EEpptYY74UwR0giype4mUe7m9Spl4ViLtbGegB7xt6rpRHJ
+XtdXlXES0g7OP1v2nLtBx0rZpZrQ+SSBk625k/FV3YPq1NidqhUykfIPkPwe0KOWvxQinQiPZOB
GGo1BrgGG02hFA0ZLNLL87sRjGytDizYfLVjRhP9RJn1OyL7YDlzqbGRq5Y/nDjNXFyhkk0B83Uu
Su8P5jGP1iaq2AhuDeM+wamB21Lq1hk/alU8emVRoQ1GITYaZXosFNw6VUaIwazLdTbXOlezA9P7
wG7MwtbHOWx4eZC02aBEFEYKk64jxV3fLkrghzuqrwBy86p46Ac9tM9VjCogX+FBqWeHIMm2bhKp
aHgySa+Jg+5A7HNvaUYIW53xRH2r6ulkVMoaF6xvDG8nFZOlOYn3orqz2MkcfZBdzHUlnRe2k4+D
0feVLjz6aL74Lc5VErqwgd4mILtsMpiV0EDGaMTY/motCd5PT3+Go2xTYi4efk/2hARJOIg6FSCV
uBsQ+nuWQDp1RoMjegA2E8zvXlRy7szdMzwE6psP5JZ4SoMrYnnA58bKRmIFlSZO1WFKwJC6aZEt
CiKj2t0zffVPhRAze+KEyzhCpC4BknOZKk4K8R2j6+4fRgtO55ATKey41KtMaaExjnHWDLNsPuP0
XWboelni9NM+arc2o79pb6MFOjuf1KGt3d6FX7yS6mq6sTQddLMyUG2TaaqE1Vq3A6fk+TUHDfXL
wUyKJgKaZ0+StNWQUz+/ipWl3sbYfeYuL/zkCV84w/lQe8pI7SLRF3Yl8UTatybOgdW15H+rs0d+
OMEoeXjxYHxHuggTB7pPfCArflVHjbyUvQnWRoV+nc2XEVVDpR+sWluCFGPthdAvppwiM789p/B6
idFkjf3BLSj6lYe+U3uTy44C1Lw8jqsBk1zDREYHooFquIpp8HmAFvEAnHZ6GGbZuW4YEKpIlw5x
bIweGcQVbwCOGuur6gQ0VP6DkPQFRa6Oi6oNTZg35hQRLgS7P6LF3+lUznQYvJ2p1GfjPjDArzFT
YAeMGWrakPilDLiR520ZmF+3vFIFS+VjNFnHmyzwfVBZV2OWzz17xkeMcg47NTw9xY4E0vdiRdHY
vEM/ezbnhFncN1y3UQv4WL+9A08JBh/tjEC+JIO8RfKEMEQbHfLPqhsUZkAm8FsO+bAWOfSzBEpR
9aK0zUR2/9HBqMFZaVzHXMhWOLE2QUGF3aZ+vTspT4P1HHqnecoAGXQAsXPRNWATonlXw8PYcAZu
Vjsn9JrJuodYcrVjKB9K27WwlDvu8G+R/sl6f9UKVpTEL0ejQ+Yia0M/GGBQhr5RZO1BYkCeB7k5
TD1tTGhAwZ3k78usHE3usdkDUPhnnPu770U/JGS/JForD5E2zXYyXzEZbGQnaiFURhHfnY9KVAyL
4H6MXx8SRvX9XHW+dVRX6qOvvF11MRBp/eMLB0wPotC2tkTj849UloQDAmCIm0CxF0C1KXEbZuvV
NoECrYaVWdVt36uknpbOqc1TF3prRZhY/Jo+aPkZWiOnNUuBcy+JP8rLTaRb44ztmHSp6GpGfBis
MmHFcVDIzN+B0qOyulOxmVR5sv9iPPgXSU2K5GsrFAAWi3eOyzPJq4O7UjwmaQsrlU8aYxFnoy4l
aTVVlgLVLOD7Tqvip+6Yq6LyRDq9+/hOMjmMZZ5j2VNJQG02xCrSqTInZLhoId2O0aA5taRW66fn
I7MyT9lI8lW+u2q1YyfmknMVFfa5BJExvYXU04bvhyqHxHY9JU+JR223LFJ2w/B3SZNsAYUShx5m
/0oC0XGXaIRz7mit2hx2O3w0Roz1/iCJKhG1veH0bDBTJ08+w5FyRbUhAktBLbkcx8pFKI8gF/Eh
NIqdJToB89p5cTOF8G2Gu9I0zmaeF690iESz1WU3f6xEuBN36FS+ijJ2vZOJfgyW5RAuQfmLG2w1
+AWs1vObd39O96t1dtwE/7vKFLOacApzZw9tDctWEBN9JfX99Az2LAmowN0I1R4cPYu4sG0xvI64
fF9hKFOWat29eCfhYDLuF8EqyPtpN8whEzEj3I3u4sxKA3ICCyvpKoCW5bYKGx5aowc2ebLkTXGl
fcWxhFvhuQ0wuf2TVYlnbhJBTiBEvJG7pfFpgI7qqYyWCgAtqd+dsmdmpYJq2Cna3Bf9v6lZfgGv
2+pHbUwfI0mb6ozIRXAgdqnvLfU7OvMpVxl9Wgdju8W3H3qyitobtCvZc4phOjMmjbSb8chUZCMK
VFqNBVk7E4YbPKLjv9KMomUt/RcWyyaoUPq7uk2FrO5eRtZXwGOTZ167WiMA2YkZQoINZkFEQCm7
VMrADnE2ZJo3oLEjikh0+gCwA3Y1YGkVCXKpDJi2thH78oV/+wWFCzDf5tWLNQAAhMb2ZIgjg1Z4
gsZ47wqQEUOzoCWcW75rH7AFHugiODee5/HmfVVbpQ1RJrgIk8Al2plW7bMBIG0Ekc4mwDRDwJ2l
jmRBbedckjYpmyP1wqHgGsGb6vyBYTRgAFxLJwdpTtgYxNrAkKbwS7JVO51p6kVV/aZqo13KjEBb
IlSvhtbluyMsmS1MIvu6P3rjwOA0mbkGg4vvDK7F0EJ3uNNQkR2ujYATyjyfKXQDlAndUrAWR9Jh
GxBsTbQ7g9GC/GdAQKGdVX8a0nskpdSCa9G4QAYCbehM3aLi/LwNp3X+NVPUl+5hDBD8llV4RwN/
rzie2z4QKv/9elp4bYRtYu39AQuTN3lvpjRUba/2+o2h0j112fFJhALbQBL10Z3luhOA+SZ67eGz
ZzVfy4Exvhd+RMavPAWt/2S/dCUr6c8C5ONj7ZOTcv8FXSI07huqIouObhb9MvZQdiWx9S46yEtr
47sUxP1VQy05Brfba97pTP6ProuLdCFsNyu+B8vABxyIlhELpZl+5r9DqKmPalF7zPRZOxckE+Gj
tiUg28WoNzrzVK3Iy0ql4FPHXmSFf/dlFfnJ5KkmBNYQIl4xzG9dMgBM7g+wCx+49JpeRFZNCjDI
TeTJcxnhDtQ7/8fJM8xYhMRTjeU/aXxziNK3AZCJ9ePvQ1QoFbzS07n72Y7P6qN8pD0hx+kX6OOi
pqTkpzROSDhcrEXANdc650DMS+11EryZJyefhudz7hi8dBzuA0vxAq7KV8L834/8EGy0DFjrU7du
JZANlGIpKGSTQPyATSdCQCo0eC/wGXNJpyvVZlfM74kR4/yVQS7M1QsbsGVX8PAf9PSRd8V4L87O
Dp8BLE03Xx/c2W2e7oU9KcBhCJrxml/gDZovKhkpY+cT6b9xw/29+g1Wm17sctOROBJiVcIG+Vdv
/9BKxo0C+HWz6Q4ynaXUj+JViqba08fHof018+aQ/Ykl6Jdc+//X/D8ThNQGnW5KyLLfCWNFnxSb
HGelZgjZGT4/aw/KqWnw5l1DygU4E5HvVkLhgZ8fgGyssdwyjjFcqD8cdM4GggcGKjurSTEeAIBh
Ltr2qtIlo4nG1xGXOrf66cDdTXp9FgCOSuqxUS7VbJY6P1LbkoGCo9K9Snp/8Sfo/JKHdAzcTxXP
DEIrDXQAyXinlRKDgw/jWfriMYFWcJgz5bpZ2BQd9YjksgCA+iUbEieCAw8m4FSszFMc0z/DznMq
2aoUJCe8CTirYk58LDWYC8dFTKhZrhMVL4jhRdD17Cm4VE2TI/Qm4IYF1gzqTjDsgYB7JE3cL/yi
CDTC5e7JTlCy2SYMDdggYK4AlPNXzsQLyG+5AAVczptZ0copPaZHC+4l99vabDrGR2PQo2zRzSIj
uL/2UyHwNnNiXZmN/W5B256RW5mW2Euw643xsIzCEE5aq0XXROPiQF/gqvQXrDix990Kk6Uo4QtV
K1MqTMrJzN03S8rIVECCVkgeg0UanoFpiIF2ZL39aw2gYjkigRcd99qlAqSS5xiMXESSuJNndBnt
DxTqCG7RfdRP/SjHm1Yfdw3z3lKBfJWrt4B/eg4MRCOCzgYPPL2/PuufEG+yTKFRR9KqebWWTB0+
KCwPfzbtJrNyAhv2EnDsu646zSm/mzV6ofCM+t+toqBaSFNQC43OIn7j4v3Ncj8S3NBJtcQ0LcfK
it8p41SDjLt0s9cQcJHBRFrtiYfxySl2nXXSF6A8SFMqSv2FlJ9brNwdBLAzQbHR0ktt4tt0D86r
ObI2IamNkW/WG0LDESATo70Tc7dVftLwsIouoBTeQTQ6C1T+ah3siv2cqBshSgCn/qpMM2D4AJz/
mKP+PBj1B0t2vUrvp8S+2MIaFxPcmYsgHifAF0zs6olWXyHyMhMDEUBH5a+5JzVTuKvEs5lKyF4O
+oUm9OxuRk4ow+tKhiN6rBgVDwAdBMr7ZK4MIJ2AHmvefULleHNUpdVH+ktFxZfWi8yRTM3w9ZaQ
AvJrguBEOIw8zgh/T26hBb39HCCQAhZhDsExrYL4MfgU/Yl3uX9Rs2vxMGd2B2D1zfp83gDXzZ7v
nuAr1uOtjlpsiAYf9hoqPhKzBdDn6c2K8D9cmYRoQrP+zIG4mZ1NbqQx9CAN3CBEXp7C6GK/icxF
hPde31kfLal9ZZeBJN8xKKO0V3lfbkFjqIBqVBPhljPbLpn/XWp9+PpFkz3gTq1XIujcie6fuun4
iuRAc36aT2zVepyoRdfFtT5SYcCsnJZjLtm+wGiqBoyGBBgbw5GaTpKQV1GLs8bXgIxxPHdSxRqN
WqSyCintLcbly4EmQk6gxDauK5GCnJv5hvl3ri83puSsuLrScrGBnCq6r2Dlf6kPPoyylaEKqsNE
sWDBqOn5BCVWosjW1EJBHsixaUYat8qmyk9jMR0PhzWf7Der84XvIJTu15HeG0j5XomX7aOR0LWd
Rx9ZrpEG+WSGLad+Srs6PUNs3Ngl4wCSS6cOOs/Ppk2e6Pj3voBjfkfVFZ4D+OupdsBXkH13qka1
AISg2b5cIuVP7oc6UFxI6snOMEQITlSrEemB+7pL5svyAs+kEbtNLlpcEDEnr1jnvTrjK+3HFwzG
/e4h8gI+r/I9SoYHxt3cmtBXcjZPT/wF8qlrOUyL1XhTA2/3rxCmamhLwD8M4drPfXc7dp1+yQt0
PifsnwCWwFN3ylXFlP+rxZEk9yBtfloWYIPRTPnRV6BtduDPUIKdJ+0MosbUctmoaZ5brxvXNhrN
/cBzYh1VYRlCkNe5ck6l4KILJyHKYgO8ob2bwuizKGW7lNj5ypgazxcKIw67GHLU0dEsBgh7EgGP
Dc4+u5RGMS3RALenD92bFrXtLhVaKWo84+u7Zr7ryDDzdC56wg4yMT/Y1bOL7duOKf4aO1DukiTh
OYWJGBk00/odSEBH1EMeOQpXTG8aZVGsDe3JA4ok1yldsAZ42VmznDISqjDjW6cG7D7y/ST0fOHd
cKjEJHyOacU8kudLV1U+9p/xk+ymMcjgOh+skCKImhGv0F9OMreF9UdIrAPsfmAIjAI4oad/AHQt
T3d8ELrr+pLuxwrF6syhD6b+c3ngZnrI2vua5dyOBs/HvSgs7qao8GbjjDi+QWeqOaVcyauya+vZ
tUlNKsDWdh+MMnujdlUfeUt904L3u9dG/rmONo4GN3zGQ2SFiUqs8WLxOzP81/1mKjdGwj02NBuG
mVypxld5PIhQKXGEKHRiJswQ5tIo4lfoRkvF0jkvQLGZilcep8zkFoSVtCttpGX7F3U/3UTfXWty
+/CgyoweM0bjoYu7MBQB3HD+TulxS1PolKMdpwNJNjTwiObJHocV5ub/lIeTdAp7osYMV25F00no
lsMH62kMeqvhleesPMhZU8Su8HG/blfZEOrKxjyRwmE5gicw1QV7cTOGncCJmclycpzNkG8lE8My
yJHJfIAnQWN9ZZtY22zvmNMxteMUgeXfqDVZuxTH5yUfL1NIqHPEtLpQQkGw6iGZiixA4HShmX0B
34sBf/Gv+ggO0thAJxAAD4mIZKHmZEUIUhGw1PVA9Qk3HUUFbTn+zp44J+tp0rBjqACPo5LeX2er
sLhbt/WJPMMnaE7rhs/niYuOopequE7R5I6RwYuKdkCYo34cxhYVUcpODaWmu3RLAUD0PBSWUbud
8bkStgS1PGfARKGOS9JTT5xbjyrxyTmtax2N0N2iph3nwhyRcEL5ydi4amh7OkOv3XCBn7XCbENt
MkF2KYIk6IijltxPbGGjG449y+b/hKeDXy1fMduyB9w5oDK/GmroXo87bFpmBbtDoCTlvD12jvAp
fxw81gxnCykFXDQ0KLd8iJFoj00xLc0V/frV0xHsP39mEPjitv6iv8NABj5GDDmChFcNXbvLlPGO
87aYDQB8vsijFpaBhvIZVAELnRFJs8r3Wa1gw0wQmHEceNPtEviXpmCFlNO0CyJcJiC9wCUjAPiM
3WXy/vKks9hEIpMb0v1WYoGBl0cCO4U2LP1JmJp1/Zu2WNfvmfzkzCxLNJjUswO429MtT/iHVowq
uXBhsr9JupKdUgmgKB9HvfaBhEHu7ttm2E2fEbkKJdvHb8Xpb0+AfKd2/VBtl+QCZ2yR7r/Uyzke
RENNn+clmwIMfR1DMtBUjzwgcxMyHJJq1n1IwXc4Qq2zVwTDZ5d2PdUX2cEr/V9KUDfyUC1i2E/R
teBIF1UDhWBMiJvNwDyXO8Gs/H8MY1elJTxLI89OAfq15s3SwIVgNZxdFucXdIFE/EPbtOEcqAh/
BEkWK02cen3tCKIm6flxFxMZO+amjkwsjEXgrv4VmFr+L1n9rhDz5E1edj6wLMm3edDxFwoyLD+K
lib/UcL5rE/IXs2gZ41146c8RShIS+tq0TqBcizTUSSNuOgCo9xDj1DGreV1FSv8O5t5lIG9XKlo
wWELaDDzEMBFH0ggb7zrXZsYUSLwhzk23lDlp3wzQr45LaJDXKfI/Rc7XeW8jwJ2nnH6jx/rgFUr
11x9l72RwiUgXvb+smuFurDaol1LO/tezoyqauIWwR1YBpDFBJdWL6oLKJISKsZDDNrhyy9rliGa
UFU/+I4L1jP+2q+yPTxgSgG7dun1jGK3R9hYFcHFOUp1/zMPcULvTNENB8pgMmZOzL3IUh4zV9Bi
/qPt02L+mqkYUGEPBui3+8eof/5OZFfnMctR4k0BKestWzgtrzkfR8hi9AA82A/5t3W5iVNh4ry8
rUvb1I0skzbblUu5v+UNJqOrP4u89ExnjGAxTfp+31oyLzf4PBpzgL6awKWROrf83R6cTxVhqN3T
FJP4TfCzyVoXb4DG/R6x2S/Kcj0SrvLxCUioda5I+fU1PlwaUgEOB/KwttPlon4Qcryd4nzOsQ6p
gWPFrRQGRV43E/CFAUG8y9Wuck2ifSBklqlI8r+ipVcLiaS/3UtmdoL/3VSkV/q66SEq05Kvb0ja
A7bVIs6+Bmydv9VT+jyKh+BZUVO79jctsN/WEB317Wo33/NaRUc+9UO1d2grlBygtzMdi4tY+Sv4
ultmGzRue4zqVHnknkOHfKOpn034d0alhQWxlo3NpX4/SldHP6Hver8zKJp0vBQe4VwX0zVmzhsl
jZmkTDYSC1HOzODjt2SNuPgXXEml90XzF2nz0R+eG9LQ9j90Ass6gLCft8xMkDZNWzMNyP/PU8yz
UiJ+ZaBGuNXEOnRtPXCczrM8DxN3D2Cw41k/jtjuxhI3hoWdyv8tjArkQ+cxnqLbC0l1fDzj87O0
7vNhMilAEXg8A84twXtLjLmWgyV2AFjVOZ81zY58B8sWV/BfK006HOsSFkst0+EI7S03yabfnmVB
FkrMwF/HBR9Uaz6UbDZX1TJBVpPfIpWfyPQue3ZZZNiMLikfvkx4vrH89TjeJcsvQ3GSnRKydVeg
SgGBaisFo0DxV8diL/b1JV3t5Ka2yx+kV3cJjUnexHrVrEOMjMxGksASp3cLMoYi9dYsgadI2zRc
xnpqK7peES/XdwzOBKZp1VMv8Qkl0lyyEslAVJpb/9AMwRiZwUI9RYgGkJHqJLqc6J5/p87TR+RH
LSd3ypLJTjMKMRygXRou0Tjz//XrpLD9HJgboTiq4Zm9941M5u8wHc0tZ3zGV4Mkz2DQVTaURYUh
Q5V9ofKV72e6D9F/9n3A/KPX95EElmkt3x1nCaGKdh8kGgXUzWHzApbU6vP6Pl9NVcNvLz/YsMtV
wZdpLqTVVI5Fw7epdkyjk6wJGrNrSS4CnsF1AAE/BrRevNOc9iJ52HuUd2PGdg/05C1aHvGwXuct
B/vUhlDOKnqMKsYOB7iRLwq3nOEW/CqZEIN8baMUQlAqSWjJmuFfxEJwiJyHaszka0CUR6aaZ/9c
KSgjwbrvU1/ih0MnmYAyhStIul8O9oJxwxkp+nCjIRmCcLFb/hIm4rDHV+YTcg+fY28nwiPkTYdy
LGfMGqXeDYazHnFQy3YqmiqH4rF4mSgBwYq+JQghCqqJQISxsb1VXujHILagKIcHXNPHy8JnPPDs
NVKvTOIJnhBFz0qrVRhrwkhkvz562pdLmrjsfBpnOAY4OsR5EcC/ZNYUj+XMkGBVRSuWaVsIPTcv
fiJt40e8oa4rdGM68ZvsIKfs7y4/NwU3O5S0ba76sEl/0TuP8qhz2wu9tutvyKzcxyEfSHWB1zTn
+VrkAr/9l6F4qMESoI8K97EB/WdhDP8biKlQYJB28Zb1ZY1N+wGuPvArz6Rg5iLGbQHe+webOmaA
Vug/Y7FBJoPR8CbH5pP0uIDfA5QEXZr8Vg+gNIcaqDYIijDOdPSdj99Ox7NkfQgwAb4MsnRxk3V5
Hv1OhIbqVoOUhinx3mhvWH7aMDEpCFQ+138aVya27SXOBehOlrwIDW9zx9Lx6J1R318zb0cBE6G+
C2X85nC+hPr75BdvOnWxgQC6TLF4NQgVJvGHGqDt8yTCkghAvVba635w7YB6LKQdeOs3DkA0xw3S
DljsFg3bLMIZ71ckAYpdaa1V28pikbd7m3nXHLXlUbHNH8XdVrf7dwvefQo6eJguTIKdA8u6rQ1e
39eF4vKhtAq7kAB8H+HN16n5AAFN05038/aplRFvaEXqNABvLKJr+zrDC4O1ulTTvZb40XmM4Oo4
smJHaaXa0nBSYCeAxg4qofjBGwARad4lUInZcyTl6PFV3Zz4BEImOSSVsJnkFImL+8Z0Cpx5Zy33
EE0j/oBp6B0PCHi+ebcmlMdN1D4hjOvycb5vXHUPIAlOUuM4YbL8pkDt1E+LG1N7ZcS3vLZuNXwy
QSxYt0yhROWtN4dzxeyxznjNtJjFNeqUBG3tAWN5U2bkAs7OzmFSZ2IAGK88sKkFO5lvsGzdxjOk
8+DeUDaCYCV+2s8Uw9GZn6vcjDo4yB/ukYvreshe9tgbXhLZaSYkzquxdWD/rXGQz/Im6WNdyWUo
Ry7Z2R2UmsPVBdzkbucyz+TGYI0HG3G9IMbPne+ZVVDmuaCBmp54X1hg/xdPdyee36H5XeKBuArQ
Y2sRJ+ohG1RzpToNpkGqNVkMobuvdrT8Wwtlrwy9v1RzcmDoiZjyoqwn2uIruwkD+YrE5xjAhW63
UVdbwxtKlal4cMTsHsL+BW2rzgdzW6KgAUZDl+3ldZHlna/FuLOB1d0am5pn0nLP7ZjeoROWxmRV
c9frbENXspfRBUc3jD0DFeV5wW4mJIuMZD5tuFsgR/fxG7qBFDj7lFGRTbeP55/FtyOPd7v/TPfG
1xo/nE+JqO42E8DrW0jjxiwxslV4pcKJcOM1vaCI7lLPiB1Ft1tF0fviTm+jzwh3WdzNSjNv7bzm
WeOl5g3n0OcGXwgIjdHHpX5ikUkRpdmxl0K47yMzFWDoOTUn1L3TBvIkiG/LbYCo8v1RlERtk6RT
u4+1SuwHzbBpMEXQPU4F5DpL4TcC1nyNJq/ua0sLPWsUtxnKLiFelpIh3jbkMYTtpl9TNqA8qzLz
mAfm3kuulIHEhdttkJTiFKedZ5C+IvWXK9RFRUR4Yd3J4tWjZloTxd9JA31m0UlztahOnlJ1qZCr
4Bz78Ig7Z3qOiTcTc9+rsbGaL/xZGj3J4C1YQTUT/s9/GLk0B0/IVYaonLpE1ADk/WMClDzHysjk
/vK/T5xt+6Ye9JAPmQDnd4UGJgDhPIehvFtGTsf9KUizbjao3AWnPtUshTETTeUgw56Sf1KKov/4
QlSC7jVeYksv/A1parb6uRwKcy6AhJZIBf4uxpg8/T2qTrlbzLf4gUN7ApeFZCmNRc4vJZndeWuU
fnITfCCx3l/B7sT5/0OkgXQUe82lBSmhytARLLsZKRAqTstM1W5UqVqB4omEQRJ8ga9TlpqBEkyh
bGcdTihejX3DNd5PxboDPFtF/BYCwq7851GCIkbwojCh0oaK4krBaTGxAFcxxM2ikY1x9llSgtNo
+fhf0DXpS1BgjQkcNlHzVb21Nz3F1mMIs6gcpYymngP/tV+diMGQeWR+Flx2ndKPcxR9PZSMcHai
PvvwSrlt85URq/kQG6ILTUA6XHh4UI/WH3COcg6g2LHUrR/RoM4Ut7aSRjdddL9qlNOeuiMbe57A
zNIHXdygzw13JMdWx1PJZWUOoF8oFGvoea6zWh0Sp0jQovGpjjfHpBowkd/YaWinwu1uYtYLb9PN
adAonN6Q9vUXpa/eS6HVpgUGEIurEUJvytHB5H+mcuybxBaDvAiORyOsFM4Nghtx60YvCpC11KCn
qXpWKwVD2YZqczU/7YIZLziQ7AG+c5XzY/ZMA4/7MfEmeKobzTRJrPaEeveyixDhjuKjsCLD4+z2
kpMYF6eJFy5U64xDcjMcyDbhxzrQfFyvgumu8pv0Rtmf5U/El385bvzFDsk1pYPQodG1imYjfDlY
amFcCZFvaux0up20M9v29Omv9qpUXuUeQr3gwIhff9rV4I5pFIImPZHiWSlcy8CNsc0q616O1ARk
ahLMhO4I2NK23HFQHGvGwUlvRyLj46K6TjCAY9oQd54Rb+s9c4pjKi3xbyyp2fZRzesq8pwSyGwA
kQ3phWHchgcBT7le9iKidcuL5xiRG81NFG3lGV8FalhO6ZnqW4FAeyKmHabpRMOp4joQ6nHmlRYD
3jbW/uuYJRWNmX+L4B/Zh+bCuwF0lTJdRx6JFpb1Mu0Eow7ao1Rjic/ThfotygmOzaej6H8y4Gvq
FIuQAwNekjqAt6MkKPi4gzltTuVG2hlIHF8NKvhCBnMDregQ+nDWXhpMlW1Rfm1Gd21BvV+JPIir
fyeLB+qWxPlnB3gQ6j3GSJVzhYaboHXWGccPZAcz2mxLBTsjIn9LyNi5oEQ5yabdNnY3Rge+KNCI
ytPvv++dDkTWVes4zozAxuC9MvLaS79JW9CjWFA2mcYtThDHLJQjzrtCM/tU3ZExgkwJkI7/Eh+m
LQkudiAAeVGAnHM26WiLViv7J1Y66iHiZgeZSfc6M4GMx48h027Z2iDpoksdaPqPlj2riORGqZEi
Pof1VBEj2Xyvufg2WMar80b6a8mCpihgqlK1lzxcCZ2epyNdaf7oNzgrUcW0trXgY0uNQkfO7X54
GaDVsaQVOs3wYJfTmYY4U/rjCrUsbuQdHYWSKhd4r97MA0vr8fCwWg2h0cAw+HUBZDLkV/hfURtR
nC9URJxKPO19LCe8XwC6mzCVqMjyqaML9oYSV1A9UmYRUsoN0QIGp9821xRZcbuxODkDhKqRB48g
D83YEgfTm79SqPF/WzP7i3mS+X7dAZcCJGx6km9npLD9HAzLfllezZy/qZhgqvFvgA6JV6c6oX+S
SuuZqgxV2nQRqz6fBcO1eVJxZl4WOcLZMWbhxuFDbWfAItPmkDGkEpafFPhUQCZ15+4EzgIXgx0g
zGrVpxzogKyjG0PyEO4S4cBwLhE5FVLpcDAy4Jb7UnhRGdbJWx4VUx2juBf60ZWE69FwnlnbMuwK
Vyxh2Uwta4WpKJzwHNVKI721Aqo5U4ZQx4kPiXagtaB4ABMXfhGYOwVeoUnVkU7SPH5HRUY6Y/SR
gfGLvPHDc9nusKsqPEQhONKk9wec3psI+1rDe8/Gcr6NflMY/RkV1C9xhqjQQGoduzfUslG4S9KR
721yM1brGOc1XjpdH5IWkuCTM/ACgWXkQkMBoMrdIleEor3z6YrUA5P66GsFaa1uSgbb7eAtJGPG
Zciy1b4yXMjStxiNi0lXSUvncOOJ6oB5zWIcKjZejmZFfEMKMZizTTAmPqjEcT8lCz2BE2737fe6
TWKSYWbT6dIRifGP/NJsz38Ui/02uFpw0fCe/7oVIriUMGOKw2amSKkLF4UtbDPAK0/PUAgL5VG0
gTZ45A0a4LXJI8fZu9rlfMjUwZrYjm7yw05TJNE3sb3Gh2bayPG0S8nGwvAyrghlVVcxxf9eKLb3
8J6cbxVAfHuWo79EqMGoMHmOGskRO2TI5+xw7aFSn4PbV3MJhb1M3YQjBSIxKiZS56V6BBvT4x88
DpX8aIRRvTf/Im+QSxNrV6KPZg5WNF+zuOp2hgaOCdZMd26MT+eQ8TEWhVD4BNdwKV3iy4Ku7U6Z
y2Db8Vo7dTPC2xVXX+HYmL1K8cmnW10F+mzAiWVr4+7haSRJ7FG4f9lZIf+wTPAwoPXqvzgIRBKp
hbIE0mRGDGGDMt0x3qHMT8sjIKmW7PPsgwYYadcNHQGCKPkW2gLHaGTo4n6gidR9W29/OhwnQ6bI
PgQEDehbep2SMrvxAmvbc3rz4HnHA7ShowVE+/fKj6zkgFxzA+KXJax6z+LzGdJi5zGZwl1IScbi
jsbRItluZUqgQS10dpH4Cb1DlKeViKTnAVOSRDbuSPdanD/SuUkLvR0j4B1lSs/2ANqoBgWPEoVX
nv3iSh/GOPGUb2T6kBY9/S6Vt5w3E04pYxxTDQXetMFloFEoCgq0sXK1W9ULEdj1/b+M2DTm4Dm0
0xSvu7jzzFmkjPjhbNDt22xLaIeUKvaKgVl0P4APcPe5cixA8uyVqKg/OZXx1AL2cyHwuLI8l8uU
oyzwBLyUNEihchEfGFoGPy7l1XxqWtZuPTmAumHmuaZVl044rbR0WfaAmBaw8B2HQNJbQEHmNasd
q3vqYXyRYkgfBhVUx15GeZ6KKAG9qczhsQ6tYzQE8/BA++MCHyrH6YLuXU/DB5Rx3keuMkn/QOh5
eC5tavkeQi9ZW2eHWh6IMVJ4yHV0tq0VFOU4aqgeLUCnjFZAK5RfB1WaPyVK4cqScp2S+0B3nEle
QdD+uzFEgjcxoGDjxHO6SK4huNXARWzKQN2kcM9Svdwx4sUxXLNyvg07zbt3lar+/mXyZuLACiZ1
8IMMvxTfRkSi2SSXX9N6+910YTmIUNgjGSpx48R8cKBX2lddLOL8bi1PDXKiz8M17SihRXhWum/y
5CKpzIgdaAKgkRnEy6jMj81kXNEPjCvCo32iJcWteqiUHdH0nX3/FhY45MRnPVl+TwNcMENmuDKU
RBx7BivnCIFiZOsCo8dwxad0Icpte9u/ssqAfmUndBjEctw7qXwQDtYPZ4EKibFCzrCMtMf/i8oH
E96qfhphdken3sa5Ak61Ut5fwtP6yEWI5rSbEsQIMOaZrZxrTrcPJsIg8c9YBHO9NHaW6i5A3rI2
kdTzauRw9CsCQnlsnkz7l1tUkiVOi3IbhLMAWGOI6E7ZPmXHeQw9yHG0ISK94bPaIE4HDScVaYF+
WGXNMx6pTNJRK/fUgP+oQuY6RmQ4QoOuCR1eDzgW4DJQk1inwineO4tjcXfa622EG5QkUnu3lptB
dRXPBgFDWfbsx8lV2GQD34S0VbJzvrmPYoTXwQ8x1ja6hHUgWvLxcb1Dj6t51acRQagoAVz6ykVZ
N/88BhY9DnZfzuKM1ahJL5mPuOsQrwi1kb5Wrytodzvgq4R+vVGGw369+MB0Nosq9fjK4G0qh3JF
cNZvkKV/UljHZFH1leCVuVhVscU/bQIMJ/WRUQGAEo7sW6K0hpA6KTb9T7P+xUaDcusTenmUzIPn
aEdL2KxosbN3+XF6YBlsvtnbzY1k8JpLWV705ESCIAkw6maqyMlf1PMq9yI6I2zkDPJnKJmv65wZ
L3u7lwscmPEbq9JisGD5+49W2P/DjXPK3QXy8/CGZ7aLGCLAplKd1cS0P9O8D9KvMEKZBHQvUCBF
TSvSGjAeuUP+XO+t3eb5ekr92eBR2dkWc9ZhuY0sqIwjzZHQK4sVIK5YVlyd9AQGXvUOOczQRMjH
ExdFb82I7A68WIfPLUiAdk4S2qjhFulgA0RKB+3DqMKoVzIgeQNdylYj/Y3Un3QhlKNcd5fjicWK
WpdYZ9VV9LWacau7Onmzzc+JTu/wao/LWSYCWhaNRlP0d+ye7i1peerYx4cX27phl4jubT1XdOXH
UyQxMGefYTSnacYEjuPniZlG6ZhrYTc2Mx88s+xgsJGmpmPuV6CCzk7mmPndVy9AY55gDCO9hgSq
M+ZaRexl+8d9qWrchsPYWXyhi/A060AaURp/uePrqpjN51zwEGvE1gDJWea7xT/vg4Wzq/C8IcRx
4IddtfnBROwpKpUN5wMesmoB9OCeUpA41AvvaHZh8QE9b/M7yOn8bOeGtAS4v6FJ18xnaoyo0udz
cmmcIjGzgJFXpb8teCNcoQDP8WXs/JC7xHbzb9uA5lkMRXgnCaVJmT1tKbFVVv3Mrwjm+ruTPkCs
QOaG35JVQzsh3EEPUbo4TJo2RaSYx1fIalbjzbXVxh9qRIrS4W0Fa2gYhkGacpnJr5j8BgADJgA6
+Z92aoD2l4vt19FTCoWid+9S0+5rsSYIGne9MkmJ8CSEShm161Vf9+YxbXRSMharXGI6eOlFQBe0
BOsM6Mre9Egp88z0qCudrip3I0atJ2Y+1/1iPA4PvH6knfwbxFQpH3e4siC9F9GNkvNJ36VJdcGK
ym5w3OiJaDO5oK8YqVrdkvwZ9fRE+BDgwhjyPJCx4+VK5p95bJfAVGpherN+9UmcDyQyLVK7mZHE
txYFKzTU76TqEXT0f4rEppI7/N++JTlKPf/kqaiNgZOXSqDCxfIgId8No8IZwc6YDD2wSQcGYp64
5UHNQtQBKHaWhs4X1iVqm6cmpJ2/SvUwMbrfcbKFBZ9yXGE6GquOO7ZiaoHOoMF11dhRauNWqJVk
6BAbd9QsKok8//O1Kllc+RB/WVsnu0ei4Ei5bYlVdOEPauH9Cb3aGphyWt2A/cAFJ6WJ+lgSMVaX
o7MIX/enUq19sU9MR/OEIEw7i9hSCwTXdbq/mk26cFF1gwv7XmBFKHz0kp7utaq6kJWSy5+r4o2J
st8ITQFIQscQikeF9vG2907GUvOUkI8Tkg2mfAawhKjrR3rDUYwRqyDtQpKqgoVNTXCJJjX35pnS
WfuyrR3rq39mtudvZal/r27LTA2tZN75VEmp7b4PbPFt5v+i7FQujsbCt2tMaeJ3jz/O5PjCzQXq
UrRLzqGWt95kL8E+X8OCCZeLU5JGX5SG9fj07BvB3A5MTyYJZT2GKzXmdmAbRH3jwv4jejOWMGAh
Gf63MNfs8LylHLxn0YlUOYJh7taVTT4ARX5FcZWTFFNysvbVqSpHRV9Ex2f7Zq8jVbb82VHfszb3
Zy1rZodyr81CXaagoH/ncPjnFahEIAYqgjw2IyrPnOECNDayDU6kOEkDDJPZm0jPjMWwUfwmiV1a
GzJubpShhVVp+bJvX/YOMoHJ3B0K3cQZV8WdHMDu5CDzDFAHc/w9waDYrzU0T3TnHSKv7owYvd59
0J82KaGAIsCwpkRWTCiZX9TU5LIMPefvvX7RT1hR2KnxUpI4wgYkOtRn6wCOh/fiHl1MjcB4YvBj
qhcenklrij4w+gPACAdlItkWoTjm2cnxDh8u9yWpubXlA3fVFw2bIDl3bzTQ0ntyEgY3xswnMpJy
pgApDitTHPdgR9iBkcVmq7BIlRYzj+/QSjRpc/u84FlVJOMaJ9CfFc1PvMQLQcoDkOd+0vx/tO2F
Ju1utSpDDfHgpS4ANOs/mBURsvafio/FRzrVNbUFDB2JkIZtNZuOQEjGcOZulZc3FFq5U3uHKbzQ
24cxcOgOyKJ9ZrULegxa5gRnITHju2wMBXfBZsitDMcAI6sFYJ23xj/SjcFdX4YD9qx1HuMb71Bc
4+VLqnvKa2NUEllWaKEwzTuTGlzjmNGnrr2oOjBrtMgpUgKFmn+W2KPsa2PMAtdbxw7bk9pXIi1k
xeeNBj1DMlcEj3b8PSLYFjLYiarv9G9Q14KwWy5bwJFDgUxtReGuywcA3dze62IqjVJm6ozUdJli
q3PynA9jXG5Sz2Yj252MaK4ZcsL8lG15pvZspNWpSnLncWWb0qr2VFAJa7jgx7v+8H9D0wjHv4II
uSKApUODpC9YGwYZU9E3M4nWvN3yNud7MMh/Wa2h+Yc1ySEabQqeuemt2jnAJaAPWwspFNFEEL1u
gZbWScCFve1C6j7RSmup5KsIC4VGynaGE3mVMPpIZ9LDC/6X7ESCsUsXU+ACYeIXydgzdSdTfcSU
xXRK1loDJjvqQs3QOD8+7ESXf1JtVO1mcZwE7vGwSw5L50TN5Rqq9Sk4hWf67Kf5DDL4qcm6OfbX
IAAmewGOI0VXY8a3CAfIqgT0flx/mpkgSy15Iu+JLimWBcE2ZwZpdapYTS3iDTTJrM6nuY8P3dKF
4fc6ZsKeTx/g+CO7LAWPsI623PXct/QezT1ouA3NwYBwrCHSuGwKIw+Tcs8ZYEzQhw4ITcoNKic0
5dlM4anQu9neyQbWwJCjICMmJvaP/Z++yaNg/vZal1aS/Mjp22S1C0Zcgop/7vtWrG73hH/ytXS3
dwl8sCp8SAbIP4BCtArqLXYQ3oZsGO8rVc0cduPB2mqMv+EkFWeQZMrZQXF7tB2oHHtRlkl2Kgde
M64WFpGmIFVhalBrjrjyvsw5zEwUxBxMvLJ3bVFJ0/VbDcZ12dtjoXwEcKtKKZNGdTsx6VdYnHOx
xt4I9xWx1NtIsYG74MgEmoN71Mc2eynOkj5qoKaJpXp3R5MhPAZDMgCx0GVOJl8QFIeni0ySjJU6
rmXa4Km8Zw/n5OrSRczomiNkQ+7ugkTgqsQsGm8bQ2uaqIwDJaupqFxQtnMPBFRti9LbBVOehFbl
9822EkkZYpBxPu/mM/MrGN+LwANWX9tqgcOMjaKBSmgBOQ4A5uwKizNv1VWoXTt2o4SsvCKszbdf
GNmEDRx73/bX3jfWQmmxQN9+GUHFMNtKV8HmosL3939BZ7pxygrQkkBJ9pMKe0ImIgvxIMIDf3KE
0CU4feM8vNY0yzR8Bbrav9/YtURIfQDWs/eOUReDQxk1O19/nWKOqsEY1dEzle1lIN1EJP9EFVg/
8eTeQqMj+BMNUve+wBuLlvK9YH1qXtnGvK228mBkPxuMQq7I4y3NXl72KewMqdae7FluGOLC7nUy
04gnOL7I+MOj1JfWEq7UR29pnbyx593obGGQ7RsYEGmWRDoSZrx+Q+11vcvgiyuwnsNTLpKCj6Ku
PozYXMzTy1iMS1nTclBGccTqtbtZUHgmAOdZhpim5HGaH6U0AE0olvJ0WnAzljJBhzn2Q2ctUoeR
8G9rw2Spp9RcxRaZFs/HwaDg22Kombl0cNUp+qA6jcDXz7eEGGeMXwyYWoVw/Z7kZNv9gkOXTw8b
I1M3IF41yPdCzVCAFSVJqvspNIVNLMsqIPHLitlZLhrTP8+3AmxaiYAGm6m577hAYj0rHHeK979i
oc2a5nmR08m7YE9A9ZnfG6ovo/03A9hqxG2Jrj7ckl/O0jgcu8p3uxEcxJzaZBrNptLQwaxnUK0w
mvtoszUz1LG75limRi8r1PwbazZipT+Ucy3258qUFhBndRpSvhJzHoTK6GotCHlDbXXssL1TMpSP
bbNLQsGVFF7GGWFe3t03bUGo0F8SFzsUxzTcF3CxKPvIiAMaHhOdxiPf7s18Zwvc0Ya/MXIZuqZt
eB1GK2YtF30UKph5d4E1UcdxIXf/Ln4F/EBjy8r4y4X/Sn1ZrV/Sk2xlvH/9WH+OLNnKHCdy15OE
4Vt0kkiFhCy20yK2YmlP+kNYbYDdyIOWn/FLfEEhBRgr+EgsvEgpo1dIvP8t+29vRx8cm81oaceN
HZ4NAjikx2WhgIIXoQqeU9udEVJVV4pDEuhTwjmgd50AhQaUvkqXDS4qhA5L6ZvvbcsEJBEC/OOd
OOYnoSweM9XQRRA1z4bJjrJpY0XmKrXJAriMEaDCYUFLfCNtr36oI3pBkLKU4MCDwo5VzT462doX
Orp+hjDBBZBMz7FvVLP+mU8urm+WAaG7Fr0kHSOpw7njIfm8VNsVNMvIaQ1oEcq9ucfCy5klY8Pr
VidnTNMx0XAEGE5dGDYDU4h3y5GiGlAwyP63js2fJZiVGCQLC+9VKVFYOwRNo/9F1EG/0EpUCJ1/
JldScEj1X/rbA8vVSe8wDVxEZyIipE6mCIC5jSQBlorMk8u19eEkwNSwk4b08agi++uvUfj+Zms3
/H6t2b378FQ9dGlt00ZQrsp5K8t3Qp1qRFhV62fsbqcZjQQzPacfkWsrs3Dl3vKNnQCQM1uhOi9M
N42nWBQEtYvzaN8phxqDrXRlFfS639Z0TIZXgsfcObQ7RKPQJbBIe/3QxUdtu9dgeDW9DJWz3xCQ
UDwlXbEG/oWEoC7S+HQbmFpmf/GGCTfq+3VYQnQXXa+NHy/zVxNGMpjkK/ibZSLyECt0wKXCctvh
XCDUJ/5fTjBiof0Hf8bXpfKYejYjA2sJBzbwAOtWtM+ZLVgjWX41MlO5LJpZ2gPuOJ1+n7mcQArT
F18kSO8gG+QLshXDZ/1Ocxh+7DXMtPYLFQbLE5GGYARNOiFtzpjA480WU1pS+hezJY5iSUp8dx4T
v9wQixYXBUMYRNmErhwdH+EsxhZoGT2dtEgttRGrdLWWL8Su5PoS7Y0TYPysw4bEuwfsGKarrLFC
EubQGxeyy7zxuAkeguj91vTuBc5VcTFHu9GL61e1itZ5YHdWR0SCkYsjtvEE5bzv2ic0pLf8qfN1
wAW/uJSrlrheenFcvfw2YHE9P2rB793LGFpN29YJ2BMLQaKb1lDVdhP5vXZDGrRBdGIE9UBfi6am
nxa4BxpQGp0D9fLHEFrZvfE5xvRdReCFfJpJ9CspkKhNRvrvOAClGQbHOTGRtqpqNlDzXm2yNY4v
AqH1LkL8TRiUEBFIgKLJmL/FB6yC1g6hEZhXKvbFfkEureDufY4I9hfAYJpw2gnhgEITmA4n7/t9
Y5JoJvF7Qnl62NpIMwjheZruvGhJZbrcYrP3TVZ8OCyuldZPj0LxyVZBl2DTo8ll4bdAXSuOXg9Y
7D8yknS41fLdp5Vdft0+eGH244MaE9zkE6BjmkZwrhzfGwh4PIpTEItbUBK3P2dNeSDQMxQODMUO
bqZkTVKS2A2ZBaU1+1Zejdk4yJKVpxt1xJQVVm3LF9S+UCzFJL3Exeu8CFa9QJFvbamYQDx026gI
x3MdvsQxEiGwZn/1QjhbcInAIgdPehWa9L4EfR7dyqUbmooAKNSiyHKHIlUvEm8eNab4A1qPPNxk
5kEpfWK3RXmaSUaR1wHjGmoE5IPNE22BOb+xfGiOVkJlnJbzd+DW+FEiyprzWy3boaJ9DWSOdkQv
G18RIhPWGM3h5unpU8NCyCoEJNkj1dojr3GbdtIOdsGes3mCJwsfOLxoA66twYy3EiU/GD+XR/Lv
6DvNsf2iLNezO/LOzdVIFdoJS7kdjMqDZl++C+gVyQ6tM3UOI6hgs5VSHSHfjW7kS054U1gd0Z4a
5Pp8dwDw10mle5A3wrxzM8D7Vi+SCsiQ1CSVEM4zK5qsINyvPUzgK6XmjX+M1nMvUL9chc931uos
6KFDvdWW6JSWJqVS20jHmX4f0EUQs/lBnSWppDLefGpa9jixvtRh5Zg5lftNFY9qSC7s9TBh27mN
fUQj/DdpAiFk+1+BaT9k5BHAWhxWm6X9lBo5iXEA6LjMHW0ONSyeL4GGDaNh39Z+ept9PmxHxiq4
gBM6PiPSZtKctRCe8oE40I5ZcRwb5gqJIogPZdc6+CzOQ3uN5v6EJ0TSB7ukW1whQaZXCLSq2Sw1
fGFoQWhTWNpa4kqSP2yHnsc9ev6I+o02DbpwSM4nutVx4Bd7Qu9vAoJPNvURFxOs/CTuZVA4uaFE
AKH6n424R201gLT7xd8SxYNHoRoUhEG4iLxds769OJLoyqQXeUKwoh3Oc0Eex0/tDUt62/04UjsV
eXuEAv+/SqYbvgbI5eGS23nMBwmlJ80MItXPOjc+uZ/xymeGKoNv3EYbmf8PRR5DbaoNkfn2xIPi
uSe6KAXEod+HTy3DHGSTqM0ox3dF+BapYEKu1prd8ezsnubXKi8iJBvxVgmyGk9LLtmEnR1zo21J
30FmMebE1nv1d/R/x/sI5N35TXhuMtet14eY7g6ONpxpsCc8PqOL9H/eE6w+pO7twLvNg9m0eCpw
bU6LW+jflxxaD3HcD9kozjIXA1pPkUkdNb7mTt+z//+o1XiUFt7pWbqgpFBQj+2HTss9UL9SdKxU
abBE+j+FgXQnDE2r2ConIPWCaLJw8bcEyxRsuM1zTFaespB+82WBR9NcbrIA0MSGqQOWFIsxAbbg
ML/LcrHshChL9sKoTqGzywryctPi5FhSDvSm9SygL0WXLiy60f/PPgPb6dOZVOIFdRBSRjTk7pbj
uBscT7WyoBxKa8bTt8t6SHSzPeM3ZD73EcWguSMamRIpwd3Uo2bS/7gmyea9mhQkwtY+C4aecqJa
aCDQTmlhYS6xvDep6tdX7xxc1eiQpspYGIIDKGYR+UZZ+mSe6wKeItz/8t8yc7ahM7nznx9m2du0
9gk7D0Cl9Y4FyxmkdDNg6wl/NRCGdYBgZmLuMkF76Bti9OP4pC9nSRlCV/NqQqyfAOBQkcEXnTSN
gu9D55kjJbjx/hRftg3EZLFZnB+YOnSKFdmj5orztbOBz4fDny0w+CtRbulUvh7V8i6cQyU6sVgL
QQoHjyDHEaMlaJNkZ1YQV5m+DxPfn/r7n/L4PBVltrZCTEFPDl12SX+/nQ6d63lXS7iJHk15ZI7+
fS/mZp/SdnFZ7dugLI0GNuMWHLIXbbxR0W7udfjX8TEKUN6vJSYp1k8W5zdhKMRrAZe5Af5/d60Z
7ibF8fJNJlHp3d0Oq3utZ8tZNc8n66AZj4u5D4RGt/dapdAjs5q/6xV11fKhSLW7sLMYCQBniIE0
tK1d1IxzgRvmSbYVI/9XsV6lXCzW99I1ISfO7ch7qT0t5muk0PuXygbZ30lnReF7p529H0FSQE6l
hrOTuSoy3IcTik+JcLArWn2Yit+XcRmOPPoBP9UMUd+nZSQF9Utk6OmmYUqlsR3SVzLlW5U5+8Vc
J5uWG+8X08S7W8VAYxBblVDuipaM1Z1cSPrwjjmc/h9DsxuFK7kt/jVkGJDUAoM0GS17lhYXmwoW
a1UU7d/fdqy3dHZhTrASgRa0SBDHk6PvE/NZJOzAqE+Ez5RkIgGtjMwXIf0KFdbm87NGzKaq18ag
m3BUCguThKEqdmk+XQ79IoAeO13+xIePL6jjfO4Hv5WwNMApElJqZl58XRmTIRvocb6pIO04McHE
doX/2nOSf427iKt/XeWmtOk5f5gbs0XrkhvfmCGsuDRlBYfAEDMH0seAmC4CreUfPPKhYohrhZWx
Ofhb/3qYgpzR3Ib52/WXy44BP/shF8tv2B1IBHXNcbVzHcAgHED8GualaHs/V3+tZNTGzTbPpUJ3
yEApRh1SgH5SQ8svaiJhHIk+ZCvxhmlmTlz5OT1NCOpWfu+XDAzBhHl8HCtmjQ7MoibOKP0rEQV6
icC8WVx/1JUVeRM4bOtbTY466+F15eExhq1DU6J8F2cHqxxJ1/UScmTw4z5sqpPbulXyfOUdw+Cb
nhYHa3opiuV/qg0WIoRsnfXGnfjlcjRvG9DFd6bGUWTxIu8c8ART2F5LJOjAlpqkAwtw85K5vX4l
Z8hR4xSdO4MNeKPzD2QNhqqfFWXGWQi45brR2TzqIOV52Qy3/9Y3g78iUMfHHocEVGVrCgtn99PC
2EwERrKxQR82dlI9B3HN7CGrm9K2oNKj0P8BhlDtkNmLJK5WKd44htHAyGIJ7yB791lbvWTYj+PQ
eePUNBxUum0DiH3mPmzksrwBw8JKkzTx22TIT+Sgq7vXPtmayyANTC2IcbLzs04zUn46zd7S+RqY
sDPg2Yd2gS+qqOKHvqi7PYs9Q1jObemDuUJWDsGEgS+9EataKbn/J7j1NtuOtRnOkriZk9K/T5oi
hPJKLX+NJqxWnWrt8ZjB3are+ofeK5qErmO3B1/x4y37Qa+Cwg9/8LUmb9oEOuGW3xWpedHk3Fty
yCZF7l+bQV0ch3b0c5IgFPeeprYMVgc2kDCueF9nKT27JgwpuYFGBKLRDkH83hzqNz5UtcaLYvhM
K26f5y5zDPMQZvlp4bh/WHmM1Wn/WKNa1VAIZopXECn/L2LI5lXcqdFLg42UZG5r1WHzjFGlCXv0
u8dTxKkT9gnXLCaSK+9KChnqeY7+WH4INmMZIz6nh5oGdAVn9nvUn6zDOeWBDIyUMAIMMe1gXqMh
j0T3dkZGu0G+IYKJtYWhTWOZQ2TLTtGKy/tlKIKOwP9YhQkE/qTxjyQ1o8sTM5zzyxLCCuz6q6wX
MNxkQ6JYEZnJ1m6P2wTgAM/J4m6PJsMtVHhZvhOEe6WsXoAixN5iCjoBq8lZeSgexSj/y+OeTv/J
S7qzV+459ghUfsocJxwGkUefpYBzfNW+cTWq81TSdBnKRMEWpCXYEsuYd9E1FZz3TBMLp02lEgMz
VZQuJNEMmWSWhP4NPiTnQYRqBPvSPNof+wGVCWc40SzVyl9uOdhpeBLD80bFs571Y15iCXzXfjYr
W0xN8VyVERgUAQ2g1vubpeLE61B+BZlRPaDCM5FgJix8KHDgbP/5J0UoQEiuQL3I342iehLaS6CQ
WzlP2CwOYaruXzLC55iJcrOlvo6sGrC62hbHNNYCU6aJ2siqpg5FcLURDfrsdzNOionJLMTeMUXw
lipm5VFocrhn0PXA4y6w/X3AjwxGtcFifBVRfneWUZ9Z94wlgg97BoirxMvhoYtvyLHcu0HIi4dU
l4TQ8XkvkhcBM2SMSgjAp/8RlwosEZw/Z+z3qCbOiFoY7jfFhTky8WdT19lsmmeHyrk4/x3OExAE
jRoXSRyBJ+FYyh7Sy2uI/aYmYi5QbOQmzTE30t+zkWLf6pNTa/vXkOxEPMhfM4HLu8a9o/ILZSTz
52GNgOq3Twt3iMscraXsLwf4jX9UfBpljmfQXTfXgVepbaauPSz5nKCvyOgw/R43gV/SrjRrK8LH
4xk7n3LntsUq2Y7dq3ad4I66AAxP9hRInBSI5xaXFccrYvBn7YM4/SRVfZXPQjGTG1Cdn1XWyDV7
10hI/dTAGJgWFUhhihzQFp/sCDF6trWw2KdmBi32bXZByZyecIQGi8MatYgR3uz6x2PM+pzuYpVg
k/tKT8dYiGrCjWet4j1/aMaOpXV63DquTykswv5FjtKZmu1O/i7i7gnz98Wtqf/+NcQY4+oIe/Xh
2g8jIbc5XGlV/qf9vEHu186+QS0FhqqAvWYnVIO2LnCqvtVHEUcR/+LzEnCQ5YTFnNB9DywyIWYX
V5qkp4+Q9a48Ilt03oZjCNeaI75xG11nH+/S2nh7PgDlgNFC3GiAgQ61YrUDgFsH19HCGo4yw2iU
UoqX2753xsSrNpDujVzNdlfh6KFbXc3Zl2+FQ2dbymAA2EVEg22x6Xsq9vUpgWexvVXrPzsQpXBf
7AZ664mjUh0k2osD1JH3KWtN0FXKI7qCdN21hZCMRK7Um2+ES9kn/bQOGvTduCMAuvZV0gLMGsE4
EglQuBM+3NAUFbdmtzrJHJQVfrlR4vLrcpfwPoUbUMix1GVvns7NtC1vleWJoo4SG1ByK1Js8ZcJ
FN2JrsMwKD/s0p33Cp/LtmchHMRwepI+/HJJthQUukNTePUUqwejYN7QdQRrt30q3hR7z50qQp9a
ZMqpdBSKm24GYIeRmGoQcU1NABmQUrOFRAK3XsDlzTO3VtGenBZBlQ9/IsEjNrFYjg4JAbP7T2tz
0tnn2kUeQ+pziuhHZMfJxFU/QbhnxKxCbQkdviZ9DJOR4+RzavpsCKv4Trgr3jbAS/dKh4njcLcV
WRkrNp2iCdo1zjOtFZnCQMYESCR8SbmCBPwwFkYhJr/eM6TMngGtJHwlzxJaijgV9WUyKE+EFi0J
cxzX7OkOXdv6ZpmogjHxJI7TzOx4zNivBRNsvPyftkmOKnl6OolycSaIiER0ip0NCkN7SyP0uD0e
PRj+1eT5wLuLw50DNZ/KEC5tinQGnVIN4q2Z51MSYxjWQdmPBVcO7wS5hLTnXkP7gsbP+mJIFEA+
U5ex5iaGWh0mSgaUY/NT/Q9N2+m86UfMwPJLEpvlsLCsAC7ma7N9WtHCByzPsT3IhOYjqPi0pWtU
H+0/GZkpmaC+8++/4MJoDNRKGwmQQkJECZQ33jVWpCQKs6EpbELN3ttSPHo8xV269WsSOteUJzKs
2P6lgWwzIeGTiQ6/PL/Q9F3jKjPVG3LgCOaXBG6w/6xyaPeqrgNZ4GHZypU77rKcLJvNINYWOaAH
gqpp8MoyiXPr72405mxGrl2PuJa5KQYcmpBsEloF51vw7ofWa6jjutFVIvAj2sqpUGqo+mgSG/YQ
QdNhSNzz2447W3RbrzVyQEtKsPXtpXLr9SKNKMntv8XX2yhpivdcwI0E9kxRjfGK3iKJiMfgSgQH
kxQDW9vn21j5gE2l7U4OFCFX9BDswLMUfhCADhxW4yZ9GD+2I8q6H/+JG8dgkwSB0ag2WXWoGXeu
V+E4t9JRtkU9uqcPL7EHNrHlWaLfuVsBZhfdwQX7ByDjzYSv2IumOdxCsaUiv6kBaKpiqmLoqhxc
MeRMwkNu3A14b9LPWIOSNU0EydgwXXiGomeYxYNsGNjnZR/b0vf5xfdTZJRFjnxzg2O+rEYUiv1M
osA073OQPaFtdJV4HDHDNtNYxVhGpPUw/qcBu2KBe2e07hVMG6hd+RP8kRT6wNasBvNiIBxa+F0h
YmpnWmKIYvpoFF83PncCBlOY2PGdQ17jssKLPEm/2O0o7B9U3ITiZlPuzzGTAVW84sx/Zpg+Um4U
vhUA9c4+53VuMz/kyHKjf/LECUeoaoeePhxgI2p7dpJlhtFB7N/OB6rui+FUyzPlTOzElDIaC5b2
nImzU3zSVRvk5tZdmDBLUhCN0+EwcNXLAtKmYcc++aW7+zNQLreowdEVHNK+ib5ot+ZtnwEaM/IK
Ji+PKQxnr8u1TDzsUy/hm/KgL3V6ai8mGSXK9OI/5/6iKDR7C3Ot6F1e4+HzzO+yAcHezDJHmSOA
pqEdfOvu5I53z5lAH0/PO+m2wHkcTXG3DtqiU9bbzqoW7YeJcdaDPyWgQgdVmirvJ67OGagb7jJA
LI27jqIsiaA0MfhbUy/sBHg91J6lIfdgaxR5c8sgWn/J4HFHZ6YJBGiy6O9Y+7zb+KgayJPsxYx3
9vpu35eJvLuavHbONPxshBG9cmv9NSFuvEOyfOyUsl7s35IG3DWUYgF0JHObakogmLfOGtk5OPJi
3/OA8rPbOs9pomYHJYsxLVYxy/v2PyWMa3nXok/bv8tSeuwHxvC1WDgCMYGLlSJ9XpI4lcigvO52
rNrGktSzpkUfjG8PcdoWqHt0jHvqVUl5P65uHhLmJ8+NUTqfwBalPYZLoQUxTAMb16cVsgRNrtyW
To2srCPcmhdcCKLQ4bw8AY3VxoKkiwJyIESAlKxpwyBvVjV5Qn8WJNeIPMJpa9O1c9q4eFIDFYTh
0JyH0U66Er+2qn7ofkNIGgQ+u3oxLa7Z7OFDIn60wGAarQvly/5yOuvMEclZTWx1IfDWvGOIrwsT
PdZZ/bG82yg5rcexwo9Yo+59Jh7BgGS5ysKkAEWMtWh5xROwfBo9IXvxoc+3T7xK/TwiHQ6QrYef
n9odqH1If3X15ytqQgQHpH8OqwI/c8IoUa+ZMkBgFyg7RgR9VAu7ttveDdh2p3ID6DrO8Ez6oUdT
U04Fct0VtpC14X9XG5lcV6eKKzHzN/hSd7klVN+AnyoBGYdJHTnGD11Gx8OYpJIJ0eBtNDZ5hICk
gIBEj11tqZGVAF/hKVQaTkfPozUbpgxSnqMat1OkOF2sQz+HmM6Pa+p/XfMChuKl2hHRPr6H5MTx
aJVuQJpwWbrN4l8JwG7jWe/IYceoKZ3h2OHI3H121POJBuVsX5dUM/H74jODzoHTYUpkikgnP77D
yzo6IADFkdK7cymmShinoKl7aFR7aa2rY+i9N3JRFsznKGCDilk6lJqZwNl+K++Hd2zAAPKSvclX
P1x5kvObS4TzCnz58ZKHDxgidRpvYpKFHZWgKmXOShUV70uUSJshcfi938EzRa/rPgAu/SWpGCOg
0A8NRFZbZ3CRluygfD3XobfJiid3kiicCfJzU1frNIx1n12yXmiXQYIGDVw7EjOKqm5K1RemrU++
ZJ+kDttb+n/dhSSv0ECnghm+rkviHAlvJ3lsafZws5VgRQpH0vtrUbAReYmCx8b9FUEdmqcodOBA
IhuqFImMTGb4ORTjnER2udmJSwDYZYEI3Po5j+LnPbunMKos0uwSEzlRxtgslrAMZylXhJEc5cX5
Ni2N9srOmFRoazFcbJg2PZHNmgV9T+gLIYIRwRoqO5/LSeB2l22DdDXfowxYAgmT8wCnC3RENuu8
RuaczvyXNbLbyxXA+rP8hR9EDsTC3+hYv/j4wwbv2Dm51aIwIElNuFzIMeqjQCNj1i+Eny7OvKV/
5/YP7ayY0CahVXa8qsAi2WstdNuKgzanHhputym/20YzFxJXH5dvlTowSBRZijPU1CfeR9ed2OJr
xeOuanQDKceHlUkxmpktUKuJtjH38g/SRVBpPAuRy/o479HRuxNZhNza8JBBhLwZUFYY0wwNvE4s
02XP2GCVwL5ZYIyQ3cGXa0cXQmArsQqBG8NruzYtw4Yf9qwmwigtsHKtkALF85k6zDzNIHcDbkly
2JIqqsFbgkvJUcXKRPN9QypbK6CNfCGG3o/T6xf4jxopDERSl6oq5+vPmIMiEteeUI45UBzCT1A9
wjco+Wr/EjtVkJO0zHlr/jkPSidtIIhS3D4VtM6jGCzrsRt3JpQk57h2AJbNTz95DvbOeE6RGG9I
DU7iYFpDNexgIolU6tH87haZxMGKstYDPlDD8CAOPGi8spiZSiJtxoKecmrY25bTRg3WM+Y5B0LX
nINYB4ERMJlBNNreTtXOfW1efQdt/d8Fr0rmHx7Ewxg4eVFU4nHz6581PaRjaFoURYBqqGwkoNP4
XNRVWaPMpuUwHYl1il/GuS0LnL+Z4i3zOQE2c4+/gbqopiZgggVbMQHW2crSMTVFQqQvAwIemYxA
TncuSGFnfI0VPY/GNrbz6Y92R9IeTk6EXe860dbrCSRtl+YIruY0xQppAHTYRzbdyXJZMlAE/rbz
F32KLEI/RN2VUr97sIcNjuD0WSbp9E7edevDzoMQ9sZuKM4Vx8I1HO03C5d6jUykCLh7ZvOnnDOi
OlsAEohQzFOjzxdhP+x0XwSmS9V0vE3WKwFdlgtdt7iNbt1v9XMtCnfCellXmbDkWDSurEJpoxei
moE5Wgf1qEaohI85d7pONod8iEoS+hX43giNb+redr8g3hI7915sppYRqpEM5G4LHARd+QShvYCE
HDnynuoA17j5Qhm2NuMKN+TDnHZtjBfz6/Cjf2040sB2sH4IAm7mGruBeWlCraQRhV57SNbz7Bez
8NNtc0iFiQbmeqRg22Vcd/NgB0Q21BtJsKCaA6axkPaH6sVAkq6KMXKk0o+Eu/xHTg43mCtsUt/w
ZKyheMdLv2j7N8oymDbko4i3xWlVOCbAACc9GKI+JqbksNnJPlGrnmpWOqsy+q4InK/JE8oz/Ern
5oOxl9+x/wOq/UbNXaxzWc0kD78AVanIgznOAHc+9fOGivZgKSQNHDVATNcLgxjeK7x8mDVoxhU3
qpQ8vm7iN/RW33LICBx12dqZ6j26qf+Lpr8BykkSVsHe58+udWZ/ui6dDLXdaizQyaFLkPIJxhQV
LZOOiQ4bYMw9lHfJeoPvyC7rVfebVKWgnZdlExn/edtmQeNpBiontgqaRiBTRMiQQKboxdPR60Du
m6RbopZXrH/NknqZXrJQBcjgZ4+LvZWqNNK5is4e0YHp/m2jpyqPHnu+cph+EdcNW0DmDAOn/FT/
XI2qo0zAogQIfwmLf2XCfOxn5/QGo+rJuHb+uBqklSUQDi3klAlyu+wl1VKBBJVxF4NJ5hawBPWa
Vnm2aW8KVNSSLlg3Eh2QrK8ZAlvOTiRyC9ijxDzrgXATh2zNB8sGINNj752L+dwX9Hhky9Q5au/h
IGQqzk2de1wnp72hR02e0TjoxqpeJkdnfd23tZRvwa1n5aZReVfepaPWXiDC2lbLSjZno1+iffGo
E84ppyfCqxMNR79j0ii+N6nMe3DsD1kcso/RcXtL02ig1EFchwQv+mxNEH+DcE5VCCnh7KlAntKj
QEXqyQ0utoHC4rq0GxvbQmo/ts6yF2GTthX2Xyc4jCFk3rDVtvGSzgrO7bVdBjxnUUdkZ3q8taWL
/5M7JEomztqCdMXBwPv6OWOuXdYvTit0pYxzLRLe2GAAVgKmlEhu9+O6j4aQ1376yG6wOPuZ3k4a
bzQBLmReifRe130WkEaxrPCA24uVSLHdNH6tMEpbbvwXOtKLqkIH8HL1y+zgOFS6UQxknoWDPb44
rguSH3nmD5SJxPOPiQTrHoFX2fhnT4sOzPkaldFHgJzYpmmzc7SHYQqw0QFHuuSPHkc4PsuXjltI
HveVehiYylKI5eFSppMvkTWE3SW/XSMg5xRN2l0f932VL5O/ChcN7JyhWLwXnjZHZTxIDTbnfmzX
PNgsthpDJyeCTuhAXHnt02jg+KxN/MbQC0lvlwaYolRU7Kc6ut4UM3YemVPuikD5mcbnJ2fM02F5
tDUH+W4PE26Jf2VoNvn3wSMjqQNgwUtyFJJx2ZSTBjVxuTZvBzwJoF0rxhqk125AkF63NguJDt2M
SlPu+VowUXyaYKGMi71Cx+fa/0oG1qZQuIlKP0QCftAEpfuTbO9CBLZokQQTPQ4SmFsDCvd6Lcaz
4lNvJhh3jy8cVSqkngzCxXDUB9tuI02VqTEu64XRAN3dazF5fN9nMqUyhyJb8QcPfftdQh8ffVf+
LZ8syGX8W2GkCSR/HEFJ7tytI1NCb5IsPZeUYX7lnLAv7JB6kj4AkbDmE8EhGg/M1pYpXTstQZVX
QqyIuHJL9f56oks1HbkB6CJSADQJsVquHuvZIXS0Rxrkc+RVi8RayPP+nimUUsWtcz3FAIawI6s6
XCNqYHHVYNN92I8MTQt3ZhqkebJ4Y+hoKVN2pvS9Ku77+jCk0Sj7EYofD5OyO+4Fd/5vqYlOea3W
RP2GJrUSAf2FMJs8+Q1MtrHgaMkKfwyjfDMz8rDYs9K4h7HZ7VrRA06SmAqpVUfpchfPVxVp9m1d
e6gKrM/qE+71oWdO+4RiE8of8s1OyjRz7ZLYazZcH2xG0Vsvd/w8791CILXLe1MVHp6k72XuP9w7
jumAJDNyDIWzmVHA+IU8y486wSDCZudAFJF2cOXod465iK75ixTUrWP9qkdjrlQ8Fpsa/gWTdYRF
hLH/TpFX2E1J68eVwrGFYRa2H0SgFhgqqw+v3MigeP1t7vyER8RVg5T7/yCNernayb0LnUQjnXRK
8+eSBPCJnrr+6kA8rL6HYA20rCE3L5Q/P7+ht+6G0goWfuv+gbsq22l6yr09MZaBPdJ210F/Xvg8
3Qk2B8/SnZ2lwXuvlARF7ZSvTciLyJrFuUpSVNSTWW8rFH7Hk3VvtyrVTI8TAWiKmQ6/VTjhJDWW
4UHF7RznvdXYfyUMiaXvUNR6+geQRh9/NlRB9MqRZHdUsP0tp4qVThlfHqNkcNygtsupNPNBbvVB
d9zvX0ZZPNvPGTzkVYZv515ZyxqcAQOdATutY1mY1ypfbIV7NsNnfFZxbSFWLJ63PWHKri7P8PQs
S0gMzKXdECDzNv/PRbt7fIW9AjrnV4UC2CwYw+ioaIbL0WkIkIk+FPThwb8peAF9ETgVubQKVgZC
s5V4fm1SCjvyz1yNCuecul8tkVRdGgs5QDgRmbIIk+N3WSiyeA9B3g9hxCEvjd9/FGYPNR70kNv6
UiD1fPpngyNyQ6oFnf79qjgz79RZptJlfk3R82D8pSDtgBkLSyRXGAgUNDIBWIwnaVuuN1bixvBe
J6ix3n+CA57FneNk8HOieHwITJn2Hy4n7786YgC/o5icIq8BpXEKK4mhzzz1XVnsDVsGDDbm+H77
LBuYMoJQDkgmt22Gz6h+AmT4GebFBOkm4+F9KkZZxj0rjX5EGYXi6HrmAN64t1hPDISgQi0myLGG
8LIMmkJWRnm/oa+YKogKRrmdVUKiFbs7WWWskDNwxLmZVNQKqathjw1hlE6Hpqga7zpXqVxko+Kc
5WSSjVcAoPJed6mdbAnwtsc64cy2VLbNk5aG87/ngonbaotaZ8nTUQOmv5ukGim1ziT5ClBgtF5B
GIwldN77ZZhW4fhlDzn4BukDoDazkS2GZRqoRXNiP9Xkb2Ye7XRi5tUgq2Up80MmY+UnWEIdDuJP
7d/ctCsyPQysTiieEkm7N6s5V/NMK3fZzu/4zub/diyMFIC2ooLtMmG3jM/bD9zDLraGzcA7BhOl
2ljxbZR8G+8KQ9hHODM3mVda/RDITGOwpkJAqB3fZZr3SC6G/6/WI0hj+lFehaVhi9ARv6dJrc6e
eRwGNAXEzLft1WAveewcTqofOVNg8It1RdQehw9plImeUC9Ly7bCBi8RpOdKcoZnnNjUfWbZ54DH
m9kYwQcOdtpIFioouV+pGeQlB5lH6E/WhQ226Ex4O3evQ9UqRjwXgq2CqlJ6HgOKJcpcCuyhq+Ng
Pbt5MawjATf9Yp4baoRYFlHWPNc4qdXGhJNx8Mx16H3YnxVgd8OPQA6oId7vyJoZ5hgLBZgh1B9Q
Yv5R6mXpB40VYCRBuuQYTEMh91gC/hpknYTA0paOEQ9uyO2FzJ3DSBx6zKA77j9dmsFIx0cT10XS
22Oil0lgI+9PK323S1ZySIYzYoPySVS4/P90HZPKZfuNmW3pojUL01H6227tI4pSpcg0ia0BhWx+
jCu38EyX6r+RHrJbkeVLj4JJyr/08ClzsmCl9i5Q0PjFq3RHogYa+3WDyqDNUn987tXkknZ9j2dn
sxR/ztogFwpXIAQQPWMtFgIRkgQTJK0RkruAZXSP/kHmuQ1IkYpiD5Tvh+lttqlyk4U4GNh1LCT2
knk2BHpcQvyiAyDnXJEPIOgRYVig1HJMVE47SwOvPxEM0RPxoNI7rVohvA0sfTfJmPyXt5sNwTET
FQlDj87bCg5YxmjiDJwsHXEP5YXeP1fjVzV0GQPTorqVDHd0a/nmuBPR+KWTzUVhwCtEYZYP9+mr
eIYU+uQaDZwfmBjqI2UlLuK6U9qKOKGoORpn/Asq0Q+sI5UdhGhhnsT29xooL10iIVUeRjWvAATI
IkwIybNBrRvbUCQJci/WAoyayqxUUGXOtr0LRNncIU+YXguxalM+waoHy41D3ljTGMedbtmqzs4K
PToK9n17omSEWayaazOPX6KMt7YDmhjcbHooAU3rWL9N3kx9V4nvTGLkkZULNJS3FRtXzBXbs7vn
YJuZpj0lwtcqO5anMv4Q4OyJ92EHzWf2XxKo7jMPB/lN2bz2md4mF3lqkXDf/8yLSIJh2SXBlG41
AjThSpUekaQD9DnJBaNDP3yesThUtu4Fsxzo1ofv4GDFmFIWkhrVyQp2BXf0iYB9+U2DqzEze0R2
k0mJq4F4wXU5rLk4x4mEPzdW3IwdW9kxs4AiqgglSawWVNp3W2Z45098HY+4T6Dg7B1IRsOfVdcQ
r2au5qkacckwVW6235M4q/Cu53W7UgQy7cdprNCADzgXTEPoms9MKXxhaTZO9JM+RDVhyUB6Nhpl
24JhAYKiwThAZ+dsiV7mRtiBH6xEbzmUsJby3GSAklhUiuBYSI04E9fK+HyzVRmsoW37zNSVfsCQ
Wxh2yflgBwsw4VpHG2VSMIa10/D+DH6A8seorW2UfqeuPY8KSt7gQym9AC2JMx0rUDROWiZS1oeG
Emtw9sMT6zZMQo16Bp9rXsVIUPpjGICOBteFdLDgQe2Up0dKCUQ9eN/mm44rIxrHcQ2bYs7qiZB6
uR8VMDCC1TAV8eBS2AIJ7zwH0WyFKYeW7ieTm6s+voa2yxX1HZ/bZuuG2c2C1OMVXOvLWkgqML3v
PNi2f2S5Ekweo5RtT4QIm/I11d0voW4yA61cpH/Q01mpZR1aFJ/cMIYFKC5CIYNRN7EhpksH8xl8
y2YIGd9nZrwdp8kjUmK6ALPhSOAvShWrJTSoCEZ+urf4P5OB35WGoCQPH8jF2d2Qan67sq8bn8MT
/Yo/qbnMGGMMMVYTCTta4gRXkAGukFTvwrBmCVL4f+AWuJsojXRwkN4ZuL0sZiKJt9CZ957KBN4a
yJ17oskabZV4zHQ7VMkQI5pCjF/to0wZEG6zfQNG/ufByRXKQbfF88aQ+eaHpMkCk544BpliczyS
oTXw5s8OvtU5rBosdBpwXro1SUhIQH73r2enESGGHjAFSCNVaesUVnaGG4mD2GYoxss6BnW6Sy18
KbxOrUHkvAMrll+q6w6sSHjrlqRUHetEw0Kjitp6hbSr+gBJoUThVyAAC4Yu7EEAYHJNQ+CM6vNM
bNS7uKnhrUe1JbZ5MiQkClcHPDJp6tKnYzqS0y1YxfPXCvjcNirtP1jM5/XEGrscpb3gyz2pq9PJ
2EhmyL+tsll+n3Uj90S7vH5o40xPIYlzSXzbXVnLyJswevFrxv8fSLGm1gl9AFKE9I/ILxs9h3Rh
ZcLm0dMNG+5saBErYKCfU9NRPhlHbv+ervpAHPdaOm7otyINaym5dNVNQ+T6MaLzG0VN23ITHehK
eJLJbkc/0dynxEKaRc79BqnCMf71Jr09WBywr87vKlwvPaTNLEV6zKTd26TW2Y+7Am6PWCklFhOJ
V8OQHl3NVnCXoMt9cVRVKCNCvHnzoRNcL6kQi5lHbxkMdrUO9z7XRaAM5BbH7fZsJgsZ8R4H4hLp
6zf+Dk+63aee47xvj+k9CcKr90igh/wCCfJOJHy3L/9uiE7eNG2+mGdI9F4sRIr+vDcBLgQ2sAPH
wwgKwGRxJwsWxMWwZNp1DOqW/66mwCBntIhdVEmG6RESuZv6LtJfGvHKAmm8XnCpmG7lYdxH/R+l
bLUaACm+3HbGZ1jvw1WG7BgbvRMtu+c2cTPdFrdol3JzWzAH+TfGJKkI0bXFvTYwOZP2vP0VVCcZ
X0qoiQlVFvCtY0la6SRqFvvPgpghhkfxXZHP3eQtMt0TYLjDbS+8YhK4FXB4NvUACdnK6966U+Ts
lCW7ubGVeBxqiXo9YMTUwCUihcWyvOEgUgAcxLnFgsaf2IPEcV4XTlzxLN8TtnLbR4n5KzWLrilc
hGhF0Dqkho5gAE9F4TNUCiDwegDN7lqXXuK/SEZxAXJxU9/8OYMUzcDBFDN5uqJRiQXOvbjNAXgb
veXyosw6uxjYfcvbue6qbQ1CzlIXccR1Tz9UptkmMMNxvCQMwGc7mXXqa3lTMw/HLt1El9zHXrB0
gmVsSvAMNQ3BYFBtc0gKcGNUsGTTtiR2wPUrcwwfAwMxT5Ux3n5Ftt7ThjcxA4+j4RPMMNrMF5ya
ia6esEIEpqD9tiON/leQRjKeAbUERuA4Z95HNhsoMZElcso9D+0N96vBeNI875M+u00g4UsL+xsf
k57sCytjvKbqCzM2Hz2wuiJhu9Y5QpVK9Tz6EPB/nVPTznX3hNkLeTEa1hctLno+7w3hmVMHfJWe
z/vU4XkuXmBsO3sw3rLQ7V/II9Et5gRHA3pbLig0Ve5SSp3gtzf8wV0N05nkEOT43QO1V9r3UpFg
bPKGlw1SlgJr0OuxKwJgLpypHGP1wxL3dF6jn6nloJi08RyBSZE4x7WtU+j+w89mzPTiiKUko8EK
BybAM0mqQHIdMC+nJA+/ZnqgXjmQBZjIsRD+HZ24qGmn8xibI29nGDnaZlz4rVdCF7+xv7TW+/Wc
I99XX2XBDzGMU9UfchCJy7t2KvFIRrdU0h1K1efncT5gCs3agv1Lb4/0jLrXf8zkCazhxZ9WsBpy
qS7tvLDCsVHo5EJpaySUW280WrOp4FwBPwyIctGK/0D7ufXyOYb5iPlkN3zmJ9mIV07GA+l32p4J
0IEpRKZbJVEp94kchPH70B0722n00h6igJDNm4ITl0H8fYg3F51IbL5g9FDTMkMzt7Eh78ul7NuH
SpFWs1JaI7I9ILT8J5Ix6DQPE/OHkYgwQEFE4o5qGO32xsYNG4bbnyVqJSgynzi/KKWeMVYZFnn1
dziLISNioZAwTI2wskOyqyBglX2a5hK2gkryvYyMCfwasFSI7hsf7S54rGa/XeX79ahmqgSVJ2RC
swPQ9nhC6/otmjbQHR1zZwufVGfclRuC2tUUSfhIocQ+fM8i8RiFRNYcu4GnjFgMjKPowpmHrHM2
1VWqoj4IdQGESQJfMN2lTViOivgxtgwD/sN4oo1A2IO0YWSuHHHWAth1wTvhn/XNw82KdRaTG3Sc
hGdnVtnSJvzEBByH9AceHWkMUISamssTkdQ/+B5nmdPI7cChcFc4nkXcu5XP+kfH/e0oHaLf0NTv
Dey1soJkk63Ky4jxDZO7c+T+9HZjWGMqmDUns8gTVGJt6hJ6MKJqz/8xZcC6AvUJcrZ4Z4zgut1T
N3Ents/eTXZNOn5beCqjSTnbN8bpcRoSsIbw+Qqm2m/h6I88pBwAY2g1Mwt8M8DfKoCL8w1OkFOp
KPEArF+dGGiY2cNQz6OQ70GklBqLDWCA2g03bvQ3uoWI/MT4/vx33r5pTUF5ICPIgL8kNs4UjVJB
HQU51o08iwNO5jiZyMo5oBAo7ZXRkfx9A8JJ8ChLen/905Gucq1N4ikSoQwqnObE2S1N5Hm6cVEH
ogb+xkciXN7Wgj+F6+iO3oo6lUjaOufzzC3l+zJ2nB+BOyCV2rrl+HmPl+cvayTXC/dxWA28eusZ
Kw/YC0ASvnKA/LKQIFImvEEBcu7dEtLLlxLxs+F+JdC6DvgrIl07qQNXLskCtUJyI1fEfTmPpwxj
LWx4uswsCJCW4mogZ7IGixV3zCLfkwKQzri28U/zFh42idffClW1AfqcfIOpFWQcwcBIDROJQ0FS
gqTk2T5E75ilJDLqrIF3c2RHZ9cCE6Do6LcAKcZTXg74/hB0IIEC58kFdrjf76LUmvVoXnnA2xjb
zCkRuKu1x/Mh5B11mANCXBQ71Ez5nroHJVbFSOZlAHm8a9Re2grY9TErUwBo3/3Q9t+MJXIPl0an
iAqXnzI+v5ISelQ5iMRtJQthJXPpoefYWGeYN0NUxW1XpDVQq8kg/BthMOkDVYoWgTRbG0SnqpdA
2Wk1Ge8Jahf9wP3+IUTNIQP4AR1FtRu0o1cJXfUAAJFONt7Su52d0Ka3n1oZDM3eIy1yZDIWRfba
4ZzBm00UFuq94QRTQ4CSSRUIvGSy9Yc+wgHNI/1wvmLpFE011j7g6RkRbwZumQwGqwaI19N2EWSW
fQXJd8z5k/N50S1vUX6oTyKvkW2dtAnBOsStRTZGibkylxLXSEp7q5xedp6dakY69UsHw7VzQF4j
05se9MCR+Zd/mK8A0/ukkcguzUuvMlvAST9lhBjC+HzMUu0A9zxWcZ7HArY0nlFCjfiCXzXgu0YW
l0t16P6KT2VdlnRhi0PNDhX7UrnA/ulUW7KM2ZJZmBljylh9w2LcstXYWfZYEMJBSBgPg6No3FAh
QDgBbg/g+yfB+EjiFW0sxQUfc1VgMeJ/ltHMZdOJQugPfh/XJVz43JbXwpq+RmcxVw82erWK5LaZ
MyoYT2T/SrUKjrUP29uzAI/XuWBXGKEMOxjgmMBhVwRDnffbr4b/vMeAo6oDI2/Uic90vgMK2uKF
8Pbp2ilaGlnbXp5Go1wiKqxEPsM9GxkcTVbMR6Q30vgZvg51ae58kRuD6ygEZOSM/q3H4fvn9Wpq
PYI+iIgNKrp4AAADzRg2MCNxAxMcg5O+nAbnMIkI9/CyMV6RohOuTbRGtwpOUfImFkWwmnT+WhAJ
gQ2SWJufkX6I4PXk76XqxUV/RukSII0A+hcvTRgDEtQqwkZhqbtWKf+BX2wX1NCxZmOJvC0q6EhS
FOkDCTC0bAD2t4eotMSZY3propzXRGZwDA+O2y6XXAi+NTXqI8OLV8JrYAcjl/68mME3Qwoudezg
LDPyB5vrD1m4OEQh7EL5pXpKCMtr8LqVq3K6RNl03h3G5is0ftDhz+F8keU38ScotpP3P0YQBvGY
Yf7d6SSblFib2Bj84mb+bvGXUcbQQwM0eGZsYOgIqMgRtzNwRtAeWbG1ZuAHJE9URyPdQSfkoPsh
IRcOG95X3IyKPTVXLnnE+Sy+Uh/+78/BvqcZBkWhKUJ6XAn7EFlGJS7zs3ueKDPYK5fAYwi/PWRd
5HqcvXuFy35SsUVw0FbpSz+/+ugTDDl5JYf6qR2lgVJpCVRK2c8IX9tobbftefWEASj12YVCTOm+
TALzAzU/KCRVilsrusiQIefhzF1SK0liGD4ZezwuYwN6jQe7eyAXsvh7hKBHRjqUtbJ0nL6Z4+gW
VRv2GqhU6/COvgk4qkO81AsxJiKJk1F3E5kKJ4Upp1rgTclE9fKJIGPKPSbU1FjR9F8/19aI9Yap
WU1Gef78nz4O8vORTymAvwMItFcMeIWHJb9VCjECY02KyuneO6ungZa9KhJuqK2EiGUL/tyhpXyu
1Y/kSoLz3EaR7v4GBot1WQu/4eGy+f/rKhsPaoIwLk4naVI/PO+huLWVgzOcLldytv3m5WMwTMab
/2JDWxl5IdDiE/kTLgBs7oq8wpP7DxoG9CwZYnHhbLq7CePt5xYNIL8BZ++HFZFwsLt/CYjlWuqR
qtR+Q6m0bdSmUcqoXfKTOJP4EtDkLPtmnlNa96TkmVixdfx5UGr2qX/IMaj+vAqjCi6i28nZj648
/wAciWlF6NZbumgqUodVS6NBuVHE2J/CjAbz1cQM2pUnMwrOchGKwIaCdWO5VSmboQ3xnU2eeMdX
C/XA4ZliBQKVgakarpTReC0Y06A3wTWUk/yJc320FxJjSTEeWo3DSlhmhIjJqp20bjSec3s2DOxR
PoMpMRwggjaJ76Jwnrz+x6xweuYZUZ0ar18mdapm0/PbfgfYFMArryrtqw1TAJTGJyZrZK87IWZc
iYAPbb6JlUu0btIXheiqsBHjJ5Lg+laf7xuww/vdOfgl5sl1uiLoY/cOdtynrT6nc7+lDYBARQrt
/DlKLKsoffBVlFdMjbqbVmcXUJ4XvJ+1yjKr7TuwOyBCmRsgjechfXM07k/ioFchD7G65oSVkjEV
dN7BOOCDDeOyn7/xJs/GmK6jpT7yS6TaXhhWpVVsMO5cgxupNmVZFu1Qh+r5BBjMX6nvK05SUAUc
rPoC1yyXIBzjMRoTjtRfczFsT1K+cvPjD+XUFJne7MSqo66r1CUBwMHHtJqH26LFTW123EdsXI8l
QOtpB7uy1k+ijvceRogx1Ba+1mbcqW/TK59C94cMh6KIa9trBqyctGAcxmOYpp96gG62fLHIltCA
ynLKXs+cYuTHMJRH289FiDtoqBqnZh82vHUjF7N5VQOTLBL3FioeyPCIOexJR/59G3ZSj+9x0IIK
8c4IiKrEAyLQHu1DU2v1ywmOj0tYhVLHopF3mvKE3ev1j00/q6ZIXMhVE72Dfwzp7SJlcqc41Egz
QeXGy7Ez0DVuCjYdkfEIzvjT3JWx0MSW84Xpiv9eoV36OYHlyl4mDcxcySSR+b7UD3n20y5IIgY/
g2ki0rbdj4GKTHyF8xB0i8LVFipQ8UhktnDWgjYXt0a/y4nyw90rhs0Sjp3tQC0weCdHbjHAUr3E
67oBu1SK66ueL88DGZe4iIgQOAnnlQCvAY6m4RJYt/eZ38Hlm2nq80Gj+YrVLmaNhIZOBdTsiZV9
W3eXVOk7YtPt9wIC45lGSQlBz0ySq+7bcgHltp+O+tM4sB2ADZrZpl36FAqDEIM3SqEJWIWEpjRv
aJvuGm5npbKixhKvUgBBDvXO3r/JmfFm0AX7mFYnUtJW19U9L+eR9EQb6xTrIleepSFL1JMULzcK
KD728tuO4YCRMtvm8BBsAjQoJnbNRy+4OUEDtl/teP0WZf7KkJYy1C+uSYTVxDtFqPRJcoP9z2Ms
Sa54A926V4IF29UmaeoVQIZBwrSZreNSGdj5OLrBTG/zdDhCRnJPPVg+5AbRTjnCisc58zsUuMWU
qspJ4twFsN1rbop0SpBvlS0koYX8e013FzoL8F+XaC+n688JZR8B3IKv/6CCPYWHUDUXdhSxzKch
z9PYWx3J0LXyh/wBZD2Tw/fIlarEi70fe7TUP1dAIaNnm1CcBhnHblQkCm/AjFX+7iVxOC6IGIfV
QqM8kLeNGaPUk1HhwreaNLtzlZ2MZgUbimFsjm3M20z1Xze6KPTJdh7zRBtEf+sM33lf+EHzVY9K
JpDM8bFNARWTjhkm6b+IfMnB4QhI5mnsJ9J8DB1w+CHKKY9hBuv+h84WgvzWX7DkdcjeSd5C3BIq
gYdOCIM6Oh0uc7Zrav0XxcZGdaRR4dxExhqG3LBv85Uf4NNVJgAWpnf6oV8ro3Cxc/e0U85PFW8/
lFIAADtTy+QEjjCQIul/Uo5CckGbgNBzgGL94yX/lBQRrezC3hUgpLbqez/DCfRmwYSf4VXX1LqQ
WAtql5xxOqcEo0fhybSkrzf4xkMDd6fNUcie3tQlrzx3p5mVtUb3bOMViVKd+Pf7zO2bpvqKKv6k
xRLoyjsbLU6FnycsSRRHyxy819Hai8RI9Ck4qFEWXmGcnStWyQ9+owk07wj2PDVWB4NEkXb3X6DX
eo/1Yv0X41Pet2KR8x5NnZuKv30oNQhemnq8lMadKrX/5QnWuCLieFoZm72PW5BqMfMnncyiyaD0
leUNPlb3sM+UjOfbUeV8mCQhov9T8U38/vhkit57rP0f7dAaVwjAunUaN0KbRR0re6sSkPBkaslg
fGTWxYC2nRFOQqaGT/9CFRj+UscyaFA7rcNi7CG87MxdCNnRzft9uyi0rIpIVIQV6z37jG2TKGFT
p0iLF9AsYuzNouNvb/Iw9U6z+g/KzbylCgL7LkQC0vFAqfLZDRiCzU3zJBWcG4DZuQsTgZseqolM
CUFmdirUfdtrlieYI3dlAYtx2DB3M6mCkQ4lDxvrjQ/MI1yRriVlP8LeOkHq1UwQv4ly4bFTevBK
gTrqtc7HdEzGuBMHmtI2/4+82oCXfwaQZlocdtqCr8+MGsiaLrCbEJmJlMsHZ4wPdtPtkJRlw51I
0mL/6k5WjVyNGZehra3Zkp/AzHwULQUvHICRLgzakstGWQtq+Q/Q263s8BGIlKR2doBDhUPaA4hn
NG7UUh1O1qWUxsSIO7VRQ2fsbmmFNlC6+Stps75mfkVTpXLR4Yb6Pof2MmoVSLGra0b59N3TFtuY
KZwY51aCulLf/2G7U59sO3kwiia3fY4WUeKGSl8NHLyP8J+YJyDju4mMBbX6lMqumhex10zK/I69
m9CSg5iQqYOs+LziBkERRu1Pxy+KC4ThHUpJJ9UrjVYTsms8lybOTFiAHQu3GFxOt+hRcnBpqvhG
cOktJMb1twaahzVZtePrY+i34kTGP/VhV0TifyRW8Moq+U6lauffbUx7grkh6GBTp6GQZAkqz8zj
A5iI+y5Jt0GPNjQws6R4fpuRuUq6/Gv6hekoZjCvzg6MTqFQ8NlGG++o+fFnZJQL6dVwUP9TOuXU
FKX73V3DZ6PKuI/Kpdune/iSVEaHZlYd3yRYFdt8JryCzXaLUsFM0zubDWXKMnXYAC4fsvQCiWxr
Gj+/J9+j183zU0CsyweruLRM6pQXZlin8wrf2NZEmwEL2k3M3h8xFIANa5jId3IySy+/OSeZFvM5
SYQkEMKRazII2K91Wd1dB/ACprDaGs57xELGT9Mi3PYhKvwjDkFtQ58zRSl11x+O4U6IAJhM/+LZ
vYSSRtp49/8WNpFySrZ9JhPVXEPIDGwTqJWr0Ww4oC+58GJ4HWUvy0GTNguubT7uPoBgkojZlsKm
CyFQbtYS12N3iJS9XdnoRM7J3xrv9DKnDRsAj4BZN4+j3QFMV6Xa9jABRoz3xSSq+XoxKXAAKKUw
YsoyP0y+ML3AcwmgZKZiyagflX2n4WRJENcSvM5hnDVzwNqh3IiUGyuopdnXnOSYOGlfaTyGl2Mi
J44b/u/ep/0YHdmpfwU5PzsogxJtOR+MhqbxDEaQZp/22042zLr6QA4wlt2+ZTTG20eWwFOu7yh9
BwMdIRyIHbaTaH4Zr+4nT5GK5azAoOT7faXMxihSoZ6UYXk1Xj8r/PqswFYKN92fpTz4kS6GCHhn
/xwMMnPCgPDuv6DNgZqTrxm/LfZiIbtK9BDm9aXzEZyto6gE19ABeRNuZnnYW7jYaffJuPuUFo7X
NWfmKM2s4TGY/GFOid7PrwLLZO9Sv4yicaKaqzRdgjb13v+X0IWuQqDOwj26bQVyKK3/CvAisP1Z
lulFH+yG8r+hyOMex3bxSj9mPxtwUUwjRDPzKWkWfu21PwliVVBcKfSx1/ddOQM4uxRjccCKYKk0
9VBfJzD4zV03AVva+9kwUYvBk2KxvCu+r3Ua1sdITcmERi0cQag5kMJuA80bD6X+/LDIx5LmLwwr
LVPElPl+4KHzT/A4psY/ln+HNIAzZo2rSAgT6u37pWx/EcBQMD84h2h9kNJVe9QWNjk0vY1KLQMg
tfC4HNHCF64NzSy25DBa3bHj9GUFdULgAh2gYYcmZ5xQeoNxUYCrbb6eZ49vwa+w2F2vKnR/2yzz
F+aKdDAErVeQQTqyA3ecHtH+C3xfhL0vNh9OfAQ8CKT0ulpSw2Br/dxoLejPFgVvQi4gNobUo8jh
NF24RHNCGXV6cWnv0nldB1nN4f4JECxGtCWZm43NKzSsNKxO46+7miu++QmUOKUKUodPWH5eaqo2
wA4BNISRpC+xd0RqF15QJdRhuh07Sg5RDVz5TbElbBMC1Qq7Zr8Ygh3FpBzR6HP5pva47DqOdcK6
azTV7tHTJ6+W0SU2tN1ZPKlCde7UUpBMtzwnFuPGXk4xNP1IEJxJwkO38lRSjDMTQ0up3MqCyfpK
o0hfaZGmRYaE/owni/ggRzVOoFbDGQzVFUJLxb0gJlrvpjB7z/Pa5hu7+bqt4+NcGUl2S6jkKxsy
T//zdP1G759IMg6Wm5ow5M6nhk0gdTf6a8T2H0xVja6+mzHPNzqk9Nm1rYvqSQj+do3fD9Deg79N
cp7iW6mwdEGYym79wM+F1K0YZpms5xrSOhmTydRRj2FCXwp0unaVTmH1zoNjdvu5MJWVkb25Kwka
reDRFRrylGhJrCeOPQ2nlb2eHaD0lChvAmMb0eMCYHX82M8lYk6FwWSVnEI4VhEhUhFOapab8exn
pA0j0Iwac3m7Kf5Mh7SwH8Ktq8eSEVHW0CCp2IsfByld+MEIYh7F2JxEH1iM0vW0dE844qp8RfHy
W0dFmQxfjRDO0OZtQdl7/4FyCakuv9Hcq9ye+ahnbM+P+/CJ9dV8yrQSuHaWi0Z9YQr1veudK7Z/
ToL8IcCfN68F012IZkScRnHn3/TZRWIdUuJskISqGgFOP1FVOoOtq/EgmQ24MmpLhL1JN5mPn/Eb
Uufxa7XPXCM6JgCZlhvTf6EvBGZ9ugCmZ3HIetqdHMFkSAKHDwM8hfHSQ+F7rI4e1RSnohC93LEa
sjUr3dLtfwDuzmDilJeOV8O2jdo2I40vaS7aWi7y/JpjKOntyonPC6ySNceAUsEbf8ymbspbEdpR
1SMPDDcQ7xWxoBrfcfnJrGw/KrNuQnIADF1L0Hy3ubzBBy7wiPFzKDegJakJk+B0v7SKk3tpQEIy
/aaROru4yqiWtQ1hvoRplnba/WLVFDGsnZfS045e3vdg6hDQ3g934KhApEGrENSfqvy1E5uEA54R
VEAv81hCfvd9iDHggABRXvYFW1De5M+PyWbjshWdivHFr0E+S8DGeRSTYziph9XIwzR3AYHLnwc0
2ErthmzraP4PUOuLqO8hUbZTWiNnSBMajOBmoDWt9qqgR6/P/H7hN2fiu7grhk1sSyhNrOv6uMaW
ilLHjIsLV9vN2LoZIu3BKEogCPDiIOwWqxSXzUmWwUK5oQ0bejMLFVsqKorny244wfY9DnGCA5B5
XDFmEYIvlc5t56ESVIUHCdTVqbHN2kUn0yJhKlHqIyIaqY7gjFBLCV7sPXhlk96byFOtNsUK7oW5
lk7xWSUBHVhWTp6gTzq8jU17aFw9WHZ7wa8JebcM/GkPGYfa05tZ4lt+pYYvOn+k8fpMtp4DiMLs
bU52LGQTOaKteo0QYEehY8EF9ejx3MfG3VZwGSqXGmM68IaS5GlhTSlemB81O0gfOkskbuycx9S6
fkCxZ/+8/wPmFEB+1/jCC+AuBCfqqECNWPdxLNq4Ax+gERyJbvQZDsmiVD3qaQb1up64fXezyAp5
15svZ3TdENCmlYrvI5yIld1m68fHYmVom6VzZhkl+lFGJx7dPy9tr76QOkf53/MxCGGHbLqRgooX
NwDxBlk5TjMo4HU1Ia6i7RT6BuSbgmTSDMSq0EjYn2W9bElc5FrNyCOyLSPbjbhj21lDyOdUIzv/
MpkUwCfoBGSeAXdaomj4NF3V+tdLbB9gwUoIFPsGj2XJ2jtj0ld7ryVDpzele+7WJTqCS6l72GCK
+4D5rYhI9Zb2Wl88waIjCXbth7uNShXhNAD6/fR2/N+KBtSIMpLQtYrsPlQAYjTJrJXEMSPdPyHS
0PIOl0sAh83kMO0mbLNk5T2h43x8ywneP3sOrsTyxcw+BWt4rbxBem5JHVpJ1NGnZ6kXrEtfjmTr
pz9pYQ50UG/EQbGQfYEWUFXoXLHqwgPTIUMuFxuiZS9JEZAL48K1OCliI7WT82KlLhD7mHZXmjgd
b9k1b6D2/Co1nebQOeEzY3Sw1nEYzrZ/MgFcCBFKP6PI3tLArrGNMH6gxPni4LU2X9TWPVtFI9Uy
cIJgkwGKecxe0z4JVY1BjfloPLO8VPTrmwqGQcnT7p7ZRP4l0ddhW6zyERZp1cL8ycvgRTkp/l3B
oUgE7oV1H1rnUy+9xT+NqDCZznYv4SMDNgoxHxlWpBxjFeFeX6UHP4+280z/2DK/e+cUBRA5WCpU
O1ldqDgoAiuG/pznCgb4K0JPM4GZjiVzJHpnqZlzvp48+TGva4RkN9+ljtmbUqzBfhXrxvefael4
gHwSSxludgL9P4KV1HkF58YMcJcAY3ZV0nzYXp/vGpY/RO0UYel6DpRPJqBOxAhlAlYusTWnhNp/
TYIDTXH8ZzUO9wRcBRuVwfakZMDdHxhQwKkUK4m68TeyuNesrQPBR370KXPOUNSIUnGfNcCN06jL
kTKZ8vMj1RJouF6tKQe+9elPi5uMqF378J7PKRQ+zyhOFx9WOKBBfF8HMdjKFE/wgG533sn60fds
QWdCzgr3+NFozN2b+TTiMO1GOOi9Cw3GsJy/2yXBVFEykUdWBOOqwdZb14fAlZNawAno2zG61Rjf
UkqT2zyUOEbZY0iDXwzD9hn86wxr7sZy2zli9/xWzAYnClyE2kki0QY6Y4No/oVAPHGe4+LL1FBh
mq7M/34f2PtKpjm5k83llhnVu5BXQZRh3fG4VHRm/i9f21LgxsTRl2yddVV+xtF84Xp45zrOraLL
vsNyY4kcbNaVdRaInxnEDHyABPezvbTLRrzQEMzh4NCLlpptZa/UrPJiB34FlLKkyNPkJVRWNZjD
G7ytj/I7RBgBbdnZDL6/E1dWxyeY50Yik/gE++YrwD59WDxRl38Rd/wIx1hRZIKUC5aWhy8LV3C4
D1e6JQsMjxWn9kOa5clHAYW1pICEPBqq0ptOtoN3Mkel5kd8CssK4bF5XZ0XJ+dQsSVwGYJXCPa9
hreCbh/2hXZesz4EiJNpX3wUpGEpSzp4UYphcqI2GxWQiR7qULyu4fjaHSgDapVd3qywW/X7jWXo
8cDorfJmHtnWsvyDe15Bf4wPZD9e9hrwqBXrYqpa8tP9KsKdRZIs4g521Oi0dxKehpkxpI/1XYE5
ZeKLEdQx3OtQi1PYJSgymRgpbwLnaEVlGbmsc/26Y/C3EnOsqOBYXL5yq5P/iAuZ+Wgi15x9L7tl
dZ2Bzs3sAY4FH2S3i6Coki5qB8SzUkHrhqeW7gBIHjC0FWjvW1AUCYQOWkJEu2EXchXgvnkYSmyn
dmPuIzFYK6qFS4Hg0h6tqdYF4g+x1oy5g5V2OzxYp3vT99thoGkWrZFRHw/7WdzMQ2R/JPinQc4J
9QHVoB+1OaCpaP/b2onO8YJR2DHn1PdyG4AzGEY+hdjDjqe7+ett9HDIhfwkce3iGltidk/hHOE0
Mw3xYslDfgZ3Nch1V+wAw+bzSwGtRvmcIrZQJSVFniv/tiAGnDSFotluiggUCM63iFVRqhGlCwiO
GnqAadUdBeYRS50Me8m9ktSA+/yjcuRuEhpGlywDNgZ03wcTfnVP+pOLdwzeIhWlM51jc36IjE+v
ubmlvyoh5aziA7YLteGeQhwxIumRvO4hQV3dDnHIiVdfOTrpUGFb4nlL8Sna2tsvxogSmheYjS1V
7TZ3NcCbuCflPhZWlBEwU6NqwyfRspcDaE18pgdTPJ+JV4OMlRS0w0iRuOOucqbftlI//0e9Hq27
38ZyAruV+zvaPVmXoKWBt2+eJ/WcUAnf9qSf9PUcbgfLHogznUq3OsjVvQPJOnVYXw1F8z3RssdM
y69SfjQIBW2IUAL9YdrnEjTDZsQto7SCYng99sHOzetFI9kbtUeNTc6tFjNbP2xHgT2qc0WqnFSz
AMI8QjDcmVSsbiit8bsbHdIoa0cXZHbxuON7w8TBq4JnPRSGb8SFSkwWlwGOdCiYGHWe4LPCB3XH
X8XLzZGijdPRCuTz53tieaJvdXUFfyaB/5dVBKIuSnPZNv6rUvwZOGUO6vKOC4FPzHQTjuCB+70J
qR1XfUY+BUIwatKWjbjikr7QgtNHyGwMjPfxLDee6LUQ9gDncoqjR1AMKUcWF8StuRub5eVSKOJP
3NEqQb5XyVUE6xxTXk+gfsxLU2JW1GZVYFafPUUdcANnP46akPaMoG7GcsmE6RrhrUC+x7J9eo5H
oZJPbldd0otZxx22Q38AgzTyM5eTnaoBDWTw1wfjHE+MvrABTsxLorlcTHzIw5h7fM84sKApxz2z
vOXi1ef/P2en24ZXN4lGGm0MDjuGHumR/904S5naX4yOt5TcrQFTimdbZfiYNeJ0Ez13PiJ75OaE
qKRU5cvgisL3Ui25oKRkhEnhnf1baBrOaYpRNORA7/x137YnMCTsklRX6qn+JPyomu/bXw5rZDGe
Jywz2Wos0sFRP4RwvLTZaDnCXfHhlVW+77HVphQb9WeCVMp2mrmC+Ye2QpKoQrvB2JeEI1ln/dcS
XdjMbarn/10TGSOXtDMHzjH2rqj9kX00JqIeiIxIU9bmWJyuXdcMYv0Ay1ai82c0tqA8AYZUc8X4
JtBXh7HWPBSkafv9JucCZ9DI9HVyfG5pwZ0v/WPPCX2r9tVOyOYxrM/yDcEHyoXllByEzhEC0nsy
33p1JXoBAd1BxGvpbeqHnyScdfQBM9P5PwLU3dewOZP5LL8TwubKMTRszX6HdkOO7FZYrcBT34pf
LEYlyQOuWruJRLy+bDvlcHuqcEHzDjTd79zHrz2xypLKZvf8rm2Hpn4S9W6f5+8u1Wog1+l2Qp2Y
kTAa7Z9cZgr1CfigKQKf1Hw3GIbutRErCNvl3Ofp9GvGc1Y0TmqjdWdYBxTn7F8VKYHxGcNb70vX
3haHcUvs/o3yRUY4r7CyOEvPr2qv6eWMT50kmQOkDiwe29rPGPg+sT/N2SWFN03uSoB7ziewPDDv
B0813UIbfs/fOsOe2+jsgrAk0LbIXPvzLgZ7VXDHq544PEUhtT6MRhn98KWOjX5AimasgBusRMub
4pA/OKX+DHT8FClGyKuXeYLAn7o+LVBwWPOG574YU6qNM9anrS5GohlBBrGhfPgemidkXSDdXVBO
1TZ7QlDji+GHA1ibp/tODZLiqtbj3+OgXlQI5ZWTmxH/jqVw+PLYlJIl6vbV170TGPpH8NRisIOx
s9v+lakSZfdwIUM/MZcuk+WcnkMoWmLsE2PG4eM2QWM+v1ELdn7karHjUd3Uw+WtDReSoa2Zv8bs
mgmS6zlUs/18selGGd2+D40EY/yOeiTSPiGrtZ5hPaCJPTsCHGJIv4kpqf6jThXaSQ1G3txVrvo8
ORRCPR1dg6vKEN6L4NRmuhufg0ydB1hnr8MNwtTe1AHYsoa5KmDDcn5d9FK29vWMPURXbs/McjMa
MfaURb3TEa2a8EAq271OQpWq6kw2J/ScoevMnTsfy00zkhaHQM1dIPUAwNnOBmEBkelOTUtvuXuL
/0onpa6N5ftOnqyztPToxhrYwRcuGvbg5TAWXNqEEYhIchcunnxFP7FE26L9h1EUwdnudorqZzeD
M2l1Yrbb62hZyoKmSUGUo8ba9OKEqxOott7xpT0QDWG5/KIXDJgsbiugrCMdWPhaONeCqjVWa3/B
+covYu73mm19CCChajRDfEX8djxB9bEAwxmJaWZZo0uk+Y4ZgDGc2J/BYrkblcRjwgaAxGQi0j2c
6YheZAoMTlDMkVZi2yahVgJG4bKb7vo6aWMDR26xmXgmq+pUMFjOspQHbrBiAeQPQFrhwX5MOXH7
wvPC+l2f9z0jVW9B9rZHR2wOrGsPCdZs8KN+uCw/l/oaO4lfKXr/SZ8G4ETtpFLnsPnVhjztWqwx
nMFRDDT8g1T93lVMDD9hdd6Dq3HA43k26MukJdE1gO8rPWByDz1rO5aQgVWNLSPBkhNnxcZVZCq6
LXgiq92JIzIqUGPrZt0Jo5/lIv9RTm5qbD7U2EdeAoghacCyqPq8aNMf2whtq69suhND5MK0ABpw
RqGTZJ9FEvfl40f/sPBbV/tvVBrLZ5okTUpWVGd5T5AA3+k5QFVid+z/OH/iVWe2LDbtRw+xt4Vj
DuC2O8DsnJWcD6+1F7Oed32hwnqNedg/Yl9pXtyOT2+2T/sNZ9DcFWTslu4L1nnYgQy33ph9iPfV
b0JvGY29Gtp5stn1qkFgRMSkl459CogFdKvtMyTH8LsocyQYAivGtc543SJj290cJUscQFF0iq0v
jH20kO0i6e5WwdXNHS4azLjRh0pi2j1RGuEmRZHz9VfsDBe/oFeX9w0vfxH5m7//knSRxIO3d9Gp
VJFxasa0C1AFPf9tXn1UXX8JA2ySq6ax0uPDPE24qGCLRLfCX2rIDhWqh1OV1iCy9A9zdUV9swf4
RqSuyLQTf+hGlzMVzmCU2N63+RnRjdsWQc8eRxHSNiMVVEESe85Y9ktlKHJ+Vxlvm+IgzOHE0/Fk
ju+gaydwTnRJGBEM2p3hk89EobO2SE11lM99y/1QwdmDxKsYIePfbGEZPcjHxHbcuWuuvkHFuqKi
ZUYm8u7ZLVXqk/T7Ftt0c2HkNa9chFrMwcjEkAf21GPDfRF3Ehl2m8XJp9dW8TemVV1dW3qWg64B
QMZDyJtAMjXEa4Wya1jsMemIM2mimd88869q5ndvGVFiT5nDs4v1uSBe7W1v7eZCO9dIRH8xH/ax
zu2/VUOGCwngevBzQO7hnzJtuKtPMRX/Eft1Ig3Y/rea+HutBfyx4HVON/qlrbuacspgw0npNICS
bUPn+xpar2t4JVv9+i+o/hsE1oYAtzSVUxlLw2n3/taIZVRPcxyn7sKbxthXeMqbK2NuQNU/KWsu
JgbIjLDJup+FlT9tw0YxVyfh0IPSMb+OP8IM9xwlzZ7zHArrOG06ztid/NNNom2KA6YFTAiXNKq7
OLWZPLcSitc0GqSKDMpTNVhyq7Q2ank3+AFefWSiWKL8uHgzBNlcg94g64eieNQWm/H7zi1xPxvH
RUaPR0lA4hreTc+oF3JiFUvOmErCxGvyeArAYhImDwKWVdNp6u8eWV/WLyYytKg4W3WgIKcdkM9F
5RPhLarOjM3ISwdwX0zpavlUDg3igX6Z3yX5cFwsrfMBO8JKrq6ZWvkmNhkeaOPwICDm5vkkw4fy
umOOsCDBJqqVGps1nd3PYaBnlAwo7LK2/VlC5Zbww2rMkZEej48KQBOKNhtUODo1O4oTx4I+8T0I
G8uL30aSLSNuQH3FmwAGKZkGmJMJuq2CyujDPm9trqCt8AaI6SkhVfWlk+xs0dMqMveMekWMfds1
RF4yktxfsrts+7y8NAY75+omRtMUY+dmtsH2MQ==
`protect end_protected

