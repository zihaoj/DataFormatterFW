

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U25piDsIMFzypXwCunxvuy0o6hoR+co3yf7/JA2KaAWusCEEI+goaU8wI4Q9V+16atavXLS2/buh
ejS3QEMuew==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jsnsFusZNbbG4y3ibEA35Jyb1F7ZAcSlW37QVLumQEP/49516LdYfPA1jrs7k1hiLAW1u+3fIK1+
qAMys/QVHzYuzGCCF0kQW5U9XEzgYB/fW6B3FYf/5VHqfscu3JlErCgXT2qPTg0Fq7Aj1Kq5v3qP
6qkMtBzoVYocl6EmxC0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NoP6NWMp0rPpBfrQ9uc3i4A3LxQ3dpltC3rHIGekfFdrcOmczm9WdF5SjnBRVA8oIOXmMvwvxYW5
cGqIJvfJBAWBcK7gINu7Alez+M39QN3P6UxliEsA7rOXvPJZlfGZ729E8QGXaOqVIg7n1mPg0Gv1
lHT0bDK1IB0AJRBy02WKJaRnZYto1VfpXn6rIOGUZkMLF/QyvQxBz0I9NGuVVBUNxAHDQmID5GJv
c2KC8Qhy9tdLuWhn1QL52AgKMfalsABudapR84zHnnP5JsIe/MNPIFAyhqt+8PHtYoRFNuu/KRsI
Z+LZAW2MZM2LmxSSb1rzX83GvmUk99B0dpOaKg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZFj0qndET5Qb2QgXnaS9wixRp93pcdd6A3R8ovmdrtZh/NBxjFOKcXDZlI2aqXpeATG22liISmxC
fd3Cd/rCGlXnvfj1T9Fe88rjahHwR3OjhMjb1OWT5lgyRPB+3x/TrwX5m2fw0WHGIfP+/pY6Ag1F
QW2uJMT0u99CwVBgv1s=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oN3wP+CyfJSgK9oJXhhhW9kRRtVvo+/oxdp0oK1SasNc5TjjVuqBVA+KpkTkpsDApDXGR/c6Ud0l
3vocxPsqA5zSFRbe4Z2eVtB4adSTDFfL/+ZLeqx7kZcBeNt8SE2qKJq4b9+xoRrGASQeMgI8ZZol
MgAzR0jiT0X/lEQakMNmDWJol3PITZYLknXLm+9HJyL2S13yEv8spZiz92QPm9ZxyMbwgpShZP9k
XKu0O+jt0jHjQun8RvaFK1W5Q/Ka0/YkvfPXAswMKj2aOLTFQKtXmHhX4yWETuYU9yRKZ6oEPRpw
QP13P2oJrFuiZU1jHSte+uThieUL9yziCmnjOA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 144176)
`protect data_block
AdEs0bC5ofk4uG1x6gVOo9N/sStBUmsuPTanOIdoQok0jtsDZtlZi0m+Fxun2GHzgQbTgaN6KUHx
CaZj6rSG2rLQG59PsnbAJE0ieZFyyhe0xxon4PmS1Qh0T/UNqSXKdJkUjOI5ZNsO9qLPoqND14Vw
oonUj7Zm9ukJI7CqBNsqDXEc7QQPHYf9AaQ48e/qIa6xUQ4ncglJJoMWwttv8aw0FoBt+ByK/66C
x2JZUXMezcVFbU/yFG7tugIkmUerx0tJ+VuQ2/mNlOnnJ8PKRwBuANZzt3DF0Sw3GHqX3NLn1QZQ
5JnCANvdVurGN3kZaFHQTJkbqlr2QNfZVbSztcRa7BZHVAL09PxHN4u4XFucCMsUWsVYD8HPaHO8
Fj25tfu8/8jTaJtZvk8vzAf91PunV4B6MZ53glGLOURlRdmBRA7xpe61IiROCmZb91+O5uO9KNac
D0VFGbGYGA4TqS2zWqHC26y/17QbX+s8sQPulvVuMh8PIBDbpXK6PQSiEzNkc3rKKLRyYQLAbgRH
0uhs3G3vMSoxEBf6r8gRtndDIEh7sKJUmdJ4wpXEBgZqRgJ9pFHaua0NVVFfOTRxroswXmFlo0xT
QDJ2bBnR+d5BdwlKAUE9sQ+JLoEL+TYOiEZoFD7yJCLJ8BYmrpWEpxbzkkZc1iUenz4PwSBvnWTL
x473xs98v0q7Dyp18j6Hsnt7suy7x0YT450BeZbpREyomf8W66KdotyUYwFU/04pHwlavln6YT8A
NUPocuehZAcNFkq12TXUTXfuaIKQhuYJOksOJFW0OK2Xj2P502cEU7STjTBM2AeAvOFi18GvhX0K
nVio+mocIeQSbj4Z2P5+UouC+UYLSEUjzrqG769i+lvAI+01mC2dgImZHWRM9LMhxSisg2Jg67wQ
RhFC/grZzB4TSabjJ0pMsUa2IwnzlrO46PcSjeLuVix/sAGj04Xwd+yhNW3Q8Ih4/AfEkGWGtOKS
b46diUWfmKFi/bztAdgfR+HCl4GEil2s7oBZE/mXi9gCZ1oqn9GKteSib3xvmyYA+aMuXSQCGXd9
6WjVqPU+5D//opr6/7qMtqro6aHU5ZJi18LHB6OPLBPNhcibyMSTiRMSnJjO/NwakqVBCuPHeB7c
q6d0imk9vYucBHtUL65QdfQ5EKLxohMH3Ow72IOiJkLdOm1GEM2YkzM0Rl3DSaF1fNJ40zfemSCB
yafll/hfBk6rvLk8WSsOuBQdnxjX9+vqqBP9Ao1+zaqBSu/ci3K+6oFuVzD0CG1VZ3I0vmvqIoJS
RyEncOEicGboBAYSWdByDislhLyqvCphr8o6B7VDl/iIJE6+tKNjUYdK85RZU4bY0Nm1V5A1e47J
woXCFztBSnQ2bTpmxL5HzmTPBkyfa0ujNpTkRnVz+7i0f/onP32CO2JLxTv3/lO5zsmqVG/GOwk/
BNHSqvCdulTggdBSEWIl1q2nbFMo4LcEuOO4KJa+5GNrFrF1Kj48hMpdCG1Ej44LK81AIdijl84E
RqOhtt2CwUdviDqvDRz2FTnPyfJg9je9nTXVvE4u8zy8bMXWbAiL1a2p38tD2GkqkPw99k1ZD1/h
PJeXykCE17sizZr75AmmCflq/DfyfhYjYpCbcxR4588++bHzCnCRZzNzru0JokD/i7wvDvYzTU8W
KRqS73qIekVNknRalfFh42uROkhbr6Aykfu8mjxB5GwOFLTlQ5ZdrikC6WBg2xVjCTGYC8YAKcL+
dv3r2cRjMmjlayQwKn3rz8s+t1oblO1NafIV7mrHkFqBaFAF7BQyPCThuG7XSuzxkdigqAhqlj9M
tO2ojgpfupzb51PpRCBM0OAD2t7z378Fln+KprfzHi5BM7AXNVkNHIzqbQQWlsvvaijp7gKkau7x
q378S4QOkvqzXYsptUdOFurGj/z+orSgcDWGAiR4hYQZc/Itp1U9UIWL6yGogSntKdPrIpzvcGP2
5xxhQ1xCQZG7Cgr+rQRN8vut8QEm0oNLRtPzqj2okZdmkX6iOZgmMRC6iaXfhbyKA7tli6GR7Fke
AY0gpUfcVk05OSLzrd2m6tADgOlBQ26EIeso1J2JdfE1ydr36GjUNzIJ4VMf9txlVm7qF9Sqvz5l
mGty4h1AKPwZRYddrC9hGgZ9p79XaHhmYQr2m8Tbaojkkl0p1fhvYn9nm67avt+7Kiprc0RbdOHu
6lPc958xwoC8pPB4Fphby1EzFs56pyeAKxLRKudq44gO95qnKoQX/89diWou4AJrNxK6yA0cRl85
XcnnV9zD4F7Xk5UAWJMNdR9MAK0y2adfL4XxgRwzwBl45A+xo+kB1/LyBBRETAmKS/IPhFAB4p8v
ciJvCCMhRTUsNDlRwtOvINhfm9zZWJeHVOqu/+/HbCfkwhlZxgfX7onYbeZ/XCjHkf4k/Fruace/
1uNO4IX1NZZjOlQzdqTowGYvBFkflFGrBCgSiyqy/78AckCbeeYq2gHQvff5JgRxN+X7jx21PVgP
xMQxrjkzb3H1sS8vWJ5HWDxIYmLAAuSlOVHT8gLdg1/zjAu7nHoXhuNxXtLsLBUji3ATbZopP/F7
++sH2j65U6o4rJx+14xcBfyTYBdB+TXpugZscsNmdJbY9d6u1NtNA5rGxqp6aFDRFOuXnqFIfqyZ
8UIF667of8aSDUdDlEz71fLt++p5lUg1w3ciANR4SjtaBfon5p/zRsvk81UVw7e3K/RdScoo1V8Q
lCR88n7JwPd0uOlIcQtgZJUZnQ1aYW4hskEwPbKeXfpXqOzGKJ2iVMTyRtNlUPUJHfErHK8jug4Y
oONcEn0XxxmibSElEgahSX0MWwB0vQuMNtOTJKI2TC5SOjgXBPJbfnJqzUgv+23slDgp/sSw1lnR
hj4XPCICBU2DrdMKsxK1M/dJ8GK5zFwRkZWAKFtWRkKEb/aNrkJDGWkFIvIZS0ctd7E5sL7rdFHy
0Lb2YxDIFeibnhnSV7YdkXYFeH4xymdDJZCCCKLQzjjTevJ+6e9dsAofUUTrpauD50mbDB8f8UJC
O1iWmZ2Ng1YhVnRUQy1fcnBRAq39Gsh7dbiBF89tX/pCob/hJwwbh1Z6TAKoXvmsfyE90gNOMeZx
gZUaSXxp3H3KWVZeuhhsz3vy9sXWKvFCc4mxD2byd9VRpi93MUhMqejtlY71EwLZKYON/DWryzwO
wptR9CHFG6vygBnMgnCToLq0XH2pXZs3OQyyJVeeHisrKDD8tibXVZOr5atrOITsOF2dSF2oZVMi
c701hIkMWt21OTU6OZmvb7nqPNumlPUu4dUfzmpblYNM42Kn5GUVGb3W4ibOdPYtMIkiczJ8M43I
Thg2CHeID5wTIMSMgdAK90LSBzYb1bKRISHfUMojiD/ZOOSJuhvXQ/EC/9eZDSlEm5gb2CcVmBW5
yqQVYjjn5bTCk1JgMX3eXW2JQhhviYdJ7K9yRlhBz9aoGt6UfI6QsYKuh3Tp937IaoLhxcn6TLWh
OPqK1IJpRs/LnYLzHWFL0wWRXD3LNZFInULW3T4BkErQWFVpXijp4PxkTSdmpxVAKZ8anY9dDmb3
4RmBYpn63T08ZW/m3C1YuaO1Gi8OKt09zxiGhojRStH6igtv6A6nqPQN9AU2BiM4VOEimknDFgDH
sV/ZjR4Qpk7znanMRDUs+HGpSrBQuwMVZk5s8t/H0mJsX8ZJcdOu6uJIGZBL4mR3bf0k2OavVqGI
6l6wg/Q/DZNC/fhgHnNs9bafc9XtZ1vPKMemAMp9p5xW3pjFNSfWandIdJ1DB8kfe88f1fbVSe06
RFP/1rzsTH3ByhRRWwWV2AJH0axsWmYb6ypnTQyuzmVy+P1834KUE/4ph4SpLZkwBXVcdVh8EtXT
qMrbeQOSNHurHz+e2RbMmPpDa7pYi5RniSEMrTb29ZNwm1aH+dp/VYY7jTM+cAnUjeAinZMJnRZ0
Rq+k6HAoU6EGkGe+cz+x7qqzakpisvnt9Bi41BS8aXJuLrfYoOBj+hAiVkFCiSB3DKeNcZUZ59FV
f5Tj12Id3Pk7dX4YTSGiU18OYiVZOT1SQevSTP1aB3YfWbVW5LZOf8mGpnFZOS20qjIbvrBbbyFc
jWWfKyQKelNVDAWskGI5FjeHXaiyC0/9DLojEmHwKjAKjxSBJmJN5nXRxppumm2pntVV+DePcjV8
+qhxqccC5Wy9ca24o9Xz/3PfWTND43+cn6csa/Fnb8M/G9bHbx3u7+1fqLUg89o1rdngbfhJcIJI
l2dW1wLYzJy8r/bU1/y0UNjoo+NX9Q6e2RPTxPSouZQhAgnRtaZ6sRt1X4yjkH+evLh1AePDe6FB
Ys7ECRUKlM2ebhuDRQqjFvh+91B35p1GJwiqdnp9L8UzWYnLKVaQhfsr59HCkPnmLST/ilB2dSc9
HXQM7e/uT3TC/BqK687pJ4Nd+FXdQl8kReDDWaQKwZ0ZP6pMEgGA21RuEMaUG/YmlqQQlRQZSt/c
FdcD7S1bfGL8TAI6n6x2pDaTdzwgE0mz01AH/0z3BAdqmQwzUW+SsRyVsIaBfpJTt1JdajzkeeA4
A5jMrZTbA+ypp5LBNr22XXpRvHmcaB9AlI8Rz7d7l4PMAGLQJcP8qag6yAnfHZaEZui9ItxzmiVM
T6crXFtIASmlwLQlsIz0tqlAJ8OnkFxB/0nnA1fdeS6G4Jl/dzeEPdsRt9ux1iirt1i1TT4SkL73
WUouregvxuaR1937z09mrFH3x8DKlML8BMYUoo9e0etu71sLQ8UR4WB6iBhQOeUYI98XkRUzYfP/
5lFssTwJ0TU2EnrhsVqJX5i/uGHRGDVeAMSCnGKrLni/lSEGv1Hul9YiGngiqayqPLRjKJ+Q3btX
7CbT+Jfa0d779NcFcp4ntb9ETTJjV/HY54dv4+Da/BarR7IeSSsNNYg/+g2H1AvtnA0z5uLYIjA6
ftTtXUYyPVvc2RqbYAddeW+VlRfbMmiAP/chGMyXTXQKcNjGxzuIWiVnIpVlqtKL+/ORU6pTxwDV
o6d98J43NEdKoE5iiZ+d6P7mMMCX9KFD88k64GIMZGziqyuoG2M3Wu7hq1rsWoUPWC3uLZBhLAja
43bhGdJuZcGQ51bzvg7xGSqR5bjRQ+uSXG4XsGVBjQHd3gjhUUiGdt5QbwPBi4XATN3G5Wu/317A
dRmxSZ7JgZRXJVxSsEeEB0gzI/fAK/dl+aAgYpEG73j/J0kPQbFSN9VxgWkG6/g1brQSEYGs4i/j
/4qIUawEgwCipxr+cRwiSjxQ7GQu+ntR2z90HLkmTuWBQkDzVqtt4VemurhhzoyTkZIFfbq8nNQo
8n2zNw+AdHL4XHh9YyH7WVmPs7Nl7yKVVWJ4YD/nBHotqrc7+yNRKF9UlSD2SbY9nSJ5e/11JaUv
OCijyHN49yEbgUl0kSwfjx21jfhjhL1po0qNx9knNMP/h6BIGd4AwuN3ZhMy4quYCLGgFTL3nRCa
unrr04ra/rk/RjL2A+/MXlf5MBV/XTyzCog+F2dlHCHqoJhMUOKklfutim+pWTGqEzK2ILJOZn9z
9T5xhasNHdlXvHCAiDNaiNHniI92mStUkbBxvYY3iMNwqjzniTCfeCnUoP/smQEj2qAnihys88nS
mByY8woo1JaW6AT0WnPX1OUz8upgjTQEipdBLdndxmQkmQ3v/t21xJC0QWsv1b6nzl+EMQdx7JIh
okcBcfdEeN9BXfB7r6kB9VU/eXa1xwKc062xcZgc0XxHGEVjWuxCZriUHbPberk3PODv0SfTD9qQ
BEWwv71fw0n5XRu5pfp0XAGfBtMoir9ff0gZRGA50CRVyVYCHuF6zyuO3/5F7O6NhrNLLc+whXv6
tlI1J7DLUfrUd1IdJvV6QBm8B+KDaT0QlZ2mg1QTx1obRN4Y76inD+SL5QpvBb5/giV0SfB+QbeW
icImwaKgegVOOYyUhJb27VyqJ7VXSF24KDRNKzejcwAJYQWKUbmgVKlZS3wt1IKl5X3wCTsBtQMN
0pM5mOJ7uNpuPnYUX0vMRKBTtvh/T9aojYQEYL9Ehx8VV+ow57p1QdcLrFrnz6S006+cfumjV/vv
xXJ5hhHMZiRYhSrhzroh0W6U92YufEZ2QdoT3t2xhnvEmfwXp16HfuoEUs8r7O0avO48pO0igIZK
H0xekVh/DCEHp+6jXnPGlggsQt1c4detL0Ixt8qEXpb1N4dPdHXJcSZpUoKZxV3KWrRZTX5nJFxw
gH0uhFXovastWu6O1BB9cWNaZyciz/3d8LzfpRhDSnpLi0hRmUSOcn7RFKhGvwQSGvuLz27xAG4x
op3vSws2LJtETytWAqhncoJ6uSdKezBPERGVVT50A9a1CzT5xWpfSamFVTz/YIBLGGfxm7rRDn0d
tVeoTpAMxxrGz5s5pBpQ8JEABfYYZD6RJR8MrFT9LpOivvTV1nssQjPrF31ekib+T35A6w5OErPj
4U1trbRZbz1kvdC6RJXlA5IA4EhfpxtcdoFh5aKsk7HxuzUz6o90xhW+zGs7PvYPYYlWvgR+J8D2
NeIsUubIIlonTZDR1GJ9BjGc6fEBRmW8VIGBrt36rnHG1mJJcpIpg53c27J0pk72hf9pxiTdbCys
vzlen+lqbNBIB0YE45cCYdGqqY/nTODfAMMbVR4k+Oq7kRlJJfv4Rche5ZYgoCIktbfFrrzG23tl
8hPwO5gvNCXYeJvP9IPWtLGY5YpQVO+Kx20M9/Xc/sKZC7ZRscuC8RU9r/iPH2XQiNYwZjc3gwjf
eiorLwOkWRNxt5aYogfrH9w4Swlr5+dBhnZOo7wlqIVwzVU+MrxfcYop9NemNyoTD58+t2sFflB4
wHA7DLJpq+m3y1JAmE4Cd8ThZs/sL+DXKpkjhgqw+Bs2AEbqOjXEZ3R+NjTbyB4/6Yj1q4JdxSdy
fGK8XpdtDOPg5CKjzNs29gvpBYTWZp0K3MZzwEhZTFjlYW+GHe4Lr/IZdvRKcDRaNWxvQb3K1CsE
bOlK8i92gFisoky5B4pO/t/Ayb8ggmfNduXbuLFMHaYF8C9ovBPWXRP/wTEwsEFc9zHLpt8GmF8Q
oELfH/FjnZS38JYcf/wB04tyP5ulZdz0yfQgWZvgPubLNhQP7mxHSGCi9aQDwUT8AS09n2C+rrXt
wJVeaethQqordb+HgiWwUnvDWF7xAMS2WxNlntVgb+QzvaGgpEtlH6VRB1/wvA/gciiQObpR9L+S
oXrQ5mRp596NE7XakYzw4+ZI5dMryU7wg1bKQgW9JndGPWjoxzlqlX5OfI/9u8v5XT7j35Bmbbk1
ljNdOFaLbd8P6EqFWfGcN5wyWxKuMlJKO+FUR1fxjtBO/BpY/mEvwhvz1kMbvnEWcVxx2AQciezy
mSHNDrOFUTnoiV0KWCpOoiT6xyIPnvPvSiuJlKvbc60+TkVrFMk2K4qWVyGFtdFjvvfXmtSFT26R
WJ7WQlZyy950F3kwsgZa3ObeWTM6Gdc4poorQ+C8y0TlyEJysYnIehxSsJ9wCD8U3v/B5HTz0/dj
u7JAyJslTfT5wlpqyCNklntjvonTZHlf3LI0nFueX8u+UK2BTsaANrLLSFor0xwAkM7aBSOayRlI
3aXI8CL3JbJSfaWkn4TTLggoglSe1LcwUCyFfxNM+sMuSqDvFY94Ua4uCURW7PMt9vTm30pI+XbT
227GF94nYXmanJAaMNpyy9VntwkPuf/ObRAal1Ycj7v8nME4j4j/N/v+AX6EHHrVj+cxgeTkYHgt
ACRt8dIiW3IZ1YcyEXRV/9rnjF7QFdCpc7VtWpaayD+9tKjQT2kMfo9CKJH59m5mN9BFYSWNttrH
Pvf9wagjy9gcuTlOlc+8r3927Prnu4u4WS3YmH5eSxWTtWWxU8J1kQpbCsseVbXkLzkRFQrPb+aI
7S+SI/hz2q6f6ZD8JHixPld/1Gmh6izB+I83vW8Yen0nB/KUnciMYwlIOCHi9SG5IenrwW/16khS
i4cnYWzqZF+S54NY9ICjbs457gklKgzgJS6w4p3m+dJ1FWWpYSp/cMiGN7I/cyo3ZxOjzZtyrmTS
+gWeOKGgHGEU3B9k+xpt6xEo3uo9ve8Jr08yy1dXA2gi2iZqmGydGSGmhxwKafT1m2UCC4xDl2lT
4MUkp1GbdBReN+ScZQQzGhlB8qNUxetQsnzECR7eGw0BByA/Ceqz+3R0e3WrlB/VLQSp1ynh3KAW
TncU3ypWO0q1HM4x2gZyI2f1XkmGPFCH2EYO97lr4Hy47NI5cX8eqc+PSVQ4rQQsSaUro7GtPx/e
gILFGqLcuIIkukybhwZeN7zWJzsj5iulOxNj1UGgmWgSFiwNsXfXXvgKVX8OpxDapqucfcAnyo1e
x3y5yCVoLf5HBUM707xTJYAoTottVGgmlvl6YoDYAqZ+Efv4WN+lmF3Bm73s/4tnuAWsmQuHTP7I
hZgivRU+tg6AV+tBtlwSEOoZ85ASf2j7rnHlD4n9674WAYm2fzbNZwD7NFW75X10T7PxRMs/wBs4
ZaJ0yZH1LliDFxvb7aZIRdmUAitfJ7QaGjpsx0FlkEPswrbf3sfzkjb0l9iBEO2e8B59brUK0mBx
Ft2NpVPQcZq4yVcU5oU1sK0dsjwztnqXLAx0CjZ4DhWZsr1+C+t+edjOiN9ta2hRgRdutAOV8BZp
4WzO1FV2Fkfab5v8iIevwsTA+DIJDo7jkcqnY4F+Do05NMmfvEC0RG1CaaXP0sWXHqRRVVI/XsXN
kohKFTIS5fCYz24PzGgGl/80L1qYwQudQ3qzuRtS9MvT5aHVdBtm37Qd77Az0MZ8VmAKsDZik280
fX7zjVh9oMcWcwqDlp+cAb4Rd6FoIAMNtJEuOaFhMv3ZhAA5aZ0szaAzAnzcug6L2o2ZgY4iKbWS
BJELxYq8jscBOog2DnDDhDTl/czky8W8N9f09a0r42DkXS0Hsh6c3tUMvkx3epBF4yqhzFjP2fHL
0aGtuvvXq8FQMQId+8rhmBfMQjls91G4IKf0WWeGslQ73D0kr/amUHtG4ZSSwZCQbZ4wRUQm0pCD
XPhetgNuHnGH1nNTz2NCu9G583y+CCU6KyywZ6fjpXeucCahngmK5fodPOHqFABN8IbwUKLuOXpY
+HHakIlmROcfVUmUAjrhrxTZg6qZKrAGUuwKhu8g/FyfAITrWR6kqMAbz8bZP6Zf0uJSGF77+fWs
E+t0QE6eMtevkIzuGLS5eRZS71Tn9+kknYyRvfb8WmPEA1S6mSRXT3NuzGKeV3uvCLOf0jxFp6zq
R1B0OKaveAZ1ticXU29PhOK1KW/BRulPIrniR0nG//dFqclvW5+rGsm3WV8EGiBesmkMtA3dPFYq
bvJyv3NnRXPBfRL3xfv3H6S56Zu67d9/K3yasLUzKHiKA/s4ky1GYE1YSQziBbxUfLrSK1lSY+KT
AMtrUGQgO4NXZqLzoFTUxK0EQ5JvsOjWlIMTBZvvLf1oAcj5xN1H96be1dmCmy4KJAdgj5nqVqxa
MU/WtB5gv1g/NZ6dvKbCGMDHVIiANeXPsKeyy62Ue7WE7N5mwwXje6E5S7znElewSKqEtAuG0UVm
mskkokR36zjJaLTxQ1MM8IYV8IqGNhX4zR/LmFW4HvOzvO5i3qq6n4kP+uE9ncvFtc7O+nYNsqoE
7nsVomC+GfB1LnFSppAXSk2uKo+T8c916ao5HTmQ8KgSahDjsxvIdO/TJr1k6RbiozFSOJHgTXEe
94FzzdXQ320q8OQyzRg7I5I+Az9no+PTsB41PZ6XuDigmjEss+v5YBq6OE7aQ3pnZQdm6kIF4b5W
B5jbhMIxkWoy0KQ2TfOTIAV7e4rcxte2u4hUzQ+1+yxHK/QyZVmT0HvoxucQTAym2f1uX5ASmX+u
YxbBlmNVo0jQ9lXDE58yqegiznwOajAwMNpaZ2BbK41nYNmOIJo5TrnZRtZW5x+p1v4z0dDnIw8j
25Qutw9hNnVYFdmDh0AivQCR85A2PCyplpnjM57TmMyzc7tkHgKsDd0VRoZMIqp5AnDu4OJiHW3u
aW9JwKfwM6N1pLREa1pAY7iA6ynRg9umrSgZmbRJ7WDdo2Zw7urjiWPkYl9Lrh+nSzonfVEf28sf
lGNYf2J7ukKuzKTYT/KgQO/YJ45aujOZyrRZyiWrdHIl/5FtKQQ3aPNVCDXjG/4Z2XvMvmZVKT1M
JFG7sRpMFj1kqhNwfFZ56ToQyHaywfeCXEOuyemS149vhXWHVbQhoER1mOKIO20nokJBG3KPfJP3
w3z1Hdahz11dfog8GaDTDMyOmop0P9p11PFJVn20mxBKyxLFjudkISE7xXLgalXRCrbhcQ+NYFap
i2Z4MhyYJdydNwq7S2WitQxe1kmyR0z6m7ahrJWRxTm1AUi7/IB2QHRKNBWqtEjMlS817kMW8Zy6
rr8MLA3IzAUCXZN5CE45WdiSmf2xWLgfN1I07FuIu+ub2ZT0zXiKqRSp3ug6K3tq+UXAQ9A00JsJ
K12fP/Z6vno6uTsf65yHuUHooeQ0daiLwcUV5ZJZqssiUeX5jZFQvobOdALj8byG/Z/nMrI6JdFf
mNbOXyAAVpDH9VpPi6x1ZVkdFZhVnt5EWYBB25D92QDZBI+BtePqnTkmmHOVyyAxiSPy9B/r+sCM
tQ323IdQmh3CJzYgOL0ba7SkctKCq11a6x3eiG7vZ+o0OXMliMPSzau+Z5pb6TTPKCDjIlmyIsz1
vZJvHSQLQ/9rPkzdH7720ugS8o55AW65EYS418FFWN3+FBzuOzZURjjKGQ/oZnVOWrt76ZapMbz/
Z2CZgEyFCDxT2ZQSuyM5pedBB5N6vKyOKaj4AIe8owt1bj9lSmOYsF3tHlvlBDz4iTADkL5lea5U
dRpiH1FVeisSGPllioJudwlSuQEY+38zr17PGfpc+Gl7IeM1voF0B+2+fpUMxrZQeBVQs/YXYTtI
JMOB+FrnNBDupjdHzjwYDMhRqp+1fkW6SGrSj4VXe46EDBX2AYZ9b1Ckk6hz/RhzJZooWSOA6etS
egB+cvg4s5alcGayEqEI+67M/3e19AsiaL90eqgxmdXrxmToapbkV8jFe1n8OkVQ7j6caHiKFBCp
wwKNvVziyPLsZFVl9cUwU/62DcINeE53oCpxrnsg1cMHDv53JGC0Bo4kzMRCfgDEfZslo4/PcQVs
wNz+lueRe7S6gHm5ErrK8z1whk6tokgFOwTTEG/f0VfqbwI8jL1q1xH9PkaC+WRhPSk0V1PKGOs2
Ngp9CW8NRR7/wuf2UUN67r1u5ksoZq6MtK3nPTWYdq9DH543Q9Bw/ReGhcvclQ8/122DBtrzRfPw
tgRWMM/Ng8ihz9oYpUCVJWG/OojYLmmvLXs1sACSRR1EK2SL4uxKjlJl2atnGlNhaRj6CXpiy/6m
/iskZFlFbYggeKgjtOciAdC6HX0d+9d8/L85AnRTuLwhQI7rgct1uqfCrZKsLv/hF7v0fPbVk4wd
Uj9zRgWNHs+tKNi7YkghPN5d5xA+goB5Ei6KYojDk6R9D4Mexsas+YFGfME5nGk57oimFAtoz5g8
bb5ZiZmHN7pe5jhGqaCoovVGLiQX86thaMTcL8AofMq+UY3bZNQBRJH0PApd4TiqUOVT9LXEPXcY
dWRQJRWMxxAk2bKdXJdhSSw4/Pe0JcYKh8XjCJSlU26RUHHo1RWJ/LFt1g2F8jqWE+CXxmblg/4O
rUqwhAYkvo9ndRQl10AkqBZP2gYxqPPabMJysHHzqI1guDDgb5+/VFsaF72JpOoyp5WD2TP1dY7E
9LVYGSUhtOOKsLc5j4BU0zDcUg6srybzW7GrwIYGte0LKeePDXadlZyxYbF4GZVooX59YmFpNG1T
bP6FBuloMoY4U+tDRGkJUdzEplqHgvNmhshgoNh/Gxfoj7+OzUhnfSMuE0Y8HyvPboKl6nq8ULYX
DUUKRqY3iGthcKynP4Oq/hrUa4jKbK7nneE8usiJILysF0wW0VH/ZC6vTQEKVpmcTDrW9VGiRftH
c6WuPK2xZHU5M7ZSZ9SfyC39qf067ziE6IWjElzdm2GMQGQ9ADqkIzJTGP+0hvOsvT4LhOFUR5nD
/pFCSSBImz1jYPBD+qdfXFj8+ly69IYqA6SwUBM2oz6ZxDm5SZQtTLfOzGjqEgHbn3i7V2gzTN5S
+xWDbIJie6zj65fv/eWe5I9TewozfEVXRcCFLM+34QTCymLzVL/pqREBm+5aQV49WFHtTNQnLmub
2b+lbH16eIFuQOjTLOhsoPdhjeDBRTKdbmXZNQ2pryX+PKGkfEvSxWCXXLpnB3D4CvWdJUHIfXGR
0YH16kqHV2NuT39BMvWcrBafDw9O2WLwxOhqqTavSQiItRl0RtfJqbzYQmwqxKpMKm8RnmnHCDB9
iMEYQUBXn0g330BjgRrP85hQqbu8PUMm/i+rtOdXso85dU4BJsIf0HV1Z6RKKgTH7ayErh1LxNwZ
rZliGLccz+LkvU1h9wTWoDLmEE/k8evDMxDy/9RshgDl5IFAaXr59wBy93iaTGE/TX+x9camCzsj
uAcmQsHHE5HPxrj4QvFnL+M5WTbaOz+YbhshkMGcd3NZo4oiz4qvxn5hf+abfmvh9cH99+hoi797
O5DIf1rRVAFGiG8Zsa/6TyqxuAAkmtUUPEgH4rFkMhCUXvRiDrC9ZzlnglXn931Y/JWuXVxBQreq
VA1Pdex1kBIS1g0lCHAygfr84K55OpATSuwrLRgX6jMADV7JFzDzoV4RlUCKL4oVp2ZxtuCt90uO
C7DcRl8BgmXM3geOsDvSYgM+HHLV4QiptqHj9DMxYWOD0SfRY1M4tq9Q3BNh+wXYz6Q4BNxIWsch
KkJxhPtJ5GD2j5Om3c1V8oqbydExNeOXF8Ep/XC4qjQv4Hq8aOLjfqiq+LX7EyvjPJ7VSWkuBM1L
/eujVdLdDeLbJG0cP8wa42xoji0KX6QIL1U1OCz0NvVdm5Rghhf4CE5zsWD6TPIaM3w/Emqj6fLG
no2e0kZOH02jr9VZ2q24fsyC51p1+sbGOl2awHY0ZShHIGidNF1cTluQovNZLMPbey9JswzPvrQv
lyMLn0GWG1XUHFIeXlPgCJ7Gy6pqxG69sl757ObQvfR1YXWl00JyOdPfM9yuHp+PbU1lYzlrj7+b
TcaE9h3mHO4feqHBDG4HN7wbzNIOxd6OB5XJpq1XFXkUv4lMMZKLePA3ng07Bdib99dSctQjb0PF
DR77ZYkSGrDfTHhsgzle7DfgRmf4uoxkq+oLv2nsZk+O6d0sttWPs9hHoZtrgAWaeQthNS2Zu0Nt
8Gvmdz0HYAIjuFn5k/TD5/tjXJDiSasQggYmRRjWCXFBgL8sEHbHvrwIayNSpW9GDFnroHPOVO59
4a6bZ4irrYYe8EnskGPQSyCghBIs5WK4WcD91Mx/Ib1uhTMEPafG97F84syfEpmPjxe93gir2AVi
1LLL2uUPeZFlfgAPLRPgYcNJnRmkFyjudze0E4I6T1suZPwXjMNkJOnyY8F10jZAVhBwJgpOKjp4
NWtr/MGaRedKI0Do+z6Yim0ELUCEE7Fav/4gBiHfZFpQIpt9elxcT28L7Jrs0wKhwPC+iNXQ1+vN
/BgEhMlmN+0qZXihig6yqiiASC7EH+zVsnvZJp5RVO6jyBTiiS+xMCF7svx2ceRiTlubJ/krTMaI
+Z8ucwLJqWQPUtEhe70X9tV7FzZN5k6LOfTpvPCsNapz6+vv2KeuKqFCXNpOO1ngjuCebW87B217
QdOd2nQ/ZZcMbGrGquegVrk1aUan9uGE4Q6NYhwpKgR/BYkIP76+sC+kVSp6ZGuhL6LENUySovIB
GVFzhSAtqDGnMyd5PN+7/OSnGfDGMVpy65up1WV58cYFLrop7FVF9GlaJW9rv9eZ50lw+MmspUts
oI/fGXpVvZcNYKLDdhiATCLkWclruEl7u/dnoOcSVIZvCUhhDgMT04bANI+GUab/Ox+DV0wsu2mb
KKEyZY5tP8/fvyriREhsV5k1NZp1tUG/6YHhlak6Pt7awcdKWbiW4pZTVZIb7MfpVlUSBkhAqJHx
fdzwx5HGDxcMgi0DKTFx0dmQEA3JBmI9pK7ICsyMh3inaUHKJCS5GborHwO5NxafzETXIOllAfXb
3ruXSElThDSvzfOZJQpxBUjyYbBU+ZzIhO5FpzotE5T2G+E0kLKs0AdQyZzQLtbCMc6dMWIVmbS5
MCgRM1zAnspxvAWIqUjC/8GnE5sswy7wUpX+L5/7qBPp3n1AR963GJElrcw/fIriNgYvxYTlgFES
3ZZ5X/5GgnH6jTxUltQTVSIy0iad4ROb99opPXPAXngqXKsiz2b8Bh2Vi1dMKSS+2EE+e5JXA4mM
w+rvvSFpZ1DYm+4oqGDqXGNvVU4V3pzBIBdJRnXrISRPGn3H0ZgbSCfbbhP9pFYutxohIPS9bBL0
GBAjr0o/uRtYOIedbgCoiU8t9lmLLd8GBvFvnLoN8AyUWOOXXiLaoZpEIqSNz6Bd8gISwoBqUMae
txc6wtUGDLentZqrXtuKffKNnpCAQoq/UAsublse+p0EDEGjDSFymuZ9aCpuNEOKgUohrEAwemwu
KXBt2jxy4nBbeR3lquErbetW8rZvDlROYEfgDbNuTa7W5QB0qBEdtiEqS86Y5Ob1YMjD2egDr23a
kslL8niF8Lf7+aVOY3Q9i8DOe1/QJ64296Z023wKql7g+4SKjYP+WwKp23VPDDKpZpz88Bt+k3qF
eLPnJAoitzG6YPY9V7QnR2AxzT4EUZDcxlCyq1r/j/T5PeHdTHITy2NzvTwa+ovphUpflGvsv0ym
iX1LgbjwIpYV05HSGurMbAK1r5d3sAc6gMvEqPQE+0j3K0G3fTZ2Kh+CkBr3VXp1IrczDpOGCeGG
WtRpCpGiPRRE3WlMzRJGfuQxzn4QciiyVB3DeaSb57lwX5LEU+UMK8r/+OKC2/szQMUH7dw2OFC3
0Yp4/tYcKKOYAX6S47yVYbSoNLCjc+0q5SfoWl7yZQ9j8nv1tH9DVArvefnEWBixN+27W01ZF05T
G95UCLsocDqaAmXspZnHHcxhRUlfVhN/0NOSq6OQ10PuzQVZ8VELpgxxJ4zw37mgUx/ZIxxXHis3
ZJA4NVI5F1YTqzcyBXpoqH9IRgAc8QK1nPcuqUUYt6XvOODH1lZJxuFfkWJ4L708+fJYe4q57tcC
3qCiMHwhqfuFrLKwbew4fq+qKsu2JRmBcfwVOHY/XCpq81epzNZO1bykw8Qppfc0XN6/gOcsEpT4
8jd51vYjP3px51q0HtaxrFDc7VW8NYyUPnw9tEtCANR5NkzVK1NkN2nZ5LaDGiH4qbLjcAxqI5XL
jk11du9LRToRjetKkv7lOrIUgdVCr7/LmCMUXR9npDySC5O8cNhmiYC/hD0a7fCsKw+mY5DBfD2w
cj3WPDkf4Xx8a/gNHK00DUHxrmJfkPYTu8I/LPCkNiZOZh90lmYS9sQD2yzRr9ewva5fCQmCLTz/
aaxtMYYzVneW0mo7DmguwDlrNvwnrmOeRiQJfkUu5Oj44z351tK6xawb37J1h/eZGN3OI4zlsW6S
FKspWX/CAQFwUCtLreR/sNxxaBilj+Q7WDreX/ectiUup+IkwsdiCdLvZ5y/oiUeDN0EcSzv+o/9
xjipsE+giO3dBz0rpgYaH+pXeP7chgvt8N0xneLuuwo8VJdJkvIS/XS5AP59g9w6tZJaUx8Gda6O
ae41b8X+0/3zZfdvS87G5WraCqEiX0yL4wp/i7eeRKnVztYnRUWw3VNMLxqQ3g8/T8BmtQ74hTxN
RrhX3aBMvcJrajyDD8S2Zi0yfomb2Bp85/E4+dfIWp70QsAhMRCfoqjwj0rnIJmzOou9DkWYXPvt
5v5+3k+82dxZqSvO/7Uy+a9LNkSfRg8wBjkluzV6sGerwHYIS0GSK+arVtSngBLAGa8UBK9rEl3l
WZ/QoNJ6MeHEn7in5eT4pksew18aNvcc0Yjc0rqjFRGmUKzERxvWPFjKXGaT5Gk6HPG3xAga0OYO
CetTTKe0+KWHQyLsyH4ur/6zfSMvPOPkkqMqYy01W5n4mPh4WP/pw4/xMoDv9dDDUTt1FAsS0HpS
gcjXBeMlNgK13WD3R0H6dMdo9D3c5zdxsXIFwJOwZOwlYNgnFgYCNVasMjQ5g+OhHoHqZlklteCQ
7GzOQXKJq6T7LzMFU4ZafR6LAfAqrmCyTfZp28jhBXCXBDuxL5FUZXeeN24GnXRc0JZ40CVLMSGh
PiM84qd4RKjR7FKDGzySVKbAoDe6AVo/OMoVRM6TkQxT4uj0eyug/TBHauQin6nn/gWz2IladOqs
bnv7AJKz81SGJlEZAUYmNrBFntpM1fq8kNBylrS7PnkqdHcFpjoFzytLFUplu2ymclKJTO+8fy4G
L5PANHd760vWqYHhgLv2t4sigVBI4lNoK4qv45o4LOkoJSr1w1oYDyiIMD3CgufnpyxgLbD8mpYI
RCn68NMlxW9NPJwS5u//uMlHZmPZg3pYCuWNp38mFetvH/M4XgQylY/Erc8W2zSinB5Kz+/1xE+W
LX9e7lMnJh4Lo9wxluKuwLs8MoNIWxANkR8pH8u7v32WK25Qsyd2m+tMXhEFw0IrpmplYLRWf1R5
bFrpwtXlfAeQmkHsd3hvO0Qo0G9AtIofRqJYCedw6PKVwj1ZPc+jLAFTlIPz2yCAX4ZRfMIHdWoX
81eZU47dNG/vEJU5rYe1N5Hbo2JfnJmmnM8NbnLxTI3WUR5/HltdoD3zMCHgJTmMGzOEni/bk218
0fDfGZsX+qUHsoQc5Z1tzvzdq4cGE0EO6+ZIaHLH9oP22XA+7YCMYb5QrztLuHy3wCu6XwHS1H9o
LEQcxmqKe16gI4Rp4z0+Of85yoa3DNbTIALxyHnXDdhX1YP4AXYM4kKetvzYT6cZmdfha3nOiVwk
QImP2YSa+YfIbUwzNPjwwzYg8otx3vOchzXIyGWTaDPCjXnOlliDng2+/1v8+hxcdSZhi3K8F3OY
IZetdy9gFyYKti63cMj+q0ds1tth5RchgpRib/KVns1bavWPBCN/x0YKjVw3zZMybY+78MJahoVA
NIiGtpCbS8J3UdQMjSh1zev4hdSZqYO5zPI9kcJiLQnp84LgAmbLu/5FYvlbWu9ekevXaYf/+0J6
WS7Uf7Nh7wLEWJct1oaxKq0NT8aQXX/JiTP++CtVe1FK1Gy+It2/+GOBPs6BVq3XWhg678G1Ekk2
TFSB3dkRlQVFjugN+dYfGHLE/es3tBFit13oj7iqxwkoZWGWr7RMpQri4OU/igynVt1UKKoUW3kE
ZDTQlECTfTQW8DkPXUyEZY0jV0z2AH/rHVYH//ZekDtklXY1RxVCRv7+0m3rHEXlAtier98Lsqcj
yvFVoSnDLFuBofxkn93wmkL9Ltn4qPCS/T1d1Hfl0FsWFU2y62Fi57ygXVRUIyXRvqKvqThMg+yr
lY3jWnOVnr0OsBWuoWm0A2PebNS5TxoENQuFZME6l6rE9NYOdXdaAX74//beRRb3ucUrpu+nNTWV
DMRfTfjlJKKC897CyswCSIzvdrfDOfB4T5T40TSNXiwkyhCOU74EWoKiR/Z9A1ygObh5ReWJeKC8
fsdbUfylQfrBHtlq3KfrUgMabX7tdIv0Ll86WrbcblGzsKXX0TEfUjydQY6QB/x0cG7mL6GYvb+G
b3YXFWzWn0TS6L3Majz94PojFSW5R10c7Ax61gW+mXcIvIcKcZp/RzmM0MefYzCoyw3LKrMAddrv
LUBKjVjl+yGwouU6ghKKxm2hfJIr6EC5FDtWTa/KA7NhZfvPs8Gil/r79QX6loSUiXKG288KI00W
uajVr2C1N22oQIWwuPbsliBRtYKo+VtVvnwMMDBGlS9bDX3oozEP7QXbLdvH+DpK0qvAKInZWzhw
xvogOe6fIjdXQsAA/pcfFoTgh7WNwUx9yBRvcXS5rxfzAxtI0X1ydOIW2+k1qKdbbgXmXBEdPtII
FqDA+aJC7fbSmDOXeT+p2tzHrNlHXjeywQypE+p3EJsWZsGbGYkjGRDHOmSuWyTSUQgxa03WjFes
l3cUwk9ruV9edJPpQh5WmJ1EX2xfwCy/GiKP0xp8ZyYkcn2evRijomxZ1sU3p3NVQLtLh8eK0Kzz
FtcZSL+QIGUKkwvb2PcJpgvkkcqReBIYvWhPH5fkxaeJzGPQ75r/dOFhv9G1v0XeZU2SGoH0j8d8
XBbnMlvGKFv1547XYqSYzgljrxv8NjmwvCXoffyzBF/cBDwOLxQNGGMMUPMdd+DLayblU4RZt6s4
vkFTQKA8yK33rQ64S34TuNTP+dr1eMEj22z6TEZjSBdFuxVOze7VVjynKgykJ3FQVvg20OxNLPDa
FUbDt2dOLVN3atpIOkDN7407GEi/TgdBwhfAEzJI+aJLIt7f7yBg0Y4hbK9F7QYwtCzZzbToUu2W
SUPBVYfIPzKVSNkxHMWpkntVad78yyPyPBxAFonRlG/1vxPK1aWl5pCsZSHRVjMEz2O7pAD96Sv6
VMqZVEn7n44HYciwLLgIIbh1KnPkfcFfX5HLPSjHNABSYk2LlGlar7Lu3ofoj3Fc+Q4gwU/rUbud
u2nUrvMdfUnYIxbyR2NivhWHY+UqcXbvtHkLty8vzT/lFqkiDC3dqloF8EyNhZDuuxD3pEFCW6fC
nz7bKNOE8qApnbZmuE/vMKwJa1HidEjajiDHhaW41Y+6BWDAGwmYOhltMCUVqMFukxlH+AhZK5C8
odPHRYAVrMCUo9aFRGb1JwtvYIgs2YzjjKEPTx8w5d6cVVMskZEhmkDfNom4eh8LYEpUFOma0wzf
mBSk6MN/27eqPtKFX0zcdqG1rUFEc3LxBpggX7FxOAtiFx5jZJDaggZI6lsCdRnENJSpYMH7G6yh
vu29nD1NlIPsxSBjT5Blxa6EagLZB4qN9YxLpbI0gVcHsBle09dsBmCYYZSdK3NywMSZ+1qXc8YG
luEjxTBL0Y6hPE/oPLCRFtQcnB21N3/244N7T0fiihTw+4rA6ZPE/zlxHjtdV2uc9UKtxclokYeL
EEZsEGaLNkXsvZDyDbWjzmgQ8EExiESTc0b1YWP+o9ydNlJbbWaGkjSaszGIw2DsTsw9K4p3i0+x
CerRaX/I6qwfFI4jF52Tg6wpO0T7EyEy9QTB0FYFJ9SOd1/rqVrACbFpVpoiDb42oBwUKOHHoiLs
fUBuxkdW+k612P8RXupFnu7ErRuiZdRVxKGFkMQzfk6sFX7IB4Rubkxwf4IwrbZcNzW+TB4DADPv
eY3kfVJhLsY6hFwJ/QGIxR+Fn00fJOqJ3VL/+AEg+wo8EqzyPnuYUhG5O6KdoMXmccn+Wc/UdxzH
grds++oJvc/bowXHwQjf5dmpa7Mc+vD5ReRj1zdvC7oa6FXXMJpLa+tFDB73i/bSn3ZoRqYkXGAC
QFUX2mDlwDaqfuT/7uKOx+lwyoxZAJ05xw8RQv8bSncrvh/UMdujjNSGQkfxskUm4viaMJ6QU95F
iIBppFVe1izPzzOxAh/fuEUYQQehd5NfZd/F29jcheU5mFYCrBfIUSkLB/KhwqrM2pzrh2FSddp/
ufl4aNpv8L9ikIpAO0UxLDmko45yIRClLuVD/1Gv7UxbgHoeEGLbWM4/Q+iWwBM7qqEuYvU+nlg2
5ODRofudq3aewlXlXvA/bMADA3Qn4Ay1UFLEdopr6fBAc+Rx0prHpX7rF4FZZg6mZ1+laAVzxrea
A6np2n7vYLh769WkGK9s259O2WOJ/11oJPAz9A1BVQgcE9bcOnymD7fRIGWDTUpBOW9LAABbiuCr
07PCRvaZ5UVXeMsQ9dzrgTa3ZDIoQMRxPy9Gua1Gy61fDNpSj3G6gAd3/TWuRaDWQ/k94BPSGUKz
BElwXoHcFaULntMRNsI+Uuk+sJGF0ixA8N1Hxvr5pHeHx6O7I3AXjvo7Zq+o7UhMxqgUB6xT+/sY
0fh3HF/xHj0CqSbD/p7mb5Fs8uqqa2y44irLJY/50V90jFmxiGlTmVTiyGkcYQAPM8bxRAunKT0/
Wc+OwjJZHkYtnMoUAXNqS1cMAuejr5oiGN9X7xfMCdts/syXlcj4t4feKjjwFQ6ZlMvilBYUXnD7
nJykPxyzZQl1nw3l4zfNJe3RWEF4TF4cmFVD2MhIyoKO1I4DcbYGOUgjcFl3VWeVSJ/muxmEItTQ
HHo/EkAnIGzPOGMyyttTVEyOGcxcpNxAmITxAiUaaxGriadBB9yccDmGLVNK3FfrzWPZSEce2hlT
NJSHmkFeHcteC6/4tsx1u3xjwVV/JGGzcmKMNmvuoUOgsxn46AJ0+WBBJPfYUt/JfWFxKMf0YXgn
jPh+ZhFit/IN9ETTDTV2nsCm0p/w0WEhSMqtBD65jfypOC7iQ00d5HzqaSBPqExasIRMthfANmPH
2j61BGUEdRjwk1SH1Ou0ZbxBensSd4um7d6PMaILr0jI4YMtleyQO9IlGkSAu845i01Gou6bl5Sx
rhYHuzethHKseAmXh7lowW0S43C6xWzuPKdmDyAnpO/cnCsHmGt5ZUMmctaNfTP9N/qszZVGsdU4
lE0tRnW9shiIVeKU87y2FL4hZfNP4o3RpDdgqoeNOUa+/MhHk/mmovZDa8up8w7lMmGNGg5JgU11
TJtB1P/QcoZG2lSXlIfFsiVwxzSmKnP0bqeJIoa/GlYti74t69S9g2iCaaoa7nfJ+ptFyGzX8NVY
bIJn45iGwE0YlWtIYLlTaz5CPwXESTUDkuJaG3YEaw1UD4niTzprujosf2+Ke8WqLrBT/ykOtjmQ
F9HBKgrwnW+YAbcCmdzoFKLXUqtKgeJTrWIFUfc92APSHjXm6Jm9tWoCNaNM2EYOvB1++2k2zMp5
DRdAkorB5KZ+BBUUG/sWHec5UmhnyQBncxqgenjX/U0ByCNqbROtv5fI/07PZqOGjPDLLtWd2uD6
RrN7BvqH6JDDhfAk/a0VQIdxaTeLTOTEJ6I3+NbgTohN1IB6772RLISGfJHGroYzoYgZNGO1jiWV
NADXxXjFCQtYUI5NkS9NIWzy4l9GbKw6RAM8mQ4rU4/0ZHhjPcTeiuOF8bFy5fzjrv9E4G46C723
PE8n8Pbk6ceWyDoxfvt22bzluh564MwnDc7rsnH1wTS8IE9KJoNX3JQdD4EWYEDaOnB9uJSoltD0
DQTU3Up/ZPR7NBQSAOX5bap8gsNyj3DoAj/MhxV7sJdCuCqkMCpDlFGucsMwvD6Djtmox1ziyZOW
x/7MXCw2Y3NnjU5FiPWzeVZPcJKU0MV4ttu5JFDpHW2C+pnuKvS0fAocEIkDn5ktFwkQpQzJFIh3
z6l4Y1tVodvxrfu3GWqlahwPumBcsqUU/x06pTpr4Ty2NcosO5oMLv5TrFIHNdOUuP+nx62I/YkY
eQIWTARo9WaKlh30gERUQL2J5WuheqA2FoiWfZepTVaVJFOA+jQ24s3tFqDmrS3nsgL5/LXVytu2
KyK9zamkt7jFZoKnyll1oW0zF5trxb3cBg33yT0xuf7spY0L+GswYNlRwndr9Dya+MuyZEthDGzk
+U1NP2k3aFiriWxVeuFmSZz/JWRhKa2fpzWTTBg8O+p5kh2sZZZ/qgt8UnMoMEzl4XjnYp8WTLbJ
AjLOENcelxDtA92v4YF+6nIbNjpAFUchdQH7rt9xVTdT/TdhL0XusyhjLz8aidA4Dhfvmys5oQm9
QvJY8skfvl5XHVRu8y+QQqDRIyvCi394FTWtBrFIfXc90Nz0Xb21a42qPS+sr4iuNFJXa6KL5F3n
mSYqxwwfi/TnHXEiJ/WfdpNFy9X6YD0nVolDBe65hkwb6sEuAUIQur7X791n4jU/ggSO0PniyaT5
rVgUkZukIBhUywihns6Rfte++O75PZSy//ryYu+6cMwTeCtVrnW2u77BgsZNvMBcG5spaI53BB95
T/swDMUbWRQMhGiYUJdwg2YCi7sMPGKSgjjbNdo6XPSryLX/tlH9V3FR8nGhsZdlqGhKODRjcdxM
y8BMCoMWXFnYgWyXC1RHOFpGK4gH7lEkX/YIgDrG/ZwGy+yTbOPDeijOkN6mpFWT5SIxHWdgb17H
BS/2FyS6SSPsWPc0ec3wyyf5+Ha5H7BisVS4lQEz8m1a3Bi2Y+qCVNId/YPQaAVAiFhwhs5Hdxlo
iFN8i40W2eGf9cMnch4oStga02a9815U/feYzN/tiDgY2A+QExVt+TBhWctXWeyixFJ90/qwA/eD
04LpVvAPJ1INYRFAqoNOr9Te8WhK9hDRrxBS8sJg7tjG0m5XydNu1gMXOIj15HKopNma7YiKudyh
Iq2sQQ9GwxJCHJ5UWlbg/2SfL4OpsnmA3s3LIddQ/Z2SUzAKnWZTiJszS4kMPw9TIgG+bXzGGGGU
Jhh076j8aSY8fIxyX7Kn5YsTZBCDyY093fslv/pKi9gCXu7ckR7lAq+AztnRSUsLUWoClzlWVuMI
WQLHIFMXwSauB4iefhUS6JizReetVXWxZNw0kh1L5CaWJ7X5oUkI3o1EqPHCWro9zA2LhY5vNgkI
5HW9+cNOAZf4Iu/2nezX/VNJb3WALDixoeOMa8rxV2I0NpcFhX3qvaIbKREZuHhPb1QDgVxwd9v+
blwIp62ZI/K3lA1xVgUkHAe5iwdaSV7W2LnGnq+iF0sAt6wPaisMmviWNJCl2v4vMbm00vx5SiXp
FcJGT4dzAljhTnY9zCR0k89Pcx+W+YvdBCMZUfmDJPQnAYFB4wVTeAdZL18KdanhKk2E7IhvwuMT
/4F+Xkm04DwF5Qhi7IeEi6lwvsGq7hA1KaqMM6sr0snwHGo3OM5qJROi2sDnfGwMuAJBL9enodTP
G7nd/fP4EwiOUBAimRDgC3vqRMBWFBn78PP9aHc4ZAIyuz/S7hlYhMtdOFy8zOjofLD1XLXMUlqJ
j2laVhR7BebkrmP9FDuytSKdugZZF0bpvfR0dNOP+IYxtKJrRpsfHUIYfHs7IL+r5pqd+OIkVwbN
o+qPBVupu9bAp4EeafGc5GvF8s1nSQlM4OlC11ePASXkkZO2Ixos6QU/CR3Ks+wvnVhMxmXIKVg3
bQjdcHASUFAMEtgJf3zCZJuKoPF91CUxOtee1QGSHkrTiIW627Lb/7tzzIvLMAJGHCocO1xHZvRl
z+0A7DAre/698hMEUb6wVI0gUhuQpjg9tXbGc5aCrdLJHdFrPjJDml9fIeB02Ja+OVm4eg7m5rJL
Bw8xuwEc0gD5pXzZy9ampKDBJns+nX9FM+6oNSBifdEL3Fn3aDLxL2HSbyEvIHnXsZrraU8GcZ6G
EJ+sn0k+RdG2DAxA1dN/Mr6Yt/HGV866JAe8G3tS+e+K18gu8Gs7dcyE4i/GAW1rf7ua1/gjmPXJ
BVHmVshHpD2KbxeZX6psShrJqBNRTagZGR/PSF4qWrd5X6JPMzq/DazwPsF3qGZOrGDwPfiHpHnK
Wkh38C//S/68I2YrqEfA8OpjOxX+QkZiAV4BwdrwgAShlvj3/Oe/mcs11G8VbRmAaeBmXWu1swR9
7xj4TFQR2w0xWoZavWQIpCuOeB13m2qtDZW3b7pprlOGdrQcCnHwsUv6K8QBNssRxlCKqzPl19RS
xroD5XokkVtz+TkrNem7r/0GDuyqJ6lwU03jxCKGzQUr++AZ//V1pLu1bXMpvIi7okCz45eAtej+
5WhVRTGlxbape2T2WP6REb9XSUw2VSgxHoXWKaG+6lZI3DRmGbvS7FUY3+9ytUuZ5I8Cwzi4YVy9
kaxu1+HlrzSGJJHj+qxhnm6zLu1rfW0ATQCZ3xeRYIEAgG4iMctf71JayN8URfqdRDDsnd2BxHkb
pFyMsqfbgxNLGTPD2qSt0c7Vr6tRvhRs1bX4pcBkXP1KxuSZROxyYzzM4jDjf3kuX9EvU6SAD3ao
UXfY3nX6m1ee2OtKsJydFJlbpjNXD2pN/ykbou8pLaFNJjCzL3t7vBMlcBjQR2I1Mn1oGT+5beRv
ivaYbVtAM5CNdmy7p8yKa0+Qt+IW5vm5w+1q6JnhD8FfNAqz5N2ID48ikbT66xgQFrLVlH7FCOPc
yObcx/YUmGIAZzYVcQjrb8SJPKPCzbGlQRnNo90lNf4KWpFApcuYvqNRV9o4cK1pkLVUJki6F1FL
iohP0AEwxfs62UyE2VRDxsNi/Lpx4HcN3j4Sv9b1n4zM7j6V+rL3Lxe8n0NpZVzBzde5+9RPDOou
RWiGVUdpdVBIPrJ2RhQHlXqFqXlPslW3nsijVGKn4L59e/VdL/JVbf53pwm8Hv6pAFfydGsKjzTS
89556wBK4fcIgChDhlE82xZauVHl1VZTkSyihcqyTEwWqd/ZR6bce0hEanVgnw0H0NTpNM+/AJAU
I5J1GGR8vEv5GH+WIJsu/i4e1flTdycAlfhMqLEJ9GAO/SvVUMfMGtP8nBsgW5W0/mZOIRvWVzNS
oeYgEQ5RMseLSAf/ammv9+AdQs/2yXcNKhao5BT31hq2R8nTW96YDu9TmkaLDNwZC01xj3/KGVAm
MioGiRHWNfNAuDjrRstN/mRpIGxMk4nRj9ZhgDFnjGQMYey+5rk8kkdWgcvsjKFqkPh2Vp8IlIed
uDE1NI49uZLFPF9xwrHdeEnu8MWlUdmE7rg9XZQuv2rJtpUjoGuOR0MyokSR8mnuCLz8esHdBYgj
IBCaNZiz1+/D6+UmJ87+HZc1pn7f3EUiZ3ONwMRUNYhoU1A265jYB+aC6K+pmXZuL7E9wz1+sk9Z
iN/VaHbnQzSEFWaBuxQeTmRqoWPu+tO5gJpNwTkT28bC9aSZu8aiyQ4OjtqZ2H7QVGitR1l98cyt
Qqn2HlhUzc47mes6RuqtoKAvM7QmdUSuhAJOnUpJldNQOrxymKIbigZz+iGzeT6OHYGIswa0m4Sx
RYEwpCzKm2j2Zvo+tGpyhJKReRJKQUKzaSUO/afviBxh+XIATuTFHSS2Ezi/LJ+KJ/AQ4C+kPVV1
QfjZYsLJf4b8p8Ro/3FmKCo7GV0CY7LuepNO+HNuCQL8wqAcZAKI1Z3TwQ1F3hFg7oSCsBVSzV1l
uNJz4e/IepRvnRwmoFcCMcq3Xh9WBq0KqbKK6K17K9YqqQhUf8k/CJxTj3ROYG5OOr+Xfnziz1UY
f+DqgeA9KjFIpa9rhW32XALlIaubifXlFgxU6nkCtt9LlVDiGdMEQfbWV6Fef6qASY0JkHEupxEl
JH9NnlU8JOnaKZb0pQAnsk7884R4HdreBtAkFiqzpC4SGJ6IPHoms5u6tZryAlDr18NfyErQEPxk
4NQEFwvn59gOEuOWsZJBrLU2AdQknX9y9T4gj/9YJzNnR4T4kdmjsVoEA5567jpnPUdg4tjEKcjI
gkkH4GK2VEw8YXmUpYZB97JyUrhjZQJOmn/7ccKL7CJLt9oO0rbDI0XnRw4rUJxn0iXO+N4G8v26
PFZHqwBRgChVolRzEGkSpoRB3sJfpGQiuYtwx6EXahBb/FWGfGm+w55WPwTwO8UpOuIJyrTOJ05S
KTCCdNV/c3Cl7U7Z8o6zxngQpMMfrkwDDcUhbDK4Uarwn7SwmiYE4WrRk1UWBmzDzc1nbp7scGoG
qqbI8wVnL4DMpqvRBd4qvaLBoG9rNzpTzPa4FfdgEUNSEdnuiGbwh+GhX6Iquk9mNrSfRtzKQiRr
3G/JD1HkHFA80h9zSl8D1KhFcqexQqUhX9WY08EldKWwUIRBzjgluelRG3QHUSI4Nk3M/Agsx2UI
DfQTdz/m61BIgulxocv9oHYUGnpjT29lu6FnYFn7zL6L32dlFGB80xHUs2J1Zi+2JpobVziiWQAa
IFCqUsuKFDfDrp7hBZ/bg96AvGtB/USM8DzqO2vIzaocuLoXbzmIQGjlcu4bRmFJOaI2vBuqNia/
wGKzBBL228Uj26+kExMK9tc00UKli2KSnYLVITIzT1HmorZkM3LYqk7fLneQr3E9KVsENFLSSoH3
zJDktvw9p/l6EyS284Wx9lW9QHTa6fVD+fsjD/Zxhkdbgr86/z23Kk6hHGPUpkzXgBmxsVkhFl74
t5+OK+3wgq9Fsb+NsSFaWwxYzF8URHcePuM5qQxzL1DGM/VpL3SCPHQzqwfhlJ2hyG9jwynkzNhX
6tF6nZ5fI+x1BbVOUsgaqX88xzoErmPhWHnMxLOdAujPr7DcWw45qqNRIoM97YoOAuEhazjv5ktE
wIzKeko+0yDtyNBPtZqk8RCMTntxWbBKXELyM+7gJLqpSZcEZAjG/WCT11bx1DWA0LXbnltX8vJy
e5uaFmSV5nAztQ3KxwrO8nYcrHlHYRGWTZ9O5VSoMx4dvgTrM4tz6cmWb935JNrG9K67W5prWzTK
uNtqo8VmmsfvJLnVmcYDZMokV+aOx8l51Eg8FdXZwJoclNZTf/mOIe93VOaAh4HPak7s3/q9aZPU
tQJm3gWlIpsMFw6P7vEq7ZbTxdffmMyKFjBNE1rt9l/oXXy1lcNrfZG4Iq0JjfHyEtqEyuRk8704
0OJTQHR8FNT0BBCVWgAOGdQZ6QqwE+s4OEF+UoOEaYjvWcwSer1R6WYFjyck86TK6j2MJH8qymUi
yPes6W4OJkxX/7dzK2E8ZtXpESo5MkSskhxkZcquBzf8bKXtbH/ij/lQexoMjOkTcWZZAm26mf/F
84JZYruMjSTbjgPQJEdw5LjizW1VCGqDxJ1FxyfxtDEQaesfvQfwvGJG2dguiFTn3JpYukl5tVkD
x5Ofk6riLeAVncQaQkcEJpA2vpPQ7IdjR7C4yj0B2nTP2Qb/IuvnfZt2AhQ74RJ8Nw0iojBsaHoX
3BxDKzLG4nVXBxHBNacN8c2aS8aFBWxe0gqSnI+86TOF3JG69I5RId1TGufvcqgYGVLR4Uwmt5hn
SdSCQ4eqGGIwXOHqv/oEjdqPZanXvP6xc95EI1xPuJfd32E4ZDZjT6qip73ilhd5fxZ2rgYvp8UE
Ye3ldGxAwyEhLGbFo4LwGYm8uvkeWLpxD9DaIrFyQAxmMZ1I0m9EaRfGcUTKf8DdwVL1NsZL6x2z
JunVhqnS/hdm+tPWe38T/PSmcMEU7gGf2cVMJdw/wKlOjYjEgzHtBcaYlVylcFCtLytiP8iwcgjy
IDznvOgdFImYIYLsz9qpW/tC4Pdj/Qggtrqmz2pRrjZuF1yXvHiLLLH8zQd6WDbWQCVhYK7BQytV
hqApuQHpU02DBhjRpGeLGZ5DIzaF7Lwm6kPpau/IDsuPpkA1B/aJ9Q5Z/ZL57t/Mhm8vFhf/7Y3a
yWKkt0TReC8pqBcaMqAJjpBTTSmNXHjdwb6Tdd4dp0og/7Zeow1uPZvSL+SCdHUEX/irEstxm5Jn
nVFXs7RjkGINTazqi1Qd52Av4htobr/1/M1ASAiDMTepQwezxo+KBiAGu2x2ehmSHGf+YPI13pod
wdLJXUBnKK/YCQI20xJ2nL1wGTkgD6fugzNZuFVTaiPoiMqklKC4CEWUUH76BHjcw8lSPkHpmUmd
G3NG0BntCO6gXxLui9vP/vEcV1ARIsTFkFE/emSTmcmIyreSpPHgILcg4YgcyDAtcVca2uhbR74t
eEEYZUOZhyPSEQy5f38mljAP+AGFGgXWyT+gF8cwr/YGCfhTjBul3b4Z09SFMmZi9wmPRPkbEai/
MopENf4kHkoL8XIrhvNM3bbnKjTCiu+XCGMZdPt0eIKcf+s9kquJOWSVAI6n1/hGatAzm3dH2Fae
Io1DmT+YfYWOP2w8rg61A9n/nU1FQ4mHn7eNy0LossGg3BAOVNhmLng5/Rrc4Rabprr7K3DT68sV
A6YTLZ5gKEtnnBKLcIzj9ZhG8ivk7M+ZWYGEzVFBkaI9PD2gADLjdsbRsVd13zYmw0TskWsf2kDD
+l2pstPSV4r176qwf8YpWs/YdQ78PL+7H9E5uyFd8xX5+DRyIe4tDTuoDn8mFuaTjgqfH+W5apdo
1LTg2oHpHwpuaRhk/9GGgiaa9CmW8DDDxxb7mdWMxQn1IR9+UiZGyKkuxk5QRndfY4AFLFnvLl/a
thilW4XK+lMzmtsSxwxSWfB4ifzpbXSSckeTygiij+3k08DLP7k3LtgnP+hIrLN+a/dPT0jWM7Og
XrveE3u6owb7nBrQdtA8uNNegVjDYX4T2vcJV+PKfrx+qmJ4giT348fmK3ORpPweu3xWXALxhf88
+kUB4LkhsTeJYQJwPx0Irw+WF2JAj6HJCGMkg+EB79ufToUlvAsUJvrYCi0Ma+/rAXY2HC5N/7eG
Y7GAvwi1SOxEhTZq6prBA+haO4cW19N+tU9s/Ov8TLkRLutlrqVGJ4he8EyhJa+sqoBaz94acl7z
q61y0JlCPmDe9rF2viDgHwLlhp/KE9q4XrtMtfycWsWvLkzQCxMTTczXS+ABNb4v0ifEpb6A+Y9T
Y5URfCQHCr/4wNLemC9Q0lsOSnekqH0ynGMFxqGtbEI4K+14gBFdQAkauISEnhkOuhAcaS26eVNn
We5OsEm+1XSIpzeq0USAWez2ytHwHalHncMhmPunWxffSZJIUHkL13tXG8GqdzljZNANWQ7XBuBG
3OVQcIGQfhBlqLYlnrLktNUhva5HweoaxddosbL+nSDBs9JiXzfLaP40W5BBZb89EyU95roHuMIn
K7vN5QiffGCzwEoNYM5SXQ0ZBJ8FET7Flq1b9vvOvNESPk+biELCBXUkJaScDK+M6t68Z1mt8YFG
kdeA9ql5osZn4vSV1YWrmX9aZv4JLpXF2JHxsmPXFYxltBNzMy8mCmT3hoCDCS+rvwR5/avbeAde
rehSykpw+UkKFGDUHTTtHgJ6Zg5OqAz/izDtWAfDx40xMNRCPQ0g61NzYjnsKF0kqbssxSWkCNH/
RPvIQJybztAJmhela3yCYrsVFTNkHCfXifGwA+axqLFzMOzpsFbWtgtGP0IBcrca/sXCv/WVE51b
p9+R90SVSfeijYs9O0OMXD+Wp/NUJQKLjme9QF+AxOBvrVbyXuLbG7W9IRaTwnuu6+thyun81qsg
UfUfD9jWiX5hUjmQj1Y0yYKJ7lxDoWB15LQJ8Hvbh+Ikgq283AztB5CnepXR8NRd63ldJMPBAB1l
IWOvMlxb0IbOcHnoQDesInOQ0RCxRJW1SXFzH0JaI8avfXB8kVxS1oeLE3QKOeTTdCs6gihEtlmr
wBmYGTIm4jWv4Fy0DU58GzqomaFvro4qdUjdYg+OpnhbGLa6OCE9ihFHrhlBtPftpDICO4dCk9gm
gNlUDjJ45YTT4nGN2rLh6ZsZebewHiwRN8I+jbIqz/d4QymPU7z9HksVeKCucf68Q8V4zG59Grmu
nd8JjK0wp/xebwvZ02WK93G+N9R0Vz2moaoOsAYk6uDifUQluS/v2TFPWsubWi/0kLDmDdjV8tDF
ZCHLaHGW6/81Hf+57gQ0EZGyfuEw6CNZ7HVMJ5vooXUWBockQ2NGm8jxa3oaMpLsTGPVXeaDGnXV
GY/kRrf6u2iIz5xq0y86GBGquh4Qa2E+m0yMCYG8svw4YjldS3PbD26MiprwPttbzVxSFuhSduCG
KTmMxXKtQalpGKXLA7Rk5Iak5CU2vbHyvfiZtC63m/66yGceVb44PDMq37WV1lIkwHeKCNP/Jw4l
y4yYkj5CiAh0L61n/Q6c4NeEZLwQT7Lw57uzvMw/2KjJOVMlbPiDJe6yCydTZWG5ybyUtXzDFDZG
2K8Bq8TItmULP5S9v1U0t3UJzWtSNaQsNcTkJBAkdaLDrm+viNjGAVr4oymoE+Zk3bYC7SnoRCvd
bHqdp3wOsAOfr8f0lBuj3/kcRi/AQLYtHswwTQSzLPivOYohllIHt8lOWfy6rvGooAsnIy9+ZoOE
P7WGnbZY1OXE2l1RJ8q9DA6SBUoe+ifpfvoBa53/+5utFS09Xi0hli2p0la5K3757O0aD+dtKkp5
c0Xb/1+slCYodFW39+wT1c6sEUM0YaV5/Ov0Ry1JiMB45ttbOJgR5YlwMghvhTaA73jRpeotznqt
A20UozY/vKVc2MhhykDXgms1sfRvsaRHxmq8SNEAbaYblNO7/UfZSgWkxOdIdKLbCqMDch3nXaF3
Vyd9irllm9RqSK/1eXDGiE2FlLDQQ9wTkPdeYWgwFtyj7MXm40zUlm8ml4yqpLm3Wah4hFHJt1gS
bIKWJlPyi+Q/CTQsvA+Doa0oqmEYSkwgOIt8+AbY2P7rFRCc0sPpYudd8fMMviVJ4SUmtJMx9mL0
+Ltl3uT+9JSfGpwxMaGYPJOZavXhf/TIagmeSZqJUqEgjwY40L6UzUFi/iEY3UzAP2KdMAgo0NtK
RHOi3O26eP/B0zEd3f0YjbT1cVlcOrDhS8CPYEJh2WoIlOERFcKCMPmbxRPyKWL0xxf+sqgeN+od
7hsmZY8Jhm4tzgb6TL1ftOr20lnlvFsAoIODdXuIb9KBGkwXHIx3+c7F1MGm9G0KKE+nE26HEAXU
qwptqYvTL+iAOhsVean1i3+N47JEcKOyWutTCKul2FtJxqcOZNxV1Y/psgyrqHVvIZ+Vqd8QA3gp
D2OZMjR5MYXDXkLlUWx3aoTSY7RR54iwg2gOyRbCHYObEgVlEnOlDt2xPikv1C3LXzl4c84bFYG7
GQ2wFpt7alt8F3KpZuVIOVAG9OwU0lCaiQp7WexNORIlnln8nvOEMl6b4Uq9kjeox245L6RbtD0t
Ae4OAPLrRguQvV696Cb44Ut+YDdO4ZiMWkCVuO6xTU2H8QPh3NbyjmQEiU68A3ZiYgUqtZUnEX7V
UIMaQVgPEDONJP1pdi4A3M6N/EnOWCvImKMnnC/s+RcmX2LMQ3n2N3IBHJbm28NwJI7kphNArEb6
MPDJgnVWeLmWzT+iw8xLSqinrY6itrMS5deqMa2jbAN6fQ5mjBpC4A/OAWdL1Jk07gdKZdJQv3OA
+kIZlE5kYZDdCe1Gf31rEuZ8euptG71Qcp5eZoq4cPyGJs7gB9TvnvJbaQkQc/PvbH5vE8r7X+A5
aTcpND6QfY3gqSjmyliw6oMl5PSVXbWr3EFVAxMWdJReJ3gapUJLDtfTuIJ6FH8w0b/gKECSjEyh
tqzmxJljoQ6ylht3AhQV2yiq6hja5D/tQgD7IteUj9Qj/wmJfAFu/pkrkwqwMAWsSHuwOB1cTN8L
GJctqGGg94m5gG/vhnWMEq2cWxos71sqiIUyW8Tq1Ms9QxxWRY8VhuCVyKoFPgpJPReRsKUFb7mC
QZOrPch/V5WE6i25WqV5qmS/49Idpt2gSF+XWwYcTvv77gTZMNFY+r+aez2RtJk/JsSGy7H+nx3r
zNULnQLKH2DhO4lr33DOCwle+TRQGHP+jxfRZLO3GLYjy8BBgLRMA+5DSmUI2RX8v5jqTaFch+TW
XXSiQHj6o2FsFKvyErRM3XKWss3YvyFfT+kItSWbzP8ayKaKB2AxRvxM+fukGpfdHMw7sAumOSY1
sS/sSzRRIsdXutDKppBFxw2Uay147HSiaY/g8avzynIeBoDW7ZsGh6XXU+o1VygzuBBglnM0BN7w
RmX0ZGv5Acy4M2k/7ee8Ze/nFIDrcxZwp/Il17TEWJLXo74ao5OrZswdshTzqz2lBrv/JKd+7KsG
Ne/BWKI97ThVs4ADdveVeigOK2ZvcNT2gO36rZvv2Q4b3Kgza3F2L1ovbGDSU5e+QdiX7McCagad
DLrHGkuvS2UobHU+u7xfUVu1m9fOSzfgZ6dBS4HrhN6SiyIgL9p5OrrMRDH5RyarYSso1u/8T6Dv
E7JNTuoeSEkBARbvfvUVqmylYAFYvTpjZd0Izad3p6dPRWdYk/qCKPvR5UwrWHch81p99NFXW8K4
MGl1euwF29UZFyEX+l/UQnRDHqTukVHKqzFxn59wD3DHaaYuHNnCtrM4kyP1U2Umn+Mg8t9X1SCs
ezpd/ZhtIHGM+af/BXON09asli/1xWUTh9T/DKxlu0nD+4YBZZ8QhKBuBpMYsAkEX0YgmsrSeovE
YLje2d47BhO6ZdtaOUg0Jjwa6wYojSGzryEpH5H0W0d8kXFz23r0pLMLOjfP0dF3NChaNsaZRw59
kd+hZqFm7YCohkzocsvaxmJiXR9dGhkHw5btFBcpimaPM8RJL/2QGt7kwQ0aaO3cZ3KRmm09Cz79
MbtzxFy3ivRwKJRi8BuzCe5KiM1l1zB3D3QqN5RXaeQbSqgGzcosR9Zn951F8qxXjLReEKN2iAmp
7wmCBNtAQTCton4SOVvFYz7+yvAbGWEgBN0b346VwdAy8EMS+YDHzxysbH4Rczt9WUvBmVDGZqnL
42veKcTe+GNcg2EiMoRsA6euqRglPOBqJfbOtZgbZ2zNK419X7k3Q5W7xZQ+4hEUYxohYTv2SUOH
D/+h5czLwIKmLHgJ9N62QD9vUPvf6ZHNhN5bTLLJZ5ykPzavn9fN45//Cvk0EfjDSwJaVTFjgZOL
zM5MfbBe4A81nITRAflJkonPZd08wy4zZ9ng6Fo0H6VxO/+q1o6xYXRLaXAH8KwnQNNPbbGS3eW1
NdMhk3ZwdzwNL8BfBOzy0EUsQDkasH6uf8BCo1VtyNNpX3am3uainN1Z6RzifRnQbYCunwJj6U4B
/ZX9mFYAWdrg69UwHwmy/RZMvnymgbnboCwTVpjCouyeEgkpbhFi2erugj2rWI+X8EHjnt/9C3rZ
LOLOCSvEaxDksNt2b6FDuN4B4/ecy/BL8tsPaYVYhiuMMZqIYPczvYXINpe0Ve1QwdBM5qLq91Ng
ldZZcZs+TBaPJqFKx5naCiKOkczFuf82I5tzcjzg6vfwizaTa3WmE87CJMTGjJqPTEkKLsvlNTDP
syodxrgFDsNaqct+MnBPGQSNKR3nU/lzQSGbTs+TTjbkeULY418TF6UtQzRQZ7qKxgTAX73vihy2
IQP9eRSTWaHG69XG1FdKCw7QmtXOGWn1zgDnJY3YxYGbV4Vr/JIBm8AA64UXBzrHz2gdqdsAKl+7
XP9p263rygP+CJRxYMKAtbBTorTuCq/J3y085fzocuO5epe84wenM9Rre7elZsJ0fQFYGjBTdZd7
jehuuejkKvfQbcAU+mBD21a5Qw5GD/FeTvaWah0S7kHlMhOyyejaxzt4l9ZJn+wgX7BlWfc/vwWt
TTbuxLukvSab1500G1A7DcF9X9xb8FWnPE+YHPxV7lXZ1jG/0fNDWUmBfxor2r3ljHtu5DF0Xi6J
MU20V2thkwY8np2+tmd6naWXGB2uhvSEiFD9s0xwNaLw9uAOlQv8fYjuGUJ0chnXGoeppTBGwMrv
IA1VDojNBPxV34jOaMeliUYORRFjttqvDdnMQ9sq5opI1XRb4166Cz4R4Lmy4T8NDsnxFuHGneXo
F7mDnTEBbGqgijlgH2oOj6s79H8B8DRwr6EbMpEVABeafC5l8HpPeN7gOnAvet9OZwhXAtZNd9rc
Hhfjalf0j8565HxnSV8y3JJjleWsp0HFmHuR+DDEpDG7zx3+5XXV/JygeB2JVzcX5QPld3aBmUf5
0FK+0/n3ah7KP3lcP7StZ8QbTSfIUvpfn9SVpChaB4D+m1mzRi9E1XjnMPuRdWm2KSJETeY1Z85u
ZopTcGJbTnfCaHOAMEAaarg8qMNyIoYmsO0qH9mr9KaG78jr/ywQbr50URd8zZ2ZL/S8EHder9/8
BwDs0yj02LG/BCwMsT7eAXzS6o+u9bIEbazu9MMdxy1fUlo0X/L1zcprENnClDxopTEryzxrEJzI
SbovWZL1dkgVm6nrqIWjhtFmXc68R+qEOheQKgiUW17+Z/2MRxodc2tCjtJEvA1395cYcS/MEI20
CYtu7Y/6Ik1foGKBOoNzK9k8rtICQJYixkxeyG3tKM4alKUMXeO2sv5bbV4dNvA3NEslqYzoT7lK
KRjvGfzIkLlywcw2Rrt5wNbUjoFY08meNziJZk/oZ/qpl8TG/fiAnEDsG7Zzb0EhsJnnz/sLDc+y
u2BgB/pMJKn2Dqhz6BTdsOZCjeJALhGuQznCf5UZOYezXXz5xTpwXjAB51ndL1tStOYbFTHXEWbc
tWcRdI16r4Xi9HBOoG8S3yAEi2QId4soFKuij4h2Zk1A3LyaNHeGI6KBy1hvAX/0cHEw3BYwtUHV
KAQbZd3x9KG7CJPzmTmKj1PZrDHj3lO3ZCwia5OJT1n6oIm8no7+LzEiFpNmS81WV74dVktEnya7
DEqwHhwTbpShScdeCGNyxBClt+8l4HVdaAkGNJanPlwS/hi+vsyqgzqpZUljv6xg5jVXD5lIQ65s
r9Mau6MpneHvDHb7YnhPUiQN8/FgvUP1lheAutmS8hHwyO9SBaM4miI0u4QNqPRL0wawyl3rWqVB
WUmDUnTygDk4shAaj4gZTdjUavx/15Bi5WyGWSHxQ5ZEIVLqdbacDX/me0wWfUJzYIS1t/E6F2zF
R427pMwIkRZv/zmThcsD2n1Zn3QDO8lttncuuIfQEDGSWleW0gQCSg19EfwgpdbjvXUKfmbhFR0V
A/AJwxfwY1cZM7Na5P/nBst5IaTDPKziHnJtMAAotRzNAPbOOmNBv1vFcHUoH1ryqGcezvwfRSLk
YuUv3qCMYGJgix8QwA2Ow+jwg8KNjHyupWErvm3Yvos+HeSh95beXp0yJbL1S3h4HY0lsEKP6s6z
eI9qjPuoqHeBoqN9Ldpn7CgTTIr21Xr6dgWQ/FFK1b77g+tHo2T33j/oPvr7roo4AVEk347Bk0r5
KCrJY/P746LevaDW/VLcFj3V6x95BlV0wxNuTDJZykT/jPnUFm8U0JEORyrzi7keu466k4PBw1ZY
quDcRwzAQUIFLigczNR8+qhJaGEk5Hfo6Ga0dtDSd8nCmej1aIqhnmBCRp6hsJyOhAbGuHljXI85
OzoKj6RVYBNjexm9mIrc5X5bYHucsj5r8yooA1ZsYUphhIh6hEprJUFFM8rfdiT+0nLMrWB8CHvi
q2Q2FZyWgVij2rNISCzsPd4al+Ntn4oOOl1wUSgiNw7wFbJwzpvSF5f7aKrzhTDDVm13sUi8s2xf
o0n3ynAUGRbRG8W3SJg3AKB5h/8bGuHNLS/rf7OOk3UnGgTcfD5fECu2MGEh8YIzY40pfrUB7lO8
ia/PmnJJSNjqiINph3eMDv9qpbh+MwHV/YMifS2+ogFcnCOGjlNlVtVbCOCsXvWV8jW6O0lErIoD
xgsBc4AGRDw+8Xm69zzzxal+NO0/4f8VYLpFmOwyvwSOk5HU+zZhV311CFKR4znAN8I91zCVNm9Z
KAlCMkbIWgq48gsl7OnZoYo/yJGqBXHoky9/Kd63qMRWWy2P/QWqFI3lO5nAxIa21CcP0HVbbKAY
KiWGDFe4P6BXWiMCu2nOwkpFVCAOi9ho5Fuz1Qq66Cx3bZ4tsSqU8UWajtDAyEKoT05LnI4sscdP
C4enZA6IlFXjDf/HMncTvj8/O3sZfjl43yBsWTXJasnkr9QVlIu/WaA3M815GmMYwlQyGrurAAYl
qiGLV0pFSoxEefgKKurIdOEnNKOT+3QymEcO2zRRga8ysjzSGE8mQwPVqEgamDxveyBQHrWQCRCY
CxvH/WKEScKhCrF7ubHZk5tHBeHWO0rOtPA719ViN0G/6JPW7jlitWglVXBonVQlDDfx5jU1wIxB
BbZ5uFokmvdAtalQP3hzuaLpbSQOhQ9tahg7uJBp+pjFIq8/3oz/BNPN3exAemBKnWMfcSJmKyVR
j/UKRBSM7hZ9ZgzzToAxNzO5hEVMuhVk6qCupuASr3pNdHUTnMi6CkHUNfafqylUHhQCMHSHGilf
lOzcSuIYag2FWJhRIDlNmNJfRa44ydpkLjpjkgCuke5Eagqh43wGlwK6OJhbWEX7itcEsfz74T+7
hQIV3h8qIHeRiCqt5qug/Yfdu5VozdarPgyZdusGWHNTbu5s5LLQaKKRV0xZLetkFHCBYrHMGRs9
maSVGgM3tVFVVh7fg1YI+GltTsfln9cHeMcKz3rYCxF4uXDvxW6U4eznAfo2FiFTOc0Je2SQ4yCm
MfRDa0UlObz18vi1HIbunLHAtfqxNLoHbpQ1juo2TsYmE4MU8hmO7jnda0kqixSZjqmjvDqvJ73w
NWiHBXDnS2wntMwWQA6k1sPVi7da7RW8B55NZvfcgFrjkzq46Y1mC0dxwWNAfaG9KwSW8CSY+mzA
/INZnEM9fc6OIZGOweuyNBiN8LzA5pSkPMa9frI8XKl9+qbYb4tXLtkgloB8qJjT0gugyi2TdQJk
WJOguxFQKHNm5VBR4htMPJ4xZFKmYqSCzPdhcmM6swN4FNYablFJUbHQf1fm6S2rXoqILTIfxjV/
EOX/gJko7AcfaJTm/moR/VcsHnjcK4XL+ZooPFDDAR1Enw74PyI8medGcD/hgxNAuslvOSGhn0ZZ
vqM7Pl8f9oSdfvxwPn5qY0L+ZgE/h98skyeVrrWNHYxl/eHSBxOZLHfBHsdq6J0crXfQIaRvED9R
7BhN0tOOzz5nxFp1ZM5SkrqaDbtXEamOb8P8Lxr7UOwBRBKo4eQQwNd7Fq8k11hj8FpxaE/hfPTJ
DeSGAPobrO46GcYB4O0Kwq/GN05MP1Ty4VIy0FLfCucHdLRhn+0y4uUh3U9atD4VQC00vFVUogfJ
3Y1Bp5/ESt+mRivm39Ap9S8hVuGuvdFijQVHR/PBxo4Zju48oO6WBLjlmlxlTkcQyQSmxYmy+58n
DweFCHAqMmdmU+EaxIQHLo2aUbYtBCskGKIop02cqNtvVB1mtJu+fLXO6XFEcp/Zeme5qzkGQ0ob
ZRhLIyreWU7R9SLhXc+XfxfjUgCUg6Mu5eBeyteNh8+i/5JfVKsi44ypYtyMfG9VCwN8isWYZLlt
M+pHuQWJ4Q3wDcxDuXBEkPwVTw6Bi3LbPaO+iIEINyILXmeyCLlFIJeUHsQRhXL7u0/TwSVvoyzx
0/RedI2NOr1GiVveES/mP0mbMBNx8DI+7SJzzW6DR5e6K9rW96JLQ3yjQFEOS85DUdd8gKMklCEd
I+/zum06NDUQQE1MOCjuFQPpzfKYO3clHzaFoN0xuL4Ow7dcBz1UkOwae8n/QHvq2AcZbpKKgNRc
aCH6o15TngFOFloOA/eYV/1a7Yrp7EeoRrFyc46X/CIiVE1PkMDkyEpHxjemyhFsQwaqfZ1Wr2kQ
ZfInC2RtN3pWmR6WSWEyotRXLB/AhsINm1+pIi8YDvmGoFUhIKcVenur4Ka8jEi3ghvIFMw/NMGV
b1l167TszHpwJdFI7smJDz9ywK8rNu/XpQO985Aa3uticoueHhKnAkrf8iGVdYjPz3rGNxfx72sI
1Qa6mUOBhDyzbtB+SwcClgFHC5daKK34ladHIGxWELrHMISON76/TSvi1q/fuoS4JFSK0i4/ZC/3
pxZYo/9R8YlaH1DcKp15BQNP8UnevpE+n95e3LGCQfwNaar6rrR1sXgwil+ypGSWJwpCUcfQVENb
XB8O79xwpLg8isa6/zrAGiSsR21qI4jdU0b6IfMg9qruoqp9RGctmoYLr6f53wFdbfAL1kw/h2dX
Hhjbg3h+2MmUWDwC7EfQcKHg1BFOPp0SswUVffxvoZbZ2zPWpORyAatzyArh7dsmbkQsfo+nJQ6g
q4HUezjS5y5meAZlUyffw/10yf9rQUflOzISBsCLBYsvb/prZ39+QVlPKfEnfuq7DDAfBX3PsjQ7
8C6uto+ER5iZJ8D+cvKXeBO+ZV7F9uMheGXOfs4+sdMGpWwM94yEy7n4Q6ZJeWoGMsymMMr0RZ3u
ejcbTeKH3akmn+GlXEWjSxivtEX47wgkIdrl7ioGqYnPErhmfvrfPvJyHIOsuWoEjeQ5Jo7TvRtT
PDMP2U1ztd4EtWXrJPdVYJ7+lw8oxD6yfNsxyc4OUYuF+EzrzszKu3MCMlKqGAjcic3/RMhije+e
uVWx2iQsQV4UoIf07SUCowghMAZCf9YA32T6LNXGB9tLmRym/oC4sV+zB2DSKdy4YvM4WIc8UOuf
dklzd0fES85b8CxljTv8jzTiGnlZ4INCShFn4KMSiAHMc6nStjVKk4WTZ2xUgGsLmOFcAbhpgiD4
3hwbRZCV7bnkyzJQ6li6iZYT+y9GExVNTV9crtaFJMKXJaj6nekfkel/D33QL2KgfY8yv32Pbssy
4Q2pNpg3aOMFzb+gga5G8HiLr3TsNaiQR90Bx3pivNfOWhX9pCL73MBDweOHtFtxMyLmjKpc2hgk
m8znqktQrYX7ryBYTi6OSUHTOmqARr6k9ScRI0nZcVRkPRnbTcCRlzJY4XHHVXMqeOHGjeXh82VF
ACot6x9rPbqBuf4W0h4E1EUw0g6OLjiUzrdTp2uYrAiZyq3RyWERibr9DSg9boCOIaYBW6SuWzfl
Dx0CKk6oRSI4j97pxKyl8kFuVyxIZqf9lDlgQFA9wZYaEUnARhg1VrGGYBeCGlQUo5myaSXcf7DE
lqP4PnuHcW1bs2qRhxn9cxlblT5Se3lJPYkaSHKM2SIEUyr4tRYjYL2hxcf/ZoW18eaB0cJjToiT
q+G717Up4j7iPiSrVuYGWJAuHU9+J9k4wOxcsMUpX50txfTL5KOpWuy1D61aNdc4aKpP4SkmV2Yc
OAYn55am1wwlxgTfLrow9qFPQVR36lOOYMB2sMmG4ne/lWqhA5alqbrp5g/rmrMHhXqGI+NwN8pu
N7o6LUA2awUJ53PaQitc7q8PR6lWAksB8aZkGh8qK/AlOY61KwkW0M1ZKHA1CIvt+FF7Yd/XSlc9
kFvZ+qb2O45Pphz1gAOwvZycRz+bld0uez+PQZbVYnnm9t+03U13r5QIgOUkbOb4NHvuTt5grcDe
XuJ0AiYmMG52voxmiKc1KM1jsbUMFdqEaHDYUB00JvWfL54IX9nzXCa/32M44d9pS8obgiAhbyQK
T0MTsV8w1y24r4qJe6wUPRzHgEi7Suo0CQylJYX4t5UItKabhTaMg871IIOjQxPCTmYW4qJNYXTu
LG/Y+VlAdoyFMrtASndFolptb94Ow/5zXh8rSGx+rgW7mVnZaoCGDlSeMO/J+vxKOzkqSIJarnv1
QYF2WKrA0R9dTTaBb8ycy6HMn1Nsk7VW2Xnym+1br1/2jOYGSKIX2s6x9+txBxgt+P8sGlvHnQCZ
v6u8NcXmDjNETIB7yh1UKmdZo6FhNhxBbtCr7E4HxbSOHNG1Wex2tkhCw13gg6s+nVS7iSwlkzSg
WMJgSXaQnTyDK9tm6dR7cv6regvNwfnjI81H5t+sj8qCKjASlt/Mlr9OieXH2091w91CFSRtGULk
dvHPvOwtgLDcAAwfth17wmaDIvbV99wrc04c4OSN3tDDAanwzuuWcluwjXJAuUX3f3sZBMIEozSH
Zzl1ddbn6D0ftVpeBbwA0iddMZstmqPjaZoQ3Eojv2rArkahxw/IVRv0jMJO3ZPFpDxI1o8QcNZJ
o1cPXCdg170qbrLHqANwMk82R5fyzqFlmZoWmoMxI9KwNR2/MV0m805Cb6bctd9u2+wzylw6Db1v
H1S9qB1ypvTFkMpnbawYRqup7JSxatrzYjfIEc9UZCtz2Yr8919K/jEwMWzbaETCrJPPYOuPveOE
IOM0Fm4ghTRpDCkttx9U1q1x35I5bs5jTZBqcE6B37dPCbi2fo96iNOwmYZmwcRUt4d2hnnHmvdD
k8DaiKISgQILgrPlZwCPyCRft3fMxSDP6qshQTGh7afokCRUMrWWsudy9Q4rDs/gdDveSGfg+vDI
Pf1cCkHndyg18bdfcfplcmVCwmDL4uQdu+mqy2Pz763uLCKf/l8t9qsQ9cDeg37sKw83WOxQPqEO
9NtVYjMZh8tf6+y1IyVnBDZIyH1i3HMZhctT2swb4mCNlfD9526SXVI9vR/I6uKjekGH4sXQmJ/A
LQnDL6G6JYPJ2ftPloc6VM0I4yqwlDcORYubJfIOxo31utowh+J0w+AgiNcYERjzLz5GGOdy7Axg
oUojNoILf+nYBwOaI9a2WYcFgF+rV5z2F/06AbkZBZsXmcuFY7i79eU0WX3HoxqwqmVLRl+oa3Rz
U6dffg0VKoBQyGS+v0n45k6UwikMYBz2paTdqB9ItIMPoGjeMJshAGLGZvKXmiUcIXQyDUnP0oYS
NC2s7PLEdZbLPNUeaDcohV96/z+f+ReCkcOfAcSY5BeTwbmzuzhedZcQjLjEFndKVrziX/tnff5u
RwEeVOSzFPVPyH3zSwZjyS3sacJahuEpBfXJvtFZ4ImGtZKS2S+6slub3+QTy4i3SffIvx8SIKJP
+/p83fHPRKqzAslgd46YYMaLju1EVZaDk1VNDrJoLKq6d7seegN/8q5tVsHHY6rPDBLyKZnblKUr
Q/4V08+nGHx718io4iOmw/6/xoq+O6vxpFtsqbV32rGM4HoFzZr3ptDP1aQK+bOgq3pMgsla1oY4
VgggtXEFpWSVm3R5U1gz7CTyAtHEQZ1kRdZXjdVsZkicHa85xnTz0qFDYPLEyG3UOoFqifgyjjQZ
QERAQls+mkQLfwctaekI8a5ABUCZojuQJc9c25k/fwZjS+CqwRNWe1CJSNngwSEVNo7Y9aGzwY5P
wp3Xt1iZCUp3zay6uUIBzY74/ZS6CfPSirtWLYbjQQZ3cZ7eWCbrjHJ0ocQPnDk5NEoxELDcZww6
Ym25X6BKp0qW0C6cPDUbK0LCe82YWwQAXBlqAg1XS1yVsEmFEdPY/E0B8dhaiwq4mzLoLZcmSmul
QBBwXkUOLMsQATzkUAaHUepixpcVm8wXPWGIs6Z6aJej2Cz85VxZBxmSPZpyeF5TAalO9nBScFto
isZjYCHLbThoG7ZDxPYbp7nrJKmhVC0+1mkw1fdCyJCQw106Ukbw8YwCow+u6Y7n8Jo5h8CnkiTm
lD03yHNKlAAB0NgxocxKxVxpQ8gfeUlX1b5F2TvVQl8d4bW+K4JdEn/rp/NkZo8GbQI6jSU2GSA3
FMFulkqr2cOTyXR5ok0BnT5IQWPNRV/xbgGbMI0rLPXJeIYvJLHwjrJgQ0NKgEIbctUqbU9yMj3F
TBrFH6HVilG3/D6kZzUdbEL+MAv40OSbH7TvwHNsxEcElnDiaRxYrObv1csC+VJQR+wo2Z/1A23k
3q9kmJmYkVbda7wBWuwdKNImyuUWbXKNUI1jt07yS+16EbtrubcQnw9PTrCbuw8djzVGp3tH8r6A
C0u4bV0NmQ8HaqZLO/wCCNDwmfsO1efxPEFsSGCvnoev69bxDq6G75KXXOV8G1cQnU33Yz8rQ0Xi
A6QDV7RNsNqYepSHzqWHyB55tTKeiyqyweh29OXnzO4q3C1Jx9i/Xk8GHTN2h2Sp6/7HbCGZVvl7
J650DuCwTUIdwWY7438rFF8GQ4i583lpDHV0rZuJY14Bq4Z9/+rhGFrSTRpRiq8KZZrI0RZyhd5f
E1AR4lVO11aNQaAiRTTZVpUZveXW0Qtq+eOWfSo/2707sIlADiedddglC6HJSjfZiguknSLf1+54
Xaa8Pe6Nmy0gDHvTvOpAAZmNpA9H/fF+mFF5lPin/CNmTujnAisXVSKQ6NWyJNPwKg37r51zHGsz
cRtb+xHPUrFKIbMl6O52G63QW/NJSaSlWcvK4xmt2Yczf+i3uwVr4seZU+ChuwLnI7b6SklaRMVM
CXxCDN/SubPqjyVRdLURDX0f4pYNKwW7gyDD5Ka9m6MI0TguYISfPpAObmEcp8jZNFtjlyixEbX9
ph1vOHfvBIOIX7TEatrDP2Lk/qvH2Sc45s757aXpjSjhYYOouYok9Epi8DjTEtf2KccrxZH6ZLkv
N4LqKpa8VGaE5TZkuV+ow0+XU0mbMMl3QuaF51WokKz1N0KTsAZHP7ADVHjKCI5Ti2RneC90zfBc
IZRlrssn4+aUVVWeW4qTmOxTiz7jUvuud8eZ3eKN3RBgFFJ/U4dOLnwO7iKtpTwjT2iPdXHYW36n
1PXHS66snN8fLWJ94SeClDnd+/v5LA0So3lvFdZEDfb8A3TXRwZ4NCJkbC7vQAklwOiJWUt/Sl5c
MoOptnanr/21mPkLK5hXW3fnk4ZvBIF/sFJbWkhpMI98eU+SDXSnn2MjCjE1d8zm1qd2ArnQXvRO
enA2ifOEcQevNzdA5v2GT2/mAZTeDuTrg33gkG4tF6ygKZbGIpbF2cVFfkMi/jK5VqCbQBcZI8tV
zr0D3curxJk8/Kok3wHC1uIOqLiVUGGFrOcuiGvc9jZo0LIm65B4qy/sSzKzNMKaTGD89zHsihVM
cDln5hhBznMUTmbdKY5c4SYqiYn5oqpK+ArWibaMsJgHaKq8/FuFxvlFYGa9yX/d0+4dagfQi7o3
vnICWxdMiuA28Uh4H7LKlL/cLqDpHyqlwfWBI3fwaFqeep2DOUJZ9+A7Xt2BqYtj2yW+yxBoxEUx
N/3R3n+PxaxmTPJlznWlJZXVyOJis+h+FV/VBdamJDa/eY4hvfWGqt1/qSr0mu1VlppshdF0FZzt
QouyP9ndn7QCG95srHME+PPNCZf33JRdoVRGQLmkoCCTrTW7NZh53HtccJdXNVEte8U49duBNMD7
YcaYihrli4NL5SyCKwpNQbRkTgUPOlyWX5rbqZKG8M3cFRv5AqaF1+vZdgl7I+otz07LM3gRE6ri
v650XKbiWCFZpZn+cTFNolpDa6glb3N7diQBZC0RliF3LrXCrm/RFjsjp22RGk/CmT6FczzbptUu
JFjNXuHfE0qGr0E01zWQwoVkXtGVVRqGmnKAA4z8eLbJFrYOIw4prOTnPqBB4VWmZdtf9qTYWAkO
C+MSVlg1XbBM+3njkf2bwWyjWNRJ8Kxn7ldEsThEjJrHZL1fHuJh/lm/1wcGhhSHeR+xWOgDxo0J
gH3GrUW6FDxKe2i8RIkHtGKceW23umut1Vmy9/gMbQr1wI/iktt4ibHoLdvY9JpS+k5YRRX5qYqy
HnxiVlZEqMb2vr6TT3aVUj/y8qFb9F4BbBU/cM/23Q888uZjiGS5v5CCZjCBYiRDO6rymjBq8D1S
tcXgxzvTFoe6jRJG5ZDuzil5SXJBJz4sGo459JuWemEFltcAIjt9N8wVMGsUAc4xF7npcyecCodV
HClWxNXiK8tWlOY+J4w1xUgXfD05CkBDRO2oO1HDL1t6zpEph3apsU84Zle2U3Eh58jJEey7dEdV
E/1PWqrdumRzMup72HDj3dQCQ0dXvP/T2u3nxpAOFWXUSv7cEWUz+0YhYmCDQBcpKzCGb45WkVCJ
i/7Gqmc6+FfeyJdqIdnxSuGvU4but1bncJFUY/42oJdfzZ4RZtEZwp3nKC+rXrNZQnQXD38EMTnq
YfLE96CxjsTkczmbXrL1NYbVlKrnuinMKzGkA3iQJDbBE/4sL9FSWKWDEYQOW7rwcrqrln8wDzGH
o1qjRZZybfE4gz8hus82e8VQBoaJ4QC8uFd0I2C1Y3SEOX6bCgBP52jgax78f6ku7shwdJCiYH61
erdNViY1sI6sX7q8NL+2viaM6gIgCuhoKrRtKpLDMObs63Jeep37pLhsoWk2yK4FhT7LK45jTa3o
J2oPSWRBr+z5mB070z2zrPrJZ9c1jixImbk5W+048AcEtcF7zhJI20GNraa78cgwr3dEneZrFxaw
vVJTuA5giTTJ2ZNQPwSR9K+JV5zhjzrSB2lUn/4v8dOtqVwgB3ClVI5zJYrrxRsD0zP0j1DeKrO3
xAdfn1MLs7+l/GLFmsE3h3ZAYVV3fMYnPF6gL2SMJQA9j/KphZ/a0StVrkRg2qkQnr+fnQ5VFLqV
sq/EX92OjC0mHbCbsTgMvhjhO1cnY+xqflo2LYxhSJK4VsoUIEq9jLGaFPQlSg2mnPGkEBM5DHhz
k3QisnvZIdRKGkAVMTi3eJpEyBUcYuEWg1Os9dper7ZcNZlSRN0t6QeU4tOMH3q9JOOisQL8SdL2
bp/0hc1KLRomWvJD4433U4EDuOx+DUInT1G2m0MgL+0e8fp8sR9VuORwvG6xoCA9Dus893akpqDK
5K/TF5VWzkVUGetfRw1UAd90pFBa+Ju4hcRK85f/h69GmN/Tb8YMV1JNTvuyu9jgeW+Fd+ypeAGn
BYgrllPVTuFf4HiKDLAz9TbH/ElDZxS+3MzwS97JAY4CcrE9+ASRw+JbDd5rGm1czgGscGvvTbYg
ROURP6DgzEsRfsaD/HcoSMsLFRgpdLa5oY3NtW/ecfzyu6aBipvCvg65r2AhWaPnDLKgCItyK9pQ
8TuIV3YyT1LEYIOGk1/aZtyxyztPuDnqkMhPu1z0KrO/6MAuF1QX4IoCRGCnHbsxZ0KgomBIGlhr
6woYohWBS6nZ/9Xbc6iwVHZbWdL3vVNG8wICwWZiCuvLj5knG6SQzfEvfgTWScnEK4C2ZQuy/en7
DaNx62UNrPA0ImgFfJTM0YrCSa1ni369qZPLJO7YWV0756MKo+y+aMVPnw1iFantLQXdrRkyFPI5
gkm6++roll7uPUThvlKVZi7atabtAbNKSw1KYP+lcPpWEpjzCmsD+A67HVYl7NEKTgo9KNmZgVYt
Zow+IcK9HJCqoACsY9QxsslvmENqg9jjLJWVE0Womy/knycKEzmfvzi+uwCkrcQXCfzmvjsQ0jvs
4ClB9rvsME5jzpu7h+3ZmJ3rumuHbo+UgZIiv2GMkPyT48uekhPSuzk4Lsm+7Id6ch7Y74YLf+Xe
v0XDxq0ZZQehVQfIoHDSv4cuB8RomeGmWp50E2kmqB/TXkKkbIM5y2j7oMoIqDe0XuAjHx13W0m7
kbEFmu95Apsiyi/fIktS/WHIjKJpdYjRUzU8+oAuhBDyf8h8hyCx6Li0gUyHuvyoyJ2gdsi2JpUt
Ovymc0ARqKLc2EOzSgXJtkHlqvgCLSFAgf+IxzWUEdLujPdWT9eXkd/64fOmCrSDcoaHxbEJJQVX
C7iVIlR+2yOAPfnj7J+c7w2orY3naHG/KTkwFafPZwsc+nGpC290tSttO9YPbTh92c5qUJg/OxHL
OobhL/k2y8W6VTmD9Nj1g8RYqpe5ytBv+7CqupXRZaq+ENIX6ZBoYSZT+9ph9ioPMhYnMMNBoo8B
iLD2vFYC21ZtqBQgfQqhWCCXNUeYZ5YFgSMSxwqiBRljsl3Rc9E4owIpE4+acTWg9r/yQFUj0Wz7
bVdprKbdgtEFiUwgbcQThmj8MeMa4D+Tw6KqJRlJwVlmb67G2U+xmV8FWijeh6/amhXw2uhDvRtg
C0WgFlF+l+HsFjjvMZLbYAn+L/FunfwK1J4wv0XluVZxUSTztrx6o+AxHv9zmGQ2hU1clYpmzdEh
8nfPsHU7Z9UrTBBnqFDnBH2z+ZiNSvLe0Tt678iPclonKMIPLgLeGULVMLpQXoAYLqDNarHO5McY
snYRFadYjDf6D57nf15+xBfkUschZPZbot0jbvECnYoQL9ukOa1DO47a28/BZ2TOAuG9Rn4CLo0Y
iOQ8R65vIVh/S/JdXdYgg5nvpvYfIsyVBJzpBCxkffuIx6rR1LKYi06kHQuu1YZMAHsva98geKFg
eQBHDLlyitf9PWwGyDnydQ3zyjIj7L5NVr+Z4Uz7jP7SX1s9AWUEu7zm1o6zJ4xGE3691Rdo2BRR
bpL7vrFvbHTEegXC0F8MZWMi3t94YA+zSemyLEMp/6Ak1yE/wd60D/7OdG2qCzSf0DEf51Av2Zfq
lwIQPdYPrGHd+sN8YZ6XWVjXJcY6/TTUJLKo/dVUvf79M6dLaUWAymhVmjCFU4AKt33vq6h1NONb
3pM0cYDOtp8jjogcoEYrtTqxvboh9EX67m8OxW5N7JAOjgoaOvjCOsWnQcD4TbLT52MAHI4LoKfb
OGOPZVLm+VogVoPFnYoeG5rM17k0d95liGBwHSnGAIPdopCX49As2+SHSq0qIW+u37pZzSSBZzis
k7XxYWoQnppw2O9GVw5rKaauCPs0DySl6mm4jSOzPR5I96qJhVb2DWyzReanCsmLyzR+LsXm/Otv
u+HaMJPz72c0T8/Qssz1XbH+QcxwvretRe52OmBapzM3Yo0PN5/oZ+535ihbsdFH9KvqRhPpvMEx
1ROPjL7aySUI4KqRx40XFoP6sOYGhyB0+/wN5OqgWA9SRLhci8edbCi6blm9n1JqIDv0omBxL2ZC
+miB7D41MeMFtLwM9uw7lbgB4r5uwThTTPJ5wkcNq+Hu72xyJvZAW4qbJSJkcI064VXg2M5+WYes
NnzMFIgzNHm6IILt/lmXEL13amyUwEJy2FPbrKVgc3J8EsIAeVSqI0vy9SIG/HUsDKdCYlqyowuq
pkXP7XqZhheyxHX7zRjldV7tVDN6/aCmio6/7TeyrQjjFwrfjGEyHvjKS0cir6pnzzovQEGcCldx
GgfpoTNuTk8ighvp/gPB/0IkU2QsldYzNw1l+DnHKdSqCuc4mlUWw9yLUWev35PJGkdguYaz7p7d
7vR8v+1sJhhFZLDVwf7XSF7LoPDRLF+19M9gHOB1Em/ltl1CiiMhXznMVkXSciFHRVXCAcbLkSjt
gULlD2nMDANCX07edC+RdvAod46vwgNQUKqt+M420rENfIL3kIHcnu+KqRO/8hPqZqHwS7l/5X1g
Z+kqeS3hQjPOsPa71bVgZLDpNzabWoszlWrl97RMQ3X/OIJ4J76zRNA9axPdtBN4V4gP0DyxYAp9
920LNiYjYVXAWO4absELAHwIGORDAzNx9JMZD+zDswtl8Dz3H32vZVgZQP3ZKAhoimQ6S0Ejn19o
7yw47XNrMJidhuRRUcrppmqcnGXIcmijUBvI7/iBKdgPScU/n5zrk22QHY407EXNXWjCEaVAp/2b
X+M3PDL8SEtMKnfWj6DfzU3iXgSajuSPBW2EgXIyvDRgjuUXWh5ASuhej0JOBxqQWEw7hQBulATs
ZjgwMN1rVtSLixLMSReIPg4f2yJfnAFgeNMYy4cxlPOpy79a6JVxWV0fTXpSONz75azWBfyaUWzY
9/FaGIkJNt/bOG6hINRrLmqD5gpnw3SrVX4tol3gX1Urxqzshws4Unlhb2xdBrJ7qxjlkL01gU8q
S/lr+H4nE5VBk/vtZFD1wK01Qfb1n9Yh72xwuM6GuJsyu9g7bzcJaZPV20E/lvBOSFjL63zerbfE
qnx0WmPba1frN/RI9Fh4HVX/6sZ3+hxxWlHIsKcVO+qbIwuiDjVdwz9RPaFEbr9DkIDnIJ2FV/oV
DIdhdOStcTJf9WrdTXIQ4UpXwDohMVU2lH+hygbNZ6RLbfKA6Qk/HS/9FHoBXHUfsWsp+5WpSTY2
Vg6Uso6APR2TmpZWmuvgmwiX+a2z+aQZz8NkUCxYRrV2Bs3VVzMvlOYYjiTR6XMdkKD/ViN17n1a
UEjbq69Cm+hWH8zqoXZanAbXku+nqANxLb3p824FYvNFxEvMTaW98TECjuKeDczt8GTVrCDHKTLX
6zR4XCGWueSScChDzvtYzKWMqeCmM87lbo7fNKtdrAQT6lpwLp+dkh48CWGUsmwLH7fjWPVroaoJ
2gtWJmGDWxjBcEc4Zj3dLDRvnMC3JJi8yASGXsqb1j+gDww1HDFcPIsenLj4pdxeuVaExTDaFg59
4zhs+vlORLYhpff7SeKQEHXVsD0PorOyeIZOyQYMs6QbL4g6WAHNIp7GJffR4g3wYrofzL011VtO
tKPkNL0PxUlLos2Qm824w8JZk+MFotOr1CKaHCtmkaWq9ITt8q6WeQBfHAQYwFUnRgWngmIWYMr9
YLDZ6nsFNhqXYdwnNYkRhzcrml1XmpxEK8v6YGW0osJAr2V/P0GFO5BSGQJHmsHdScvq7sz17MmL
RzODb683rzCcs4PERz2xmuTAxSYY4C5t5KjcP2xbktZf0fWMXjIJgLvkA6YkSb1E/UvrJMBY9W4t
sDgCbnL1YG0vyWXLklK21WgchRUPRSbASvc90RTDoJ0v29TD//fE3yohLylfrRvsyb1T1obaALvu
wjysWTKCzIeshtd2FpAbSS+X4vEpk/wuQAqVsRaRwKt92zt+w39vCfLnHQui8cp0g20zhUWEEWOH
14HLkv7nvBFUZ5xXO+T3vc4rA/5ldPp3YxEci/Pjm8F5LqJ5sOc78cxyoZcR4WJltgm2byh/sEgR
tWPNEJj1N7lAu7ITn9ivo5j2dJu6izVRrE7cyyrc/FHf80aRiJXrr59Twvea9N4DD7ngoeKp1+eP
ePdN7PLYZ4rllLNZyVivZtDRL0uFUGn0sgljtlRML/7cY76V+0hT5w8GcJISUhxlYd3dE0FImS70
ZLK19aUtsQ5sG5bu7LHkR4lvclyt/06Ks7e43IgM5Jz3+YbVk3S0o7kv9GPXhCQQ/fXX5nFbBGQN
8LMNJyyJeseUm/q0Lpw9WJR9VtnKeNTLs2C25NsniFqFTIjqW++rBa6btl7dFf7z6FAykCYq5H6A
T9gMY3hYD0HJQ6dgW/YXOJly8TJgECcX7NRUljeH/jETY8ZJ7BkNiYWWatxZluz0SZzApp9+RCv7
2xv+OVmymBHNW0Xw9unRHraBwPsh1U4FML4n70ym1rLrYOhKycIH7DCsIoVzKlUi1P8cw8Z7m8P1
9YBMliYbohHbNJOsyBcJJyUWBGg97nYylIA64cXYV1UH7RP7QXSrt9fD7A9Ebb++DaubxT/Kgbdw
eJEd+fpi2DzyJQeR7o56dasyZhyCuxPNo3WaFtIrUsM06kVOR7mcqAcVblYlewz9mZXzKW1bzCuq
FqCVgrLEwzuZx0zzJwos2cJ6khMh2k5+7/1h8Na5pvuQtxj8g5nEKb6ehdas7n6MOXcaeVBIz3Cz
s9jOCNdxAGkJWbIscQF01QZRxK4f0Xsakmm+ae+/4fjU/4AAx13isivKzMevDNO+PQLgLrKSPyVt
jOeNBRclWErLgDh/x4HFAM3ELkrgCWwlF/VZeA/Ix1ncJjWjrEihS1roJKWklb7SDpgDkB0Ak056
WLUdNW0uYflQzBcw6f8QHody5qdcAYsyEpZCc1SplrQ44zpwYtr+5EmbUkpvA2SvK8mEH6+P0rsV
uQ3VmtBEGr+ajfUEtcw8FtbNautUNifs77sAxJg8nfhjaC2DXz2wqqHVonnS4qbH2tCrdw/kIw6Y
qhsGKRwj+HfAuQDBj9fCvTviIWswj+86UvLtN+0ELlm3vh536G31VoaPMPhiQzRsg6p+DJcdqG4s
jzL4X6tkzvTr0xUkq9EklIjNavNbWpXOFBPTAKSYQCDH60FyHs9eh75NXbVW9EVlr9X8ztcduSSB
rzK2VRl8PHS2gJ+G79MsZAqr/d0xD1Tflgnxn4rVjGGXOcq95WEeimKdscEBNxevjN6Fkl3XRMNt
lAniixlHmHseFiNY241R5suah6nLw1mS3ck8xLKTtUeStt2ZcWG+lm47EwgPX8UgJP9zdtcu9kYU
VKEyjWbrJX0IeD5os0HYXaBEVn89k/9YpJx8i6z9yxFHD3UtRy0LBMKDB9YF5kwXUjlZK3owcGOr
4+Iu4RCBgxKaxozalbyurJhzWYcGWE3z69+88gg6MTzHy8ZJ3CS8IEfDSCxbaPhdr8mP8uZ1vlyp
JDbni1YvUtnChNb6ndKPmi5nMHrDiOBgkrRetbUfMevIdWMZuWvhERD7faarJvFQDLTJX/TLiCCy
qhY6Ag9dy0xN4JaExuv/Eik40s4daeS17r+uHAQSj+Z8oZ1YJGuE9HCkZyfCXNaUmYwMpYV02FuR
4oFNVb7CWVbcLgiLAmcl6CfDewxuCPESMKJ1T5ubyCYMNJJQImoO8VBZuSwSmFoZBaFe5IeYXY32
Z/s7TMixepw+yNIOzjJo4w8hKwm30xcOxF+gpcBefGW215BVmWwkuQwcvN6ZhAEfvCGN+v8GZHK9
Wu/4WvPG8icnJ/vb8peRsY8xeZrs2W67Qs5m/dkVObbRB/pNMCEiKGD+IozMhDbtwhbcS2SzTC6y
5ZoULjiG5XozEcPfxYHSKFTelP1ZHoqRRAd3uJRhaRGpRzt/mnCxwsSQBTlaUXCGE8RvCRnleZWX
bXNkw9GnG54Dwi42z3jwdNaMDmvDIKdnz0fuek44z6sIqUVZQOdihx4KNjTybSB3F6aTusTfBDXL
ihmb0zIrWGQLbTt0rR5A86LcGfy8qnJAqtV8f8/yp6ys4HBYLSXH1Z8GTl7KtYZ7YDAN3f9pQtQh
LP/dUnKKn4Pcfp3Nhmm/7levNGqVqbw1fImVGwPD8G3qbd6ngyopPbH7s2E7jOIq44XHVm2V5EYB
Nth2rA+ATodx0BHyBX8kuxfemkCt2D0Vn0/uftRtHNm/FSmItU336yRsnXZqo971T4Zal+MTOO0n
Iz7sdL0iis8PUeC+n39jXckwNQBS1eImvXofplB212+4pf32/qKdE2ntDfVwym6pSjyjtg7/CeQw
Gdc7IqdIlJlKVhrDJxqIVaYtLiqrQfQT0JOnvM7TELrvyf52dpPvwVWK2QzZDOX/QJeZ5aQRgb4O
EODzV9ayu+wtVt0zFmCSQYwSeq/4PI/tYGpmXXAe11pXA9JbbExicnMMVQNlAG8FxQaos+Ztobwa
5Kke0aUhsKid9e/0ZnZi9kjnLK+RcSjZaDrhEKwuDaacI7H/E2DdnhIQgIdsabXp6eazmFoQDiAE
8e3l+51ErbUZyQkRk53ZXQXU0c39jVRYfpUOfTZNfQ3Go2LJvTyQ4oglQE/vY02zFGhS259fJK4v
M2sVV4SByaic8OYTKMSFglgr8fY4m8O0VK285WCXKWdIoc6/422M2XaE49rQPO/1GYX8FeqIIPrV
rRkXb2F7WEQEcjKyn7xMyvLOHc4EWWiiRqBRh/scaeZvv+NtkGvB+H+50FdSH0ZU5oOtfEgGlWoO
itBS80ture5uHetIei9khPmQpykI7qaVQRikL5YuBZmAfbErwbkQNoAIkmPH1u6Q4mXQahJyT207
A2D87nz+5TpKtujxVAj/DlgxGps3aHgxMmX7hTtCwJr4gA7RwhQW4l5BBFfP6d1dqbSXq3Oelt9J
OZ271O0VPEW30EJ9BvJd85CipoJNxywFYw8EK0jjB1kmcFmXz3zFUyKlVtSJ+ceRSe8vw7aGSzk8
H42c4maskgUW+uH1YTxq+8EdPK33jK7Rdoj32YiN1TAWRqG37xPq2692DlRjot1ddbaBYGSlD9PF
pMpb8mmEkn/CLyfypu7e8HkcINYtshOFwaJ/JDY/wSmJIEI7M9qXJxhjQYjFdINLl9rZpwB20c7P
zWBbR7O6cd+jbUbpTxU06Gxm5+Xa1u0ajkWrgcuFW99wA6DYDttgaxPBUDzArdTEEizU/PxGKPpL
GgmRGv1FxxSj7+ovbUAYbkrb561WFUI1DuWK8P1GD3uPxKR2khYS2iYrAopz7jP82LzWWaF0l3FN
Arp3fVv9exVNSvQXrnY/L3lkp+H5n+LqvWBnM2s8zRI7Ypb5He8dSpJmsVNhFEOSW9jyw15fLJZl
kN2MAv5GnTxe4a/Y+YX7n9D7KkOFqgElZAuJBX1/lWSvI497hLORrurEazo6mfnqxsnyCIEb1l7b
iHs712jTwhY2vNe2ZT7Zvl1stcx/ngxOoZePYD7UVmHJ0jsKDXJ2TLUmS+JSlA+EKorCM1ByWmlt
f7eQ+oMPeYiNNkJoUCwAGHtQbQO5M2bcf3jN5aKoYdHviIl1FVdkJlFWq1lKIs8o37hJv/vi5v5D
qw/dMVsY6MAGyLr/nsLQqFTCDn83ZmmHsc8mb/NloF1vpcNceI3Bq1V4o7J0OFGNGs+XtfYFaV50
ysOKjuJsgfzwCUjB4RFO/gr0vzjt4goMVi0fwmBZz2xayTRCJb+b+klJFGIlziXBgwmPtdwNG+uX
VdLoSWtWmt+Dc9e1XPmDVpfdbz7mztSJr9UCTtOzMLFh/XHT8uByk4D5b1piIVqOaPs75TC4xGYF
2teJZlEeXMLeu5Lg4c/bnZd/SoD2PQJAV/sHPKYAb3B4QQj21KMdwTSPHt4QVFQjzkmOIPj0fufH
SPicK7Yg1ML3NcqzCo0KBT72xpnEBSxa0B2hoUB4IafU9VN/IrLrIAiCf0gZr0OgmhmPeKblgNP7
98Yk/npgEAUHAEvH8HhSPbkN53AMNITCQXU9EkJ0umBABR4tncglCi4rTv9NLHpPBF9SQ6cdMBs0
JSyIsgbQsu+RZPU9PNGt/c9yC+1CXayX5a1ZD7IHqheLcN4iDG2dSNiZgIASZgCdTVCQ0cAXWOFR
BICIncRk2wPtKQXDwX3SfkmuN07wGI9dh9ili1Orp2NaAXXrnnLdCvpZ5aO33BGDkah8NXVBYLYH
hhnCzTGXWvC47u4018nHZJ22LMBSl8IsHQbcInnCauQWP8WH0ZmkGK54in1dLD6N/cJWRdMm0J3p
SxJBAMsSQh7VDe39S8OYvE4VAxdKFA4dMVMQ2r7jVuVSYFxPPBVv7mpuNT8XeXkd0kQsEhZKo8xh
zHLkeC+2STyK0sV8Catxq7wem1fhSQdOlmtJFXwCQHJ2Qrz3ON1dLRPa3032EJPpZC+x6k/n4p/2
BT7au8SZE4zOPIH6mCGdQx6esv7o/AiAxCrnkuVr+QED5al0E09iFqYQLdVFau5qNnavpovcV+Xa
a1dpuMOG6/d4VDz9o4Qrtedk+v1vuBi4caA2sT3ILjdPFsOaOVModGtMuY4xPeu2yZum4T2kqbwv
L40u7z2Qmae+xwIfiMbsNLhbKH1Aet4qCnyP5cgS+iGNdQMJZyqf2fQkXB9PM8dXld7KHh3sYD9n
56+N9ouKqNhhc4+wkQjlXfNammspg2QQjBXh0nilAbE61veqyG7Yudkra4QYy7rVp2UGiqPFdyN+
LFgNkPitq4xHgRjlvs9ePDr2+ysvzd2a1Gb+CmTkmf5wg9LcHwXS/HXWll3CfY2370ZIyLo87zah
aZ6EWEdbBfLwUrzDW6LuN8W/jvTDpoDVg2EMEUJx52ESP3MDWN/19gJ3I+/Z2YzJaVvSLeQ8LsSf
MpuSoHYCzBl3WiQQ++lwRr0sNGHnAWpBmHJciq84k488dtPk7cfN8xqnw93ZlrTzB1mEicBq8Pmo
/UWxu457CWvum7nFtArzd+F0KUExdddGqu6zpHzJfkj3ptb/QdhvmnpAwXb/B53LPI4S4qOdHCCY
AVvvWuyBgVYEa8tRhSaTG5pAgBiZGDnBsKm4OTUlKu5ciWtaxgVlsYma+dBMosb27wzOZoHMHW6x
KzE5H1lY3CBc4YKz17fNebLCx1Ug6Nwf9DLYsGHVWPGNmrtEzBMbwL5+2xf8xmqd+Ir5ccTCyD2e
DkG92i8502KgfRfo/3ZOsKFoyUPfY+ybqBbfv7m/IFCTpZTFav9ZgxOSEtsXWH4VbcVZ330D3moa
MLVwGP0ZuP7ljTeAYCsSIRXHPjZfb47z38MXTpT3FVq/d5VOJiNauEobb5+fnb5bSo8gA96UmQvf
E8T8ibUXly9eD2dpxkZGc4QPFc/geRd4po+fm63RW9VZEF1So9Wwl+hL4qoJ54XOt/+/HIgLpApz
5gN+Xkf0mbTx75eoysn+j0IDWxhBYSO5twdEublJWkD2H74OzPkMxuPn5+WMwv04J8zr941WSurk
AhzAXqoh3ZsBwZYAM6rsGAWrJj1zA7sSRx14Lg/k0FlshFJSBtvIy0pCaxAFwoq0W44ahvYmrLg5
yOhZw042uporwAf9LDlwS5nljjMJ9gvfD+cPvIwessnzPmF4ampoce5lMAdnJN8ouNraTIGOrszl
SVfNyUKSnzwZa827MJp8atloLYDGIvBbtRZXAv/AX2Z0qm53YvmMBXuZh8Zxv0CDKJ6vg5P6Wnrt
GmB7s++ssUhVXQzQka+VFQSJ8RrrmFAhhuVxkfkZ7vO7P/gT1cBCn9UIkAVPCCQkpZosPTT3onLS
dGcOXgvJGj8cciucny2QwBwj8jsbj4IEjAjNFSnIi8S8FI3p3DkfhGTN5Nurlgp5Y8Djykkw8ADg
NdAt66umbQlJiqxHI/KrV7jVGUv3MaWEP2AbJRbc0Fy92bE3TlAJxZA0PKajuzuT0WoCiqZlU3dm
/zHe9WzE5TYEEVeDvmEHsIMsLrlC8d4UUBbteRXXtAgJJBStrUNTBowI3lEWRAhGPh9L9XHk9Gy8
VaVNRe3S5Tqj30gIU9uIIkBNr4fTqwqDWs81GONMVpZCbduVeft9bCEHQUSxllrwBTV9bbBbcQg7
My4s+/ip2JuqxU+Zo3VK/p/oCrNalrNAP9+7vvCNLvT2laGbzx55Yr48pyWGzuFFGcNrOJYSkKPz
asJayxJRzlNzfjJVbef6+hra4oEL+x2WPRQ4lshbs4Ui+SERWVwnNSFMR9lIAAJbLDIOsuBusmAM
ReX1/Ynx490S2f8VqTmraPczrJlPfJb7I7VT6Whvy0UkEKmnJ2v6GciGLfie1cy8J+psSO/5sVxF
/DIIitqHWxK0YhgMtZm4p897U8ehEKN4kCjSFMG1em3sV0cIlmFu0sDJtvOJC2KZQoWUAUktWuMr
NL2lRa1HoRDpQ/Z0pOfr8p2Fv751gg9e5qRt8GxicotWUgN8e4pVOo5XSG+uCLn5y8ephc4dfGlj
c2owT6yIKN17BOB4j7X0nzahaUQ+hbCtpLNIjGFfiIpJB9kvuZHKQI0N3IxhHdd3oX+SCOp+ifEs
3WYa8XKUnmsRqgxVvUUM9Cs1QKAHKYw6oBcyek8RsYeYGnvhaUYCIpdyCmRNEUd80xUGryKSEjo7
wKBz10Y+cXdTI+11wUbio9IECkSJdfB6iTei0y7ydyKW4WoKxYY4dcaI1L6CVl9CdkhSdG0w6qca
3+M4i13Z0ZZipDQxPxJvWdeXh9DcIJCnqvD3cE/BzOpRvWd4qQvMyISlph5nBIg6qvUr46HS509n
KLxsYRjL+iU/t01cIg29FO2p3epeI02weCre1MtDGqDJRSSrpHHB9GBEKtRmMUWDUXqN7nLatGTG
XyvNyPcD7uKD2TeGbZ88WNXll+JckWnK1NBs2/kK/xwi0zoI8yNvNFTnkAERnKmQSqrjdem7n7ra
MsR8lIL36SAIH3vct+jPGRhW1XuNxR+/gGdSdAGUJqPB5eHFvpo82mA+jetXu4L9o2ZdYSdY+C3p
8oD6O1zeWvap9qv5nmIUf/1Dg4M12L1VR01lZ+QNKb0DMPOgo+/YkI9IJmL4DUiLRZkjlHV0gIOZ
W60SR3J0ITiupqLzukKNQMwblPty+NpvnXLZIv6KgBLQwqw1DLssd2zInWubCmfIfg9iWTT5lH0Z
6jpVqAJxgyJh6iRlX0cgvnS67Oh0YzfY6Njd9bPaEWKT2oxHNWFIjighkdrJ96z3GEtIf7VabsGH
ZpS0UhE8qPc9xAyNfS455/3AWvSR7MQmi9ulYCz1WD+Frxgamzx6QC4sWKjdzCs9YLTEvb5wqAyU
qUpMB4NiPKjN6ELxUJi68Mc2nDvieJcTPPNdtnawNG4sMsjDPtNbKkzZ3ZkZXtzheMWVZ135cGs5
Nk9C3jgYfB2Qq7R69K45JsTEqmZvUvRI5aiyW+B0RHHBGo7TwgTATyQhhLTHRsE1UWJ6vlT8ddbK
1uDpAHtJLTSpvq49m1vXOodydBJ3cB71xnOzBTLbz3hzYDOfafPTffh7w6iqlyBFrJEXx3PAX5Aw
spIZRuklHoR1D20WhKu+kGssBcg3BlmVFLj3JG2xMAUu/RQyKTil8w5KrLTFJfSi2dAcf1FTD1PP
NeZltDzjCCJm2gNZjMfg+v5GEowYJ2bXCwCDRThxHmCEdICVw0BEOWkQ6us6vkyd7FqLnhrSDTp8
9VbF3VHbjHR4DOopGH9VhnOOVKo7LsRL3sf13AIVtPB+r9axj1JzSQVelFq4Ij8TghUvQYYeuoDI
MhAtRLqvpK17RXFRqEM+jezHNnqVjS+FcG6G+Kfa6dTHaSYDrTS8PNXDwI/YqJDZVEtNZr2K03VN
iKNqANW8V3Y2F5wdpTx2y2eS0ILqT2JmnpCiQvKh+9DCaVF+B/bg2/yo7pq3tos0aUKIy6NL8pht
ebbAdjoMTOVS7nYrqzWGOYI7AkY6m8/2kYIQqDfOjzc6GHMCggJsy/8reNCrzBUVs5SJ7Myqktpi
8qSwsmJ9BqUXJGqAuqdrbNOE5pkcdmc+KznbgoA0FLiKHQird+8hl99mTnz+1XQVfJnczPiJWjSF
/vZgY5YsoclCPlh9lNZvJ1lXa6UqxnNjiDUGWxdiCcAp/VN2HzP11TDwebU/Po3lJAohct0bf104
zS8EVIb7iZ9yFSrgkZeNLjl+EX3xY+dfK6X7bKYA3Ly2hTQ1J2C/zZ1H/OuhFeqIjTomr+YvxDoM
d+7MQMhdtkOt5K1hnKcIsGNzgub76yCl0bn/Dk5e9IgI7v3SAQXyrRyrn7DMEzFTsnUud3eWj2zv
UhM4h2sCZsPs2/01vUtMbj3ieOMNBhTuPHLBLGLuH28qITG/PEw8f5O4CmieHIZvN3bdl3wh9sCv
1t5RzvTnFq2KaOvqsRRi3GspPhOtZWiB3XSgR1iWBaP/qXOXeA0wrplr5MaxBR7C2c9gL2Rhe1lI
nfD7S0nqI9lqby2a3FNwM86pJIfRGkTQa4f3EPSsMg2v0PcCtIyVmBfrmBNSUjH8eA0e3Pj4Sg1F
FkXfoBG8vhVk9SqCrA+2/BI1PhOuQxYMEe+tXewMaqFXLn0KDBcOfr+0pFc4GnZ+Hm5w5bFmu+eE
m8ArRUdBKxhTnD14t8ipNfp4viSvNawtqQyJtjxn0V24TmNUY0Xjh26Z/TuBrhZRBtaDPIdXvBLc
gcJsByxVw9aJnD673mDuqlZUmQ5Im3ZVvCjPE2KS5ngJmhPvHRtaESZq65Ode6MzqfitdurBrqPX
hhx2ZuL6KuFLNbcAMkIOhM+UyCPK0Lb7D/Qh0iQ8qq91pPSvrZhq4NkybJW+Myrp3Pon79KuIEzD
OUZO1z8PhMSyFSwO/ZPmiTx8F5GDbCIdknTn1fHJ8nq/fM3OpkEHhL+6VBTgH9mtNb6AXtmZsAJR
zRV0OjbOmtO++IKnQ9N8HwhU/XelMxwYi5hg4S55UXSo4GBvQGI8aWa70fakB6Gr3Ojd53xiVQ7r
5zCyVuVIYQR/oKZMD8EXhl043Z3xc9lj/d/IMu6jo9+Fkym5u1nKK4+VLD0YHeB0jWmWIHAHMhsM
JOpa7ZImUdxj0mFVrDkub2L6dBJrZYCBUgKOMFR18ZwQW/n+zJuq1u3J/OFp8SWBWdumSdL4QM1I
hhdDqmi+ACscaKujJNY9qIPtbRqyNFK055MMM8O4bioJQ3oGWy+1eZOVqzWYJLwT0c/5YrTCk+Q6
Bd8X3/3zMpEq/oT9njRFekepVxJ4sgl+lQYECXGMPLv3sIFjuX+3EvKj98pC7mDsRpmr8eNpIFh9
fdhdqgqqjUhzs9+51smfX5roFHY3uYGNJOwHNbJrXSjyqmBYye0B9KNWA/0Q+kmc+AgHsZy82W2U
hXuusCVnpZC6eE0Oep1Y/pfOspTvwyVpwdn9uJJW3sPpH2MDmVo8Tu9jJRx0YBHEl6HKKkDu26d3
mk43I92cdWs3OYPUAnVE4n490TgpZdKyzBUfq8eWPABUAh3MRNCAia7x44mpfHrWbm/K86rUlB1O
FVcnCNoy9QmJAKyj70vxj7psImhm4PNnKIOZZGKj89zxJYbqSBz+1IBBySzaxk8IDOa9NUpU7do3
/HgeJHjoH/CvJBu+GwyDg/K5M091/8iAmqw/BqNwyCNeQPDymX2//u8CZYlLwnr7I15+cX57XMsM
VbTaqn6t6Z7h1ANc+QabV57EaqX5zAzAqNG4Dgev3sbIHeIgAIp1laaDjN0OdJ+eLnAdujwaDzBU
KTwqYFY+58hUq8ZRnY+hODjegQJ0Fy2XwWPlYDADDueumI9lHA7GUoUPhfhNi9+B805D5noUk6rH
jXrpmt9EzMhYqw1Juc3w5LXjs8R8TxW62Wjt6L7KDCtmSOJlYuSFeTc/859Jfu27aKchfeDbFK3n
Uw1vzlvGssgFD6ma/X/+EhEiftW0wLXiF30JKf6GkJq03zTPkJ2DkatD/vS+3EObxhjROLoDG6bE
Y33POqeoZh6R2eKqsO+TjQ9dua80c/rhFCTjlafi9iMMUGioLNtCGvOH7Lc7trgX3cCkMcmsPrwP
fbF4hCD60mFWbw2u8+g1YBTtwhv1JKKQxCEcKkSgSuuM3IPknfymxb3zI0Ys6t1tU3s3KcK4aNFD
/Gmb7PUkJLd+mey/3OU+CMxx1AyVXyXfMVlqJyakWTMYuxyr2ziSBTelayDAd8MJWslN71DgOmgY
/mCQJTNjsmdHe/ZoOvQ1wcXcNJvSfYmd4n2Xtl5uJiB+LA4JFa3nIz+IbAcE3xeJRsN3VcwjY6Ll
Sxp0b47cSKuBKZBgvqReMrDh1aWzMs3RSRiEwxOnEbHalrWA9D1c3+azr9GJswF6rqMgxZ2X06Hk
j+rdjMY0syNisqeV5C2yp252ZHANIJjeMKaH3XSgvUIBC6xXjZvksA+2CRFXGio7lXI0PxuAI/Wv
YcaTFwfMicKd7XFd9Yp9/B22y/pp0T/fEZkT881V7jA4bJoPCfl1NUyAWstDhsphMivK4jl4sLhM
cEerSkS2WTfXk5SD3LX3oIOboGZRGJVlKf6hbHse8EKBmUgnPh3FjSoQ6e4MdL0ncWpAERw9QKBp
3omYVBltarJ0QTT7yoJU3FbDc608EQGP/PfLkduFUM+JIS0fAfJV3Z5un4ycOU/mDug3StwjU4iD
pmmL/H8PuRep05voedDZ+ckGzgjBpp/2vPOQdMZQl9g5Dk1L2NTYEEa8Qphlk3dQIXnfZq+6Bi3o
3EgYiUvAgCvIeTml0lJYZMR914j1PYBKCeNaIbRbmAC/+5pQpvjCxXC4EpTAD+bGMamAmz+zVB+2
nU6iTTJFfGICx0hzVXTooMSE9fcLDMo99Uf46GsBu7ofirUeO7WCallYP5r/JX5/CifyqbmBySvu
ihdtgY5x2MnJ7cvREddGDDLz1U8H6XVhUbhbucYibS7gf+Wa7yujWX8evfbE0yh3yH5lGW8OqeH4
xM0ON1PN5ScuMLQJzYV7SL5BCMG33ZJL1aaqRlCXAGYF5SgZC9fJkHbUAdeoUR8a0kkNmGRnFV42
r9Dv2nvtBeeAVeehR1oFunHCwdPtTUfcg1oZ+lwxedrXf0OgOtN28hyXxVcVs9CdvR+Z2KtE2rgY
rZZ6e075maPxpZdYSKzB94HL0J9i9nTDdBSaSD/pPfKxdKYeqPsh+Gb5AmiHDjQqz2n7QXLqBt1p
0n/AKL4McZl1i8pcfDvZ8mc4xJbMUdHTTVSM7NZIBmyrlE/vrm0udQ/pg8ZGyZk3EyphKzyL3HWT
0aug6v0D8weuI10KhL4MJ19wOncwuTpEKpVkyQlX6YqCqFPDX6a/8yLVDpiZ0WNyfnKVvWxhjO9w
vcvX/73tqdNxEIzk6r0ac6xpBL6s2Ob/MasX3KUO/y3avPJ4MGBOlRFbDDnnboEwfbZBxE4LVK8A
R6asfwpNA8cu+xSt040n7Sx5mD3IZfPXaknL5NQ7Bjt7Tq7lP8xkrXbI/3KS8TRPc0kCZSyW27G+
bI6kg6OFKyiHQMf/tkVkimumjxebKfZs34LlhslxcGSFyrp3/tIaCFhci5Yj5jHEXlitaCuAXQfX
raxWe6YiyB0HeolwjV/QHFL7aGHl2DqzkNVyVvCbM0LpM3TI7s5sJ3BTXC2NMd9O8yhs1NKbqJQe
VlNxMZN3iiq6YH1EDBt7m7l3V8L9z7/0/pGvYhODJOK+xqm7xkL6xignPHBPaOGZMlrAoN7VB5hg
xSH+6EekKGAFW85EWSKZ59leYr1VhHk5hHJ66LQiybsarvmhR3u/0cIQBORUA+rFT2wanp9PzLq9
wgKnegYgUtwZM8e47stQXk7Xj6WQbHnIwrUPbxvmZ11sercItXFLrOah61zH6prw1/pkjITMMbRX
qK0LywkFWRsywjsVdpdjztw5Sy2El6JPB14CzQ9uA9ui18owlvTPbYWj4XsxvO+3QXynKNytCSPF
9JZ/a2v8Ucjh5z7EuuG3E1bOncpYLAcdR9wOwSHc7D99BXTEvLEYA0PoA8ErN3UrQbOKV5C/BKDQ
6D5tTTs59BSx5iQwaNpuYarKk2FOB/d44zVRwBr4utZRraVgjN2/qwT+DFUTKOiKAMJBMUsucMaO
6hDw/rx0p0kH8VjE+tkmyKUVEGy5S0d7Bv7vfA1AcdfzcHverEf0qe8dpcPHmIeo5EODlw5Drosq
kt7eTjHrm6VgEXE//GfdsmU6LDXWcxk4ZhYYmdDV401n/84ZOUrnghd8nLQrls7G/PgYDkyeS1ot
m4T4N99qS1oDtrIHuE0X0ZY55RRLnX08qe39KEgXwdI4maVzsa4X95g2D1Yfur2p7xW07p6Nci9G
OrmEvqbSCMa++H4zDcOTW/0SOKiL12xNDacAuWcONx+WlLxwDkJuBmpzZTRdaH0BD0Y+m4fem53k
TWCBVQo4kWwbqyzOHP4lzmAJ8AfK/mvYDIik8KiWwBH+KU2DgEVVU738z903IB9b0WbFUFx6E9M6
TzQH8oLeOJAOTCGuR15oV4pGeGNG0eHZNZvWbhQd5HA4lE0Mdh1LoNjphX4mCE5Qae2QlKQz4tf+
VrYKvbiVfCnyOfYd7AD6wR8rgTv5Jt3GioVBilUfo1x8mDJtUy4+o6gFl/3EGvInMrAGXndD8/5y
VncKYug1JNbrrN/tkYGreoKEab8cjnwvweTGeG3J+ie9hciNRYtZjl/VCepx80c8qVvGsKIzMxkU
DlYcyaG3BXVndAqu+fn8JWgGGel0nuHKcUn+lPRVD05TRHgdEZE5UA13UdO0P8fq5NbKxFFEiTIb
oeZNI1aZzYUtxyFa+FDiKDsfrMkfbW6y0G58+qba+VqywdaBAnGJsY8ZnN+QDNaG2hsVhOH1+dtL
HSyPmAly04V36vKQszc6ALPMYFKV6Oqy9pLT1Vqcf73IyerjeZj7xW20fdKn+e58X5WO8wLvgNtU
mtM1sZXrI8Ls79KdxlDfLbFCuGgkHADhD2clI9l+u3Dg+eHRKOCedML0Q5MCQOQTo1gX4TtxN3Xc
cEbYTJXaG5KVMpA3P+a3MQrvKFLmyMUkdZjksLfXCJXKCN2gex3/hsCYjygJyh+XlbuCLpZoTFEi
gwCq2I2LEUCsfJQm9QXysRrj84bYlLmsK94U5/TzICZna5CBLCzv3+MPQcj5RFfg3hcbipD1v8Qf
f6TT7ZkusfYhreFtLcJ1sYTXTpRcdAK+cU1h8f2uT2e3Y7aCfbpPwv9sGWdNdrau4C3wS5TPdQLC
HwJVoCccdddkJw0yXpyEHOG9INfzKlnDkRzsOphqVXDSpfA295IZCjOfCYRuIngn5gHWHP6RvsHg
gbP9dEd9LrqK7PPSQK9vs+TioJ4C0yZzKBg5yqglyUMPHqNctddhyypPNmNufZi37/BoDEEXmCOY
aQByxTuorOJWlo4FRzPH/Q8p6acqv+Y5vkBnuSyx+cawFKTVT64+/TmEcb8NLvHGdf+XUHWzvD7U
tApqRQDKB90jK1CTH6KsobeuZtrwj5GMLZEFFureC988swbam/1CIEKlQZgzYETgkazuFTAvfMgb
dfxSFrxwPTwkWx1ihLZdv1SAXq3bslSua06cHX2rjmaHCt7FuCwpZzyDDg0t/bxoZRkRcbBmrY3R
ohmkiVu3BGV1RziZ57q8x/d5a8oZS2Fcalw5MsvexydKckVVNlzF/HNdv8BBoS/bH/+Eoiw6/ee3
+cH79ul+U14iAGF8bvLJIcXu7vMyY6MzHVG9Va89WGzBjc/hGP3ToeGiv8D3azKLWDe7OWdzI+ye
r23eveiAgSlFEBQ4pqBx5uAsX84eGAvkDHOwX3P8YAKJbqcbCUuS3Cqn6TPCGWE6eCBK6QLegBMX
SGaofy81+GRVb7hltPqUR+5Lf5gz/z1EOWC1Bai1X0o5GAQLRgZEuDTV1GsCbuIjNuI308G9N9JI
ROA1miZUaEh4ME7jyYxIgl/063CVyogfA1x8w3CDOD1/6PVHdGXJLbWbAP/PmvKtxK8ZSvT3iz48
iUzNkNxieDUB7YwOgN2dA1QnLrsPd+E6DwfER1dIg2QSjix+hVaDEbAE1bHlApnk406uEacQ+B0c
f2VuQT/k8vKjC8G4N4oQagtQMZBRsVZcrcphy5KkTjSlHbYePR2JFnZGOE6M7xbwAi+kz6Pvaasl
iaamLS7sCa69g2sxSIpCEyHacE3e82jLtwck0VMDijjbOxx1STy9mD4SquVqE2I5kbZA2z7dBctv
ok9Lv52eA0XBxT3x03yk/2Y/JJneGwZuiBJCVLCGUmQBhUG3vujiB95XmwEISH5Ht9e9L4gGtzuS
xwQMxTs5VqI9ULzSa/ZOhd1Ya0Y01pHgv2rKZSEezB6oaYvelCzEobMs9tl23tDqiVk8supB0Kv7
/gMFQuyti8kww5WkgKLeUn0cK8XTKeT62tx0+paLuGxXrUvdo7I+T2jgkHgjWQKuFFvzyi76tTd6
P21nM+TLMndXfm+aMUhHriVRGgy4vaDm4jujW451LLl72pzj8enQjVj3yE0o2UwJ3JJmF9PwRQvu
rc21JwVAyn6XtB7zBOd5BwH7LdUmUnK3FpSrl+nzIokO5z1AD1lW0RYyD1YI/w+1E3Horbf+oRsI
3FoD/LSKhrx36S5tn24YFdiCOses1XlzdmMRF1ZxHkjk42ci3yr6Dwt8tOgBBHLpBaME3h8L9/t7
YWRw9GGFh13C81rkN6erd+GTwubCqpmPdx6IqkGTWWH811a0O8wWky5JBo8DpdHtkNSTETY8vdqu
ODqg1tlLKwK1WUOMWiUnAkQZeNw5ua0fO91EKP1/Ne7iSKgGjv/dO1z+LqZG65lG3MMvFYgQF1FR
QPxlWEveYjv1Vvt0f1q5LLgZfhFspyJ2eYLHJX8La8HM9iO2kK25FraOMRdTOvj2qSb5XpTjNPDg
rguyddmDheQbB+aEwRI9DQNuOPmZBR3NgXtdqjs9orhqFqKG97WshpzakdHAUfNEXZQpNWu4/A9/
nia7aT88EZCjgrxnP5cttdIvysN2M3tDpuaUHsKfq4EgMD9eZL4Wqes6SCigsXjuNmdpbWLXlqaf
W2h7CjYiEuVTXnSrQZ/U3qYdoSSOh+FVBxvEkjsnOuuc9AoSqHF6FeVDDMKC8fUk5QJ9yVd5O6Vv
3TfW9La30rw+b3hjvNVbzCn4TuNJq/llM5wfO7weHZCCA72ChFju5SyvY/Ozw7iNyOaoKcO2AoVg
meyzG/YICWiTjSzxFDWCnuwKufLgJuQXtdwhekEIBY1AinGpW3g4KlwVIVAsyftKw+cjY7N4Jn3D
pneLufO9Orlnye8ewF+isA2W4MeToYtT/yjMPcj92Fpd0zoxQc8LX2rQ54ArKArsSGxNpqfhO5Aw
ic7Doa14DKihNQH62ezw7iaCQINMLk42VgvuUnTVfkWNOv6/HJyhQcnqm4nWavNRChDQARv76yyY
gyT5VFiP74Fw6z3QG9fi8g3ogb2iYbjNuORV0G9pRbRFvWB2kyESZnwpjN0hRmWeGboR5ub2Zg2A
R5lQ6BIeKy3DObQEKbAxpC+KSTvJivBGoBJUQj6Kvz2UJ/E3Ftb7h/NeW5us3tXxXa/7HXThzXpu
Sx9l+zBeaRg4csxHDjdutXOtkz30JaZOTYo0ZmO+LCTJm+SNb+u7wVw91/p8PxFTv1zrvE0odDt+
a2L3tWz4ZQzBolzHLodLYJ9+QfLWAPbyb7gT1ZWf1/E9+nP5+yJyFeWLpEiyP6lq9hJDLahoGjpf
08srCJNglg6xLgmG/dbjnXRjBRVyzkt3Nke92ota38O3+XHKWMtKty7zF3OZA9aceQhc3vfNwH6C
zRghH0i3dfnD7BdhA94pkvx6OIF1t6fDgIQ6e6fZEdO4CXT1kq/lUTQvk/d0H6EaYnKBGJTQgv2r
Uts4pz+4fHSGguCKYYdNBspY29MOlvOgTr+cuPWdn7CQcnV5ZvbBomSB/J/NkgleuI1p3haeNX0D
cEUPU2eddbC9Jf04x7MAZr0wMmVErU/sN/JXAQYmwlwE00RpHofpEzTa0vRWp6o+L7T2z3/3WPqV
Lq7VO+XGq6Y6FHDSx5AekWy6ZtO9YqS4Q7O6aCPGIeZTnFGe4whmZTdGovZnOqFpm/8VJK0iP9UY
wtSV88vGtD665q4pUy9xDGxxRAvTeNjFNWsCW+1RejMERvJ/59CDb3X56vVGeS60XuTlEMbbdHwc
Z+ewcYRchrcrE/w+eM446lPRzWb17sxcPP7ZED5+dHd9ewoyFrDeg3xoq/KgCty9qaHGcTfFHNSK
aKBqdyAX7WADBMwabetZPbH4+5/XuEhwC7s2wbvDb707pqilIDa4KEpiF2sg+++HrUH8eH8Po/Xd
oOx8LchwPZCxVaV/c08olB29tAoI4hF8h/rYp1Ky+GBq+VoBQt6f8gvCmFak2rp9nTblF3/CfWDH
ecO3jwbNGkQSSOPBH/RDTjaylBaqxhpM1WGprRMVzHROdIwXCxK3A+9y6qRdywVLLvqPwqElI+0M
T9gVxe8OXHeOPo0slAXuPu1wSx7YX5/OmPZ3caAC3o6tvQWc6Enl0sTXzizVw//nASGg4ZXyQxDt
Ml8WKwxaH83BxsrSbylWy9pqAgOOZaEBsw9m6/3J/XL9f63N+agW1ZDr76SBJGHprSZq6aMQnPAK
oKmP1hfqaxRZbXMrC9IUUFDdH6FOLGrX20sZyo0DS7LXIrYQFmN4YI/1KwTf5SXiz71aP5DSZiWx
Wg4Oh4My1r7GXuj+kSX5fNahG2nTtFuoKROVB0uxI4ugHGh4MbR1gc87lqG/8mAX9Gg0ZKXB5XUS
+y0IAwOn2AD8lysii3fo6A2K1gW5zwfcJuwLxl3IdkGSK9Rmyn9lQyp24XVqiNhzEvFtJ77YCLzc
2wdx6GFYqqeZOqzlksunwEmlClthhLD/tVQPz5IEOMA+bGZ6IKmieeEndKjjK2HtI4sOk0gWOhIB
HJP4ES1ejcDJeYlgxvioUOes64cZA4VvZeY45wM06OG2Of5E4Fcx2zdIjbHCx17CH2f+7H+ZKVhS
eo7+EEArwkzCLJ8zG8YBKtjYAQxQWfOmGW/nKegVQ1PT3iclG+RoiMJ9nEua+5ia61jAmb3lM0Zr
2opLfrYCHZLvtB/3TLDpJqS+eYvzrckGzQ77/XGC8NOTf6XjgQlaFc93bmYEQrkwpvQ8oFqvE9tA
wVRvMB+P97I4bK4bJg/SQ0RMYVhJA0C63NrR9Sk0UsJnin9BRc4GaK1lPKHl8bj5vsywp+xmHebJ
uk8X65IXQMIE8eKPO+gDAxS9H5eNYMGXY8tMQ8opYtcNmVlmW06LWpyemGEFc9WOSjNIQMzKwHdw
fmM00VIMjD/hJTzxfwAcAzNNF+Xh4fphMZKnmqGcpGPQaebTiKhUIAQQphMOrRrCj+cctOZBemV3
n5vnbwOQ3cj031LZKszvbH41N0mJOW0VJ4YeK9zHTCT8nO/4k+n9oTlV0KjEh6iqmAIsXsCorY5C
J//ko3DsoJ/RErQwBK5GVHONIgpFXilZdsTNqGDQKkxlQwq4FEWyB/7TmoZafzeU9MyTPPUCcQNc
HeO0Lw9CPAwE3JFx0gtM31H0RFlO8cra+uDbYbe9sNlktytZPy7/8ehIX9H0nLpfXgXTDbgEfkQg
mhhpvof4RaUpeEnarNrKIjj/i5cgtkPSHr2r0HprojtqcPNJOGbwYFq+1I/tc5atdwcFXExSwGYs
Ow1uwj1m/FaORe9h6H5nfcw3Ew6WtQwFddLocJVADoYQ5ex8NFIlLsPhXhk6x7WmzsIobuY+Fiwc
0phOrgqtN3dD7Np0xMiXAIgv5rbVnKrOtDEdQ3GYn5urjmV4ZnFz896TDZg8LsQMnaqkZi6EPHD1
iJlSdLBCLxvpxczI7yeE/8OjCJAZ2eSOqFikJu6gp+tUsqotgzyH/4evwpTEHMmOmWta6j513vns
AkEOmQCOr///eBKmUiroztHuOvwA8wesVFqaxDrjbX1T0/dOfjs4/BxLbQVlg3H9/ZARqhWo0dBT
axHqtLoxdWUyok2Ipv3Yjt2EdQ5+y8FqLPqYGLH72ot5ahy0zxIPQP7dTrOIXd8WPSvZVnKlrTBL
XoAJDGiIVwaOb2SsMKzpfYWoVFYa8flptz6U97jZfnt0o4kK2PnQr4fwaDEkilp2kgqH/lH+JA2O
t0lcbc+mJp1YSAhTZEgZT5DUDJbuceem+CyncSHDWsFM8MkfYzUoeAF1V+27k0dc0nk+jACLSGZ3
GVVlG1mdP0yuxK1Zkqb03SXyk3CPHy+PvwBnJZa/8PbeIcDn4EAFiUWlxgThFaNmjdcvAwOeVC/8
NtFZ8sY7bIOdzSPOlCS4APKW2WA1v2rPVqeDYg/trFBhmLI04Kz+h6Pn4tBYqxfOrBwcN7poTh1y
DOcrXxdBdbSwdL0cyHCLyX3zNCmGzEpDmTvjJBCWR14n7nl5qhR4gKrfE/MmvcT8QHsBtz/cGz73
pJ4MntRvRcJFIWlM0jHBVEOQLbTgnoNAypKVAVcfnfU1HeLRX4v16vISTeTH3ihhmMqtyQNjvK7P
xwznj45asyoR08m2gYwkReq0D+FaNWC6x+DK69SqE29x2oOZgGlzCmrWm63pwclXosJ/ghal9IaR
QORUnrzFwut/8wLdLyeGk2HvFwsr8TWkcjCVflRCcQbhbk7GQI3/Z+UX7V4I+NK7QDVXXV+Py4r1
VayN1Im7CRsi4cFdcxn+KNCfPtWJSmJlrjThrAUhxMC6l90/d5KBviLqdAOzTn2HegWsUFSPQusd
SPxqLY3chsEtOCT5SEXMOJbHUNm0nqymgq8GoIw0o3v4wp3Ngzx7AF8/pfL+xd2Kjf/A/cIiYIZG
IkRsQp0BLG6rNwBqKiEHEo/HY/xX6q1RZng2iptsFfiaLHKpZocEIzUnIKdwANFPnoPqEr47jFTX
fSpO7CT081SnYUNqkyQvUQc0d22xThxGeavrzOtje9be5Pszc81uXSLGXK2niQkI319LPN2S0yqu
F1qIofR3GkXEcZhX/AaeVNHwb2wakUnqgiU+PmluSmFfIisl1arZaqzA+/1+fl+fLIGFkjAKgqno
jjm6Xwd4wCdfU8ZbV/XZRN6nJXchbFgr9WCZOUk0dDoXkfJpzi/XM7w2DW9C1pZiGLvsyTRtg0da
O3nEE60/VsUHOMtfotn/il8OkJd0FzVDPbSJCoXoHbJTMQpq2KSHnBvYlzZfbsCZKEy6HkH/vV5+
zU/+e11xifzd7YWM9skzrQmixvOTFqTQpmi1pPC11R8+Pclk4rfRLb96J/7BzDcJ1coVARDJcY76
EyH+iTNyEyQ3q+6na+ZSiWdjNefunWATxqUvFqSpVn7cWhMmVzKK8A0qprKyT1MVUbw0l6CQVds8
37woX7w0/8mSs+aj/lDM3vVDDFqtZQywji30byfuGbtxf/9zDpkvi4ZQ5/KQo27pDSGvKfYz8qsh
6ZYsC5G/HhsKxocBDuGye0cfiG2gjJgRiFHGFw8Cwik8CcBUlDFgas7GxwZLi9ufKVz6ZtzGhGWU
6EEGuTf7ToP3tBuvmx0qjyczFC3xXlsxB0fPrt18cUO4oTMx0jba1GtOVIG/JrNoAw7BGE3266qM
jvVOk4g3qh/UcyahCc8g8LuGbwPP8974vMC/e05z6dqB6PcBUjGFqrw4BU+jkUWJPX1KkAmU9Vxb
MWAsVmi7Pn40HtzhachF75T/QUnnyb8ufdBz5XWoJxKPgi6QVemI6h+ImUBkPNKgmECL8yMQO/GB
AXcxRilJskHnqU6wKXND47nubTk5tkFpGJ90z3/kEwJ4kzra5UOkx9t9E2FciE4HtBh7NGMzRHeG
qAygc70qI6Wm1NofL1B6yYarg08DWOgo8fYXyuJHoAmaVXq3q6uZv1dkU4IA4L9abhl0HZWBnmig
7NzKkJIxtaAteKL5FoKO90OCQunnc/71Z2B1hhriefmLi9jsOZwaq8Lnn7hmKlqzKcdPN66zf50w
4Bb4xX80Z1aFCg7q2Kk0gP644UhA8SZEIca2GKxlQWAIOGQAEkp2jIedirCDDWWOj8FF3PeWltii
O7OTiCWp6SRA4v+es4MlqysonWTNk5aqpShB7mR9IzpgAIluvLHK82ruyltY2lj908e+Tya6ilZb
8Us2QYLPyjLCkk2rGz1177D8KNZ8hEjcZZYEkib8pY8QQi1jbm0Js0a+JiJ7WQEtw0n5pUai18yD
I21xR6Uq/14uoUTd3EQ+oQz691JgEZ+oQBZclLgmTL4dC3R/qvtrHKsbdUOIjLyKGmBeJAvrWEE1
r8C+r1Z9miyt7tZn3Ctu5QCs8dDXpGU/AEKRY/cIiKhseptXjbs4DFMBNmlagKRDzOzXhyUdPYrI
40U+tAXSWr54j2BFWcAOWJQf1qRJ20Fv+hJ/c3P/2W7b5MIgdgJjZYJUdv+jesPNB0S/+hCrVBz6
hzC2ouSk31QZMcnXcsTX+P/XsrfdO2oEUyI8YBriOkP6TWFeo3zXIeBUKwOKGRrjfcfhG9iLDYvR
5P7v1di/DrImViX9zEv4VrPRRNvcKL6hLo/Ai1D69HTyiuTFVm432bz3Rgbw+8LhzdEsP2FIXKB/
QMGNV0UHbjpNHaIunrAD+7ueLVR0YIiXTCcrEsOa7BhQc4ADAFH7OR2It9XwOJJVBV0+VpsZTwG7
P7EupGGMsyXeQH7zGjVn77uIQelFAlvt70WpYgdiy1f7UEf5FhOCv4a7N5mnH9yvrtDwlXJCRF3M
Ga6MpGBi6gKd3U/uvsi16Im/4C1bcwRN4pFy8Dnh3PZRYcUk4QaKuxPa/HhgSceyR4WyLxDYBh4/
cHrvVGTfg3y2eGd9b4eIw9wt5mBX5YOLd/1h5C1teprmNgQOAJWMrw7Z8XtFVKAQu98bkz3bW9Ep
7j6CpHTnMJ59wSv3ugy2453J/BkKPQhzBqyBC/1zoct4XprE6+9eJwjYy9Ddh4IbB4dii8pWzfMJ
z5k5N4/4ac4SwbQqD3v+ahwhjeqL6tfk4SS7eM0+/ZcBn8gZDsE8HD6byrnZBtOOI5QiGLZPAoz1
WJ+dd1GQRs4ZAXspzSgBV/NLQqgvcz5gA6Lt32Xi76xkPev423H2oimRCGoNiGQNmlGbnoyHQx8M
6qzqu4oqBDROF9deo6EyB5npBtyn27788rThl1DcbSJFaiOdmzW23qjDtNNI+yq/hV8VtmakkQe9
eQ9k6xMmyRJXu3mWUSm6nlPA705HJm3U2NvPSe3CmxFB6t6oirjyv5jJeh69YiVRhS/wfrz7LgRq
tVz8XQoVurj/JC6yFie2NFQGmUI94hkU3OydJQFbbTh0V24gBoXoHueT8/fnyTb3NsDhFFU+kh/M
L9j7az4qjXwou0GHbdgXOok+2atCsiw8LbdUzm4PaLGGb4WtU3wLXXSujTnKfRVS5dLL4/jqmjZa
ojZ3KC7ohgcPtiL72dHDVCeUS/TFlPBS4tSk7O5e/2TNi9dbzCkrF2sE/h5cYql5FdmdAlNoEV9w
zUPv/bjcehwN3usdk0NEbbETtveeWnl1O4sFpVBMq/PZGVV9j5zF021fIh59/2a3pYizf3eAuhfV
gLsHEe3Txw8F3UDpDr2Eouvxh5gkSGFTVABaoC7+ZGN53pVHlyiyCJ87KrmogKN4E/6xkN1x7/6w
3zcyS5/xh1FL2JQ5f2ZmQj3FOVhmDKZDPsROAKvSqoXCHM7KYSxC6XIWgFyMURG18RbA9+nmFyQK
F+aIQm2O+9Z2y+uKzaIRhrzaDot/EWuhoXsUaJYpy0vZG+k6nJR0peVPeACh8PHkvY0sGEpzgEna
c0BgWh8nfLScTBaBVJ6N3qxLFHIbjs3e3Tfu00QZ4lP2b4rs3CGBH/lEeQeIzytBIKPwmmG0xMHr
oBFVdGhuwkChkafNPUNZe7oepVOacla78uWT+UIbnnZUl2uudPCMP5z113waoj+5+zUYUAqZl2Dm
qdqu4ll3EBFTKzaUBdEmZ1dCqcnzbMgWqrdN3X8pZmxpL+53FHpI+UBOdiFWEDixmjUK/VXok5UI
LAw4tAYHcnTqP6LJr7eHcfqRUh2SWAw3TRczwdE/b0ExzZqasaxBf1xgGXEAyViHQ4UekPdOJIth
VOHJiWEHwSk+LAg75v6AW/2BVMvzGPJkiVFlbhA8dPVA31bmXChnNWzNhkM6WwF0ncwYx8glq+Eb
8/2/zGLHwgJALlWCIEOjSmWfINE2UaF9e3b4JoTlJu6VBzrGsprQv921N2nx5DVfdTAe4gVhzPQv
Rbu/pC+rnpN4XM89s+jyuvbJbZ1G1NV+7GGmcKK2axRIm7qi1b2VDe5yCb9dk0sDAiJRine3+NC7
LH0d2x/JvKgNGGOA/Flx6prJjFPCJ7poU48tEXK4iLvXzoPN1/NANDpfZkXyEj9cGJufuIM53reH
wAqgtlnFIfqKlxVGQNtjBn44qnKJg30bQgN8dreID5bQ3fH4j7uRL9+lqodlBKHvR1s7+/sQx6dl
dvcvjGGMIaN5FgLzaUSgC0IPRbrF7W4j67C8U5T5v20k1Quu+JN6D1uinYtUg2g9mE3NXD8Rse+3
pXLeAHNcQxS065PRvJ5LqHfvAj1vUZboGEwwfFZ0N+aejhYLqQpLpV5rwBwDkwjTVkg/MkWdIaQL
d92B272wA8U/5yu3yGIN2gjCMItFoeDwKgod+ofqgsr5AnHf0RzXuM7ZJXIVcgKVF6wlCLHAEkx7
4whaoVuMJfAn4vhfSDX3Um2iq1EvPDXvntkFV0PEvR8v19yMdIlHAAwoWu2hLYokAFfhAJfZw6+A
eJhOK0hCfhMC2GkeiIuca77UTtvqHj0vhQaqvZRV6jlMLxe4nweG55VBJaaSOmLPL8Yf1kWxh3qy
0Z2zs2oRPXoublurJaxfFjLrkhpuwdLHxU41aBuuijAYoKKVtqAuFvFNZ6x1vzS1el3vCai0mpBW
41eYl950Nu+PmJDw14c97b/GsVth/gGxLVoVRGO/uFK9b/36zRGmkStK/TSN0TXlC9A/MNvTTLJo
9YARuLdo65ZzOHl6oGu82NaxvpYCvK/6/1v7LRiFrG39dA6R4Xmzm5KuaVyQshgTbQaArua6fPh8
EDqonPn5QI4e0jaAYWejq/jrSD7bhNJMID6i5ygVb6P/I4g8guwlsewiAVEyDjUQJpqp/COHJEb7
cdsNZoDbkx5EdnW5ZVe7IjL6Di1A3XbiG4Q6RR1oUf45FGptyFY8QBocX0Cw6wsopadIjKuImhuD
SE2RjMt+g5vBV/VhlvTwppskYCuzgo2QObKZkllSnzyDJjqPxB3u1N3gNhtN5G2gMb2DFrZkGJWs
EWj9AO8OsycBHatw2Xx+sspod0D+zS56y0vJe+APoGooTCH42439bV6j9OURCbLiPM3D3940FQKs
kgb+nlDIS4TFQsqXILM9t4NpeRT02KE17ZYGZtRBbgqfMxE68cVZwwTzFCCF6LGNE1Fq2pmqMWp8
xY22zTxlP5Xjw+iO2cvgzXEL5XiSLNYWoxJsJ4Zj1kwaw5N4QbEsrbYVwEo8vCmwCXnLqAzNSsET
ZPXoj0t+F4OBuTnbcmajjg8BXmEGf5q4XdVl6vRCiQ97pyMpFvNaDjlLo9M3tOj7M3DgZQfZsHiL
YP8ai3wo6lURnxcPma6/eaf2JH+fJXhlPQjTKiHy8G2LFWGdy1O1Wj7tTxRo7Lfbnd0bKuWcixvd
fMjuNTbfhjs7Q+bTJ/EbX5d6VubaIXHl7W/vWTB9+tkcudOplyw5KDmV7gjJQ0KkUw/WXQPqgITu
EJp2ysUC8256oyAqPABjd/a69pQOdJgLXekTYTQXY6Yhny2lfpU5FNYyQJAKKPjaKtQgCn0kZN6q
M35rwilaHOaqC4iIwR1eAdTSSQXf6W2kiszth16HYJyndi1oewlcMizYnYiL+zMPZSvstwop+28t
SCpNJDiNdhbwF4jd6thzwwm68rrIo4GqQameCvXZ2xZ2Nbfym9+oUQHt8I7kG+A8VCF7lkuzTEGw
vdELfV3j6o851CvnR8ZshnTV3T3n4BuLb3ihS05/hlaYNEiOwOnEmHmMjgslTuOlcb0opa0h4ZwJ
luYEqioi9ZBNsPso/HHfDHUvoISY4qRh1UZAxe7R0CX7DgMUeOiVBQ4chU33J9mEgyHlMc1K8tvC
OZJ3yQqOZxlZHeaE6eOUJNKq6GWCcv/dkmGmtKywWWt3KDuBJhTSkIPMcfRpNHxdht1QpJQaSKdz
MLNVbmiypEZGkEy+blft6vAgJObPI+o9USBL/yP6UKN96pkGFMRzb9gdtPeocbTZWdEIc9f3x00X
BvX5YQPYkrSgt/BOyYc+ppnfuJUuqAIBtdeb6Yob0soOy0QtC82kVPmiaxe6A7bboxYCmDr1I/ik
E8OXhjsP8bMmPAMJqKs5wnDK07C0f1fuXfNSe/CxbSfyBmoa+FvmYmk15z2RPYDyeZh9eaLGC6ws
3rs0AYw5XG5tG9F1mK3FpdWPyk0zdefRztmTDtrzKYOMvJ9vrXqYtza8Kgzbi4zzn073JM9mJlyQ
pHBzqyhQVe1/2weLdsPPkI9MuRhpLdnVsQ5qYKxzbKO3vxqLqT934KLZApY97XN3paymyxO5wCQv
+8BsxBWwEAE6ygRfIehREFggUXMGfU9Hfq/ZH0fsgYCRUFUaPhgt7bB62elSXNO7KiKzMfNtbRSo
izxPHZ+4LBWskZtG+OakE01LwHbso+R/tdTXvFfju4DgmVK8RoIf7/iUP8e3ya2tVM868mxU9Omy
7LajdaefmvaUkRY3RjtJ+i7YULohmkQtoiCpvUMVWvZCoYIz4tmkm61DdJOMQV1t9Sz8axq2Crc1
O8UbCcG0/iNOt6ZCzXOCTvI4HQPLMi2ZDRqv7fLYlHqVItoOU7vJwPBBw+EINFhPaiz4BmO3f2rI
En48ztxEnsFcW5hSjXC5x8bdVvmUi/dbrSOOnV4y5mOZrKJ6UR3wrt9k4oKrE1nqT8+R2/TogSfp
VUof+3e9biQHAoMayUbv5nqBQOKmvzYKsfNpsNBrDe1TRXBufZ+/NALLM65p7f2oPP7xwkQ5ozuY
5WcES+3PN/HjXic22gRkKSl0Kas/NCKZxNVhjKjX3E+adDIuqtm1U6yFAHnrL/JWj5zTas5ZwgBU
rfCCcvbohMwbW31/JA8Op6xqBLf6tt4/zx57Yn7veBM4ELvUoCZeKoiDkqD41LWX83yjBvDA6Cqj
VHpmCkDcG4vlFXxCml6Fu3i9sQPx2lCWZZvMqvLyZXODUMBgGf2ZNxhhktM4mU/ffMkWVn+7uZWQ
fm+0CLTUxVWOCnZe9UxfQHG3PxNge5J7LRNjU3wJb9yJjavxKTlYMATBicqgGIn8Wcnq6oHnrOiZ
5jZHgpLAgB+mcpctx1v4VFcAgWe6XJmx64c/pARfzNhPUsqc/CxpKEhgJopQccXYxV1RvcHQkVte
Xn6XGZgvrbaFcX+Pik2ulM2W2ShyXOtDMv3XqI7GaPvi8Im5y0eLyBp0GxZaxeoEnLXzGAQyVAsm
w8dngBoiPRmzOSaijl37ImtafRMJ+I/Y7ysdMU5TRlV0IDg4xc5ci+lMMXzD/wzbdVY8c/U5dNj3
fOLwphXJNv6GmLhiHLrFUJOumUGqYFKb8vsj1Li4u5JdO4v8Fonny47EON5lCwbal6hb49d7OiD8
xKmrwNm2Of849udFC+mXbi6i/HOgRHcF7MAYw58BpZVE2TLYZS2iffUxnZyr3n+q6KwFkJce+muJ
kw+h/qZdu3B3FUYDBoEnbJ0F0/TQrorXKHNmobyoH0vsEDULJ4msHUdq2Fh9XoP49NeNHPveE9zr
o7tKtEKT6B5X+ZoZrkar07CfY0RAZzlnLPFoe+QBMLEJK92qDYSKRpKE5Egt9CxEqx/7Ml08rsd9
zMFWyUgor+aSOlvT/hWGouBNQCl6tVvoiiInUb3YI0zHX3tu7V4bovWz+LU5wyPhdPpELsoR+3tn
UYNke7Qh/hJVYREBqfJUBDvCVHpNo/ZLz4fBHdZFOZWIaa+cjAhOuZCssncXcu0UgKb1v7QpbfvL
NyyIHmWviyRU3EzdFZi9Xr6l0oVs6cpFAArwhpVoUh/rKmgWaAGABoF9VxBNhYLiw8oTCf+YDwOf
LXyV1pnKSFlCIeSw8fcdS1UYolo2W1JXJHjlztreXQYxd+zrrGTafGuYMdnn1igTz2hFxYv9Fedc
fnsyTGQ3IOwB+C+dmbUYLTPrBtGfBJUsb6dKQC4Bra57s4EQ+q1RTzku8ySZJ6cFgqoHLLqkFq78
gnoS+DvCUxcQAbxUWxNnFMDwD6X3QkPmHLUUFYordFv4ryNTga/9c8G5RfJLxp3EEDQscImlBnY7
lHLJaGAioMZz0ZnafLoBN6V5UmkzYbEpQxnwl4nAWQpthAfgTB1UOvbraOGW1uwTOSbEMhY/SDcT
wCNihXXcmxzOMH9j0t3SdNQZW3pbdP4ldYAY3AsOlTFDg4XtogYxAi1KvcF6tkI8xeMClUlIfOjs
6i9J5SVH5G+CgSwDqR6xypfdzRhEVKMHB8dMaY8yLkOVWoDNCIJKi2SU86b1AvAjXuDd0fCBEjTW
n4krJT8c36GQf5wguEz7b+BGg7JgwttqXJ/T/ukNM4t+t9L/seXHkOMvJ7fkZv+Jw6bjB7B1zlb/
Ncyp9ZY0Yt8GYphjKRD88vNaWZgtPmUIlIWaTTWucQ7y6lAMV36WBIVjPx/KknavL4ULLNoBGT2W
rxSq7suQxJcnxXDa5XhrblZ8Mm77lynevJz+zb+Of2kDUuFHR/hOzbpXw9HaC/jygrC5vC+rWise
EfESAj947fkjdpwTasRLjQrKJaPRecIhXwcQnktvDahC4rTVmOGB29BfaTbVAQh53uMrKuL1OGYl
XYyq+mvr4vA9nQ+HBJ+Z3e+LNrA44zvh9hmwlxV6kaC7SItxA6ZujaM4aUxz62CbX8g+C2URbm2e
eGTn1HILZ+G2IOYgrG+gStJG5WkctfWZnD39k3dEDgNUEqwpsX7WJWoXZ0qWejM6YR2K2KFdJBlK
M4jarDtWHC5/PWkRNgH9Fkjg/KH5QBX7cdRlZCUubVRuFDHzRugkoFC3hwQs2WbnHjihl3+2axrE
qynjGLun1hNv02CuaCxw/ELbua+vzNGZlLH9F3SFyhCFaX5eaxEn7umvudlJb+3Ase5J798wN6Q2
fusKRSzTWYVp9lUOtv/qbr7J6uj3nsIxkEquCBSqOGO7BXovzS63gz1MLTUbAfWE9/EirvNpqIz8
osvzwX2HbWMWBbv9QmjHNzyCgZKxa75+KYtUSt/Vea3bu555ucdLWsmwNo/to+zA7AvXC3VIQnhh
YTa8bqjXpZMgKGsFEVejYHMFgxT2HfqFZ6K98FDqbxTBXn7CvVQ86YaiRDRtssPEakvkrOJP4A0u
i5cl713iDRdrbscqvS95YjM/f7TuwPe0UQCJNkaUoPXhZxK7yw0a+pJ8XwTKpUQwUAvB+/2JTXlL
asFFx0O+EXxgcUkOw2yH16NSIt2LX5hXCRlLWjKALDY88xQhmr/av+XTz/fvgdDwFhoK2aS5gR9y
epkm/jv3Ol3qdmoSwlx4athHQ4+pttzUsnkt1fubTPQvjigOAn4zU2wVsT5JD9SARQFiTrI0P8+u
1aYNkRS7Jr9bE5YYl1R45rsNdsBLMGjTtFGgal+abA8serJy8Umztgdieg4x7M++5hj6weVyYhwM
B88Na+7pfVkAqlnxihVu8DvubSqSR1X8avYmT54AIV0XUUu/GlqglZcfRBDbs9Ul6V13ceYI2PO9
6j9ec9XlTpUbiel72i24paW+MEaR+V2jxT4G5ome0ZxOI61u1Ec8Z28bDresxo0470IZth/C3BrA
o38o1fvP57u2Oc0PJYhpdS3vRNE8XSNpeVsPDCyQy52rw/W05uGCMk6ppalg+O6tcaR2PK4UBr2k
AsFaWgEBtbwG4Z/VNEDxh7LyLtlTSNYMsvnEji0b7PaBqpD5r5Yja/SqUs6YTdDcjP60gmIg8drr
1mOP1DwEnsYVeuh+Szt1B4M/NkL0wiGmG6HcrD1ixnWIY3bmWKhXmcDD/5h07XIgJoIgqptnQ2Fg
wPeKdRrdPryJG2evnfEeuXoZcdtu+ZoSS0qy9+z8Qxj1rm4PakJ4ECR72QSEjH0Y1ykyU2LzqFCo
rR0bS+x5Ibm6kz2NC7bu1AA0av1G0h/gAGe8Fu6JorHvi6IdX0cWU9EIxWYCF8ZYPl1hPIGdHiFK
Xu6Q5jvPeKLw02vPXMOmMeLA8568HqQOjaxaiNzNkmG2XUMUUD8dhHtS6AREA9AKWMcZRT500Wy2
pux+yNVrs3P6jH+166YD68XjnVM61ur5K4FyL7t/d1zPCTNJL8dOamBZdCy7zgINIrSM7A/6VKGr
K4PZA9787K57v/FISUvBWdpa3C8qwLg1TVP9X+qC6gH3YBToVUNSw9ypWNLy7htd5ecL2zkqHz1f
FpXYbJTrxAN6WW3h3shZCjvOOxmCb16Xga0X8ud6Bqx155rPGMq0SoWXQh1JWkOgW0pmfCUaFCIV
bMw5/8oBxydsDhZR7+D5c7wv0jVitZ35hcinkJt44SkMUrVEXimupkq3Be0NVdwi6Fmeg0Ll30ab
ozcnYnOmxD3JlvNNb9jmukbFZgBrMNc/xyisDRdVq5bV/uuAY6x9BKQWDsWZtjIFtGY+Kgz8/xZ/
iGuyy43f1G15fyYDVg7vSKILp7CXRs7ByZ2qlFFIygpJGg6RGJUIlwpNjlS+aTEroz/0f6kgd/y/
LT8KqQFCeA5Qw/M7xFPJJnkCXC1AQEsln9skT9hYDhBuDpBLr6f08gcPRuMwHx6u2zPsiKgkdapu
D6QEZSLdhIVWoql7PpLTQsJ0S6xI9xmO0WINvRdRwWzyurW8UTiz6lP0vjENMEwLWekk1FfBhQV7
q3gKPMt4qVJGndO52Zpi6oFPB28MzlhdcMWe9w4/9mQ+wWaziUHvlkTb6TGzXc3UZ9ZFtuSWC37x
93gGIBi0NPVLJUZzTW0U5Ze1s/gR8MyhxoFxzdcDLophFxWCbKVrUY1tBZiHCvYLj/9Kva294vwJ
KvobCqzl8sNF7VVaqUPeb0WbA7Brbt0OhSRYDsZ7j3iQa3tKTftJXJZw2UKm/yivP5dHtTo3G5Z1
CiFNPDb7Sdi/zFP8Yxq5Ek3Z+nvsS1UFryQ0Rh3pi8mPBCzRZsizkCYJ5tkPDWEbbKswZKt6fnaj
kL9czaC2drrn1Afly01/0yDinxa6H38TiFYhULPmJLcS2TFyOhgDvg25pGQvVJDoW/0ukh0gemF+
Mn9AA2taHmI2HqVlb5S95GrzLGpKD1h/odrDwpcD1Rvb3uaWJTNxblKGs88Dq+2X/Woj8dRqt+al
YqU8m15YQi+gj4a5uNwTrXX1n0jEYFDwi37AltozarrHotmcNNeI1j1g/GhgGI4EafMFfZKcyf6H
3LY3xXYRI73L2K6trxwXZEZwJPwmqdnhEgutq97bz0KMAMUjhojuRCmv5Zc/aYh0r6MMhrNWIgOp
BKIvVsVJHtaqkWj4FV0xKunbYleirE9Ea2drrzs5YSAqehIDdQ+VFOpuCca2hyzBk2CqNRlQ/zLD
Tqy3uAkaLAPFugFRbpAKcnlO3V4/sVdb7JGAgtzMY9JywSOqfS8kNdm1aVAJ3/jphBfyXj0ZUl92
y5UErHyXo9hzLoBjUuORllRNepO5irQzs62tSFAnm9wbzazOItNIueSoYh4eCeoSAwhbBIX2Njnh
nmogrWKigOd7vMyGgFEoViFYwKnOy3KENPQgeQTgwcB+QAnLuv1Q8gOcL3YO7ivu+PrptDRzA3os
SFKVC3DoFzOXYcrxAW2UcQeLA7kTAYc0LOd2Y69tfZmMmYeeD7VtuIs6CUOaAyv/Qfnpm2RcKfYH
g7iH3kZPLz3wSn8Qq/xfwBw3MgApuytrQVNXAxesP/cKtOygZ2lzZBxPYRyNey6SgdSfordis9lH
52TAvkyFqM6/OEGjjIXQiys90OwSdz0Y4jyAO7WLxcQgROTnx7bcX59/yNFjVPqjwK58y1tbpdYA
uc7D5LXE9yfg9Rm/Ffb3OTd+q2d7trPepshhdMzj/NR1r9L+TrH4uRebn99Isdh34g8567LP2P7t
QVZ3lEpCbSZANYKV05AVuJsYSNcDx1pfYcGesGidm/jgscJFPc4JrEm32c+Mo+4/KjQZypBM8fgG
tKTvfJOEF0ZhZ8Z/IwNddcNHBiHEs8mqzyuBgxLzULm9tkik30+9Wvz/HyDEoh22s/QpfDOE9WLZ
HHhpOA5yNeD1TOPk9yLqLagF/a6fC7p8m3RIXwEmv+ZIQQeHVx4ltX1LdzjHpoTUJMDaO0fwuma1
3jADSpmyXB0vyZIyUQETNMsp8NUfAljKBOFdBYCmYswxtQIK0NNDcP1LkXbvdNR91krRrje8CjxJ
2lal9rJwDXbbNyHdK1FuRxJpxyrBGlnccdEBPzjWr0tLzq/FLjccuq5HBhmDKzanTm+dy5P75P+H
FvB//L5r9JsWXkdCm6kUN2uZdx29WvNvkLJGRlT0Tn0zy6qKnx2D2DN3GOF7l0iDJjK8f61LyKSC
6QB33/d1jDsafpdYBgDIJ0XivMxWvufMnXt3RdtqMW9uWuPflbNpJNh3BLfcmrGjtEKumKyuHXBo
/eS/WIvPWJhnP33nJigEk91t+QIk7jp+yiVlK6XxyolTUk4v/+VNNo2CPFTUGhf/U2ezlbGjTLRh
IrPh+v+hr1HkC4FLgjCxnt7czUOx1lf/S01vIdZef1OCjigN/cIhpWCxWeFhVwDZT1sTsqcXAP8D
b87XpS1CTXzRt0AW0wXRTNz2vXBvAiS8WXKR0TQ0hSrbBp6BU7QZD9ypI9xs8i702VXnJ8Hg2Y9U
CZ3BvM2xW7SO4McR0Gl53+m1QMA+ovGVmqIsCF9hvdtcXe64tA75RSUOxznga3VYwuX6PTPpbtGB
+9AVWpRIfwYckEQ4cK/9w2fMFJCU5d29rwCsb47FBKrtzOtmNYKVAa9J/CEmP1mAi+TLYDG5X3u+
Axq0D/TofPO3AP4WKi5V8KRxXL4fw7e75DkTVGhHmdOp7XC4ABw90IK1gwsa7ADHQCkYIk6+1dqE
hPFSjAYtjSghEs9H+s6+mOU43txisZtAO+pKudEwTpTEUB2YCPi/Z5RbsaU+OZzXgudjCep8ZWwG
CxrbvLdYXuJQiNpM1UalKiKbrcCERDD6WdQZfLeoO5f+B74CGpuPpYQkWvWBIQtCidN3ZTY8+w7D
2Azwzol0l2jbGBKVTsf/cca4W3URjwjRmSNNTaA5HptvqEuvE8v4u9OFXWUUJg/TjZj5xsVvHcfU
LySst0zhhOfDj3w0OO0MSjzFmerRIQVpjvzuFtnovdBAD3TIzS+wxON6+5bk1bSeyTHcS1nTvwmQ
SfOCs5Tkvs+gxb67ftGqOqBH+KdpRhqusPzKC3SI6cd/WRyDmgle+Sx8kJw5Z06qdRfr/ho5egpW
fFN1nM1iz/ICMTTxwFC0LQKK83J0fpfeRpQb4PUg0fDUipxjACcu3VUsiCz9ktMddvv0EmIQsvLq
re+1HTCPRNhyAjt3wEKaylLJiVS5jlUSJWV9gwL09f8cL8+XN6QDuOZFsGIiS5ctwPnZmAWsFaTu
UxfsJWMQ17VozSP5+3bD8bAA88szC9zqB6yqlFRuacYIs9hURPg253X950Rx3O8eaD1/A/h1y0us
SdIePLJ7FgCaFyM8UabR1AowG7TyJDp1UVWL8EV9Fu9d7yZDaVlwyAqcdQAJGbLs3YRkpXiiybZu
1BKJXlmyhHN8vyDNhfN7UF6AgupmU2TU6H3LFtQEkbwFq6byt6kLOJhc8l+nx67pU280D8ho306b
aV75Im+J0vknlvDxVIJdHgpyg1Jt0g5rDNjczzfTcWpPwhV49+LFE8QEeisyu3yCpfK9vU2H21Yd
BBPqXWNKgVI1gebp9i69LJx2kzx24xZ4TsV2O950hd58XefsezebHgsrCpk0JJ3/gPeYrRb8t6Yv
KZGdymiI1b2LaTlsMCZRNYnrrJTLRN6pnJs4soM4ZKMvg+LT37FmchH/0H+1fkuzbcZU4dtoya/Z
Ka8OigLLJKamhyLi7KfieCplC79mIj6LSm8DXHb/H1xLUHCaoYUSeaCFxLeUW3fvZD8KKvzN9tIY
BTD2lGIZzIOlhFkhs5bLNhaXVr0oLcfeUfwMS6lUd4d1Qi6KInUL5DmxQGJg8uSCfgvkHL2DUggP
JKh0diHCPbhQ7nH/0PPGVtNz9F0rzihPclWKcrHdroAIVcImnDeQgOmk+9myiDJ65WSOftpZTgoY
PICbM6PqDtJLLx00O/6fak3CU5NuW0mtNHtCsaWAryKkjYAVIgJUzl6cQvdbOafXIcLm8DhQWR9X
QHzB1aKIqpdavbk7n+29MPSBHu8rCYMzaNlW9Q9NO53nLJxmc3Ji6SeT1SkAzBZj4B9xB81BsHqD
rG1y0tmPhJkDM2MA/J/FJS4SjyQ7vpo0zpNku1fGZ06UIu2Xr7iXcL7aRPvdBuQlhR454sYuEr3C
ltL+HEZ7u21JxCBoTBgYxshsWKOMNOfS4RbspvJiB1HujiXFXKfCAHyE492uCnhhSXL7O+yaCl21
4m8qo3jM4Knsh6mIJdKRQjUmfwgZt0iOxQd/SA48ckg4aMsOGnx9FmfasOtJDpMgeJmfFpgjUyBl
4JT2bdVgbyGMdIDraMSDZkDr+rem/DFpSg034xAHLNDbCp9x5mkzoCOQSwyFgN1hyA2JkNyk7g6j
psg+pVG8rKNpmiFFuWcZyjPvti/aHzyUZlZs44vPo5yoj6viEfJVHcSvK9s6y20mHTXElUK8Wq9t
eSoxespfvgEXDJAzUseyF20bjlSaja/a8W+M4GJCXK75YIWhJS7BfkoHQ/lOUiqjssDkJ/kTfBYf
kjAoLIsl4pvEHD+f3Qndsw8po3osTMHHB7jXM/Pwpk5uVWWSkEmfQ+IWOUOqZIuYMbbQiNGKghye
zXD9tvL76Q1qnuPhTwrSz/zA4KcRNozrdj1udBqPGzTcmiAz2w1AVx1/aPN3qfM8rFWd+FudCGIp
G5HuiHFDZ1El8EpbsGNQasv0AvfAYy6iz7OpLZTetUs5wkMIuB/sQmpIW8jG/EjZrE0hYwhc1SlU
t9cFTD+/YbLd4eOEqWsa1NaSbQNRbtTtL3bq0Z9hFf3gAmiDqyuzSe7nMX542RYu/Gxj679hQky/
5mjjQLbq/fEmR/o1CJiD1wXxJpiRvONiF9N2zA+QBkkscG7ZeS2KcrJJVcbYUMncchFMkFYx8qFB
aWIt6o5r5qGO3Qb78Z5z9XLLe7/3+SoSLJBC9pB+0ucGb+aMZhtmGk1LNCdsbBmDAXnzMoutneIo
s4BaLyHm9GpQ9yKisLGPowodqZDRYevVd7u1SkqsBdtJ1jMCSKjInJ14ZvS6n+oq289GIpi+9Y8b
6LsNJQX9HFUs56/z7Mm6CN1C5AU2S8gLGSQ8TYtgjFbUB/fs9/aUeunZC01Sexro6N5ld+qtEdUW
yTMXjOFN9a7HjXblXvS9g5Ujg2p63Xgyc1TN//QnIijNiTWKsaq97znVHAwsXD7szRjhma4rDrU5
Cgk4Ltzu/YTqgHYB+jkwTsNPKLhnA3D1X7kO9jxrMUgTX0vTBgpGWJjJLUKc00K0D3lSYVFC+v8O
/wOL8EPgif/R0g/fmIwmKTVlXYVATbsHOpWzgjaS70B1GEj1Xa29mVMo/OIIoqo/IptYzGAUoDfe
ZW1Uh2l9kaAYG8RzuRI7xz+9brf0/ky5+VRf/M0tEblCGGNDwopvZWoMTrx492Wm0LjARP1rleqn
WhxhBrt4133iO5fYH0Pky/L/8EjLeUfQC09qnO+OiMItXRY6HSctoSRpx174fRII0TP7EK+rvuZD
GC7WXJ6jusF7VqoS+9p1pZmH+Q4k8X7RK0TQtStO2EcsXgEtgLOW9PZis0wHC3vDVLHqXHflMdKy
uYkKXCWkSqiwicpWz8xA10ewm9JomG6SIubSMQYfx2TF667BjcmnimCFYQaX3Xq9RcxrOwESjTQk
xSNiRivbGQDiIrhpaYEAt7j/l4UnFneCsU0+dKjTjamVtUYcPpia/pF8bULwqPnTKLahkjtVKxbK
Kh+1MKeLA9HhVdyrBz8y2iqcMBHVHFCzj9wD84Lj7bd/Kct6F2mUAZUGiS1Om0JHWY6I4ZWYvKZ3
aY2SBP0ujCLydTr6nS06lINdJwsEAB0yPIcGKvRrqAa1ShWLcuhDTrTFrSrcHKP1FAnH3sR7tO1t
oXS0bS8S/KmobEnVzC43RC79VAIHAeCOYM4DIVCGFiuHvvPMx3nKDviUpzgRbfBRft3sSNFXZ/bv
W2p4UZKsha9ithWROWw9V/6gUB2hnuFrq64KPKhD/JSrnHMMIhMzYgxsAfZf5+jMRHm4NL0VLF5K
Kh8hes3pP0YrJz1zxdBmfHgeT30vBgiuZBns0GLwemYKA1SvBxROFZCYcKBhpBhl6USMpi8y8YL+
4pIeruj0vBAVRt2TxkMwq+9mnyvf7VkRws2HzW7EnXEcNZ6li1O2zRl3M5PlyvBwMG5//Ns8bXKu
wxY+SWcNYGT8JFT0ot+Atg8EjJNEHwNArKywYdeflhKRXfe/kkQrJP5BnopwQnzrBTBccyAOoZHm
NndUpZatmI+/7V9fGlXVMxBhjYO51SfAAir9U0bQvxT7uI+9QqSVS8EHU6z4wmsoUYwINiNtJz1t
FCX1ofwwDGxj9oNJczg4om9g0F/gdpCt5QyFt/cjU/i2eaDtjaF8tMkaQIz89SM0Rlv6HimD9PUj
2ZKrZey1HJNKUI191PuqJkCNoVVbWQOYDEJ8bb2GR5wpTy8n82vZVelGp2VS5wTxe/KiS7vynQij
5QOfnJ8QkrKMXnKyrXH3I02pheNhvzmjWrQsA8J34aAuwqejuNNghCXoIxmytZerCw5pXowTXaej
zLZF4c0x9C02UZfYBnlxqKDN1m1V4Gi5aSMmNDvRSBSRIZex6uVdIiZYVd9ZBKNR7VJQdVDRmRF2
cvTEOfvmLLAAvZRAQZQ1OR+0KkHd2IJUdobU/cHdFh7AT4sx/ZUkeehS3eObhOK43mgSIYoLrHfE
ehvWIrKCHkRAYZX65IZC9vQLrmFak5Q3cpBuzMRIaGMi+5d2wQlhwjifvyD9d97NvCmgr37jI6s8
SXnV1ROZTi4xlkiNVg0ps+/BU46FlQGbxHGjYdn6F90hJSUQb9nxVTXutBVYU2aCEqsHqzZW0SAn
hJHumlhRUiE/Kf7DI+iIz6Gm2G+RE41bSgDI1ToQgqvvhJzPeurVeEuECQB7pCU6t3TTvfz4Fqp3
7eUh1E1VBAMhp0My7Ebu9+Yf8QyEEXoo5cDrYYwkdGq5zzXOTqwLy/rsFVynUPaB2LyKAV8PZdMF
na03Ut/QPx78JMAtEx/1DpdbfKCq/ijGaDXCxBrtlx3NEb3zOFv9nVHeYUDyFZP5OsCdU4ThcuIC
XftmftVLwQtD0FzeA32Ub3lzc97b8M53+UolK1Lop4Z1bw7B/l7OcBqzQEcs2ML5+xiWSIApgfn/
mNSpt8HgmuP33gSWXOb0rdt72bWa7D0IMCxcdfNPptk7e3GtfhfW/tRkB0lZGykKK9W7Ub6NCHlM
xkWemB6W0Z7dwDNJnXM8770rGpBas+ICuOwoD+nQYDLfYAgf4An0bNLo23FZZ/YK7hAscwhlarId
7U6Cfi4qPnDNmfVhNLRapZTrtvqYCifHLOJFRO1vrS+bEJwWViUSH7QBsBoz0e4KvAj7R1B7/iVi
p4GwSIOJZijp/Xm7OnTM1YnH5sip6wj7sZwZHmLALG0ofVfxQB/Va1QMrO9wretnyk45HZR3MVnf
7H1x/3uHvcCMkrNoqnChy1lLlGUBwBj6SQf6ODWD8C+krVC3brCtpyqjg7lY96faofqNS06TRhBT
DLwEXWOpl/YtqRJPvVvOZXYVYZxZTZPjRC//wSfAYozEORSDNDGkkCMwKLyswoHQkS3dKQgKYGNT
bMsyHDYYDeErIK4s1DFltlEIcF9bXrmRMobjVFZNiRH7pdvv+2vexGPU94kv81ddEz1qbhaCmYEU
Bo96eExvy6kRv2qpF4dfVbXivp6ZMQzk+dljbR4RshJJjGS442ejDijlJzppiy1kis+qLivFUPuv
/Zu78K9VSC+z4AH9ir2t8/sabzXVNowtgJyiy0gjsnidnaj7c6A79LQtn7CZsZVKt6tmeePC6TRO
PMcnySlTRFi4zCD+NFGLFMQ4QIS8yl9OD68DLbYE+oZogaF45g/UP/FPpv5ujhH7MvM3QAEG2Ua1
aTOeappM/bhVw0Fy4UYv20SEroNsY1n1wzMPB4S9oAenc6Si8tthAZj1dRxCZarLaTmDjRAgWQ0D
w3vW3ozXIMdpsAFJ5VtXOPA2KHI9fd5S4dRGfi928MDmn5uwzva07Mygy3DeXxk0XEe6ux89C3ww
Y6B8u0J7rgrb4t9HRWB74ms7ehxpkMbTsg8NiA6zfMdXQCYTDYC/jftYTEfPyHSItdg8CkyitGtm
VfOSMpKFe2vZhCfGZKxz6OwLrq0dPnGAdtc4fFIaeIAqIPbpVsRAhQxM7UTlXCucDVrFrHiSKmeN
zXIYOMm3aDd7gxO5IkaBxgcNWlUGwRPyuthsy0BLbxfgj87cK55jj78nMqggGP0b+NePLnucJn4B
FlyOEE8f/6aA7r4MKbUA2O89nKMOOs7FXLxAEH+tO9ra0dIAvxjywkO6DjufYdD1Vlr0/FNRLubU
rkI32wCzNo6VV2Y871Cjj34JhKsMjGP9d7glSgAaugK9BfboHCNHpVPQtp9oC0vPLY+sUTXBEkz7
0aOzYzF6+ieAawSfMZy47HooTmmho2nscH1qB1LzDHaZBHHRcbTUq2CT1bOjAtuNzcAEUev51hMc
gde4TKT4M7Au5hGorsoYIRryUyEBB/YmkiSlcmSKPpMgeasRPEXX1TyykGbC/4r3iwEJGPee2dcC
08aCjyqbdVCy1RNp5h36SJKwbm2seTKD/+uZgjVZHCRy8mRWBYMKnxtau16F7YzF/a6dLNQMoniV
VX+KpmyNj/9A6v55Q8gtiAsZdObo0stCuBvFAC8cUs622aF8sKyzjd4fvc5KrVWf5zO7VafD7dvy
nyDoFCnDfOH+TVRhpRp1Ve85JK2O4F5URVcIJrOn8kUqt7lDxJBTwzeQf86itU4uaMprZwLIOMKW
Q2c9gdXqdos44zS+d7VPnveNUq4p6YIe3TS/i+Mqp8os2UEEBjkHZe14MAFQs8MZSXpGqRvU3328
g8DtTIM6YJnUj5hVESwHYN6Ts2DU41GxU6TldYluo465tbnz51a8jrTgXyWMUDrd+IpKeS7EZWcl
Jj/XoV74bXJbrSXp8Wix8OT0Yj3nxoeMafNWH3y9U43aDZ6rdvkmGdwv7oVJMqjcYf5+ceimG4sl
uKheLLQpDtXIytrFjkNvNSqO3FawVVk+BtKeuA5K6l/9tT62EPPMmXTf9Mtr+BSoAUwF4bn0kYLV
SPXCVAxbrMwXo3WavrVuqj/LKCos4SmjNYXxIhtw3g1bGrT4un7isZo/ImI9r4SjmL0M4yeWsCQW
asJBCN4XBJHIP6te8MDDC7/v5PBBaeuGZDGPhelQH2HmkOcqTqGrzjiv/WO4FFTwnf52/mQpTMzF
1l0kPchn1ut0Vvhhg1c51WJbqgeH9skY2K4vpHRw3vjgiWDuXmtycP3U+kIYvbvFH2kwZrLbLSqj
jlB2wMCvvrQ4yCiwM0LSlHrI0h5ki4J6sfhSABxXYTHcymMQrckfmOS1OK2nnlSejo6yVO4+P1yO
gQetg17x6nwV+vybsWJX2omvr3fp0rfefUaSRyJmKwllVmZzxpLpJH9kPJXZPyUBvAQkV6xs0OJ8
PpO8Ro/iWVkx67gbUPRMqSg6eCbM1HwDxyAtYAvb0qNfWGl1PlM6SKIrvlSLS9EUmQLVKZ7vyI1m
RaHt0pUG32X8shwK+H0HJOzuUAm0CqRSWhyTtPphpF0HXwnEyPWaFVERDVKehLoTEUrMBmyIVjaK
1Eg5AkGxVOeauZANPSVQ6t2ps6JqUgSZ8Lj5q1YUwRyWUvTCAtkMdCJ5l/JFUAEsIHHMJhCMzhH9
Y7FiU9jFR1Ic4WGU5NkLCA4Kh+OYC60Pa9A1lieejlKR9ldGHA2UqJXeLyfmE9NJiaSDjvwLtSc4
9/+epE7yvKrCdpPUSq0X13jpVJbKFCz9+OSfunRA/1hgtBnZpgKHniSPJ+vk/LBHsrkdRdrvJh5b
sMcMFhST5FOjCkyEvQqPsRyXoQLqZfNetwgRplXDYYvWLGxP6UKcNPc2rYGsK2IzfCE3DWmhcmyG
4a3/W9/kf1VwAe5fTPkNz5/oZ3/182DZq2fXq11WjZJFfRFDdagAZldUIZSSSmll7ZWwIvu/f4yz
jvORRX/nGEeutJuC3cLoH9yTH+y3Tohm30hGPa/1c6u33CG3SHUARcP69TuTzq39yiIl8nZ26KxS
/QEB5V3ti21MpUEkuwDT9SJ4Oc1Ngl03FoyyhMzc8WHwcu29q8TrCqPUZnfUi7aoUTBz22kJwitr
Y9DRejAS3XtRoxi957yQXsB7T3+4/ROLZwQ+WYqe88O+WGlQfbROn5MEenv08vIUl4H8C4oMEbAL
JmHZrtWzpBITDW4Qi6+sWKpdfw5o0g+EOI6SSOfCSz4Kbnr0z9/6btOTYrGOB6k0CoQy2QUsvDhr
cYGWjMCnnAYKJ1GkWHRRdb8DFtmjyeS/vzpfCmjALtu4GKAuSNcWPvh031xk6o4Wn7wf0i9kaswK
AU0S3a5NdY5zri7nfRhhABDopBgtnqr+moGDwmHqZOdbkkXB6EhFBzBBO8+kKV5Pja7rwUrZcyNv
WEP0rkiFbAQICcUD+A+diwqN+HnLox1cMXU/r4RuwCZ/cBX6tIQBt1A7weND3GnDyBm1J00cxBs2
CGhQdB4AEyvrveqNaO18T3Ko8S/8Dq68AGMe6HVcaQGjG9LFqZan9qIA7i8izl3isjwrEDQ4aI5+
ndJ1Gx/caxEx+OW3FS2Dd6oJ340eEifn/37D85RADFkjKOMMrQ2gAZGgIelCNIrY8nE2pC/o3Unu
RDO8OkHieM4bchS/gs+CmwEKrl8A4UZSFg2yJKHRwa/sGHCy8g4Ft7meEhpF5kFMOV6hA7YFLVc8
EpUnrvweSUGZVuS7xv4ODHo4dNqANfUSq651lDt42OY6evwqrze/Vw7Bpx361T82gQJzMGaPp2ao
SkNYPrC+wlfpNr28mxqudbLthp1VqaHImd811k7j3Bp5+/522/ybrVXni1e9gSK5Oe7wFSqERbre
XrVBs2C9AU+DlJUyFOlgweEfyQQrqJm2+Qz98tjLvdiCNAytopYeU+YvEMDUJeugWjhcpIZ+Dox+
phQOlwOoOe3ddJnV8r40wxYBrAXkZlxcoNPLLSdW4dTtPJKdR/KFzq877ZU01kAZrS0MSORuDntY
UmlKXu05SzAa1WlvrNv1RQGkIjJQ3btu9YBoTLX9FTvDiZH53VfqKeTcoa4EBksBeBuiqtfKRLVL
k7zNVYITEqUuO1x/PkJvin7zCHreBgDRxd1npzhHWM9aNKkh7MFQAGU+zKj0+GF0xmu62LJUGfkm
UEQzWDvqzg+SRR++u8TK648qc3rsvFiNkPzb3yhzGqAy3v0jblCthYsq6b6ZsiSJ0gOCNxWdNQil
upGUbv/l8xbKBH1WC7oHTmSTe63gOMDp1AsJCU/cHqAdDugBU+UEXvFmW5eokgGC0brgHTyBxpr6
tZmtCojO/1zssub6q5bx9MHsx0T2e3wjVSdVWI5Ue4nS2ttQcFRs7ETOq8+jVj8OGz4HIKAZG2Zd
UiJ7e3KBtR4SPKDwqbNVy3YUyJ4FNlEWqO9yZGNUekqnVQiPnT1jlANhSZrjKEdUpCNjNZsFuEmK
donF2qZBIDoKEFn54JYjAP73vWQQX+V1nSQsStS4bccUhftD461Ny5dP561lMpUiF42+GvmLwXiQ
/xcqqG0+lkwqniPm4M39VYeaf4DyCdWBj9WLf9/jy6tZbQq/p4Wn58Bz3Jva+G4cK9hir0GmOe0P
mrAYYxMUvRT+ibtTkq6Mhzuy0Tg8iVFDINAc8cO2xZ3M3JWpww67sDR5Y1ikLt5Gl6zgVU58kjr7
J/3lA/fWF32RXkzP523TOz+PnriIMg4ZYOPJ8G3cRTlAUznqRAPm4NkCR2q3kfgFb6YUJkxw2IuC
5gyFNwsAL6BqDWDhiGVLn1M73w/2rAMQHa6othx3QePTE9Py5wAZl8MvP/jfdZJLA8qeC1LJ/byq
usvmd8j+FxcK0ujcwYwoWJWq28m8UdNAQ6bv8nGJDLlecBIiHIYfeNaNtJbO0RF6wojFtl12c75c
P4sF59CGX2AQZhQ1yZQ0reKVVsw/mn4G8GFxh7FFTMSf+Gnop/SvCN6wAqEj1tkmCj4Yw+/BClND
f92n6vyHBbTr6e7C+4vC2CgT935MiBg0ZZQ5pnonjE1IsCmobia8ixLVcnnN0LriAxjR7fmMACN7
4tjkNGN5WrOAtJsykjVd4Z/EDCHImhpNWr4BplyZq+bgoil+aPXBztA66cr1TjuG909H7LLlj8Lb
DMjYYcUGgPrmbDPBopnb2Io2a0UtghEdllUggl9slJfKcRf/8EDNWzIub6cGAXTyrDarsGnrvgxn
wp3NPDnyp3TXFgrAw9r2mA6cUKHw23ZYEH+IkxC8Qt5R1r3+lv50NkIFpK2w9h7Sy8uW3O5xscq3
dtYzTeYfqXwyxs/V2oSWvl/faGf2dd93yCSlZCowYlHCJe48fFzjcn7kZajH7saBaYSJzGCDlMp6
GTqLXHE5T6h5laljwvXN2LRckpi+M1NGjNHFi30GZpmemer3/SE2YensAOYRbGxYepq1q6jds83b
E8OnWFQFpJ3qnqmk9FBwFQcstqjKIKHXcw665IGsh3wUEYg+Xhp/PY2tYMHaFaUma0sjnLCAcokv
FnfXs9WZ9I3ooi8/rYGhItGAFF3B4iQkWH4xkA3rmqvk5+HNaYbAx3eSBk1DN/1F4j8jTAZF18Y4
jX6C2cjWuLHU70gJ/VjqTyxNcMmEM4vDVvpMxe2V7egSaqRLjhvIYHtlSXTT2kvTdkLJL/53Kxcz
e6vU/oglk2/xRu9RnzNCOma8muKKf3p0yr902olnzOidtOwKpEvUTPwCHV9fT4ddgJsWGsg77o8u
zOnEVZw3/+4HUYMfvMyIrip5sVsMn1gaV2GYwB+2xC0oikUon1MZ5PBtxIHBOnW5cd5I1HA+mFi/
x+oRKGd4kL+NbAEjfKtK3myB/S9b6tDjPSAByLWIMIB6YEqsk9IOaD6Q9SSvEbmEk6FP36cIN8WI
floAaKuzBV9o3umbFm/pYdXXAHH4jdnku4DmLkIVok03dJsZsoOIVMyyxy8ssqlJta9iJTn02rPB
rjKG7L1YiySr/9tPuRTZahXAwyEheJ9L8vEL1/8hdqD5I0PZoUHwWZhX64k8AD6Rro+PfyjpdG3Y
o+8O+wP45KdibvaLJCgAWY6WgjtCzPfG5izk5DcO9LLl3V3KLu2vtFpjv/0MN7G1qBa/egOfe9lX
7kdWJOm4Bu1e3g9FYNrK4DWZfGR5NjXmQXWlrxRBddiOsnb4sEgclacS8ir5N7PWE6Wk7+vQm0lj
vnHAYCjjFyT9p75Jmhu/6kWOV8NAfmN+7bctoV0/RTOZZysBhyQWEh7wHQCOejdva5QmFk+pgVMj
+euZFSrL1e9L1eoy5GsxhGc7sXq3Vm0SqQzmCIPRXSeD/d0ykO/mJ6rbcoiSPiE0koPOdX0g7tIc
JYUaogpPxn+e8OD+hYl+oB8O/UIk2WdLHAzRjJwRUWM2yxi+cwBuUljxxo9Awsrr+BqUgLlYkGSv
D1eqzPY5tM/NhsYMMWefb/KxYGMxdtU3zMU9ZP9kKu0tx2a/yGJ9gp2p7vR/89VnfT+tA4N/ovGZ
WKRDyuJltRa/WlGLGFT75i12iBYktAO/gtgwPIq/9057aXdkIlh4PVDn4o9vbBbZ68TJKkXRRAxf
11BXMqnacG/d986QlVC1w82BTdAqfdwfwFR2JHmeyBYDvHO7/sDq2zbTSbxZx8n0JyZXVXjmsIc8
UTP0Qg/bw7H8sYvZb+Jn8d1NEQoLeWb4/5SgOG0PfklYm0SYGYpsUpKT4OPZjfB0dIMPx60ZPNYN
N+A8IAxvYMVWLzcBoMbkQc2JzGDe0FJbGruMf47B5Jv1Box0kGgU4W24wRb0Hfp++Xep17GsOYDe
c+yMNi+b/+d+bU54713KoR07FAzFf4H13Rfz0W6kRbeytMaAL2dNYTaiKwovTlTFj+VAaoD9Fs97
pF60/S5fLeQX/hN7Pudn4v6jQtdhjaUFYvTdi2SY0DjyN3IaUScCTGEtNrfLQOHFPkNbkzY08g86
j0lnQmlzn4Q/g4NCZOnJnIyTp+/Pf32iMwixOKYcKnBAaqX9SwuIWXKXpJSu+yUJou6rvW+1fqkf
iBoVKzuyk+fKn/I42fJyZFPuImFBRzmAUeuQixHO9mYHtrU1I2B/MIvKf0OMX+c0BUzoE7L05BU9
kpXqndHTnHqipIzWMyf6+jHOt4856nqn+58GTBnaMrQclSSjyL7cRUWG9v7QpKAoVGQOwux4WKao
k6g7v624ndAN9tRoQq59QG22K0T776DKAYnQWaUzlHv2GqJk4knPQ1gifh8EUXk6LuuetGOnDq5J
mKKJEPRbzX+nC1EUKG0oIYQiusl9eU/4SVxBQ9BCjighJBFY4Z/1rb8rLj69rQARFUxScXorD5K1
JEw22LGlJok1Tj/II7NVmYJxxpt1iiJ1RbgeEEYYuBmjEPKVLnm8byKHoBcFClDCw6dSis4IaVdw
WZUvrAQY+hRo2JtpdnAJ/2Wv9jJfgacvX8oQAyba6sgfNiv7Zdx0sqyLHpDWXU+Jt8flgTS8BEGz
MGRfUhaAh4GZXL8h7FuIGHdJfOvnGPqzChv1g1gmy/uGjF1e92v/UZA/YYE0/zORZaHFP3RfRKL5
BKhhqxIIkxy/bRNXkWFMRob6SArIJofCjRmD3Xcbpvb7Atgi8VWOXytfMmCA/VcgQTRLeRFB/0yN
bpKkZrv7RU7iyjA4pdGUQo3V2j9i2bfnreqa10SWjjkO6IXnMU5lRih37jiIZJqPtK3p9w2HIPrH
CrXj8EDvuNsOI23K118kxma4rSBxiQtLzGgO+40JZuoOgHSKWbvFYro/A0cYIfw4cReHEAVFV+Dt
LrejXME9oDAQPpeWx5rPAaEzyGTYnkKiFlrrRW/KIJ+bEHmrK+nniG6oXZD0s9/5zsYQl7TwOUfl
emSWhf/AUnz/9qTJx2vDlORMwoHnQ4YP281xcrL7rjqC1Tb14d0aVbzjIDu7/6LDANHNTMDqrL7G
I9SJ8GZOwtaAKlYVGsHQx7EhROboBV1ZsS2rMN3xcQjAaJeXnRrtdWT+6v2N6JVAQbpltWO8Zq8p
1GxD+AvnaOq1SpFYq1xYKLEOeF+tOeO1KsWuVDcH14nmhHPP0moA6fkP0L8Bvjfmqw/9zevWHr8g
XdJZkYdZMWNMGPjbR1iRaKgWfwYPpB327dBGlqEmklj+Dh4EmyDbX72a45Jvciu0vLEOjUjZxD3d
5If4WzrtHIArsBww+w0uiNVWXlsqqDFq73cOIzM5sGafLjzc1IgbEg3KJ0PiEPegMBJ6iE2FXQcC
wrvJwVwqwYrfeOs62EYD06/QeHEXOoPR3Q+6YmyJ4t4RObx899G7D4j8EYkB37cHT5axfzoCpjyF
3CIZOUL40SkcJKF9Mt2oY5jTeFxLi1Fs1zJJGvqXKQsD0/74hLiZ6Zc3mBaJh5RgYZ387KAGltG9
VfAQ+JxqmMr+PuN+t7uAzr+1k3bTdLe/Kj3tC1oPUKnCJRwoPSLHqpEnwaE/Jb9So8+Yuo8Ab5zQ
+7RTP5k0ii2a2nfcZi9ASL5fid8DbxujRYTLepJwD1oK14k1re1JPHazEZX0lXqyn9G1DNoCmkby
uK0TfgCQ9/LfgA3sSdlOvOGoEvEw5wGNBKSyovIa5Gsl7exxM8pXR2OCHTT5D+tLUKVYru+EcGN8
AHJtn7o/xZWslBYvh+tJXTyVo3aAxQHhtS1vGTldZdlYAhCHe79/Wl+aTuqz/zkdThvBieknD/CF
VtuT94P3VdLd+BHmuQYEgimP64tpgx78csZDrI6+X10Q4nn7lUq8Y4pcok7Hog7c9EBsy5stdtEW
t6uk60SMGy2OlkvEouPHjgwinbtggXKykVhKun3IlMy6p+oyOhKhQTJGGrgryDcmych82XxZ21a0
0KHoU/F9VyknWznPL8526ihrBZwN8mfvQJE/RS/4sDqOnlmRClX2Jx5h971r2MAlLbPh9jMIE3y2
O1BtEV6rv7NeIq+lU8EDVLn9I0i5TFgE2FTLWE9SJLtVtxBt39RY8W4ADuR+19kNO0Lv6o+GTtIq
8l/PfOj6EG8ozKXfMFDFWkYf6Sq/JlXLMoX5Le26l0DcUlOIeQRmhmJUa8L/p5RsybYf9gWC0AG/
IE4zPgXo9z9fEPOfr5MTN9tZNCVQvVLqEu9Ane4g19nhotLp4DBhocswaZxLnEjX0fZJTvUMO5kt
rtRzhpCLvnWI3n0AwvZf6x18CFaCrC895un6rDpU+1VrL1KMaxnGx6lSnwg7VSvWoyIF0wcdpfXc
UrW7Nwa8KNeiaLKEhBHa0jPQnkF+H4ymFEszr3C+IC/K2dQczKEu/kUolwneUsg4s7hZOuxJTzwZ
41NhG0WFyfyjn4JPnChECauoxMCgfjkgqhae/Jg3O7xJ80LD5i+9Tu8nN7bWjzEvgw8T7SW0CqR8
qkMNAKGeZ8U7lBCxXeiY9cmXVJdZ9vCcUE9RNWaE6q3sdiUD3Pb9Dl5DqR/39Y6G2+LTuueAOLqz
lvak7izRzNSxUAbAaScxBJsEEuA06f4yPEITyt8j63MQfGPLJxCxChmvZivO7r5ktOIpoo8XWIef
gP9EAX0q4D8lgmcwBUKefxtc+GPXepfhbynTqHG3fDXaDgB6+ljaQOeIGvp3RTEKpHFnXfvp8N+5
ycOR+mNXThklBdqiglb2xgAnm/PliVjIRamgWq3XqhLs8NS0Kv1mJzEcKPfICwrYT01BYu+R+FWj
g5c917TEl4mISvmHgxM2U//XQ1jdJVUsnfj4WhUEj+GRaw5simzRjnWo6E7SmPjCQ5j1JvOtXNCX
f2YO7orvUJ03fzFEs+B9LWhDNk7V4NAwjq+c86UEWJXsN91NNwKc1ReriBfJzO7H9ltvWHbFXJm/
0ZvdVxUzSZw3EvKDWWtxMjQMrF/6fAsTc/ORjewRVb1AfIkFfXCJo7FgArGPxBtPFA567Dl6k28e
RSJIc17vFe9rIgyRyT3lVIoIdt+KIxHgAmdy3thgJc/HsKqSqQ4igGiANmmjT21pFNk+gnFgEdKU
iekzT9elIqbd6516gyWbCiHhvF8I5AMhaaCJJIRisYzYTza7k/HFlPw4Ed8+wBfFszyCD32e4lXD
6e3y1Pv2qa9JOkxa8DybJIyVNFMCDArA8xMVd7MGsG79PXiJ6FBUdmsxKRHkEHUt9sap6onqttvb
HFaiKMStGvOPqGHh4UJ0Pz5mznIMA7Qzk8Jf+TsCYdX8RfFOClZafigSikFdUgjZct/WPE9WhXpr
Odz0ljPtMp11B46rEcgLuG7NtXn8VtJb29xGkD9yJ5BgZzIZbr4L2L5Yfk64Cdx8JP5dXuXq79Ce
lsH2lUR2co7Tyuh1wqh6LcUIRz3/zasDNQiOTey0dww4Uae2Gt7Mj7R0ce639aoGaLIqWr4dAKUV
ww3bxUcq1usegYyadXpzOHipu9WBJVbUNA/dFLlDRxLfqwXGjiWhvXj+zdG6S2gipmH1+Ee09P+p
xVxEOVXMPuRDGNYMJSF/Ybb8oleyyzA4kxTRyYi341DOUUxQ3I9YZSDIGzfNlciYvCuoJO2GzKwx
Pol5cX/wAV8vqe7LEiQ48DovM/WDGXmtNS4Q9BAgUZ6PdcEQzFe0Sse0Whzlg5GUtbbGtRpSeCnj
sSsd99l3LmNSYU98zWw6FjnpKalndp1EypTlULiU9wuMVE0wXKk6mpuh4ytyRKLg1fiU4fNrXZO9
NdSIntksmviN/6u4BB/8FaSQTeP+nz6o05NCJ85dxsnPorSYTYQGpjUOLHbYz81mkjOiWZZpLZhB
5R8d5qq0q+nnShrYUsqbSdu0lHZIT5YjHjVKn+A0WBdl+WZTrHK0rzcIg7Wkc7F+b/iClCrBqK8O
latIo+gTAUayk9KKSJ4wk2JhhAdzLsIy+cDJqXhmUjI0E2xNtuMQPmLgs5hfAvmlcVtkFZZLgexo
dnL5ztIyZ+HZYJNKzUssMHa9Hacuvof4HpFtMxPCO2gQ4mjRXQ2jkYrRnoyDb+gQrw+TXAxrGGME
Je7SkjF87jJkgg/pBpM/Ib/+O2YBWcABLBRC0iG5/PTgNX/7NVGO5i2HLWsYstM8MF7mjpddDOZ/
pwhK6koT0MaqpiPzpDyq+SpUWJrlWnQD14y0lH/CZVHUnNbvkS5MJrEApOUTYn3Wxyi7M8HQxyyi
8pZh7iVjO4ZqC1OI+bLOo4cYTBu/D812JvyxlrNgYc3eYhfmWGzky7K0cevQdDISw/copEG7oSf5
gHDJsxH0rm0WMBbbzBfWFmMqNecl9TVpLlHNX+t5mGQNFYNyb6xDnj6CuKnDnyuCBSK+q8y0Xmvy
ooFx62VEQTdjlP6FB6ntK1nCY/AKzH4We5rtBtN8OrJrgCESMItxNZMO21kTOsGVMh+HibC7UuSK
8OH8E0aTLYrwV5UdImib6FQW1VsjtRWnGNV15mZce8cF8S77K92fH/d4YU/0eLd7b6Q9vYxnJAKK
8PEtfa2msAXC2TtLIHzqX8mTXJoogLyeK99CEbMHLF+gwXoW+hyWY4fXBMLXrIo9RuYpawCQY77h
slVX5x0BYBgSyAX8HpLuKkuAAKLILAlZUi26gEAow/A081KV2Wkfyd1140n2gzfPrP4DMlArIXqn
IhXu9Z63G6PUP0JiW8s6ehFlREQ7hrOWsPRyMXwMHQRDtJ6/R0WmGAMvC9T9CnSG7yoQ68TYhjxw
5llb1ufo4ECFJMM8kX0JIDCkFlpzaYVwo9HODgEr0o5iNbofZ30lB1Dm9bM4Kk5EIbI5bkVeqoq6
HEk0MVl0gVTLDYsyknpMs3k2CERIH+PajCSBBitDTTjvZ0rKFrl6RY/rhK8Q/Qep1lHMbwMN6TS/
w7J/zG1z1EnJwiet3WWzDvA+FDlNNtrCF+xumQG0fcVun4/pGm5tl+WZhiEnghQrTKeP/wWFVTCp
30AFj8/ZVGnltqd/TfxQAuwT+CcztYSX9awQ0MXerD1LO4n+yxJOdwj/obwMBzjhvlvY7IK64M5T
xBgoqoSXO29GbCs1XPYgw9I5yTd1EBXKJ9WgYaUtvF4qMCWqJysJwOtAbGWX4VbQ7poeJIMOzpuu
nVCh1Jx/0nP4cflYsWoyDjrZwGt4H9pguDRi7xz7g0wMZkkhSK0gQGTipHEgSIQc1n+q4pYQxPnD
gVNePY5efu5bpge1H1+bf/Ek1ZcVsNS69A9Ksl4jRb+jOOhg2WEfXCqnl2lh/l+yVQ3zvOck/CZC
obUepWgE3kVQeguKaB3vsTbOdVvjf6mW2b+15USdG2meSp5ae+vnP6WjFKjBW0oWQ0jhX9ysXzHb
JxUeAMT7HTUhRh2SG0uxe5Ry1xPdCOn4ENsfreWQj/qpIaNoOncAhmllEkaG+hrHwd+COHntqJWS
cdzUqm6Gha+29GJgndTMfY+QRI4JwzWt3YwNJDZDdmbqfrtnLmj5p6jSU+Ojt/TmHbJtWkENk2+w
YVYQbCft1Lo4pjLA3Ms0q+Ph+vccs0fLbtbza1f/z945QU4PZ34vfmV5q9wC6GnLNYQak8lQDvgb
uWebIjrNkdkCITo/Tim3v3fEK8Z5BLULqSuxsAXYdWGvLrwkwRDy5h4rcH51r1fJv7ZgsNGMnEbM
5tjbcUQN9KgH/3xbrK70/lwaI+lOlf/bwE4e5iMvgUv8uK4BpxTSP7jHGMcIMmT+qp1sMV9u0VpM
X5i6UaNjauWdgqTEilBLwCIYRJWEHYskpyZ0ivnl72cg61Rj3KJlz3GEOwB1xISQH2w0Y8qSyDD8
RP1ZdM72be8lX5qPJx5zqOcjYEEdGQvwpHGZBCyqvV7BRG5ZfoYuCJhKSFQbBRGm/N858oEwF1SH
IKTWbJkwf39XWQbuNQF5ksWOVedWqIC07J5piteBNihm6lFPtJcPbfl5NGwB+ejUo8FHW1wksoCE
r28hV537ghE/tt6qHrqg0axMMN3CqcxwhNr+Xs49zVm2sW3rhZxMTkUUt6BZARhIC4uK0svnq14A
RMfEB7MPmWr+MolBn+o/uyicFWLRD+d6ut4h+mEzUbu2eCymoJENbKg/pHH+0iZYozWz0E/gpwZx
GqSolWVO0wKptmjH3eh7mqWhPVgoL6PlA5CIAoDS0LR/4QuNZCTQbTKii28maB4H31nCNvJ4Y7dk
VNDiz7N8gdqUXLQdG5i6XrP1oDe/G0N881zhMFGeW244iNUS3fZUz97wzCB5dd1Q7GsTybQZdQ7o
F5MAwP7T3yZP1QT9c9kgQznYC1sVtuzYRiDml/wv+R20qRxCXjc1RE0Tl8yNfQc3DnQRnmPzpAER
sYD6ch76lbIb9PRP1lwtqzvBV39HoH46G+p5bfYPyN9nTrHWbtb9xhg+FfoCUxpMzUeMvSE9hF3M
RnPZgoqrQORdfRzjcadxjDilveDWyUSTydq0Elj3OW6VfrDfdDvc4ukfFHwOqg4I/D13XkgyRR57
vqu0VezLqsJAWVJguh1Rh263BzFzlzqeKLhWufHHVdGwjlLOaNOZQ3yV3Q+oq9vmP5Fg/dw6F0/q
BkRCbhRcrd6KGRFT6OFfGbK+XSfBBifgnjQ07qYhVkgL6M6mcOoSL1LyRzIMCNTLAqXucB8P1298
TfBJ4dvUhTFZop4+i8whwa1E9f/3ZA/r0I+DMb6QfC/TgyKAwKLD0f2766BUm4BfNkFwKmG9hpZz
37g8327s2ytKyHpnARf1XNkeYCEplzN9y24d0LMWYR2FqNdfpgUTd0SN1QYZsozei98YCo8/OZGU
k9EKJfRsyfgK4qRyuUfLJmePPpvfsi/GOISurPJpNqcd9pww2uK+3+13RWrEW2yI1n+b54ZQEPob
03cDET0A+yf18PBbcMaBpkAoLG+Gm96co1UO3HCaGAAYyGLmH7mfTEnudjeb2AqWt23LgXo98uJP
XJFwDb2cbaaPeBHHtYIv8JrcgvxfEaf/cVLa+pWWbegTrTbNdlBcfw5Tux3v9svEdg3dJPP4srsZ
Zu5nr1GH2nSVqNC0OYFK8H40p1ZheBz28EGJyX3Q4XpCWhDFA1iVuSQvbLStWs+XNQVZFJgVg7I3
2S+l9s0jxtC1JlsXH+m5kbWclWFobJcGIETiQ0Qo6kBgOJZq0uHVdHSy1Y7GRZYEasW/nJiMztBV
KBPELZ0Qx/j4jpKif1wi0rcD5rEVYrkRacaIkV3ra5wRLz8JBAm7It5R3ESwlw8rXnnyEDv68MyH
JUGUlBpSWcdst0GMiAyrtnRYzKyrxM5NEs+tcF6h9ia9zxxTqjEP1RcX46BU4RjmcfNNgpjPqP4n
sdHtWBrN9ysU/gcVGMqQB0kfNbc/57nZx9JdoEp8MEXQEMfIuSwBfj3J/X9EeW7DDnZrMxVi85lt
x/5JIzAiDac0aAo7preskBF0LiPyCpLHqFyz0ROo9FErITiSbOTII+FGlP3yakYVfvGiunUZk/zb
wjV6N9qHa0DRgDXx1RaCcPDcToczLw6Aar2X/UoO4Dca2S+DGgMH2NSG4hnUGF3r8nxjptUo/A1B
jqieINdkOj4/7NW9HuMsdYmvOTcSWLXHEO4cmLkNMBEglKX42DNYCw++sKugzfZU6IKNkIbYstDl
oJq97in8j9OM7utATgaWtsaxR0Wooucha+/ZUnZ8njlO/XcGV1ncrez3wvqjtmZSwSka0dPGEwZn
nFWdcOLj3T+34MbQXVxrNzmhhu2EeCQdltfPsls8iwg4fUZX5Z5DclyrVPWWk5Wz9nPHYiclWTnd
K3RFUwaChRqg9JLwpU4+8MWwrI+gsVqKYEsOy9G2TmIXEiOWzP9lipEcH5QmeIVJ86Lhtvc+dn1m
Yp1XKZU1Pjb1Qs/71qVtoPP1Mu+S+abGtnTfQjizN0YYXichhdk56gPZY6qpAJKambE8Yq61Ihlo
SRL0Bx9XcrnqU436q6BoDaYfLAQ+bVF+L5XtWkMOdB4osAlyTuzQdyYId0+AqCeRh4Hc5f+C2+tM
BTPMARPLov2mwyCgRRD53vOjWetKn/i93nAghzSWBflJLwKoiYAk+qQ6OHyyeORvPv4gJ4JVSpZg
jPv+gIdM+P9yg5UeZTj1y6FndXh2mObAs508fJV+a3ttX1rJ7wFi/hUn/pWzwRaws5rdaGA+IGf7
UXpDw4P4k/iO5NX6nQODcS4LSJ6IBwe/SrGJytOsN3nVog3ip6Pr5S87t+QVjjOQiuJZE5JTKK8C
qEmk6bQd6mWWtgaaex4DGLLVuZkE5rY8B3wVu1tNc8E+XWm7xuQe1x4m15EgAwbKElMWne8nvkiZ
1C6DfewR09yhCSB0RJn+EbLpELl4ZED8Kh+GraFeMNyS1ETU8VksEZOvzdzha6zuzyR8W0zopcJz
COOKeDpWjuGbMG+1zJ3DO5EeeTlk0H2jwk83aWdeMrCXGmQCfqoVL0FlMn8w7PZTXLxhRqyuXkg6
AiX3F9GmvX+MlAwPgey0gQGk1nDky4ufz5wiV+Kl24VrCrjeRyxpvI+y+kZutDjSwhE5dGtyV4fC
uv3oA7YQTtvBDTLOK/PZSK+qnn5JfexETulrQGoao6lMwnIuwXHmAB77f9tNQyo4TAbqpRxd51w+
9kQbAuAdGw70ehq+exTwcrw1//Khm7A7KH8b7AW9287M/+Hb56uvS49lXV3QbPiPAAXCjgaxlwEd
Gprp9t3V9gz4Hb1wOqb0fAs/bwxrmBSeAWPhsyehWR9VOd2ZdvIBaszTlbus17bdMitOkpunv/7a
Zc9tOMBWjvSqGTXn8N+R/z/Pv6X9Y4gt5bXJPhHWGVlkgGj+OG8Z9RunTH8See/2CgqYx4GxKX0a
Ay12+s/mPkMNu62Ed23VpzbVHYzlOvDmc4MMsSck1YRpgaeGedrINo2U04+/zdiIECZsnqVwgTLi
zwqpeIFYhNwj8uoCXmwsf1dvP1+AzdkyMQBEj4N98vmiYXJywViqIVmoHuePsKwNg0lCWalTEhGg
Tk9soxjoe5cMTj0owgQLfB8duhh4v1bZ0au960DfZunclZAjBNTmbs7/F5eD+VeHKQVfwgxs5/0R
CJx9EFq8vDWG9NF7/3NagWYw7kolnTcAAAoJe1zxt1+vIWztEx3V+9UtlU8bDBHueRZI13h4pN1n
4BIU/efS/tkx0G6rWUGB+JOUH0gYhrCoadmPyfMu5jMpoA/Ib1FoVGSIq6aCq3iipbE8BRCHe5+g
L6MLt89/dCCLRH4Eeoaw1LXp370u4bxBVwRXaC9QhpEe3K6KwQvqu4iDirdZ/tZY4f6PP/H904t8
XpdqOAHzQ91FC72HIIAAftHorwU8u8ONZaxwJji3kTp/PMievRmnDhUnp5/KXBT+pWDpEmrVliv/
TwG3l/xHfSRtVHXnmZYXDWwqp0VOVFHVDjmtOtsr0spkCeTutpOmh1hGFmNIscWnJ9sW0VbAFNkP
djI/rs9nENyaiM5cEtRfLUb0l7GXD4s8y+dMNJi3qXBQ0uMsqCvrEUU202+S9yBREOJPb0iCIHOu
DNK3s6SI4bOBPmIe5ztFnV7+zDuGxI2kKgBd6DasCLeRu5C6iBPkNgg4KfArb6Q1hNjOS2zTd68S
PnicMkislfSxxZL88mnOeJOheWUI2zTJBQjKn62oxaV16pshsRptVrudkKTjRQdkl0iJ96JcaONl
W5qoH3H/tQQsCl8q8n+3c4G2JJa3Ca6a+jayblgr68p2ljHnTw/lNSoWf4n+Rp6ZDcuk+sbQaxpm
wCxUMb+SQx4Npnh89ttLJ9gfOpz83dga+bLogf2np/XiPge1POoyOK42LZSDhns0wUIFJpHGTx1B
jm0gA12MvRkLQM5ZYEdftdr7oQKjYItpb9fleTbqEsg1GkICo1iyHrzN+ErzBbjGy30ks4TC8hln
8zuvSDFvNGUpFXENJFvfu2Ew4QY1vT25J6F7J3VHOKmFwimVmmyfQn3FwlmO6JvprTeVGg4Rx3gh
w38qm9OcXKgyA2fvT5ZeKJZ+KecANY62WvrCuYjF1m8Jx1F98ZxdfxSfrcjtImC4gqpaXZ/Okhy9
IaXNeNYtGVzsvJ+08VO/qoonDUpC4aTmOA9IdxRL+zDTNjP6+AYxuB/2IlsyDaA7AQZFop9l4MK2
9G/bx9VES3umt4JyiVH2aOhwheLIYI8EvrVXscXeu1y0QJNlzSlJvmZb2iw+5igRWKlFKJebPiE0
x3xRfnf6U6DMc+U0FlhQ5X+AU/YrpXmwB9ENbHSrezhvQnePifDwQ6N9mqpCRxteXE7HA0mkD4D/
cs+3WFFGnJCrM5Tw/47ve6RPZFbyKjcQhnQ7DjChnOSRHGY/v/GNK09uYV8kKWAdM3psB4AwHe70
mS0OKEtUvnK9Rl9cv16SYnuI/T3JEDY9IUIS/7yHDgDIpeS38xwNtaelU3RJ/8MyMod9ZAVCvJb8
jhDyYb7V5wWdEpNe+/j7rbMXl/8JR1H5POa1qMGTVLdJI/HpE4bsLQQuPARfzZf3BQRAEjNMJBjC
Lj2AK/sLL3b2JR84fakHr64C6oWvbl+dI+v+D6OUtnzYsws4DM4/B4R6VconG9rk140su73//KQv
1Cge10zC7VKDWrwr1RfDC1EI7aLOP4Sfe0frqPJdoTYGEQe2Hb71oLsLmwQs7mB5GGAJsqo6nDYj
RpFybkLSkcZiTOKBfTy0hGlAY6RN2Lnas6n8jBpYbNIC/msXp9vEMJYz6cEOLJhLH/fMJqST1kSH
RKZw5M8Pkp5NT3Hbmh+CM1rOYpx+dP2Qvcu4t7PeuAvGiMz+1MCEaEcjZZFZ8IZJmHCILCl+J9jX
+RnWXNgwUbSQNR4YO4+Vxu9X4qkZ6Bnp5Xjx1RiaJ/MyCEDT5qmFNfvQkLD1dXHA0Ke+gx41PRip
s402+wpohGz8KJybotvV+CM0QPFVEHyaETALdvMk8U23mAhx+fPdx6AOQK5QPizPOhlMYO2guft/
ibaa/oEpRYw/E/HhCNgIWSf1+1PMs2gTOCHCCWsc/vTCMRs/tBLiaK3yfZ20gvYS8L/qxWqGbENH
XZkGXUqEVbXVGMGqR7NodZ4kUYQdg5Q7YnYLqMUHoReLcmLiWBZeNOGv1k9VtU4rghjU21u4eeoF
WZuFJaU+7YK4CBnAvgxG5ccQP5Ny4EJq0pot9+RrnUnLOCy78KBoDpa5hw5ALem3OB8ueaABxPBK
cTnVF2RLuSpatn1CllYuxr/0Afwrb9L84nQ0p7iMIwi0+8Y/+tdQJV0uvpIXcBuqiDY9WxGvWEU7
ZLC6pXV0keBtV3TZcTZXHiiUsfci3WAJmvR93ZiFnlAGMEKBAJcxaJEAUijzeniFde+R8U+7UyKv
D6YQ1dQPB4lqO6MKL9egKCC9+2ONPGwfwp+//pIot2ze1DcNTQk32vYYSrbFYTy2QAcHKaLGDKgQ
k8wLDDYvtXTryZq8uG68KRra7/2VAya/RPMCSR+vabqRY1RKpbH8TeCeFnT35nIkRmMAVa8KpvkC
V+li4w4Nq6vZ4mhkegv+9oYStmCdsl7xKZs2QNe3eLqDv4e3gTybw0dc+omfBvfqYGZ6nmv1cAoQ
4riM8Iy9RLjMuAWz4lLL0pLFWuRhBEjyUtvDWmZH+xtcmYJ7pweSLFBZqYKMITqVyjpw/toBu/zK
GQD94DCruw7VV04z9vbYElnFo/LpTN+rMFT2G5oHXuCIfUpEQ516/t3zr9nl/tlahOIDxySfVkNy
Wfshu2EnlZATlUfF1o82HJRa6sEN77ZbUeQAs7FIyuoh0wmumr92o5fxlH3TNXfdpPfA3InKWk6G
7CXN32/fsq42itpX0FBopU9dOcdfuxyVcoFnQ4mXaXno5vNtLtIzJ2J/W1Y/qN8XoHSODd8eBfgW
3Tym3YWVCykGUyRq3vQykDXe8SxeT+NzmWXSLJ2+TqNKcDT7Z8I2iDreVvuK4mVudfEqwyfKmUnd
T4HKDXm2n+LbBYzdu8IQMd5XkERjCvVhBnUm1q+e7hDla2vRYsyc79SyrpbIvw9I9C2HFs0XoyuV
fLUc/cF9UHVbSTpiI9MrTOzxrzF3EEq7VSaw5667mTLoesAEqo/5TYKApc+BObp5xEZsyZdZeb3J
xLuROO53evE1UWHZoP2/Qf7KMzOYzN8uEH/tEIbJJxeYB3PmjQ1tSlgZde2QOIJKQFqXFGNuPms7
MNdJKu3p2Xzy2UX4IL0V2AiDRQ4Bi0XguaVlJ/PLcS/rFrOJd1gQyrmmZHiddOWe1r+APAyXvFOp
7zp/EX/AaUZo32U7Rz3WWyu1RbLOEYHcBgz/OKneTjKU2a5ptyd8GHRs+MvAELSm485MsJptIIHM
StGf6v+fOgKMkKkhC2SiNW0+8iGwFvOMMJMkqOGYtr4T7JX1KaYQrfwJctjQfLcXy7EZunfeEXs+
KIn7FxIMih6f+8axaP+3kWScL8cL1d2CGQagjmXn/ZZh86iib5YcHEtKSwnmJ3dQiWncUmJBO/OV
7Ej/zrhb2IBu/dRetp2o0TUlMxJR0AR16k/3N6oyo6gqwct1Q+lCjoF1tMshVIJz7hFKINmvz1SX
YguSHNLgEw3lJBHtcI1+D4tnCLyiDAC/oobc3+yKgAWHDCc6aild8qtcif4RTvWbEbrAmuP0aoVD
SSXcTqOKMiREjN/F337Ev/nh/6wAjYBpDgB8B2wApBgqsF8FMs0birLzzBWOorww9/eMz0UkK/wf
6mlxojGFU9Lu5Si8sQI2RrPy5uE6Qsrnwa+fBYLFEm/25UJHlhYke6UXCLlZoSDVt+kS3+kY3IBq
sOjXaPV0wHhq8vvYzZ6rBsbEOg2SyzRp5amTgPl1/IgicvblK15bxkIzvIcAKNyoyfKO2bJZO+P+
TMqy9qAz6lT12PFjXeQ2UYGpSmH5Vk+omy6rG3sReR8hO6uVa02ZBv8mrIlFdqiidVJzOVHrHzao
yyHS5iv9Y3F3yAdHiDuh+49JIfMQcEkqFxfW37mO/FEEaJO0L5hL0CO8fFuSdje9gR4RGCkvls/Q
UEuBcHvJ+NP0MczXOwljUjjiYZno3LxCQBLZMKkmWjnMH2KA+YSTE3Q9x7yMetuJtrqAkJsq6iiF
gE3YEFZVM+VawIVDqEBx+dBMnc+nF8Wfcn3n2hiZ33AAF/uysQGLUk0uJRMvv97fguWzN9YR/XEt
i6zZgqAiRyr9UqGTSE7mZa0fJJ7CyA0ZE8H2v6iNFbHwsXzP5rZCjyDFnkgJ79tD7IHN0LvO8gtI
GWJHsqrl9mqK9FIno+azQ4u7YN4vcbahhWW1XtaHtrv4UH56C2TPr4VVS+eKx07DeGrDP3jySSgP
1gKYbzIipmiwRDdo737CL3g0yHqfuV05d80WmlMSMEHWTnn5a9O5wGtv0DmheDckKVRdYKBclsEC
KvaHqUM8UKsNVGU+l0DKDrNnR6YTk0fUDQCWcCTNPyEe2JyuxNzyMOlkQeJgSw4ixUv8IdDe9txL
isaEfFW4kUYWPUiWLxjhNwkFOBgh8JMUqq3vWVhq4Y+ob0Tr2iOeejJvuHV8N02YqgoEQ82n1f+V
Jv/smdDm659lKzxcO90gPUrGeJUKAJk0bKYSVeoaHwfejt4Q5t8YIGFwRXBmfLWVrvLn4lgVW3oK
mGRSGYgqaBlCz6moX4sCP2XiZfPv54pgoBifDpcchSeectddG0A8/pUfWAEhBJLvB0oE0iwnoDXg
6iWivFpIYkGF42rS8veA/s0i/OcXfku6DEuvAOoBcBMsdCc4AaO+LbKAjSk4wf0LVC8mIQdHNeq6
/oV5C4ABoJm19mPHNPTLeTLnnArK+Wyx4GibqhrWS0WMkRCqPbLTDlfVXJf5F16L77UqCef3vDOs
ZX/rrjihEcAoFx/Z0z6/At9uihpqtkmSLlEhFYVEkF96njDgOFueFHJ7i4b0Rs70eaKHfC3y7G2h
cQTrk6n4EODT2G0bMmicbByQfyE+0vYxposxOBGZJy8Ht5uA4sjk21uCc8vA1gJ0RbJ+Q+34DE+k
6nAa+6SrffAWOww3TE4+CHpB3jj3J+84gBtzG6y5Kp+j11GZDpUru6SC+MlJAZcPYYOjNvm0cmLn
hrebybfo+aLtYw/2PrzDSeBXfu3MLVzzkq/DRZUF6Y6WM0+A5cXJVscstMm8B3f7wt+Lti74zQDa
g2yhURkUCfwpgmeEQIzl3Dcl1iApp+v0+viReoNqJK4YH4m9yoMD1c/cA4GA3sNKNNlyRktcWBx9
GqyFYYhYmaH0BqWfawYcBQyfUFXYcTB+K4zZQMwkcGxDDK65XQnO145SkMt1mtv5bEHZjXHQpcud
mktay3Sel55hwv8K8zFoGSi3ggnI11gq/aMWUKTz1yBiM5FrktMsZNV/BUvwNQA/tK88QXM7KJg4
ysvT/dCuQl1+bo/RMXpu4+3+7qqdcAmXaJwKGft5FrVMMteTilet29SeRyRsCAbSFMk116iCVNRL
TLCOte8feYzZf0WCDChBhdrEdyytE/0gJBnaWFh4+DuWq/RFIAx0s9LWnwdonNYQRz83HE8rzN85
5ue+NS/xBt6zZVb+eHciwtw2aYhwUaL1vATKCPOcyQtrDdAYD/tckMxS4tngEGZkPugGXA87dSTW
TRqyfl6CCQrPM5EBdLVXBub8rE2WMTr/xBAj6Ja8fUl40XhAPQmHkUjH1JiOHDG/Rm13KHpPQnR3
KRH0yLo8v+1ws2yM1JwFgP08U3+q/KaiEAaj49tbCdFmK54U3ezRYl86ukgnpBuGogpKp9og9WTs
O3Lq0mL3DSOE0iRcSSKZje/NoLW7Zsbd7ThmndsYsjSwbgcRpXbkImZ07IlOftlYUAJa09ck3VxV
vWs7nb0y3KqxKO4VwW/J1LHcdeRsy1yOACJgiT1wB94rfaT7zVmi30o/uzmlTEh2vQqpmkxEeIrB
w0/4s4Yg5jROgoJqeOYwecaAdonEU2vjilLmJeo4x7ytThJOCIh33t49hreobxyAu5FaUCxmS74L
W5geCmGRxCj0nZ2+/9xOIH+Ox7FZx3ZGU5Lf1LcHfs8WvVf6Z92KkYghw2GQITxC79XJsWzVXU/N
WALbNZjMTdZF7ccwq+lO+zdiPiyeCW7DkuxTP96hBpXYHGEUYD6aagoCPyaQ4W7flo77NAvtEWEv
2J5GoBg18IWh0Ty2WgfAJJSeHNJrBXtRPG4aYrkthHG9/1RBf97KNo4F04iLSpDWdHtqtvF80ica
Tx4P4dI9fOXav4DejmdDeia8oKDq0ZylzfTgNdHK4QSM0HW6KE9Lm1AQAvoG8aHLtkkgSbNDG5uX
+oPmrXQkMkodbyJr4EHEXi1SuzD1kVLzyJpAHSD+rj5VMC2SDNBcVt9xQ6/3VKH5dsswp9TmTwl/
HrOJFlItXuojdwsizKfcVIlCoYyMlyFUkG7qm6eNYQUer0cj/eLPEEe1IwwgxghLG3X7UbSPPZdi
2SMcp5bSuhnYdUtb0w30inyITHWFSKrGxdm80eNLCuGfIgzqWc0Sp6E4n911ik1WaHWCTZyiVSCq
ak1TwXBbTfMQ6orUfmeLHOOna55+s/LmJvjCSYIEH3hLkxRUTXmH8w0vkQCPXhq0QtOBu2+7NLIZ
PmqcI0JGfw6RAF5YgQf6eL6H+xzrHUjewRSMa19VXN8V8udnONLCp0muMWCdb0/a4O/HIkMMRLZ6
JBFZGjer5jK/5JL7I49xyYKaPr6lcwsAUd/RLLgrTKjXS3bwCOphlDslJMv+Y8ZDEmEEtXe8Ex4J
yCKkaqfOVw/oCV7gpj530h6W6rZgAO597Y5kAm5TNj4h8pGabf/MDueZOqOpeJxkcWsHfcKQTILW
9DOAPUFb0z0+fBvTCiccjI5Vxt1KjxMMPMhQHN4NxohMynMpWNW61CtUF9csGf/sfHESARDbGbvI
YPxBtuk8FIY337p9YIti1lCFMfB84F9v4j8IE+civLn3RPqnNSndY0wCa4lReOkNveZosI9ErlSJ
eNZJdWkeyngpJb54cQGN5wOhZYkC2h5FeuPest5ADaDVqPjIYf8ncCqm+MDZGtnN0SpHWl7zm8Vx
AcOv6i5fPkOlcVAiY7cN3LvpsvgqkdOGG3P/K/WapGm5U2Y4jBToIL0+gNyO5+7H9pqNDGC57mWz
KHNG5aJt9enKleviFtSQb/B/yNPM9XBPGcAcsX9GSbxCkrAGUwzMjEjqm+9nRgHSrKM5+QL/D0Xl
CORYeKIeYkDxBpft1ptkyfHmIbg0kIWoyM/UOQ8dQ5xeSfz04dgGTeAEphuzj7SYZ029qoT7iMYy
/oJHg6cBKIlyyOgU2ALph2npHQ0poZynutFDMc5gv5o9RvKJG4dauMdWSYmlBqPiGHUWakCnH0s8
TwUv1nT7c+Y84w5s+wYQBvz6R5han1kQfeH0FDQ9mFAQz68lNuUoclB1OgoBMvSF/nIHnZ3qojV0
xpRZh/qWQgwGQydJZ7TnjHfbHV94MQ9JNGCiXMkzJNEGGVukMAiLvwPap7dVj33KGpDiGpO8gsGy
E9XyBVjR4ojWE5y0eCk5IsOVd6IpzriNs76EoXbqPnHyh3J94gqpcKSuX6BkTbBgQmYRLOHJZzG6
NpprTX8QOaI1UmP2Y4Euz1a31BXDQ4BgYemm+Py9I7xIpjQrIKIlnutCCkTVQDhprxJLzWCPrCj2
wChjhlaUysU1G04oJi1xHR2YyZdACNNR15FzfawoTQOYiB69w6geVw9NrjrHZUb0AYch9rdc5wUw
diFSWfAf0fjke/+7MGSYBDdVCr0gvTPC3d5GV06NAYIMFmQP52EGsWDnmwK7lByGItGH2JMuO4S1
Lc39yVlBIFIEOTCZZBp/ikaNtR3K9EYMM8UgboLpCSXWUugJzfePtbyF378WTP8GfIRD6xycu194
YBi01uoXvahJRMdxwI2rURY+Zvp1WWtlgpibDwJKaeO6+QrElk/v0bhXuEc8xM2/GXmexHb9gD3I
nupku4iAVlqvJv74njNMHPN/MUj96HTcZslmgufj+TezAgcv5vO9MY8LdLFsN6JBBDBc2eLQrE9m
g9hBjL8d15MCS+jyPIF4ctZa9XadNQqgBPeu2JlJSzxaG2M+2fp8rR1yriXZC8zdPkLqo/yR/N/B
/BS0U4juYWCnrPEyAv7N3J7dsjSJ3f0jHH32VF63N9Mavu8ZRSlrWMB6GQi2O5QLS+gXWO9mLTra
TqxOC84DeoP08rioudcGCDz0fbjr6F30TlqT2qBnNLXaOwwn1FORCfCzZZ9yRdFUw3Zymy2dpikf
4Rtr/gHQwWRc3LRlzMMPyBt1stPs+RTJ2OlYmuFyGgYrnq9t6zqz4K6PYGt0U8jZDvpk83e/FXiv
5WzqEhrTdm+NJeu02Jj13p7NQ10YNjc2aIUoPIMpXeqf6QFjVwZCqPSUTOzdv2yUri7s9KIAbw8h
8VR8zi2LSqq1RbnpN17vf+nGfHBMghX6LqL3Qz5N5nNzH+EJwmd9d0CKP26FHv9DwAVmPZL+nkkF
AS5Mlp/Q4UfeUpVSUK75azEVFeKGBHOvqqMfta94dJt0WqDm6Gpm1bj9btBD7GkGZTfmBeLMfWO4
CbzRyCd6a62jnKS5XxZ7GzomDpAkCekBNToUzdM2rw5Twyq/vXEfGujWHE5zgIHpCZsp7jiGs2yv
xxYVfVJyjwlUxBQuiePZM138q0BP8tmtOzE4hdLvzNevHuhO7Jzt8WKNWq0Kx6l5wU93sgDvSD4h
bQGk2kdeFCbkFWicWs2Dk70ou7La6o8oc29ABcTXaJjqf+XV+V8hMyZcMgA4v+4+6qy+Ot6xbjiA
lOJMx1s7VX1BzhSy4x153qjqsmgh3jSPk2qvWjnVXH5o7+QKms/1n9FGd5EpLlFvuQc8cR0GVFCD
33C8XfUmHtE7gj5XDW4UrJynDqA2iASiWkzGjMUGwXntX5whczrxbsri9cw6JRSLkod9WWHeD4vx
WhFtbCtgi98sZoet79XR6Q13+FaoIq9ZREBAUQLthFubLh4NKf4ZOUKfF7RT4DUFEAgZGKEDrqS9
OUe07RopQaTsJy4Sm3b9ygTI6Go89TsH1cysP3ufLytRxk1fh8b+aKYLNFheag3hXBCTSImZkCeC
7MOiGrAJjXCc6BUNSGqqGPjem/vGghjZBpILcidFgPuJjKDA45a8ZnXAH9v3h1SMXB/WL9RMZhq1
274w9XcQlfa1reYlcelZOd7rQ6He4J3w3YFDWx5G39+5DeEQ1IGqWdDrkhbspBP4176p00OiDjrZ
woLc/kzgtb+I67ZxlrEPOY7yFTMyrs+BWtxJg0nbMy6HwLpZ48+wrvge8C7zCn8zQQtKN1t2HPme
CSk++HdFtUBeozc/Qzg8tcp/ARkqoKknThMXr7qc97U8DTeujTBxnEBSmDvj0ZXj+3LWAJrMp5wM
5IdttVsannzlYobi3sJx6zHL/7VGLT3it2XK7rWd5QAgcfckjTbL7A6rGr5zpHKY2+fKvm9dZrU/
zk3cv4KNkvFpYMTyxW4Q+VQwGV/Ce9XFVeNUnIpp9TzNN8jyXUZCrgDmVEbJE4OA0SKVh92z7ZZd
0iaeeAvR2cE1ezCCiKbsiF2CoNrDo9kO07M6+K9f4POZdnElTVXtJUGQlvVeFETeMnaIqX6TonB6
SUyoyxrGJKIFNkY5+yA00hxTmZX56KPCsfMoe/Q2dc5F/5vIb/HmFrQ1FjHLA/avBnTxO/h4/IkD
BYpmJ2nXU7dnq9DeaoiC39gWigfOYJTEoEbNazyc/psEO7vFg8kLk1uuv3J/e4fFy9vBndnhJCe3
myC1FWTDmHTmxCAdV9DvqvK+FJkyhBHkxl57+KNxfH2qHRnDNwdRLglEKvX4xGdob6DX0FoJJd+Q
Toz/E4xkhzza9vR89aO8JmXipu36D9JObx6u6s/HkFwj9KABM9iOgwdDN1e0KIALGyVtQCpt0khu
tG9x5EuHPdN5oTaFN/voweD9EgTzHFsoH0buphiPMnlra0nAt0Qf8YZHaMh6RtTDfzeqne/YJ48y
rCdFOdhPtzDE7Hec3SzINUZYMCYFB0RATFf0sobt6fFOXh8KpB+SIVPAF/nta7YJW5fvi5fIQVx4
O8Sp9frZwEEg+x9pLYg5o/AidIg9FXtFRjtpe59CtmC0laZQGhOb+eSuO547zkDJDuhacpoLYsP/
BdEShMKADVHJzjvBBuBA2Y5etKudJeYb+w5eyCDqPbZjO5OiwFADhhJ4byJ9f+Xq3jYlpigBxeRk
7iRVoQaMH2+FKKslwQ+rLcpEcpkqsFGGO0s/seMPm6YNBCFlR8bxFKR0NfaTvwmOEpudgnpGY2Gd
tMpW7vCPTfgr2HXZ78e/nclj8QhqyNYmRVvA4Ny6OAqRFTH/IyCTm+12JVDitUWQrnmqYvKEzZmm
RpA/bP4NWmxg4lh0HjY3OoFzfi3KBLqPpQA9WkEiFUh4JLIQVwBIaMnN0jiDqFzlWf1qmcS9FedF
CgfNxp7wXfFq3Fo9Oo4MJfEKRgIiK343re8uInZ9LT6t9Ydo2rkBXk2fJM+3saoQS0aA8jRw45IP
QGQmXtlhQsdm9AopUjUQflwi54wlP/Ryrhj023lCmKNJDQK1pOixjBWj+klPyakaTfulKbNvyxik
bO+rWxGZrHOQZOyHpLttsB4U1JJtfedeuW/4quEUpfc6uCdMx2dF6sZV3XGQXBvU2h42xNtrUpWC
Np/hRXPVF0j9TuZwAl1AZTMvTP4Omjqz8BPd43bMN3LQW6L073NDKlRySFPL4uSWhjcaxwrEsa41
WhwgvzZA1c/YCtlHqwi8X5SxktP8jRiNOsj68uynrKFgvJgy1LIy4tJ4J6MZZAW/0VP8VvbgoYAs
5fc2I9ofnrBi13bZU8rx5R4K9sBIpSlrGt6+dYE4vIAGFQeXDdph599yaF0TWKk/TettJBEDMk5H
2HoG/QfkVPbF5cFsYpeNtNdm3+CZJro0e+hRRH5aZv33+ivSADdoRb4HcmGekccNoX1pjsM1+R3r
2qCfKRgF9YYCbXY32l5LO0Qox8rTJXgV0/FusWI7I2GwAN6duEC+ATW6cuIj5BkdqKOBy9CDXfTU
pwa4rJJve5tv/WZlt8V/9Mps1erln6hWKEydoOsBTMENVSDGiuUHs+kg45xIsFuLGvTX/R+qY9Nw
Jf9yF4xfD86reW0U60Hq+rXweCWdOLXGgoRZZgFdnYihs27qDIiYyg0vzzCPT3/pDHygFhe6eosk
cLwdSTIpIckWD1lS5CgXljs9gA1jhKelvhFTIAjcuKti7Y07C+MQN61dgq2t+g4ntJVmzizPUOEj
BCxOHP/KohZae6qBrXOJzhUI6QbNXeCps5mBzfc6CZ4fU4MGvBbu9Qqv30Qk3hieVeeF/mW/3q6a
FYSOiO5fGju2ZHBe/8N3LBonLdt/v78gns4p5sej32JwZhw1tGvkCfre4g1Y6vEhK5QUX87VizCB
faCNT5La9Ezzmi7VcviURyPk8OJToHEd2t2vquYqpqOqacY/csLwLqsXkQYuuRuOEuYbDoyGH2pI
WvkB7j53fdvj5StkiJPjQD18K5B6xs7MbCVgJrzlrd/0hqaKpy+QtHCaqZHX7vjv2PNBbqG/Ci6e
wnEdN64jtrgv4sBKm3p3YxaTUboHrfSbcJlS4TLDPiNSKT2qo7ZFozP6UXJ8lj8YElbPRuPrBPgV
vaglj4d8DWJB7NTofySy+WrctMOFoIQx8fi4AUTnKS5M7S09SlYjUB0niNlO+6VIvNXXaYa9T8Dm
nyRQDwSdGrCO7uzlIxQBCaU4yFjjob0l3miENF/k+EEIIMltq7nLt/yQLFqmo9rO9Jc0meT0NYko
s7ApYt9tk6brTohH+/Ecwc/+ZNQghutWhF7hlVvwQek/fJXjKl6cy2XwFv6js55pmwcHuBZTiImq
UcLB2atm0883gTSJ5cm/yGJWI1Gfm56M+gZeFjel555FDCSIn27aY8j6ESFh3+PvPGppO1B1WuIy
xP7WdNDfY6P9CfL7ZCHr+LLNK+Fnz1MHfGaT7wO1i9W2mWpBtDJicDvfJQntRejxrTdL4T2Jx2zy
s7572Chtd4cgam+lyB5Xe1fKT/baQlNkg5cntTJToxJElV9wSPszuV14aIGm5QH0LPN3r1wY3bvQ
KDuEbbRqBjSAP5qKwUd/pDsdkerzyOhOM0WAjSCdgIYqgNbjIDTHqJo9VTIqS5cHbHdaG4VMAmCA
8TU5LlyjsFnUL916NTDMdLkBRL6HS0P4sF7n8JyUNpDN11KlM89mxGxJ+AngacCu8BA8dxn6xKvZ
HC4tN3fxpOfEn8N7tmaKvBmbj5fzhV08eEnIUkcP9V1rCWnDTSTV0d76dn9BydChQYVARUp0fcgn
33PugngGh2Aw598r0Kh4tc20hTRjNk3DskRu/EXGPyq7XclZDDQtp60ZHRc4C70JjnRhP9QVmZDd
1o6XPwVTLFfI4HZVNsmm4y66tSZtklkyv6+Um4em84EMU32IGPNH9lsif1l1undgxj6NqfKEQ3ll
hexWzlaXig+OclzbUltynDFvkJmx4q+4jSeUVCflMJXZSdXSRw8ck8AhfjO6lJ2jSzR6TG2VMCJI
ZW1xwGaEHcorNmBpiHb35hfVSlvfjC3BaOPrNfilEpVx2a5EeXQdjAGbfuHkzuE11brCgqjKJzQ8
u5hoTYvd8+1wCIL+o+trWAZ4uc9JwSkpyB7KYd9A8nxzacBQj70kPJtUNrISToYmiFeUHVc7MBXb
/jFdCiHxTBMyw+EDnKUXXHS3RjCbBOmEruVMN/FthAPFDsntdp9+Whg5+n1/5OboTKKC6ZvPp0nE
sLNro8uz509HuGeF5jkBbXnFINWBHcs51HW/kjvXgU2QLZSP5I3D0qkEZsErkOMQHusEnf+RfAet
qI0CQjLTvbjudTjWfi68h4twZi8mhmhxcPOqtU64RoOOr8nAICHYk7dvzR2is7jWaM8wU5WfBkNa
A/TYrecX+aOwUZ546iohWjcKVEluXtF2eARpJJ4kmbU2u2o3xflhJRvvlzGngO5RWbJxqD7W5HlV
yW340i2+srUiXsFS8z/GOFKv4L8/N7qxPyw2z+USPFmLoggqb7CLnhUTVJD4a3RLUFqsB/N6hinp
6FL7tHnW85dUbROXybY94ygPZIgiRepoMB8HE2xeqToFWoll+Sw7R5nTIg4WwlSahxj7GUWMFT6H
0/Nr1FdXuyO2eIdh5SzpIXzEtYPmRxGVAH+jZN+v396+CKhg5VrvSeMbFfGA13e5xrxXLDniFCdd
Rfga7U8wSng0jKQAdsamK+o6q02awWANvaGRmDi96JNcxuXfmuPIzF7rf+Jo9BabKj1yz0SwE1nB
ZG136TNI73PIWepoNz57FBIv/U3WkQr0x13aWi4UwSc+HJGT97mGUC9D20To72MuaF9D/7HUpV9E
pB/TBBjSaD2cLOMMtcdqfgD7Q80nEuw5dX1PCo8Bxe6c9JLIgH18kO8nkOrg9fOcNMfhxWeF/E+f
L1zRvQ+rkZ5PmzgkMvi36x3U2fr/HE/zHhXuHhCtkYIy285L13cxQ0kmyg3MxXMOCWqBJx2sH07l
nQ3j12XWR+zxrirU0xrIwRaPM21w9GyQdOoV158xdtXlvh/gt+VIEw/2bL7Ydam66ctcIFKMGIqA
FrlgBgId2JZgjPFfN73eeiuZ/MVR+GYaq7YVN7NGU7ED0ZyIIjBrtQ3n8OytNZIYVPAxOVyhn1Q2
dfQmn3IczEc5Cfzxe/PZ7iBHofoZUMdSVK+ElNRqS6WDiTGHSt8WkmbdPDJ2eijuO51bpEDfcALJ
ebBzNeUdlGkCw25IF1E/EVv13y8/XjjCSXncCe9wRnRMhdWkOD2GbwcK2zxhNI6LY6i4N8UOj1TP
/3Fg56Hmko+bWe8JJK30EJ21XAXimSiH7FSuOC8FKfqhBGw4kSgSunG/7zWUrSpZJ1J40gDRLHF2
kJqQ/Yp+ovyxJteKF2HnrjhyCxQOV2vgsJcRR1UzYGvDPth1W2fNkukcq1QXyDgY1ngpg2qjwXMM
UaX/3CtBMv4Gy2bSr16/yWMccqZ7mUBgplqYdFFhjvOaizZGOHxLjKbtGAVtHBoQ2PkqW66n7tdc
EVWtRJtmcS4ocl3zrHkVzMVbRVMPT03awfHO7vt6l+zYjNHWjwS88zlISalinhH/xpTFIxlfYO8l
f45N29d3cn6qxMmjNDOFJl5/WF8fhrpccrzgpr0VMSHM5UZuQZfpTClyv+CBjtbPgOv/6643Ijhs
DTzomSoLVKwgSVfA3cmGo3MANdCbm0Cg3DscutI/61bwyDbQdrPSb7xgDEWFVMyJCxjU0xgOcMQH
DwrPvfnO4f7p7KTFBUSK95HHDG0HZly7l87YqPcmsTU3KoRhEj1iOB7Q4OLaYXUqGbZ3Cw1s48Ho
JTHOa552O3StBLMg9v14XLv4LTXNXLnISVIkyiTYVjn+B1xVfOZjpOz1gtN/z9rkdi92vJjCDa6p
FGgo9qDEtRlrR61RCkeVARZ9mobZEgaXMJxwpce0mi+W8q4mu2mXVBtfj5XBoP7c+4/iaNCmvWWT
GTSzOhAz5DmPJiv4P5vh2fzTz8WEKZ9kTBUK6gyre7wV793A9ugeA9WyHhIY+sDC1BSSWNAkTiuj
6+63rrsTom9y75+xEAvqowsXvOU39jJAUoh3JZvgrEFMU7G+PsrOLF415tq3x1uV8j1S0HM6Hv2M
rOfR+eqjylVFpAogyNLV84+eNkM2m0kJQlWeR4DQ2HxeH0OsGdB39IsnaMFF/Z0ViNO+JHu4hhU6
7fvIsDJpigZFPugXZ07xzv08IzR0x1Ou6SOjAgB/QxUrdN117sLd4HyA4NGY7dj+nDBTBwOls5ni
Ka5EUPC4LAdxI+gKiZsATN5mrbB2CY3q2dBzp3ocB1C+tU+ujEXYlLsV8QSlvwtWPvLhnihiAs/7
sDT3Gcdi0xl/pV+PeL1+jE5kuSWuVRnWeasVvHmm4RCa2U0fD9O4M4iMXXU7u6qOnYUsA9vg5rxG
o0EPShhINSvpJRycMqMni7y3psagnGk+8ksCJ0XTkE6E5jkb6RRAHq2ZVAEkXSfCNxMEHGCO8dSJ
pMnoXxluFyNfulVoPZkvhsbqeY7YdwRd0QXEaVmK2QVq+o5USPO/af/fR3iq/Zx95S3cCGYohNCY
lhk/1bG4eQ10CL1cSPplqIpP1314xH29K0C28Gxqq3cnwjxu5KwGI21SJ5uA4dG8MF+CLVz0M+Ma
JYUEby6/GtphPA4GXzjKoDpmtzw69MYSQsKMwO1aZlxYrcCzS5kiPyYOZR8Sbe1VCoiZ2yPPFoCh
zfq62x7Q3qy9ZRXG4dsHXsI/Ia5gXSYfM/PJ/maHJLZ/Yo0WtSro5rXOjxH8ta14V9T5+zXV3ZZE
4W5f0O+yTCLaT6fwh+mwQUk7LxVGjmIYqSQ6q416DI11VcX+GOTbYakuUu60urQf7MrABJ9uaZgF
C6ziHzSUHE7aWmzC9H5HpF2imcYf/y7qsNaY/iWuOyHnE3oLfJyIc698X/9bWlqsj2vYItG95eYq
n/kFMjH+yPdz4+B9S/LijDrJMM0KxnZKQnhBduB5aKcsIdCjyOSNrizzOX2bTZM9oYHJx0pAfrZZ
Ow/aSGD3N+VwxPoETs1jSkbicykep5hFx8bmryJwlK8fGcrYbfTA8yOKaD3Em7GY4BODihn1Uj5F
0G5z8+yuAejMO7X8iwHOWRsUwCeJ+DriBnZ6GRmh+5MfyLpOVVNzo/9btQj8LxreNrzMvODiuRVB
QIUOZ4tGCB8BJv/Tz2kWQdKJNy3t/X6jzuBXXuz8o2D8f0lnBrY8gnn4brsWU3+pmNzafcP7bZog
UnWqEjfFZweodtHPiWA3Wizhmt8wZNPc+SXCx5ilISH6yeeair85zBFEyZUTcZ8tDD8q8PZZsjfG
FZFDdEZ0l3IGXSuzydEJd/7oDnkx/4aPI91VyWi7ss9kB0VzRxav3Lcer8VDM75tuAXDjUvsL3vu
PTuA3MXUacIkhLeT2WhC7wsmgzolSDjLez63POuQI1CL5j79kUmHLXbnMc+Wo7axJN2CcMqfZ5Fe
xx8Ioq1tJo3Wc3Y3T5QGJXX+YuWZQrdQYvAxs9K38ZTVH/m16pjIfE0N+mVKJAS1aNAO5WcBrQeu
v+z3q2eCalEAPh7q+RMzFBrbzxc8fP8rAbLJkT2/ozb0HBIQdjVan39aqA7MsHLFh9Yt67+gVU0B
XT1JDv1JFZnUHh2I6JuSI05wtdqiU0N4ci0LKPVBJ4s0x7pmFpaJaLC4ow+YyBLW9vAC0ovOXQU6
h2keJCxjxojebT9FAOwYzwMBFGAH39UjfxwbAY7hptoEHe5Mlzh2JXxVHCcSaTYWEqr8KLFDbDsj
FMEFMGgDmweRRPa12jMi59MF1pVW/3Va9G/ENzzIeLIdFPZ9VxdnWYetrdx3vf2LCYNhiSrSgK66
9GNM4DoGMeJh4GzwKUw8w1dKTIgvXEgw6Uuwf1ucN7Cbqlb77l+s+MCawsz0N7PDQF0SJvhp/VQk
7+Bv8TMUYVyaFUH1gBymtFsRe9ztEmgwsFyxRgnyz7Kctpwzo8ZS6Z1li4jnpGWgl8fB5dBmhnUS
QmIjJ/RF8yCZtT9gN5IFjQr3z8Ot/ofu3f9mhzA37Kd1tRUTcsM9pwukOB7YyCRaVrohhQKn/Xt9
2eKOq+upwt9FIxLVJSMcZG9RQfUtKoQn2U2oz9QrInwhb2DH98URFVRiOLX8sQnEMaipRLCvyZ1e
nrLXZdojHnpsBi2RTWhNTRLT5Hf9BjxkZ7g1e/59ukRkwztxLhhthETVVa21LjgCWscRD6eC5bNL
UFpA7Jn7NrvA4BPx/QzYzN0h079OsZzjTFUE3dFR0fsOOdfNauiF8Y4HtW6qvqpbtL6Om5IOL555
19SsS9I3WSxebD59JyoGFI/xxnFNw9mhCIiyqV+gQ40cI3Gncwvbg+Xaehp6plHtCkiURgj6hINR
MiMdCb6rS2DKn/vpR8zM+KaCaTBZsm6kNxyi+s3+GxIT5jYTcZb8qNMn+nLC3j3hoVkx920M4eHT
eU1qgJ6QUUdbCY/oq60PwvmATZQrxBtKslCcBEttmOoZ1HymsDRU25YmaEjx4ChSp4clK3rMdMCP
oJsN8yOgDlmgTTBuRijstfAcVgUYJsBUH3hRKRm0qdNl8GRaC7Wb7jPkrFKO+cYPDknWNGgdY1+G
OkQsVZkK9tgbn+a0AW9bMKhB/u+2Ayp6b5HmkKi8NkE3AyUH6YET5wx8/VValf6n5JMf9cAVoIRm
JD9zvilM2zJvVMFgJpCOGpl6bAMT5hUGtwFCWeJ4YNKiqtFevQlZcwL38hXXI3owuSrqi7vN9hI2
3it2QcI6N8PorJv8/a1JRc75J6IZ3sO8+7GsUxbx8ayOu34hxN54GhIO0tC3h2W8SY+LC9VqBVvU
0mGC7a7LM8oSVFzPvt13uQhKLJ8q6QX2GYk/DV5kVDSeF8P2iCUzhW0nRH4lki9itQEykpnTTtL3
gDUIbU02p/sJgH/mvlI3B7pS8J0CZKtmUuXqxifldOhGxNm4wOYJKvxz8dlxztiXlD7I1CO+Kmci
TWcjeDrO9vN2K2ga3q93eoLEmU5ArcudK6je2Kp85SKPWlZoybJm8cl2wn77fpfR4d1PevNNnOt/
t3Y84Jr9gCmzEW3by4k+gZibJPgYXib5ieS7tolCQBiPlWc4no+Ij/Ua+87iMrIuBGMgh7XI5vF5
MxDX9PW5VmPw3KTvc0x7yPk49QVyZPRrmF6C+10RsnBQJUoQoII8dTsXy9NfArn1sc0vjw7F5urI
bvL9mzZ3F4qsoXavnjmTRAPKeJnyi4yEqbHg0+iMttPQPH7yk6SXy701nqVUcT15avTjTHtVtA2E
pbYUnhldPtcH15HfL2NkPatd9GollAxQz7LvtLIrUNiiHh3cq7BaGcsvDdCgUjgQdIVt2rmUCcuo
m+rx+evtDUTsOZZbRHwIFP6YHcLlx1m+iE2PYW/Fi6xjB12CHMh8yk0AI7szqPF6cwkne+ySjPiz
WxGmYon1K56GuQFxF7DtYIdsfui/2JneadR4tPyoFnjn6fZ9CmqMm849LkEg1xKsVsEnkWNi3G9R
VEngP6/CmdJaTCOxUYEHzS+Kf4b+2N5O3SMh/1c4lD7knEMViR5lWn0J9AB0smAcDPUbMwOVaIRG
qCGf90S6Q9GaBo/NRNypztX9sn04Hd7WMbBHtIrsccRAOA9JRP07rsgAZuB8qiOUcShlOm5u7z5k
vLtr9uvg1yzjvcRtBjEbMVy9rhjPHJtMpK3c0PgM7wB86lCR3So7flvEt0u3oKwFPCEHXrjUbbvh
4PHwEQ3xKnUK8rPinLZfjuJu5jvMhjN5k2lp46UFbO0VmuQ39VopRhdkLZDNg4ikCHzN8mIu2CI2
nyawBq+HFbLc81cREqcfyQ8ZGRU0PZ/WZlNPOIGfTj3liOXzvOarSFsoouZTm3pRBaUDBCu+ZPku
Gr1FpWp6aQ7ofGIHUA/EBH7dYRf44nFFeAKE/ZBXRVMxJoYr26dw6f6U0YVyM9KyFeCs2cs0tL0S
rxjxYvnRE0VkNg7OL1ZGAk9Tmi4DUAkVmZdvNkVniY8dOpyvbpfvHdFfDqrDyIYLw4g/+HTT3mAt
WtqqCjxJi+lgFQmuGVAPWEGdwfwljhzkrib1c9zQxnUhLYGivypp5ZXf48SRY24J4LiEL1Hj2y6/
rVYacmzSeOl1T4CCLemSPi1VjTqHP7jyzL/OUQceJ0ayogdBilK+oNoQbyTcKTlScGg0Vptsfw+r
sb8/beJBtCp1w3PmnghLhHZejoREjbUL/1cIcvuozXbfvpQ0APeHY+oxTAeHvN1irYSKVqweK7Xv
skuq2vGZqC724LDdnsseZ8vsw/Y1hKMEQ/95EdwelBGrAIbkA/XD1M8VnMrmqcEPaBkE03V1h5fQ
p2mC4M6aoyEmhoIOgKM6buZkmlKBd6M2XR43K1ejch8VV5Gs5+T30gCld7KN4Vtht2LCItZbkY4H
3SR3aC+6K/l9WtyVznr2B036T8r5TVi5/+od1xial5fXXU+hcZUuU5f7Q4OyQXbogz8EejOznThV
uzL0GTb8eDG+o1+UXv2LH9oH41+y8oqQSVpZ1WGgGrUkmFS4SdOsk82L1acIix4WlM3NCQHuMaRD
k9kDu5VtMI3vWTWa2b351j1RfXInMq9s2HOOqb5KqhHzuXXHAKXG5WTjkB+52dBfyvtjz7Quy8Ql
9H6PHS+dHq7tDjcS5J6+Cw2LSaY6q9OURP3mZX5ck05Ql8mkU2vKfaIEEGdqEo0MrCUVEDO3Msjp
x29oE5iTYaV/w898xBOXBRypyiEl/Ulw/WScxv/WRMxNsoaYqiuqgtVMTMm1dVZwOC2uapVf+/ve
8/qDG9PicsJ64A5v62ieBTztw4F8jDRtGrSvUdN09Nmvt2CLBVMa2giQwafPlvN8mHwqkNtQb9Fq
rxrja5Ttq+nG33Aby7qriU5Dce+NyhXfJclji1icYpSz8B1E5UvxeWSjSgKxR8XXcGTe/czlngM6
acWeLWt+ScD22oDE11UhIomtFNAFRr8EYC9Kru5KjTH6ttYdB/VxXaNBSg2e9FW0adiDwGSNnE7e
eRqub/7yKbibgTEJBdb/rlAN6WXwuC+DAYBgNNxnNiULKCQ1q4tmiCXb1tjCU54jRj5P/ZfxezSU
TsW4XhiQzEc9STniRHCBC5S3S09Vwjx2fgeScmFNQXuvT3jW1/N/duzBsp7K7Kyd+vCPv1M7b4lN
VGauOaECbU+sdWAKDOyY1fRgp0w91aOZcTT4dH/jh4vJ+F56uFiDJigmPG5A3UPAV4kF/A8AU9ff
DSnXSJxiUSv5G6pY5hfc3jN0hTxxn258g2bjNE+o/yfEypYl6Bbci888J8wt9lhdA/4bXsZLlzhf
5rJl4n0hWk/AjIx4qSJCFhLKg5IonZpY2FKWReytoszD0ZBjqGY/8I3e2vR/WYKuyiA4hKBdNg+0
uJZHVl+b6/5ASufqj++kXvZ9QMn/eHj8cAQu0PkeI5+SOTTFwuo2k21VvTllbb61e/hi4YYUoVtl
PYRxH4f/fWhGkS3x1DbR2eW+VR7zzRPwaRDynEhDOpcZb4k2kxbw4IVGDp6Aue3jlN+fJevf7FJA
MvbTkWdp9OE0zcZtYWI0RB7SnlpLn74iFR34WjocMUDJTG91MnYpeIkR1tleErxko7c4wDpNk1Nk
a9n18CJuuTfV8pryBg+uaBoyRz7PcTBAuBIKpWX0VTO8v7KZGQZSBjfRKATwsxZOtQa8sO4llmSz
m3CedtM0h6A0D3NFAqpGG3NOfxlfBQyn18tPNg8oTo7VPPh0QtHWMo66GZtwoZxGLg3Rt5KiMy3e
gyQwIjYtUC+YUQ6ftCOfZQPUQ901hdmX1BNbC++kbad+icPMdab2XTsVPpPK6Gi8JwHqyt/X7WIf
nRd7PA+OUDpOpO237VmSQH6g6C70DduCvG5/z/Q1WRCh1sQpe+09t+3IbhumUPC5yfB6bpLTMTOg
461gIyAIK16MhEQNHieOnjnh4D6iCpTSnfK9PrGClcLcIbguvEztpU6x//ngIRwIGSMbBCzFayKn
8vdcTJvckbUmgSWqmHXX+5YZNhY880zeMA0+7OgI/idl3I0e6pWkzh4SZ0eUe7HFTRBHAy4fOe4K
mRl4vG8s/w5VjIOErV9OCBTeYioZ1OzRmyh1pl7PNRVqY0k7OeWSLQgHqBce63o0BNm7oa0W2Sxk
E+S+rBf4/P6DuHcCNs5Er7Av/2xEN1cZlG22god16OctqOD4UeNQBk19AjgKNrkDSrTM+Cy3+lA0
3iF/CxIOrO5TJQXzBWcBJ+VW+F7MEV3xkhMArcK26cykSDbritj28z4XpgpBcOPSoHe0NTnyW8n3
nnjNS9SWAoDSqexGMcLvzja2tvnwYfLf/oSsrDFuupI9s0IQY/1EFfX+CWeIo/U3SE9xybm95aXf
98mFbD2K1HcEJ+d2KgmM0+410autIA66qHsoPpbmqYknpjYngKaoUzoTHVK3/RQv6d6AlusJcJ9t
k9QEoCOLZb3stFV/zP+4j9X14D5InR0Q8vlbaemLMf9F4h+NqoHaEmV/1cxdtdvPRphCAzU30ir1
q7OSiOa1en+IqvAqOjhvwKUSrHfyrhOTof5iP/gftFjZkPkJO+6EjmvzJ8edDBuY05wTTfYKeea1
pYSnDVwzyxpwFiNBpUCWe4jcJZ2CDegLGTcmD9H+3GYMopnjLjoGI7sBHjgYhbpWi0WXmm1NJAAy
kAJadjqSUDAFPfvEbUUK+B3EJ0SqU+NcBjngDmlaORPCWdw0TJj/4PCOX2f1UOcO/PwizBpERGGS
2Vz8Z4wSBPWJfdZAeXRBunCtu7kqbKmut5WZ2ZT7ol8clFTZdUR9ykQZ5uNyzTnS7WrGg5GIgJCY
pS9LUsLGzFIVEjpsYKW3uwp5AcG79hzWiRU9+9gREGoE36PdUkkqpwh0WahaAzOcCr0qZyFM7mkS
GownUeCdi9cvrliX+T3hhOdb/H/cTC3sHGSDhTMyMTKPxRflOpKhnB473QJwqF9GKRVAH0Z7SDTr
e17JKNCdUbIdQhSoCsrFSaparLwg1MDzlMcDFrI+Ns+wForxduKzkKN1yp2IlF72qRfuYuh+twMe
YaO2FMgvHEavU0T7VGegvgvvDS2HFl2GyAUHlsQVmoR29Na/b1xSQgJLXeEztqjQLecmFDQqPNzc
9D5YS0mxenuTd7duE/ERL9hoztceQutSSa7YMurp5P+mUiiJquD596T+drHWXPc1XF2Wcb2RQ1WT
XNJ0ESvU3YWZBzGHUPSDSvDu+RiL0aBBhLWuoajNSfzdUIZrXhHjJoVP/M8h4wc9cgh9J+c1Zfkc
sRnXCpGW4pGMUqcUNj5zgGsMooCInEbdFrPuKjJCRtlzWfLY6GtY499jVeJrrb9uQ5SDP+JM1Hms
Kj6Z4Zn30fyHVsR5U+UFvAwt28N/P4vceFqufFNxxZR9+VwTu5Fm0LDHRE//npwncGUDlyfBbDiP
d/McuOAklX4OaLLZGLJBzgSNr9IgnDgHBr72V2/BlD4ehYM52vBwioUEMbk5OS/CRpHlVWqlLe9C
kzSi+CaLW8DCeS5jkmeLyQUGBNO8JIX8K/AtNlx3YtL2NBXQbgAQ+BMuJ6ybNowyJ6X37pSiIftm
bFeMZMaiPp5/oVSXoDF6iuavah83xxJo5l+BxaBuLuwRBOnZNqmte4lBdpeZVc/GKwbTteRgZwYC
oQn5STvD+qOaDj8hNW+ZDhgbd8isRNbEFe2WYJfGoJvYikFcZ1eTGttoXkO5lniheLhNDl+2qjx2
tvY71yLrMhMN/lu/lHMqWHL18eVnrDYW9f6Vd+EqxTKX6JHDuXzsdaRT/TQTz2Fk94kiixV2c9lf
CiI3wQEM/a69NPupGZVyAwaDf7P/a+mRzcGxdm1bY/EbRcoq/BEWAw47SUmnzRsUDEncjp3VhEXR
MQ3fAQa43qKICD6e5S1LsiKXnkqZMittUc/C+pewbFj+T5gjhX4pNn3ebbiTLzUrVRbsjQkpJKdk
pMIbHoLOwtwuMGr8JqiO7+RC7aM0xWjYVz5msixhlFi+ZVQNQbE8a+janBu14nzyTN8rzDezP2Rv
x1r6l3TaMCBBDwwsimaJ/2gUGSEIvZqbi+8+SV9uNDZGQ8zZ1IOJsm5/+vm/DYw2sse72+pC+87G
HEROemjQ0dLPgbji89YPPAJ3kD6i1+d/M4g6q11btGn1BE+5rUl9IXHJjioEo59no3Li1AAtORmK
TENIwk4gZZeadhvtJgvl14iMK84CM9ibnHcxHr+h5fz/ZNVVmVUJeD+fmgtxe3Sb8M5Zh1Wa37I6
R9QM8eWAdS/mhu8jN5x1ntzyFtasXxFG0Wdq5OJE2ohwur/9jxkw7a2zmHdPIQoRBSr2+/nTpS2V
MNQKxc8wdbEJQjgwFpiLFe0xeeOox3/tx3J4IN8TRTY03Q0T4l/FcDJda3p4wPwpqqszJ2bWp00Z
OI8e4E3PKqZte+79B2WfiakPgvvEpNtcl4DWA7toSI+KL37m8y7XPN8o+tB/LEtvDHY5tvf1kYd5
nnawyUYYucPi6N16buNh1488HU4RT4nwKzks2heP5qLN5/OLhnDjiueRw9Xl18IaQOKkMVtVQ9L2
ChSpdc6sith+5P1LwBJKEfvsmPNF5vDN+7NBqmqr/LbVeuVNxp0/Bkl5J224eXtPaEdYVxQs/qfr
hf21v+oFBtz02duAV2V0F8AyuplmVa4F7iym8LScL3oAnumBwyTsF82Q5SxpdCGUw/WWIlpEzrUN
95GVtErjLr99NYNv8DcEa9n9FB4T3qZyrtN/qtNjG6+rsXYEMiF5doYcFOOAn7I9JJBG5ChG7IoN
rwXaEMfOf4fg199K9FADkkxQ9wEXjQRt+hFryM4ohrq5XmoOlyo1B1HDGCgoGfm0v1lvkpCfUXMX
AjYOgyZG3FGPWrkU5mmbVLhaPu1vvt/DYscQawufpn77oiv8YcdisNLLvtZk2LZAIunRSJKXokhe
XMMahPIGMZ8pOnppHMNLJO7nhliRnfQ7PrXjEN306L15bYbVMY+C3tXPY4uCNKQ/CDTDnkYLbrFc
N5iqSoHdpO3wXzLWO6Ka+dBSWqPItgt/p3IlNiGEqOmQEh9HSGhSphmHNUAfxDo5QYO2Rhmy14mW
8Kd2n/M86IY55Q2bk8EbBI0npiOSIfhCltiK5OIjJqeryphB16wJkGkk+ozLunBsNK8TflXOXIxl
JEHAqvqUW4p0ebQoAtQAoU84UyI8YY2Ht5kIdVD7WNWsfAxS1tFeig0QvsB5ilXLzBloE5kkqlwT
mPKo2nvNRGzggmIJC0eqX0T6hABvC+7CNzOt8EJjRNWAfy/6yt47+D18ebvlmUV8wSYaUyOBq6PC
yl30jEMSHFo3ft0x54ZZ3YPtOEr9B+F8hpRoZrxebAs9u7Xlx00I94lBVkjXdz55imlzKbkxpjX6
b0gYP4Byvvu51YSgPf0pTDWsx69MdLeRbtoclu34Cx4wglCYxLalt06NcVXxYv6mQodNqPRsCN2w
2nF9Xw5yNtxyR/xZtXoIU/kt3TRAUuJJ7jPsGaaHp+hxDU3oo4EVY2mA7mnHJleFnOtppTQeLi2U
U7XMf1Wy67Jgsg4rmB2IP9CUrHZQwFSOig9Vsy8xpSucI5UMsU4Mq48gZ6FdeM6WTzr7cRZZA5db
U7EOObgg/LVlZN3hP5cDYMOTfOiKpogs9B1Dtu6yYQvGfcazRh9SceYPDGgSO7BRukiAS9HWNme9
i21tFiaWmscl5m1boFITuYyIqbgbyImyzdHwYU8ksl2P5o1UvidrYkGBKhZJ2sUqnNxO13zIuFq5
ZqHDLkZXrSwVcmQCirCvhVDbEnwG4WWg/5aBelkhAvSLMmJxhZ0lsuQFw04UkgWREzS6017GQBhh
z4A/E7Ca0WdWJcgz6uN02VQyfPcQrhPEWDg3h8rC+9Gv1b+xZMbG3oAFTxqILH7TXNie3Foq3Ys6
QWYfWdQtX7SD1FrczX/YKX6uBcMWWgSIRRb2l5gYvkIgnieqO/OslDmT36Z/0uJDP0oTESX87epD
VcVA1gVbkMFvuaZ85lIPx+yQHU12zUIr6ksscuQ+8iAvxpOrrZYT3z57zn1GerKYzrTujiU9shMf
cuvsdkiusY8+5zkmi5IrPnk1wWWsqcHTS7/0I8K6qEBciqMvyS36dcI2vI/I23Xo+8A7Ii5CJArh
xkFRPG8W76Wcv+9oMKc0QDFVpS8dBHHh8JxFfjoni6l0awpRsm+927NTKivAbosiRoBYdD+Ae8fL
tlbu+uaxS67Nn1Yrfm+C9bjhS/Y4EFi8vFdJrGpgzHUxALY+sU3ERSjaCMFdFmqPZIY74Z9LlzPN
PAQhLkzxz+/tQLFQ99R/y0GbVcaEpONZo2hN+8xaNR0JaULnXt9S1IQ2YbIk8Cyb+fU941szQ9Lw
kMvfs4Q3RRyfJXsjX5cIkXDZPHCQwYnnEVaHKUwNYpOXzTHMJ9N2njsqfa4SPhuy8UXmq47ZPEbB
6Ea7ynwJWzzaKiQ5yakAH6DRJ1HiE+CBww46aUXE9sV5YZjQwt7ZrbCFSKzLd/TB7qoEQ2TMTn1E
Mt9ryckHVnlytwIR6rrYYTH2A5CyYR4gdT5bIRhLKa1Am2uzXXCWBRCy/GWaOWpYRZ0XxlrWk2ed
1aBAl7XlTWb3NAM8NyP/cNYTmBKAtiScBXVYHdn/ZH2eIEhfCtsdeyvS/p2KTka6zhZKWzlXL6sx
gXzsMj5GzpMYou8XTuL9Vdca1AZIE3tljlyq9Niiya4AzyRGXTGsv1s3eWNh+65UgrMBylUe2PEn
CRw6Pf9WS6X0xgR9jTgskVwZv7fI+ZBmPpHAXcBnbEostYY6/+grCtQFzNfbE12iZOAFbMrywmj9
79tZawOievDWp9kcFRyrAU4oWAMqCgxSM0T3TgvNLJQ++HVL6+izhEeuBAOjt7XQQEhvmYRsQnT5
qbGPVKU/yxEFQn4wGZbs5CWDbzoHe1cPO4GHv/wJ86aUTT7G7KUc+VK8lr6ZCt60oNPDOrHUZnr6
EGxS6t8KyAf5+kcs9RGGckiD5e53oJbQaOWjy0K4QUj+HnX8xD0PnoLT8Wkr6ceYgGOsnBNG2GJM
JmlbwAxWcRckWCXtW+hKw6VpykhQIHFil3AjGxZLa09ewdAj/2pEysYYYWW3WryMHvv3nFB0ztBn
5Yr2Eo4lK4hotUxueYEPLpzG7aOJklHnCT1aIIX5pkEg+EBqnYrPkpRroyvEUMLazfZI6npYbee5
HzT+e4l/ipvMU2PYT1KYNzTbrTRCuRFmJXER6oGh6/BpPy9oCQuWZZxt5cASma9apOTqFLYIQ3ZA
ykx2TI/3Jnn/HZACfswz+gB8PjAnE9aTiLkEfIcdj7ESs9DMP5vBaEDfK7rIK5+Nax+cQrRL+Jiv
UzlsndGOjfXlEdXScU/r+Ue1EooIgq/Q82DF4xF5j/4epXeYeDrxSIiMmGTfEE2DVCJSxHz48uif
zg1MvA2QK0ARjtmqQeLoHYzj5VPvTCW7sl+ulEI3osj0Zj4vW7a7DI3+r0+/yjw1nC9Zbuc7oIKV
MM3EXFOhZFKGlpgHdgsMAEjm/hz//lOsof+8DRMbQzqbR0vSKWdIE/FHEMbqDLWBBnTVEI2jk51J
z6nKVyFVwDftdsTImaZ/qp4NYaksfcegGDIGHEvzuCSfrudEEgazWlkcowgm0yncdrXgC1cSsR4X
HUXSTZWpz42cMwaag4r91ynQTg49qFbdwhLHUJHiZ5VIkDJ2yStgO7mOrnMMTv/jbDjwnZzfhbwf
Hm4dWAJbgwZa6324+gSSRr8suKjJVN3+0i1Q24m6MZNBRXvO8EzW+DXOlMyQr0896PxbRrOCeax+
As676AsvT2UndU18vIiowT9Edfg97sCSw58O8YJNOrlcjmzYeWBZ0aF6cnzd/iS73VbSzjBdRQDt
1YR8TKdr2ONw6YXmEXTGRw2u5xLoFC+oIpiPfL1yrjn2C2eo3BCs46rl/UcK7IhlOC0iTMNlPgd4
LEWHlAKxLCXWqn9TI18veHTApLDYTe45WKemsKm+Csx9cByxiXjP7WDfkFUX6dF32nl1dL2QbVU5
YVkx9s24tImD1wf55NI+VCaj9/d2eR/MWUWs/XAEuyoC2IidTsms+zaKAH5EqgcfdVi8bTQPqMfp
XRyvVyLU+ptqLsSOU0GSNYeFwpN92UJSE/xMi/meIqf4Bx/wr9nM1T50VcDTTOjZPFJYHHKHw5I+
R6w4S7Q2b47pfQFxztzPk1vG98ohgOVvhTvWMDIf5ghFY4MZyx81J2yqvzqihd4q3UjupWNnuoWy
Feb3pBEP0QnJhMllNPaxzBVmLONlbiCvP2/Vj96LNUCt3CfRQco4dnu/wEgIYhlfb7S0lCE/LIES
Sunzt0wnyYILX0AG/OGVsilXies61vuo1HN6sYN2KF5a6yMyWreFuAaIOHFT9d7D5GKgb7QZPEAj
jxA/RK0tGtNltH4WVWTJjFoF92QbilcMDUxHahYqxcBLtfSOx0XupHesdyBZeqdY/0ak1RZACUKu
dcizvWmVdLKWNfRuI9K8XToCDzkZn2efs0osSrVx+wlwe1UTg+WoT7VyR5bqBegsjtJOxHIATUvI
bHIkxg8wlbQpjpjJTMNpHCV/R575jY6IUYQBaLIZMA9v34oZKcmI++jMJvl5hT+NyXlh7M5m1via
wMa0OIIW0a5/em2rfNaHpJtrzZLY1yHH7Xy6/HD018TjnAzr8++cUiWBe5O1vPmMWvEd9iPLorbP
pyK3BcD+boJ4q0FCyXQZZdMt69JCd5nXZyWEEBv8aU2tk2nwGGh2Pc88Z+ZZwPirKx/bBiZq2NqW
FiOYDPHgliI5vBgd1y6l2f7iXUdwE75FeH3rlQ1+ryPFh0hdwsp3SBv5wiLUze6jltaG4hkSzznZ
aUkHLV3B8H6MNhy6DkcoN/3Wj2U4TSrfSaEKxDq7TQBYJ9ylzcGaZ9+dYXdHqrPrBhBvqpSSII+7
ZtgIIGGxagIqr3juDbe6NpgYslD1KqmuswB3JvHTyvmfnwTzPAzT08KsNaMBT8uScE951dp2SmXq
4JBVcQFtetdZjg0CVpM+TBOVxF42s9WlJBC/lsNrYfZ1iRTEvqyAob7L3Ei/RegWNahNNa4FKO5N
6EHW9HVS7dE/xo8SdCs9+xb/8f81zPvLE5pau9BhWiIdNqIoeLzHi+e8ZeRqGnsAp8NfFrYtVpgu
5S1mbbpkjNgtb4Zwv180Y0exmUutkVM2LIsBq1C6r3upGQhBj01HmHZcn4wEy9oVAQsDxUIE6wnZ
A1KUVi+ytAj1M0FruE/Vl6XCTaU+dsm03xe7NnRqkShVFK4j0jhU/W4ewWBPPqg+htlzmSwaVHt7
UqCHvgzUclPb4kRjHD87UEauC5xlPfnw3HNAhiZ291HFPzNUWjL9d5fdbTxahbzAYwabWRL+/X7n
1sDrQq7ibd2/7I3H7wJfznATdSyyt6H5IW/zSQlafLgVdXG/dkS+mLQCzPTzNi3CvriOQOniZ50n
BIoowyxP8YGJNrh3pAyZWuLDNIEfRD87G4tepeSHxGxSPlVK9QuVhDex/5txAmQ5+a1Jl0NyTLnj
WSRVInIB9GnMAoTS/CqDfvF1Zoka9jLhD+wGZiJBsmxidHTvLliuGtuic9I7HRTrhuxosx1LTSo7
/9KOLt8XFr7hPtsQMfo5jhu6dKrZwAh5WtoPZL53Jgr2uxhmNaRvfKmhsNtANZL17x2TcurQlcV0
mOLlcCxTnvC7rRuPfhf6zntD40qbEmr4Muy94KbEYsWMOecBTxw0LebnKXL4jNZvtqVClRpGQLoy
ePJcPU28CfrmwSf2M62bhhSu8mLWl41++zav5+z1VYqoGa0oxg2vZ65tkA4g+TQS57RLmdcJgeYu
NzW10u7CJgvX3t7vPyHTJ9M1TIhPRorpozBzBATlO//i6XvGoYPTB0wGlCVJUKrG+OaCtAbCTcbL
CtGbmYSFv2N5SUZeGsYKxtlIux2j0nFKRBZ5sbqGFmKOq70fnHsOGI+QheDHTzXWfncR618pWzCX
rE0mThF3NVd3FT7SUZQhDPRa+ID06fpyKC7nGj45OmMJfuDiansIlhL1Qzi2yTaRuPWjSa17EL6e
Mx9js1pU5t3v1irVBeTlioX4FTcTOXnzEpZu8uRTOHJNnEsa8q8LVFAWIQcTW6z+TU+ho790CH8b
W6LnphjJtr64w1m7H287/1PRcV93PvAEkeIlqDJtGCIlYfc5X/GqHRWNrqj4dvD3QQ0ood01rZ21
5Lqq+dUbeU7Lxx9dT34xejEjkTDwHvv1pIay1fM3Ga0k4p0RS/n84AU9dEEg+rwYuIxYiCZnVT7r
E/092UxSBvLkAbK4zb1zPAKqqtBYmTNhpzc4pbeTPHKWqABienLRO4Dn8wL5TgDDQYYLKCGKCl7c
ZTR4URbcBSl7UU9TaWBDhUhl/NrRNadOGftkYhqCDWSPZkpXmWKUNh33bJN4SZwNIyLOEjHZ2LH6
xKcbqykFfpvN17AtOcAs6QSqvJs4v9ZipiB+TfUqeRT1G0zTPYqog1ArOviqdIjbLVD7wa5kOo4D
Du0NC4uwkATvee7Frfc/a12BVAkavzEf0iaB7Qox6rICibaMpWN8k0OgsQKBCFt3C7w011R82rDt
CMFb4qrk9mXB9AY75dMa5xaZY0620uVWZ5o0oX+/duApikK7j8QD6iHtZf23G+zzQUIHFQBz0eLF
3DDSXebwaC63ZOfjr/NvdwrQWYipwrC7lIAHQWafXKHlyAilj5id7oJ4QHFg6CVlo49QuOsC5Aym
9P6B+aCGSHCMbgMmq42BFXI4/GrIpSvEEcRab+YNM5C0LrzTIFOLwOC3B9oVKe/LgN+H1izPVvCc
IDr+SDf9VF/fp3/Irg1sOawDWLOaxfoyKTOxZTe1Ze0QlsVgc/avmExUQlvTrCOCUvJfrdLIGenW
CEK4zvka10bv0Kt8YLJuANxF/+cT4KIxpBd6mrYCSvTW7643L8feoFs4Y1oJZcJP/wPm+exBO9x8
9V3bmxdxixm3K3oFLvPP7AmEgDkPzrQXYNwypi/smYIaYBkeQgUbAdtl/BBhPXy3TLKuwP+UY4kI
g9ryyaKpkLTsEs+Sz9YdNp+RRP7OzvE1QtaXCwukIyQ8U/ajJhGHJurwkdBpOc79FVtX8a0UbFLz
kHq7/6XpKSuYSad458GE8mf+j4jaz1vScIpxLQsklcrx4kSnQaX06oXdKsUVCyLY8AEapt+rHwCs
/M7pQnnKR3EbCwSxIGdjtGMl9e72TDc1VveI9+7QOsCwVkaPR508BogxVe83rryX7Gxb7ktJsaDp
h4ibFYbLALFUTeDu4rS+g55Fj3X44WBIptYL0zYRVrV+8OEoXi5A7PFDtwC5pZyG6QPf/xZFwgWI
oJ5jLbWSoIDS2LXuEZoRe5qZ12EigIbj56qUhhL17HXlIhSDzZEtYtoY4kj0ZbhI0fzDFCSogDa6
m7tk+TzFZ+4u+r2eh9T8YRxs9zWCM6PxZL9H4QPWvWiuZHKVm8/QCyT0MydVllLm5hOfAv4Co60Q
8sY77+zk1SzxSsLoWBRC1Kl5xbK4gXDxDS3iwHIi+P3iOJ7DJmb8yRWCFaCDVumlaVaE1mJMqnKi
6oBnd+LsH7qxqIsHNbuoO09sJnwtUOUyWq18gr6+BigO+NmCOoAEr3q0KGFage08nvMdNb4UqEWz
O/dme1PLmdk4GoELX1fAdw3btmr+LGCx+fDOI3c73FHokzBDffBJpl9W96D2r3jhp2aXCMzDiCjn
NJs5z24fCCAElS8+BFSzeL9x7Am05cGd8TzeWfl5rceCBXlXBawlHRALMooF8qX2G+FjCZ4cpB0D
mrDjHbuGqPlsWGgCs2idTtkK9GDtqVawP26GjgSHLrDTUJGUC520ZTaGgnkNYcgxqPKmG/HIBtIG
wUeiL+88+r2kWIXoTkuJCXizw+/wUtGbVkA2DZV+WvWAeyKMsH2+6k9NTyiyonasq46YdrVJakMV
RGlW9QmSvrnJqt9uTeKh/AkNaQP9Or0UVQLofL6MahOkS1BLzHs0Vx64RD3ah9Nvqc6507x5Cr8q
NcsQ6iXaJ5Zr51leQnxiZpt3logp9Jkn5vcwaXrNjiDsTHPnPV6aNXb8D4pX/3A3po0bNvqIXP7e
Ia2Wd3NAKQ4btua8tAZIjDc5aIOzu+AkO8satbZLGOgs4NTTyatO1YVd1PPFeGFqb/goARf2ncj9
VylyZBM2swaRtqDNhWIRkEm88/2i7j13TCpxhvw/LeZsYtPgmG84Gvb20PbyOQuTy3GkPIeNmUbp
mbf7e2XhI6Gb7RKdF+L1aA33bdnPZ6BVICsa+af9fVWqEhNDtKgnc6sKUwq5j+GJvyy7dnfWwesO
s49rVPdl7Zu9pJ2R/+lMsFq1KcuIQaU97FSQUDamS9PjAmL/LpRqwp8Gg9BuPSTxCfA1iGN/sDZ2
olZ3Hi7GGo3uxJzrRxVeqLNv+cInPr1Hl+cXBx6vJyioUBxTu+9vIHP8wuugmT4gQRQySta+LDlB
ocu/yfnsjfrshyeQ8vjGynnS50tCkNQu2dIGMUNfi+d1wXV1rlEYPHn0h/HMfzZBhBRRaqhUTWPA
x/atJpQPZLY9oWOTGjTVp4EdQAI6XMRJ2lt3c9b6hMc/L2QtBBdSNnI4RHrRZtxOqIJdNCKTVvVi
WtJMCUpQkdRclazAyaC9ItJgrjH3DwDBCLMkUfimq9RUFtwxFau5PtfxSRWOs44NS9jwt5dRNrti
GKk7ZZpol4oVeHzOpeCwcvyDF5pue50vm9r8s8KNSxSWK6cgA/UYL9ZuKrfh8EFHhPeQiMQUi8Zf
vGqRFfCdf0oflDQ2VbCayzLJLZU52qOZ4lKe9NuJ6jlKwTuIX5Db7KKnEBm9juTBoYycC7NSAxgw
4JntUFhVa2Gsvftil7++78BeBcEdPzDutlqj0czlSOJIQEZ3n1GBJzY0Slzj1nLJAx9ooG8m5ltM
J1us+S2xuiGNtLYl9bldjP3k+tJiYvN8Bncs0s8DzSWcal/pOt4+ML7MGpcKIkRwvnHMISZQqk7H
7CaevLcHzo8duE7UFcjUirXfCfAIXZwLCUhtEanizP0xTpNTnYOxuy9B02nujFTvf2N29NMVOcWa
vyqGM8IY2jAHJCmg53NRM/JLRPvYfjiZFwx9csvDJA3Boo6GN+73nOLmXaDBkltPGeFIIfk9kZAC
GU+CvXvKrBbT7vqEQYA4gAOWia7yEYvrJUaxqP/eLI5drn932tWl+TB4SZX9eqiKypp3p+HFhasp
TT42KwB8r2eeHE6P43644vxp8xv4MvThDAxdEeIqxG2dc9/NLhvVrnxHjkbiBN2TnPLU24OyPk7l
euFo8xsKRRQE0wafuJrtZtMCM9+tSQrNSN9sdfFov1ZDRi8SAZzRG3SNOZHGYbeFoNUIC6IX0qDr
xLs1sKmZHQsKdIceRSszTchzlynhk3/VPwkRmPh67snPI5H5VZyer1P0aVm/CBGxTAlCRwEw/xOO
r3lsTSCwh/eCYcVMVFaahxNvkJOVerm3IYzker7/VtJj5vhyt58QeyN1dNsUacSOBpJbEe+Rv/UJ
O2yFB02XR1idi4B8yY7FS3SEdvxdCBsRtix7n1i6FzuhiYu9gu68+q8A5ldk6kMMcNE49KOPLa0e
7bAzKoBW/oB942U18wfwcFQS/dSo40hFzlcXq5R4rh5PgDRbVESt7EOjHLhVhtOODFbh+sbKm0CV
rlXzp4dpoDwWRYeMK5uaui/CWXewnT2QXZvef2y2p61JfkSbnSOeM9baXIsDAPME2lYQkLBpVSYB
1C1/+KSt58v3qIkca0qbNjWCzUVgA48srAI1w3gFpeqBm+sFL+CUE0xLfANIil260epStDMTdRfH
jFshVulYCF9PkEYTvTFj7eTCS4hq86dC1Jy+Mo0g88cCabPC0knA6kwA4+DVUW8zxv6x3sw4f0rc
3+jzVqflPAk67mQfh272FI85x6vLJRkoNmsbQd1XdEfLjm+9+Y6Iv9ns3TmlsSn5+vw6xt9Hz5Yl
GaQkSDTxtx92GcNmT35pLgDW8oJvVlkWJQllnKqAcAHffBU/dmv49UKnq/gX/vkAeKn9D1G1at9q
9uuYHoDnDUlwVJlADD6J9qF69BULPfdwmI0rWKKATGNq0fW0kM1GrVYa1HhQFhWf9htZ+7WU5Rae
j7syWgsf2efUyXz0z/NH4aQrTzREev8OjqE6EPPgnX2iichG5cdKVUSMEfYDR7MQL0Y+ZGbIWZ3i
bc6wTkl9gc7hSPenCxbCAKqkZlpLswJUwBGPXCRQbsZzrsK58PetjXunMcUQ14zfDMhU0Ny8zLLO
+XNh0BjehKS3bJkk7XWBmJjmaYYdlDibdwehhE98rD8UxJoSHdwovNQ7QFdJnNnRxqIoPZ0hnLCZ
sK921Xbn1h6pN+PjjO//X5tMr96+Y0+uYn0GjwTNtApPKBJL71Y7/pyzkkZX2FJ4bsTAEP62Omdv
s9vqk/c6lRMrvC9hdysz9jax1r0spkTBP6hZG00+cKv7J+S6RzQwESjigXbRd9XVaeTYuAAObQTn
u2rcQd3m5zHQakJFBzjglpqv6P+NX3NOWyXI99mLXddk+Eygwo0NYTEaMNvrJItumJpxjC0nYoAB
AoFrNJ6J8sUuF5dK96aLYO28YU4LKiCtJI1CXs1hn4GRDmfiHemCN12U3Xv5qmrnNEPninLwsPK5
Oh81Hl0QozpDAXFm4pQFqM7236Xbk8dpVneI90WHOwtwq4qcHE0phVcP0Ax5iEjsvg1ih1AYeFIV
9u+ArLN6ejpim7z/1q7k5w3W6b0IjyoDXFAAJ8rwmZ2J3aYaR91uLKX4/J6NLYAufHyJDcpr2iOv
7C+8khNBxfOEMxUPdSak5ITbFa2d+wckwWFAJ92tbls2xalv019R2tuQI0YOEp5m1A2AmpqR0Zz6
FhmEcRBNxgoOwFqO011qIuBlybVOuZzV2LIqZJoFv5zhtD1Eu//tiNPcSUKISqS7wsPikMUuhE80
N11jpPybHDApwQ0eHKiuUUlSNdIonXNnekmLJ+O2RlRKjFGS+zYkVt7C0GQU/cs4OKQdqiZWlkxO
58ffUIwHj8E0TYKVR5QF2b7aV6pUxY4kP/q0Bz1RUqSi8Xna61kbSgd7ap+UOEnx5HOnIVnNwtm2
vl3Z/hoQ//44Csqrm9a3GGKWz8ayIShzsIJc71CCgdmyNG0uDS80Smnqho3+csJ6I4GlFIi+Wv0T
heNEQf+FZycl3eebtitvIyVYgHudTShidi8ADXzXN1Ej6Z5PhnQXf4J/jv7Wsl/4ilZK0st9PtSt
gJxxGD/VfNAg3H/qj3gNCunbn/GEWk/6famDMjRAVlJxnl6gLaSjk03YOXwGZT+PlZLUq/eLAB5E
ZAjprJC6sHgzxtmMokmFDvK90aTqO1oMGU4AgwNxyGJQ7Q9z0Par4WZocD2Cqegp075RU/1LBdsM
gLPdmHVhl1Ur4f8AOd5AuXE/PnYLQywNrtf5eAE6f/TeHFqA9qS0LDDiyO7GYIh0qbZVXYb48BI1
FjIpZv5nt3rppZfTlRQDwLSon37vjO+gbAGsxZJx4LF02w8kbeKk4fKV/E7acUpSo87+ZcO73lRv
CRio44F3Ridm3I2jiwB/KkvBDtEVoVCetN2hLzq6lnyoRDHjmvglTGuBerpWKhds5jc1k0KMt6Vl
lPNMeWR6mKuR78ws/xp/UQtrYNk9707JteCabpvvRG6IUTw+E840bIewbA13zIEXTmLXprzwxmBj
Le5tPcBnPJzztqLSDNxaEd2kkNNii02wrLrjqNU9rdAe/qeIcIGXNo5ITjGXwRjWH7a+XC3nK7Xd
sikm2o6g0wiz7ETfoR5CTAmCv/T91vXp3ZsBKY94rQ/8B6qUx0muWuYpdsusPnQsG832Sn8RSKA8
RG3D0kpeIDs+zJQTyBY9HjdElzZyllNj+0v913yUadZcIO96UZyKYuANCq9xzzBsrAd+GRxK65b5
iRNxH+rhtvxskiMfsu7MTQw+QSEODmSufOIopIq3Ar+Tg8RffNCMjHS6jglEjbfYC3bx+RFYLpjj
tAbzdkxqsEjb/s9t6Ukyz08in7axzmFByC+vngZDPHsJ3768SE2drEHiJkyXeaHG0mvRadJ8GtSK
N9wiCEqnuNccji+Kjg2A5hNyZza7gm5bY0Q3iBGot5iqi/cl+m55meOrDoIAlC3fs6yaxQlnlo7k
x8Ivw+4zZJBvtdDKGci5BV5zCIzeNCpYCqvV90A7ncvXhor6xgqW8P0Z40wi0rOdsg56BQruU3aW
Jt+J9yaKUGONJAja21ftYfc+fE2G3HuL2vB2IrchMOxqrYUFnXLv1XdIGXNOoGlF3QtxkPJAy4MA
rxYoJwUKMa9pjbkQFQolbuVgShrfXZ0R/0z/bIfraeIxDXSXlwazqQ78pTLZ2q6t0AYLPeGm6gKs
Te5tUwq5WaSPHAjKjseyeHp2vLQfDEEmcs99KRAVTEOvHAK1YH5VFEnJj0R3XvO5O0N7howjisNi
WKWAfT+e7n9KC8mikdmWYlaG7jWMiKqkQWhdfjVIyAFJdDMq8qTPK5nOHN4Iootqs0hBgITEIkJL
6pCUM9WiLLLHhYa5UV4JS7xyxFzJKsReFnapLGtOn850MckkbfwPorPNngjr1BxaTEl/9I1Barj0
Qo+cfYrZJBDGpaoIYRv0gNsQC8Gm6CY5qhxKVkJkzNuITnvdK+EusbhdmAkYTzwyI1Osf1vqNe7I
8sbYTg9PFnVmNg574Cs3MnVTY2GRjWjqnfRPiBXdoLggauedT1Sq/LbQLXT+DIKWsircSDt/wDtQ
uTk2W89Woj5x2Bfo0CStE7pLGJQVWtR+z5X+Lupq6GngKbO5j1EqTMcAP6xXGZ9w0EdU0sK4ZTBB
pu4u3A+NeGN9uNfuQ6CZlyoQiq4qRSM2q8NRigJj9IZ1UPAeW9zqmVkejmCkK6QOMX2i1LwSwYeE
dqO5sFslRRNJIl0vlsNQ19GurOTqwPfbGugP7UmD6rhVfj6syAaIy+3CswmqJv5nMBk2i5LKYnc1
bWtR9kUHf7YFnHUMeTSwvlYqVNpawaoQfhj6JvlhyzcHbxEg09+0Xj/KXu4pEbv7isIlnIEIX5gi
pFffhevIkHsxVToaQsokOEvAGoVD0N+zZDvtddCJQpNEMwvWEe1JwbRFyDRKTne9cfAJjzDBvdgp
qSRzNNBbQVIphANuGcZR9vn4cZe3mpp484makiE9YC0t6v+7ISZUP3WJWOC2vfS/yGkbW3VQLAQ/
WHPVXcaxXpRAizNiiHv9IVPW/XdK4o3NnYc1qH3JKrxM3kgvIpu62RAeDT6XvbcaMr5cKvUpm7+x
Hk5Byp5nxdoygBA0pAsfLFJ3ivC5C5aybLpaHJRcDoWA7yllF6idc83WVOGEYBQ1lPae5CRcPgHu
yHkLhQalJX6X8CmGlPwp9MyyEZNMf/ADIVGRvv3IJsewapPKzz70Rsfpurmglw+gPi+sGHi5xxZ+
4eO5gmuf86vJMGBlkl4VRs7dKtRg7ywGXW+rT0VrJrHG5puUhwpUX2WkwwYwu1MfQVatnq17rzGk
IEhyTqCf17Oip2+IygyqMqSNj/uHLbC4Xc2BKNFhgM1toP9GJ6bgOxlUCrpkI8sWwNxk9+9vXBg4
Tae5ratkfkNtFwQodil8Y8tmUvGdTG875G2dxPk9K6vPMqgggye3mxFECkbKpDJ08RGcvQyBPg3X
TztzGq7Y/S7ffvM3FdxHt+u2NlOqwmDq2c9rTbGWa9TPvumgd2a+An4w10Q9iyLCoqr2YvA2MDtN
rxiXghWXe/IzIpqEn5SDH33h7/YHAdpzSojKVOgM9m3SWM54rO+THgrXPdygeapo90SNme3mK1wZ
7cxRs13qikk27oPpmYWdb+NW1FfYdBJFhpjxCzDtu3LRLob/tFa9r2p4VeVglF0+iRA4BwS7Xcz6
oUdFBaj1zF0Jgn3li+sJzMhN3Np3vkB0MN5Fq5rlscvXsmFfXk+HxJUMzU0k27A6Jd0WNu2UjOEB
miKWbDSFugXD3/hz5tlN2X/TRETiokfw1HrOCQf51GzHTmg6ZHI57v4fECYShhZJJD2nUOlEF+8B
EGwDfyMNqh2NWXFsWIPTwqFoTUVVbS5JRg8gXN755AyY1wM9cJCZcV+9APTzSBw84w/Hcb5T6G8b
hF0q1f4TyLpznUz6mGU0OV3MITryjYyIdtdz2sCPSc65r2m4Z27IsUcslsABbtVfb6gOG2LvVBXf
1aOLkTJ5JFvr4RpXPtRAbbjO+zhHcR8WuDJQR2kBHg6rQgMxm7FrMq6qARe3NiGfN5EKKNkA1nFY
2Vgwbr0GnHEE4WH8A8/UaGg+YpeicJ11uVNcg4y434A8ok6Bv6lz8d4JuFqLmjAIXeeOW186Io/N
er9+i/Y3Kfz1bMKVn2w3NjO+lK2dwiLrKfHRwwKF6WMiXCCQNyGSEZsyfv7lwRZ6jkC4TC+uJQT+
YhYw48yUoCgReYvE/qr0LJuBGe3i7Nx46w17u/LwcvmvdQ7AhrVfnJc/o1lyUqw4rjvvxqAmgiPn
xdVtgffeHL62N3CK/PxPn9YmMqUnoCUz5AXe7P5WdycKOexdHG9vsbdiBQwil1CPv6m0NuKM8B7V
2n2/Lz8n4MyFkK5B7///87U9I2n3hek1hkY3zlkGnzBWqXKcyFjEJ3EB8Dz1FwTRk8oye0tK8Yg9
Npo3m+yHUhzhe4RXfkI37/4irTi6P4bAQAsiTSi2We0m/YLt9UMWEMzhVydoPKK4KDDDVpDlk4R9
KGqhYVMGozhfK4yBDqIw/PZkWHDJ1gpxhCozuupmQm/8/+2jlrBU9amHgFLZK/0xj5K8JvAB4a98
Ja31Ueg9RYApBR8LtesRXuXNLgnXbeT0DO22//W9uynFXWFDhvGlaU839h8ZkImlGA0thNFxIoL4
PlWXK3bwj+m1Il6ZPrcAQbHrvE/XfQhK7rDkwysc2ENAIrmu1PE6EGQ1sIzVO1zuB8cvTjDxEEbN
15SXwRRprDhs2e9VcMoPyW+OFwpBM32i6t++yYaoIsBdVk+vsUHXq3xnWhF51NnluXbQYM4qcnxe
EFJd51D/6p3HuqZOolbZh76zN/9wnFTZEv0dEMeqzdSUnqDJZk4JfAL6C0HS43M89bwK+fgyXwwY
qKO27k8Gpq3PGvLyDgQfSD7oFKds6LsgwBIWun1xKnxwDHa5+2nE4tkPxHedcUcfJTLVNgvfbCEl
A+THiVOQhli0SBDG1WscVqFzb65brhrJV989uKcyCFJug2kyKZAlThAxjqYpiYN0C41VuazA47X3
hUYZcar4t7Z5+5kcbWtdwG14PUX7cB+tNOMRM8rxkrv3bl6GHX2Qu9LJ5cYX3cv8uhqflYURQ3xE
rnjEIEtpTlSmfhObZeOAoe6IHXKsf+sJL7pLq98IKOOziKIKMAs6AeqKGAXw6gYYvFvsgac1pEl/
y5Ekzxkvs7MnQEoPYDRb4+3I19NlTI/hSlB4+Aq31JjWqNydqTRtoWOCtTp7BsqfTlQAr15ye4yd
0U6OSw5OVmQsUR9/vlmvXdvVNSP0OdWqKgyJplIEirfrx5YY6Opnp/euNL3R/qncG7L2JC26rpyv
9qPC7DbB5F3f7xUuqkDJMANqHo1Arg162BPGO7T/p5iy9GBP11iTSbbG3ePXyNA7FfY8C9sjhJU4
FqZd+HH0HIKlVhdR73pxcqURdFhEs4nTlC01qxkpw+F8/lXDD3QCyFUMTtWgLG4yirEiYXflbpsm
soG5iQcnw03whiUf233mh4G1xZFmmasTkCvkAMyQ6cy+7g681yxv+cEdxZ+DHrXBytdgVDncU9Da
9ZUeyNGAjjhL23VzSOH21nEKW9CDNFcafPFttqT0FofxeQUMZDyiK7xNNiOC+T3S91MmZaNtKAFN
TW9k2LZEIpa4JlwtNWDFwByt1wDWUPd0h/iZHOUJpEGvg2x5N54BvzS0glIcRBDIJUEKxw1Vmmk4
DxDXYIU+kVJVc4fWOVQIRP/b6AyeQRl12xBY9OZza1AhXFct3s8i63h1RnP3CnSTxWs/XT3S5cn4
CV92V3l4IUOo8MDgiOJk+j0otTBDjx0JgT+ZBlnGHaY7vmg4FCLhkvfG598YUb+83nu+k7J4QnII
1jiH95PvE3wXOwXs6ddOHRnVNOtttmWJ9ADqmocNR0jorp6cVABIDuy1LT0lPVLFVeKcLCBuytr/
OT/r0J2flma4EaaSq+TFFDgxcxvEnOK2pdfLHQp7hbHKx0xqVMyD0ulMdkOS3uKTjFLunJdM8T4+
7aqpgSotIF1ArTFEWam0/J7yYE4toRBcVTS7kdRgcXnxRXPguUiq7/bJn+bXR/DELo5m5ZA/rjg7
FQACKGA4G6CW7O9iAoLZYNJEWxXmn4bYrcmz0kLARbvPRvLqsu3sM79qYqQCipym/9u7AdVnDpnS
N5JJI5Jffcx0IWsdUiHBY31Hu7hyZjWe/DPqcaI32dlbYnJ9dpIT/E5E/xtw3LEDXeVidorP/vWz
twER/xYnrwym+ZLeFMUfljEiMc6rGRut4IauAkOISLfhvkg1JVG3DSWPE8qI1atcTE0ENaBhLa/f
tjiEdS0uA7GvHpL93w/5DI+ePqktvmHIVkpF5pQP0QtDXRi4n+HYLYVsqEzEUU3pD3aZhtKXybq/
PQEV3P9zXj2gz/wCg9wooM7wNfeGdpTcQ1vUVUMqv/7kIR4F8kIT6Kpo+YSt3HKPhedgVw+xiYc9
gru4QUrGTaAQvJcHVnTJqyOvlERi7POG9QyYEJTD0KZzKn8H5gCYEsUJPKQKUtcz4PB13G1ONgTi
ff9NYYBgRx9qhJv5EEnyn8y7yMJHkX/MgRjKKnWhaaZPdHMnILWujyjoXVd2cq4uJ4Mu0rD1wJpb
YsaDpQOKA0mZ9VxoOFZ65foOkBew39+2mCR8u2gUWrPJrV2H5GHtSj6694ctshmETGx6I/0V2DU9
8ZOzu5JaGi0dbob4XKvF/i0AFGREYRzygDdQPgVceLCTGVS9ALJxyRq0q8TDEqaPa4pFmsSbFIQ+
WXNzW4erBTAo1CzAg+vxzA/IW5Qt+iuJZ/rrvgrdhJtv1QHfQ9eHZfYXeA6rKT6exwoFosxMgHjF
KqdzA2YCiGKdv4QK8o3N6x+DL6XrEB7JvvamgwRnG9aL2VNtrHbHCj5+C2XBWw6fKsy0tg3FDcoP
KP+U6yraG8/WfzO6JOcgW/KGTJLPyCj/eS700LWLF85rI8/KzOCDgHvWAV5QT27G2tawyaHJ4nNZ
umMrBfOvxkZZdcc849ZUUDM+8nye0vXTM4Wd6XDyxJ3T2rY3x3XJGfcilKQbeN0riJ+1Tel3nkoD
3fOQcnKVkI/Ctpvcm9UI5KN1c5mStlac/vspW+beECn/DZj19l/Cp7InhBmek0BKEjtVa7Nzr5ZD
TadbddLGHHkBeMZPF2dio+GADF6aAjTVx9ZMw2H9VJzX7TcX4hkCSRX3L+WmDdiO4ymH8eg1vwlX
Sc6GSQK3NdU6X6E/ONoJzLdrgKtrUDuJCHK2+QdUJIWiQ58X7Ou1JxauTPsdPy74Sf31wbqHgQAn
arRndRzNXSy5Y9mC3Ed/JfNERLeVBkCsCwLvMJbRiSvSeUR2hhIGarw4GCkbiLyn9ZWfXuvQjVxX
/fj8UX2u/KwlGKZgf2mCkRZyaa3hdzz92aASmxCp211WwRmYfm2R1ZVTp3klOvb3/gUGiKT4jJ0q
BbTqMvVC0gERCXERn24fxpXIBHZpMVpEZ8Uzi5piXl9u3RCSg96H97/AUV7kL9VIanWwBh20zxIu
ExNGcA7TKm93aN66ztLMoSc0REnEUlLG/AhgIWeQl6snDjBbADZRKlb7r9oyJAN4jG0LHpnqBkbH
yYFZO5OjGqshHI4nkJd2tgSz88n1JLw5CsjpV3kSpIrG5snshqIr1nc4L5IzuZoJssub3cw0rQa7
DuIj1VVAzJVYQ0ejt+QpvpbM7qASW0q7NUVPiwzW38v18tu23osVMXg1VPaDLmFLCxX8PdwS8Dzd
OeSV1a+N1/4+SB2PXBh/PvvvITxaPIwJiGQx5d9y7imS/jaMXqUbn7UycEq0zL3K7+IBu9HLxwm5
hlkUPEG0OkyV2i7kc92LZ2II+KqOMkP6rnGbkJKASN2A99jLtFiznrJ0T2uN4Z8AeCCa56y3zLLW
PfNTpGNW2DaCT8IHOysRE32CzLjQ8Nf7R2xWvY5W27l4dMhMeu25GuK21/6QFJOE2RInvs0AdDOw
wHw6iblvCWVfXAQ4K32NkgQXaI6KB6ws1o8KHhXAmkgOLiJO/l4+VM9TH9ZjFG6b6HcMILcL94Kw
PvJ1J1k+dacLivMxCK76jSy9pntaLU0VOYnAdy1ydM9BxttirywWtKEs3c6j8KKf7N1hvzxurPV/
Fd/6Ufzx0eneU1K2LGxAadsld1i15DynpGh3rjt8osxAWFj+WjpwkSTZf+EM45CF61FmtojYu7jd
3S9HElU2V1hWyw3SEqOnzrDwDqz8kmPWBMmduALYbOeMJ+z+BgOQmBIVFaXNcsFuh72W6lH00eDw
yGmxO3vNRzHLQTtkWURWfoLJ/fIulPrsvMpYOnoOOSQt8aanYfG5976eiNOHoFMzVY24WNKL6dGa
7rPOs2ZeB67IW+8Oow1LXL18t9yNo9QLEhSuRYbY+8kHaYrwhIBV7uCZ7VwXj1WOSFWdCYlcjWc7
BzOYaHagTkg3Z2xEkc8k2Iklw9yXMtxCYSe1/vIqJK/O9IOIe+BgoVnKxGVAF1Narwt2Gw/AHtUn
SKwDDW7CKF88ZE7j9c0v8FcUmQq0WsJtvVa07N7j8glHnOvsm7yx8J/1K2ABXuqUIBSu5yIghS2k
MqhIEZzgk4Q5knkAuBMCDDAWNVTlKPMSuflOALNcZsMYxm20YEon13xRO4P6SvKZd5703FtMrpMg
JOX+w0+aY7HFMLiHaEX2Qo0UVBH7l28MnaXGhqSnOdYrxV2W94RwB52Dgjb0O05yYCEZfhGcj+Dm
Y/ueK7sSHzj/2TZOqiRiNtyugC5t3EKoqnCvoQ0T3Nmc5hPXk/FhhOHvLt9bNgu26MFDtTcRPauL
HF3QFH5mXEAY55lpwYQ9vzz3hQXC9BDHmzxMzBnFaEYKjpdeulyRJssPWSGjZgceVAtTTF7XA78G
KLOT3KxDe11v+K3/kA2Gtdwk9deRZLoSuNHrGBxS5+MF2EJ7pK8azSO0mCMN017URwWzeB1Wn3gg
XOXDUFPlWNrB+m46/0gghPHovro6vrc1Ipcgx5POZe/mGmPAIdFkzJqJjVvT89EBtRmBFxAvq6Q/
wxeUh5uAXYG34c2rHTfSgOhbW0SBL6TeKhAcMaL961bJfPyaEjrvKIccT3GcRHBzPqpfJt+F5Gm2
DCMxYmu181ypa2HNB6FdEautWNj6OCVggORq2MMzSTqOQcjNPkeLdPB7OuLY09Q7YZES2w6cWiyZ
NCi1qlr8wmQXg1cO5d7DxZDQ0JrmgUPVYaPy336OvvVAgQx1I2owDqPKZyfZr0ojZgWKIAq18/aj
KoZ0VIplSrQYaKteEPnkRR89m9r9N1MPFK3YeVSvz0zM2SHWMHiGepcO1ar0H0dx/bgUyL02Hc2t
l035guF7fCxBlxzH6/n9vIHtKT9Ud3Og4JdZwIUmKiX25d2BytmDAz6J12syG+ce1gIBETUL1g25
pmHbtkengeGwB5no2yDrMQ6scyZ//pkMeWeaP+TeYA6yH9jgjItukLAUzJruP/xC2eSHK+ZcS3gw
IBjNNZom1xlELvU1ba7V9lL3mk5FZNfBW6n1W0nUOWHxGgGRDAkddu+2fO3+huSsHDqdnF+axqsp
9uaibepK4Yyf/0QryLwemC3Ubf0JhPQZHbDXz1AgPnoIdlHrUcRQMLOJ3gnyEhnVBcTN9LnBL+9p
i3A5EEyzuEBNKUtRXYiLEXq6hlWuMckq0oNP4lzGRElOWIpVIQDuGTO9vDdlhXSEdRd74rw04/sW
0iVgrCOw3jxoO8uBMEdYX306KV8zeLxWJOdKXlENBckS29RIGDfWAfwhZRX7U1wvAUO9uADtG89y
s6loO39xE1EYFoKyOpW4SQZp5krKuBfME5jlAuL0oKaTcZ4W6RGGk9FjH2d+WEcGZRHegwJZG7+Z
BRp7oMZPCBDeMsS7KiW6/+roFYaXh5WwE8RKBJb3k7X1iHFEbfVmUtyf+A4Pjgb8E3fjbcowazLN
whgd1tvbunHq8NQFYaiWa0YfU+uVd/QB70q5FAtRfAlj3v5YHKZSyy8cTN8Ieq6u+MfrmUSf4rml
B91UiSk2vmheEyxzi+FUYmAcEBRRskDuvXlka6tYOzTR7g/PLMuMJV0tm3perQnzsCwoxl3kHz7U
Z1MSqxutxtuH+eumOHNPtB3lAZ0NfJwpf2ms9GyVlU7miXsXys6WZQo90n758FIQeZgor8fmTLOM
3opQdkpuFI+okH7MlXKJZ3lehbuUUiN7eNaf7WnnSnTE1k9acfdkmgPZdQeE3i+hc76UO5w+col6
cEn4MuQ7leVFCbGrdwcddfzVFO5yzK69Rql7o3DSZD8WXpCD3P20Xv/KF6hVg7agegrGKOB4xJdB
U1hY2G2nP1lmZ+K9Moh4floY4CI9UQYvAWa/8DNVxelUq4kW6lOD/dlhEkMJLXxMTNg58KfErf2b
J4ezBgL3odUm2qPJHWigja4ISiIwe4cUagZHbCCvGXWsAOLiKfiZwNLuUtpm4sTTGj8ssSrVtpOD
/qScTkFeuW1Vx3mD1vnTiFiE66w1E66nbn1FoTHjf9lFUPiD7aPuIIyJ1mxbj//BdVot8st+VD6U
jZxWhCcnsnqVGZ8zJpDvzUm0/BhMdz9ELwiYm10RCslxc4WdRRbtcKZVA55AxQSmhsjrs1Bix4FN
xpkIOqObMYL9W0+54HPIe/7mm5tAu6tbFsx51LlUzFGwjd1dBCzHwwDlN9yZXFAsz5jZaK0CYAsl
4yCuxjpgR+0pD9H4tZx9x6OpcFXBC1GfOzFV/tFEov1v82zXgL7/rcWDYDgth6pnVbp8o8PhK8MY
7/Nk/y6QlbjXSisu+VJGRBDPonaqAPC9Mp43HtYJz3xzfEX6w/IVN8ecRWuXUDgGzB956jgyGb2+
E1fetMe3OYtD8c213FLDqt67Z0e6As67CMvqusPHwDbMQeLpz4T989hwsH3+VtWEC0izYCbJM9Yh
90omwT3YBliDik1Gpax9Nk83KCv+6M0e/C6rILuu+2asbHs2xBI6KylRAcEsWWNY9YfyJt2OAicJ
fVtB97DxWr6cCpDGmxuK9C5CZ5toPCstM0+eXryMTSB0hhe7BNS4osig4bmUv5+xgZE7GA9IehxF
/pHXybjF4SfgEU7QNMmhehJpG9uNtqvrqYc64MNbDRmxtWj8arfqmTs0VhE0qm9TlqL7dzTAlo2T
1vCnwfJrrk8i6cFuGp/MNC3IXZO6MHBlBkuDriMmsD3feAHztd1F+PIjqeEl8V6vxGps1O6sHrwa
aSjVK/2KI+zMiXX0bB2S37KB/iDK0AdAo+dbgGm80HI1hq6NZejmSaMwyOc+1BJy5EhQpgX2x9rv
Pb9a2Gg0RfA84g2XlqQe0b/WfX1WGaWOdadXA2VQ3hHAquguJtFebviSzIQNV2ixSFdsG6je1PPl
IF/FYbBiUlgBhhppMFqA+X4RQ2I3z145M9pS2y8nZn5bQH3NFh3kSVDxYmyM+Z35LGlQoLIH89LF
MezVua5aqLUzIEAnijJHkF88IhglnQ027ckm/HgvmfWgAxzMJHyulzStY0L4rh0lUNf1TriytHMg
xM+8MPcltmspeahleXA4UxjbJg0J4MDvIiheIGO/BzTUewgTsZ+d9s8fDtm7eWuN4LxroM+fhE+I
xkYyaY+P9jvO9k47cAtpIX0HLcZ+EIPrOb/+mb/ODkI0wyPSHVNzfd4fptMCZ1rHp0Dr65STnl4h
ZNdzeHjEOATSydAauwgxUs8btPBpfUy9XS4Ja9Tlnr7QuDTe5vSuvJ7T55wPsmQeHeHCFN0Tov13
g7c6LDhwbYJPt6e6TDEUqAWOBR8W2wIR2nGYg7kwuUsCUv95kfJzaxrByJP+A3ZqD7Q5H5m+9xHY
l6FagOpfDUfzTrDIT5bVPyt9LHM0cgGS9NJiHYF4nPdz6MfdRlc+JBpq89YyGY12LMQhzjsqrThH
h4xag+wzOrud0oApwjv+/R3i9i52QSFN8RgfasN9ZkzogssVwNQ3rDNETOlCS4vKKJq5oNDpa+sT
Z7VWmCmWxuulTvM+jnLUGVfT6QrXW1UlrRTubu9JZt+Mm6ltkrSv24/JbYCqjdRwI9QLk611ct3k
yO5ex0I/14+HLrL5kgW1CCbylXqEoMoL2P157nBUlKm6cIHcyVoe5NGOr5rt0Htn9etF4F78CjD2
K9VefgH4oHyDZwKPtAhTvtXHgmtGw1z6mYCK3RF6im4JOkBvntNFOdO8a1sZ3EB1/NSWPBRKdbCg
x1bDjvWWxJ/z4AO5SK5iXSOyiQxAs/CorHVfmci6TXQshwRR0dCNLtefrVjjA0lj2kdESNxabaYp
vjwQcWbc6EqKLgksX861guufC84+KUtB4xx/cwI9Fne6MuJ8yEuGtR09dqtVQgcl98EwmvbmfKDp
GtpBXz52AVPuZ5DS3zKzg6RlGyf6rTxTjWsju5Mt1drAkuz3Kw2PQtQcu/BdcNdFsBWE+kLphedo
iHGuKJqr0oDzTZSXzu7i7kxqz1KxVQwPHt5n11oNdabaTNRZK2cGjgLS1eNltMBrUlsxuhHnrCEx
kUeEb8qvLQKxs5NLep9cdRev7CplxiXFRAP4irMxpWSzzplrN93GHS33eBNHtH6mAoQbWVuqFlF6
Q/wIVb2kEOE2Tk0E72hf0hHNWiYYx33omHyeZlH6m6dY2YvAGR1DyjD+Hrq6VpVK07cucFX/CUNa
momsqNztKntQm+Mzdr3kNDs+JK+uYd5eOTAI5NOZzTg829Vjwv2+IB0aRiGhC44QDTMiirXvaNCP
t+OwW1agKlXGyU25t/7W2Ep1q9cJ8yOMPxI8PgxcY8pYmlKMplhbHuz7MB1uJV3XgGzMYgHmy2Uh
AQbZxjKjA20dmGpiQAZiF1r28IlqHtF193idnUNG8GmJvzyjzrxd3WFNHvRvH8hoKpGJ53Tr26zT
gqyAQw8Vx+2BiZKXygNLFHEmI4e7Ww1se8Z3/5g5hNF/Pex0w1vVutOb+HuTwh0xUAetceN+zG3g
Q6QIcIsdMlBLuZHcLxDG7SFUUl2yuDE/ODE1QRHjQuDaCDxneNlCBlAlHdocRFl7t5Q7+RqCtwO2
S2ACobz8soMBKYT2rlA5b8LowieDs/+rL362PN17xJz1b5Wifi7Xl96ZMRnErfpEZ6/1obWccoZR
ehZPAh/TwIl4BoWLaXNTfQwDItmUwQxRHrtEPsQLep4bC9dsdIN89Rlq45OCgEuhczCKeCws6L25
Wy8zUqpSi+J/E2UO9rSMnFEijYFoh6UX69aiDnO5ok0tT/QV4G7shf4j6jVf7B6mXIjtyuraM7A+
P8C9w3SoRWh6UpsaV8Mws8Ow3UCyETEu8dONwEUwr74pFnKU4hA3Hy42b9FQHdYIgyyzx6N96gky
PsLk1BFVIxKptl6vk+j93QQgYTyTh6a9cIVNiymd6ktwcxHCT59iBRre6+SrwkP2ofBRfzjtF683
9BXuV0I7QCxjtQrv663WbT3BfgrQv51tCYDREMKYGoRcPifpBWAGGYj+MNJNQ0+Rv7ytA33V4gCo
EAIzbMOITtaPr9brDJBbo+dy9SbZpkvLXETEdDIXX4l85N2NEEo83Nkb3cFaXJtoThFYQ0Aexdcm
ne5bmnitvFX/JtbFInTO7MJX9YA0SvQLUSedyBtAJktivil0IrKLSF705lYtfryhQcNeXdJ9YTEC
jd7nv4lkz1VXTJ0nEus8FaWQJcEGlYNGIbsekJcUeFJorvef4bXDmPtlUOeVunArxgi6rIL+dRXv
nNJN6ffMskiWvkPGIP9aDTRX0Pl8mGLsJs3e5AEoEFF50q1E11fJLXPEcI4KnofLAyJRkWjDkbNQ
fNA2G/SoHdj+mO0FgofpPDgcGhQoA7VAAH67fi2pAb4lDLdGvXURaSK3O5dpvvPmEL5iRvoP1cnb
58/j1P2wuXRHsmwAzrve2+DiJ1W3pe/e5lz5ZvYF1z5lKH4wLVCTp3HkEKPwH1AVVOAx3pdmuc0H
emQgiBFiAGhVIPUo7kr0y3CXDWt7BUjy7heSzVwa7NrIxgt93cUz+77tbBty//30B7wMC13ORbNK
+FGBftI0hECf8xcLJztMbgq7vtx9weJkgPkHbVFIUDorMcbWC2dguxkb0Qsvnd5zEeZyrv0i8nNE
RQRpgrQRWs6YJ2d3+JQhexzHZcyxFeQYQ3jbfwqb3VnQ+4rhPOSawVYX/LbYfCJEnoxYNXI1Zqsd
tYpgcwu6LBBvWNVjrScMOE9ZcqPOpABhR78sOHRLdhwfd8GGBvyDdQjzar0/JQ2YMo5HbD0sB8ga
SR8umsi2sCMkcb8epi4VIeR39kPjMHeeet9TsaPFDvknENvTsNhBy4YLjIIpNFUPfOlh769os0ub
q6h36wKtaEsW1qWjRWFs2xwhYbS+vgLX7Kj4Ntye4fwH4TvA1iBJBOAll6WUmt/iepHZRTdUW/n1
JGvigw2JxfFLvJo8Ofy5EeEcbqVAs77k+BQpzVdT9JWJi1O0SGsmi76H9ihWB8P6mYbArup/SU4u
t8IRHWfOwv6grzzvfBNiIMgzR2xkt4Uq9K+5WlbLPVp55TIsmuSHLoEpKWHCy8EQIvCbSMiC+YL0
NN9gULmQWyT5iMz7+5XTQjLEdtOQQm7vUZUmJVzZnChPpZCxL5w+aotDMExZoeATKNpG9KYafgVK
68ncMZErpNx9QnVKydPobsSHbWujEoV3Cq5Bjc2ki3oNBOPa65yKOs5djgZ0/5SOqSXfYWu3AKnX
AvTt/fQUl+370lA1HTQawDGwoJCwvCk75Avd6cv5AuaQT379QzFYoV4zdT5aX7gE231X82TKTR25
3tJIoLs/qPTvQtoEZTgKjmjzbHMBqEP6tTOIo9dLJ9cQCiesryx0yN61UWpLCelAvy9X6j2yPlRt
uh46l+HSLIZEdvVi9v2sCLXj2tj3nANXk01mu1ir/jtU6rcXTmhzE5wnumkneb0OULGFerdxjnmg
+ov9nwc4ZUsHK3arWoR8ZiG2WZYXdshCIy6RATIwIoOYR+aeB6JG47kZPJcDenrvKcAw7anEV2Ua
uZCJTHhXXzlOAQ3caCj/b7khbFJ9kC4aAGxNPxpPQ3vIT49uppR5C3Q9VCwwK0gJ64iP0R1BduHF
MsA/5/SFZaG+HbWSKGdA5pVTGMh0OX+0XdiBab1lYK1E90quwmDwdr7mySMvryQIHHalUguUPC8l
eoF1NLUfXOG2m5NUGZefkOKwxW7inhZ5sdj3094oCtjJr4NPfDrgs+76OQZFLQAt0ys0QV2uRnZf
lP0C3HVLnS3k5zBD4eIhnRAOviu2I99k9O7NUwItO8RHoIy/S2CazboEQpPeTl6vSoBmxqeXxzWt
+t2BlB7KGA3Ek5ltVQ0jeM+IHmCpoMQJJC1PzRsDQuemlMnCGvXNHvuoarLAT31g/PkhwLF/TzF2
qHX9a03etpMX7U7ImkPr20nWmqPwGtQWn5kzdj618L1jUtKV8zovAxsejm5ZKsTkAL4iP9oKHuEi
/BoFiDf541Udgf2V+Q/XBC976CPb/948Q6hbJsdKSyJDqHT2s1OnZyztca4AsRMooZvjmy6j1ed2
F+z8ljvkj6tRT9dJeT+/x+eJT7wOLPcXIrbP/rJjRn6a4nXZNdJfj+XrA2mudGY6HLM+yHNPZj/J
66cBSW5PxodN4FXkkzaKMnHY43pQFAiMJdXYgmL6xcOiG9GkA1glt+9oYL2lb56WtAPNB4TSGZ/i
9F3UihAaSNOXielPWEBa6aD4aBYsDeohg51ttgSoEGU1hNvHndUf6xjgUcePI1B0JzcTtA4gYhPL
XSVSPdg6uhxxQtMzq+T7bPGqgQn40gaTyUINELf3B9CmJqbLm3zPPn/yB8ahKxEALR5XQfzy8bxV
+MjR/C+NMp+AtL0FNOjqlQYFScpo0SxTLrcYt+dbzlcE3TzrTSBLkFVkd0DIhK2t8qVedICIXavi
Tu4LMXgozJId2UhCxKjkOAybol7O1EGwphJtV8bDaptFA4dnWh/rAKHzOh0iRZ2v5HwULLgyfUcv
qym7S/c/n+XJPKdNK2RrdlEILQYtFwvqJwdV+0Vi+H0uWFGUKDkf15r496QJBXs22FSx/x0T/4ec
je2rmhZTQY+qbeBKFo/7TEdk7WA0Hb8j+m2z6iHgZcA0VcwZ9DxoFWnC/OZjJOz19zqZNBbXWAfh
qVw6mReyBB3yxNkltARZIe/rrSZybKXxL+BTUema53f4YqVOywVQgSW7QVbOA79avAO6le7XlY1D
SGu4SDYm2jKxmAHaEpFOaEdGEQbjCKwpSAfahYM+G4Tzc/QiYU1lmKLWZonENnYzmOtQz2ouKTcO
Oop+J8NNMhiH8u8A/7YSVrRXr+ivf2a3QirIRCk4CbM9z3UzjphPNK4yFYfeEI6CvxDjhNI/Trqj
K9f6i+m+/57NSfCuVjH2T22gVf683/DgSIAbWrVK+cuP+DR6q6es/udT8hUZsdR82Ei0aEuzjBYH
8mCUHRo1mk3aGexJjSMA4z60nbSpJlGioBmfpxoxon4M0ZoW/LL9jJ0TS5eXDQ4ZPGqT7U1fSIUX
9zzeYVEuGSV0xTaqO6r2mcYL10wMPHWYZlyC573H9tJpDWPKQFTTyaYO+i3hZ8j4bWi1cK5o2N1O
RXrsfwGAcCGELm1GZttuZVvX3OF+4UetRncsE9apJoHxHp9OCu9RwRwwwrAK20e/lgmxwoixOvrp
WljH8dlHpKePCU8SVGI3wVE07ySdGL8hQiiL/XAAwmG52INUu/sBRIO03MDee/G6cyUYde7LeXLr
9fekf2q5xwHC7wE2fMd07sLpIB9k7e4qM7tserTlLszRWgvLPbmuhwmEgKwS0yhrfbFYHhUd5vUI
Fgdn4N7oNNnWN1OO8DzBuw5Dn7ELfg5VuszChEr8lyrHn50YdgOOeiNd8SD7WwoVG57+1y05eIQT
1vdIiSrAhk4k5zKJbHihF0FqaHGO2oJR2sN++3fXVdeSe4jCtYJljr6efigA/RqOuayWjUfAH4J2
TNUSyy8IzVnuYLQXvgqov5FrfTQE2mYn28shKKbu8pQZ8HHmE1IV4aRdYKzKU8fdNoadrTD+0KJ/
0617BM1Ai5IWy+eTAwVQGLNcFvegNroDOPA3poXje2pkX/db+irQkizvJAE3KPro5Gn8gzIf1UTV
2Tcibxh6UyZ/JTgeGOawQ8UNxH0Mq3VAJ59S2K8WUmskFQ98OZfEsT8V5voFZ8U6pk6Hai0E8LKQ
gSf4E60CWQlspndmpX59UXC2DSgzhNCxtSrzSTSPxVlCw1S9Dd3o4r9uL/a4/XaJaWT57oMl79we
f/KYscGqiO1wadcIOmen2nWWqKfgi/9vJUGhJ/4v/DcsEno7wbM70Omvz6LE0p0GXKmgGZ9LXjGq
3yBEoIO92cyeCTsVOtUEuApLd/ab+4EOJ2OyiDUN+fPgbQDG4ioWkfHjBDtYRRBO94djUtFhQ0yo
iABursku1rrmsz2pNVYctGVKMvk5dYk0wsrEFy+x+yicoZNhK0XjtS6Y8T6oVHJctujOm24JEapB
ZgvjLcZ/+9ce9baBhh/NqAIlmrfCJBPcDpMd/DMTNVfoH5cCFMWPr48a+LU70Rr1Pz1ltihlwz4t
14599lBknhuULWFfKdLjapXyhMfRe++Yj62dDkoVJ05ILWrVWkmWzZKo31C43AoStNIdtCHRBsjv
j4choyLH2V0F6Z7NsUY3mXQTMHkTGqa6lzliQR9lO4cwwkgvJ7X7Flsd7frzOSsBKgEMTjE8PLBQ
W+l0Wb5xG2L9sRJ+m5+U2xKSUf/qYl8EUHRrgp9HSZwAxbJzbpwfWkO0gNfDFbohqugjDxeR1EA/
fL6apC+mvF2zvkrQVtYhC3v8FSbi36hDVx/+0P1TYqp9RMMxHcQHcryH4n2I2sdE2SifzmvdJMgL
zE2E7/FpEbK+0Ulti3m9Av+AzFGWJc7kSjQxR+aDkmG6K1nfbUB7A34SHRklpwesCfqehaWHWd5c
rFxrKetNGxRlbL87jfO4MAyvY6qUYR3PL8kE7jPaic/VnOlPdLi0Am49ERsXpPnIjRyisKFXzwFh
isWvo+8QXeAn/1/NOxkZ9nalrN1qa9hETSHuLhxzrxNWwCrXolWYLEmV27McKdmEC0lm7BIWI5W4
vx689PZ1kJj8QyjD5ldhkPbqAHvbFpZD/HHj6rDXOL7kljSqP/skGmajYnLr8um7GU+VeHJ7gITJ
rgOpJOkkNMkAJGE6QnRh95EyHPFlLRMxu6XhF7FntmK6rQX4eobErJENavpoVDYH7kq9tpGKwiN1
8QXzjYFjTJOhvOndpqOyPtAu1yzAVrfmjaPoQSVi2OCE9k5GW4/SbOvhW/2Ccw0JfC5fqasRBWCE
d4+jBTz4fHGBeYt8P/sxMi0BDaFHiVFXku/1QjmfNxNAjgLilV5rO7ASgNSuGo+JdahrMVXstGu0
vF38zPSeK2HF7lyfScOVkWwaamMl8wGhkh6+ToD3ROLBk26hX3e0gIDe0cpcu29cLlPocQmMQ5ny
Ter8anwnqfVjr0I+jMNUf6iV1hD+q9JuSn3hTupMlPwrtx8Z1i2lI0UTd4F5ph+9eRatVpYqGzoM
1I6gj46aFQvaplIp35bucONv4nYLt33iJs319+r9NHQIQSce7wFMhNmFCaHZr++0n14WfW1FZRjp
MCyVusl6KVRvhJnpZJihx02w3bftEm9MdJYDvldyJMmHZAZg3xbXCbGvYMRjOYlUZTY8hlD7rGdH
X0LMjpQCH+UEalxEY3yCsqUwhCYq9Jartk8rN0VhKtZ8JRLU1nK/0G6+Bpa9kLz4aii9V+i/F3Pt
piD47woumZfZzF4KpVGYZxV9GCAO5szKtOHithi6iMcTTdI7Y4y3xgweRaubdGvKePB1EX33qvlp
gI938QQ1diHFLrHtQZsPIaz5oecYrZsZJwsPdE0IwFq5q6ndKOInakKaU/ixda4BZGwze3AlI85D
ODNeK11nVVcabhIwyhJIH8bPP5qTr0AvKZ4WlKtzVlFniIoFyW96GKfsxhiu8AUTY0lBZXqqQNBb
gKgoUaIFvAYAyPl53G3e14gBnAe/3XxS8VLWrqd1GfbL7JKx/NuDvQ2vBemfL9HnvE9RUULertw5
78l5jJ7Lp8NTx95RubeeR+hMp9txrSAYTpLyWbDhGgN1UgiV1IYVlDhiS4fZbX2MWUWGLBL08+UV
LXe6CBsZcimX24QJl1JkOrbAVgaktHC74jFxucAxGZz2gbjkqkY68yDrA4b0wVif0QRLULPrCqHi
L8zO0L/vcKoYPs2LtunZ2nCX0XLMZLKzLwhzaTz2JbWHLeUBE+MvBt1cCqMyNI/Th1u1FV6B/syf
IGBdgt8O6l7k64eF/dCrut1Mvpq33uWguI8LSMZ1YzTKgavCvdy+2aJJgpwTAjcrqTOtI3vb4Mmg
a52Ppbihx9DH3aEAPklDnE3lFRyy7hrNPDEDrroTGTmR+rXErC/aTYIhGBRcFa9x3S5CBkn2exnQ
sWz+3Z70RYSj8KNDUHZRD6FIkVoO1LqDlwmxG/DStjhhDNP4pvyxChzoMiu/6u90ZjNiKJKrCvL9
MEOQyxWGiaSSLSHlpOxmOEjaQvMNnvtA6qyIILc/xOp7R1Adw8XsUXWcQv3uWC7Ly0cI9TXy0IEs
8jT2CDtCFtEd8t/0P0fP368Be9gk7l+UL+V4HZwsye/hizFU6crbyyj9UD5SjC3000VgMiVJDFD2
rr7D8f3HtpE53bPZsX0KauqgceZYi+cYuu25YctNBjFvbFAclJl5Jcocs7E54ibaGyZmJ9vOUBdm
M07uyPVWQh+69MDI/nJ8ywOYPyxCZSFs7+NKwJcMxRNUle34ixWrPSpfQ9QKltcECWOkpz+eyCyF
dalZ7KKDeqe1U7U2wpZxgSIgy/Vla61SG/+lWW34yDwyVgZCbE9xlVFta11DQ/gAzOAdAaVbNHqL
JTPioKYcPg+D4pISyQRY0I7C8Z2m/Yedh5bJYyXMP91nnrjly47jt1Xh5rJIqcjLxTsf2A0DFVa7
uF2Cup/6I667WMZTnB+biXX3d1JJumZNOkxaJvXKOXf8lmtzTZqJA5CX2iViYR68T/q88p0XZZxY
SZ1iXvIXi9lWnYpVn64saNIdV2U2658wM+1IHsHfl7uoY0HSOm7Gtost1dOg7HG3ggc2dH6uH10t
45/I3BF0w4SqB2hfHYrNa9yOd+Z3b94wUOWJoHPW69kucQV08dogD+d9i2F6YnvPQEtjwKpSuaKa
s3wpzwG+hW1olqsmb/g/KFnY+fZKViFi2o6MOW32K2RtmhyCFlGPdRP4xhhuZQhXAfzSS3kyXs9C
sSb4z8uK8bU5QLeOAPY7XnVDntTK4IEi+8En9stIwRb1YjssRbHub/814BlfLQAoQHajbcxCgHpN
jlKWptNmxkGv36evC+dCNHyaMzd28qKcke16tNMYSTtVOIbi6hMPYOtk8doWitJa8Letgd076CzJ
E6SFN+4WXKqAdvxqm77+ooTYU2M+XJv0XkWrGQnxvLAOhBHjwExH3GqkEPh8G9kMJxDWtyyeYgtJ
NVBoc8PbtZQRAHI5rmIZvpMEb3VGYlh0LWVXytFjoJLmibMABln/DOuUyHEw2PYUAMSCLKzY3DTH
ltP1ABcXXit9D8rINGX5z29WdVSv20RtWjC1BRrwQVgKC+A0SIjTfJ1XRkkfUIgBuy4o5mnkGVRz
D+yRcSZlIzYCu2sFN6i9d/83PZcAIbfJGfytRkTIzb3FEaeGXivRMhTIo2vRNOETpLe7BovkXob2
BZLNY3Eiup+LGIG0+Ze9eJdSfshyMRMtpV5sjMEFYF/Y/oWfR7gDxttHnH4gc0NSKWnt3p98gmgu
iaIpIYly4EnmQyCBI4Zf/2bfrCt2XFzpBm08PhLDB2fVUlpTH95USZ9XU+XdIw9zjYkzq21Xefqx
w99m7DRd06dkzYvOW0Sylk2SmzdlutEu8foOyEBo7WS6sTojhwqOk7QoSjPoknAt5PekPNtJ2mZy
o5HQFOVd4mizf/UxNtW8Rrhb6SkRBeQbvwNGhbBIdXhY1riSGBDFP46Ou7ITW9Y33X8Qmccvp+wR
DuTzdmaZ06ibRIxgqhKRKx27mL2bsfQiHsvOUPM/njCQrNiY/rvESSEn2UAMG0MybotsOXk1yT/s
WRT1VoqWORmBWMcauDNqZ6/9N1s3S3H0fkOZCEByK5CvMwYIkiuD0ijhfvjQkAqW0REeK24D6K8+
8vhfHXNodJ9+ROXj/nW5EY+tYOJPNccIkfN7p0qpKxKZJM4QSejSmPEWof9zdYnufhuezmdvbXIS
uWIUrdr5OBZebTijlIP44fQiyUvX1BFH2KtM024/LA7DFkBlOJT9w811UOv7WmS/fNvj8gFUdg7X
x1VUtNXE+0Xcw+YCAf6+kSU54CTd++u1284EWqpO0+ZHa2bRfL1wB1FvBCWfR//UhTqwnWA0bL4k
xx4qUhAuce3e+EHjgUIFQiDCW1lrrh10eONmcnOVBu4V5hPHXy4FjHESfXFGoYCN3HKISOBe41Xm
hRCkhyWjZqDDBAyrb2kCT8U71guszx1WBz/i2/ot4dfMQEshV5ypA+SfxBZoDfwgZ4YCDbEtiq0M
J5+qB9w4y4hrLnefroOTuLPBNdtXdC585xERBp9pyoS4SE34Hc00ZhUhsRgtAW15ImLEdYhFBELj
F6xQ1+fvuf+J0Ze+Uri56FLL2YJUUGynH5E+Ct4LWxG1a8kAk/HXnOXUQw+XqvcbZ5M2wu/al6k5
8vZdjsobEhb8ZDakEwfjXIepG0sO1Pjj+G8/Nd8nEY/zeCx3AX8jOV4jdV513ykmfwstlEgfLSG8
mYceuokZWYmGNpugScojGBilqbJULhl7/8igHPWCO0MZFnI8JgZ8RKb2R51qEc/0PQSBibDAp0hO
yYY5M6uEQKEkS1NTA0DrtC2FE+JUBXJS6ilFVC3VFbQSCX3DmYxkTSmmaZGqF9p79SqqOCHZVAK3
GcZrTd2jdlAwLyVsmn+VK08PlVn1INTA11HDDXgHijtqb/cUQvWaXg2YmNVq18iRvhdPX3bXQAlW
brUZqYbVGCVil5VXP2aSJ2s4fcRuCxX4aYltNujhWewpcNMwHKyyDR7qi5VDLBJujDX4bxWXWXR6
E4nMCPVPrq+U9XxGmVDSe1Ih4RH/lQdMR0xxGIFH0EwqDP3dr2lVrtRi4g/oQkEL5idY8n09Od/n
PrTmlVnz57vpBWjxOePW3mPl27UYsmCUEZ+k7juHkPMZsnv0fKouPXXJlgSXmVMhohn0Nfj2drI7
+70CAkwwOaxuebleYZ2GgQTCu1TQYLkuGJd0dczaxSEa5pWtjErqiE30EiOlbo/2oGPiEUlZjYhU
Ej2LFXD38ypm0v2uDBCFtTxGt3rBXqxZz/9mbMB8bVjS8dNvYnL5aQ6mBfbmP7yJD7z+jby49rM1
jXyu+pjXLjowVq/N/Czk+GA4w1pNVeKjUZxCDbNgHslMQQ9vvRQjv/hudSQP1Wd5ltb2a1U2EZz4
dxoc99TVR3Q7aKPFLiV9PPeTLYfwWWPf0pU4ErIGLGgMHbAHYVoEyIVJLPL/FwFLJzkjz6xJdlPt
a1n1xztGqnIadaex9WAZLDUQt1Thi6laB2W6bbPNC2CQHOq7D2XPQGEb0TeorYDLmFZYf/9zeLxN
RZowRMoH1l5dUFB2sx1roK0Q5Y2N5Yu0gEC1GvbjLZSHPGaNjj7GozE3GCSxhcCSwXsP0hbzg0q+
V45808FKUNk3nEaCXaYnOnBJKk2QVLGzZRNgH6ur+Y+emyPLq+l20TmVGZoEkU9kyuIrXU6F/o6I
8bNH9saGcM31Z1ukzWN2PDxBgbAflhNRpRBzOMF6tqpb/g7CTtXZKlk9dBl+Z7IQbSGe9LOvXfn9
6hCx3iXjkBzpXBKQ5TCcotU+stcrusov/9lwKTCc0VZLvABd7YsWI3vc/1/dYGQl89yVMiV1KieT
mzOLYMbeuZh9XT9wVANaVX9UqdO0AyFJSx72tyLqYJX133uIr5rmi6yEz3iaVIByb5BuV3gxyvZI
wM1Ka2lIFm2CsYwY1Pp1cV+a+htwcdXFh6nwEsV0ep0p5n4cJUN3OW6oPYBWlud5BkmgbSatv9Kr
pvNoO4w4UkMEJZzYiV8ulwqbzgazDxbNz5jccjM44aJDpIIhjBWr4rXHrJ6bLXwkOR6mqxa+VelU
GtdjwxaEpAsX1yacWYgLLV2kfLcFdaxS1MDVxO0IIt/3FJk6+QpipWyTh8/KqP5gibugrRF96pQt
2z0/tNQl6ad3w8z68cx84UZpXXYaf/1s/KOThNISW4Lwmomu4YOOIXpM3Y/DwTIcV1oJAjquQBZI
fl8wUSFGpsW7f+fWsOcOYg0cCVGHX8QE9xt/pxxYPE1ve+6X8wFfdsXJUVDwAHkZNIXPU+KXw9mz
bHSACqnklNuzAJkntDQ5x2FPkfAXPwq2g4Z6aqu3RAYEUHF5awm52/Kst0hr0QYwNg3fIWcgoy4g
/j129PTfH/OgrFZn0h6OGBYWi9Iu4XRR89FMhfurbSxILId4lUg4uAwnpmNIymbLGm/chfibj3MP
IIYSCLpk0wRVZO1vhWkAaimaxansovPWbhS+fQRIQzIlNKaCgQ6SA8mm2GxYSgO/ASb4x4/fxDKM
x/y1fr7ebBF8NzDpzmAHpQ+CnOpXAaKA5TiJoldk6RY+p7NzdrK6DImcnsOM8UT3s3vzLxIKeCl8
3CPo2j09ERNv9IZx7rQnZyB2mWK301WkB0J8eF4PXXpF10QBM+nfG54EbVudiXjvSISb+AcFKpuB
qf3hfMAb+bji0JKwhyLERP6JZSCNv42G2trxNeISPxdAz4OLCm6ww6FiMpDcxOgc6h07keToDfYD
QsZvlpKhy7W1jYiqYaUvdvr35AYE6vN4zyhTHliJmZnMNn43EqSqRgOm6aiYH1MW8led7w8bmeGf
u9It9G5rLY2btsfFCDja0ziwQtdPCbxgLi6fiXOdLOi2ysvmpevDEHMf1LHmjiSbjAwTRDH5X0O3
ECX18RprPntKNPdc97Phu7Zva2vFHmEKvuYur6ADET/lfjN7PONzzYdAVNYMyPkJW8PMeiAZc2q1
p6DHtQQXH8I3dYTs6LbST9x/Idqhw6zMaxO9Ky6iyxnzHIdUAXb/pYEeqjQbMCAId2JIFb33FPAG
wzgkdzR1fPjRONMdnL+xyPEljUk0qrXQK3jqEPmQvt803qdLzixYaj5neTnFXyM0hhDBBQHhYYx7
5WJ1DzsmtqzW0Nz83ph1mB4tlfbv+/JAUCk9MeiJ2pn2Mic/jwuDJO4+evvwLHTBMOTeTsCj+OLr
SH//1rH6ieVoL5G7hiICOJRjIuiHtgLT6DFJ8jGSWq1d8l6+cgFtA4AluxRRtcri/+8Zyb5PFgpf
/QJzheMlICz2tX22eMlV7AeWOUht5I881vjzjgkWDwgSmFDtsz3b0kmkDwMO4Ku+RslkliKEGvtl
VDsACfAKH5WtQ2Y7aiiZqx6kfTMIFUQGnBb14LOVMFCXN7KxPLhbLqlNCUglJJU6h2aBqFrp/AoJ
P6+hop3wOiSovSItA8z42q7G6L/dv7xSIIsUooxJbl2Snxcg9zcP8cLfHIHNCRr3SJZDIJprpYrC
kMrSfeNjCP+t/+kmJrCs80cpvCIgJIj+4GgZ818jf8PlXG+vczuuzserQq5yl7AXzM7dGuva5s/9
JL+Ia+Gl9tMEbECO4+JP8hSx6baNIhbN1nXozKOER0mrxIBVmjRIBI3BbQhr1xJyavKF+QntIxei
JXNpoYy8mL09LCwdIlrCFoj9Q2sFxEQHyzko5zEVxbEil2THAnpVarjvdbmQ2VYsybM1u1NUxNhG
RAOi6yqs3EAkzNeceH3n2s2DDHsXoDtts5qe9DzP/U/sUnivZBTj86I25Q1NWrXvR2nmXJT3c3SI
2ullJgkZ11WSWWH4pGuiZxcGvoJbE2/XgSgde+QKhoghqxcFg4vedxgREHtW2U2pfFzTDaSAz2GJ
NSEYzn64cA8NzXP80vYwShxCcFH/npcOd0bn02sAWp6HNEW+DeICGRc+DmQ3pNWc2yQubyF9HEOz
dI+8OmYraFg8ayWlmWAlU/GJaHxu6dSooOpG/wCMHfD1xOlNnXTTciyobXH128BLGYgRqHe9Fw6y
yisUb3TpZZg+6RycJWOtYu3r7U5PDKK+8q6o1vTLVnAZ6QyDN1VRRxEhVfwWktsWhMfqeBe+WGjv
ChZocX9k4ZxmWlb7LT1tzSYToEz9KeMXkhp/fcoTeRMWh8/wcl+/2kbqR37oG+JSwAJqXGmNzpbG
FINCaaCntArnkDWjP3dYi6+RIe7LBzSrRTajNtpMGZ1GefNU++dJ0Sw3f10U/Ov5qykx9/x6O4Fg
SgxWTAYkoSV/xDpeAkc9hpjwCssEbXC2+xEAvGyt2LresHRJ/42HuyAyUks94asD6Ax1gwQq8pag
9m+RZ+PAJ4tmeoGmz8rMcgp++7pC2FFtW4uL9+l6r1lKFIDhtqBMxaU6iOaiAOXpv6iavrw7laCC
QDYMRcfkXNhhvcxg3mbNM7DZMuvuKVoDVKat6YwSCjnyT6fCx/hNxL/z7sQ3iAFAkoHPKl3goWFv
ofdVezPrq3O4VuFAySXe4unqeqqz4S93t9w4nQeMIZtlSMZH1MIQAmXXucWYOhgKwViquay7sTBE
fu0Y7SjG5FR8u4nu2KP9UqZFEDH+6Zt20SPOFnxlEYWaAu3UiE9TylCU5s7vjNcAYrh43pwJyKn4
O3G/3jO4QfPc9gUSD0c4Cp7vT1P+lYFpDa0PjQqh8GFLljvQnGLPTLMf7Z1FUb8PArhn92pF+2p8
TYf0+QeIgqw1q5srbTRMpAmiWq92DJCni+GhySiRQAwVHMeX9GTbxMKkXGB0X6UrikISjqt2kCZY
HIkB3HVgMgk3deO3UjjwRM9I4j0Nl9+Qdp+WOoBKJoEn9z0HFxhm8MYNF+fTlElY3x/Tk55wzibU
1klmF9WJ1kBi55bTcjPx9tnd60cCqjsGY4P4ttO2rrRGTrTyPazXejqfvoJ75mMou2JrVZKpPQZd
KyuVg0ZdTL6Z/sbGXh5Z06SsCTWDUOBeuQ2/FBnmQ3T7Oq3GHrP4iuhgjJ/MTEfdWRxxHJOZNhnS
NKiATvKlv/Gb5OcAQVn7k37CkihTB4jNBULuqahrh5AGgk6KeAgQvShntPo+oxDuefZ/SPzVibXH
sj7UdJPQuqa+WB0Rbg8p7yxAk0y6JzmWOBXdouJGWNjv8AnsqAm1BpHy1FWOSNqgu4A9nc7pdmDx
gbAH5tzPbOuBStIS/rfc0sUrT8SBvUt4GGi5RJuqs9bDCpgZtQ+YRwl1TLIWFVKQS9YWcMq/l8LE
FyK/yMzsbgGgVg59NPbHc7QES/C9DZn4pfBVbwqyZti3Zqjb5MdSIg3NsW7eC+RWf1z1+hTiVflj
C9Vt9qmlHb/ZBzbypxJTfjY/y3QcDh0EyjzT3AWeK7qtmiIaPSjbhn267pKU6G+8VJddXr++ZXEb
/T3i6gZ9tFUkSCjpPmJ9GLaIFbsiA7nLuHim+FHlnvnz54VjWO5/P7fyqvT5evzLIzGTIwBayAOx
S0WVEPJOdHkaWVwvnY3fSNpYj2SZ6gmAhzTfVe9hSfHOSZbDwzyhF53bIAAz1UmnlaiuZHxBOn8A
STwZ2yEGnrOV/yaivLCqbhgHXEBlXvMXKNVtrh9zLQo6O0MqVU3ww7EfhJc16r1ezLDGluSyM8GZ
spObTW4CJMAe/plO2wVnryEIU4HleL72gbaGLJIg84ZFyEONsO0da7pVr5Puyd/X/1wRB/j/99w9
6ENp6yFw17H5SaX6kiiNt4Gms27fRkLe0beyPuDteZIMNJN53lX2k3ObLKyNh18yAxbIvzzRMKnG
8VYkZvva4dMAg5X23/+Mtfus65ubCNmCrHrrKgD3vOwyP+J4RQaS4VfdsAUeQ1fI/up9cdkALe5W
Rx1RodvpH4ZMs0Dz7fdVH/Vn0b3VYcbHuPnBF5ZMO7smKp5UkeCjO0ARMK97w5oHuDcZhkX008Vr
LajBZS/o0MEuvAprATHy1PAzVN9TdbspUBpPbQEtqaZwLeMERXyeo/rWhdLpQf9ByNY8RxLtdyPa
3jkc5iik3+1Ra/St6mlIKQWHXTy1Yosd8FgaOtMXG1PJgiuiiByueSuYH4vuYND3YtIeb5RsGygE
rVjtNfb7kXv+35zz3PEWj7/xszAgsOsFCK/bYwivI52SqZM4F1abNDlaWjja1P94VeHjHHImnpm+
Of/t6G4iVO1vjCnz+Fio+kmNCwMMsg06IAHRUS/G+40uIZZ14/4WVqCxW7FCrONZMBw799KWIvI4
dIoLq4c/PQ7x8eWIgsM34D6i8xt7SjBgt4eAHQfU0EyiYcSRL69EOCnmne+E7oUDi6AJXXRycAjY
VyoY919MdDv8QjTOwle2diairs4EuJRt5sXYVpcjPNw0tT7dw9QplPW9q3c6g6hTjGVeZWsau42C
lq3UzJfA5LCGqCRi0aBxsQO8BhZn2EUuUWvbkjWe3AZmUwFOoi3L4nziSI2niIvi+n+x/FTGZvpk
wlInSd4sS6CngdfxBrR9M/GIL4VK3JsnDgAkDY+UlMZmo3nbkag0dsepaUzP2CxtGRaUUC9ErADR
Gk4m69Hg0UBMtbBVaw64vjmh756lYTAyfJruOsHK1h5dGZZ1XZySVSYKvDpgrp49UWPkWpbtNM6H
OpezyI+FJ+QnDqd0wudgPxZB50VDgqVGno1w+JiR3bYCfN7l+Dbs1uqsN/WU0iTlQl/gTWWS6ZfM
XDdKvNpfcTUKNIatZI46t9yTNbSuE0ws/stSrxtmeNM6uPJevEKPpxGeQJFJ6kNIRyL/nXHMWDOn
PZZ+Qkm5YeQFcUet9nImb/AbLy4AZUgy3DUhN/juipu4u3EBHkK2tBRD9m2/J+dD6n5izDA2GA2w
Y4hQQTIqacZ2t+tiwVUef43VwvXtka5l5bjhq0iTl3DOaiqtu3MZHZoHsl8zKlXjfl2wn7v4Qmc3
wNL+xmsijG7+zdd7g1sf9pbfk+p7VpBN0AXt9pkvG+HA6Me3AhT6SDaasILn1MR4eaxRcvUZpWyo
HjiJ/Z2sNem3g5xV/oa/jvc0CD/ISLPO389NXL8fwNFHaJ15F83dwTcrLkU/9U2lkdDXpv2s+AoY
IedKDOjHiQ1+ybasmREfOKN+Rab0/f3STIyLJXfsWDWrhTaXcTBzAtzsUgZyOE66stGbhXOCzWV+
A/CJMJmB/p9OSIiC14/VUq6RnMK8jUxDClMcGcHmwJiixaCQBlQCslCeKsZs/uDWfPFzApKw4Bol
tu+xkTcnwDnnpiy03EKdk9kKbflOlQ1CBPMxHdjm1cn1SmfLdzAObmbDUXiYInBZXJuK3+hFy7aY
+VNdaAJmyCCFgb7tLX6fS/kY3yBfsZZIBFbRtU57O9QmicyAYFbI3EfKefpCMzs90y2CKblZ5SxJ
/odQyDxH18m0NP+FvFJslWETP5gsdYrr0pu+ff2K4uQg0w80PqTAZqSrSYLMbaaTKttKcA1HOCAa
SpAWSXRvkrgd7rTTz2EI715nkJllgM6xnMOdNPzIkgYZc3NVMTg+tox89I6JAim0ok/GTfRLyYXf
YOW3VBQE0n7hkEEmlMCGID6KQ2VJP5X9cYWyQ4iSCf1e6D8lRb6fUBRbKVkyCLIQJ/k9FZXRW3EO
LFtMsRp7lycE0vkS8zFTEPzFFp7HSNVFGJpY0WDpSB9+MMLdMGLgWoz7UwqUIEbOasC0xI1m4tol
ZvcWzB9mnuxqs9pc6NKb0fqk1tKjKUPzjah8TfZAMDS1oNNzmpf5v7iga7di1Z0UeZ4onj2EkTQj
w60BwqmPPQNHGu1TV3Qoqqg9jhpQPavgnlZbld66893IJyGSMQg4aa9msRslDNeXpqfdLbjV0jLp
AjXCWkxAiSG61RsRka69+4v7S2yTdk8K3YzftCEKAWdVk00MzLMQbxLBKQkGIV/+a9yPGpO0ioFR
kUyV9SdLkJFteXL0quxsJjBd0Y1g3ftl83937UoprZ3kEU4emn8rwDGD0ef/lUGQQ99f4yn6bMTM
BW0I6sMP/sGiJ77qB+p0w0isMr/3ifnrVdRrpJMiJ2fxJPdMRidQBSGja4jYf/M9Ko9LdUP8zHC0
rKoITRSOl4vt9Uv8N57r2lGQOBw172zUDApKn3ZQ7JGxQwsvpKFVZA9JRRNOU9U1ZG5E3OWoB5rJ
zZdjZ6kmUHv4L0NTap18Tu6eucGNe8DH2mvbgd8a16L3eh8Wm/Om6WsuH9M7qE9SnOSpMRGAxjJc
7n2vjwZLg0HNrkxnA6xvky4kX9MI928iJV3yG2jghX1h0MR9pOT+WoarbC8NyKczeKgeVN3TC9KN
ZArhCxefvu6zNNVEDJ9xvU+rwv6uBBbffYV9Isk/RV4Si2bexbFmp9VjULiniR5Q+7avVUN6+uNf
tfnjX6HVYEbvBgA0LjsstVYDg9N8F++VctFs+xAN6fAXA2+q/1kVpC2DzG76aBvqFG+UYmyDbzl6
Enfoxnw/g6hq99gexfq+URCI5aWg1CkQKnWS196KgjyvS0nXGEgWLow8QuuZZlkbNxmw5myEAGpj
PzUVdjnHgZUnBrp2oyE+FJD/qvu0EvBgbRvR5nFGlNGYqGC11VD3lh6UaVpkj3hk5MuvjMUHnjTV
mPKDFXXlggh3GLi0ZT6af/Tx9aeV/7RNjFeVhitH8RcATvxpZ08C+7Cx5uxj+qcZHk7nkQVVQHfB
XxVDPnY1J7pocDGNKfHA4yJajUmy8IdThz2nq4iVTqYh4V2azddPgqk5nbrwb+JlvUOD2S5zEkZz
QDTlbc0Ffd1DFG9ygfucGlN0MuKz7vpTKgSEQidVVujtZmMCz5kgl86Tj+Q/gpYA9dSORTGSuucU
mrUTlGU9vNf3NbiAdjO7da6X+deBschqc7DBRp925rUAKeftCwS3JKs+7qK/05srWvtZ9nNNiwni
X80ZCWIid9TvWV9Se2l/fbgUtX8GO6XQZjXam8IfODHKnyNNTPVZEFzLNPo7WbUi3ga/PO0o58pJ
7bbyXiLgXVak5yQCJHrtw5ZO4d/5PqDNxAaXh/s1BCBAKjQxnRBeAEzJn8KswdVhI7W0L8xNvVyB
vTzlsLuWfQIBum01L02LcJWqT/hyC3ZiaX5VbVsQkfurYLsOoPCnSCVZ0xt+6Xq9J/q+cc1Sxloa
kMyXomkhzQIYRIRaAFgS2pBeSk1YtA7cmacto7oQDeXLPZLGLhxQe7Fnvery/mkxsKuLNC77Sh9k
DcZ7rulgftU0T+vWtHmgbblHU0efwVICR7ao0pnz3BjZxfZWP+3+3QyzshmklRo8xU0lY8K7NPLo
QhoZ50AXj1Syj3A8sCqHuYRNG671qb2lCZj2beMRBC9pLaV/2gaxDzn/o9Guj6jUcJqrtGBrK8CS
VboFvUlUeNKOFH9AqrkfKL7xP3gb5LkTozby4mX/1lT5VpGnErZmwWipUGc+IEEPQYYVXfp/1l+N
j7Nfw3s7c5b0r71RyGAtfZySwfe7ADI7SpFWy7lcauaZijdSILThECzBl+ImiGw+jDYebuYIZYEl
pORHKVvywxvIaSIsble+5T/u7DeZhLvwI5l2vEYBV/rrwFMCoE7BEyRgrUQUzDtiMAQ4ub7ZLGrt
AbtQ5NTJjCNKPUXvKjVT2UM3LSLIsfY3Dkh9DWRGcaHi0g9hrI/Tw/emKosa32tpABZSFF8VfzL9
35PGwDPreP68EKHDyAbC2Sp/cHgoB9ZpEpgBi6q2v4n4H3xVJWvT2pwDyj8skCK1tcffF2cunmMi
MG3DM23m9r9GnMzWjTlA3aqn4+/jpuq4SlOKcmXtKxtQSXOOsrVEcNC6eIzauKLD8eLpdalqM2Kf
CmERFF8CB5IMlG3CTsh2Pp9oY41RxDM4Lzqs0Ma8yzJuqLRygiDLdg8OcKXscuInWpsVBUK25FHb
rCgaxYpinorL2+pHsJKNkXUlnZtgMlGI55uMVDZJ/tgVz5hvwlglg/AAJf9IKNnrrMCiOfYnug7m
zcyPsfi2xrWOQSYJmffThrOlck3NQhkuiYfiFjHYkVnsZrarG9ggZFm3/pCXwhDS4zFxPubsNlvM
TrOqHnfwF5IchSjmrV3NymiBVOH/IiC+qCykQiXHpSqYB9Y7jiJYiMILUnWPy4XBMNGpKa5dDVm/
+qUo9vVBMBOQyUQ5GFkw6JNs6pSGQlsc/+o8LVr0biYzBZsXQT9BL+fSLi2lFGSWNQglR0gN6a9S
nBsFNgIf6ndenfKnc6RuTVF2oWzhQE/ZMuf6JhHLCLJr/sWXkYEFudCP7rH61KeYAES2Wt4uaENh
re8yJwImSsY0D5EXDfcAjQaH0oSO+oEi3HsAlEUqN8/N7TTQotN9+pVhtmNfa1G+VqyRmEE+NnbU
O+IV3l+pXDx+4J8OodJgd7/LphNvBYsMPaJM4Ew3AlYosQCCcNZifWBKfOrcmh3plWF1AhjholyO
Z+0SaOvh6iGa3wZ5p0tihEhGLSZeevJNgPhPDe5fy3hfbQ4IfE1ubV08aEoKfDzMZTgmC78ls35M
fjUhzjDV+/Up3kPNFt2JVaZAXT0A/En2S9Zn3UjoO7XB5iDM31Soli/Twkbl63p39A1/gBAL0s2P
oTEz+nSR/y9KYuiifePniNjjXDGrRDSUH3XBsNEHGAvmxRgROsvQvsiKT1Rj8QG77/n7LZCBt/fj
t3cXVyElNMUKT0auebyKnQQi2/xDqIcaB+kwPmA6eR80TzjsxSas/SN2c+KGfDhlCWumPXgNQrSp
BTCweZP7aX80z0O4LJGRxkEdPX4Y9zv7G+WOntDvJ8i4pmZafcPARsvV74ZTaP9DiTJ702ubdv+q
z72T1ZUysbb8DtcVE8xTw1uRO4z6b6FDNWex1bFnyv07btqlQ9K97ZradrQn4suK8Hy6hWdWoyZn
Sm9mIZT2V4d4W8khXcNWp2YrpXBg2yOgW/eUzR3bFQorilsZb14x7ab0ZPVs3kePfEOXmqSF4H6M
QalPKu/hHZ/N5bxPzxD5+IPLCFsBl2rsiXtVBWvhChdm3UA9jfAxtBo7eaxocV6FjrNMOI2B5xis
LuHhBCI4omFBuArovFtWgc1pZyFfvFtqq6UcLMHU9GVkve2GZ/uTZoS5ytMaUm2DFUlqoFUR77mU
HuS3pzy5uCkzq4uNf1Kap7Ot6D6QZHmn2vOKdnMeiAleh3rNXb1GVO5NRnJ/Kb20GHARGkpQjXfR
lc6kJ/CTn2OgHUqCZHutMkhunZWw0VLJviaVJdE79D2zgY1l4c2mYzRPv4ixtqNeNnC8scuO+Jcq
CVMh6Utq+kBaLUwHGSdmTxpkV6DD4U3ZbHpDNqH1FicfzlJcLSHo2+to/8Etqvx/meeCsOIS2Z6w
FH9JhACr2sUhlxB47wcsvwubN4wLNvO2xO7vANoIDMEyV+BB3IBRil/pDlHNWmAndA26jcYv/nyp
Ht9I/lH8B8/MFc+Fq9xmO3ZEg7/oPR1nmz8HEZXYmG9rYg40oEtO8zEO2gsg9nJnLZAOdKgatniI
A2IPvUFldPiUzU5bUHaFzcRR8x/nCZoDa8oSLmvftmieSkBu3sZD+8e10nu10AAW4CKDOXWvce/c
532/hvDNQN7Y7JMl+g5c8/GgcETV9GmjnheYxM/+E+mSHAGN4TUmio6RpZ9R/7fsey2aoInjgnow
u0XzFXBxp5tYTwFBiyjqFNXfYPbCDrFPSqP4w8I46rZEnAG5jl0MgNd9HucoAtCczSxD9XM5Xpc4
Kw2he9gj34nkqoyXFmvuoaDIbOyHeryfdIHFQE5Plw1VGjXWDqWGXeYU8a1mNLqhDNNqCZVFL1an
uUnhRBQ54rx9RpvUdcW/fV+0Rwj4ecdVQOBEh0QjPP+q5Uj+D69w2iWr2qez9vKCkjQd5jleJNu1
PXZoIzjhmTVz86uQ36y8z1tW8b0N8rfKJOKA4mUmFVUDlquarVzWnRts4H9PwnwJbR1yYWGopea7
jJaocRV9+Hama2r/bjLgjrtrmvxfCArwCtbP96BNYg6BFl0qdxUYMyrzH16DiAYDXwibJ9VvmVMe
rpu7CHR1SoV7h62AabDqb+onhh/pZbRdNgMaNUJeD0sPryPxeN0GNYizf5Aa+0PC37c+OrP4jEwz
Wd2kPca4YuD5AOIsv9cDRKhMpE1GiEwTViYzA2WBlUV8CK80sWehH1wtu2UM8PXwfgVBXVuo7fa6
T9wZm283aRXf6nhoZZy3QMlzwwdjVKOPH4huAO2h0O73g5bqAw4VpamlvkeKkI1Uz2DxtZvxZL21
GXMVzwJhvefhWmcEs/sQSL3AeP//xs5vheD6d5dy9o6QxCnaHauRygYMSUTDpOo17CdTxgSZfETF
6ftXOgbpbzC8kL7flhqu0cTW7yE7Zqj+yIq7w74sj5Y3OCbYZPn46XGTlYYZHU/DDF6I4AFr+n+T
ds5LpYwcqTbidAOxxjaUQEhsOVnMUVlAIdOq7LYxKkXxNt+7Z+r01JxrSsnYPbfQcpMAHVxPy8KL
Sg8v2N0W66E5WTlRS7hS3qn8UwyTw0xD53yUUCu9SMYtVZAX5Rgw3xsKhXJvP6bonteCnAfKqMPz
X7gcIgKiWclDTjZe8Sb44wzbKtas0GgmlxPflJPltLqGBJKlLY+C88HKZsF/tqFcFJbguklLYT23
wDk3nSVNvuvtFIPrFtarM/LJK8baPUJhNnI077cn0YURke+ABCVmdBFzNCPTwKa0KMIKROWxVxqL
ipVRNagSr2DYocKGdUdpQ83dH0pNcZOnbknQqy792wALr7epBt4jalJ9PWBWv1vb3D07eYqcwpjz
/A5OKx0MlmTCHMP+1V1l5aipYShXvtsk08RLPh/VvJ+yXu5hdYNGVZz2lYmj33LuFO0TtCIMpSQ6
kGoslpnX/HVZsqLeFb4C1re/VYYpnnYZH/VeElPVz0+MEVezpLkzdq7ltWkvT36LpncWdvJuxxd3
6xSYzbTrgDTXYLOqoqjXV/KPY9nIqnf9zuMKFOx9XT39r6VhdO8/umhhHlslFmjjdwacO7AVk9EQ
9GVvu6HfevQoNPW8ALpnoC0tAPq3XMbnByfqzXcxI0VSGnOsWQoW+PWaVY6TN7G9MkRsGSDMfegk
e18byj5L1e3ITTLEgAJtidXrEAhmMuqIhjkZcGicXOy7KWZDEfuKEuec4jVfFPQJjFAPhofE/y/Y
f18hpjeLQmHZSzeWBdzymNZquFnDn6ut6tp6P+gV5hqmJpFJPgG2hC4MnDZwwXQ35xAsjLLYJjG3
ACsrQS2SMa6IdTRWqAA4GqL6+opsXykqDqn+BkAFyk5CLxId2Qa1RU+uxFJjxuI9Fmm9u8WJXFC9
I0xweye2sCanBjYkOiO8kTy9P2T3RPAPn2ncehxPj8n2FcEgTQInIXrqqoNBpqrYRrmH+xBR99UM
gTjaw2tiWemiwKSqgr77L5158I8IZaSP+hKilmcRwIlS6JUCZUfKoMFpFybVDJHrkwigVxwAxKrH
FvmRJjOz1ENDYkgVOdTwhqPnCBkxLw/zUDtqjy/Et9hzaZgPWVd1qOPEMqLVGbYt2MudTKfa8xj8
Ha6dLrTfqaWW002IBstd7z8YhoI7AwaXO83ryNY9mxfcZpk6NpRad2zsSxFsv0uJgfrsP4JzjlRp
PI1pIrNuWdbzHyKVLr0AMtfwqzEIT0kaYi+PoNvTXk2pnrMYp5FVsowZsIEAV+EgXvTZuOKBVpi3
NfGYRihc/NY5UBzK0YH+EYW01zLxh0C51Kl4Vi1k817c6+fWvoTJk03gIt/rJtBfa+Snw3BLBfUF
LRl0OMy8vzQuQg+9SoLaL823a7o8Xvou1LftGhEssvmMcSrqb27y9wklmZrHXS/BOSjc3MIU+p+f
nCnz2aqRjvzX30xd/qwpYxAbuId8z/JIZcV0J3Mx0T61h9ZrDv0Go1mLGpmyVM4ekrlFBt4SCJCM
SSbxH3u7H6wEgzot8dRmtcXscXKIIvxBMKPz2egZsw7z/iSPmpiFKaUA7a2oRyCmoqjUBlO9eCxT
YagUQWpvZaq57ipsFdlMbE+P4s8ah8hWQqF2+s/6oKJMCf6gC6lVYdd7a2NBngACP/czooqUXtT5
VxBE0bMYNwjh6wibQbTqaY6xmsJSFyLtnOGonH3K/op+oFZL7rzrYh6DPechCU9+aRj1FRN68Onh
yhpQBXu6xqPoA7v30u62eixmq87jOJqVOVBMpuTH8j8qHVaNiUjBaHhiCSlx2aoB4GwtP7DH6RfO
tP8izwUckVn6+fQfGtbUmpJzETYdYNmAvkRozj/QUV6P2TdVYt4zH1cSHRRx4djjh/YTz2VfvyVe
Q8WqsWd4uuFhshpRKoCTYANDc180KCn+YyoLxy0WGZp4CUhhyIUVGn7KOiyBKjgQDRcpEnez0/uX
dZPJ7ERqpz+SZOCp6FFz7Xo/0gAZ4L4ZqnmxhOWl7sHd7N3aRazI93uqAnrVquqJzsUpm0TOdhzj
kBH5MYC8rKcjlQdLQEwWAJiaMjR3r87lvYMBi1J3urKNIM/bjrWZ6sKk/FfvvazixYwGZRGTEZQh
kDrcMH9kX4Q22rV1hstnROraL2FxQJnfywp9pxnkfcB7RnO3MpYVJ5hlIHvQE9dxy76fwz2isYnW
yRYgZdsqVNRkurwqesIKMeSs4t3OJ2wONMvib6dtmt0jRxdpp/8siptkAgOP38b3XkXQHqBfTURN
sBpRFx3lE6DuUIEapV6nYKwriItAbZ77XhenhPRcJHnJdpe80vjQzrMf75tTuMpRKzNuv/lU8xp7
d1KTWy+IyDpSviz61KRWwGUYeg0r/VZVXdIWxO17NFgSys0gaQH09+i3FUkCs0CwNp+WXiMyo6aI
A00P8xQBUCIrjsJWiy1421ZsAsctzFhWopvdAH8GNOAdsHX0OsfSmq/AXNreCFmT8HQLx87btrRH
4si5eZWyGxOsUn1+qp5HGvTnuHBbDWljRbkW7CkYOzHhR8NZ03Turj3wN/ffL6+RYZ7oa7Mj+u2y
BT89jHfuptOge4lppgEW/DVgJm1iHB0y+CpbJHmb6HJiCMUj39gmIWdh8D6ye0pFinh+VDxBjTtx
4x9Vr8FidRXN0BdGZ1mvnvDaS+pSZWaG3P32EwccBZMmzcV9ZzkXmtdWVK2HN44o15KuzNSWrkka
6irOkKZ1+gbIHEkfbgJ4DszuRbP8eTB6H2mDUw69X9XJTOsg0zhNO00EZAbfNr0cw6dQelGm77u5
C9VUonH3kfZBagWpJyTUkBxdscSYc0xE3aeYWxLOwfEPTW30qXfBYWPY5kPfZVVbkQMyiEgPsk/F
HjVlDRAOt4Cj2PlP8sItqS5nbW521picw4sQ5T1uEnlwqaY3eSbEwMDKToIWu4I7G8OPj3L1vDK9
+PgnDrGWdwG0WuBeKwREfKr4SV4jjjbkXFyS9m2Qa0GNA7eWHyRUwL9pWLXo5aFiqVKmQECSoaRj
8yrecxV1SkspJgvCXA21dn9peI4NlsrgsNPpX1hF0gd14qdGl/kUfYa20GP2hKJSScAdSGs9jZ7a
8M2ATFgFJXikk8IjW0dfLIMm5njAmyj19XbSTom0c0g7VRTw+DoDWAtkFCY4zGybyfIuhgbIoInY
VtjEBUvoKiSX/aU0n1S3kbs6RhprJ3K+Owwov7lafVAix9SUfieJ+RFO9O8Fv0TG1vFgTRQOxkxb
FpbLME44udZiHThOSc3IWkc7/iEkCSu19hz0w27/mObC5yapjrJLlVPJzeTuXk6pF+GS8zLhdHml
r39fQp0QPLz4xJE0hyR2DvqhnP3htoybaOipQFYWUfWLrTX/C0WnK7zCDs9dnEZh4n9GckkrURJl
CuqoZbnyBsNZIwdIKqXYuRrv6iFOAOEGkgMagkz+7p0Ic2DW1bbBpqzlKBEKdXylqR0K0WyGIkOz
HSxgIi1y4zdJWFIBNDpXCwyG0FhyMHTAHT46Eb/Ary9AedSrN5bUTOJRY7wlm84EZqqDpICWbwtg
xwaf05tM/7vP1bXZfApUSqE8dvY8KkE1FNHISbkeSNCkUVClRA5ClSgA1smfcoU90sEofYqwp0t0
y3cponEk/BKd8qXxoAjToVBPMsQ8QWD0bXEEKdiZOMRKwW7jDtW+Fy6KlKF5bjo7O7/MaZmL8wyr
xNWyD5PHVX5tg6xFVJ7k1TBN2AFqhbwtc6g25Bebd3OMLhX/7L2RNcWJol+OM88+mfehZvGdfaD3
LUTjrP5GUs7q2VkQ7YhamKJcrSIPMfvdBaD56BYouuJSooPXo0KyCMRSvZkiYxndnRlUxBQXQwau
irpGR81qo7jTJeIA9jcYJkQ+ZOdb/deLEMQuY9ABZWhMCatF7VcVVG3wgJfy31cXiz5oaWaK1iHs
+OZT+tZSzgeDd5n1j/AwdZutcowL830oFt1F2PfwUvCfGLZuhUWV+P5fnATfn2yMb6wEwdWA/X4v
gZ6VhY9sMsH8c6rJ6pwaF1ZeKSDAMc5rFDNnDGkKXLZ52HiS+hN5D+HYezWEUk0tAuGyPTMsnEob
FOQY79lX3KSDA6E8gvnhD5QO2fRLO9Hau3tImutuWNRsZtmHBEPN+128g4s12R8Cx98Rz0OX9ZQW
lvrW3k/9xVfyXPWRkRZOlbxR4+8xs5dwoI4SLElDG7z9a87TP++aSYkGR5ZNTmwmwLXWVbga/acp
Ua75a8s43naTEE5nHXxbso6wRPYtMcrqXg1uyGtXAdDKABZSUlqS7FOZkZo4Hqkiwod1kGRWKDGo
5KzvpwPXHDmmsDFGXRAKFJMCj9RerBo8ZGwC0d8P3JNZs0EJVuCwoRjC8ZDfzZAteI031/3EvRgj
y9AQhtUH275YYllVf8j/dTHeMI3TOt0RPtL8lCocYsgCj+egNF4+g3wQDdyymmgNbeXVwwjbYxqP
cVBH0XHM5g6aDN8Xdm50rdgaFGTnG7Ya2NZICBRC0paL15MxvnOYY1Asdmd9jmfN5rOeBEk02hy5
CX/HiBE0IxPL3KUALztZEJ8Cm7eE3XISI6YznLHQDaQUXSNHxxQSW/Uor1z9ptHkC+HtsrheYDwa
lAmOfhR7PdQSEYJYLTQ6hcwW1U0vM/jgrfzvnt6PMZYIOnlK+DCjjxQONRinWRz6u6O1eToXTsFE
0nyzfHdKq0maqXSTbmDJ5qu+VeP0n3tpbaGHVrVpcKYAuf4hA8+GHW5RMcsbs936psXNGE7gshuh
sVGwn4NKTEhhwm5KJnTh1XG4HDd482141I2F5aDnqUS//9OXqyCQvPemV00UDyylBSDRa5s8feIi
cHpETGl+7HsMN0aJRj0keUfLQM8pUckDmxAoZAPejcryjplOFwJyPVW8YZuXpiLXeY8PqS/TVGk7
d+e6M1NyrKJVAcAlD4cJmr+eNoZu11QPClMQ4Ti1NxyFqnOZ9QI8k0FKNzYilqM0yEHatx//JeCD
y48IU6OakXpRDsTh5RTAhBHrUIs9bu6fTPSYWwST+/HKlnE2Nh0rJSNQmaSWSXdBZQCGszMxk16b
6thDjOKIIQyfGppr7p83vav8nFjZ+ujz3LvyQKB8w5Gr38gC4U52PNEzb6xQLm9VOPgrOMgskU83
XUlx+c09lzr11n/EXC01OBxenvOwizEM001vRqjsDVlU8FGSbOjQ0gx0+MMzjwVB6cjK+VpieBRL
56d49U4Kh8m7EyQR3lqtAp/F1VvlFbVDQuy4rsWoDBZjVrv3nnT/iao+Up6nP6Vwy95HzQbuAMHS
yDupHsBqtsEnKvtGxFKaFndwDH81R28jn7JG9uw78+NvClBLou+UyDETlwHzcqqdP4G3/V47NzBG
WISQ8RwY2qtKJ9P4vQNI++X/BKu6JRE2Nm9LLGt55IYZBCKCA2NjRm1DCHQ0lgZH9tpov6LMRRpn
CUHHP+tqZ0f2vKC8gq04cGVOonkAXW4lSm6lxSo9IqMsB2A5Af79+OfIjBNfX1pHG9pSEcyF5svh
mKD4yIJ6aOY+eUy+HgYGhuIQS9qecxJoXdCBZx5mi2XYEaE52N7j0tBn5QGWPDtae7AADpT4Fq5Q
71P2jBx9ultnYng/L4OdngX1Kj7DoheHcMRytswrqhq/IOhOz9S3dkQF7EtqNTUyI2isKxXBVZJ8
CgtFUMP8uvFReaRiEvUIXsXS+NeVwLP+qPCDlvTTc+Ww+1Sv22drFtdaRRD4RbxYkkEXkHzFis7T
uPVeXeZvv6WWCEJghHaU+ijdfM/U5l0cy+42IbXJg00tnnMwwo6YMp6KZexFx/hZBMS6osF3jA31
TZErh7tH6khGZ+2n8A6aZsNHw5d/5EZBTUsGa7Ln25TbSNTkdDov/QiXB0jS1B5RimOsSaPpvIPq
3tCnhDheMFlAHLPsNWEH/fIsT+iDvoTenL7en4P9Lp2U5mZ2B/DmzkeUGTWmDzl1Mi2R3t8asGB8
uwcoznDIR/cxx1/sP79xihdVEJ3FuK3LV1Wpxbt2iR1DaYKa9l/097dtDsOQf+Q1LYn4gbq85PJm
sCbKcd2V1VAN4JTRlEWv1EN4v59jDnWXgIG3f0Ch3UblzHdb+7rqCTrfkNdZ4pipD6sFidjjBse6
j+qz4dvkXRp3oVTkremGTuETH20DVgFYdB9JL7FcZwf+tlFH677O76GZ85dgcCwnLjzSgPcXlncm
HvMBaD6Y00h3B8HEIG7zzIrpdDA2E9sxtqsEXQ5SWPL68YsRndzESFNbdryxm+cE+q0QPCOsFCuy
QgnB1iDG9pASlkZtuLcxZac6CCX33RnFbXPYgWN/AcJS0b7SsPq87pBZaK+2aGv5cVALNc9WurXJ
iHN8st9mHjFNQm7D+TYOYmu1WmmlCXDUoGpqWiXiCxJVuzpojOwN01lVxcNxQRV6dfFhuaCyx6zl
DRcIsuN2pFKRcNB07sAHvE6TyrmHkDHO64/iDdxDn5/uOwgSnHmRv0NQlqRtM8pmC4EFZGggclR0
+IabS+vFOxxDKVBTTAEYgK1YLalvZsnTxqMDjFgbqa2WPaGvrdSQjnBdd5zjLsxP85jsOntwPhHM
3qdX6XYiJqLof5jv27HAjjljWOPEWec5PRDOKgLAx30RibPBeWP2G309IQWp3WNEQXj9vfgenNhU
eX/nRf/se8beYdSgMZvulUwcweoQpfbKOtbE50utmGO1Q8PRSh7rGhurasUV06ok9O+9yxMaSMdP
8kPVvPZt1BzdbhuRIgT86X8OsoWM86ImecW2b/Y9OwfisBibTE6SJdDHe+ruW3yqljZ6dVYJl618
HJwbM7D1dQJqx4yJCtQMkSOlUyQWGQcyrEsDfCfVDH5sckTnbIreBiQ48sSiDnuiZZSkf/V3euDn
AaTuA7ToQYFaRU+P69c2GBfyJ3bUbl/7XQqFjwaMhsDYHfVG7dwogO4WrIhy2wj3i91Cm107JyJ7
rtUDxRfR+9gg63lZcIAYeJ0KGTgcLd5PiDHimssuZHBU7p+7mMSV9UQwxMuGgozLxClH58ojLmHZ
z8YEwiUx22ur5hOFQJX/cfEbim1Ru/bIPyxgYPFKmSiIZpnBgKnWhhpXNJUymCbVg9Cq5aVWgsDN
F9g2UeSrU1+m4LudQl4Ooyd/ypTwzql9ZzpEyIOYqT58iqq1Ebs08EXBIuZr2QXySfrAMLq2kxUU
UX4LJWG+XhtO6JDHG2u90eG93T9WYdB6Um0r2cDgMmBtZV1L5nCmhZ1sx6i53CQFtUYHUaPvghtg
vUXCPtQvRLeu0My+pa7EksIafoHWK74WegyAgXPXIy7FaP4eOFJF1d84OnsvIBIdsTL+7H4YbnDa
qjCv6cuqPuVbtGYwOI0ziwz0+e8YFoVxwYdM4XWsyecB06t48Qi/ejocpjNMTSd9p/dihVbFTb/m
BQDj8tVnwvabHakr9xscK+a2s1UCmsERNLWhxASDetJf5vimXsvln3Dier0S2rUVG+YBB82BUWH/
h6GOpv9WgHykzzfN40hG9CoK76gIL2zhs3/7Gf6Sxw1qOnR5xc8uvR2NaAZ0M6Op5al0JwqC4j34
r0ZSp0otlatjQ0P5wRkneUSjGC5oaN/geE7h2uk7qHAUZarRnI5xPb8ZLvNRa9lLExtB+Y9mpZm8
oY71u9g/sPfy5oQDTpBcdwnTBrb0EducZBcApmELd/U2+8gFoI6G1W3es7L6Qbgbee/zXN7TrL5a
zgZ5teQN3+TzfCnDphkrUmd4bRcEaUbCu95+/wBL0Jf3uCKh+g3T0f60R63tJ4K+pv1ccAR9jtOU
M/LEhhJgeq2X71Vlk3/ytQ5ezRXBrdPyjI1OPaRozrCMnCmK39osL0UH453PE59eXAzOD6yTqJC3
vbqE5MeGsS1QFh3RtTZPYAEW7BSPUm9k/mt6u+5iF+zyCQprUnbDM6reH9q7riXF1atY2Xq4awKb
OXY27JGC0jGavUtZC2lZ6YJTTIwdCWiMz44SjivCBVixVkjogNvnFNsFGeaQp7m5fjBrBoPehVB9
LSjASv5Qd8jVEFtuNmBXMC88IouREj77QCDI5JXx7fe4Ba1PJqlLBiNMvPyWrVj7AWn9ov5S8m4q
EQ/N2Sp/hKqRnoXhW457651MrvKhsrhEYg1+eVu4Ye/M7Qurz7GyBmStM4jgYHyeH4ewi0RpQFet
2M7pOX6wKn3CJc7BTo32Y/mJ3mdgjF8BHkeUMB0DRZt/tqNd82oc/IbPP+zRDDQxzDpqAXaQHqxO
ok9J9M/xoWuLKS5Mo+FVcD8iSU2bgtNcSEGJF9f6O5IQC0WfzvUMaG1AuAHabzqyQK2uikubB3uc
h6AGTeWV3AE3tAAYgdDYegq8ZOyc3QW/94Xv2l3jBDj/h+MfMuCdz5BK5AC5ZgxLZ/k0H23hhBxL
dQ+Agb0RBwGaLm25NP6A+2qMlZCC2IImDJMU7b/CqvBZHUlrQmI//G+pqLSF7hIUQmIbz180kRwE
NrqUjA7LdVd61+fMjP+Ad/Wv1oQQopC2z716tBGXqIPsrrLPu74XYIEmnr2J/tSOMQ3NZD/jcZL8
qlT0rpUv+EzFZZhS/X/NvvdcoQh5ZdPgomoS7Qv70IgUuztY0aPyMrTDWl9e0tfcqTop+0vf0KEB
KnBwKuLxBo3iSa1fJjHaRfJZtTFnKtCAtWpEE0JCuXvEt+3OdDc3CjtcgqzpAb6GivBE0Q7Hm3Ud
TDQ+RkAvyBi8U0dwyJAUIa4sf/JiGYf40tzzpBj+JNaZGTn/9VHy2nAm9nsVgUmwJnZgpQ8fPr2t
O+19/5AyGerGwE5yLKrkFS0d+EHLo55AEtW+AgrTpjP2cnbi/mr98difqKn7+2ujfSmt7bBhEY/B
TeWuR8SQdsmwuqUoAV2T2/bNmily9wP7BdIA/rFiCV87w9g1ATLIzHm2RrF40VoaYTTn/GHTcEoE
HtDlKeViryrZwOMF0vWfGhwePmX/PSORJgF7IsRzHg0cJWr69BRFe0+KqSgdX0s/aqeLqtZuNQXy
46llyvuS5gwWfS3yijTunpprkhH0DzIMWXGDI7/IirHjYJe3ZeTLaXiQVu0LspW7hpdDmFIgUR4o
OFg8hIxa67ee3ar2v3wA/OgmdkgooD6oNkLlGDezmrJyVg6Ge/h77duVjc/tG1DIjGsclydXn9zW
eEf3xjtG/dEJ7Zpv7ystFP1iaGI5uiEd/4Yvc/FeMkjdair9fUHntn/99hhUWSeeTuQQeGOgRTYx
l0rLbYcIiQT+NxJvoafWMaoPGgd0f0bmWEjIVcv8FwHPKdvaYWGoZM8MtFXUOcYpgO+3/JBVhaf0
eMN4gQXIgmGT1aRUqJGxA0QbkDwhaEfXQQiMQysUbXdxy5PHeD91ywYZNVAfQm6r1SvBgjyg3KDq
Jm9WjFWO4Sq4r31o4WFqUUcH3/gc03EnZJ/xLZXTf349UkwN26P44gayHs/Ybn5gPK5MMYCZHEAq
kJi5iBi8yPEyzW7RISSZ4tt741kggOa+/+eLWMCxv1wZnej4rOMhjZXgFjz1Qe2RS6OWYZ8iqWvq
bMvv4orwB5MdxBAJZcPfvMs9IQU5nDZXFSj51wFlbmLAGYVNTG9r+Qrl9adTgguesKDCRHrWjJxD
4vUvA89F23jnCGHurmSU9dc8uxBRwrRS+tPWD3Ks6rjIZLIBOztl+6PBFZuxg4QxDpDrPBd1FRqu
riIFiRUXLyzdgd7SHnGozI3B59WPRx8yElZ+DRYMqt7n9enqNl7y/1pnLs3eGfLfhH56BOvbokUG
QIASTS8XCnSYY1leEfw06nVQNwtcaJBIDgP4i4s6Uba3ygJwFOlmAJ2svu5FdEmpR7b91u7XK+2w
DvEQ4Igb6REwA4SSTfHk8zEFkBzXH1+JYQ9wd9FRVHEo7VH5HePbiN2xVjWtkzLGRwl3nOftyCHc
tnpvz9SVejsYdNiVosNhZqdp15hSA9dZ4Vo23dT2ZTusZELEFgwmdbG7XvKIhwmgSQ9q8mbwlwC9
pDzYpG6J66+S0ykWrf99UATFp2ERiSVQuk/XeU9P9m2MsO59jTWUTMFV6kwq7tLHAOVEzoFkv//I
Tj857H+ki3DHoz7JvRVaOGRB8a0UceV8ObFKWvHK2tl9i8UI2SBWpsIJHQeVwrNt+iJ1xWTTy7hO
CbQXyEb/CRkg16FEfRx1dzmXF5Sf317Bru/fGQ5Ki3UrV1clTnb8bouR+ZCeav+A2wL+ryPuRosc
MML3V15Z2BmhA0l9Hh8501kzRP+5QAG66wvpkOtBtS2n+QZVUbo435hWJHIHFGI52nRrr/GK1RGT
VsOpezruaAIixIrz575RAVONHP+5xl9oeY/4n6WfIK7MeoeLTR8usIWJsK9NDkR4iyplOyADOEjE
8dRXlxr/nGQrXJDsCadFWLuX5Vd1QYsB+QKKLpVq8s0r4+juQgj6Nq9ibZafrMB6Be5ygpw7rQgW
L+g8xLdlPf5Vhf36K3aa2HAqVbdoMUeN+ZbcYKj2DWBhbfnO40vUU1FOxQYVoGP0fvw+8wx5jJ7O
7KtKQfs9qeR2Kz0QwmiVww2j1NkAfbIR5DJv19gBOjcsxXeKG68eo/NcfUWOVL0ghNTes0gYXkwW
/h78ZjqJ8AY4I4yDikkjPuJh/WdKi9WF/smDo/TADX459EY0Nnic3ydh1s4jLYHcMHb8VZP0PWSS
PkxWAzjtgLrLzAC0RS1NwnqrCT/ypKq7rW80Eym3r8NVxuYPdIT/RFM3p68TPraEWlPDybt6RMPs
I4yMtNA9R+v8VgkCYh4N7v4mAhA+goQPO6EJKUYEywJrycYFyOHIrvUt5hBIer/t2IVfWDuxDh7w
fxzswaBFQ3YHfjFxJNWNuLPazJw3aSqnoCicOyccSLGFXMaloWMzT572Vh1XjQ8mDiKIr/mmn0Jz
GmrK6a7yoICzz2VG1oJ7EHREcxd1D62mvaYeXfT864fx4a+taKUpWcGdfbe1SmVZkcudf+rMUYGW
LtgA9Luj/IkzxxEK0Qk57RRXzu1uoPSS3ha6x13cPkSagsKnKkr/ns1rlrcc1j4U5nQg1sSAdP58
bzQ5v/O7paCwZRN7QwfPn4Q7PoXoCBdwGP+QkWlh7vVxjFalyKp8F6dUWHFK/ewjz/y5j6b8cYbK
3CgjdCyvu2iJQQzTYDSELScSL24yX8Ko8XrigHcha/tJdfN6QSPqTUgnH5lEM36QIo/NMSPmr2Uj
NRiKyXnN7v0pXgDrVnaYGhJulTkni4UWjzcxABJv3A1ERZ8vLuZXCxY8Yy6YV1lhHSniWezlTV+J
Jz2m0f0EFN8l+qlSujr4Sf549mXsiceN//m/7A12bi+r2QQNTPwUAXroITH+Eq/QA82rzzhNPfku
CUV7xCmvSK82mIW1aHJ4g8Os14pYSQJqNiU8ZDeJAI2tQxpRMKLaJpE9cfGl+heukmQxpj5AcWmd
E6pZumtL32hNOQ3s1isd/0ZxPgCnC1wD9r16yNr4Y7yzB9Akji9BD3+5Qndif8hGBZ02LE1GdwLW
JuKM+0AXwK8tEWhZ8jAlVlGagbKaQqlQGu8p9kG6fRmy7Ov00sHU4rCok7BRcbZI9amvm0aaqLF/
dQ9uSPxj7P5O1lpv8Tqv9X4O3ASnUJLJ2fWH/38sWLyTls5IQXgtCe3373daToQh+OrwZjJluxQh
yiC9/Y+MTHnWby4uKuVsNZQjKJ0Y13m2IMTB1X+dU2o6jwEtJbxdgI32yPgtZ63ucuD8YPDS6qG3
xeKXHW+H7+jGRhUQR0VlBltadrzxMvvxsxmfYwbQtgtGzpYNHb0YfddLB68iqu+7wS/pz6zAu5cB
WGcPREqj/HZK8DfSZ7/Na2GGCLReBvZQb7/wk4Dh8+h/WHwLRpGVpMylapbi+HzQTM8N6B9Wlwrd
4qNfpPWEkkZpC1NWDO04YmwngMW8h5Yf/MCla/Rrv/Na1kydg35BhO/h0Dzcp1MX3rcRdefCDSVG
9ueVnkeccAfu5okabBontQk3m0uNnHMkw0cnay4WyC8rg+IaM6ZQIBrU6XiWtFUaWyidCFG7Ro1P
xy8z6HJOV7C5+TZMtfdNOtnww0FY8s4RYKkIjJXdfL+xGPglAejveApkE1FyAP6Zcm18JFPoRpf9
5dL7GMa4GtYXZfU6RImTNhfx5YVwPRIpqjOxfDP23oMjRzrVuELXjxnH3yzlhwI29sK/XDjcr4ba
PHUdHEd6XRi6p+RzRUqv5Lg+LaU5M1/zx+QpEJitVNRHpqhCpWvR9fli2L97yXtvStHeYpy5J3bY
LqK6nnaLk/4xzz0G9H4K0ikVxdxvVmUXXVMzBJiGlz3oxOzBLDiSVUeqU13ySME2rfKju9rLt28F
+CZifrC+0WgzlMEu0pvbbupDqcqXN2OrEUMdhfwgRx+V5Ws3HCrAhZppMn7pEKkDCfgzgtUeHXLz
SbdTDvsp9UgGwRJ+j8C4/EllxX2kS6U7nxPnQQyhOnI9QVkeT3Ye7O319pu2L8fseTNaZ6j6MJFu
w9ubrQSxIQc16+vHxcPLY0RJDpTso+0bXoJbE2KrOtcO9iRvFGFIfP5RoQCGr44aztl3N1YPEYSb
cXKKNpZrhReEI5MKr+XxDhsSaZO0af+w+H0RajLHKR9IgQpLmRrfuHfYf+ZjbKqEIS1+Ko+/9yEC
f0clSdsk8mJaXKaEtpbBv+jfbbgghr67e+988XUvvDB7PKMHHN4azkO1i6p6OrLCgkQSVSHqToaK
sOG2mzvwkpBgyvS0tPEG2+6x68jB0NhE5o5cY4ut53BG4Fon5ZjK/9QWWLjZS3aV3NVW05obP9Kn
9rJZ52LH1vAz//Zd1JxFB7XxxprEajapOalGLElpD46GzJ68TSW3Z+b+IWcnntSGq4uouPR2fAB7
7cJO8kt0dddB3rywa9p7+EmLDdhU/oSuJkxwlnWQuO3Zh2jTemeiSRFkgrlTEU7N4Y0EbGvxC4/t
FQpbi6kr/fVgt5Ael/QJF4red5ZxNQIaM7t7yBkXCYTvjEd4oXkI0wIKW8+feo0Om+wiglkjjbTN
XO1GwW7CpzqvgMDEQriwxTxhdoh4cDcFIwGh5KQp8XBcag+NMUbsut6krZ1yHBFeUZjlN+03+J2P
hyl/x3a9popsN3/JVvf+NB7C69IEUo9KFDvLZvCQt9LO7LHQaNxFu83u6bpjVwEHgOT4Mw0B+7az
4Re26RVIFwKaTNGwdGSd5nq1t/kdCbWx7kcOsIh/lS/65PFGcgf7RCRO0glEM5yFblJPh9sQl2ce
xocXngTJGsJnXDjpwwQDnvig+ydwBQStYxJXArSEHtQTDZ8YYwY52E83cyTbYePeWB1/PGYrDIdi
U/iCV61O2NPFSBM0y1SrQy9ZgfcXMBQax6aOsVn5Dfs8tcchQhQjKqjKBEEBK+Kpth22d63+SzoV
VjZyMd7vPGoYa9DsVCjdFtTiGFKbRQ5Jp8iRfY3T19mZjcrpWLpKCQ80Ra4Pboaguoh0UQPrqdcB
3cNdqTaC1FEPhmw12D4F1W30rY3PsHmWMFz0qsO6R4sBL7/yocEBWPRQ8Xoks0LyANeEV13wHT8u
LcYLNNXOQrnMZBrFbRTd3lr5tgW1qz5TOxtZeG+2/zAhjXpdwYI6n7+xBhfJY2pds3sROxxv1SGR
9+IKtOVpGOevrO5mG1D1b11kq14f7cRPV5+XijX41TNrZrk4BrJPsG1lmgWBSegSI0cbDCpubsbf
VHaomgzsdtQ6Fi5Z7ROM2FRrcWdxuS67SxJguBivh9VM02zxxG9BGaREAdacz3F5MGV7LWGBQlhv
4huSLRBRa3fAg6auo0mj3oP+0gp7sEDBrWq5OT2+mkVkE2TkWoMoGrAMz+o0+6o/mi3ojcM1mS25
Co0qFOejINqsco5e8IGUssauZhfRqGQrxpLCcc33O2N4VmZQaNTfmAIPqxX9JRZC1uHxOhYU/I7y
53EJWPZ8Q4L7MvWIiBEldKYrY8qSCnmBfzhgscL6buY0EPDRknWx2h4YpbBqhwejtMCUu5Pr3KhD
9/JGlpeEx71eVB3USiQ4t47LoaeFC5IaqdUUr0o8rct670IQocFgOOusdjBhfJz1zfUd/4HFA9z0
Ix6LNVDG/PEBhfpno/HX9oVNn/Xp0n17MJiLgvTcrTxgSnJ/Rim1n7J4D4Ul6GpdB+AJGq1v/Yyz
wh//ynoQJ0P//8LKla7fCzOMCl/W7xTfcW0VDzFlopWKufj7LI9HqPVd/9Wt2cVSH7TnlHnmvS/e
4u3SQ0DJut/u3dhg0xSWWudUI/o7TtH7gv96M2sxMP64CY2fMVZPg5kOMJ8EFRlAUSIkFcRoB72+
lbzW10A0iYlydb1IX8Br/JlTNeKbrbe2oxfUOZi+59NU7OQCiKenSyYMlfV6bL3/b6GyvV2FooB6
aQTZ5RDt8NGf15bqbdSbqYbMOH+I4H647eBfN2BoOA5AFht55nDkGR4ksl/9JDjFFb6+49IuxuXK
L37XXT02CsJsVtkgNyWR+/1p7x5/okCopqe+0OYhrDA7lCcd+LDhGB1W2attcN9GqWoMg3tUhp8w
7A/FUfNloycI0fjqcu+bY6Z5wPTDOYfXnTaeykYD/zYpu+oHChVz+AmprGB20zncZrD/yEOR0gGK
iAvaGOjuEC8zrRXUHuYbBJTaxHMe97Lr/ySKtWXS1PbseduLPN9NrnBxxGYAnrPVNOmZBDlX9JZi
zJnDfDyH/hbekHiBAq6Rf4eSCVsh3bHhnVh4YLdPCvUlKjpVgQ4W8KKn14l5hn5zagwhi/hYZKj3
VfObOj2kKiOLHFThDs8qxcnbMkbbwOaiSr2MaFz9/xWmgbVkATET5ubi5l6npY4HSgWaLBOTX2r8
igc4uKGfrg3NrKQXVUl9gg3N6+c5m2nDWyCAdzea+EdVGhNqKYJeDA5HmxEdidsmEUpMGjmvWSOX
c/nLtlNsDQ7cMpF74JC45oBHBvEZjGVEmIkDk/Prm6yKcMtb7ny/TAhGNLt3wVO0e61wr0W356gM
/nCRZTrxTLHAxangSwZSPoNknlAW0Ghl374pUKf58zB3gLIEdAckJGhRmwTGVHqROZdBR0BWnYyE
JfL8ANZ8QvlvNeMQJJRp00nB6XxYXylXD2GRAWMthb+evjq86M4jk/gowR9Gf0Yc8H6T/XMZNM2M
eIR4ViQ40UBlY0nt+k3kqwjlLVXXCN57RPcfEMAtvNLGLkTC9jpmZoMIpi1ZAfwBdLpaolsXXis8
Xf0jMAlEKav1V0Xeoe2lglwOJWtQPX89PNgzF6zy3d7GZqfTQZzXONxTmpXYYzFBHY4wb2Mwvip+
F4WP73fM6FQZ/Uz16HXCxMJ3HhWdT+8LnyroYMYKjzQeU/8G7PDR6P8OTYZPCMHtA8CKsooch7Dh
REMiYBnP+0gAsWs0HbQ7fQ6rYAlZ9VApdQmJJYXQCh3z+4qEkJOxjTFaSMDzlcgdcH3y83RHKOs+
6/xF74QqZ8zHAwGcPUaa15xWIJl99gB9ajMnSDs9K7+yh0R1WL6pZVc2RkyeueH3cRT2K9Mwl9sd
YDJ0XujJ8D2oUDA/6X5KfTvN9Z9eyxMf8oxAs7pCpKHPBB9/e+zFghBxtL101gWKgDogWIXSA7YT
TztGwvyal7xVa11K1ph5RwW7fDCW0cT/8QJ5HFWupmuwshieG6rmizHI7R0YxcSqnmT2mtRWe+kH
Ga22DF7aQY9o1SRxNRplapNQ2SiP1JO8hZ2CFceU8rHoyOVLjP8PaLrc/gsFhTL3w4Kt47oHePlR
wVmhYoxZBAkMoKhoxZo5ALHdXr8MMe0wEYEPWXiGbpUHu92qbWYDuLNosEvOv+YezYTWvZdTKmZz
1sbwkSI6cVSP6yrxKUfhwYP4XtXI9ttftsdjBM/29D+mqWV2Z3+d6n5k/42ndRNi/uxF3+gQu4Eu
m2ySplBEsbhZun5zW7MPcFF+XJT2RYAFkEhIlwj05L1/dBBVQHu+iLUbI+oueqzzulbpgcYajlfI
kHVlpli4UrlbpYsIFUiz53emtYVKYhMoBv+AMB1qdbf6narC3toUn/fGUqkoVuc7d6aVSmUWKxMK
THD6hXrZ261xmV980Qgw5yVjzVVkivkE921h2RjflN8jcyheUDerKO42xMRFemFmrHrHIT9rzFue
acOOpwUvmdOtNFomcMQU37UOL5IuIYKgUYRLRt9gKF6nsZpmO38EDmIoy7MpwRbm+dPJik8df7sd
ZrJXtKNs1Ds0KmL5HCLJuB5Z5QVlXlrpILgaH5xmZ+NImkTGnrdcJMXIGEgNnFBsR7cdvUh0ty8w
/yJBIF5Jq3fBIj8X4bvGHtrmpWH4QJJNeJOOwzbielCCgQr9hD5VX8+Xx/332FsMgOCenb3qomxA
0/YJwedHr8h2RzxjufCQLmFlcuxnuQrTgwrZov3ptLJi/bMYdINBirJvdlhHKVFScBvBd5VadQGO
3yJFL6Y7zd6Hr8zWgRRExeSfMtORd+fGk6z+z+WTaWkQcjmSuacn/e/leBBzdYllRU8b+6QN4h8q
xcDOBzi66KagDYlQcAuPcbpze/0DUAZiEe2jaBGr/L2QDpRtN5GVS8wtMCwmK4s12tcUxPhogJ8F
rNLecPg3v0NKFA9JSOauOg5/R5wO/UtiPRN/gz7Ehga8mP1QP6jQzJOE5rur+HWqv5bLKB97DGj9
rZBSzCD+5DrFN4PCB4pJ9W2vQwqkl/nDjjm800FIEEAdvGFsw2AEcCrm8adr+NUvBeTmcLQ0H4yF
NML3vn1UGZtTb2RQ1VkXE6poeUkGc92wxlFXCaYUAl0qPW3twP6ZcxLSC68KGcODs1JVpp0xX0Qb
cL2zpLinCDHRXiunIM/vwVeY/k6jD+6H2D+1zE/UcpRGufGf/Pg1m0Yyihp8SXP4CrT2LNGb2Z+T
IZcEe4Hh2HLs14nAxiE+1l/laZESxA2DB3mQCpG2MIlosdxn776rfbQtwgpLTHYK3/ftEZKTO3wR
HbznscCul+xMdvy8ojkCKSz650lA4zBo8H5bRxgQwgMI+IHE/HXurxovyRCrbys7EolH4rw2ctSk
Komhhp0U6hEpTsTyNDbM4v0+DHUo9JS7KMgSWYyEFhrvRzF3229l60fq5wO3hXj0DvHmQlB9MINB
Xmo8Yux0gxHpKrp/EMBgGtJx8CT2N0RbmSSdjx9V2OK3NQDE7Uie7/3i/3CrSpADmqbSiTPvcynz
1dAvN3fCNKHv6Lo9w8nvM7pDWhwDJ4vo/vARUxF6328uK6D1WVe9IzbOm2FtJAgcsOor9dFjvxCH
xZRfifxqBm+/iisvWdApc6AsAxWa3oBpoM9yhsdzCjj5JI+r1KpAzxGJ0cArZJhzcs65yNYg76bb
ikkCbYsnIEgl8qCbJHEiMV3j9fV6+m22FTP+mk76PMNLF7oFT6iDQZ53D4gZIReyTR3Xf+yO0k/x
N197Wa2tFT/PbRMq2djDfTk4P3VQN733J5xj2KBxkttyJFTG/MPEeH0QK1fidNNAqqyXJ94g5KCp
Ya7WcC5hGutDA1IocC24FezK6+9SwY6kU0x1JXjOxidO4V1fd8g3ICBuA4DzTNG5J/RiaLIIrGPh
x3JHBdOKF2RQMqKoCvBRHS856SFyKwd1SYFxWoq+kz0d5R9rvLZ/GlObxy020uDDlWSNqLqof0zA
JnlS0/wFl8zinR6u6YH0AvfjASAD8UXik60SkCUDX9VD99TwqNRW5E5bXGcBSzxtwIe+DDw2MSO5
AxGw7UHbx7Ro91k+39cnJPJjv2MYVHyc0GYrKzpZ2YWGRp7XysLnWBaU3Ftj/7D38CKKweeIGqzy
yP3tvSbIZqN+TXti3Vxatu1p9XU+B4BWIEGfUTEJVguwLKXcMR2MOfC5EOrooO27JfBgyW4evXpw
UvVHo+hsGWcdp4SgAcSOXvgkXOSUJI2IweH57/AyaQlWJsJHxGQjF+fXSwF3O5Rx15Q4p7iLkFkt
j6mXj9TYZw3R3zUWmLRCHd/N6jpAiERtikjUZrxP/YpMeSDGhEd29QcZPQb4biq57cNQnJ+D+JVv
joyO5Xrr+kZIMkiqw+gZ6DPGlOC975Z+V8oaWb6Wh4F232VrGV5GmTczbNbX0qTqubNuiLRMfsHX
/xfOVwqM+u9AyuJg4YXr+eW5ZnR2B86wz8dEfu2aJUikMdgeo2mDm0+mw/rH8w/ALxtfSw+lySWa
bliVKAil8lWvDx6L9EvlyHGFDthS2Ow8tRWZeeHgQ55EZR6O3lCG/RjffEVN2DRsTGNlsX/Iff1/
nnHsmTSqsNZv4FT8OgilxTxo6v6gwlJxmFXNgO2zrmsxQaPEmbSLPIELNMVecumx6PPg8D/QtMh4
6sJK+Y3bEjIkN7oEKdwVR4qEeqsspWrfI47ycp/yjQPXIuUWRzdgPen8qu28QptC0rCiPuojWX9J
wPJmTRHZeNtiWDnT6y4bm7NrHyT9hJ0/LgB9NpAzRzmvv5eIdfjgieXk+jSH0Kh9lvASgZv0gmR3
aAzhGXfl0OCfJIWlp4kIluyqspBRa+KCvfJrbyJqDURZ+O3QBZthFzOYiO9nnwCKKbZ9UaHxVNBm
Vg8kTWywpH4Yx0PHYhKYSiZ2Zn70cZT8ZDYeAE4scPveFIbkg0jQLBKEUSQhpgfWqCNtaeTNPvl8
kKKg5MQ2qBzA4FmDp//YgEh6owPfn9EOar05Ov7pG+quWZ/pA5N9l+pGz+4wV2c4WmN9lxmaivHl
7YlthFB9MZtjIpAW8UdL9wmiQ7ir5PC5OLu6pfFXDoCNt9CknxoKxc3gBVbiejr7GmjaYMEaS2eN
zTm4docTDuqe4mG9/fveAEO7omjdjQ5FOUP4MWQirS1J2MsB2LQw8mBjelHyjr9IZAc89CXOuw0h
Gg7ICZvZ3KtIUx3MW1xzcBpqpf1EREKUcwz1Q/ViKuo+WB32qYv/So85nEb8RQKIddjcP/Ls2lTI
Y9cPZnIE2XYE+J0svan0GHj/IO0dxmnaCYpiEn/QaetzfLqrNvMRy3Qko2ctOfkG4hJfum0FFyKm
yW3lNBLNDf4jxn3rZwMmzgVu5Y4rdvruhFdLP8SMi7F364Q6HabbGYNpGnzSXptbYUFAizaKS98X
2aJLefioVBJJICUTC7Z5JhUhXwBlkME9UOG5ikk3Dpmfp/51T/JkOgLR//QuKhyCXbiMfxnvyznD
m5O9TrVKJX+uB8fGYfoB6dV/Q9UjWTOOUrTjOsifhj6p7POTH+D6fQV4+6Hhmn1OhBYNAf5g2vTz
IEBVEl7VTrsBRPs5ih3Yhx4YaUR2zRrSx28pb/lkWJW6DaSFObcFxcpij/4c8GemrI/4ZKzlaN5k
slEF8MP1RqwqjH9/PIeisiBaCYeN2QXj2YpvMO0kf9RKipx3P/JTxNp2l/BHDDASq4bnM8zOVLeK
xhVaSJGzTLRsuSEQOi/xU9Vv80bkbx/jolMvUIBewSSN4iftV0xktRRCdncVz5ZMgJZNbE/yY3hz
tECWV2j9RXqmJW7WiadrL6MT/vDKFWjfN294oF8G6gsnNfO0HBpQ2LT1+L7H2t30NWABG0Uii7AQ
tZ6TFYhxblA7swjNSLghI+T6uVOYj9RUOPJRiMXe86f71/qn3h14071T25nM+Rw9cMxeui/STeGJ
XRFO6Hqqu5tshaGswHGRYOnZsMHrFKlx9EDN+50qD2XQbfU8dJocz0aGFR/KMCKxVzz5xjuHUCG9
I2OVJyJSBu0ac5lqD5ae+75VsKQtAvi40efQO2G9A3zUQZ3YR1bzTcvjHw7YV/mlejXkQThIqcDN
ioLWrVxpzazSUADc4bR/9LqJ1kp2uEiUyzxNHquEpbNvrUOMj9AA1qu2OzolzOZgsCGfVaLM4WR8
GTu3Xzee7kr/VMhsx6sJIJyx9L8ywY1NWiHjmgUllNOfdERW6kiNxTfKrWKkkqF3J8LylQ73njEz
WM9+ZD3+EUE5SAaY01zMl2i1ydUqR8/pTL7jjZLui73B35gNflpOjbiLG2fy7fyuyKHhjLIAN/BX
Gst3V+3x3c0ELo6F5Oy5uQ1tp+WYGyV3rLDzUqBWSH7GBXhdKbrB9FPeQzQo2cvJwbmjGgYp5P10
9UMpdyrMe+rzGSjx9/UOZyNe8EUp+zHfEpnltnK6q9U3N7u1R77FHySKBkzT9yKqsApFOcRgElUZ
C5QNz8OnjItBcny+OlEz5gKaRO0jb29OgEGMdvQNOs+siaDo9AgxKt5TdjqxqlJgqSz+VAS+taBs
3rjI4Slx+LH+lc/6HPhuTDFOBkeEZHnJflty7V/7IMF9WnV+VeAT7al4xXBPXRLo6fp42+m1l6yY
k+E5DzHqqdUidgHjT8wH7eqs4rVIhkzMKev+fVszOnpKMeC4qAofUbg5LS2/wIjdgWUFd2+RFcRJ
9udtnP36RwC8aksn1xmdOwkK1iSqbwTzqHK6B+/yTcNnX7njLpa3gYU1ECZjHSlZEJvoGKIAzdDF
zNID9mthuEbmSc859qmokN1kaFfiZwTqBdrov0xI2ysVj5ZyasHOIzfg30CxZ8l54DYVJLPGT4M9
n/hWN0YkNrO8tzb5lZdtHi07TSMluQ0/Db3zsntW20zCp5thbdRAlVfPxpZWx8RsPpxFEkxlDLaB
Gl1t3yYfrkb/pzyGrH6Vb+kMw+pzGXnk/MWiQYm2gEJSzB+CPmdExFiig6Tt1FeZgQ97/oHvew5U
ebOAx9OaLwxG8ekojT5yzo9K1YopQItcuYvoN1WEQOqcnXPxpiDvGIQw9He5rtTjLTSRBETuSeOw
QzVwTXm+sIhz/vkEFn9tHk6yqiDyY5Ne/13/D8LON3K8aphI9/CxLcQ9GqgF39iup/2rtqyi0uxt
CvqT/IwmMKpO4M760iBUDDWNZwNSWJxSuQvtA+wgpDUADv1fqyzpW0Aw6nRBuYw4oy9+QwICVWxf
3UA5/mi+WC1GQXVNFhiWBJh/tHnTTU/l7H0W8ejEa5ckxkhkdN7xMCikBoIvsZyjY4Cm1YD+rifo
FTyvgtAe78vEBSEG2h0rZmgPoHpgLlE2ofEh6kgPPE478rkDHupAcSL8CHso4aW2hC1Y5yHPbiug
ikZNogsyOe4gRm6d+LgxUnXk7XEPPrySXkv/I0DgFnwk0a1BjCwMlW8+KA94xQXtcUavBjz9WgN4
CCoT7OTnnfUkZzJ+ngu9PB0SVK0FhW258tHQ3BurEucaI/blF7WNcCg9UHubN7eIdwjumDehnvuD
mByKKfCuGZQWi0FzaAbhOSrnuQZotWzeYxByNrZaDlBJkhDYKbNQJw6LJ7NOT6mzKrQ7qtne8R26
Ak3Gogefk+oDQRcF39qqT9vPYpDRXWuXsp/HUDJo0zOf9pvwlF9taMDg8UyaVxpT01WQDa1V19Mn
iSmGYib5hgybeOSMjM6/lustMynPhZcsxJdiWoZ0ZBK8ZGhZHxDF1r8t3cT7/y0GnL4DJR3NLX2B
AOwK8S7s1eJwxaBs7YwB/UTaGoPLQxJPen4z52yE1Hh6eLNGWAda9Yp4F0SWvjFZJhS19aXn3h7y
nOk6QDM50Di9ZiG48hKnSbMInq9hY4mXJE36QDFU0N+/zZpmuPBldjZZA+FvXbSwSRvHmuKSPcr+
aDOOhqQ7r1UmuXyXQk2VN3kOPRxBzwBmUsIUTKgZcBWbAxEXnJlH5YbXcvfFzZaaI2n6i2sZXO5r
4GVl2a4wm+o27n5UHlX05tSeL2tyETjBiYh59g8c1q8rvt39XMjOCntiDlpuSyyruJfHur7uqU21
JF5lNHVetFCq4D0+EKSKaDtSgnpkR/0d9KEKFhyrLlpBq9NkARU3WEdioxprt30WRAmLuBfoOXXz
85NtWy8d+RIzKeiI+L3FfWul3ipejEuEHejgT7i0l7JGvrde6v5wxO6JHoZyDxcg+LfcEU40ROIz
aJUqVl6c/bHpuwrRoh7YOHAul2qIn/A5UWqfjdf2R+7RW2hETaY0EIgCQWPPFK89yZwgjdFnPuc1
G1aSw8Uf/GyV2HYv9yfU3r75YGEIaf3fVEFVVu4HcsRY23X4O9rJCO5LSrNeubmk94/KFPCZqi3y
cYiuGqcyGc904WMqxXX1gqYvP6g01ZGAIMMcf4dpqXcZdN7Hfr6eBil9WB/7q4WbheSnrsFS34vF
Vtn+dGUW+VwEJOsy5MwnzSfODU153QqSFFAL5ilRUMiaswu4A9Be4IAg4WYRjY/eq3QuYuhTxiXJ
dn2POTGkGJuFhe0J8MDBkmp7dj2oyI66NE46xN8DYOm6wFU14fD45/vTEypsTZoXz5fIyvUyc1EA
MZT02O9N3eUAO5xHfUAYx5fjkB/zTBt6jOOnhTcF3SWC7AXMd3+9x5dm0/3uZm7Xdx0JtEYZG4ZX
K5dbLoaRaKae19Bus0BsmziPnDpzdDRlhUZPz9quojst89yZZirG8jcfsyCLBXtuo2vN1A2q8Zvp
iWi/FeoE79Ym/GUqqN3XIMX7FTf1odPWueVHefumqLWbcxIx2TRddOGsKShs1WEbKT2pBPa/1c50
KVrQz2dJLgs/6/HL10S/Wa5/xgeWqWIOGPnyfwzVbrZW2Xc9ZaNPGHRJZo09uJtFdJWc1wWh28fu
xQoEwMWArHCpikCgEUh9uMiOqdMh28n6vAe031sxTCxUZwIRquUL/9KoO1PgGh4OPQBIKTQY/mvn
CHEJwOBHQIVl3MH1JtZWFthVPG+yAIvpBX/HueZssQJ1R5p+QbVJhJFuI/2GbYWDfGs0dwY+dzbv
/rn7H9utStcnq9unYC1afxnobPC96W/hMqeBpNGA3KH/HTZcVSMq0m+wZitguMDG3Si0EE0wABOq
8tUKYrzUDDm3m1cbQ+kifa1lp0qd3mHOaW5Pjb1ua6AVeNwy79GlIR05ZL/rs9V/qtGYRJ2PNbjv
5F9bhlT+o+MtlkisR4KIA6giZYv1GfAU/pI7ENE+EKvJcRQ3ZKhJ08jmMOmAHJArEEK9N03HZVn+
/zTFyMEkNyuQWf/y0YpABn5TwuPsde95p0aj6TxJa2+mxLx5z1zcF7tHjYxV56J6pVnegFSZv3cO
wGBJkFCzbVdk+/vWLT4p/ThgR8mjpVERlnys8KAGD2PKSNNHYcW/kggt0Du6WZVXbPuemCh73p6W
bkJ/j3I2Ra8k5j0qdw7D/Ag6C8/FCrkfYVAknlk1d54Qod5dxPodQK8O2EC/uJlDrRdPn5H+L5Vi
d8fnpQbVEnxuC51W9eS8xolMV3dYsJe2s29YdE4UwXyQxZ0VcBO988L/UJ0VgqC3QLSrD/isSrEM
/H3fzA5xXRQnhLbA2xX45jkOBdo3ofOUkkC2mvjfzmbONmG32hNZ95LOw/cN8Vow2W/TD6b54PuN
rPBQRh2pGCF25ozpNcmRjYtBEf6ye8JtAj3lVlhwgygMMQYJjWUdEwLyd4vX3k07xRHldTxgTRoe
Z2r6cpzEi9Fcy/D++lHllIex9GaJZl0BKWZR3SKxrzXv3aeHUuYxuFjk1QhFPx1CaCOgLA3sfE6+
GW2kUUiR7MjqVgsSEGmiK3fLywXeXdYkqFuKefOiyO3lczD6tYM+Iq4tR5OlxZd/3C8kbpSdAbts
6+bU5ptXI1gtk5vmNQc5F9gevclzl5c4SlTdFeXBU6KqmsoJKyIQQyRcOyitnfBadDMVd55llCWI
6+3snBxdJMm/Fmwp+hQbqImQM564fWJwqYs9yq5knw1vzBBD5zglPZj39NH9w305yOxTwjaw/woK
eyWIHDtnjfpUoA+MnZHpSHcyH6/JicXkXbMCIu0UCAQL9RXBoGklrYE8nBNyQkE/aOLKAW5Dl6mx
95vNQJCzIUhN3nIYPaW5GQeKPWcMBAAAdkUfUdDK1vBR1611sqIW5KrjVf0UwLxK0DAWx7hrrwjv
Rgk4eER53hmFayQEvprPJlloq+P1AkgU3s7+ML/GfNDiMiL9gkpbqtt4BGr0nBRoM4BVECOJat00
hqDiWndsOs/tjUmfpLWHRf3A9IiJtg0vtOUTShIgW7v9+2tlHGN6ue/PcjVnaC9M10oditxJ8fU1
iKR4tedP8Scht8mD5ujVIjnMEAVjQA5D94R79tTbmszzzsm+0l1S3BSde3hveZ0RYxnOcRo4ZaTO
5bvFx854eqYuuIwBMvE1zr7JQ/cTxeechR7/25PaBT5TGgLCmUSsf7qOgq1HtAQgy08twXTJyxcs
J8LbgTxhVtd8hn/rbNaux4eyTf7+hZkWg6XWyyE63EhA88C4oYfTYtnwT+zlTrFkj2Jm3ILpq06k
TV+EmxXIoexLNAfa4Icz7sjKBO3I+gz0jWiOvAR33Pz40fnrXvajXSTWspDOeZHHi1HxMaAkfWKk
s5SO/WOmqeZIsoTbu0//BnSQ7qyuqGONyq2myDuDTLSsjSgn7KodP51lssD+e/dEQfzypKsLNvuN
rh9u1aS9UvM7h9CSpWlPkLbfTJaxPKm9ruSaqcqoOptqs6Zo/4UGN1mwvNnLSuE3psFFcThwgXoL
VDOR51CSB9PyjqOrYQNHTNJk0qcSCNSxCns4lSlO3lKPmfCSIQotCe8m+1GK7K9VKupS+hFXgfyA
5WvLHeam5LOhpfwk3/V9iLqVpWIgK10OjguwG7UTTE10CaGayrzXEyDOK+KKOS8ZdlVOtno76SeG
KUtDRFVjnn4BevUZC+9mAzLfCpx0bK1C827TdmUxEq2i2lzZxicpjDnImTxfSsDQWeR9TYTyALJU
HSZPJXJTQkBb0xofHSN8b6V4Bjrr76dgoKzn62NSI62WaGnY+KwQI5DLzCeyyNRghR7DKuyRTeOR
iB5rQF+oX6bJtDG0zKSuPWdtTzmL7FdKDtbd2Q0zBvQAxVEXGy1M07shAZuz2QET1YlPo7OT6CQ9
u06rQWnkjqEwwb9UEFk+PPDcSOyHBqOE+YvYayBAtcyg+bqAqrWSO2xDbw4wtJDRyfXgAFaNXJ6m
SC2XY8c1MGWFJQxhQtQ6vDlGfjB7IJfXPpBiqszul/PfmgzY5XyRkOFpTiucdYlVVIqJ//0u+VCc
vb97nTRvgVoXW2cz+r5039MavJXcTyt4TmDiGRMN+lA6tl9Y49EvPS2RcDS+BA5BlRK6dijaTJO8
BDx/lcFs6hubwaMPXVnYgDawX+2VnF9HEIMBJNXlpPo4jez9NjAv7X513KK7aNslIZxFVNLrv6zt
6+cy/ZaXx7ich9XM6ePjp6uF/oV2RBDQk8C6Prgi/njnh4ZRoO5DWlYheyTQQkGgpwlAdJObWg1T
3pX33HB7PWQ4FYP8Q4+RBKC6hQNkMjriaFiw56zXDH8Q8aroEZknonaryZyJwXKhlRw1ISXIbHxp
3MH4mfweRscl4u45o3tQHk45z2J4ivIRvIHBmSgMpBpg/fqcMkLp4curxJ0skF68FO2PWKU3KeK8
3UkSaz4xA1+uVpxh4aI16G/3HRjbjo9od3uCJgpayx2sfdWS1IqsKMa9ttfXfNt+WehPf+PGa9Qj
eWjCYFLrPfy6vwzs7uUoTT6BAla9Tdk4A6W6Z7swsPd1L7C0lnEXX43tSe1PQXVii3XB4b44ZiAS
FBqIqa2InE5JVPcOC3RcG19SL9J6o8P2FQ7+eqMe0JTeMCzBtJf8RuPejnhM4phF0o8GUjqJen0f
u9JhgJI1NxyOJVRnP+ijnH6/YcQ1BLeAL/nsD0fqZ7IP+/8FceupLluJwyVdCpFajtbWFb8ISYxq
6Z9dDNee9/rLi/DhER9Ga2GxDWa8qa7tPanmE/RjR2MU8hQGwhz27q1j9ERF0sUGMD7oQiQpCZ40
PlQAitt9gCCUOQFR+nRVWXKx5oK4egu0NhoyIHZ7Yj5TgVAvviDjR4D+7ToxvYysT8UC1AiWxTO9
UvcHaoRMiWv3Gkr0ydOw1s6vpoSSyvQ=
`protect end_protected

