

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TPzJe199hwacfTEDRpey0Y5untTvCHMOc8UwVOHgOL6Cq0y29P5+TdKmR3bJs6CNw+Z8r38Sq89a
ki4EJwz2ow==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Drnjg+DhvQL2SL+KF7jJYUWbmCL77tWSIqOGGYdrc9R0pgnFA8Kf3gPS1ZoSxXPhS6c260uxbqLQ
PWVkxuHyrjCIi6XW3zOvd7Hhd6ognTJsTpAQEXBbU74AiPxdw4jvEYl1sM+yQfcs+vl80X4HygYq
KrTPcG1Be8KLudfbfTU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HWZozT5NQ2rqxB+k9Crrhi0GPbARLZZeH4efQ4PQb9QPZCIMPzxN7L0s+QNodrL4aygQDpi786c5
CqNe5zWKd0R9Gau3AnPiSVjrsD+MuX69q/9sY0WBR7q/cfZSBGZIx3YmVbyWPE3keUtDmNcNr110
O4u8zqFapbYYdjj7mLVzjL3kF1t07LKeeUSbO93n1VCfhG11lGVoQp4l483fEr3qPhiJsRENdSmq
wHuNzJA9YkesYjWoIezSN7aSdtBd351DDSf7hsi8L0UTXIWnRxwJt1nvUdHZGPmrdYZFVYtgkVoL
Kqc3Yds+bnW4w2g5/XKoCvlblzUEuimUEZb5lg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PpdM9DCbKoehsFWcxEdjTuRyDv7zUGcQO+8GO09CTbFl26DWCuHpm8EV8DoYagqT15HBgN17MAKc
4j3eHGyE20UnjU/j5QLshbYbE34D2uYFsm39cAXVasPa9yKzHvUPTPR/xOAbp+5jG7Bz5FglHbTs
w8l4ypT7qxfvbVKXpJQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PapJPiqoUoocuaPp/UPL6lvLFS8tFNyQTHSf/bfcUlrbN8RMO6tg3yW66Fnjr5uuUT4gweeZp+ab
bvOlvYnqgmUB0QtryXCl/X8jtA3Lr8w0XR/TABvOVV3x4oiuUMIM6iUjigsxYx5tQeU4dlvgQLU1
/BQkEakw1+IXJdvjqhEY4vwQWWNrwpILKEaELGlvOfD2KG0IqRnTVbIMfs7U6TK+tVivqTzbGTU9
dRGec5rzNS49XsZ343JXE4MoivRULUXlXgVKK0RQwg1OOLk3cpq1paS90haen7nRAKRaZc2Z6t1N
iibayS+z0c/v8eo5NU4tw7Q76e3S5HMUKpFaeQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6144)
`protect data_block
HH6CheAkeDvgpjOcXwi3ClQjeK/uRgfZqqSRMBaacOA6odgxPnHe966k+FlANF1Oplo23A+O5uKS
QkqPyFXCkp8qAOn6S8GziFZ/pyPMrD9K5ZjSIgbaeU4wmTqjxOjkMYN5NUZcJe0wAfLjy+EOyubH
KOyHKSPudeUUfVNXrlXSqbsHmxMaW1HQsWHzBQVj4XVrTD/YLe+8L1v9UrzmUpD7D2oPOh4lbcQ4
YFl5oqRPvrpoSkj/1aoYIZGKiuqHfZxSOc7dRrEkwtK4f0LQxmNkRX3tmjt79k8iIWCxr/6xbcp3
LoMlENBQ/oWM4b0wffHZ76L/JojskrW6q+Ab2gjbRXvBKYb74+Rpi6CYzI+FujSqNXpRlpKzoQaJ
jCdYPrjynlQX7QP5TTgbWEWVgKYHTtqF0J5HT9VCqSzHdNdrIArGDGSUeuyh0tnNgd7CfgDjWssv
rt39JMNtokEf0rDhFqJ69v3e3w28kSs/MrKad4nV4qrCylHoNv/dhbrZHaqwl5B23/ZqNKkk8F5P
t5g8M/bgjwllncMgdyUR9LpIrpbox1Jd28RvHzOKFgRO2SFzfsRQSsLdHDMa/xc031z3Eh8IF9Bz
CmCvGxaf5QGHZnIXBatSMPI348nzO5xjmqQEYqhYuv8W9Qaw4ywZK/TwBkxvtdjzKoX1XeVW6kK9
Bh7s410JVEBSnaaCEtuxOywAINd8iiO8uwRorP6+/6FRfc7XNS6QVANicy7GqpqPPeNtRlxkJcIC
i/Yayo+JAWDxzm2D2KWMll0R3SKhIAKe/qEOl7xJCXT0IGc/3ZnZoMm/fj7zkuTEIKH5Z5DLo/GS
BOnuuSqZjnIPCf8EKnL5Sdlpy8tEt2Eo6mACTW/ugqQG6LmRr+uo6u5y72fVQj51nsu1SF3YFfvY
JDWgzCjxZjaXWNjYELSNqjQCjuZUYwgIk1bRzHSxv4WK+NWCJJblTE+OYsOmkauKmVWXcUok8zsn
YrPBfZTs4K8grVI1rO3OCNuFVhlgQMjoXsXxtUHlhBOelS31GxMn0JQuI56o7v4v9YHMwU8rq65+
63QI5/ga0fvPJ3c0qQ+eQjEriPViGqpZK/otrHdG7Ws2WNWCDfmY1CkqTVGNjtI4l3BCqRwjfQPK
VXboxlda86s9i/6B7p8kQyy/N84QnTqa1EKbCx44qtMfxSwaIzgLM7u69VOe+mzC27hdUTCRXSXC
1QymxlPoBRdvv5OYX+XWaBvDelCXmfvBlviLfUV1zUjGlUsMwbtLMu7QKcYX/Hrzqnz4LxDuOoE8
hvvbsMmyv6b7cfCdnRA2VCq+MILdQWhgACzQ3DoYt02gfZwckc4C4Px0KJENz+oRQmcszBeJgLwP
TQN8a+qUukjGlB6/BCjEerk3ylKmyDxdkG9F2IPRWapvWnYA1UzG7+Evk1fm4itYDkxcnLK1yei7
WlyH8EG4GTJA/4QdEa7qASX7IucspdcIC6Z989kaaKR7PflJ5d/plucQBfEVl7hNnV5MZRBnbh6t
gi71cvmVPc7K7Zy3/odg9wY4qXiIasOyWw6J2/10c4DP+nyE6qXmETOFD8vb1OpKcd1lekklucz5
SfW8NYoitCKv2Ix8aj3K+wXqfW2fvInB7RELXUSXrv3K4rK6sFQ86gY5T8E+KPjimX+2h23pvfgF
4/5OsWV/v4otvXsofB1AqzXjFNkoG35kcXrFk+Gl3sNu/kJYLTe102UU1Lpn5PDq92pXXSG/z8RU
kI7goEgFjGQbXZxy9R1CNduB0oOybesP9mEZNxhljVjiyhxVrR+HZkihx87RkW2qFXrDMTRgAXqB
Ria7HhIxP1LJFDo+lnBJc7HpUuYUDHRhWKO5xsE6bH8Y6q/4JRBH3hhNoj2s7fzSEK9GruSOWZZU
rK67RWTnHUm0tG2KJDi+if8bki/g/XlgiT8E0Dws2R6WJLb779uEtV1dNjk2paAKg2fs4I4TvKR0
Ny0h/WBh5IzodD3Af0gUHXaxjRPgnU9D0aYdj+dNYwcVArDfjI8tWm3Md1bV2C3CIjj7kXFdqgex
3aQFPVCuGz1AcJpuUQc8+FV6+/2jPP/Dhhmug49lFxjH2bKGhd1wKLP2Wdb2UhU5PkoKoA8yvPXM
Ut0kw2OPfVGadloODCigxBawQUHDhr/a/9yhGf/ojFZc0SiKAHAEC1P0chxS8r+HxC+15fPUGZ/m
YfsGObfxQQMpjqJmjCGhIG16jrF9rGYDzr2YKLXEHsCWSBtUaZyh4geHNRydT5rs/W1WeZCIxXKG
hQPyxxaXK7tCXgDiXCrg5JI0Tj//jCl9IgZwADYSWl7BRkkRQAbzj7yNQZGB1aIfVoWATGztDU+G
nKG1T6d1L6SnUaXY7/YRxqZVuPVNLRWEu3hSdhYkEFGAsOSTAc84ipPVg5kiIY3PAtvYWoa79BzF
yYZt95VCjTlZzn3kun70V0FrHkcbI3C+wZvjswJELBuzpZFgayuWyipuhZXifi9fRBN4Q6fsJM+4
78Hs1HqSNnd1PaxL7IfkTS7h4psKWbPuSVoe8FjwtabRfFMVsYXOF20a+QXrJbcTwNqKAV5bw5RK
Li23sAhc+eHDobWIjhUjrUKmCz1I/L4Sxt3Nt/SZFsIDisQ2f9o2k8YZvyeG5zlzD2xiOJ6mIxGj
Nz0EUNcNXclYnDeKZxZPvmtmPCYWJJqWaxlidtskTER7znXb6ArAhIp6QmTlc+qhTU+VUb+/mBF+
0MpZAtBTfoBBsHKsgvYVOYB3dEYGShuuEgMsmoxTxlYoFeTP3zwy0muhhIBBU6KfK1kFSXYODwZm
jtTGvW8+CwWwwZ2IOJJFUHRYkuRCHxg5IWC6QMT8529AEwxWoI8HM2mVbuPDEt6pZIftABx9z0XC
O5hLaTmrHGw3EdDJYMUk7fwJF1lJFe4pra0mEPyFEy3UrvJo9h0Iqz7f+/7f/ZzdY0O/Hs11Mv/J
3gxS3o1WugmZTGdPAJ75/9ys8rm9dpYZcTiBY23Hr/+Y8RHHCG8z1gFESTo5gMEeC2xFCnImjTB5
0Irw9U/VKdSSleT6rGcoOO79Hwyha4YupRHVKaYx7aSQtDxflzlqWFVzDuITLkl8c2W2d0kcGAeC
W7qC6U5k1J4EQy5Ta4NlPjMTrsWu5pAZevJ75+I6QNwKYzMlqKtA7A3B4N0nJV9qBIeUHTuZ7K+x
1uCXfH4D7VaaTIdZLsM3dlkVSMDGnEPLj0PZEs98BXbYgy9D16M6xP/tTM86v8/Wx7a6YJmP+U3S
EvP0xKEz8ZYg0ezEJEdFPqoB4Zko+1iD+5yB7/Srg0y5edGIfL4tSVddXxIR7u6z8ZBqBeT/cYMg
mJe44utrQ8EbcHtt8n0fiM697QQBs0Rcz2oJZTv0iPkARiZMLXx6Iwmlbytfs5ys5x93hQnZM8EC
c0E0FQpW67f4HB/viGA77p1V5rhxqGRsu9fGnWcpxK1MxgeVnsWKCjSDMomIGjxBQ/qdZnENCBlU
IU25WA3ZS3nXeU0HhPGRaWJpwuSW6pZdJa+xx/+JkpRCihJ3Bl0B+mCAnf/bcB13Nkv4jVcIHf5J
DAgKGb+sWTLLiQdSHAWJ/7h2OJDRwbBiUcqSiCV0Xm9qbV9FcFZp1N1ddV70F0uXoEU3rYqMV5DF
FjTkwYiK4UvU4K6a7kzqYCa+q00RS5/On8ZApPdeWTLcxG/2dymmB3xzFQRnRNMD1nZT7h4F24ZC
aCzvUN4qPDpydBnfWHKTTUhfcS0kCasKwbeDon4s7AXhxbjnEuROHtoLpZN49kotdxhA3nm8htST
P6B22S9HTaaszhKEncEP44R4iUrOxW2HjqOMdKH5jysZ0x5CeJBwDj5mmhlKJ7JXOBSVqjRFM8PJ
hnMTSRSKBrHs0bkhal+T407nmoSK9+w8cXIDtXVB8pTGlXEOQGcgLtbX1gXZ9Q9n/tfyL48CIpce
mlmsqM1+/zCVXTscy8aWwpuDODHtWtDbm6PmKLpd050aJ1mSLCIKYhkWAuBJMmydMDBnbM+REBcL
8j79D28F2McpprW9Hxt/QefbJit0hNGwCUTdq9uqbR29H+OjEje6db25AiZEXXrmIffFwAySXIJO
Nwp8a/ygW20NYIy3OaJze243m9Nq8lY0jReRdkpzGyoQLVsrmo5yvs0OPPe9/4AswaK4t6lmNjPh
drzUufuzMmsOyng0IB0bPKmbq/a2s4ujP8BuFpjKMnUdrGTntT6AWj/HOlQZsMhM1Xa/HANzGDzu
U6ryrTwnikLOT5sQo0Yomc0rFMsaqqVveKbBFtl689M4Bd3Fk4lyQHd+2Z9RR9+gXDGSR7Fwl842
3ClSJbdwIW94XdloF1xIYmzkoZaA09JfvKUaw6SpHIsUygZwtYiahI3iirU7QvvLcR5Roxr5ZNl5
WdIro538+TnJqIXuSodKAKPMbkJ3Kkx3uB20TJQLcI+xcfR8jWI81uQl0SRKZYjfD05wBpPMB7s8
JJ14MK/F7IS9scp+Ja2/wwr0G8ElP7n+rpfS2R/GleWh05aQ0bx633IMODrNAJytxGQ1R3x+4s4f
D4ACGn+NN1UgNxaVbdFYqLfllsX8u5HxicNX0OVz0XQXKbjg+pLgKw7kMlEIKIjk/+eS6Q1sAhTL
9jAK4YOuRNKqBnwodxaqrgkBRo3eAWQvjnpAXp0Fy2IXSsqzXewh+S4rnQqeK7o43oq2oj95rEp/
cIZpusra61ad7pzoApVB4X9xGa+/W9TJhQMhd39UuOMl7JXYi3Tcwlv6iqlglNxYt5mMs0O44Zt0
MBHmdQP0jW+164pKJch2Hws2zLLib+L5/Lmbw4Qxm1Zp2TBY13b5Ezaoxfo2yvB/GM9gYl8n/BQD
Ubv4PeYhZRzGa9WFhMGzxPR+OpINGodgwYtT7lakRqKB/CmhfZRHSUv8dWElPggznyFs96ucmnnb
8vfP4O5ETJhG7WUOGwDUbUPbi2BkNYvB+/WpA2PH70rZ43q/Zve+3yXKaLuHJL1DPmeiZvxuSbtn
PXpj8g39DHaMB+m4bnDd1zIi8bqomNu+r9ORP+DbG+W+XU0StUU8inq0oji5u6bEgg7Lr0o3sbTB
XgT8DgbDSO9tWEDjBwNHrPY94QHHFWZSarDA+d43mys2yW9KE47AJMvuJuuV9wcQLLp8aCl+Y4Sg
4BZvcl+X0yRBtXbzDqUTK43c4xqe2AJTRRifnpTEiywSN9kBu+N2yUoYv7vjE62b9Z0nCCeNEe1Q
d2C+oArFeaNQ5PxoDMUa3mIq7CkmC9nvyPlkjakmypFtLo5AbAfCC7mcqVYPBKulFTt7VQgxavDn
LM3GuwLa6BqTqmBGqSSSWXQO1n3LppHjCg5F5t2okl1px9oQI67bVbvP01SxG/NH4Vtw6TV8y42j
BneqESxDRFAJPCr6HvGeGtz9GXXG1xhgkin45nBWC3mPMHu7fmLWjuQmUmLoi2TasR6YyrVfXVZC
6lVjviZS26OPWLLjt28D+IX8f6veHq9WRClprnZWLlUp6jic5Mn6YrgUAIG3SznqHoA5D8+JVQ3m
Y7Rmk1nwEDLJgs17NMiggFScom33Ydd1MQoFvPN/yG32uyTcGZ0x1vJhxGoln33Qt5/uP/wDVyR1
4z4JOAEkA5WXXI0OTYlaqb3KbpYXNB4CGrigk0lVclP58E2Lng5LhWwybNyPgZ5BY+8jwGm+oli9
NCwLmSoLGiduUXZMb5uOvS+JyCVYJXWEXqw1AmuvJf/fzfy943Iq7IZ+it27CUbns/Cqeu8VCD+f
cEW45W06HCez4jYIvHdOPUFRrtTl0Vu/cdB9rJ0u7/Z25449aDxAkib6mNnkHqx0ul18VUG72XmR
3tZpxnCo6OGEl51riLanTncFYnymVPQ5ZUFeR8ddyF3lH//cHevrg8aKTRkVmXMTQYFpCft+zCf6
/01QJh7rrr0P97llmIdDw/PK//KTJG6uiQQJwevJIttUJMyazfXOtHzJM6yDS1cLkrW6cEYA2Lrj
P5eJJB0b3hZ0jkj1/khm3IaETciVgveCBPC4rPlWbzgNALMF/mUmTbJqLwG1mS9hg/LkrLzPFGgI
La2ZMt8lpMxTkyohcx2OBYDMK0yNVXE2sqBrPB1xkrcxSBm2OM3SfgoUa+sO+13NVSAdaGDXWEdw
SurJx1cqedMu3R2ILaaQpyUKMhVmHXfyEQLcOfnDQJfSjC4MYJBMEHiWQZWpIWSnl6EthKz4peXS
xd0Js7/xrY8OF5HZ2ZI0YL7Ac4EuOX/N5EQlse19Dzt5AwX1N21TSn6n+624Xe9qfS/BZr5789bO
RmGUx0AtjR7s9vHjQX1maIE3pxEh02riE/xrjoQBMDniZnfnjG8q6ZTKPxHWnSklzB6l56Xe3dFR
OY069nuXykXZXL1iDeSUhBDqOBB1mcoMWfRaQiYtmcrqQ/GCdPyeB+Ojm2s4KNrfyQdg0proyYa/
KJA+oOnxo9pJZlFQzqdcaNJ61YERcY/TSyYz7SXJMq+yRBROiIfyUk2/iBm3bw8pzusM/4HlppzW
iGBIv6cKbQCiX5XEFRNGmUbBtWZfOavXFBLZfPaAymiw2fmLeyP3DQStYskEw5iYpxQgePC2A9H9
o1frduVNgocKBDBj2yqMStKn5FvDbDIMLiY+zyenoCnwCxcO3eAuW4qvkBzwGTSnIWxqktZbVQP2
gU+GAq6Tf/+1QVP3w/FHXf783Pm+GNIGWlfWG7/4kQfbu5qpoB4+sRMfUXUE72z0qlMpaZov99ay
bpZyF44F3l3Ajgs1Ihh+JkLFWxd1d3en4DNJ+TjKym1UIQProhooMuLkY2QcrI9SVj+lLpYuSRnq
+OHDB98uj9lvUCebyvGJS8E0APM0dpeR9Wkn9G8ZsH14oyzaFjkjo1uE/M9WeaSCVSeZ+unzdRrb
o9tYcFvFV1aGZmgPeui2oogpxs5aO4Ng8n6qGkfAJyBPZKEHISIkMabl1DrdBFNMhB3HPSKieNzL
TE3zCDar8c6FxoyaA90XzvpF8ZZNb3sbaxxHkAWNGGY3PTlvva3Z6PPjUozrnXqk4TdPWeI2XTn+
XmWpx6cdU4xRrW1uvJET0weUAZoI80FxdMbBMsM7WxG63S7QPIgUUc69YtWMDVCj9NN9L+Y4B/Q8
U2yFur5gozo7Qrm/rkzV2jrLs1bp5AJ1Ujav3a9xBrwd3v9mEW9CxFo5krCzUppK9MFS+fiNlp/7
eCoenpYcQBkwGHYG5HbJjKcdZF/Rshdr2YYIEPwhcgQrfBGS2avs8gsnLGtbTb48ikUDAiW+zzUN
ss4dsDdHzJrdPsiFKo8DVv2ycU3fmsmh0klLh+kIrT4X7IwjhV6k9X7qbbGNJ428lvDlst6zD1Nq
COmxFidVlwkWUdwASDi5AxIBO3VDhYHSo0M5MVTLPBMWQWi8WzqA9E9LzJgn8C0JdkbjfFioQeCh
NHTdABZyIFSWalX57M2mciWmrlf6XNZ5o1OkGE2iR9NoNaCoHxUtBETvzIhSSo+8bNF0d6XsURq1
/zrtPVrQhBVfzLfscrXJRlRY2YxDHoM1CSZ6dIcQ9Dl6r+3rlVqPFEmB6Iq2i4yzJaVoDOGDQ2n4
Za02rLkXHOwmpeBdYbMUlgjv7nlSVYz5FsaMOdincSQR8sX5Q+I4T1FeOTgELHEbwwZZV/1e+vLB
D6QFvJgDdT82F1CKRoTqCiCKYh5axoJjl8N3XfXxJVFqajCa6MphvoYw32GDzb6XeyeWiv2p14Cr
/WrEZ+F+a+CiPIIWlqiBfUJG4YQTJg76nCy429baQIw7fBhfSQmcLg8yg+T7FS7V5G1vS+wjMeYG
jKB5YhE5NlVXrzv7yQhi9SBYL94l9MJXtAKiBFBFZWMd97gg2X1dRFVfnYVr04p1oEIO523FA9Mi
C5KC54CSrJ+TPgd6QzivixiFO6kafIbWITT8VeNG/GCkXb5XrxVLGYhKqwIVKM9Um2m9WO3ZTslL
chFqfw+Ul9WefPRIChP0mEPHbrWXqf9R5dxLO7jOom3clNv2l4EibOZACI0OXTmRkT9koMpHYtRB
pCfDX49OJKpUU/Cp+sJYsmLd+kJn1ggridieHrZ+C1R7CK4taHOfBJIRgsCwTZBY/Mo3sJ0BY70g
IjXbEUTvjp/TJQr+xFnxiai3ELZ+QQesOPXjhCo9Rosoh5Y3qxek86TLiGdw
`protect end_protected

