

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iH5HG83MPspIMrfUarM3F07PcYUXAKsMpSoZWHor8IVHJa0w6yRGjMV2Oo35erF0AmOS2ghNUHil
HSqiFJ6QzQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SHtoTvbD8Rr6AkY+SuHBDUufituFfaUW4WapyxH4Da1ZzfrZpZyRAwcIAfCxLjL4ek5kgCHG9Ds8
7hM1binFD9EZlI2Fg8k7aEoy2bHS2816iLtNIjirfZxjfXgEsuElVQvPWXeWnlAOMuhxMSWnMyYd
N9q4mBvOGTJvgvxQdLY=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c1ftUxIx0mbVALHhHbTdwFeSnBbihw3DpK04nuOzYbcsAfDUjxfb2+E/O/2gV8bnGiPIW3mcT8d/
V3kyx9qURbiXiSRKXFiDJuGowNo+y0gNTh42bV/j8/c7t9OHJhrWhvBezD7IoTPU4fW70WC120OM
ZDGuPlehijKIPsl8Ct5zwg7gq37PgBo9QqrGUtZlrQG8uCOfYZuOoVzbojKLqf3kRxbk8tbj8CWr
95kdxHrvQ2Ml4y75zcgce6ocRm/QFWT8xGz7TcuYZiDczD3mRRoLgvmUYnFbd5JBkSxQ4YNy9Mea
mQGvgoslhjpKD095q7pfcHjJUfLZzF7q28Ae/w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
0mHr8sw4iGuOu9vFtNEAckvbxTPHT0+dBl9QbXywMNbiASfgyFj2GZYkHkkqLJrcCqa24pDH/uDL
OQknymYM6Z0VZlJoVdKHwvQjfop6KikITxHoxycj3kQVI0ztNKNK10fTthaGJf/71CA2OxyvBeEY
7GVA7XeEpUeYUDd5Ehs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hEfvvlIb1rS1hdfMSQ+Bz5Ud4uvVfrjo5HlcwJfSqFWMcsqyQa+aGBT1QDWfR2gtZOmtfMZzDbDD
fJBdtmDbaGzUb0zG0B/0BZqbcxFZMhnHKXBviyutkpEISPDNEvaYQWHtMRFjYlNJLQOHXnnsWUSO
6xETrwrpNrIIPJzitaqVtSRDe7gPWOKgTdlyPxdzoaqUJe0lXJLNb+7eagsxEaSlOvDZHpbMzsXd
ucQPzYY3a5coux2DjRTxkByqOKQSEVKz2xtIgjp1tOb8mjNyUyvgFHzVIABrnb3LxTAJbNuX82PF
EikZOCqlEC3xL2Krki8wGA7T4JruCEEnAj7H8A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6224)
`protect data_block
GiYXjMKfSjINOmyRookcRfoyVV0QSrnBHxtLCYofj4kJ/9fnSja20WqGhuzcQokmj908K9yGiZMV
cgyOSQAMQFWDkb8j9lYdcQUpgfNVI/on0zDfmkKAvWZmOpcO6lZWtJepR4N+jY7Ttg+3ABoPFLta
qEC4OUsWJdpjfWtS6L/K8GcxvTsShomP8xJ8T59K2Pxcvemf6SGcJkniEOW/OjsZwOPchyew7XjZ
O9yYiy5CqKSX+s3igjhP8tSFL/exF/6TcHEvrUKG7RpYeRLM+NkctTA4fy7x8nmWl/E3mH3r+Njk
4dAyPyDgivORELrH1ghw5wMI50OVQISBgTQ8oKUsNNY8lvxYgphtUuMtvQ/zBJ/dbEBb6+LqgbFy
d6QhUy2RHUenEC2qNM6DWfmCIUOBIA9hoPMo2m8rww5lObM8QfB6hmlaMxVzV/PFmmNZHvGzAVS+
Lf8pVq3gLjsjGJ8YRw7jiwOKC2ZQaY924GS4hlcqpK/9KhSAkBqo6EEjREQqMVd4VW3BElfxNlNJ
YQpjOV1IFZZMqiSw7RcHxgM56CAT0BUlhlZo7wKupRZ/MxIL/o/wdksTfiZW5DF9tt9onUfJ79xY
6khWbSDgYGUK1AEz7fxbGk9kUtW+10r6/fYT3PEQl886v3RuR9vtS1r9zFvykgNw7cmvxN+bEKk8
YjJQUVoWx7evZgZP1FSTLkaShtsMu6OMi0/aN6+BFZTcrDiCv6FbPViKEQovJf/K/GwXEARP65Vi
2FYynMWc4CBE6x1rRV+tiUMC4+bv249sAQyCa9RHIOks1rCutIdPzoe3YiC7vd4Qh1isbcjOekhW
Jy0evnrYU82eNp2FkMttHcb7i/GSruMtkflRfzqLZ0xiHGLzLbL0z9XegwHwKJGPu2R6bK3SYOjt
GrSH9/Vamm60dZUssnFjGT2R5ghV6vVa60P+U6gsf29GB8CRbLa3fUIQ+5bJQxybQxw391RfgYPE
5BG3izUdvPotXE8TUL5O3grqdvQj8XJM1baTV84kwk3OAmUYwoOJ1+SXgCgcnVm8/r8maTOpQNcQ
NDA/SMPaxNwNlN00yLMKbcoscKcryWLa9onGihUMcUZRKS2yfSNqushN+ooeSLSs3r9RAFYDiSA/
g5U+7ufvARzS0LXxHBqi0amliwiebEtbZWLqUbY7gYI4/SIHlqoILZnJcNWgW8LN7oZd04V0PDMF
et1MKNFx6du5Q7dBf4rkcsrTE/YtanLu9fb+fLbuw5/i6echbHys3NUIDttqdc25Z30/Rgis4ZzL
sp2/1GKBumrSlS0nsEDZkqcU+PP5hiQFTALSBgFQDJqvIFfugF+eqDNlPc/1RC8Dhcggchgfb+kn
uQ3efP84nfPepi5Ldpl9DzJ5A5AKPjVAE3kxNSoI4yzN4ofGWRZH3KXgbKrDUjzfk+0zvaKNYdnO
+2tPNNkHIVM9LdkJig0cy7ZfhXv+yP0fBq0SeD0VIaSXdfkb6K13fU6NrU8UMcktN+IPkK70cXAE
/2DBbqXjPpUMGFiPchbVM0X7cnQkEIYiJS0EdKspo1OYhhGXj1mdfyjL3i0785/3JKcQCOgnt1C8
TxO60LwW0G4cW0PJ8vfTagsMMfADXqSmCV94tpRI1mDgSmEbDauZd3nQwbfrbAlqdLne97raaVd0
eZBtRzOb4UhNJQC5YN1Y3arvXNGanmciUxPECts7pDPFCFcp6Hj40IkK83aD2gmHJiNzHBt1PpCe
rG+0Zcix6V4RMOHezR1+BuaI2WKthTpvr18C6yyNekwkLDNBzv0j8fNOjBAkTtb27OXBrCtPitTv
01VH6tM6H2t3M0hNSxDyk8DD30x7RidyVwFCirVm1CqWpy6sWmWNvqSF3UZYalo5CBCQP89UnyMR
wVRqI4g9bkpwGpEJ9ezTJgo2zIZXFB1+84Fj6JixRa3CDvH0hY0XI8gNZVK600IcH28rgpNL61dl
yAxQEA4R20hvEKSpTZOCHhOxfUCiGwicVRnmrcBFn+TPQD8zQGusn8sHYc8omRaGziP7vtRmkR94
9td3NLham63r0VCRu7YLWfPftp4XmG70wqnEURD74F0K9xs5lHF88J/AR6QwOiHRcMX6Bsw/HXwj
6xtmwLCyhbgCrV8qcTAs9KRGutSMhw2yseAh9kYk99696ZCbiQcltUnXOJ3PGPQFiPwi6PzxlVza
P4m17jJcfC0myT6sTxWkuvpfkLgJPZrlbnWCdYwat/x/SOMMw1cKH0kdrAg/mFKcQOWzVlMGY6uO
Y0eOlETQDPPOcsYA+50ppMQ7xXUDiIXX1pHdp7WOcjIP+dC0twBrCGBcA53MmhGbREmRMj9FOecD
h+OYDxxDBbIxj8MyIeW/qpGQdVW7cEtfNvAQQAZ+oo6Z5EbXi5YUsrohcEJ3h5uNenHU57ijjL3e
PcmUXBsHS9VHO54baHHTr3VKwjvQPYs4LlUOF63NMkfKadnSbQ1xGlcqAgEfu411hZOrxo+0YF7d
daTa4f6tNz8g7LScr+fGgDHpxUXU+I29JwWbxNcrpA15QefRWInrdDIHz631ikKgrvsg26VGl2Bq
CvYExUGuEr+Xnzrk9mUnPC2IlZSDBWHqk1V6PzOYj5Jhk7q5NXyfbXSFzjqlN0mrU927WiCUgpTD
jooFlxwH2q4jEkUloSQyxFcjxQHWUnihQhKauw2qOG45jN4NOOO8JqP/Z0eNzAXNQK/WgM5DfooG
AXs2QbNhIhStfd1jVGgu6XFHJGEjKYNp1rwho60Em8YQ/LLDHy9s1FAdGep/7X6WUVX7KzdiM/+z
WT3D11xge9GBdsw/U/YeMfUK4rqtAwTemP80x24PxESE1uqgJTcMvgimdFB3O8Nm6upeg/MSoZG7
8cmpceTsdnrMljnzqlrSzARtezBy7rWzRSYM8DYGz77tYbOHPrOAx0MaOqxl9RrBQTkDWJru/Nwq
XPVSzPKa1lJL9cuRbYGoZdGVNdkAf0FG7ztR+mL271JVqwVYc8+ZWb42kZ8xXZLXfhKqbLqkh7R/
P3f84BmcwV+rztPwQ7qdM2mfzgnSsKNi//KcWHpWxf+zqb3E44R9Qaw2pkWh74xuWnYvKVN08D7n
zxy5msgRghrstXMtu2jSvrep6yctHJAWRrWSGcSOhkHBY3VmcEf12ikW2+FrbYAe6yzhHcJfjeYx
hh32EOl7RqodBgOFw09GCzHmZmoH/DD49p0OyCw7zVhnL64Q+AqB1QHW+CMK8B/iVBtHH2JY9QRY
3aLH6cjjVnVdB4GLLVyFehE/vGZW4U6INcNvumh3HduyaZ9k9+DtfnCq5cgPBCLdGqJj32AsD1dG
Q1tr318HM5ViZFYp2rl2GOwAS9C5BPg+eNnTQ7u4nMDYT3BXEyhQ9U0R1Ue+WYKWMVEMU8oceDOS
Q3zdhJnYItAXQsmtHLk5wtNwxNgL6TmVIQJGC/Sh6nTJx3t7VnEyHNQf3KUFWhwEnwMT9en1ilFP
/0qaxAIOBhBEa6vd/C3gFO5T5tzkaR1xo4KcoPLwBktvmMOHtQ52pBwtcNh+iQIUOAAg6xbU8FTb
2o+66BgGupOVXMTCHo6qYLYELzPOAxinE6aWMb7oqU+gfNuOxeVAGh2fkkFDSWGSoaln5qjHOF2k
fCARRufTZpJM56s7liCsy1n/WUNt7KciWDkeTKUYV5FryUFXXT4eJFxEypANw4FPRCtjODa/DDL5
kmWlmEvmYvcTZbzt1auFwq7smVrbBs2qdNadpGqSitxFypXbnE+hLVzhydll+/vfKzJDiq547cwX
3L6ioYNWgnRUmN5OciBLHqvbL+rd+fY5lsboIWFKeHktSzKp8BgMvk5vgcLfHjUBTJoHKN8K7vlo
l3XIlqLgasmmWHXm0sPvVPzfEPIN5uW7v5NtDgerAfV8wPDdvYcLPJ12NYUvPDnk+gOg1AmBJG9u
AXL4WTFGlLl6XRaqz4hyOBr7BIx4F4i/Fhp4RhtgkMGdcDf7vAQVoCFkR5wRyI8yIzn2qlZfP8Mn
x0gHGjOI3hn1pNCAxbYh+6ERaJE9c67NQEQQdZFrtO1tX38FNUDOfrhlfF7PPPSS/x4JICPCuRMy
Qt6FaPBnz2a12i0i+rlQUgj9kshNwNvsenB9Xa+tKLOvlkzRarXHG/I+hPurPl50HXVIJMLdfBHn
AUkrtBc0YnGfsnTAxB/zRT2Sim95K5GWN9C3o47227dOfsXycJuOhatfzTLQONggiA0wAwXgQ+vI
uS107JyGKD5qSAemZt0zhCeWjnumczytLtSfK5bKIRMW5uhBn1DEP4xB00dJ3I4CrPWaH4TZcFqO
I7QU1h5pxkPAd1ZNUsIaxAeAniBvToPt1Z0x+pumc0XN8lvUmMGiW1dHsURcdcGhrrQjA1u3SHmw
TGiPZO5nJz4f9BhK9nFBWLPQ5tvM9o10NixtSWauu5S95V0D28n0bkDOA8XzZL2AUiVuDXts+lGr
aBgYNFUSRWZl6NtulHDQIDtCK35G/ip7VE7r9F0YUzxBB0IJsq6stwmmCZOowAeGK3EZ7vtHnruI
WBQ7LsqlfkA71PLgjFSw3HrUFzNWMHHYbVwp7JGdE1VPyyDYI6SvqaWYyxwVbdKN9Kq9TwFp+k6o
IEltV777RTTWdpz8F2gtsGw82vyayzqjKG7lO3ie84eBzuh0KQrc9JWQzzFh0o/KLNbTRQT9uKBS
rTgxx4Z8dox3l5aS0rSz+ptFsf8PlJKq+A0eE1XnbSnKSj+bm0e/k5Jl4Qm38lgLt4JH6grDucBv
NnL5nKzO0Q9GThwm5SULGR6bAKu4PEz49EkEC+TO1VvyQtLHEtEiCSUeW0GJzh3dxZgEFYvuPhu4
R0samI4xC3W0P5OTlDNqVybxl7K7w2Ux3/10HypnaM67iyuj+gCDCsbXmGcMljMVSHQMQ9yHQkfY
0xj6tc8MV1AxNWekRkmGoJ29qm7tC6HxDNbkujw2lK6ohuGHisR9c29im/SYy308Cv1Om9ysStLZ
42VHGZtue9BRQJAFC3GcyfgtAx3+EBGFBVjlOfow/EbHl+yMhAQ2wXYYEsZgHi7wFxWR7sPXiLkW
0KJfeqKB1gZX1mT+Wde11hzxd8dx6eQ6Luy0Voo1DBfObKeu7Q9DTarmcpAGO9VQNQgT2xC5svE9
iCHIOQ3QkPPod5cqwcuMnh1TQThUoLis/DnH7OdWzDw5y+ntYkrlgbponzeBq0vHmt6VPt/jTKAc
zS7gsEgxpoLVY0biei/TijqXgUDhr0XC8Ba+dJ7c5S4AaKTmtb1xi9DO1MaE8lVF5U6kXJNbHR0D
UHeL8EpihJJiAoMdzzkelpMgrLv/2CfS3I8qpuk0qDT33Ul0k4DYZQEDQptAnS2lqYQ4L4oiX5mp
9N0B4s6bEqytH2NzydjQduUob1xZ/NO6bkSFCp5tlcwsyh3qPVzlkRc6g2JsIgZ3QcjaGwCYEpIc
kUIVVNPllxaNN/hCBbjR0GQSblsx0FWfycR8tuxdymu4q3O4Btri4k62hHXqTlwjKaND5qA1zWKO
QkHcCdc7w4vyVifY+x2noR8Yb49/bRHteN7BwRqFSkCMhuskQ6M1pzWYeOZfE/Eaw11k7C3m1iAw
SYVdYEBe4L6DQdNk3IEw+Bh5yuHjwd76FTCRGUqNsc0iAmX/kWvV3HoJHW09zGK7ACTA+Wt9QQBN
lsJhny01yJVZC9zqfCUn0z+Mp36Ym8i3qSBMfB8VklpwFGCKRgdiv6OiARkjNHYtvn+mj2ctlLks
uFhHEd7i9niCJmUuor81XwJL4CDJVt0Yt0KNyrvb3SCHe16P4GLTfC4zEdVOr2PIwYAdciT67p5k
cYJ25IHjWh60jOPF0RaESw1+/a4AYQJ3mgFfjOdJicmdHkfjgWjVxr5Any5+fL8HIPq6oz0boj7G
4rDTys/Thhi3YdRki6nw33LZzrWcgSLVy9vl1VoQk21ZRzv7P12aLqhQ3HOHoeRb6U4MRwRHBmmJ
PTM4Cuc/jSzKX7ZTKPOEF+lmCwEjZAlmMzvP0ilNXEXqCyqtleghevFQP6wIBNxBEZAsm5eiU88I
mjN5phAat3xtAfKxgWt7SFj1iBjLYyaVVlQCEeerKOHtOIPzTRRF4eDnucmYPm9cm2F056TkT+Cf
F9XibN+jMd7TZUCgdXgGED5mcbSSAXyj+RqnoaktuCf46KXpPR06TbL8cIGApQ4opzUrLmognTyh
Gr61HjatR000WpkUeabnURdIlMEsEobLkHqRxkMPzRh2Z9IjIZqv2a0N3n2oy4QPdklFEkVLnj4Z
FUl9+oDCaYJluRKb6LrZq3HiDE/cA0KxeArLEOqSAVQ+m526+Ba6Uh9sx+LiGG6CaiQae0U8hf12
XaoZJcU6bPt7C1ZjAefOqnYSi9BGDUkeOdxea06FAxlmPIZPpzbzQPoR/iHBCTBXUFF7j4hMtRvg
+sW/PBYbqwxV0/EhFk+qqzSYPjC61WsdTiDio76Y4ZsIXr5JZxL5hPeXRC9ccBL6NEfFI/r7zolh
74qukU5h42zJiUSvE/LmSksWpxwAfgK7J6QxQvf7mxXLTgoQodkgjHArU3DFe1oBPjnAbAJJnQKe
+Siisyjfo6SSFGyVOp89TU1vxZNqGvdNkold7j1su53Uum8MyKSg5wiy12yRoV2HjSn9MAvnRi+5
umH79NB7sFn7J1ORsdiE61Q7dLetHPeZVbPZL0reRs/A4p0YKwT6EAtpAtmZUgGHaGSmQUiPuyuI
0cIDl2t7ZnqO6VMmdn9HwOC6C5kquG+Lulx0aMi7gayVnMn8rBwr7jMYbWnZKjaOv7ySW9IfjCLA
nknEtRftZCCHu4aCDrjmWKMhDYMaXlHkofmLPo6UEZHPSVvKCezHyhfz506hXJ8dTetzJeonCA2L
3tH0AxLadNsbUwlR+6SaZJXZb3GAjmIlwxBpzQjWIZwFKgdbmh0DqtwVL4PbV2cycmQFd23jYK0A
9zkYOExRD9mxkc0gn6FjuF2UA7pjFZCQmj++VnqC16+6O9ek0sILoCg8Soqzfgase5auXXLWi59n
Bug2Hz8wzn45qr7e49926TGvbHHmzlPH1BhImmhg4+BXqmCeeuZAs89/Cdvicy0Wb7fNoaqPewLJ
NAswvBA9/gl+3nvb+Pst4sheYYEnM+46e2HKGz9khpOzwBQdYjl13zZ1BHoKvVzTW896lO9YziuD
Ej8+vjDImTtVTestuiO0umraFZxBH+DAeMTGAmu2qVZq83N/7XT8+eULkiEs2VK6EGj48vKCeyCf
jGj2KIEuE6JSOEwQpl+z8MBK0ZD1uV5dA8hni2cJeU/INjo8yPZTEhDUz/Lsc5VAOGWSCeV7J7Jn
V90wXHxTxYc3NiYHBG36Y22i18jmuPc50Z/MMFxZvTbqpA4RGbHAb3xrvs//86juWvy7koFOUWs5
pQsjhox636sabEbNfd2Q5bSstfiGjBBgXY0SvEFvLhRhmySCNvjilbhCr2GyLWuqeN5bI1VzO7Zr
FKBabuOj6Hn0NaXxbwNl0eybIPaIMHl6XKSdFke+0JHvcM8rPXUPjABCqztfG+d7XeafUCEaXivl
C8GgEo/9hRu+DtuFmNfipT2t3PvDIVaIuAZCDfpuF4Bu+d2ITkk2CFPA9oaXONxUJWwb1K7AYhs6
QPOl+wPm9LfsICEsxjaETyV5TSdqo5DAhYI5VlYzZPiYLfklq/daf+/qDPzXei0NsbuUZXuY6Vdu
OgTgqjnhMkEsEC3DufA7tmU3n9XyH+JfP92WnSKqNac461clUGrbDbKC+EBW8FHUWCeCZuJTnp/L
yv74heXP/SQ1PzLsrjTsShZqCGKlunNAZFyZEjNOem50ZP4BTlHH0BFnJcrGnkD6TRoWi8zBSIHN
aVqdofSaNsRgAs6X+8frrn5BeqtMoRV30cKQOPcVL4dN+SgM7qyaPAiDYI3wLRcxEuog6WpVxRLV
b9dlptTD2zvg4nYGjC9PfWvUQoeQ1UBMkj0lR4O9FOlShYRKgbhmWoHBMb+w90/x54IiPilW2P2O
5PZFcEtkJZydOrAbhPhcXgKIsPNDxhWKdeYF3U/Gi+DfKVs2tsSoFJny7dIUG50LlEmTzQlOfXgk
Lnbl+jzhM0xzdGmS2zjvdVptjlXjugRJIxXq0B0+T7u4JlBYbvqtDc/RjOPvdTtUmk/DUkqNVoJ7
AYUsVK2eEFMMObvBsZHysqCF+oWF1r6eGghsvE9g9smwmrwKs7WNiMEgHXNmc2xGH70pS1MAUdWW
GI9W0n+wQInvT18=
`protect end_protected

