

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lEHOI1pWkEYCNgH1zKudlBPIBffO5qXEABnZhCMvMp/N6o2CZJZgnDgsgQWia+9OI2uUO2BGwNCP
CRrpixVTHw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IOLqqZHFVZBENbzvNW7k0Z+m9/COoXnW/wg9J+Xfsu8THYyQglMEpOq/sR2Q0Z9JW/WLZ10nARFo
oyykiJZ57oUF/WAa2Q4YLbK1a8RNXfkYvbVuoe+Zcj5TkD52vzeDe+WHRKoIDxlYux4oixsLvJ+b
zajIEu7tSuP6AyV4ofw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VmUyzXwDfRPv7i1nLcfQ0w7vfltu+dsArRfszkUZ23l3rWABIxgR+nZwJhVXXAEBTkwnBEcW5a2q
bHtanBWxCPVCjFkBYghRT/MFAvCHkss9PMfSOHFgWJ2lFFPN4na/pslXAg6wFnUp+9HR4OkYM9T9
s5F0Jv/WO6kRhhwx9bG8JWsGsvQFfffrXGQakBqm/L7ULb+Cdl5Yoo02d+984ISI3kqTLgbLwesx
8ZR7p1Maay+8T9JA+PVBV+z5G6luEKiuqWgTRYPU1eYCRXr6hr+DHROX6/3981m1o7vWBYEejtc5
KqHPUynqTrVYrtSb4+Nj8AhLqJBKQaHHxdgUbg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yUPHiVOEEjydr2X9OsWiPuJh3k9pHY4gmpZE2C+NpmSqYzRqo+gBr5RpkbcehcNZxH3/GnaVvUfa
oUIfTYnKL8EoO3FIQQPxxJPtJew0QYOmWJHQG32xKti4KkQ0RmGK+46xV+mUqC5qOONxkeurqqfh
zvgr23bUJO5WAkPvbng=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
azZ7mr9aZkVJjumDnv/aCErn+nV1rO3ffumyZKKPGC1qZfaUlh9Fe3WaTjJk1sB1z8/ffPd+M0OF
eoHBym1JP1nSGSiS/YWBHRJ/CYmN5GJXt5y/8LWoG8LS//UEDIqV6XuH1ZQ1lsUBRO2PpX7bha30
JXNVjKMdFbcyLCFxWtYb6SOi2bnF5nyNJ9AB0eymEkgMw1nEnJFhw1H1E+YEu8z6tATOMuvuigtt
RP9OqiyqslRiLQXPGcD2xuIlNWAgUfOlCNfKHqX6cOcg/Gb9Azhm5IZ3RbOrHqKOX2cc+QuFl4nX
vDBf3zaQrfZbx3mDksRFceqQjCeQ/VKWp5MkNg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6224)
`protect data_block
IEzP4bC4th3uGvNMeAkbEi3ouqaVnK05kbbui8UFCWIKyzspuXi44YVDaKSJu+OxBcztnSUeULJj
syzZA1tWXhcdllGN/pt9Va+F3kGdSiAjqBgmQIH/FvN2QwzxNfMo4tlOECqNR7uHfbC67NtnN+ba
Wu4i81pkJaDTCYdxc6YYwb4yy0Iv44Ot5id1tq4rf5bES3GAG472f0g+gCiPSAvA4wGtQ9BCNyM/
6RzKQP3knBL2/Oh8fFmJw6aIpCoXqxOEbqPf6EPLZSiR2l4lmfrKyzRZKEJpKugf8LFnuUPkS9hK
llouhyrMhqw2ZJfGS4x2sCxMV7fW1HkFl6YHpcRmFavkjEvFOvxV3xTNZeOKcifcy/iqQ51U8Lzs
1+SgeoZiSLD0nXGZJ8wV5ORkDJ0UiF0dalkGxqh5aNg0P0eYRfkfwm6U4eQlfJ/kFLOb3G+qeaUh
ot/aaH3AwbkNklZHde84fvZfvomTcFn5vp+1ald5AYEZOo1v3NarwFElhex/sdUjTsUA9RNQqWU+
DVf/qKHWKCnZKIyjnKIsHO/NH0KFWVlb5jhi1faGImphfAjmj2zkYuv0eKsg0hnStdC6Qofp03aj
/IfhtzNF54CmcYB1tXv9+UAXl4hyFBENE1mxOdafYXwXcYNbcNBf15aSpP4fQFsbb7ArXk8x8ZU6
ZNiTFIzoq7S6J+XfZOdvKRXY+LhdmJ8vbU1seIzO9pCWszjnlsXnlV2ZGI2LnzyOM2ETY6OOZLfX
FUDh1+Ntx2Hsy91bbKrPCEOIc4UU+TSriFrrVozZNVN5yWQE6KND3miRNyVoQareBGqOUu06oNU2
ujYkrlL5o90yA2OzIC3S0WJ+UeMTEntO3lr7BwOJ0wxy0DcubytP57aVvA2y1V5G7LmrAyhJWabs
zga5EaHnXwFjXWpL4rBd3AoIat1NoA3rjSHRjODk9tRtWsNtBHngyZ90K+SefbBpNUIxChV+7/Ez
FdXKRBigRrOT/wSDxHN9mrb1bSK7B0ZTJG8mWKu+qpkYsNWL+Bd8gwtOHuSyg0Z48spiRdgMRAQu
kMZTF/x6zqfYiUliIHSZ+8CTN0vSa/gjKnhRbVk5Toyxcdp4DoipuiGUiolzTaJepXCU1Hci1RlF
2LmQtFNL4Lw94/YJ+SHvxckvzaS7jTQ9NoFo8elU9aa5gTAIRNyfCBhQMvRiOJrertCJ7INrJueA
YQXsBAcX428p7p/wPoE48ZF76g2yhHE2SLXi1a46OZbsodQZRO/B2W6vHLOyF+wJpfxj0BVTfDRe
Iy9lljrjAu2TQNZAIxvqEl79PM6Iu7hqX6i2GdqYC78MHggBdMPpJ1Xx+yzEFKUJfKGqRmyqNPtt
3JmajdFqGp7XvRZ4QyeLegBSgAkn+HuHcJfWcO89ar8+K5TP2h60reCSUyzEIB8xmUixKa54p5MB
QocyJ5GnpSsaL6eaUa7ZUfEVFybub1h373aMl+h4xFUIySavc/OZahxe8Mw2AWsYfc5QEyOY2ohD
1GvmV7FLt+wS8wrGcvMsAqbHpoAx1hWkQysdSA/bttmKHyfZRcAoAtITUt/YordztRBt/7ZFKaDD
rr3tAenk7uB1AGrWDxJ5HR3BnebiUe2uyOeCT3DyHIhgF4WLGuWPjgFaYiX5TmLy7uasiOu4PH+i
D5mkJCHBEaCQZUDpQhjjFbxAOHBbpasoMZlRVWeErzb7Q63wfo70v+65FawqYThJZcG4QvXwssMu
PN28ScGgJC3blvWfYSjG1Is/aObQtBnnawl8HJXQ4dWNxcwXBL7YEeP5qLqOlyG0rLwHATultaaZ
VHKq42MesGYzxewjjLyKQOJq3+bDpLt7uBpu3VR6IdasfCePSRuTUxc6B0TYmxQA38x8qW+gw2zH
iqr3erhBYrtOUCzVsGpnqfRgYLFhBV0eGCEKUSmPae3pVdhAAByyVshf+B3q27C4g3YuqetTezjr
lb4M9wpSPBfFx1buAG/TZQ4KGc/CX+vPjI+fn20Ymwd+frFeFbM9DGyMF7asNjq2gL9scWVzzWla
GdTnA4jynmur9FrLNh1lxEDvbWTishaI8in08G1zyrxw0LoSrs59aJX8bniIw/fBXWmaygavkmW3
PiKw4WMGat03Q7KhacqgP5lQjQHpD4/L3R5o6s/kvojakWVJcUREL5aiyqMbWemOYq0w2e7xssm1
rRaopXcoImxNOjpwyFKiDCCWlkXQ8t/Xp9wt09SLaGCzux+qkZe8a7KUuaFJ4lXShti189Ybaa20
9T/gDG5Pb3D8mwjBlDNWX2SEHAvN1tntG/s1EFQhH1MWV0q7IgUfd8FPxko9NbkwFtpvDG56VIQC
oVIddctS9QlsrPrP859Na04tOkLIrUjpCmsSwT56CkJGiqjk2XlLv+K85kXK3daTRjcWkKkyICQ4
CHBzDlIQDNXZODfuGHKZ+fu8twnkRbangAF0Pzig7OXu1Nz6wVLXrNcHzsR+Gt0irJoD+/NjdyCv
BWyPnTDx9MEwIYQhW/1ehDdD0Mgp60vvp6kFLeMLDENvWQ9wxnSvAE4xNA7tA90umFZ2biU1j17O
iW42WTD7hTFYT6XTPr7MEmc7NVB8wtwwRI0NLeOLF7fDZiAqadbz7aRDsqVKJyYqJgRhVD+roOa6
9fD2hNJbgLG3igg1WL0xuaCTctatDjtU7UfVi3SWdoiJ604RnkaWXTTNK3OOcdhXohD5lD01wNb7
utNW4q4jAu1sv32Kglp3ZGIlgPoFS6C0qoitNKs49GkfPBNVc2Xiie+2nMUd0aduDHNntATZWGNc
G+vqdZNtOGZ6RLH+hy1XavQev4kDUMAEQ7SyQNfYQPZbKkMpQznxbrgmAKYzSxY2A/J1Sm2CMjT8
VYLMJUgqpUMxXdnCPR3Yt7nNtgreqtVu/FY7aV1SlDGVTToJkuGeA9h/Wi+jfIjQWWIDlzoOtey0
3g1MDB/vrC8yDXGxDhQWMcXZ5BRKWTlmQ+PXl4dlkA+mXpTGQuDU09wBYoQ6QW8EoxJcoVfpd7Iv
A4Is+0vNKX61iEbeAJDeiQbJXQ2sKZKN6G1Tu8sga/mIPgoQpMqq7ubBiZgxcKEVGJHUFABdDF9l
/To5uN2/QWIQzFhKoLMaSdvKPzU+GxyclNEuRt8RdIaEf8/chxXqgr+s0Ikvii52ARAVFmK98C2q
udjG4TSAHYVRUMQIZRcfdwoR9MPT/KVTnDcHUYfzUDwbcxx4k3RdtFBmvCIgN5ymTwVpphnHPnGl
YrjJlPKZQ6g8eKCP3TGFY9xMZb9Zkjavxl+m6EGCFTWHH9X2y9P8pEhvWbEnqF85vwo4/3V2GGiG
pPiEpU6vJY8a2HryTgZguZTIMACOYZSIyR/fdbkgGx9shKYqEeWixvoCzUOAMXzToWSGuHFNBDAE
nq/zakSNZdmvV2BrcFJPBN/dTydgUdZTMcA17aB6IugxCmiNcupzzkl40f57OJGrXrYFI3wxn+7l
R5224rK4RCZovzDNQ/lt0d203NRq0N6ZekCZ5RJ8bkLaZgKx9rvjTXNWGNHT+u/yODCnqySGs/Xa
o6ZCuDIeCKK542WwBCYeyNZuqNoyzRGUHolrxQI1o84h/lSfcd2QdRT+vJ1n9K1/gQmWL4GApqNo
qBLeWGEvYK8YT/GUDd7rYobwnRd8awTKeEfjbMEEgENfY8/7gAETmSS+ARZsDI0EVUT/OzELT2Lh
QPpjmB0f+ccPJjkpNGyjKYruZHrCp7sE0QjPbMCt7bH8W1wYNCXH2Je83JNlPIe+DncvJlv5otdI
YerM7wRcgXEx7fFhGusFxjsjUxWoGs5tmiWOcFHZNGi4U5h8jVEz7DiQZtrj6fsBgnyxF6M4Yngi
b5iipKs8AwNfQvILkbrzBJdFhamo/m1AhLx6H6cQJbmOCkKxbjld46DC5YqR0T1DkwkrMKMebIj/
OyfEaU91pHNtKBlwkQCI8GIYk241657nvfXSG83Qz3Cv0ZsDmVP83/+DuUXXw/GBmUUYueMD5xna
P2ntqa7xFAZ1FQm7RJSqSWPBlmGViJYy1VL+sXmvAKwE507JKQjPY1Lhp/YZDfvuXSVvwlBjI/jl
vKNHAQHeH4Jw0SO9EICxdnJKD3SqJ233afh3F3eJamcJvCO3E5/FQHwTs3e2fNcWBS1pBPGz846L
9yNes35OyQTc18AoFSC4OwbKcpdSGvz3NxoKakQDVTI4McH1fQtoSkrxG1eFxTEmtVF52+p3eQrQ
VTWr1hchTdfAVXfE8R/QEA7IJOM7DpOF00vGu7xyDI0u5Pqx3aEl7yo/h7S/T31DJOk6nk7auJic
kf8B1TXRJfIteuSBJpcBLwwKDMCJSmhOBEc2vCbEzr4ipF45O6Hq6P/6NjX80vxFRwtid35KJskT
suNPdggAsfghdGDgFdOMjodoWAao8dvbwsPCUUMWSQQ/2rkyomUDeV6cKelozJ8Cc69ubbqBb8Ap
w4469YOIeQXjIQYShDryEzFVaKAi+fIUDtryyhX+Gz+iS/vpxL64Z5yja1w7mmF2VtulW3OhAIcw
rk/PLj+iHio9NzprMcVNmIP3KhN0tITCepEGitPHZZPyVsAq17MF1Gyqpc7fk4MEnIyVerThDpOB
EpAQTA3gcQxkB/zIyZ6SN18Um4AkzLe3VHjSgzjDsy51cEvc7i9T9y9u5Qdgs5zWbRuonkCa/leV
VwYt2jd0+DtFwErzLYY2zwSJuGwVAazne68qpajI33HqeBDtMIEEdY600Kqs6+toXgqo15z3uY5l
/qm5PrDwMaXq3dfr7UDHFIfXX3PcRYAtUgBcTMj8L9SkWLP4b40f7WNIhUJQEN+BPNqq34QYSy2V
9FfOZZN2Xn7NGD8BjTpvKr453MLCXkz2DqN+fsSMUQSHZl7sd1FmyW76OwYOEpr9F6ofYSXRVqQ+
CyKCfQq0niEe5we2je2SdfLF59/C+Jkh+lad0nQ60pnfyNKfu6EM4yFH+3F6ayiYHy2t7vSVaQKU
UHjk+dRe7AUxtYG18oOdtfaiOqBu5m/l79CY8vUM8ef2I58XtMLe5zMmUfsMuNLdVFNP0vnNJC7G
zRUpTm9QnbpyLxovJj+wlKkJ6JEL2R9MpTGpl1atuRjucXOIMvPwhUCXFRh9VYLxy/ArM5Pimln9
RWKByPDb2OnfRNUs/Z86br1dtcYhftumhuwIPBHQtrFGldKs8YUa5ItMf+o3vbCKowQJCsLqM54t
70lV0zN9AYEfiX0Jwt/qxDebY6242OlSFdpm4DtuIU5sAnohxW0BQO2kCqs1aO+qXNZ5IFQNG7Uv
Sg53NpiEXJXxPlzSbn4WwhFMjIMYJx4jAesWP4O6wp6CcW8CTAiC/Kp+Kh5HCN22bYuDcApKWdAg
FxGyfQ/xJllr+SgcQM2VMl/ORiHGTu3It43ExP/DaHlEsyyLRyvjitXdI+kzNkT20fp96SKMR4wX
qDZtpkWDWD4vDEhXpoV7dDyOJtzTwVDZX8Ffiw/+XtV8Cjvl+0vzSrvWJO4DWGa4NmOqicM4NxLz
k7S6PlhP+kQ7Jq6ESM7kv5xHU8lkxnD2I3cgiz50587sWjSQvuFUaXknhe8B3ZCm118lQRQC28oz
8XZDA0lRFfA7MH6dPdbjE1hsBZN37Xzsg4Tyf3hJXtflx8GW2Nnjrj+ZuZZAljhLeNS5H1uY+ZrC
JJKd9qKyhhQqmz60Nk7hS/PkK+Lpvg433GA6hAD8ECW3tCoQvv0IK+AEhWg5Qe+UloynqL+2y232
RTlGOPHJ78NmMuhtyaSUvFKISjAQvTGwjMveNpCbaIlt9HX8QYOG0NSJAf0ZoohsEhrnM7zT9q/c
7Q91uY4DrGs0O4qZ4nuz4NiODxA2JdG5eSnojOSTiOY4u1wUSz55BrljjfpS1dZkDUOMz4IeqDZS
2eKxoG8MLBBdp8G+tOdgJU1St3RtaIYAQI3oq3WEPNaTm+q+AkKS+RO/tKjLYRRo/lwp655vY4oj
CfvQKbzxHuavWbGXyRpmxkW4ddyJeE7mMj4c8E6lSpovqbdaspHOuGeskE11VqGjbdERGWi3u9Wq
Bl/HZZZpp95OCmE+haq+NZ+fT/BbOlel3x4NFgfqN9tt7fjFHE1mT2OSfmkJl0pmUbMSvQpt0Hml
NkXi0IVRzU3+hH5y8K7E1BT1ZlP1siaNQ8hqgcUuOZJ+LkIB0quKCIaxiYiZUaPUEQzcXbZ+DEZR
HZHVnrVqKYURf4uv841OaTEog6A+UrIBqbIfxnSZayPQE8i9YIdKWjIqDBSEDyh6VMvOCKZuBn3t
8M5aYgrYi3m+XbXhV4C6MWSJmjSVId0i3lshI2zCpymk0TxbB9MG+hannSMYWftTyR9bkKOc678z
Si4BlyGr+DUqUBKrdp1a1NEQeV1FWE9+9ZHHX3C6a/Qfnm+RmKmScJTIJiEMEOMEDEuBQr2vr5sO
u4r8o2RjpeooyBpuDEryCGzQV6WyamJZ0oPfrXIQzLWYVFYu5iynmHGXUR2F1Rb1Bqo2gi0IGCSX
L47dhg/FCkLFfISMe91x0pKw6bchnlR+ABk60vlbQn3DUQ2KIvaCVojKfKvU/BPH4yjFo0OwTIed
hbvc8KX1J2HBUf+cp8o5/W7YJpTvwxa/A8xxksxNKBhBPGU1Xti7wa7cU7QgLvOypuII/V+xccUl
rkuGCp6XwNfh0g3ENrdv20KtbB/mA13U5OjqX/k7xffdP5VIkFC/Qrs9pqGGX0xi4ZJjutfC8bqH
uZOEo5WT4+HOYMyZX3+8pkckCdBBWxqFRGqjnsZu+vcZHcVqp+/RXy0x5FjgtAYOPRLxZIRztArJ
3zYK0DjHi9PNCUXW+TxoK0Fv77fEU8XLCLR8dYe+ExOiAMG6VqsnxPFewzSP+fp5yzCT0sgmyYB2
i8qdTCvY+CqcwkXSkApcGpyifuXvt7iALwCMSpBgOFpbsFZWATS3d9nBeFyXQRZoTMJjTdbdBebp
xzvqqjNbUdXKhzAEwrYxwVUo1sgtWDKH7pZ6MzK84pwUnQf5qO0dFUggg1VEvoPR4h+p/YCjjJYK
asxx7guadjP7MJJtruDjsYfaQbQKV+4DeIx/Kqn/hkmUNRICPyclhnLZBz4M61gcQ1IkpCPEXrbW
DLXl9Zxvud/ZRTyyBuV5Mivz85Zxp7qFwpZh845u9gr7eG5hS2SRHqDT1ZHOHZCgE36C5h8+Z5LW
8qfjNJKwg/Wa9RXvo2xYs1ZXRm9FwMeskWDLEYUMXJxZFl/malGF1onZDRfVnYq5H6eYxg+AAq0U
EPnqBBrUhjSGSnqmpLCCpCqxZ8/eNpc+p7tCAACZxrxf3PJiapm+aoDVHFnEhX7lbi020H8gSfKq
Fq/OXkiWHQL3gfxXZO/MJiogsGMIlMjptTD7PO4sMtQFErrjkGr1zz8dsT/+Jl51x3ZuWo4ClG9g
8aI5W5vPMrFtSAIkhW0tvXa+DtrgSZpJkZW6tjBmDhA9A1Dv1LlNrPsA4PJgjkgFA9cj2a1tuKS3
91n7fkqG5TuA5lRyhGgLJchq4Yt89c50b2BckkGkaRIM9+9gr2UPbIlF5VkeU+Cd76wkJ7TxTATM
RcaYD/VdC/SydOhrz0P9eNO9VrCYVp2E3gL7rvGjUvJOVTdNnyRRwKe8cA1AsVZIxG8qJDrssdxM
6MmEezaDcrLl5rph2UMDoJChLdv1lDIE2622rnWvRg/cIPki/GtIWnBypAbGUXO3RUtfGYQ71Pat
pmVbeloaZXMrrADplPQ+5o/C5ft+y1I9jz34XdwS/vI5PAj7Pmo7pe1wEYOcvcWDYVR3iIKKIr+7
sI6jLIYmNXGYMmyrcdCLhPu90rk7Urr4jX5o164UxKgx1GvrVr3qeJLEfq/C1uvnMB07NLS17GHv
h0xLa3lN99dCMkZY0fm2mZoeJFXmrsFx3yOQL26RgJZhmBjfE0DST2OyO3a5IjOuHBrmX7lVvdp1
gSwMUO8hBWaFGXnZxBmCNilZBQjTWGo2XKjlgCJobGWLWE0CWKhkxo+A5xsoaFLS64x12eqvtgiy
7rLMlURF1rumaWNYsoPWN3xggNgnUpbtU+qmKKYGuZD/wAHZCQ4oJqOwZxDQLduhcEr3kADMMUr2
C6g2QGdX6fwgTaMixpLW21M/LGlp+HFVYhN6xAItSbOKNich4tiJYFENKKqM6RYwsiGp4kObQV00
aC7VpMPLJdptFih9n8GN28QEEmzLPBRiMXuQF0atuQZMrRwOHk9jUKsycd8y5sYMIRMqjmTO20mB
qWq+8LPU6NqqWjE=
`protect end_protected

