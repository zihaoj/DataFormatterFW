

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
F0dLfpEqn0YUpcuwz6TYc9ZKmibaFfenDinj0DY13kDev8chY9t30QIEktN3YYHRaBSsRPUItx8i
sx+31aziCg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YWL0AUrxAFUIDB4XS03EHrO64fqZEK/v+X/U2fxixn96qRsRvvkPdploK34Sg5XijY4N8SUv2aft
+52mgzHagWORZdoqEeXql0CUk179k9eSj3aQbugSDfXDt4yzd8vNa64ViTwBMvMgbSvK8y+IyY+1
3Uuf8JjJdq/Ha3ZR+3Q=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NqZkm5CTHmRlN+gwwPhT3OlNKvzkAsIjLovjZqZsp+CYQKKsJa4nEfopvASGp2K2A3K5qr15KSyW
ZPGB9GwvQ5Bcb7Z1X3eW+IXPLKzMCZ400LAEr6ALR8sGaNKtpHnmhqDIivJGiJnZAsFN/iwvT5Ui
6+36qqKvWW6v9SiKHgxq8jgiuR2NlAhGDvg5vRfZi5L1YdCodagLoJZorOef+5GSVHQ89lA7trTS
uIWejPuM2/smsc9U1MF4LSYAxX5ejDd6KYAdrEJNp5VqA2+oj68IepXN+VOJs7JJ8hlG0OBv1N6K
bX96NkJtS94GXmobZmFCfaGSNW6y1C7GkjDs2w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iLv/smVBmP5OwL/Hwif3w7wG5zY5ElZnuhPGEQJbiK12Wy03qenYp9psKNh/ta5g5fAEExB4cHY3
eBHl8usx1goL/QXvr6Pp5Xmks1f1iMRVO4KKg8WpvycU6+IDApXdER0M0ipu1IEvpJgXExpO7AXQ
Q0K+7CW2DKKBNDHc25k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FMeHgjC28SkmWG8MKNBTIqMNBR3LVVKXp+UwNASTfvMqp8AiytuWkTUds0tPNB0GgYPX3/UWApPf
7jNIFg6xOA0tkrSJKGc25ZSpDeLVzfKXelVS56ddxTnOCNLgSFGYX1PBngWyHdxQchktb6a/XIh9
K5QPHrDrbdnhQF0kL1Mi4nFEIAUQ7v9Q27PYpELFGXtNqrX884TpE9QF+XIP2aEeJgtre5IGZHJX
evz4xvPqnUGVBBsazRYEuXdn5FLOsNG2hwmJddRJxeDX8sl06tuyf46Wq3wXvnshg6qa5BGdTh3Z
286hv4cPC+kKUZDZK04LAkFrt2yYMviRIexEmg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5504)
`protect data_block
tef11Gp3H0NV1UJhWnc3jXaGvE7TBWGbj9aLUSEvnlFryxUlgiRLzIxgEPc79LGDVvyDPV4bJpDS
VXRvgCDkMW3iKNbIQeyXAizhkLIgVWBC2iSgwZVwlbx+ryFyHGh4iv3gxKdZbyAU7cfb73vyo7r+
K7J+PCfRaOiH5qR6bC5zgTekqNMe9WLJHTyDRfe80ICMgHlPMN3DXpa7a2m2WCfVx/l8VPW0RgWb
5ZPLPDzwLGxQhPuN4FgJw8TtYM57ot659LBGu6q/2j+A7D6zWRViKC9SRBLlicWK/GzdQYyoKQuG
8Cbr/5zyC8Lihnt7W1to5JcPNpM8LGU+dcsaFE77w6vOAFGkYLorcjNqj2oDk3gNodyDsM6gUt7/
3yahM9eaedDSboD7UqUjcF0WtefYPSGRBimYvKVts9xWKOkKMpZLkSbuDv+/+Yd00IVGZ6gGLjap
M7NbtGeaq6o7ujIgh/9Vw9ajt4UI1YM9XrDjc6F8Vy20ck4PLc39Br3dSlyGHwKyz0rObo25EcM3
b8ZFz2kAaUXsAtfDBArDuiHD+YFTJUOl4RSoNULydVb8c9uIm3+ex6Ub8EB7kPvFpowKTdZheeQI
0kaTtLAg9EWCDXDFMHQBKlUFWZdsPP9Gw5m5tEL4vEUIH9XqbWoa6sjDM5nJvMWfs/mTKFxFFatp
slom3IJOCld+OVgZY/usayDyjt3DBKOheq2deq6Euq2/g8eUza16nlW6O+JJo7jBitmZzhOOfcmc
51hpJZYra5+SnXV+EPO8dQCGK96z39qJm5tVI/YvLVCO6zG9bvkMG09/Ips+gGnO8/Dh1atP9OQF
BVp9B/0LybZ9EtE5m0z+26upA8ceegWTK4W5+vrMToDUzmfYuRwTtHymS3w0P87OUaysOGNYqVT7
7kRzxZJ94ODWFOPlTq+5DToVcrrBJotxpeqEptjRgq6sPAuBEwK82SfPqHqD1hSlrSFnIQoFILpq
zloYagBZTMoG7XYaQlmpD3VTHMzuR+Ebn2FiGQ/UV6CtXfv/NjrB/F43RoZvMGf1bhi+y+fvQRZ1
48CZKRLARvPbpO59JZPd7r71SFno2kyNpEDPbE63Ivqt7UCY0xm17faz/6M6JuD1zLT45C0qiluQ
A+8FQLtZTb3d4rBW8EvWJhJNCwcxXj3PV2VslQwcSgQEMxee59w3ck8oymtE/mDCPd8yeUAYczby
9xgaCPt48SAzeo40hLImW0TFVgxbWLWplmYBDw2z4BwONYC1XHVdyLTmdGmwX5L+bngCyfIZFxUe
kKZfuPt/eIG9rLaorAbgDagum3xQkDljjQqW+XGdKiOEXWmrYDH7OBNJ7CuUO/1qkw8TP5ACdT7A
xyMOAZsUoXaT0kwpgV2K7HmRFy4v+YNFeAGdXRiK+0wREW6uJlbUMbE7I8D++xr7bBgg7vVH4Cvr
C5PYsLqae0f6PTyzxxugU2xHwTXHjblSyxgHyZTsCNnR4uBb2elkX/iCnOHC3zdfTEE9VBNSyQzu
Dfw9rrl39tBSSlDa8wvsTC5vvSVENRNytNLJu3C/BEL2llkUpG2Mcd1LxLL0MufDbwv/7oZaYk/X
tWGQbm14UNHqdqJG8KDJzYjQW6/TFp/MU0yh5cULg8hCNQWHW7Bqt4FYajbl0MVC9BXpZqiM9Lzj
8+7sD4O2mPCWNZCu2GaP0QEt4zlTaOE41UGzT8aMXXMsiAV+oAjsKe4ZEXWJ2PmjZoMYUYZVX1qn
tNVfdIpa6QyBKRL1VUFEp3uTFiwH0M69v5qmUFvhEsSL0SgUOpBb949/Z1L9aG/0Fkp8iamNvn79
9OFAYWDEyktQTM3v0Mkn5DpyLllsjccGlOVnX8ew4Hl9XpvQBgYTgfXfUYyg/5TcPaJ+8L4vOD8q
xEqT0SP9FtkTJj6dGNr+UjXIwIjgcdwfyytj7pfHzRQgqHhUDmg4aK4UfDTqU4S0T0KvqQiyDBgP
7vWUjE02kbz5lXExE7bpSFCHDeSSZj1Y6lRKU7AdSsJdrcllqbuU2u5LzFLcvyAYfJX8alnYf98y
/PogqDsrqb2VHa5STI3Q5ymV/4ZXo8CqzHdmD/kmZ5idw6q0MAV4tVm6OwGE+zYQB/xbnHnpwKWe
3plFHDKVhXILnu3xMfQrwkLx6K9mhlA43s2G9j2y6Ms5wTOSgLBFVp01mBqp5zzJa6ttFy+hHTmF
UGxCyGCcIVWqoGUwgG+dXfA7yHMJypWT0+GM7E4ZhGpvo/WSfJ0Rzs5WZiEKrl+cIG4Abfa9WtaC
yYnIsGp1cJvWJg900/Y46vSIhlr+5DrrCAMIVT8+xc1djxUvboNV7CgA1Qe2EWjoqnqWABaUuWB6
KG1mEzrMEZRawJ4HqbcLFjmYNgPSH6LHFdz9kdBIvLH3NiRrrwZf9ZPVZM+h15mcAwl86lQTpcnC
xeuP40YA2tjgx4rWBqb8BO26sPtcirHDDXxIItEr1RQPoOEM2VGqQP5JkKG0W1lnddbnDjt2C5Nr
AiN/sT/m4culX6P4DF0FEt+o+XMxoL/bmy+phZIBb5voB5OZQ2sLe8/0jBQteoFp2FsTor4QkfHz
GhYZBOinGVaV+l6FBFQPSJdFg/wfeU/RVsvbwwm7vlVm0zjnDyIgogT1hoPSqWcN0QRg8YYRWcVG
jhnRmzRWnodQIFLBbNSfkhO/70s2Bw3zXoTcbwCkSR2UMIEPPV7UZnb2iOyBtxL4pl8/HTi7cHdj
vqM36tj/rA64DIvPOdeQa4nulN4/MnEp4BKPLKjBJSo/drZldTWvADnjsPJQLfYgeLhU3ZOZHA3Q
p9CdooulnIIIhpFdET/BTveoUfUeKbGpfq1biSgn25P3EP88PB22YZJFiGszw4tGyLpgP0KduQPA
HY3sXHBHmpq8NleezfE2PhZjWVbSGjIDIcInAW2TA2H30kjvbe8dXdAO2qVc+iGVxhLBdkJIQ7lj
tSgue3b6W5w6Mv/c3iJQbMMe+k/zNFImi5/c2kwZgwpsLS/kT/J3HyIDkBIEX51DCBGFLMPlL8NL
tZm1CuqyyNx3CAayXCjeDzE5dyam70h/DzuelXheqHnge7Y0cZ/BJ1P0lq/HIGWYiP3txB+15/Oh
5TukdRNcNAh2SAPPD5cEmPWwS2PB3xtD6S586u1bZrbiCxIys8geaeHh3oG22IQZfEWQPot2pqLy
C/ZqOpMqMsauvXvAgII0jpFeIIHSnt3rMNVaTVwe9fzhrIW5VHlSQDGbz1TsolhFkViqdmT2eCKB
NFrzz8bsFvA/mwZs8HClzXULdlhJWW4JxZPIY9hBAKR1Sc3Y3aC/oYdzRe+ILArcwgP2M66e62aA
unXv8dqoq1CpSMoTpnJNyx9FxyaaFHds1mB2bMZE5VpIeDENVdXYImAoQTVUl7sNs/wD3UtMcZKC
qGRG9XEE3MHtHZC2127Fgy9wsfGyHotPs1Dtt/u9nfeNMFGnlpqXbKUruTIWzzcB8TbScqjhhMWj
DAl1uun20ja4DvAU5/MdjG7lUHUbsP6pLIdL5i/1yvW/48FS8wQ/ZteELIHsvhy4JcBWX+v1Ob0B
pRj4szoSS3E2bkC8OvbK5797Q+XBj2Ml/AZ+J7Lsewjyga7H8uTivrv0gWN8AEoqDQnGcLTr0BQr
T3WdxFy5x05BskZcXZg6Cy8waHp83Z5fbRV6HqsnhHH+QsIfO4/1Th9qPswK2F5XBrnLLClIixEg
icpU962GrfxmFBO1DMtn05l0eTNFLKkhzGZStcxtpnNKAJ5J0aiyTenjx/ROXEuXdDivZeWTbbrb
rz9v0optxzWsx9CGK4lzYOBqkdVFk0GUGsDojmqyrvwxbEsXw6SYhM54WuRMSjpvBTXDa5Iyz+g+
HkTrj73PMlJZUQ7PbozrVTcmvY79RbAAdjIzf29zbaZnb0XWFnK6GzuqCMR3CnymPnO0fR4oaqJm
5Gza9c1SMjsuu3PUfuwDF0UUQKH1wRsXcq3ANYu7MTuVS2Hq4ZkLLAidLfPDUih+xfchITFVIkTM
1jrdg7wqaQ+ZcWgpuJMHi8sGoz5DG6G3f5WjNnnafBOUAuniU88H+L9dktzi7m5FWONQaPLCPUqY
8RWzlNZFnNyZffbqgVN4QXZlqUkU6mrjjVxmWTHECRnDU8FEhI8/uX63kgTx9N2UNBWQlHtvmEbb
mzGYpxoDTLvB3Hiop3vy+XqLtqlCCzu1ALB+abtRltM0pT8nQ6mDZR2JNYS0GywQTwyvQ6saXLoC
SQHyXus3cXXPMi76CK7StGKAnqWWoh8hAM1aBcZEV2oOIztBHOs9+a84pp2315mawjWvshKbWl13
vJHqzvK6KgGrK9Nsx6R9Mwr5s5+Batb0vhuRuiCevhYYz4JJoGfWWNNCFa8fzol+YorLRKwsesDG
jVv6D4GGzdIyx3zEIyf/ZcoFMWXc5KFTGr+AI/l5x+v4pDmm67l31MEsno1DVtSt/n+dDFtdIcSB
nP3Er/MCrb8IPiZxNsjkXo3G0TImg+T7PWyPkM65pr+tFiauoGuzOvKnt01zNn5n9QEpeNpVv8Og
gaIN9oGisuJf7PL+QwRRth7txllcjoESiuiAcL1IjpXG4mx6720299W2tB/ClAVrYmam5+ZgJAZa
p+KxhefW8aYiJ6RacQsaWclT7laygpl3FfOEzrAhD5fMI3oB7JzrQoTvB1u2ZTGkTOBmhHgUnKYt
skw0IHOd1g5aAAhJu/m8ol3ft+qTPjXJIuiNJaMkbg3VuYj7Y9T5dixDhTZ74bNHEPuPY/Xk7MtN
rNXXIiW9Ia3WsiEKNkB4YPcv+Bl920xQegxaYLvqM9MaaezV59qSlEZeu4m/VY2/N5txShp60egP
yoN0w2V42pntorvrd0g4N9WxyVHaSR10p3jspr/iLkPB+jptHbur45NieX0g6JRrkakT5ADN121X
I+p3Yu7lcmorWnVv42NaPjoblWWB7KKxyHRpzh7UcKxxgFDhD1mrS06fGZXBsiBVu0Rp9s+9xeKL
uUZdbO4//tXePKmlt71b9bWvQi+6pOlrIs4OPEKm2K+sVINpcikOFhQ61+8wCeLFGp8fCMs0RQdY
NNohHM9T94pb2VuU4ikSZ5QEAO22VEfz+ZuK0/1Gt6e85saedKQaOTLAPwDG2+zE+KN0CKDgWnPg
COS1IHCD0Kz6vuDYtmyU8/PoiyHa5kdno06XED7Fuu4VP5j3srjUae8Z8MCZto6sXs0ErzVODSAD
h/tTn10Yq6yeCUSO+XU2wdJ3p0KZas9gAErEdViuTUC6J7PYsCcNQYcaEUjQBTDmPTx520/gWAKT
WliJJr5DRC/W+FdKMxWgazgN3L+7o5J7Mz6SWekzqYUbRhNrYUGpvO6dScJpOn61NqN2VLQTOVPJ
xzit2SOUd4id3BTGGfQEdvTl4UylJF9GNK22z3K2yN4UjPshIHG+nfffs/wygt39MhLGFVhM0Oul
SAQXPwm73+LRuvOKaOftUIUTp484NqIZLizWw/aI3DA+dSxlAiaGMq1ibWGYTHp5QiRREkcS2GDG
aqIXmHX8yv/OXqdgKtkMyLiiRCHm0a0hm+UGhxBaJdZrGbn3Luy0zsr1lkv7vDBoALeARNYX1vp3
gaPdn9x++djzyUp+j4tU5raTzZtDHsS6m3OEclYiVb6TMBoFvomkjfyIUOrruDUHYyWSBp/kl7xr
tTjLGoLKhndTSTVlr+uqT2S7UNhhIYkve0l1ndcAHqPtuw/RYZDGGW65kZEM8Su2i/7K3qsabWOu
xnmVOcMFfd4EHtxipfkTU5m3J259qFliSc6Ep4BGJjJFzCiU1beaE4ZgHCTUg0nkyt4RyGTuON+F
y2EUurlr4mpZmUTKSFmdeGktc2IPf3frzTQZLA8CPQlIZgko0ak68fqL0A+shwMMb/liX7hVH5nQ
+dGWWVVxVtI/rXBMxfKtaSTgMH5JBV1Ga1aYNuqmeErCnuBGbeZl/hjeAUmvASXNIgozk1f9LQne
8Y2J0qx2eXbgBE0kju6AyQYr364ig1YbnzQ7x9B7KqHd+EUeyjOsb6zniXef2qy7R6bEx8uxyqZw
uZGpNmry6i04wk6sIxU0GWjYR/8k8PcJgXFisoKlq//M/sT+6WoexmiAd2TVS2N4AOMpHvKbbgZ2
ztT4NlxntKXcW7TwBFqe1qf0l3NC3+nS4NAAFv7bqqyiO2Xx46YnoGhiS3ZnLFAzCDc06VHntOHr
YeiEAJAnVYtgw374W8fiDBE1leP37tfYgD6sTVkru/Se1WQHiO117bJ08/ptMZgWzZ70Xzz/AyZI
AtyAsCY8mckep0K8QDVWjQEbehCaswjWwSJdBQKam8upzZG67ytr7cVx6J4hOo4Bo/N2EORPRQcl
4tZfvIrYC3yipA2XxHU/n6EYEbDdJpASmoHs1RUjfwyOrRXtWNv7vF7/Gj/5KlFdiNBS8yAsZOeT
Sh/dkiMQL2nxfoFcbmfcX7o5W4fF3x27W/tuSv8QPhTDaH6lA9UA6kJbt8vJFDVhPeeZ7qqjWNgs
Ff2AlL6GH+f0lkjbr3UQPoqinkFoqELRy1Mp0hTSppbvyXNJg9AaKbvFuMfFQBB5XFVYNnpgv7LA
Yg6vwebShtJhkMfN5lUIm8aUcecMcZMoWHjwqcKOdFlkIRaRpZJ9JWF6tCl8CCGUzUvw6Pu185is
jLaW9mKdrlhfc2PQDi0aTHafhWhSKrULznIXV7JJ6AtSWQpNkV0mHB55eRzz0guqEoIKAnPXisIb
uQhsdDxdi/T59j7Qi9ATaQGP+2NqLWn9Zk6TPC9ZfP9DG9BMCettzhxip3pUbS9zgPPdfYOg9/ey
turl/69qo460sY3p/X3hQt5kaNziCXXA5Tp++GzgNZRYAAhBg7rJukrxHmDh283rq22L0F+CA5Ai
EOK8qFc6ZJFSRoaVnnsMYG1tvPqCd/TkoUiAPAzkznsnB+jzDq/Oy4YagSCzT/ExGK2MSLdY/Pk6
cuvYnzjrzXgMTpTvV3f7DIExp/L04D0yQ4taNGd905X63Yt2gPjBotZLTPHyqSSBd2X0PMLRT+On
CFGQ7nM6FAkXTQEzZfeWkU+QYByik20o2p1gHhr2Z1K95RxXkPPK1BfzZAQxwE7WeUCfulsTXIW3
/RhJH+NS934uAUT0U/lCnQwpOmFUP+EuccH4jJE7hYFtJKkyyIna1doImWeZ+fVvrMkW6Yw3y/PZ
1nWgwXRl569Hiu9x0GnmetPk9CEoxsH7W5BAmHvm+lKwu0K82Zi6TkzTJ7VgYYbOta+zjT1TOK15
3I5v2RdHox7Wb0JO3UI/Fnv1UM4AIdpOrhuHxH62cj4=
`protect end_protected

