

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cE32RSTvXYb6m77U0RUuhMrh70/RTLzajd7haZYSXDqjXBbOkMuhmdGgwPsX4IRozMfF30OOY2Zg
cQt1sy403g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CY525ALSmVJ1bfJ6RGQOsgWG5vbLyb3A85GFtotZAk5zO4kHFUX2zLKu3IW726N076aUSLr3vXPf
Oli1CD38ASBM4ws0COi5MZJQWPSLdDknMEJAKl0oLj0m0yTuNfJKpvRpKfypx4y9dYm1BaYxUSUW
l31pypDj1tlvE82HG9U=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MJ1RpAh5h6WDM7VJMPVnaH7ZiegPdJPPCSivrCDsd0xqxSx0GAxaqqMfmeUtOb511lGvdZZfePZM
6hirl35PUB8TO50mKrjpJMsCSPEsjxnu22z0z78K2WrErMFaYZWitHhHLveOzKMjOpuC7HuZ0/KC
Fbr7g5pt48elTJ9lKvZtUE12Bm/I4kV8Nb5iL2D7+gx6Z9yjuw1ePehvFreJ4y4PPE45R88eIxYe
l6aYLFbwQRb7+OvxrMFNU6JuVJgHppuGYqszhgVvA2KfvjBTtp1OR8xylerA1zkN5U/U09hhhaJQ
j/YZRr0HX3lAtGRaX3zCJX6hHNNg3oWn8RC8Hw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tYAPVapnqsddRargk5BL8V3VlXyo2pBev77Cr73Ev9YzmTYFWiHCBiCB8ZT/czUvjgo/UmF2BDY9
m7T8pzMSOv1NWDP85q4MjZAbFbgaxGO9+9uNc+L3Q82FJBqhnZsysHkNlWP9JTdyAzTlNpz7dL/A
oN8DrDfwA7C4joixy2w=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mw/yvv03pGlOzAE5woR39/UkbkuO8v0L0CwJVMZgyMdKDOL1QfsrqOcWz+p+PgnQpd89OlHw5c1j
GNFt1GcmYxLqPl1aRcf0n0yLuWT9Qrd/BheyqObKaunT2n/uAmrFHlkq/A2jl8S5hK9mYWU2+hsg
4D7zmmeOtQ9X9TfB/WNJk0brWcE25VzeWbopR0OqMQIwkm5vu8VjFWUjhEWoUTTQc7UYTGc8zuJV
uJzKkh2svTxDEjmo+7Oc+3n1r2AH3fKp7/Y/rAOIVCNjaiVHnYM4IbhfQtQlapQcmWrUinw9GA0G
4RF9Li7t2MKgZ1fVBjS0X5bzo66SEdfT0Xwe7Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9216)
`protect data_block
3S4CA16gVRAdbf7BwuUuqhWRiSJfYUYZZYY35Di8v2lSHZpH41rQGGAaoiOjmsz48qJKmsa1XZKH
C2sRkbhvqIqF+ANUgZIRCzhknlGpgOyDl3BlzhanEI8cV5/mnFFSSSVlTPx2/2s4YdkXAbTEcNev
/11wXILpnIjatw4uubl6Qrf/DqM4a8VqAxddfeP0i4W0bwzDwwOWPiiF5GsnFvvwfRH+U5R6Hstn
ZLhqQUVoJ9F1bZUKP0E/o1Mw/r5aT82/gKNcnk5fZEeEH3+wRzOio3iLGUppRtOq9TWoASVL2Col
Fb9UJ7+yanzKCfwmV0dQ44wGdKWNJMuo0BA3DI5/cLfSGYm/61yzyXqh/vnq869zhpgtVBpid7nS
zfqmAiEcUPCerLbZTBf4vreb/eq2en9CRl241A6oEMyxP0FqotSPsnk6dzXiDuw50NYDfQZb+IzO
2TP3ocAOHubcQK7DQTaetMJMIFCBWwQnuCiQL4T9xMriiCvn5fnmwttIpJDf/1CL3GJtUxIP65aH
SMm7GbKurDjmVuHSHjUskYCPhgy/3mG8aMzxPEfqwOevPALfjsnB53pebntWahn8N3k5qYeRu+7V
g8ixIpGIiCP4rsnUNzVK1rItk4xNCxAVi+xVr3gR5IoVBeia6k58XoOkKmo+t6sFHzGAgQTC5Qm/
wzzA1GkF8MDX342tchNnD7KT3NX24X8WWiJx5EISIrZkr93VrI/hUdeceCL2L11fzRlB9x/YwpqO
mVprada0/Usrd/7JfuCTgOFWT7zi1nwGDALp1fR/YKQ0CmfKKJq7FbenSbdOHqhcvmoB6PnP+c/M
BL6OFB9iI97I37YpxwL0tZOmqjZs6Qc1Q9ew/NiBrjJaFbA9hR/3u5bhL+p4RS/vxVLfbJb0PP6V
PWd0hidm/IkMTvIPqtc+kH8jixj8J+iqs2jIFyoR3sGEw8S6nyjEluapiJq6VLtupfgZSCGnDYnm
qu7hN8S2Ps5n0TTOg+32w9R81I9BXb49nABs+KyNxpOJ25D2UGZFMUx9lqFhva3Lox8BZasPIESh
y2RZC0BCCceeaV+CgT8A2wP2mGojlgm/xjNe4VeWKCu0AeTCzL4fuIIUb5SlYbg+xKZBdooXXgZ5
bz+0J1/R7W8j/gvJdme1nkJhVDvYYucU3hcYyByv11wXBXpzmyLmoTDxbuKwYBNd7aG6wpRlFm+l
ojvlzTEF0xnULr6+66DfN9uHLCFo05spTrU810peszzCCwhUgcWHUG7NmFQbMKo6Pd4YsEWu5nTT
lchFVaWRvFcdFZz8xLwp9nl/O11ByDcT38oAl1azq6HR9KZXPtb8+CidIrmcfyozfk1ST1JzqJS9
DW2DRqzKNTq6t5yDeTt+xGE8c6HmS4B5+Dj7IJEJsIDC4R/zqFhHieJlPvMvLCb5Z1R9qlha/5OE
8cq/Cy2Pe9NisgW3hKIw8FsDmdGdwuSYYMeLLpqkDsXUJ5xZ/soAKSadzKahIeYkDuomBBnBZhUw
ZyRXo7TqQtUqxjKZzUdKqJnO0ZT7z9hv5JgBFnORGZmgWg8ASAvayQlaxo1BbWbDUa+FiIkf2kDY
441uio5gAjQRWSAUzQb5v+fs8G6BRLm+3trQN6wuj/xb4VPwrsLSOosrUgB9OwoeA9pwCCorBaRr
GGQXMl1cViByE4mrD+mUoR1IYD/04QJj96dW6OKZ6KmQBqRV+ovBaatm2b1vfEfBBrFHfKfKr2Hq
zp/pvc6BYKqXEXyepTchHKCloj6ED634+0CDK0oF/wU0xbbCB2AD3JSTw5PXagvmQh2JkVOYq7/G
I1yJX2CAaLRYXD2ejBgtnF029vYJvZKYxbTi0WbTa/xR/qU4N3ft8SqNkXNrX7FOWRL+1F5zwxAt
8IbbQ5+bNrDUIIDmvbjx0JJ0Z4OnzSdJPnm2kJfhuGG8mxy/o/79uwzT7M0aolwmsA8yN0KH/xpt
vbzfXbu1dkof+7QIejPJrWGC5BwCLEAh7vtJLsVpNfcM+Z5H2P+m4MR8r4/OXA6x2hfd6VKpAHJ/
+JhSi/01BH7jxALtUEZVqVOYQathI7yNzK+nVl81ZrjcuZ1122yjZ23Gp0iseLeti5WqaMIQi80N
1RenZGgoTkgC+MciPyv09C1DZ/CANDYpfFm8/3YS5nOuHvy+rHmwwoPufq7vmXeNT7xAzoyL6khy
PkVmeFCeVMdTFpYMM2KxJGo5foEoe7WKiqXG7dPLhQ7p84DtdYvow7y7qeBY3dUCPCiBJp+YuYvY
z72Yi0OaWU9RgLJYwkpicXmvPLO8jJjQwXAJ2vx62dHcOTIM/ivQYqSoU5YdDYSmm8gunie38hng
45/CMHNZlN8Es+TWUKMUz21Fv5eAnN5aG4g+Xy51NbFJ7s0I6cPV0Wb32GEZgofYVoiHg+UMMvPg
2atiIs9Pb7gctk8cPitN+cLWr4FQeYNvHrgBIST3+ZtINoimKL2qYISrVzsrjcXPxSf6f3iAKUW7
u06KMhEg/hbZh4JouqY32JdFzXeQ38gfbPGkYLNlQvFb8Q1SGSkoE+2Oh8W7sbJo3ZrbeTiSlbLY
XLvQSifIsqXkjmgnyzmGnoH3tiUiF6xhRfwljPqI61xWAoXQDPyx6GoUG5TW/Xn/BX4yqvEYtYi8
znqwmjcX2G54BVyMMkq8CgZlglt0VXHOa+BX99nnoNs4VKjktocJ2oV7TBIJWbU3ojHBMUBOjVm6
dKwfDVdtMSZtvDqfLfvccY1GdcGd/szQhS/CtLbvfCCTK6tdzn3PSphwzDJPkGnkQNWGlh8Ynnts
hpUHwLr5PHu320ak3lE7TsPL0xfzo1uOwqr0+yvXvyqwVsz1MzgO88Z36lqf9OwQvDRYQPTPdhT6
Q+xci4DL4oKoj1ff0VhbtWolwTcoySzU1vYnj5QqpVNmTbiqQolSXzSkAx1yk6WC3CY7SuP5sBzD
9WFzyJsqPT0vCngMVzfZ9CudjJsu6crovnllhAwAgvXcuFfJR24Tex2VA+xpANVId+aGqMJxrqRQ
IFaKxdI0ZCsOJ3OranY7kBerBUrIrCUnsTh6oU6YGexhtwNVi3e5U0bJoZUS/LwqTe3+3gZMLC4+
124EsgJQMV4mNvV+ds/EuAs/48XzPYQ1WThlRxXcguZrak0P+NL+jmnBUH/q5hXA35F12TzdXtpC
BrL4NoPnl5hXfJwBmFPwsK/6g1fHURY/lud0u0vgA7hCKh2C81ls5J9D8DsmY6eWBMPi5NWxnEek
9vCcRypuQhg/0Z8Q5LUtc0wBs2Z7G+vQioKJ8b8ujUDpvwqpZGg1yyZeaslMFQSo1QOmZWHOt1fU
jYA81IILKYSlW4HzYBVeIwav9aktv3R1e+U+OvTnFeY96nw+fw5h8v4cUAVY4qcEzl43804T3oqg
Hhgj+5kTYSkbVafYoaheWN0Vas/DY2F3cfCBqXX7Me4IIhBuBYNnyN+FBAu0HCyDRL5WClNK/Pyn
5OmH0sdlUdi5kogniuMEzojH3SivRPZNVBhj2QI6SL6n5AddZHD2WHs74l3XYZvFoLxwrCM2zYc8
f/CA+3f0uVB6tF5xoNzCi9MPPKbufsmtiU6ZbQS8xDuePpCPOZjXajpyFDA6EQZ4H8rFpngS7YH3
UW249gDA/TLc+11SuHDKRGUK+U1Lqt7ml7R1lRFdDmLEzEe0IamnYT0XzocLA1hoi6S7HRjjS9XO
RcBeIXt0PsBogOe2sagKYpKkR6f+Cai+CXzxtSYe2Dfwj8kCaytdDs2Hjozbe4jTQYRa+sXh1GJY
K2MRHz8qWzHNh4trXbOCCjkgf4EsN0ORSkGE6up3Sgg/rSkBBsrOTkVU1Ay+h2dfR0rstSKu5/V5
2sMrs1X7T0GGi7GbYKsmuKt4sav9emlxLezIp9Fehof1vDBoXRX469dnXPzlFDqmCPlmS0Mhw0ce
6Agtwvpgr+a2ad/q2jsskKZRiUDlf7WVyfahlp1/6JKOMA5Tv1MkdsoklAkHmlwonwpzMJXFilbj
NuLMjxFdUK0VgxVR04HYY+zFGzamwlP9HVYNzeeLZfkRNMv2K/Q8U3gwGhyr+kNpEPs0wHf1m9AI
AYq/ouofKgtKMhUuKqiE+G6NAqMdPCzxAlG6RsbsH0bbBqk2TYXcQgd8dv+YSjJf2qSuq0J8zU9Q
8uOaSHxTWsJ6cNR6nDJ+2QbX9f28uw7l8r7e8/R+7yCZIs/unv0UJPz3Rg59U+YHEyW4iIgqg31U
DGGBwvWLDKfjSnKOqdCeDxfqCfe+khVcCuB81r4zt2GZ4WaBRod2hmKaABmIge1qsVZpneyu/+Rf
PRIRZ5+AwZGNuEWwp6D49AdylwxuXDAWSkUX+GVYMPeeoxlGRilq+xirimyV2MH0iCykRYrZNxhD
dM0ieSnpnyICCI6oZXMenqzUYL2mT4c6oQeAi4CkVFbw6lYo0dpMB6s64n6ahsRhcQ0t76Llcnnb
4/6riSEnpCl38pvMPOSNJ+MtxWHhiU7CS20DtYNE3C5wtCRi1Ly1vt+juM066s9K5q2OwtyZdLgH
PP8Tt3r99W7+t2BbT/Ym/RZ1qNeaXiK0AxI01V85K6shBBudSyFQ9E8jrkqjQA6mthu4I+GAk7uc
ULIHBYU44h5/a+tn3MxfKdPhfOrrbP0K5+tXyYGNRRQTXqUiFDkKG8T8vtTrmCStohrT+WOZSdo6
Mb+CnvXjS2zB45i4q66kZ4M5FHpUCvr2zPvsvNLvVtUoE2GEGLWZOUwHvVJ36Ug5bB8Hs6wvKnWP
W6RD9GL85DSMCfrGWRmt+4cEpTXFFELCtVKCzJS4Nsv4mU5+VFcNAvtuFMFvqRdX0PCV7r099cSq
lmggoxt52BArc3zBQrMzOldx15yBkZHO6tzm370knLmNmNCxqBYvN3gSr/Mj7anVMNM4vyVUaQnv
Au9jJHWCabf4aYfx+8CwxTOF9PrTyBmWePKPoVs0zuBCqycslCUAY0meY+mmuHqkLf5+YHxM9NT9
dRHgETCvKCYi7y0z/jQPdcNMtLYPVEDfdRVafnPrwONHtlvR0q/LUkwLq8p5ppgBFted0d3+QG6g
Qze2MAtouLrBvKmJxlFlQVf8E433hkm8MuD2edOqf6Sd6egrGdGjrvVG+qTPOCv/Sn3NGSqrjo3G
/bMrLXueWDiVyxBeGP1ZLEwKm2Q5o+vUEcM4YsObDOyCL6yqA+YNN4PeIfeiZ0Lv1Nxwlxn7wgTy
AGMWWHcbN4tbnyxXvuj0jRuNyI5lwIaHM45s+QNyXjkxM83Rn+cWLOPG6/NRKf8PEzKbNO7iHo0Y
FGPWqGu9cH8Xf2VZB5DWT0tSPW5M97udms+Apo9aB65jf3bm/4c8ljmXgChpVdNsfhmy7MbOuJof
OWxifpj3f8b4koymPqFzb+gdrLLdaGiAHHu1idgk6UFKHdIgx++lQNZE3Dk4kOMt/h3KeiiqRrJ7
90YgOKpMOtrNkDC1eRjzVsrRn3cpIfcFVrtwAGqQqUm2+QGeAxbb9yg0FY+keMbmC0liZkAWRaSJ
eR/wcvqAMcEYKdT9xC0qB6XbPHQBSy35RQaBx86Kl/zqnIsRTbx0JSwARSKH73D2sLLfSWSBXQkR
HUvTvlsGqszGnWthTWpbNS1hHTw+NfeRPLIzPwBgxznqdBqb4jgt5dZkGpR0HslYCk067yYKgOzF
ul6GNu/gz9L1DNoEDNVWiTBaTXl/oygJYxq3K+LSJuHZKxTwW+u6BDUrzAbKhfghF7dW5g1s3ThY
Gl9FbO5lyU4Sb+zAZjogueA+mCWRM+V2vm5MFHvxvwk851clh6Tm9ZPeOicGusGhysbPUW4wCFm2
9Lr0yuIFNi3C1m369WRFj5ITIpcPj0nyPpf0Iww4XzyMjXNYMa3Ukfk/Q1If66BuJwvWrbwFBred
6TtJY8uvQFCXvLAT9vxw8L/jdkWLAAsMP+kCfzp6VIA05kcA5YXntk/67uhznEY9tbIQjAg7nVjx
D8LV0Dox1al/i8fyl1of4t3+/Oih0vzsqf5oRVhSlbCo2/vcd7tCLQCl8Ssr3WrJ6ZA6XmUxV9HB
sNQXdJWX4JOhrLecz8B7YP28vcYI7FnLgrmUCxPKHU+4bO/fmL45P4O1hmKi/tB64CH25ogfJZrH
CI8tu4SSHPQpm9jMetPKfHrsuomnFphSbt1MZNQr6l+S2nTnb8jMQ7jHFvis41NDqsvhVNQjI/+y
nLdXPiwKKr+M1YKYbTas2wbYx4QPSWNAy3WU2jVKRnCGbhILi5V6SrORwmpEVXbR8tjieAds/Y5+
EZGPSIB8lbX61io7jvqAfS1NehOeczsnqO2nUnz5fm4p30H7c/4IGXMyeWDZ/pCZjuGNEeVG6QKw
M+YxdjRG7i+aanrnq1qPTZPgq9o1NZZ8rRL8AhLcc+ziiHW9ijsU2zn3tKsEWf4Tq5kyp5sv8Co6
ya6GJAgi6X7u87e4D+v7Uj2aJREiaSEdOGgNjE+QqME/TA1jskkIumyvtrqIA/Us9rsVNiuSmXa7
Y3iIyhJBki1AagGuQ+RfhXm5fzmSGPmQ91yphNdZDA85DhsWlKL74UpzAz7fut57PcHRBUk+6Dg5
zl4Eriv/3M3Aig5lh/yLYTcm+RRm/D0lk+OdFsVwF+6IybUeHjb6VPyJY/m6OgiOkLNzWj47Ei13
p/Uo60Z4CqWFsb24mtxuua+D+AdqjePhnKREcLsIIjpHNaYEaCBgc7l0IVAsubZJqR6t18dweTZy
+97cfjpvmRufM2dYM6Q3qooD+c1HTyNcta5YRjI6YV7u6JVRBUjASNRxVKig2/5wH6SEikrNzQl1
EWDAt6KwKpLf8TwGnIVKW0x/1pHJCuf1FoTdbuNwuwp9jW+BwnGCahKdg1y1WGzKX3kw85Bk7ha4
lC5yZp/3aQ6WzRs0ClmW54rF1W9rPJOL4NUD47h0tcemLdEmlRY7kgCsIjwOZBzAJp9H6gDWNXS4
nSfqCaCyyoEVaM76URx4tgsnGoVTLTaTjIvYeOS5HYy/lGUszGHvdycEZtAEG7aCDQzrPo7Xzshn
ieZlZYvscikMjdyQeOYV7UOppxy3qOVqVcEhOs0iANp9JG/Yp6NxAooRYkxjwxLC0UWLmKn/F9NB
dM7UAAJa4vq8muhQiD5bigMRLl1hg7f9rIP+Ut0S9IvLYjamIf2PrG3yJU+rqvej2T6J6BerHT3X
VISCexZgqh227qQnAdTapqZ/asGiTJecNmShApzNua4DWt55vNLOEzh+PUfT+XWMsr1OdUlrWYdK
K3eWaKRmr/cZpPv9J5g7A7f9LiWu/UxQdyLNLy/VrtuAjJ+EC3011Odg5BAQcEH5sSBusxKKg0Af
3eqWgHcsSlzazHPxxgw35fPzlBtzUuKWjYSBSEq2uwUH4iFz0Jn3XlK9juqJ8oCJsJs4uvXnmzi4
LNHXlIh1IZzwbOptJ+zzRYj4peG6P80EcahPNrPjH3kjBqN/ePnAWjTrTHsUy2HPUDG5PRL0FE5M
KG0Jpwtloaq7q30FrycBAY1tErYtQKK5KoWcdkRcsYnr8Un65ycWmOj7v53wk89JDDkQkZZmHLkF
JG1MS0I2SwC8O0mdS9lQ4qUxSxzNgGpBYXjX+kNOXspysyjw6gcRaX8g1wlF0CY7/y+4TMrlY/nm
GOSF8OZuc0IIEyu+7v6/GXUe1gjxqSNfbQH1I9K5WYWxhnsGutlYhWHkGLqKvCwQ1vRm8Pp/XYlp
PtV5KgthE8b/ZYIYNok4moZR8IsWMmswhd7Bp8Z36Te2PAxYaLyCk/k1D8407qTwADxm7ROAOgO2
Y/QIF92ivgISNeOvjdW0xO60zb5TnYkwajwBNKREmhbvfvgNcqr1TxbPWHdAp+qm0xGHcLMVzFej
AZt8aEsZu6iLPo29IIaM5x6WzF8N5UPPXRnxW6hNdJj8P5Og9U96F1Ah/JPchqm7fsvld1svUD2m
stgOm2fPFoQ8jaBnkU7kvQIcF38/y0szGQeL8R+LBMkbPn8FTZetbiu4Aoq09d7blz+9EZMDdi8y
q5KzYDXB7kZPqjk9i0NEF6RpqA+WGwqRFmuTGjf1aLlj7LdgLzYVhJ/jrOSfyGCm7JHtstu8nyhz
0wYoIoH9g8pJsclePZUGFGPI94isV9Mc7YMuvmxwC3DAzNzFFD97gtih7xp8/gveSF9u/zRIxLQn
XtMlxvDcFKOmuQeGfB2+/MZh6C/PRCzR2+erB9oL3wipx62gxS5HYITh6Sd6cBXFoMitzsSV5tS2
j1GJsrTFk7p9XJUv0Z7tE6FU/fY/n+Nih7uySI+BFkhaB0HJ5r0sPs3X9vWyRcanV8m6qrTGEmB/
Okz6qZ7IBJNeodW0X4THHpnEO81/7WnM1CNWpsRMFwEq++sMHJohLQceF8+rB6QR9Hx3p14a3UX4
rKJO9aD52ayiEQMwowMXpiHKoe0M1ccfirO8aywC/7qBKo3c3YV6BU06KvoClpEBsFG1zAMC0XQ0
v3zL4Rb16jLkACVxILPYDYSglQT49uuSZtrpPNpGhi0/uY1mZWQbdiFTVnWyZkckzsmH+7HsozyV
ISXml+2znlbV4KW80ze9K/vsNCogB17IXJg8qSO8gWk+nWiTPtcA32sp96Gr3v57a6VljZc3yBLV
JsOYeRWHj64t+biBMjw3/8ax9e9BQpEZfo+5sYoI2REv5twmXFjJN3YzPBHAivUw9idAtwu8azWB
C//KlzNLe+7rHPqSuYwhwDYTKdv8Ojmu9FTfYreyunLpDaaDo5enVoEI1ZifJEUz3cjtYinuSLj7
7NIEIJeHEGD47Slu+bar3EooZKHjVvC8iKHhsF3knPwR2kGCw8nDR9SjKC9l6Zu6J6/Pf7EgEOvP
4nAYchizXrTalgzy8v1ULeGYwCAhiNdHXM/6AOsEeuEYQo/s6+v2yQzw45CUAPfxoFsG0jE0jSVM
wLvT25OCHuRrLWT0+Iqis8r2MNG4eg0ByIwOcNw6E+pejD976sROsyp5EDyTX/58zLo4HkAfjCIK
kvsMn7td485m0DeFT31j3XKNjZqTUZqNANe2sSGHR6eLXvOyyquxBCnIszIWoBNGAluJx2CttRiC
470eueVloBuSi2sIumQt4hzyJ/iDZ/Y1TFHMB2VF7Kqe6bQvxQQfY939b3XdX6EF/zl37X9svsqJ
QrUxwqR4OqDu+Fk+LAVTeIWjlW47vcaAwgXrHWnFAu9njqLiI5bd1FANY1fOWPoT+DZHfhtsAHqX
s7uIo64H9JPOD1P0qdKnbF9BBjPU4q3Z22T9U97ENRA6sJFLdH3AfgfPIyJj5MYgbiIwiuVXoQK8
9abPKwvp3t+MgjYHuYK25o1T3Oy20qAl5xCOGanDKZGJv5el4rG9MlJlzMonkqXMm4B+ml63RI6m
6NurXIlytmS6ZmhcIECLXWgq6xCl89Od1gqZKX7sEa3HKF0DDxcXtQtZivq6L1ZYt1udsM8Gnnas
BTpN1GipOhrQpMaU6lxqY3K+WPP9pRL24ht6z9rmBe79+ayFuZ3SE5TNhHq2pH66S/4a7A0X8Tzc
eWfKkKuyBT03j1Mdv4MxTt5DvMsOBlyIbRkkCkpsDZXg5TdVoZS6qptAqV7X9HL5ZwqAQJVmmq1p
/pq1OKWdPdt3dzjVWdJ/iMRamXBHofwIBS7F9lDYc4ANAFTj654S7fWI/6YTsgJXtwxd888U8HAU
knqU3noBPITyZ1HunIZ/3TJ8P2757KZdrYGMMf7/HNlg38AQGN3BtKIEzr7JlBTsh15tnaDjB/KH
Z37rbgjwF02AL9+mOC1Tz8pikC+Yc+0p1i2KUHFAEq9bdmRiPKnpTJ8HAHt2NWaNs71WV2Z+16lx
c/oRSF5vmRyc/gQe339hnUIiV9J4d8ILWea5xzyutdNMwZOwI1VCIBjRQW7SAZSMvGSn+KsZo8Xv
fbycghmcVpN/14fVPrEVfgBBf/ASsFq8ay9x1aagfRM7P/PO8qTEV+4oPwX4EKlSHFk7OAkNPnmF
wr+RYChF3QukRCenS6+A9yL8tOkZATLKc2z+2YLUZTJND4e7GNhg2SfMjxOaK6v6EKaZ67diH9HY
X9j9w3RA45wL4PWUTR0EZTKihn9u8m/XLm6KGRPRLJM/PGgSfDur8Aqcias6/8RWWeTBfhuIQC2P
nbPFxRc1Z0KCIb+d/8pFVGYa+XPC39MA8LAbPWYoQqmpHtDeQhj+v5vL5JMQERjrjmJHhj6Pojv5
ZVVh1sCshS0AtbAPW2zWzIhaeUE2ahO3nz7e8rwO+u1KcnulNiagbMXp9m0xhJNgQPJRAt+a3k6t
XMr4aIho/UwIQsyk3bmTu8UCtAhMp4cmipWs0/8atgXBX5DxNQn5aJEpftBWtCU3tfoCf5yqH6Ty
0M+6oxBMj4m9jWTNrU7CCe3BVwFgulctNaZdc7J2sAoirFTk4Xv2zqIKNJsZUv45GSHAe2HlIdiT
tym/J+v5z8w2ygWQRShd+vOnPr1PTRB0+pRwKNfq+m/JLfNnOoHAYGnCBjG8rHm5YD8dhRdN6P5D
XSOigtTyuCmVgBIEWBaLLHJz094pyPigfFxi3kCvhowDS0PS0gjCx3NWTE8lcouOJaCn6MCLF1jZ
Q/hX6qdUK9m+u5Wg0cvWbMVmmOJges64soLnsSQWMiQ8JwW8a16g3gep8RPm3JXMLUN1kiGSNL2m
nkc/1OPUQCzovreg+kLyNt7gq/3lMdLl8xAbkeez6iSM5nN67msg1xvHh8CA34Djr4NFhAQCP1rj
26xuCtZiVRqt1TaDxsojKf5D4LPpY2MhH8+86d7C61XrR9f6J/30w90F5StWxI3TrQjSFNhqD8yB
i9/hfSNUEY/zesRhEj0antNXHtChyJSHI5Qh0HSAqauFJY5MR47u2u/hBZFVdAid+JCx7FaC6KKS
047HxrmkTPO+Z9KxHR5u5IsiTt/ZpwZSaIVawlOrDrXVksGdkXI0QM/Dtk8o2ST589tHE2sq0UJE
JxFIOnRiH6JQAXKIh8bRFjmvM0f71+tkOuyukZhydB2GBlst200ZMIP3tfIbo7IS7j+/d6Ypx2P9
NAwdaU6zMf15Az1i5i/CS/dMuvQBTKz5O2SSkvXxH5u49X0s/KFy81G5Mnre3rZ5w3fgNrBx8/rO
lppcQMT/fYsILpkFRBYPW7e+PPGu9nT73b0ylmYVZ1Loraf0Xx9EjRaeuBHXM1HD5amXwHW49ev+
AbwoAdb1fH4YSdaFnI/qBvJl5lHwsVVFzbrS+vlWJLo2PuKeTgrkHoVdcyUKs5mjlmCE8B4Swfqc
EzHCewQAQwjcHDq1jBKo/uthKESwkdCPV8uOi0pem8ZRy5VzWZpfN94ls0fZd7RdjfUZIFSycXFM
zLqOwYc+NpW0KRoRYwpBqgJRIw2PoOxObKsjtsqTB4Cq5QfvM4/u1B/UOafrszuZMZxZbkbF4Fis
UInQkkTUSMls/P+kWHjJpkDpxyjIhKQAP5g3QF+B0y5F6UAiAEbyNPWIhlNN7hRPOnDhlv0iW8jc
X7Ewo1g6VRC6ybdW1uYarKeXv9iHzQ52pajVrwWQA3RMsSPVfagdCVIOK4d9mq1rWK8Cw5NoqlYJ
kSeat20NQDax+AQZEBmkRBfZ6uibKyUJGW6ICsxJA+9VkawfX+kyZVGNhBB1MjIpI3WgZWnrc2Lq
+O+mnA8rTiJk5gkoytaRtuimBIVwKmRvq+2f7ii0RZ1Kv83jHKsYyNHzxUuYuU+17kLGgLwfcOj+
aA2LyRLM0aEuXpGOPdVLc/Ld+G0HpE4Y1dAt4hJi/8v4Dfg7IapGmIIr5CuxYqxusfVtG9J0ALBL
5dm5rxqJ/wUZ20/QFcn3TJRIrpXklZPuUJk2/EHdpasX+AJyeGIaSiEIn/opaFgEFI4W+8tVY0ST
8S0FI2NeOtWo62PZ+AMCZVJrD7IQyVRn1VCxRV2NtWENfKKOcMQITHyynSDhrZPgKKOycYj8RAr0
ohXwYTEvSK6bzWb5x2CoKQcP17FC54cAy9vG5WNF2LCC34Sfz1XmB2YmZiIRGADNbOw3lHrE6iyv
1agdQ9CENC30jmwh2m9CdegT0ScKfm7CMxN4xCQMA0h6FG1yAgOt5ZUAS2OPhuNuM6UZsFb3rMPR
dRRkjlcn9MmHJhMqpkDQuqPgJi+9+JmIULw6xoHoSHdZ+Sm6dEZVaoAhsQpTrDHH6Mjj75rJ6yzc
acLwPCYxMas7fr+ZSr0v/YtS/tOYDpBkkKPI0zWIKBBI2liwAlZ0
`protect end_protected

