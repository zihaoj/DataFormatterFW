

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
c9vsW5JBCvThyxOUH2PprRXrwDWuKZW/Q7qPv429HnbShw4Uk66yycd+J5tES7AzUCyGeanqADbi
t/NXtBFOdg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
THl1Z3bcMS4H5t6D0G+kJ/FC2Y9oXN8UuO5gTyqyx046tFrVCFbF7b10tz4zI+nryigVgXDuQjpn
REJa68sEKDIsGl5JYzOYVe9IZ30LgoXUIOey68bvuu3Fnu8lEQh/WChcCnbyekJTFEdRaUW6S2O+
5xce7Ha8Gv7YClnhp04=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KL9gEW9UR9bJ2V+rRImGqHBVYgwBOrGPetNJZ9L5EOgu04h1LECL47Zq26De2Obbv4OkIEGfGFbZ
muWpwFGMSP/qDDeS04mLx/tWX4SnYgQRVyk8AGGlepDKbn1R0w9YaYChqwaqdh3fMk+xJZbtgoWp
4ejGlCOtRuSFxFcOTPGLnPLr5saG0n7SH0iOlkdKRcxP8k1FnXr8kYqxu6g0r1ZNWNYlDcRB7pBC
lrlL52/HTgYUGboGp0/wpS3BU8yKiMyKpm/Nc0Q701u3QL3zraihgQqtTSzkLZnBFXKNrCd6K2Zb
gw1krcKarckcDY4W+Jw/vlWaBMsrX/8GffFxsQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
I9+ICDzIgzYMfdI9n5+7cSfa+M9K8Q9HlZVHvp38kWsb+jUXV67Oh07GXgNqpn7RlOPdQSyhyXf6
AZH+fL8ycTHV0MoCLtaJieiw5P4E1Pm7Fdq2uCENFjt8u7I2RH9/lcoRh4KurkxCVCe86Dtk1oWB
bacFgZX+QZ+FCZn+6nI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pyasIdA/E1o2abIoUkxhLYQwvp5B9zIwQEm/+EGPR3u06a5SPM2I1E62WIwSJ7iN/bqdRmd03/xZ
zjSCCiFFaRUwQmJJ5xZcUnw15IQqIRd/WQQ56gktCUx2rEJwJ4BBJrhOQsbLLnEDNgJUxpYVfXAy
ix6G1h7tonYt5pC9K8hh3YN8608V5TRujBAEsLi+3lAMFCMgjGqgS6cpljhaHIjuKULPnRb7+Rll
fIJqbRqDAQ0ubxbSrdH7w8ZIqWH5mG/hnLBefDFlIZJh/pHjOIOLGPh9RyUn99n5SKT8NF75l8Mj
ggHTuLkcPsoN2kGMWMDxZ752vU2X39SpzveZtA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6000)
`protect data_block
9OWoYQIn1vyMr8CK2vjbAIWk+4/2O9+5G7grOZewxUd4Kid6ZgN8vJ4zoqXw0vI9FrrcPWhOgRW5
QFAQfZ0ERJ07L1e6+++JdxDsIjK+ailB1XfZOjIQLwZyyYnjHyc31MZblTQo+ytSXJTvCc2sRtR0
oMaW3jKLlE6lUj5VGAcuR4+PYPXTmUSTN0M8ThOgpUKN/AIm4cigTVVLfbEZ2pKBfyDcSyOMEnVB
HjooQWZHBzX2P15BlhGggb5EA/PifSB+e9G5eoGgt/nega7lN49ayqrKlOhmUVBfKh2P69RULmla
dWHax9IcZHjjiJ4XLJ7+hlnDLGam4dbK7nQIsqyr1xS4p5z+/eDj3nk+eOmQcv3lWGMbYUtq6cKB
Z05XtrTgclx4NhTAWGz7gsnpmAIi6/QBBdWJrlRfpwgwRTOla1Ve2uDVQY9jJpY0uCBwho02jgt4
iFcJvUIuC6stSPgIQA6VteOEx9BAVwKhLflOURMCKb7yDtTqNn+aiRyEIukG7qYL2MC7+q/NNqE/
FuriUA+sUpiLpmmoj5XV9MwK6Q87wUInecrfT3TY97AxpeYpVyGXNb5YUWmF+6GbUwVpdQsuEjwC
w60JgTRIUg+xZ4U6l/56PruTrlXSw5a2TXfUczE3u9e9fQoScRAoY/U+F+atWAWFkLswu+660Njh
TyZWO57MwY2r1qwnJviO3L76NCpzJADNtHsnBlKPjiBP3VaVQMpYhnnqhlSWQ5Y36+UvY9G5Jbwv
8T6XlafVnz781n+FWTRzeco+GzOQkV2w8GJO8eBK2EoHlU4oxdvfjtvVwFlW2i0vCghVhMeYGb/r
0FI/5XQk3TdJe9q6vUaij/U2bMZwvp60YkPfqn4mE0i1fxEZAWBGEaY3dzALFu21h38LQexYSAwn
gau/xS2T9RNQsROGeIaaz30GgzXXMoNeVzMBuPNxe7G+SvzBSBPJOadHxKhwCZx/CuJXgA00xi7G
cnHEx6EJ2kLzojfy+Jaa2+dWu4OeyevvSb6hh3JvK1xkiSJdPquY0D/auUdDX8dTqSyKL8XTq1JE
QaXQ6mw8MnDr7kabX5mWVR43JscjjwPhGONEb4o2R4a52wUe2NLymkfEqdCJsCP9MPAVVBlmQOWR
KezZjO0JiYbe/9uQsaJpI9bgebYSUxcZQ3J6cG2Smngdy5ZWydZrz4YNHroMdZaKs7rs8AWOW1y1
sFcGhJWWH8ggQfVzRCUHZ+1hxFCSoEd/h1wuopPSO9nLE1l2PrO4Xf4gy/uSXrHheSMm83DFg0E0
qfn4jv/MQFvSecw/POpqy24A+wyZT4GtjwbY1Ej4XQAaBhMsBkv7STZF59DNLMN7Uamb+KWtlg9d
P57203ERJmO8r1ZYfY0scA+i/FieYgvL3KFm8uYixuLLcy0ksp+KJG7TFlfPLQSHrDoHWKFsMdgw
Z+J+OMyCOw7rXGWhwKg4yY0XLWeOkKpvS/XRpJemI/lZaJ7oJcWPWuHQSlUZUoa+HutTIpcSiy4R
SzND0MZJDK1pDw7/aLxOearKuidM+l5iKkutieAZ71Wil9bo96tiRFr0I8f+DR5pmoP6B9+PnTyF
46W1VhzuLE7iBw371ABnO/r+80c1Z/KBAs4wYg4fBM7MuPK1UVf22HanNNq0OrB94FtHFE0MIITK
23Hh4dbELnhVHuSk2BK+rZv7GPWyXH9IsD/B/24SecWsMO1NgCWuCUKj74hNnipQdCz6NPOrshuN
s0SbT+5Fg78xHvG1UQHAhRbgAxvMJ3eAJb1fssIp62z4S5OQ7gQubpjVVH34nAwvhweIC10Jlh9L
wnr5/eEqTTT2ZsVpXXVGMQgFyQ1Go/UmZsYbU6hPI9I+zZdf8ueCET4h6tbE5uWiwrU2hVwSr5Ga
2QZdace+5bRB8zorFY76NE30mVlV9Mp5KG+U81Fx2gZna5XuEVvTsBe2oT+wBdq9jukoFfKFWcGt
RuoIy6V0FJEs5QMCWjH+MUtpu1A5BtQRjzA5qyHl72qFA6fX2ai+2/yaP3408Cs+C9ze0O1AydmF
A6m4+oN0sAu4FesRX6toIDl0ffd+ptqzcBu3KKeojJFIW2P+XjTlLbruXK9RJj5mmrRx8/515XEj
lZdZhWUPAahRZNg95atxULdMLt9Y7IAaiMADNbYPOOXYg4R3Gb6Cybzg1qyofRucHJyHa4jIQuIz
KhDvtbt+Y0dRIvon8BN/KnkjblfpX6CILrOZu3xxDd1MfFX1iNJf42uxSvQUL+K/1+mu6fB6Gs6w
xc3QnkGXuGvo1AFx0Mlx+1oyC3ykFyJwFAhrFikESfZKAod1sBPh4aQvRbvammSH/Cdm4RYgJlEe
S6Y6SvxuNDeUXQVICxn7oHj/Koph3BS5MRguNe+TdEpSqYZMdrmoC2qrmeEfOV5heAb/LhR7pUi4
hBFkwb4Df1R/Be/tNOXmP59V3wrB37YHSZX5TRdXEbQIPxkgf8pn9IkvQ1zxpJGn8XLiV5GslPx1
Oa0hSoykmbdSmAELXIEGmB2YYeNaPaYtT6zRgm0ryIf/soUqn9l4kXGQtFSYTgaJt7cJs8mKn1/L
74XSJvAXBYXq+DPoUfPq8noEHq6pPGlbiXPzxF9xnsHZCf7VkqfxvPTVNJobka9CS4BMOgpZc/69
xczqJSLUQPyXeGFFSbDApWx/z42U/HCAxcOQiCwD2SHm4w4UAidwWNa/BGVd7+HbpwlcMigYTnvf
n5cb2Dx/FkyzVCat5PCDyx3KXXZT6dB0OCVsYLjJ3zzEOdlRJsPI8GFmcOYjF0cR6RbYfLOIW6EU
/peVLlYrJa7xHL3y2kYN6//DopNloO0KSgd0a171MqHyDAEDFMS2BkgiD+xqtD3WsHTVh4NFspiR
n4hjs1t1V8NI0pzVqryXQxBvYBlTb0h6f6kAzslUt+D/oPRqLKAQHkNkSzyMAwQMqXsTby2xW5v2
a7H6QeyV+F/UQrSseaOpWyVQx424WK8Nq+FUpCcnLPQ+3AxM8PELWThGLh3C5e90Xws9ry6Bz95Z
nVRdDXsBuMDUWwMCJu6Id2OnNZb1J3pD9BGHsiPLRlBsn39S2264ecVpZ6JTRG1pr2WDdGZLEw0E
rzigI40WqWv6y1vMkW6gvP0FXF3MRc4mGW22uilxWsUFuNBhRaZqcSFqDw9ie4nHHfExGg+egPtC
A31iwo1Ztiu4I7EP292/ZyHfDecb2UfvPsmw2vFi/uz4qVX6EYo0RfTS/w1E0sFKX6ySO45TB9dk
kCM78hJElJw33zzzZega7bJb54vPS4XV2QmGwudu1hehBTajGy6HCs04TXMKRZ7lNQGU8u4kE7B+
P4zT8k0QxUmqtDu74cfpnZVgPPaNN6xVm51EvVPpKLpg9gsvttv4hcrPViBaFfNm0X3lmjVnqzPx
QGtpwebXi+ne7O7iKShXOrORRwB+OeS6hJ38FxLUSAgyuhlil+uqYADkQZE7rX4qQyv0rx0IwyK4
v3ZExqRtJsegiy3IdTUBaYVXM2g+CC8gPyCDK63jTOYdcNnyp2a8ycOI9yQ7N5etIqTbzbHEFWJp
WpTxFn/ROj4vITaJCd4eK4FliOJZAw2mNdvA97XPLdhIoLQtYVAGZ31m68hdCD4Dz7gniZBf2JsZ
Pjbw8yumzYu9G/U8xUn9UojQwwBjop8G8ZITXqdVdwaqLSV0YI+k0Gub+McOkw3Yq4kIJfe6NcW+
3QZ5XLuCIYtYxEP/3nSxUjD888PFq1ehMpht3wJoIwstK6b7nb5YtxPhXBV8/52JpqxLrwSFySQY
brDt2cgQIXeD5/1LGxba0ThTmCyCaWx4rdgcblnMV559OblKrvIPoBTE2ul5E3kBuuN/lRGEQInE
7WrhOq3oY5exMUDBr/UNqSbTvexY74JelmR8abEL9fXqugNbh1tofdenXWIAWPF++7gb2SpZ1qu4
fN//kdjHxaVJazT57pPoYYebXeNMIcJS4ZdLifhWzA0adkJhun+BAK6lwMv1j95xyPREJhsLnImq
LTDko8WMd88RVIKMssj8AXoAJQ1ZmER+WGo1vpfzAZpcJy9sxwPX8giulidI72yNb0qOEHZ+/e3O
+0DKC2WI+jLviY+Tk/ehHofIm6Ufu+ALqVOM6/GiYTL+A0CLZbq5bm0zei0FTn7dlpl/DbyLO/Ej
EiexDGtLwWFe9pJk0AZmc9OaEiu+B0iBQgg9RHAfyFNyFetqvzH6VNWkSLmbSMwHPLDS2YDjjD+m
MmIvJRjgH0siyo7LYCN1/TXM7pPX08qZO0i9jzlXPE3GXAJkgyOJQM1yU+wUORetwYOvhTi1g35J
IWXasz9fhtXaZcQOUowm0pHqWqurX2hP3Swh4VULIpNXlN8umBpz/ZpJ74/IxdDdtcZ00ZlufC6U
qr5HwcNX8Qt9EiOOv0B9zVYP1tsxTDk2T+OPIhfe0FrlJxZ+IcaabnFYtrEkDiaKLKAEU3lZj5Ir
W/eELVVrIfbQdjvC/0x4Vz8KmDSTIbvCg+dlEuhCZzXLk9bu0UufBvPsZPwcviAItDWrNecCSDuY
9E0Mitjj1uqqlVGn24bn3f+kW5lFTYuVxr4LS8VeyuKlEFhel6gPbTTaah6sD3J2JAfXiiQIMh9y
qJv5sbGa5Tr8QLRFMg06rYA9bn932H5jwcIFZGIGk9Gg5Poczqf57iD85nk4kTpNcM/0OqGlvcj9
ZKSMTBLP2rJ+kK30CV8RJB3CrKZYEpGXTOhyvZH/FIqD3Ov/k/Ura7l8YaitTbQt62Wb3prd6tr9
m8hfyVvBWbgCuW3B5aBdAFYN95PdvrWrPzRREypl2xo6v58TlrQBvdN79wupETFKWnuUQaonL5yI
B67VNB9regFc+dw6b+PwXIEywVlSZJ2FanTlQ6XNm4U3ZbLJVqO4yVAx1I19IlOS6AWjX0MN2rBO
hNbuz8LzAIWkyeVHIFVNlzVD8PGtxKdjcK6DkRHRJ3IuKKbifs162vsQFOLuXId/JMG8o8nZ6/kU
IMtq0CFCT7Ba+MI8eE/OeLWJ196QtVTJTESrgvO9oW/551dl/pO12Axg5MYZEyD+CDk7LXPCWb4u
zIHp6zWTmkvYNoiCg5ivENLqItDjcstr0flUOKTrdjRd6QPxtpycrL0dRsjrl5b3rNbds3zAwUC+
aiT45TP5QuLTKF8s+YNlUW9MlV9rzg4zhBK4Ja6/I9UG6ffBeZFpfHSxTQOqI7eCYgjng8Ih4SCF
sjZFhBtaBBrRyQqLb44nK5aFdrSRmo02/VMLwjNxRU6uhSNKq4al38L8Kbwg1lypwCqK79ib73No
ieN/xEpC8OvlHjJclHN3cMRC+U0dvr5Mg4ov++5v2Gu1RQ+rj0o8+o/REjsota1UbilPWDAbOhKk
eg6wXJ+qptLuHkUyLSEn6mMvT8rvvwRA08v/v/fosNf0Nc9QnAB2oTSop1YeM3+cEBvI+zjYNZLu
g4EoK0SMB/YfMpssI8VOJE3115zkEq4ndT+eBMcL5sCmocGvv5xjGGBCvxPlgz6J8zv7r575IHMp
bXFwSFzOdvny7A36czE/91dsDSd5jNg7G16zAhaaTxE/0Uc/uGwZT7TUDjQsBudW5OJ8qIsYhjV1
xmBAF1pTSEV74Xas3Q1128CKlqKeD8Mll6eaXD2OhjTCGcJ9TzJEPKqOGRCaas0VkbQP32Qqr+Tt
mlv0erj9vIPJyJ2xjTPE9ui7JW9aWKNm+jJTdske2k0rNwrM42DuITlYhyYZVblRuZcATHOug7sK
rrI/WuesHW2aoZP/IgSCcPAASvOLb0+6F6RfUrBY/phE7up/ZrRe7dYSAzDvh7k9MBmAMDd+deKV
tJxo97m5MR3PQjQXCmy/2Bgcu8wFxMjGsc5CXBQwu9hJaeHqmBPjiaBpu/0Su9WQaSFBTz6Jo23+
xi1ge+P6DvUYI+S58ZVcejL/u1KGBS0PFnuWROWQF41mGCgQ2HtlRX5ttCIDwKj0WNYLLI10Pija
BqjOJFHDeyW7dKVxjDr/p5ZfDmfVXRgcwrIrwXqPuA5BAlEFlvIpu3+MFstlgYNiwSF8RMwlBjfQ
btd0tWNkRRyJ66X83fAj+E4rP5bKWrBnGya6B5E9+0Ah/LrjXGyor54Goan6K+XZysnW20e7ri6d
gnSSIGwQsXaWh/A/j7ZWDz94Q0VgFe0wEj+tLft+yZKzRR3P6+mPZdeR0KojDblKnPihl4F+LdTl
8OYHRO6nqh0oWpgBTsbbBJJuKKDyTxQu/f8o5nDHW0TUQvTK6ggNRwYXibwOSkWDY882k/C257vm
2Cs+06T63EM7PS3tU3keum45xKW1ttps/PH836lLXT+l5yf8/nwmVn7EazF7P1CgNxiHKr4oNUPS
8aFuDBY07JoMryd+GryyBxJJ7NsNR36iLhTPWJJXUkddPauGil3gYF4ri6ebxiY7BnaYkws6siqv
VDpLH+mAeZJBgltFpWZuixzMStBVwRAenAR1yLfKT6YWdrRdQE6IxFRVAfBQjAAxyws+O0qb5+5t
nZRGba9N8ba2qam6ODg/9i65XnxEEhZ/GeHggWKUYgf4+EX5wG37EysB9Bshde8kdRVNpjktI/W4
p2HEdzKPz1vRqHW7WorVEjab7BWXfvcyLNT9Yan0nkXnBqDiaYc7NfzV6cHOYrLtxH4ioSQ3/GLO
SvEaQA4Qf10kepJ6SspraUwScwUlTvm0kf9eKm0fxnBYhHCM9TD0kTao1vLfJFSbL39y8NnMjRbI
sMzlzIQPbMkF/dH7jSztdcfQfLJ/fAQ57TUgjTJ9g9YxBUEMXna4k2zsBXT2/xaCVJcfZ0RHIauz
B5yBwysc6//OcKkU5Z7qrYCQqWVvokAqAdT3I0veFKJkEJNLQEUGlahboyIJmenE0sbaBK9gkQSK
HOZItsybcuOyp/9UBjDf9i3KZ3tWInj0bmzyZIAkt7eMX6qtQ3Jg2GF2F5xZDt584x8/ZW+cmMxL
bDyCOqw7qf4T211AzFygktQmV0/psA9iAXVp5DQnxG9oz1fT2oYWTYF+PGCxc0lQraAhhTcBEZ1J
/lIYQFYaaW7/26ZTC6nRCK0P+8/Y8VplZ/7W28KN8bhDG37gdooLJysQCAxxThAJjEFUc9mg3u0w
KomkzE3uuK4Lewj+7+Eo91ywwB5fEL0ztXVun95qRQmFiwBeaPp2CH8GMG01ZMdgylU7XABuM2bA
yymnYZXT9wkdMQA+TcZ3YT5mymAdrfEHVxGGoH8xSX+8TzE7ELnkUe95cm4maQBSm5P83kKXUq4G
eg6mEY0Iq2LW8sNOkRv5Av36MhAflxjgq2MHcGYIkTyzEFReKhTASGZ0v9pKZZJTGhiNwLUBpLVo
ETHL5EhAthoXcv0f4Ng4rlTbiaJdO1ukNhuFmD1aY5FzEH1cybEVdoCR06pKNg1EUx2kNalclavW
qz8oSiIam5DbkPlI395mU7ypB3ACq34DDBc5wYVDtQZfvF3UiqOU4WGzK2m2UhlXVWynKX1K/hhb
xD8HRD5jkzc6DFBlKnMshm5tiabmCjis61k/YARWRpBwDdgWYtVmI9BCXJzltyPee6jvVmIdc8zl
vVEBOuZxe47IDMPKPkCWteoY+Dd2XJJzky61FR+2l6ds8aj83dR1ljRCna4nKLmeck8nP591yhbR
evdox2s9gEdvweNr3lBwFwPJpZV8YN61VD5wp5fWItioW3tEjD3isP3P+M+u8a4IuOyYPBKxlHKZ
lndioiC3tUU9KMjz04+y2hByeNwILzfhhseYpZ5Dz9nIqJnmmimGgK0sxD4LQPlNXW7jGQkxX6RB
TFsQVOK+a6SaKOjtF7h9HUI9TjLHrNXqTvFePwI7vXl0MNIadHiuvNejbnPCvhtuyhuAx5xq9/Ay
EzjBj9d1qosfNbgSi1/XTpxTXxSSjrib8B8+HapVb1Q93RoUAeGji3wzbQ+jM1ydZIaeYPBQoOkE
dOu9b1dk7Lvz2m2lgvtN
`protect end_protected

