

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
W00CmVavaE6xpJm+b6xK1oylsc3w9012G0NpEidmtkcnNf7sGxYvWk7hZZ/4udVcfLvZK+EwXddQ
Mb1PZ73EtQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Vg+m9KEq1D3Dj/VA/mHeuE6kqIzu1Rz586wlm6BjbXOI0was+kQj16EO1FpBfc+xCgA2kv8Vv/uO
2GuxrNbHFAH/bkB64EDnE9/zIVPVDjIHoCB3zI/pRm34b3HMUCUcP5BWmM/EgYYeAvOTUGm6JHhC
Tf/P+9Ef2oth8ALM+AI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KsSsCDq1QIl+O73zb+CIYhmCkNVRObSmEAGyyPq5fWQgZ6yxuwpPRFGmCXxXW5VLFnvTSrc4KIiq
ayzocbJpB/4bnUvuzNexfJ1boxln7QfN6A7LZPBahsghHAdfDmy8PA3IKDzmA+ZGuNX5D+DTzJOH
X4rtYWyvQfz8hsapx2NOxGGRgXRx0sFqOe6HLT6uuJJTqqoRGjiP+9MdrrqXJvlrg9dWS/IoThp3
bUKv0QodGBUMGfrArkAVQm2a+7Bb/Gx4Jyklwkahx3DxqPvj/ROjvefPz6fAD6FZqV+mcQCaeyRQ
XhEFoFLDHFG7WeZRC1h40sCf0Qod+lqTZ0I4wA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xu6mK82nJVHrDrsBncEkjFSr+C55lIRrJGrQqCRg1sh/afc/8tRMRP8v/RPTMMwluFinLaAbVyJA
qbrlZVcgPaCR9FKt90y93ok74hdhuXjw0+W6i11yQGaysoPjM+10KhEb8JoNC7mDCyu8/zl/NQyl
lOBuZbsX7GpuLWh1lZg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
p5Iixc6t1ooHurr5J4hbaaASc/tYEDZVcIxYVPtPuNc78QswHhpRBdGw3kLlcylpeH2LcvR72QdC
f227apjhBAaQ5YZ6HTEhpb+/d4ZXgkP2ZEfOkGED+x+Pgd6+OudFO0jA5rr+QFsTSb33sXixawEO
GHNFNwmdeNloXriotEE/ZYrwgQzG9VROLCTiEBlMw7lKUAY3toERtBy68/Vd96my53C4LuGk8LOK
oGpGa7lxXVlEuceoUHnfkIH8J2kZk9uo875ERmVNG61SnVWFmUETSJneGqyXQfX7E0/2GVODoU+Y
VTAgs4liRaB5+DBDSIm72W6jVcYctnd7gQs9NA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3632)
`protect data_block
blz0Tmdmn/eNI3jxGqrCqLWiMP3kHjMxzuc3AmBO+sStoyMcyTKjmOX0rwFMAylhbQE7AyKqkDoQ
bx58eowmV5L2suDjvsMfhWhC48Sibsz+ayVWWyHV8qh4ZJIc4C6htSuvGYlNnupmeYfCo0eFLq0a
p71l9RMDPUYXlHORzahdTVyjKYUjuQJUYMF4LAK10TyRM9gTHiUEATTQkKjrRiULtlsvog9LqlHJ
RswwpbRa4RkQvKHs9+WHi2VCGJtKcc1mVimhWIgwoCGZo2PiCOsnZaPbjS6q0x0Evzgchk/BMLZz
5BD40gTIovEp7VtpBr7AwcKjC11ji2lbK7MaenAuwFCSsjL8xiyUdTGqnFbbvhHVvuNjUiT5nFYV
ctKNrGr5lz8w7JdptOIZIaYoSANHvV5kzPlqf+/z0OoXhaoFKXzS9SVX10Vg9CB1cKVyCckP/vjt
nY1hUn+Fn2y8ZmxeLO1YO391NaEVvc+1witScBPrVathFmcStj8SKPggLtfuzaD3q3GCfNGzQ+PD
ugFF7AQ1Rm/OlCeH6SetfkbyKjHaYD3Qf9G3kkbClMGs5ZjeG3Jb1Urv8phtg+OzqVuc/N/R1xa+
lCqRJRnJVghC3dac3PAiDHN79mUrszvOjbws6Y2ELthAYb+cYEUxFLnHC6Z2X8FqLmAC/56uhJJO
0QSTJ9m0EUqoir0ro06KUKlKs4a9rjCoREbXx/is5E3KCPs6eG6kkRJp8r4B+FnIptubdaIg8ngT
9B3kVvVOyLPaFiRvhcPGKbFAN9epYTrlDC//MtNAEFz/Y8Qmo8IRL7VoDoO01IOmlgsf1gGEPQl2
faflilJCxiS1eG7IMvHvIVn0bVSBNTdFoF54uaEZHi1lsYmTNTAnGi9PFgFPS0/+WTH2Ts8OwSdi
+XjPdcg9mbIYTlRGHWxOJ9Cj1m1Q2GRQbc/IbdEadHh7SdTBZfm7Yo/+HVtPlz3eW49QQ+uF+3l3
ZovKq3YeHxceWRq3S83t1a5N28cvfzcchWm5ohkGTiGtCIfCxL+uv3g3rmceRlb47jXVnuC+aE5Y
4yfyyW4HcBiLav2pUFgBAtmUtLn4C87xazFTnvTzsJ/CcEritrcH75ed8Ue1+6dXCxwXVRfDQoUH
0idqMhIxYWwyVWWWXF955rC9bLHZXeav35MlDcckiC8Ih0L+Mys2i8ZBCokZiiWEWnOtYuXXMO60
dWq8MLZ0MH2/lZuBWzJoU8fWHlk7KHy6jw/G5ws/QA/J0XqEoWr8cVi0hUcqtuK1lplSsCZ8Icl+
uIrXAPGfQqoxOa0CvfoU82nftvVYmBUqpemtLXxmHfAZK59661xX515yYpA5xjRPy2amCudpivMu
TthC48bGtdRddk/XnQa1YeWyaxNtDheCpuzaeR8mPqMON0j0FAUehyfz/uFsSKBoTBbiypgnIAT1
PFPcTbJY+STt7YrfxvmSARkeCDYug4Y6JOjYYF9poVcRaL5n9etpw41g/e5ibMMudwsQ7SQQJuWN
JBnnOjp8xP/4mkYj23phEc85iWuDjAalRR9fz1o0HkJbcWUe4bbSiVrwiKM/t/+0yqoFhlbU12Jp
ctDtMLaWXTmptgYd04jHa8ehEUWXXX5IQ5Cc+7v0Eyw6xoaQW6NX7PlJ9AXN7gzcshSmjOuMh+sq
fUs28+C6mbQNoGckn7SKTNexjYziZ4WpbBGk2bdXbYk4vxg/xFWMO60twGrtZ0AXnHqt7rTG6sLF
sySPEGQ66IzsPbAE+oF0r6B6Ad1Id0OV0UdjGKO0psEh+HM5qMcRDOQqnDueqhIDlL9GEqCnZzz3
ox0IdQ4Z1Gc0HQ8ZYMCfRvcyKzl/TXLc2REk1h8GSuuz+EU0teEuDoOud6EnNwKqoSGExxXM4WCx
3wuZtBTOEXcxjZTWiM4vnVUSJznKxRmiDVesSd/rVVPG8WQOY80uW7EhLOfdxX3iQlQok5QvVs2f
QuMFaslXBRaEIBP5N1hgDHf8qesysBVf2u0vy1Vt64ehGmfyd/T0eKW9F0v0Gfhk8aX/XAGYp147
U9DUVhsSEmpGdHdzYmnIfLhRhme6CprXvqj7P6PoMZy6KqMXEtEr2G0w7vvTNzl1Ij/H9KVJQxp3
RwHRFk/6o+Us6XaK8kIBGr3EumXw/dvcn9r0mP1uXDRNgcxq3odhHq7jolWIBTi0Iri0OkFev5q2
LCqrPKJSHvC2ztrM1/IFbN7lB06/gmrxMDjbJW0LLEelpT/2GpQMWSPAeiuW1im23yKyRVMmGC7w
S+nANG4Dkx/vcj1JE8voLItXb/KGIwF5e7YXoMpM+Q43rKjMAXep9YoJFgFCOhenN4Ouw0JS7ybR
I6Aw97/1d8FbkEVsLVCvGougVw6OTvby1pIyChyJ5Znzsf3/shM0wi7WpJ6y7i+9y87YljzQ9alE
f0wVYEqI22pu8p3pLKQdmBSd32qaq0ZxwrJp8BfpvKtIbPJmBB7nOHb64k4A7E7D3EbgD6lYFSae
wgNu6OdZDmVSoN3+X9HNmXGQMIwzCgN8JwLuSwq8oarMQtju6x2EtVKQxUyuU+I04pVrruvvMxPH
HI8EDqpySxE4Vb4qFibcjjJwERAZOccXmSHei5wpUwVD3x+DVZNN/T7iIsbR36hdcNj2BPY34EQy
pHV9iu16ZhDmuH5U2BoAA3kHEXen1Z6EBIe+FjTzFFDwBxBo9juuhkPrpaJU8A6m7xvUD98/HeTs
jWyDRwSKUPbhovMDkP0Wjh4KnLgJZEM2DtUGjsq0KZbczG2JuwUuVMapEIRq55f2g1zToSMgwhZI
dd9KSU5+zaYllmeOHca2+DZjg/7a99m/nlqMubU3WnIou0xQz/7FMB2FzQ02L0hdeqZWd1XPt3Ry
dNXYNXwAjtCi6vB7oMNsMj1D1ocFnYZbxIOiZyawJhT148nqVV+ddevQ7dPzGs6APhSqF5uNPooy
EWfauoq1BJ1YHYCuLj18Mdu8ThfjqiOgGWUqYgw3zYQ9h5C4gOKlZzTTr5E1aDVjvn0ti2gMoyN1
DdAFrCs/bwE/zF+Q4Dg7gbpx6dbVaoRPTXa38b313oX2KM25czi8HEp0QB5K+dnrX6FxhegI6TLG
8wEJ1hp6oLkPDz7cot3IkxTW5m9jXNN+iJMF9YKnC49AA0Rd7YmZF+dhX6xrrVYK0caxrBHESFFO
xlzm8C4DvH1DZxl4QqbST3ij8mloJ9Q0BPvxEjbeCmoR4cPMQN1TTtjOOJhY5nqLPig4FSag9DEB
KJlihfRbyquA72vDyJJ+BAvomxDHb1sfq8m0Tj/Ll5JMbIoLO4iE+7eQME6SOcAnIP3rk3+phHw+
8fKD1s6jU5x+YK3praqSOiE29TWkwt1ml7eV6XqxM3lj/TQrpNiAdblmuMHfBmrgWHmCUEHNZAUR
EoERah5pZYvenvpTp5p8EwuobCG/Of7RGdfX8BaavMYBRfZ06fQJBpNYAG/yxuHasW9wrP9OMOx8
5KXahfLr3H2NACXOYS/ad3g3kwmeDzzawzExuwIrLyuA0MQOCziy1rS9js0fhsiNYjjn3dp0SZU9
4uWiYjA0AwJE7xDg0A+TEe4URwjyJUwIgGnyspvhCr0puG61WyS0rMBc2BZznJHsKeGmjlVLq1Mz
LQcbrHCHlxh0YZwi8hPmaTNx5BB9qCm4GRZ74PE/bD0x5yqeQ2rsS/hrz1rJmxerSUlnnZ0SVv6p
xF2szkQVZNOkgDgh6NnMJ/rqNdz3V6eTCgEmQjaLsjpHOuKaesRia9ZxBsYiiQCytDpOG8oTPASr
wYlc7rH6DiOyAcxl+G7Hvc2UoMWM6vu+RAKWUYe3guudamlSiRu1sfRBg6UWDtaOjOAoufVc4vYc
k0PvoyJZm0JTCRHjzgUOtvnPbvAS4UGMk+GE2URH5njcKQL8XELsvzmkNKKoT5kihSbzWWIGLD+Z
iuj2pPCpnZ4+uBrU80Xg/ORnBCnrehhzL8IPxRU+0RiIO54BiSz7x5/XBG+2y6iM172YQpVicigI
a9zeipiffDaYeFPR4bJh1/C39Eig6JgdXIrfoIf22lDAmGnE/3dazYwoKP4r3scrlVsfZwJb//Ks
HWjJCxlkWUFqEZuxEZInI1nL90I2gc9s3Cl2oa4SOlfXpXBYiYm8f5b9Jmyj8Oi+i0nXMKZORys6
UgexiHBgqm8INgUpK3VT8Yi979aKJ5gmo9++PHr0PRQpXELsxqvLTfkS3HEyinu2lnMzeXUma2fi
Smln45x5+d3EHXg34ZzCve/soJDDnMZwmPuiD0/ecBCD9rFhMTxS2dIYzvjW5pE0xHi+ld7Jpy+H
bFBhZKddUIKaQNb5F1G+wsRugcR3ZyXumd1FptvB4xR/TZXrSDuVfe1YYv7zL15inWIUhGLNl0tF
/Fj/PSZ+CmsHYFNql0o1zZFXr9e7PKj5rILdh+W5+RNBaboNtNTSwCox+XVB/CFzC86T+5DwBlD5
A4ICvZsNJAO1RfH878AbyooukJMUsmqKRKit1yCJdOrfvq9vFsaGPfL24FxHJHb/T1VWACo0mLEE
cFf/0nCucUoZBngPTgT9fC26RJwwsaWfe+goPViF3vbGJBlqpj85Hm1K1GQcHmsJ//shvYoegTRh
roh5YHtqhFMbQG6QwK384Sgij9a4WwxZGDjUbf5jYHmoU+wEnA0Im0sTvbaB+qz+Hmw1CBcVjdQz
UkKjqTKmoWxAhO+re1CIF8v1coOcaDuPSzrTUwvjGNwkfD8mEUGtV1QFDfHu0vhSqV6k7Vn3Cm0O
JC+W7m4+oH6CDnGDZgEEjKk898BuktmW/RyZYfjT4av7eRPBt++xQXA=
`protect end_protected

