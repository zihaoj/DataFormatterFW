

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lVwgf0Q1kLQjSR9WF5B6LMTziO4TxeRSiKHlF8IWhO0EALXv8K4k6dhyce2rpTWfPphqqiSAfxcQ
Jruuym4gJg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a6j8Mmj4cjJiKRJuQyVsLw+99gW3x2Bw3C68+j1OG/liAKFZkv3fupLUrCztIhjyGAQpoMwJq2HC
pmOjgfDv7i79WYv6TiwCgAxnexEcpq7Sv90AX1dqKbdB9fprwKBOLCP0uDEHyQJNiRV+PvSLtl0/
oIqfgRvOlln1V2+FHJ4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BNU0DSDiDry+Xzfeag1vdccODeBiun6zc3BG6iQ8xpEuyyQDlLt5mPvrYbJ5oV09DFmlMV9eFBG9
u2M628ZpwwPHB3IF8+65xpE267cz6kFMbNdKR+VcwDb8f/qepmxpCMAJKW2wxfVFeZpgV/6mg/wE
blI297kGSSYkoehXok5he/Orp0C2Wu8/2neZn9aVeBIsDLL8SqQT8jUj6KNRvY2pK5EyLuJU4ck2
8j09tGHYw3nXCx47QjJWxTgThcStrg+GR1idxRsAHcK2nDqBsuD3KTjml6rN+HGjf6H5918BS/NA
yy9Sf3oljG1sQ2IRKt5tbpZO+dHmuZjg5pbdSA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ypry9ApTiilqkQLYX3p/6ox6OVURG1kcd+spGUsA4iff/ExchqGs5aErFUqFIuBge9UKQ/637tfI
4LRe6qbS95zsyVjhIw/zYXX9JZnTH6+AOX0QyvONPDXpPIrrksq4M26dMGU/61MQ/8+NjGhxahU2
6TsZL20MooGzrhq2JhE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XQPUyKcx1D34j3bdAqnMpdeadEOKznh4svbZ3n22Ivvc1MR5nRYr5ZyNtBJ3hA8BG1c4EmBF+6pr
nwPhnw9Cm6KNofXrsaWff2kHyLc9XplTa1dAXqKnTOPId9K2weq1Cnh7CD7xyMw56GmPO2E8BcIr
GyHxHrJgYOp96Yd/Hkp9HGJN6L35pRegT7bY0bdGW2lRIAzBkb2yzW3RPxN5aRTj/DJOPaP8dlNt
nOdXm4qzNsTV+A9lt+GONf/Z/KomSDSj11gBX+K0qtZKRSWj9yJnT2w4n/kbAm0928JjkKVsct0c
LYgZbHMko2bhdEA5q7Ui43lR95Jlm6gtXxGIfA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54512)
`protect data_block
AWGFGB+muu45gO54e7QX2CyR69Hjp3U4fTpamMzXyFhWCDT8t0ngLYtlbafHGl5LmEss+Z/KXNCN
K5kfj2s5t880mpUmsMDZqhG70hZzYLVN/xilPMpkfJfzNZp6UqSkSKrcTol8QNgG5tfJYX54eaeT
kHMlWFq7wIZU2/J9ZfXNzRhMiFFaRQsR4twAK15iJgNaF7+SIri9+PrhEG8E6PqjcfZQlWnlxi8Z
AAVjNHngmwwc6oKY0IJ/Wi1z/ml2ahRp7TWBg4qeAdTl+uEh8WC2ZxFsEseYJwRl5j+tvpzN8s+b
YFJMv+QBvOCbABo6+WOdxbu4x6FRWqk8BwBOxCfetuEzkEP1X/So9kLIXzqs6BzU9efCoHncVyMC
vJfPAeGeIXo+BDSH3/NE0LEh8D/SCZosLO0jIVMOBQ2qDHS0FtO594jrpKpF4aKkvUW6JXW79Zmy
3nMBacQeFGCaBAyKiqMVPDVTb6nmI5I1RUYvqIbr/T2JTeJLFTn8ZBhhPdKLvTnMBHWfBeRsIGMe
EuCCAvgm/F/jKW4Egqs2pw/3sK7ueylr+jLaRYG8SE+61zfQi8ORjUA6zNw5RTxc9V9kJLb0C5+D
/F/bmszgThnw4MydW6q5lWHwPAxCV09c4Y2zmPzIEzWgvBg7hhluu7y5RzaoBpfU9VXlDuFr0zgF
UMeYz/xf3CWUcDYrXoe8nWY8LbA2f3GKSljNkd+LEF/T72uiVSZpuH4hFWl7Z+s3Y4MIdMxvsaMx
ShnckKrphYhape5ghVlt9JuVWBkYkhpevSmaMVqCfbLwA7lvdPPljLJ7Pna3ysCI7PBBvsw36w/H
LuOHCxq/VWvZssRzOD/eNgx2AKMkHkiDw3wFMFXqn5HGP7L+U+mRy4Ad+PhVw7ryF37w3URFlkzK
MtWh2eqaFzKhV/QgH9Rw+VjyfMPav2m1iEuK2yzbwl+r3fxq9wK6uYhXfnl4Y6TlqFoNtLNmy0vs
oIqtkCCgFxEEtC+cJpGrju96b3hPeDb/l7rPY0c9yCW11Y48Cvk6QXvJ+uRFviLrHP/XQDQdOpgc
qO+6RL3tYZWPV+e2UDVBXZ9x0tWlWncwYHp3DVCR6MAHiJbJImKaqyTW5nZp+b0D6Cixkf0+w57d
QgQ/14HpClvLlF1/uAHEq3uqtDQGOfEl0BW7/BEB4173a+hgCuDnKE4TIHoLukKcXYdM/VC2HLMC
qiX5oCkx7lFIMVEsFHNv5oqlM4BBAsyXFjsW91OFcb31rsWoc3Ag/AJ7Z3BFC417Ajgsb6GmMkH1
zxYThDt3iZl3c7+fVTYp4jI6BbOdKMGKAx4mhxcwreXgbKgEuqk17IMrLq98WxhPoH1Jx8pb9dEE
h6ibEJNC3C5A7oCaU1oaTs3GvBj26WLSWgTEA1bIIL1JX6TZsM6ZxF4sXouCSux5kUVPbUm6KvPq
pK7HA9a/aH5WqFuJP3AZITP97pnd1xOdvI14emEVRoZZs17J+ZWk2PVma/qkKZBMRaH2gsWhaYdd
svmcJcLr6jDtVDXAO1z80u5mi5w88eQIRIE1Wm3wd+65Q86f79jGkrhPgkV9BaKxbE4eSZ3N5cbY
LF1GT+g4Qaz/s6otVb80bfTWpLPAgmw0T1A9/N+pnQ0GUwASVV3D/r41sBemuIcPteOf+sxVcs8x
MP6GZdsZFg71GII4bhDE9Fcajz3L74QXN9eA8HborUj6/QMjuhcZ9aEhhJJdrcgW15sWMwaosTul
FnVyEoBBWL8HLifiiGJ4kTd1YE9uIzWnmDMHbBataUCStfKB+2zLWq5Qw1GP0pwscxWrE+lxDK5v
uPToheu5r2mB4j+gxX3JF3IIvr50HifyC/m39YH6h8j3jqOpchXsYsZ3RakSYNrDLNEAwcZmaEQb
/vg51o5921gysoU3wNCY1azyVAGTN0GvmczrZ3ZOJmJA9B3mxV7QkatWCDSILu68RcXndVlDcDZ4
/1koKB8aQ7Ab9mqUeJcH6RKmePnVVAfM2JCXDB9oDE+8GGM5czSI0CYKd3o8eL8+cVIbuhD9riV9
DWKJnGwrzMu4EHuIwOON+9KVFWML5k1ktsFjjDecmHTtvQ+Rz/H3ecfOa2/DDk2PPpRstV1Sl5C7
M8PBwLZW5KthUhiemYK/n53tiW0Hm6CbZ6pqK+RmyluVg8oX7r4o1999brg/Vvhn3mlH1pPbfls9
VUWPi5kqExZX0QV5WlsAULMPq6bjJMOOKEVG3hSvZpq0PHH//7/rQWLoeaiRoM/E9z/eRmUskYKr
X5Pjqxr3aao+JZy8c/loyR8Q/O+i8Tbj36EMgchRPDN5tmIlsut2UKmei9M5LE2KcNp88pix/5H5
gGqB08CfNiaWVvtO6AQctrE5cV43BvNXffPXS+UY99qr5hoWFLgZr/9Tes1AEf7OTVd9ilWmNXK/
O99aTi6AG5vWgrc/kVuYzIRM1VjTJGeWmk6K/DwGXCco17BQQZ9qmELDO/xtd+6fT4UubVWqzPQO
1C9ka496/wRvj1srFEZaZtGuOMX21iaDrnirGl9BI28eSAjAshprjrR3KOZu0g0l4Trhpj4chj2o
gp0ssxMaCl/7SQuCg6DTBVq0z8G3ZZiGihNifsZjMbHbrX7VLM932F502JX4ESSd1ECe5RjZ/OUY
swG8iAkwqn9ikQ8erlbBvX9zdKo/6yD5wJgt8uZgFrS7HWRqpvCLqE4kFIIYLueOfCF+jFx3CUjp
TnXSTaab5YQuuU1dOZDGWGL9GG7bvZmczKXV/wQhTkRerjUnmdOyFqTtT2Ad+RPHMk1xNEBsVrtI
R0cXMVUPI0HUfrKCxzCPdXOCWsnkLY7mLnwEqxN6pDd67lYd5GYDM0HcUqeEZdZo/s72eiFs5K6G
5QUQ7liSjrLTCpCpkaumHQg8XozRcyw+N8GXAGIbeQFQzekYFSgMGoCh2Wq7MhS3sMqsJ8Y5Wb9h
Pl0EWTuuvygjYiwohLS766Czs2IvoQlnSlyyK1nXwWv9V4593oIeby9YTnsYsypbPAwAFkMZ7VFH
KEUVzE/nuBB79c9Dm9QJS/wiNfAE0OIgXiK5y3QtO0DoYoi3DgH4uHoR1eqOaUTywgk9jCeZ9VG+
nyidlQe1uUk61a4W3hV4iOuIG9jNsr7K8XqJeRwBUeO1JDtn80JvHj0pULs/BDbw7ND+cWn2iDhs
XXbyfH9QeQSpLrzp0+5q1GqWlkyHyN5jh4wTA8aT63uTGtnoDOLY6xh14I15040UM5xtmqKbVQUV
x0PC68tcXSK0iH34xxAiTRKWxvWkjxIj6EhSziisTgPjnsZAHhA+AXddm/aggVb+b3bPWDGR/5It
KiK813Jd2omTvpKdYP0H3Sh+rJaMvQxTFnEUOMGRh959eDbMq3isB282iCSJlXKS5Ix1hez0wfWs
wUa9Pep2yfIfqbE2iOriyEdHnZTH45O/EWdWHlWOOy3KY0IlcMohfOLqVjO/7XlsLgBesgSqNxDh
sJDhzbCpKkCmPNmDPuUncIgElqdJCh14h8Pcror+hBCjykKhgFHl3intdJSVRo1KGFQ/WuW+apPA
IfpkSMpRIxB5D6fUy0eQ9zC0jMc1+FcsnB3wTqYBQPyIJYEiC5Ms3wQ4m/PhUy2bW4mAe0AAgPbn
O7GDlqnNdFyOXNT2wrNoPxTKAcuaBLeMKkuDKnL3aQvuSxJOjrvMTOsZASuflCBQFP64S+m7FUWD
RSEPMC0EgwV7yT3BN+mhFQTlXyqzH9VHiPIGrt3loUAf/IoxzUPEHxdJMgIhvvMj7L04cScjcvyX
vcylrjOF1i+IznoXWJNJvIopxTnEHqH3UCzmGVGOP5+EtmDrVTRBw08eZmj4YGAf8o/4myphlUdv
XsBqamGpM62Vv3dttM+ASC0o3F0D/jd8uQYPX+WPdKD2VDgrUmpEVDs7jh2NrDo7AxX9p5Z00iCa
dvI5GbCsjjme+r8Kn0PkvYRaMLguSxREvk+tAplmAXLzMlXh+D6BPqGInlU5KFMU/z1H97JynSUd
RjfoF+VuxKsYVBaQRXURhDEPANWnPiiDW6onFMnbiZQE3zBQP2Hb+EmZg1BdpyJmRmWrN7rQtBwo
fptfHe7yrfkcbjiJT0Z33EpzfzM2d/5J89pahMvi5PETUwT1LM40zSOX+YbuKE9eHG+3zA0ggqZi
oI/pH3veDlCFbcv3kd7sTd/fInb2mTHR/uITIXSduCCvzRxO8IrZVTclN+lRnQqaYhXQt1oqsPHT
2k5woFV/gygZLwJx7NMPpXz9NSeVErsw19S+88MhOkJq1L1LG8RGQX6W9n4/js+rvOqeofw0yGlM
9gQTQa1pgMwaUwR36KJx7/Oador/ZB+5dPykQ1YBZSjf22jepAXCgW/fhDnSPdwRNuvCRzOKPWOC
JXckyCSAM8m+h5PmHXHSVpo5WRqWKpMLs34a5sQIZxZAlk0iUOi58NbN82R3AlYgkuUa38uQuT1G
D19eook1KPC8OjyCVwUEScmGJKOPwEB+vNrDHzX4F0eGAEvmJW/mpavtUpo+S6SOPi+dtkLI2dXE
kvJWdInNw6lj7y+OU8O//FamOxaBuDGxDnaavPxlmGOZOIvCWroQmzJzZ+RcOdkR0R5vLIsNtGsl
Nn8Tymhd4/kFvONBsK0hKGzX4wbqBphd+5fV6KEBveNpyY0yq4QONOOaK3Ok2iq0B+c4u8FeUFG+
A77d/AJ35n8t/vUYxKgJHL60Ue6m+0vQ/e86Iuc87RGlGJkvZNKqaXcEbZBXC46K5BnFAkumBIWU
OsmlAD9HfkiOoHbi9xtI8tDv2ytFiAnw1haP/1IoBNTMityqDx+A96MFgAPPwpmYRHD+OLCg86ZC
CZBw3ZZC4G6R3paa745X+OvgIP2Sd8xMS5IGg38NKh79SUdVjNWa1qdB9fSVhWzHTpjcX4XkRCnp
ojIaZUzt9UfhUsKyMnTmDhWJrYkxtmVmUB5ujggB8c0n1Ci6bIhfMc1tzPahfS7QHUCtMer8zurw
kPXmMZ3gAfhVGP0O0MWCcoxR6/Ey+TD8T38eEUi33f3FaBogOGuQGaHEPzhCqWTkeyOKgyTSrLzz
Wc6wwIR0rlEM9NTewaTEzXDbmtjSoB1Z8vNqGGoQ9NK8yIgagC87ugprAm5RrkcpSqnK7UP2B9B7
QLA71ZF/1wuvxdH+hVtmTy+hjZJbqZanI64J7vuIY1oKYT0I5R0BcL47+WDduK6AvWpzvwykWbW6
BaEqYpoV9gEHmabMofEswPX3FE4jTQSXq9XcL7jHHoFQuSXa/HcELp0jMLbErz8nUNBbwCUmpljh
MYyO4c4daGkOZtUuJ6ciuhL6G+PK1FmISJ3rIffR88YJlV5ZGqVEr8dMb+vcFOS8GC9Ao0ySw0aI
w8O7mrhnxGxX6B8hfZNTY8/9l/Y4+o0v2QBvlStMH4ShpsadG5xbHhBK3sQhBXwppX1krMU8F7eU
wJbNZuNhTrGC7EBbQjmabVKgG6E0VogiNs4KZkcBZVfVVIS7fSuJYV+vnF0huG5Aj/IVJ4+atw7O
8E1lYEUCFji9Uk1fTN4uwZj+Ojc2Ok6jywy4jBh8dszkMq5776LkJeSLNAdXS4boDuVdweeIa0op
KCTldgEVJLtop137asjPrJnTLTHSagJlboAu/xqheXFMac6Yu49Z136jAtHKHMs27LHBTlPahuuO
7QwgyvT90I6KIpuGqDdtx0yRu3E34lpGGjd1xZOkjpPpzGDwvIUdINdEkSyODiPKa0FfaJx2JrD4
ORG3WUOIpBX9G5n2mnlSk4oix7rWYCRXFEgOyTVLWGMfVAFZgT/gZaK1v0MCZUrJpOpGSFRd+uXM
mYb3XDtw4yD7r+C7G8KMS/gAIw5l+INZ3BceZvpHAcOTwCfM5G2vbnbPVjKF3j2LzhzgxmGFx2BO
O7uZy999AhVne9ji2l9fyw50HeHJrIm2B3GkbxGOPfwyhXeMjyLWbvNQLt7vmUJIXaUMKa62/Fvf
40bjtbSMQgLmi5m0PM2qA3wmWglbu8vLZb1Zv+vOks8vKchsU9VXjzAV+at1phu0936rV3HUQBGr
1RPUFENrSWAEHzK7pNBHR0+ztDEEHkNH4yfV3YnULDJ6iQ7MvYco0N+lUoAKpBDrnn+NaCZrDe3h
7NWrUk8xqcBGA2mDj3FC1g1tn1VSB/NAmE5mRUIDurjPbRycP5TCl8KJBcAIeict0OGS5/DgfqAE
/SdKW21seZKduWNjQJpNFxuuYrTi06w+/JaW6lWkYyfoZSRVzdOSfSfglnXypbdi/ZgSE5BKPrFg
MH10pLERJT5Vjiu6THnYn/6cjtj7B/NB2NucBdzA6nvhaDybZjMx7WbbIfMCdPtfJI0rQTVNLB6O
YV+dsK51oXyKIIFe2XrAEKpQW6/QO63D6T+dGGoTjV5dOHZjR1AlyqeC8Lb3EjSd3ZZx7b4oTDM7
29HcUtf/WlMLEhrNOTOUE9j8rmEFSoNaeSnKF7DnZX9wfJR4xeFBuNyMOWc6SssZVdIC3ylJ8ct5
nKsUSfoK/UM3PzoxcF4Cfh0O345rY07fsE0tZHOdrlTKYSOENKCxvrp1fl4jlzJLy2czIMtCahdx
G/EcDDN5e9Mhb/Yb8vAKY3lufcSW69sjVb1RSTe4/XQWHftg+3Yo5DfmGQPDS6yCYy4SDJcbh5N4
oyhoPLrXMsm/K1S6AsmIiSukeTVUKNVIdfqZ4ZvqiMa6zzKjK2dwXvXuabb8pRJaTaO+rYH64/2Z
4fqO6URbK1x8KmxDanLH9Tg9nzNhPNvtDfza8dd2oEyC3JTswVczhLJq3Zw02+housIAlz67DpWn
95waRrgOiiiTpJYp1oRRniEcGDYRinRHhe/nHe+DjMe/itZYLFws6gOhFIQNrRPfzfjncVpwGgWD
9Weh+e1CBXxIHkzsdzWg/n8CP00XEcJPbP/swIbKYly/bKv3xbkhSRk41YyiCOh+twh1iZODJVFr
cJ4RY4u5cULnnSr8mO6Hp7Aq/hmwOdfXN8/1ReiVr3hgXHMnnEtmaFP2UUFT+AY0owlMOT42rWHu
DXV+40kM3XxRT31cRfpg8ZIyNEScU+lsHYeb34KMIBY5hVq/Uz0HwCv712sNhUC+mZakCYucWWkQ
qYauTwAEU19EEPbU1kJF0CuCMVaKPuZAI0mvZomMiVYhq2lNuRPbBeedEuBFrBb46eWMlyrJe6ku
QMkmRq63M09fiOppXisIAt5bcw5/P1Gb9w4v7AJ0B0/bHz9yxP5dsWwJAo+OE/3oJl0Lsx0IzlAt
yW9q93ZHAxs+z9zzlie/PMMOEWDcgg2aYxrD4kaMYZmi4CmGhXcdacPqXX6uomt/fsJxVCpDcP4u
EZ59S9ac/QzvbXO6BNyJcWwCxtuBCxV4kz/o3GqqJkv8GERHLcv0b3EZWUfJ4nA9uOnIvjE2xwnM
+vseS0ZqdTDi59nZ7m+GhQGhk0oh80JQ5qE9zlVDT+GzSEKtfUHjUuUeSiUb818EqbcwueADrjHS
v0wZdV5xbZrGpBB3Jb1SLEdfUS2sfzGqIEN42Z/2tnderOsDiu2aGSmjyCCEYgwtlDtwPr9nIHeI
qhO37LlFbGelQblwYlASIMLbDnj8IdOGMdf/i0zk+JmY4qup7D5e+7bC70z/Qb70kuM0dNS7q810
rIWoiwD9BFP1y0mrgdWxHPyWiq22ONJtwpJ2iT2Bq26mRKerH97jpHWMHQk0N75Qrncp7mBPRPxG
h1UWGWTOCLHX0UGKGQnyFP0jXb8dSc2o45LYj9xSHvGZ1n1fU8Gf8rV45ANLx82QFHAXzv1qpYJ3
X2E4hnOsFNeATUrKRKDWNchbQ0VkwpYKTer0hyA5nqQVX3eaQSKHsDgVBwiqCtAGgapuaEkA+1IH
K8/Rvmc8BHLJRPyec5uBmP4Hfc6jGUso+soGa/1LXNQgaeaMpD8Y/qyFJOLYxxgA3/oA2dp+HMhh
axFvh8XhYgBiCIDHEYq87V8WtdCkK1b7UOO/LYTPKQfePVTv+nDoq4JZee+E5XJpSZTMqFCCg3SD
fz1xcz6ghuVyMy9OvG8HkOkpD1bZIVwfXLFwfaKxFzV1UphCnLIj0M+uXuDfexZHpbXb5Z/98WlE
4OHLCUOBUN2Mh2rUltsrBhc/wVy5T8vNHLeQxvimlRwxwRqx/XPHywaHMqLDVhPeUaEA4PazPmZN
/NzPudt99oWDQsqHrBYbyyTe0RfrL981dlFBLQ6X83RAhfHAJrFFeQLFpvK3YG0tnX3YbREm2SGI
ElMykhRD+JO2f7D1a+PgiIqglyrjlk6ztk2/GchEkgLXxHhYyXzoW/5DvufXpu0mHl7B3o9OF7X9
eOwuXxkAYR0dAQQ1Oq1UxiMs1/ZCJmET5bYowofQCtS2A9pOxnu+UCllgX8Qag9MwLDSI58k4ruQ
68w4Ocs7ze23BFvD88C0bpk4do2MGM2EE6gTGDO0Mxef21WzbRGnLIsuZFhgwJOTRcs/GFQvXr3H
bHiRWotkdPTTn72eTBZIqVR8s7GrdroHBLiHmOg7cw400vk5TF76BRwXxCC2HwEnHFAV74f6Vk5l
5URkPAy9z5CiRwoVcpvs/D3+qYKm1BDVAYK4RMvRlMiXZ7MNOauv0hG9KG5BYEfGCtw7h8BiMV6s
3Y2beWGAG2pwGUvt09zHD4JPbf8U05JjLlkfcscmSAuaBgVIJlAI3b+L4zD1obKKTouocEvh8301
BJlDuCFDojK/ax5Ysd2oZjahXWy7eizzqmh5WA/Hs83uI93YxIyVmJdgcExnNN9DwOnQ67R0+IBq
gB2wgiXF/gpl7WlNSTQkoEusNXQV9QXvqWYcU2dXpxwua61XBAihV4/R0a3S89nGr4i6BahTrZ9K
NWowvI50cabG9jYSq0EjluNNiDOKr8YhycoaR7fjSdFh/X267plzJL3wm274sLD4w+6Pd7z1UlW2
d0iZmknJFehzxj74h3UbG/lpTrSAUFn4bkX8WU+p4k78koRdkcI4pTrwCsGWpDc+r16TPO4hAKZ9
WEvxDRYk12r9Ahd0OC3B80CoMRN7sjzixhqvJrU2fve5Si+JR+hR9K29DCYFT0mSnCyZX9Q79x0r
z7Pv/5Oj4hSsePJP22xAKPxTKCdRKKa+M7ywCQQdeS7rwIROvaGU3SeeR+9flaHnN0WAQ1xMW1hn
8eI30pbRMJ7KD9dmtyiehS0rHoYgSmyKSR4DKGl54W3mag1N7ZMrMUqQnhLf1Sm6+hae9WdhatVH
1cx8Jynu5RBwvcwpRMb4Rz7aEiiwA4SB4MZDdZhz9Du8aRhgF5P/AAFRT8ErgJzqTV9kOO7vPoBv
AQlv9ZyxYKYyVAMEY1sxsjTRwDROgabjQKHoIqA6WXD/NBHh6CE9a2CZZTynlOiNX0MxmF1Om45r
c/Z0wMT1zn5c25Iy0jcbOztf08e/nf7toj2UvkgvD0XQHghLMX96gHxfuy7SRqXc13/nSa5mhZvc
6S5EWSl33hnI2NJXQwr2le6Hn2LwTh5kdwTIPDGksyVevmctCjgGRWDtHBS5Zc/aEqVtN31y7WTZ
j3cqtJ9r8GFOZmy7oG/SuhD7qelVhmmMpOOWf3OZUMwmzhG1nGMc7Y/FpG+IPBiNjND6EZ5PMKFV
m0pOYz3gYBF6CSecLOAwGL7pm/U4EVG1YRQ8p64uUwJeTGhhMqWOLjkWuWH9NZfWbZ/E5mW2Q/de
OQ2OIVa/y/dJc5POtg7DGTdPdOMkmS/B3h6xPiTjHityWx0mHlKbg2G1lTHMDYStwV7nWMU7M2C8
L1mt80afXrfnJB/CQIboFu/1IJ5JQyjXnNNxmJZcVGTV7bCVVatPkuro0SKFfmeJB5ciu8wydebJ
+hvwFH624zSJ0fJ8hR5WC1RgBVXpIfmn15tv4LNhWmGtEwELp3HUklzpGuclT86AGy4oecZBoJgW
KOorWDcU4ZX/WBhwIBFpnOzBBXH+C79X2IzpmIW0eTtfZWhRkc45oKA6gAHhHzs3fsS91uxmCblI
71mQepKEj6itTsL4WEju7iLG7rGyYb3yVBBIa9WTNl8To9Uf9SA7TODlh0PWSD/SmRDeJPW4dFQd
kuulriVHOLIw8P6UNJd7T17na9BtSoM83TKQovEkcoC8/SjkhWi0/MVycQ9JCBRm+/G3LkuxoTDO
DafS5yaGc0X7FIhWoY4enlRc9c0h6ERbCKQFSmgUHFh+q42OerYqlTXhUlzB5qZ30ekIZHuJ65u2
vab/bhikbL3hHfoUHNTICRZxwZ/iDQ7z8hz4lEKDxAe1J5zDcSIDtYGgtFEa1gYLX8V50qveYpHF
0U13I3rmOOJDOWJKWwAXGtLKTROkkoDgx9FINUwxD/ASWSMXC8nxit0Lwn6QoId1witb48w9EsDI
OwtxJVMxIFNrlXqo0Id0XldfjKmPMT0ihH3gS3Dc1rBASuyGbyHC9jYR7NfiatS4dOnHYB9wCE+K
FXfKf91GbE1WJzWdgWieZsSRWh57s1kGGfNWUhMIcnZCJgN9MsWDGm5fxC+lAQRzF7MHOWDA7p3P
uil1Ysq9aIYjG8l2q7EWBSOS7tmhlY8pYG3n4j0gA4z9fegCiRAJ6WGN79xqQOdVII3ucjoU6Wls
Ol+jqLNzLOIUsWol0olv5jYDlirsurVRSV1bmnm3desQ1gLBOFFtJ0smNwpx1Qog8FbhSoXvoUac
1L0PmP1DiYR3ORWC716IVmIInbbH3PIt7oyvK0Ij0eTT34atb4J7SzW6XvQoiQttAT7R+Bd6YBq+
SUqckargk7yurmTjwpe24GNl4CNI3C1AvDen4t5s42wX8VTGzjENo/PFiKqWvTTMYF8ua3pJ3JVL
w5yrSfb+g44o/rR3FpfCxX/aloSOHcUrfChKekRRCHUzLJz+HfUa5V/ZnJyWj1rWfsZO0jZ66juM
egh3C5KqZHO8GA2mVE+aUwe4wz32GKkREykZrjNEwYEry63nJzaE5dNtfuMG2ViUI5ljGfNDwYso
Lp1W5q1Ng5gHLrJcAAWFu/NJNE44OTuGbrwDk69Vk5WUf3vfgg3/FtOjcxDPFyjioxXJXIQH68BX
97nyG3GwpjAKZ0ShSaRLjUyWymmKrhgpe+eqTtzmkB6v+oIkjj5Uv6PUiX4T89n8RMHdwlG0r+Rr
xeRqutNhtrBT3K5/2Q4MtmuGhgvIpokprkSUKoA0GYKmWk1yArCpPkqXjnMiMuRTXvdo1injgacc
WDh/Ffl/BbMVFf/a2i9rqXOmvIl7Z7vfmQMygypeQBRocoBWjCK7Uox3uhqHKAmE+VbUzII7hIJO
vph7ZO2c+qykMjHL6587T9QwWc9ePJCiG7HM21dg9MUuENjaW5gRZOrell4MxMTWxge2OJeA+zhz
nscqPelS4i0hZJcPa/JuRUqxnep++8c08DoETBcVEVM4DAs+RUDFNqs0ilzWqBiTZhhx4b84cGJi
FQyY3e5FAUzIRUzt4RqLC9Ko7/mz0W3W+w7xsGpL7L7B6UFk3snvaC5HGmfPGY45N4TFM7IamjR4
0OTXqdQWqkAyWLHsdwJ58r+sOInZvvzguJv5dLoyi8kT3Qv25UBq5GBhDioR4ibS5w8wk8t+DXZ7
3Gg+ncjbRgbWyaCRwdz0uJoUwhVQYtjUeSu9VrSV2uLNEbNFW13ZTGBtMb4TLyXsf+kArfwSJT/m
Tf4uBe9N6xlBDory3aL65FZKRC/h+W6KaLMh/ldLewLn5T+IhedA23pW2nkMGKRjCpNymEoVCHzG
ep5vNe2IMPjI9sFNfeYzCTw3C5CfOKxfLT5iP+qNvpzMFvQPkVhobsmiGg34+bpbyCxhS6p0pR9P
DnGZ/VX2SSSO8o7Dh/inbR0IvZmsq9Lg/VqqnVniVpFYMKHQY4J6MTS+Ai+zalFe5En2HmyERUJy
A3smSWU4/skg06gjz6delvC9qfeNFaLHQanmL5r/7amV/QMjcDE4IysXQ9+mlWFtiKh9YcigdiJ3
qm5rvOZjqeLWYzZ7rPr7FrSpPdKe1hZ4zlwkAFUFAqcs7fmRKBIPn39njFyL3qLoPIi7bKq638By
lrpE2vz1Itw19Kq/nplu+5qCvT1OYNLzrv4bL0DtpuVN5HBbVgLi9kuCRM+WLkEVAXlB9VH7o1Pi
94RWv3N6QUGLmXJ4i9RrWoZPAcAjbOVvTETnXExPNnihTZSrHPfNLt0AugmMPy9Gx/gvtJF5yymy
a4rDZsATsWdAFxQ0BFJpn6dTLPNVbcDZ+orPZ7zIW71sDraWzLV/phgOqlt15VHj0cNjkKKYnvCr
cUHDmrF9VPRf1mVNHiZOjQz6uTKKGepbApZxUI9DZoRehs7m0eWjnxdMmQDmiKDhvQGviTF/1B/e
fk+kdRZWnkKlwFi8VjFkN/w+8FYbpes1JZ3iZiw25GAy55EwtBdMrJb0ZUUGl2/s44IzYa9STMK9
TvbkwglZLkCIXSjBFjp05hq23W1ztY134KayWOW763uq524WTrDsNqZsjmkqISOriIQihht4IENB
DC2ykGZ/hy3SsNOaC7r9JsH0T+iB6qRmg7JpSasSnw4Dee2zd/adO8kSvf7gzOAbbd+wqxoOsSa0
IAbnkQyRb5CQFRvOrfnTp8A8v4il2kZWrFAvS+K7jRWPTI8MV0yCJrqoq/aZeu/NZjzA51PwUIbM
g5jfxijJonNwB7pEFi69/KZT29+oxXvjBjgygL+RcF2TkOboTiOekgbkyXAVK7zkIGGa1Qw1Wy12
qhvZRol4wtEuJAS/OAVBPpGd/VH7jFmCDarTglWrvzS2RxpNp+LeMmJ/v1greDOZL5LocyjdK5fW
ud2CF5k/UK1NlEFGj/u8A+OIFNtEQFVbQym5/U7UqsTiuZ1Rv82vIeR+8oMmfoxEwFtINXKtNuSX
hm9qoRXOGSQRa8lL2rzHscdrGx56fjS8j93JgAmWADpo9PTdJggXCY4rQEmR9ydBwF9uZZjvMPtJ
7NjsNMZTni6CH1el4/QGmvyHMEeBHvUyYopb4TSYUgLjTa+r1XPgdLqsGt4kQeNdj5vy974audaj
7vVnkZnj58kNFrmKar3zktLQSZORRExQbwV+JmAl6GQsP5xRqRc2ILLjsfkIlkU8ZeLkZgel24nv
o4dJdo/bIFE7o86MZ0F3fiF5tGGfLFibKXfhcXcVrNbWFk7inBU+VRcwA9f0m71lAgv8X67D61Wh
qNra+yPb3sSK3yqgNiq3JciRLQkBLpW+C19Zsqp4WkW+8vhXrrOhXkOy1+qROd7RGfNbg+Z2Im7r
yWWAjW1RFNRnxUpEIJy2+TwV060azQQX5Y1I8AFlXmslCAVQhxl4F6cspoWkAbwMS/DqBXURG+jd
CImYrQ/Qq5XeXmh3GQtHyV7vz35EkY/9kJOQ6cvbiLDVBh/CJMjn/UTPTXafiIng6chruQmgZMlK
tRJpKlER7diX1XtAxWciW7A/d7RpV1890T8lXGvLnFpMaWZxwNGvgPoC4g5qOO3gyClg/picR3DD
5L1r7eo/4wN9o1QQjR74BZ9912VX6Pgr7hF6J8jV9UF6G7NHtFuF2nxdhf9r8V+xNML5YdcfJA1f
DSBmDr2EtgZmXa1InAaIq1SENzwAmMM80+5SANfOvBfBSkHhnvaqtmWmN9aGanc4KCU66qG4s/ln
x9zxiKKF8OROstLtYELYd+ysUIU3zbgQhIckkW6RoTTmlN+dIAxU1F6omp9V6HSLptzWpcwR30zd
6zHYVvkxxgeYiDExOhYHl4wVTZL8FzNeFJ4jXOHsc4RqCtqMYQ7rq48bGNqSZG9vLZLEPcVubLRC
ZSBm5WgU9XDegY4RXPSjUz9jZ+R/o3SnKAgHPXhDhG5LbEfoxPizsForLqj8HhMJVOGDQuhgGl3l
OdAqOEUuJ/XrT9Cyl1M7rL4TNZ4rz5z5HTSljRTSA1Jzxln06E6nvP0Udup4u6QniajFAKWb5Wnu
Qb5xerVeZLPQAAawi/D+pYwaAOZVDVjpJVae1oER0kY95MNLkSxfLyEXABFKeKRkOQYqqdAYwGcT
uoKgWXNErFY+wXq7xQU0es+YN2ggZIzPFJA9wKM6rgDXKhd7wKVzBlLbRIAboER8m8JBKSpBRy6h
W9iKWxWx6Ejy0kQiJGbbwsBgv0cpQGndsii7/5YPET37oIEhnPz7XiAPDfuCs5UnLNL2QSiXmrIO
+Ydt7LuGtzfORSJGrNUdTqHz+wqBLOIfDZ7VCB9IG+Nd8apxv+som6cZXWyLMc0wW/l+Wro5uDNY
xHv92XdggoeNNNVqnZJ8DCitjFjJaNvraORzBniZKE4xJE/7LckZYVCpVweKd6Ay/gkxLjfxmM9i
rSbbzXXmOhBqxRFwfrYkCHMxyHnlZkmVOewqkH8vYXZfSOyq0CLVZbJVIAUDM2OtF0WfbeQrhsy7
kReOgdLwwbqvlXNVvQpzZr+boHE1jCE4engAVKPhCRtq1Raj5hMnI1yV68JaIrPo7OWeqotiK9yI
DEK/vj2SKY/LLtqHAnFgYOtJowve1YaRkrm1UUNAqc7m1Txxsf+QooEpGF13ERZJTt00dDo9Nee/
WYZu0EWeFeSV//yXOxT7oLVbLwtYI/vYo0rhlKyV4HtqxFIbDxr34I6kRySHgYHLPW5lIKLinyVo
X8C4t0HAbSC+hz9ahDoYDAsswpr1bufpvJ7TKwuqN7LJwOpOztYVmI8dcam8Qd+2KlZ1X7+AOFVe
DIk/EYxoxsgfcry1FChE5+4edlahdCIU7Hwzvrmz/9f89SizQV5FPdkQmuphktmWz3n/MPUQqfAp
Eh3DAjqd/WHfeNyMAwCjU7Uhr9d8ImjEeo3pfdUap0fOxIG5qlqTUQi8BLVp8l6I/IkOdOxEBCUu
XD4/yhVWRRjoJ3N0/JI44idgEiPxmZs9iJ+pPySB459+TaktFPOAalw7R+MHQy6Scy47EIAxaEjX
1UwjjZX4WJ6FY6YEW3Is6TxElgRBHibGzozMx3cbMmdM/8sHKysh2z4tDG1MeWbma2OzSQ+d9Lxl
KEBKElRIhkOpJhEHK+V54AChunsA9BGWOHAgEoFmI4WN9Q3hZn/sNgh0k0H8Qw9RBdirc/22ptKK
jx2felugrfaootKBMYQavt/2GcIAMMqNy649VObkS7dE+hA8lcb2YfG5EkEvtZq8WD5kP7Rb+C3i
IyKt1Dt+pWfuwLb4U46mQyt03odiLSB+ibCe30HvQ7HDIhSvfdZPXprd7vJ371q1KRdPOMlz0TUB
anoEho/V4P3+KBZT1HCXMBUHKd0vXCgt4EoztDWhAJU1QZpKDAkOXKig++fzcdrnZhFrilMRHPg5
ZvF1N/D9V4PO10OC8hXheGAehaTqzMLFXh8hT3n5SnADatOMgUtHqBmKfr4iBkEqnJnW81Lzelal
wfKZsHBF09rKK4vSJhQ6e4x0g8OJvp8X6K/b9GDI9P1apF0xcXT7Gc8Sus8657YNKCbS4FLYCCyU
UX+usEVmunr9saD8Bzv37Zc0C+uGerYEoci5BMfImn4kxuKIj//llCsnZTuylUf3cTMTlB50Ujjn
avoRgURsXkDcHARfcS8KO8/rU+zimOwyFB2GZkujTp/TOrj+uUKjq9CbB5n8BnJ6pnWmft41Tkfv
NmwjT/jZNnDWsyo4q1obCo3ybDt6FDCHW5/E5iWULKnjlyC87no5g0ehsUUJ6zSweVtZS97XEM2V
K3MYC+xL1ui+sfvzPP7uIrnJ4reJT5eXbW8U6tr1hihJIwbFANtl+0OPK4HKa7ohu0AEpgzkyq/Z
lrmBwsl7wqzFgTEgSG1SBHfC8ggP8rN8VtDpUJ3koVZA8vkRPeNKiohGGFwdBrO6mUcTN+thsy71
nzjM0DKDucfIsrn9+odl7plu2BvASUZVxhbvSbv/IKh7RN8W9xJxXrABo4zylx10UA4NZvi6IsjX
Lz4k0dwqWKQ3ObMfrgRkD286TjUOXPuLdXreuCL3J0Qy3l3nl/zSsr4vFLIqIvXrSbvFIlQDl3q5
GBJTFSK5fEbZz0DwvKhJgXmag6zMGJ0ZkS0YVszPKnFE9ZmqjPFiys7HYWzZwEalCoU/XhCvsFdJ
2mTx+IGY0WMuKsJUZEYUjWQCQ45fbyQlxOySd2mCU4rGjjX77jpewj+Jz3xZvQNTZrzZUeBDkJGb
imTKqNC0Hi3y6XhhAFYoXq/JhdFTiCLQ/d5QpeX0rMuqKIGN5EXtpkzPFCD2T3xBqLPXhJmTuiW+
HDYyQYLTT+FMUFf7ZVJo8XPmTcoD8AHlNeRUDJB3SgG7PFUs8R6221xnEt9QZxh55F/t2/limT2L
W4G0daEEjPuuRGC8w7UZp4xror18dSFzfnOugiVKyKyHX+ZkNIJWh65gCwfkm/WwhVhk8R32bKnj
NeF+jfu/EEVqdWhMvsqer7WS86Gbq+NnfjOn4B0Sgis6DoJSLaoj0NoosjiekdmNDBH7k32su+nl
iwhXAdCNdOMv6Egt/Q10Ev3W27U9itiuoKSleHj/zxPSSbXPLKBtINF8MP49fYk6hg+9Z9+5AmHv
Np5tmnvss0Tm/+nQT3+bwEsHzoK1bIVz1sLhDIuOtnEBKbHedEMOS55y75oIWZRQrpjhNWu/JNCr
AqVpMxRZhhlSRTIKNqq6TWabaSdTN3oFpvgL988Dy6yla22XXpsCNbVtHThhwIrNyLhQBNWRIn4G
xQ68pQJtbWvARY/rLpxhj8D+3yWnb8wHvGVAsgnWcQZnJiHgx8WEcfQOaPyFG2Za18WJp/vT8MTC
5MjTz0Egv8NFkUAoalRVZnnKox1V8g+TOmzU3fmjZamFG5aMZVHGCKcbbFP/ZgU3P0as/lO4bl7q
XQguD6WC+ab/qXAwFHCbVcjPjGKSgBzw4gLCxzBLL1DtwdZVDcXJ2EV2wymBVIAPsjplPi8UzjGE
JednNR+ygq1+kOX3Q+jmYdNq9UQXR6FvmKK5qUmZjwrER8I1mhUhR9A8Id5dMSAedH/qsVVNEm3z
dILjDozW/ov9/aKTprSZH5IHwKWdRJArjb+9I7XT/wSJAJbleRR/NBGjtNRWd+lurkdp707oOs9v
EVeAB93Y0joa7qLrOHjXFxo63hOEr/fg3SX04fcbH4EycwzERPZO2YbBi3ni7ePA2rNVxyauru46
0gaPBiUIiNGVk8kCALGh+nGTWbww53/t6s20dbjG1qWVD0WETUc7lgWl3TefHf+YsO7NFeW41BLG
mUzhay2L4/XHeWpJC5IDtMbTzyCvVO6xKpLnY2QF5bChclBtINfon4jkgmMBOX7vJHyU2JjIMT2P
4MU3tWFbU996bWJKvBfGOi46M5cjRRnujiF3/1+6i2gc5vTIV/u6d9qqN10HtVs9ux+rK0T/JzYy
Gj4w3Pw/Ko+mO1JeVm5LGOM/gSAQLi+etrhlsbDNSWgbmt0VtZpMS3DPHFfLVY4AAUW6QnYtepM9
HRETnQVpqxIuLC/7Jv7dIUZhJyhEwBClUOT3CxQNBgUZRn8NIfT4VGLvgnPYJpo3qqIr8A7fMWTV
3yvV3rziZPCM8wUd2JKOn0i/KXNwD6lln8WBDYzjA1pYoQN/3SrnzdwIYu07IQAm7tZQ4u+QCIKK
YcLiUYpz8rm25x9Mr6eyvlstaoahwigSwsbPo3MzEq1p9e10d5/m0vOj/4ts68GhvR89mUfWL7ZA
O/K+rIGtdPfLLy0wgDjHosKGWE7QL6jSwHNW0FbuXsGzZD+0E8QFjZpGx4ICBg6QpItMa5uJDiVf
hiekCgoFx+85TjieiShQzJdFGpcwDYbxiNfnlr5lHNJpMi+6ibisv3beZr6evWX9KOYZM5vHX9QD
aIELgVObiqnCaVVIrTfZyo60fxDtHWOWZzUJYD3JH3umgCScUtLAMK2zJaC7IuK+g7qpz06/VMfE
dW/yvbUwm1kIdX2rhCOtD8/WroRav1iv9FwGvn9Th4DJTlkHrl5W07AXWxj4upXRPdbAbZfly9xf
KHQEg0zWXNS55BBKgI2nYHbfwkuGOMHFzn8QkyLqLM9JzWGIxrZpvq61E0ksHirwiIb58rXt1+ku
f7RbolDg98CgF6nS48jHApQuE2GuYoE2+zcwhntVvO/10msbxGP5zFP7jv4kLK+zVuY+tmeYXak+
LVQj5NV/SI3Je3M+TJVrsT1QaXDxOlcmgTi7DCObak+iEMHdeBcPN1UtqI2DLqxBJbr/BAFq2Md4
xrtVEGAZIbzDi7KjKSWeRlMHworGwLVvkC+eURAynZy8C0RgBlEujta3zRhuAvHW9GqR2wX1nNRj
U43snsGKM4QI8txlSR1W6nrBj9m6pcdXW3BcT5twdWjtSO59RJVVsUDK5rS6Rk9Qb52rYPygNoYQ
N+tH4wd4ForrRi8LEMbs0huHjjJF0tP/lCphAKf2qFUFUGY7UDrC8D/94SMbh0ehVMv1f5DSuHXe
iiEGMq3Q3ViQwt4PkiT35sNyEJBqKR/r7l3uYqsVCZpLCDzNRR3XJR8rVTHpmjBrQezz8m8L0yXo
ZM+AfeQ3+pXKSqlpT2ByVjmq/GPrD1NIVSsBq9dMm3cFZXhJg9wQa5LBBkwj3BmJKiV/TBL7To1m
xN4P8tWdD5zNaf5Kr8HuStxjzEt0R4H2q2MDSh4EUuOQzub6NYPhAQI4rQtdnAa9ZvnJAKAo1O/X
H+7Nihv5NE6h7hVys/pFnCm5vebNGj7NqQUl2J+NF4QYyXphNfPwrKMRD8OA6++J7FR+ucn4Pgyc
Zz6xVgevnntANuyH1Hur+sfwwtaNO7uYyDob8M7wBUjbZvehML9ewYegr5ydTkqeOuLVduRXmwaG
95VlXvl6DHkTgIJry86RBtEB1cysTuW8NMdNWhfx/R4wlyasgexjF66Iz69hbSbxBWRAZ3TCxcRK
+hr7afkUDYCR0daddPKzPUg2vbIC/Dt2EYkAgmh517L+o8CUT9HuySjc9XYWyZ4MsnEjyDf7oSkN
4k7hsiyRZZYERTWXMAzVOirbEEC3t4kXI71PG5rMGAkdnc9jw+hVWW0ISv7VPYDS4N7BnIlpJggQ
4/X7PI7hm0aaAWL+yCZBgYiZmhlPP7LDLU4c53xIIVgvS7HmTWauLr552mBOuZLZ5SWouqsAUh74
I5yyUv9xX31BQxT+P6SdjDlxMw9N3y4/LSQjeJBa5VZ/UbbcHt5OMvviK6qw/k19Gsts4vDMka35
4+vbFlPkKw83ZsVYmaV39ZCiv2mncClD5M96KvuF25tc66sE10iH6TMHdVGAeta9ScWK73JKEJ80
t2/83AzR3nhPGHnXzzADDDJNsIZM1opTGYcM/iKsIb3gwKu7t9M7ChuVoziPgMqALKwQiX3z7n+1
GRdQBukWD75owgWZpyjlF0+mXeLSrD/1TrqvKEvE4/G+A28Vsoe/nDgqUEYllYaxyK7albid9DTr
kUNUHHCwJK005UcS6YOgPlZv/8RX+enZIctlpRNVvhq2DunS3x8x+/n334t7EfKHOIpRwWTXqJw0
m5NPV9iN6FU1fC5fRdklj2s1oruyy/Z94p1dFDwiZvZjW1h7Ur+MOWV10Z7YsLUAs/RH2+9e4f90
CaRVkEo91SV1YtHCznpykK7d6ZzJosdjy4EVMVzg9cQCC2Qglx9zNc2Aa+48v1QqJSapk/Nl6vp6
oeqHTFoLYI0WkR9LJXS9ZZyjGMcCPxFMAUkcG4BDL17nzS87CrMchtF+4XsXLCwTW4zbn6vGeCpV
gE9MUz5vUCDs0jKRXpclGDwQfaZPUmJtachIH2vcxHeysXZqy1gXAQsYcPczRdSo34Lx5jJrikm4
JmfzwOnMtpIY94SwRi+7efsCeqiZ7imRsAAKxaOB5vem5ZlxqgnaJ96boClxk+u83iaFRU/UKM80
ytkKaCX4tOAhky0B5lfSMY4ym5REpotN+CGjmHd1ov1n1khKf152xRygEAc/ncKOX2Yfbx+1QrmX
JXPN831TX0KddH6SG1kIGnF2/sUc9phcyt1YoFLW2vWN1IBvZ4+Lyv5qMNUBs/knNkdUdzq8ij4y
TDkI0CXalR6lVxFqgqJTYXIo251xNqEGGP0uUAO5sCnNb7vBTwXZCdExC85di9VTWy7J2Kvl3Zrv
RRSqddNaGlw9J2okkndO+hlkWgoGMSOYkAtsTVOgOuQ9dz5klmDHIsXG5/pcqbfxl9+PearxNJfp
kZTutpvoF5UrAnh9tGHKGqdHwfrJTayQnF1p3KOXQ30pasBcJMVrsBmR38pO+nPAV7MxbTXN9ns5
xFPHL9csw99S60yzg/3ey5Flhb57nLXsReRDhKvOFeS8nJydIkM3Itwb9e31uyAAc/U91GNQhE2/
WnL2lCizbJTpF6DuDh2pzd1oAZL6uaHNoZRy0yKE5pA2P3VUvRvQNxwScYU9JLNq7qaXby2Nv1J2
1jrXK81Lkkhty2C4Ma9iVIf37zmeFh79Mv1qIEUwPDVsBQ3FzVcc70G4eBabee63J10jvOnRmqTS
o/yCzK1Rj+Z0jPhYmmBrn4zOPel1tqqCeUEzb5oTcFmUrxA8vyKDAQPq8p0jLac93FdRUVRDZJoz
OMCXYdGp6qexgKuh9dYzNMIMJutS3eu+XyXIasXPfueWTNKGmutxI99+UUHggW9wKkCuq7fMySfI
gqgz5ITO+6Rai2XCJf2AXX6bPbwdGjN5LiBKAUCFjEdgQd5OBWlyFng2ZKWc65SQL0TAS0XKZX7l
sOkXjmWSaId+ab97YBPiL/fBjs7EtoRC+ISI6Hc1Ely/yS+Dv3ov4TYd+7+kw/ePwskAC5xMKTGq
zQCHmRlCZm4dG4uh362QvKM6+oMx3GLuaAvKTM8Om/j8NNjSpRLmi7xal+eH6Bd8HV8rWm1230cI
RUSVxx+yndA/Sv7BKFryMKrmO5Jlb7FX8P9merHF+ooATVTAXgwpSNNnFWaek2Lpa+Sff5YeYF2B
O2NczaO9jN4GXA5nYXD43SM9JBBg7B66vXSBsSpO2SWvrYjEicioEf4rUIqkeqjGEJ6akqaV2TR/
5bQiy6Gp2UoTr+7BLPj3aaZh9sHyCJxvMMtf2qNINLvGqF70RK8ch1kkldsWjJya/r1XuWZleLCG
O/NaGjae31alOvj5hr7VWMM7JYlxtrNWjlOa7QHFJM/ei3uJAm5Ehr+XB+6IfsG2I5xxpkz9Ti/X
gb1vbS3wcK3Oc9O6WcRr8VrJoINlH0YKN+gjzJTl2kIDGH6EH9MFvo22b+kGr4RlOpANt6E48t+j
SK6u11tc6cc8ILlDI9iK6otUv8fYl34+9Gg5kO38sEOo3vvlW2OJ+vgoK0biQDT4PU1uzV21E2bZ
8xNP1Uq0gLrVlC5U5vU5kDXBLwENeqD2yzH29lYBG9rrU2j41BbUhwMsrNL9O8odg+gfZyD23hSz
2FLuREYDolMh0UOt9msrB4yNFPQpAS7b9RiXqWEeqLuI7bAiRkQulHZqIEfRIb0iMFLGf8pCRC2P
RLKCNhLNwGLpcpKcY+I7Fb5PGUusCK214CyaOJCbfCa5/vVJfUSIuJbvoSrc1MugaKaA9dtfKxVJ
JBre6A6Frm16VQT7Fq5aa97puoAqnftzzTpysRxgsVTi/2iJq7nm/vtYdryfVADn+ed8yf/tfqWV
J7MQmmb83UQjCR5bTstRCEkKbYPYbiDPIa5AdyFlQKKPghZEP0J3xXMsRKCjkOn3tLWvQbtJgPJs
/xI8WZv2KnXKo4iDBLRzhNQHiRyLir5exbSy+KRveEnyTzZKW1sJ6Tr/tPJrOtrzUASBVpeGk+Dw
2eC2kT2mSH0mxHsnuvJXJLZCDv5Kn/Xz+nENurZH2XxHLgjCfQNWs/M2SejMWfBircVfMPrbTeeC
XxY1VbHHXmAmniPL+xoOWUQZ6uO/r716Yph4QrIIld/ft1Y1V9PWIswyi6rf3J025B1AnY0ACFFX
bIEYFOvjDfITfKETRnkQoXun74tSWwRF7Qn3VxlBXP24fFPqsaAoK1JOBDDma72mtCEJHO2S94UC
QW01DMqtt1AK46gXLqO+mY4felto54oyGBoiOWt8WU5cP+JJZ7zF6KeUzxEQbhnIb27WX3C8RRZd
IjNKKechJ3o9UHIsrP8JH4yTx5F0vVpJpZYVMWBYP0ZEY3Y2lxhLMZ3/47ehaTBoQdQXnwr92Erv
UbOMwEcwqyQYAlBQujO9UxfocwqgRDcGj3i2IBUtheL8tFnGIe6OkAh3bZlLT/ICYv+mWA0pRU3k
CyotIKIg0LQZtRmrOzvEpWARlTOk4JfwQ4yKNniqe576ENdvTPM22DUwpRFzMrwHNsaLiMn/HOR4
xAu0y5bQ5M4QV5twNpfCMZG3DMxIttTgX/lXAWxkzGQqj0ZzBbkMhxZvKQm8P1kdNSKZc5Erwn67
odtVtHCcOhHV9NDrMHTTWu5R+QiP1k/xQFuy6LQZpimXnRNMcfv1ZfELm4HzHedjjnfxDmQx7s4U
P2/jqvbOh3bzRTRDYz0v4kk+m+Y/ebBvIlacKFUFbE6mIHsT6iiu/kseVLrTFD/Fcnc239UbxDCW
47I6o1UkjhvW5s42gMhOsZ7BCb/0RgUHYlpSI39AYX3797Fs6pAWZUl7v1m6LVXGQ7L7MiqmcUUQ
YVusfkwsa4fAuM2sG0sNv/V/xIotutXnbYRi1LvALUd3Dx9iD3s/96EDnQUaVos7Qq/s7HzY+tAq
KWM+4K6D4lXxdwIa8WtDfWpshbSdszPk8iKxQi94ewmNVWwGWPvyr0LY0XUtOgZUYzfkHgsC/msb
jvondXXwvTY4o2e289g2KMuFB5xmHnWPWfXvE5n0C4xe4nxxJ5DvNP0RhUAbf38U9oogNvtdRQj6
xH/7LA8hfnD22Uho5R1vjckWnoJvICVrnaSHaXzPwASwav+tFe+13foxQ98+50AO4lgV6o47tV7g
e0m9spap6WB/qcJDUMGDMVuld/JR8DusrHwxVNjDDOpjE4K0qS705DHs4XciU6vqoG0+KAntbCtL
Unn6fHqWVUI+7iiliSWu00BrJLcCY8fxkQ0bF/ZKs3HtSdtgYUAs15g+akv6Z8MSF9rsrPWd6PAX
mBGFrJbAPuNZrsqSWvy0nqfeKjo4aYdAgT8v0QoLISBzyixgbI7tOAwnJhFhNKDoPuRyxe1pP6b5
B7DraV2WNI8w+VUcy0PWefgcxa+ydGNqF+g8dEG2TFFcVpc2kpReLRlwhDvQnlhvxnI312bwLLd1
IHqVvf5+Y/BVNuTom2quuL9dSnujh8PKcLnPv4k8Y7PO2rTZofqOuqXZNPcDrbqkSF2eYgcjyq6L
PxWO/fFu4Lok3xW4YmEL7eO3lV9jmYfN5ht0dzKNt09CzsVHadr9PAyTdwlHt+OT7fwLxBlKGbuj
f5xjvLdynqPZZ/R+xKOLKLOC3Fe3gxuYuwAbMts5jlAgCrWjD3nM45CkwtsuOxtiHIW9PMDVfqxe
3NKF+UjIC7QQPKdagRiL7LjoNjIMRChsSjFSQRIXM7pmd2ONZOQzJK+n5e/kYIWjWTdwmoFCDcfs
uHZSAY6auVkb7cZvbxMGHFwyLSAx1+1IvbBcicPvnzgTCFJ9CeFk4UHNoq3OOXMCwI1LD+f6cY6p
mo3A3MPSp9TuYQjj80ubSrhKSFCI9EzNrm3upE5P33RCeYjq/rV4vF16Iaiv9atz3wRP0QOeVVqF
WB+Dah9ZHhJZQon1hgGw7NjMF8lbwoJsBwnn/hKybmig5eg3N8WNMPf5Phb2F3vYwzBaEfjdiBKT
qmrwOYkdfkVY15Q8+X/ZrGvKfwm7Z0+Ip663BEo7kExQNaKOC4X+AAKoT7B/M9gNSJxQnZlMZq2+
bhlU6m6Zx+S9RqpmRrq0DqUtbGEmyBTQ6wjtOwyZRzSdFEWqxCQIWnolalnqEmheHkboI/5a+ta0
oeWXcl/ZI8ot5WHTPUj96trhhsVyqD+tDsxMWbmoQwplpmn0qa/KddjykYN0si3uk9UQQSpmMubm
y5kJCgvm8yVfKsCwkfC8nBRM1s97H6pj3xci+bDfGO+z0u7ZkUEZ5ItC2feFjYxEhpHBoUvzdlqz
4qc+wnfr/wVD56fOSE7CdzrMED+AUkOCGFUIxvLae4haoMoMxkQC27QEvlHS85XSWD2ibg15bbVo
UvP9rFxcKhCnaT4NIfFspNHAPIsruVyJASzjZDaZsnawyW9xKpsGf2oX6b9yHCEfpb5AqISYmOyf
ibRC8EchXB0GLL41nKLLa4g6Ng6d2thohV0viuiGxzy2FmVnauv851VhBYXORjHf0+7XDo9rrj5u
WkjXNHLQjC+SthEDS8MBVBeWf8stphtWc1f6BtHp2xzIlP0WkfAMI2+rCPnaf4PIMM2/woB9W5rD
FhW2so+kFuSbEZr0f+mD28vWcMusV4ZFNgNt8dSkStnq7Jbd/jt91/mQpK5Wh017ug0PSwk4kmc8
NqwAR4oxWCa1lLvJihuJZ1TMHX7s8VWkbaKUD8rz56wYlkzILtuJaqnPib8EaRD3DZDsnfEew1hk
rfR9YMRRofPrtF5j2PtvD5yeGYbStIu0sBIS9Po7OoqNPpa+x33Gy2l+hBMsApo9pg5H55WzPq16
Z0kLalht5l5ArIiqazds3OomK+qjQJY0hsysh3tMOfIHtRqmpB3a1z6iy8Hql0KfYwblk6rdFjuV
GIOAa2KuJ/QoTXq+ipWPQGEQJOLUIW3ribDIFPzmH9p/eZrrsBoC/uYKTLQ2kNWEgIB1kfi5//sb
cpG1TCd/XpreERQcu7oxP//dHz/eJOLOcC89bH39g5oWs2zlyzrCq2LCPfBbg8OaJq4drCHEp6LO
56Y7Oqtud5yM9TNTr75+4qFzQPcA6nPEklHsHV5/qoHTu1wDpUeHqxQhRnpH7ZPOWGoez5ZGcrWL
JSCx8CjOPVJZuTy0PscZ4jUvi79DyUUAHB7aV4HY1Iz/o4MKYAG2koy92ClIrJPU/elwnQNXPuQe
vy475bhJqTSpMQcS/gRkCHOA/C1FQmP4Q2JHpun5s+/2RNIboEV7mAxAv9sdVy6haixOxTbb38hy
gYWGHxMqdmvMBMiD4BKMDOfOqFc7rO6x2AnkaZh9rBzcYBxiUD65qXRPQp3YvFpquayFu/bPvUXa
cq2EM/rPve3PiBVsMyoAmdXrHgvqDMzQy/E96klwOTkhoPeT8k6lUAsURaoA8sCowCLBTUV/plzq
Ps+vF40rM5jTZhkMASRq1iMj6A1WRKHvgATEMPyYeyPGZx1dudlUlYeeDn2ifjUOhpvUZRFke3Zl
dFBy6QmZpQZ6FA4Nm4aFCiUXA0eyNY+zQqvSavIiSyoz9cxVvf1zcauOSbREpKP/S2hNm+kDga3l
2fxPfz7WuGnoN+M6YuUBnGxECnf5Wxk3jcGTsp0oCTKsKzKkIYYOQ4clG+qsFTg72w8jhmP20I3I
EMWCZBwkTyIJfnwduBr22EMJuG3+caTPOFzWQVh1Kv8LHtkZhmq5rPVq8eQkG9CPPFdOpHjfx4Tg
H4YjY6R+XT+TAltxYVgVwgyY45J9hVGNOAIN1g1WqP7oVCGDcFRmWWfkMXjmGSJBhAc2t+O7lKNY
4np+oAzS8UXwO08k/lerXU651zqwd75WS8TTBx4IEsGjXcL2l2KiyAwIjo4ztfY5BVUAiE1tv9wG
1SSbYVoVQyjYkS0yPnHjx77wMmWUJxiKTWm5r2DHYIZrWfpz2rnlRhn1CgmGNzX72ZSmzBSROnk5
UuVwDFA6uB6MMr28yjxPOcIMT/aknQJbHmDlLDfVKuD6nGju5t3ngSWNMDQVs5Tp0wgkvkKxH9KO
Y5NswaHqN0xT5dS59PjzTDn5oGPEG1iUqaO3RMG59E+hiyhH+EJlBwAfrxsHkJVNrx4EcFX46guw
kCBKMgjZg3AKpl1OV/yRUNCPzT14XKkCR16kBa6+2AEqDISL5UrtXmQgzfOGIzKIVEtJtHSW5mXc
PMGM8ZGAQbR16DkoZf4FYlTy8hjFRIP+ih0wT4QY17XrCCaXbJZ1UXucB9zndvvn4AgE8Z/skror
l8D1NvQm4EGxCVimTLTRhLxm+5pbkqwevxiTFDUsI11KRvlA685hD+XGqs0SClrf+tboAhCKBb/Q
yBwJthaD6VrcDSQYGGe6yRBISawKwyP1A6YQyWjk9rI7tcyGJuVaOdA2mrGw5Fw8N1SYjYcud228
j/ryS/ryJU0PPsss8KbGfgeOxuUHn2dc5dSjK13Ihh3LLgfIrmw+BxOTeAlVBFBb18zLIHLEblo8
O0CfhZzwQQLRlDhABFLxeV8q5XIeQQUG/Qpyvv/tvyQ2jwR3J00+BrDAGfOg/Ijg5doF2UmRGZX7
Vifsw2t6xHsjAmorDgCjbuqfkEwiJQR7gSbgI462+v+NdWdD48C+h4hPHxJflcokF0crwBw/ykxv
ry+Ie2Fad43OnYJHXRwbU44KtdXUe8O+HC4xkFuKSZcnXh0IUBp7vuKzO8HSaFO7gO5fTFQiTPTm
PVW3r6WpEiYAJ69BoREgFg5gIahsMrKldJAnar/qSd3nWsTkuwweoyP90es4AuUqhaFN4aPQGHMP
RPzC1IQvmDelJV7ZElYFHibkk0laTOqj8P/+oenDYWf8TOff4le5KqY45/6NcKFb64EpkpShpdEF
WCIMewU265F0vjLPtcFmoFSiQ9r7ewsXmXmV/cx3Kl8wj6gaLrniIUBphS5kiSVzh/a1lDv4IttJ
Lw3wUw9tUxRjJH27VVXPSd9rENSuF4Aambq5Z7jCsudEipcczFG2kvokrKYcKb6P6jMj6h91exHz
EOnCO08GlBvvpAiPgW3ku7+VjprCFrJsN2Rq4m2zM+KX3ExD71IK0A2+9R1hE32S64Di6W1hixTN
7LnZYMriX26shztYF6qDQfb7Nl3vij1g4vySRuyv4l285kqYRTs5IzL0X/fid8K41LodJ/tc7dEJ
vY7DYUMjyLLxnENGee1tOwapd4kA2nxwhKwdme3d/92KCm8gQ683zYI673NZmSEBc27JDYuggyRt
ggEuFNSksxztK1CypzhLXt7eUS9NvrThaf7+aqr87PA2yPebCbumjEJzfrQPLbX9sebQc4DC/qgO
dl8jR6v/pl3PmJwq1Kj5k6StEv7hqIFM7yLB+jNtktGVZdFjRHrsTvubSHbUJo0FFnnop9dZs5yk
B+E9JLAr1vXs9gWEhF6BzkCg6Eb9/TQZeIS94v5qf0y38eMlJM+KuPQDYOkpCWFaRTFbHLL1FXNd
7k8lKMH0l27gQm4jgTzzfP9oI5vSJIPVl3f45+wr61xrLIWBl9IPwji2HMbiTEZhlPB14XCquZD2
2dG78sWAScTjRkH/LPQlUlCf1nmRjf+07Rq9/JM7SxF8IKQ39dxDkCguyh0Yh4vmbvZjSuR1pGhH
pS1udGTC/iWhrJkCmhOLP5B2WihgfzXVETtn+OY/SVKp2xtgvFIhXXVuSCo4EAOS6IHQi6rLjI87
WazSD6yVhB2Jy+c7BqsQ1PeXiyV0GmBhwwEC+BCL2khfcNS7pkLFbGaGQVOWZp2H0Em1qtV4+WHv
w8ApZ8yxKGvXOz2Sg4DitExaZq7JgtufqOAq17u4p+O4YUKH7sJLAjROfZ4IobDuFhqgYuw34V5O
xqp95QHoF+1+WqdFBLWCQCfQmhemHxc/oQ5OCnsfmQnKzTd8RapC9mihIZv5NyEPGWu2IOv1btvX
JWPojOZAw2CgRyyAsE0VVTG2cYZrVYqaE8a1EiFkLBiDBIvC5+Bnto42Fm5dhHBxV8L1cnkpPjMK
MGJIvhUcQ339e8MH7b/nGnyy+wJai1rHo23J/saAfrXWafBoi3dRvW7BgQgmiH1AizW9OJpE4v5J
txqdkgkIXSr2hY3nB0klLRpqgGwuOzU9tt9N9urmXiVq4GauztRPvquUyt/LAa6i1uhdMiO3Bvsn
M3wro7ftDI+n3qSPCq79f5i4MjwogOWZmuxXa33Vg2/XnE9hrBoenYE2nHaqXl2skHzcdGXULI/K
edYwHA5SAdlS/HdnMTt9xixkzNMMdp2zByOyob4t0uh5D8U2V8Bq7yJwRGcm1wzlzq8NTRewDmmw
s86Jqxyt7SMYnqDrd4VhrCqhWNybr7bm6FjumGPaR1+vr38TL3LCbKyrp6K33G7RRDcXavjaT7Fc
J7G4kK9JFX7/OAgcm1I15UthgRNsIVaVvaFIkIl8D7DgViX9oKyCtuaZhoF/1D72j/UsiY4qZQJ9
BMnPVfpc6eoaAxy9afiem9pVi0iCKkihwLyV6O9/JDDKRNZJ0TOlMOtrX/ScPHj1G6Y/U47diIAN
pnyyTYdDF3suHN6+uMPqvCSC9p/8UxeBVHyoFO/lwVyABUreC2IkLnzrT2jbtczsMVeZKZyZVWL2
6VlNau8lG/Il0y0eMTiSDNY4zijfnEYPGFPZNfYXGnIaOccaFPEBv7F++7TBhGvfn2nn4pB2WS2l
ETvy31UbFdS3Ay7gC1TxhN/IoMtHwCpjBtb1AG1mn22PTZzMa31k7fgFqkRMRBFYUPFqiq7iOIz+
A4bGNXVA84z/zHITAA666e2FwNiORs8yL6w0WwBcIuPsGwxf08WC5dzlV1af/k+WehTe9Y+EIU3p
fb8Fr17aRBxJg5qIgcZRLqv+YtFlkgCTw1yrTykPfOZH/yJxu9bwTvZK7wE5MwFnSbne3CKJbCXv
baFW0+zYaQjDbL50x9b7AJ36q7C/rdkf9qZk0f/vPsbmFnTx1RsYey1JjexeJHAUcMLtaxoVBJ8V
bRlNjDsxb3p5NQYbmSo/rR/ZhVsYsFcBq7nT4R5JbtN5p8qWy5TVzcqEtG8W2Ic/oxvEULDT9tp3
ajcg8d4tRWzQwDCgFuE0V15FJYQsnJCGR01Q5wKBUOv02OriAtahFygXRCcWydllZudXis89ttxe
Zpm06DKFF03D/44b3aV3sQaSL6ecG7xCux5ZCAtMpBw6NaUGXDf3RV4ra6jG+vms/nH4QAM8SM9Z
hoe+5Xr+uKA58JcPlfONAPgFa6xAcvw4lYq/rRq/f0wh+cp6BzBvMTfuzm8vjjxrsE67ExWAgfDp
PUQ2IFLqIuvuQNi8AqXEco1yZcWErZ8IVZk8aHGjCrWrOpBKbLjkVT0K+MTKupGw1RsYA8Qx5QHp
mMldO7pVy7m5wlGezW8DCEuSt3TxajPaeJsGmNdgK9/jQ7RGo4aqXC+zUq+Z1oOkDzu9TxYAdyeD
IKsCDT5if9iYTFzriW7rAXSua24T6IyB5jMAtAS+MsLBqTPZPsUbBY+wh5n/bDPOCvbkrnNqdkUW
pRbtW+bIwwzFJybYIdH2lhx4PWK9ErR2WVjHrT8HkNbXxtXWBXlQrsPWklMTlGIcK4WL5OKkxAj1
4IXe8cURuWV/0UaUMj+0Z5sjOKygIjZlmLLzzAXoPpfGohX0WIckuCgOR08d9oY3Z5HKIdvEiAtr
erqoh2V78BSh1/Oxi4+0WpSA3dwk9FW4GZp3NmisplKyh8LuEBqi4roTy7XeXZ1dG0ECAeeDGrOq
iFjO0aeRT5jmZC1ZohAbwefVJqDJKwKe/5RsYn31577apska0GeiTBrVAHmLFEr5QvG8ZI00bWy+
BycSgUIzFwAtPc1pFkW5ce6WBhDQOOFMcmsTESPXJpvBvHZzKyMqdUobx4mm7gK/SbH7DZ9fqEqA
GZCE9Y7ZXezbsthup6yxCRhaehSFG5O4I9m3PB2bQQ2bmdTOkZWOpIs5AwoJjR8ENo74FbkL6SCW
mh4sJ9WKDNII1HQvPPjT/GAju0MEqft2CKS4twwIuofWFGkPbTRRoarEgAUH3B+nXS5SJoyUi/WJ
45Pr3/iHQLg/DO9pHe+5/zhIdemSkqKcd2twuZxtEmeJSwncm55jBjD4GBavW/GXbgVyycUmWmIe
detcLIwoTIcdlRoSKjNQ9psny94TKMVxT7E5o/26UZ1XXl6Ag8faBIP8hdvGspWmZ5/JQCjpBJ6U
rhUGceh1au3Pjaj5zP3pAHRmAHJ4LMR4HEugNGqTLzgz+Glh1uPtwE+Gxomcn7hpk9c6IyUzGwHG
HmdzqtMKwxyYsJgbjS5GDeHT2gBqQP3fP9c0/55p2alhp/bwmcPXrcT6zxZ/ifiWIwsfH9PwhzHp
iAcrKw4fOZUSONj3BrcWQoF0bwGA+oy+1VC2zeLheVatWgJONVcjssfCaSWjLI/J1UT3y02oI3Ce
8EWqDjZN+QO13kLtT3IfBztobOyXuql1wpctYHlJ9+2p2amim0jUT1kgEReRMqXzJOxSvK37fGxj
qmMi01erBr04YuN0/A9y6FclTIMoHKiN17v7AJXfZSvbvyer06rOT+0x/9qNYkjD8aQ4o6+CcGqc
5ufOt05/4JURGnEyVNdHEDFI32vZNU8PwAnL7I8gBGUYvVsqTSTuehTkPjRMKDYikVHp5jrouc4D
+Q3z7mV+ohmwvcbEeky2wGQm71jFT4NLVasQw9mCMyWUDTxQ20geBp1YpyH4T81iueugMVo7ipZo
yJioXJd+WzLc392y1MMEZtknlWL/gFndtx5AjuXhau4e8ckBqhN3H0lWiaST11iwXFFXx4kJVp3Y
3o1dW4Ol/zwaR9WaxJ1NDZoXSj9N/5M27a1mhWOGIbswEXcqFEkx+fj2YJzHY5g2H++UCNt8ZUmC
1QJcj0oHCUYCQEBMcMNeaw3KOhpgnBJNZye3o8NzsqJPmZ5BpePwqj5dVO1NEBdG8kryuwoRg059
1soYT7JjaQRuVp3Ama7ufCeXA43E9KNBKSFgEahm32TmMLoY5K01WyGhNyaeYrsv2mLVEvgQv0S2
So8dBSlQAfO83LRc3KUd1iZDPvIt0oZ5Xfhfks4QAl7lAY12XOEHQFsf5W6IkoBCqQ8njF1fjgwY
VZ+8V+tAhajAlgfPlS+2Tbj+st+Mok3PFzCdx2iPjnCeVLZ1rekh4HWqumQEhCIipUbwrsruvdJf
zXmnVrWzIrcHmBqqcu6UjcI4kKN4638BsWShZ9Ia++A7u3SI7EpHVWspSarN7hQUXuHBDIEgsOEm
mMZ1QyJAfKNEvJe/LS43wETZPHVvD67nJ9gd71xx1nLl5Gx9H/Y3KaUwQyE9XXEMiJXzAM+cLL11
DoWL91IipS7VpsGe2CnlZg75MAvaUAON8lGodVew2agerM7UOnlKQRJCpHMfMli+mFgv2he3o4Vn
mJonuqBhT5bhOPrw6+bL/znMBEmnqoQtMEsXDkd5Do1vB8eWZlFC28KjDb5FYEMnwfuwVuT6zHQ6
XNWxdPPK/kbo6oDppznd9EgLmAPxH1R+e7oFkLo/iOPFQoO2vV4CEZ1fRvZydFEm+uccrUzDzT0S
C8TawAYWwkQ2tjda8kfOxFPp7coPCdyel3KkLbpOMaGLp0ktQozm9znSAM+/AXNQxpObq4nPdBch
UDWeG0izgyrrgrRAdheu036tLuMr2B//dwDG0UKcPJdZMW7/TPcDVGMX1T+d6jo0uP4BAn9cxxc1
0xzpVrALdpKrsS/X1MttH+Rec9666BV+91/nAXjbl+e2gHz/hhR+V+GJE8BmLLyGud1Df/YkIkZI
tosVza26puKI3draK/mJR/9pjV7CE/p+AlSypB+6c4+aWR44dYFzy4cU3Toihe43iLAJQBnUMmJv
7STQeInp0N67WKSoaElHKK73L7ybubnYJKa7Ao1MH4V3nG4LLgF562uNvJ9FG1dEeIGHBlxYVHr4
X/1S85EV5C8GF28l4tzzkum0NyKJF+dVHCUWenHBK9q9wigmSE8xpjf1n3HGQbEO495RK09OQpLA
24HKT7gd5NzRmzPLhA2YghkvyttZdZU6rqjtVC8UM3Y1kLOGIj9tMzfERRnCB0CjhcGGa6sr2WL8
glpBlFlKT4wtpPKP6T13OMF2yBPV2oyqq9RdRnwLqy0uYUdIAj5fgQ31Ni9Dx39giCwHjORRG1Gr
owOsXtMWzDTrNGAjy3M1XkUA8tFUhe1q/1bbE/uROZvE8VjOdZg8Mry5RIcR54khB5TyDaGyua4W
yumX/wt8zT9w6J1yM29EiKmArnYePGfXrO91k1vKlcCqfRyHYwumIoFYAYPfW7kE2v6ErIat+waS
S8POjB0QJ1bpf5psG/REB2nXhQHHlMT2Pw6DPgxP2YKDpU6h8NkjFfeglvFC+V5VdwqIkEtUVxBw
NCVgVo0eWhRzKfvko7wIAqRIcChM6GrWLvYi5pmYxRVaabgCON0M3A/RH86ccg8zlI1BhnK3zNJf
T5ynkeEOoFANuNS+2/Sv5Srie145qHPmEHV50ywgt6VXNE7ifbAktuDr9Rckmvx56lP9xuovlsq+
zsjesGzUthwWfP77l5zK1kPP9s3C3zFar4nSxcsQoDIX8/GhVuLeZsGQPAx3UceAdmuwTeu0EJft
Tn/BNVk7+edMQ/NHBP9BbcrnEUJ4AQHhh49s+FCEzXx+KYW8gIpWQnFCwYgVOoBZkEWdYhwDv2R4
3jdBnLzDmf0HRxx1xE+o7/VoeXAchUPikNbSXL3+mybAphgxHCUT/13qUeQ+4Q/ztLnMWxevxSNc
pZvKwrxR5hSWO8FJ2Z6g5ik+NcEWkdcWX/AxFJi+zv1HG92IDklAwPb5SFUcQAEwcqO0y70XTd2O
BGoYbBX6+wW+/xEFbT0+zNEMR882FRiJ3JXImT323HAgxm+djP7dqkoZC3TZCuSyyJXIoGvBxBa1
TXDdiHQhBGQ4mwsIOo+PhjPoTW9W1qDpzb9gi+vflo6aoZvHxCrTXhu1vN7zN6JUvkSX/BtFMXEN
jeScDPkgKXLkeQ8gj9WwfHIQtkR76lrkNH7UBVcN7adHuH4ZDC43dxZiORIjEhKM/ecB2jHGdAFC
mT0b9WwEBA0wfuRjb+KovcuLwov+lol1KXjPAUliGkp4yTxBl2PKQq416HguHVInfguFzgYAIHNc
Teet+b3gAAeyXmjdyrAAtEyQchRB1lQnPqxUD/E5GmiZeTYA95aczppfTEVuHnzYvoEZ3tveQ2O1
5MU3jyF+DPF9rjz2vPnxmU+on/FSmDnWOL/37EzA4xF4RRHjJfO+AQ/yjrGrvIcwu6Ch5lnZetJ2
rjRwqvZNsNr8pJX2Pdjhq7wymnJU4te/pTRbiUkbdooD7BSr3suKUR7OWR5EnbAOYAkwXVUEMVSt
llF0DJo8QmXm5yxXw/yZ2W5gDoxs9CrRVlsWyV4oyhP7TSP2HI5dEDHeQd/KfyFfMiKzay0xAtsI
zIFBE9Y93J4/kSQtGgdDaSm7PqRlRn8Z+3vqtOkl06EjUBhkcjELBZ5lT0eIRQOVHkOMpag0+3Wl
IcfBsDSxt8Wm9N+UbWGJye2AZ1K/OTekvl6SMh1YrcmSST/U8otm7aY8vTeovnTjsYW+wp+dYeon
FRjsfef2E5rU5zMVB0Qjv+hkMShtGzQCFVI2g8pyJe+l3J1vbQmtzGnbjIfV5e+cVi2CvayPUAyx
PSsXZ58slb3trZB1zmlaeT/lwPeteNdgHiKHMCNk54247l9ae+jeBqEYf+l7Q/ch4PvYNa5OONP/
NR3nSTnYMpgDgH55jgYEUAOHEEWpBJfCnxrmHw02MjIPXFkxy38V7JugyGzf+X0h/PZT5W4XOHbB
DV6V9FGq5UC1d21cDV/RJg/aKH+5HMJcE0Z0X7/DxLmKda0WjTbvYwU9eDa4EwpTZa+M8a0PNUta
HItb9PCzKgLU3BFswkqSJrfTbsyJ+Fog6lx6VFeEs065Oqznm+tRfzsDVxJQkCxuxkfoR3HEr1ij
G/dtaIgjPWak52OZWx2K78NvBP4a/9AuVMs7DeTKonwon8uevcYk9+P1v3NP8CTUcRvYxaHLpfDS
cREIxpJjiPQ76+z91KOZq5p4nAbaKZjMCN3whUNEYecCPu6vckY48rmIDyPmI/c2aNA3HKJ03UIN
9/FyLnxyn3kzcVYTGQuRfAqECfySFLv0+kwg0+qoPEx6JkO4zGQ9iBKr5NxwNdrwSCWmqn/VcFS+
OQ/dLVheYMNdWRiPL7G+MF2fDnPXj9OaaqzvGOiy2VJsbRmZnMjiawJpoBBo4++xi1p/VEKOUrDW
owLPfyXaoE+rv6zI2bDwogPpzMwaI/73Du85zpcXQ3i8MHuPn1e/D7Kg4rlOA8wi0LV1/ntqXrFb
bLebp85SUqipwW4MMeuicGk0xW891MbfvQ9pOoh038BVKBgkbTzCxIFXwuj+Lyap+2VAWtwDG841
Q289llk1dhzHCWeDp1HBqFp9LyVFfEHu0pe4fjFCY2djv9Mp+VZpPu/IBR3BT/LnSjwb3d9eMumE
rktKQ8tGwI9VQQ3PekenC3ERzOirrZkPu+mO1HSPODHp0EMqnzG9XydqG7E0oK0t9FatVT9ZxX5h
7TD0qV1mJXNoumdNAScnxNkLK7OtE8/v4pb3d1Evqyt+g/VkxP1em1/7uypxFLxqBYp+mm5xiYmS
D/+XA0V1jqFH3DNOW4+Aeq+f0q8DOXr+0q09rc2jsTx7s6ur+ulmx23UQOpYglffGHC7j7g4v1Xe
KopTl3OIYCBU/Ge01uqvtQLUy2YqFWMqzRGy3ejHqn9GxlASo4cBKjO+lzQLAmU2py7EmO6HTkD8
b3NKlp99IAmAXFYO0K+cTfGQYjqNA8K2NNnf9gZD/HxYAu4CvYay9fwnQHg49n90Y/QF2Ff47Dvy
BB+8JVutD2jNLqSJs+l2wQFjOdEOg9hWWFfrRjS8oJVUzpZ3CupYxnwJ8Clq+AHXHS+A1xDTpHuO
M1DmR4TtbqxkiZuz90ohyIb7SlM41CPwxDOt5PmGjwMzbLO6q1pkL2Iv+YU6I3hh9ksdWKmSMByW
Vv9Gl51TtoH2Xo9/jPpHWKm7PVwjsovUUW9ZkCbZQROJ8LLM/sBCxkO5aFykEq8Lv4gyedZcsV9C
DZfFi2kfXcySiDBHxWknYF56JHWQRX/DHbHnusc/qInw3iEFhj4LVUnMjo8BS5zI0IIxwk62YLct
LsQMb0cCCC/VXTmlCfp1mxqVb61gdOpkljnRGOHCoq5ULWxJeUObsBlrVZzTcCuUcv7Lvzts28uj
Xft65CdUZJvMogVc+gcP9Xd/7YzaRHQVOCuDsrngn9HkRJh7MvfHccOWgepCnTJUP1/hS6Uqxb1E
T2WNdqhueyZhjtnI6Z1Q1fElM8jAy9dq5bmyNQ7ZuRV6EznC9tTP4NGgWD9M7i/mKvejKTVfyTjY
iE/61ezhC0Z34mRLyrQwdgcsgSRItUT4+9FavKEQwnPEaziC61SJp9pGpWhm8BJR3yy/VCt0GHQS
UoxhBWRyKc0fgs+tAhdDfmwhDZj9ZfDnmHEtitgQNrzzPN2UsmznFQKINrnTm29/5pC7+bePWRPN
CpUCEi9liWmWCH9LfSVLdNnegOuDONSs5cUBfGPnX1zGJjSebPwP2LuWou3TyVvhXcKlLpis59Ul
CKus+lh4m1uQuufr5ju6Pv7rPx5xEf4U1ZwTHrpVP352JCzafh0GC3hZ0kT0DAQzeWHmIMfj+cYM
3bcfM/tK8QV3op1n2p3Z0BoXRWEfZHC8YsRwDjsqv22PQY1k+6mNPaZ//cfbA0Ois5PAUh4yu8HV
4LV5xbYPW83Bhkqk4jUUndhZAwwlxrSL7n0/Q2bQi9JxDkjZwucIxbLPqBzdyGSvQV+70/s2aF2X
jh+L9aFWgVjLACeXPgrFBGQU6s1Lb1JSlJGzq2PI3AsYsnfyEalyZZ9yq7eC7Mi/3Qb2oG9LWVFb
B/z49XZM1w9e1KH4bWFXTok0Q/h8aN+ZV2i6Y2V7+LP1ugu/TdabgiuV+r5xwCgxunqHqiZ5iJji
5nygADT3RB3gmKdaqfmaWuR+/oBzy4pMFxjOgYemmcjUKH85tYZntsNKO9IvJYzzamMhwggB0zD7
yf4rMeqOtFQhspWFjm7mKJ7kpckJ+9nuLTgfrkvwY5jhVvBOrg2TiLcCpcXs5rKvOgOIwlIsR5I/
hS+mxjvcKfKgx+aRaRQ8oy/WEatBCMMUeIMon1NSA5gXuQCx0Dz7GN2n8ukniqKfmbJvGuDabIWZ
MPpvJVvMrN8v5Te/4ASqbnydVeFUzC2fQqG61KJNOGcMub9XO7lJSTfduDqIlG/Z+VhtUAf1jljf
oe7eBnJEMgexJ8WTlkVkqlUFGH6WaD3yQhJbulthiw/hlOCDtzw+oWId4JhpCtono7G23r4zLBIK
Guj1qfELoraY2yWkfl2B/Q1gs+2kAdU1y3COB2V+eDl8czub/UYCqJ4vvhFjb4OHIsw3m9sy/nJD
8uOC+ioJDqHamOUIosTBYArxV5K0fdOOvfPxIbtq/O2mQ4YN1bDa0C+7apxJ258G35ShbdFCtPvW
mqe0k53jCDSNo9kAG2lmyXZazTlQvQj+qY/RUVaJBhNh1AS5M/w9XPSEzqdgORfu2fvMEATx4FG2
WzhinpJR0ap5MtTtKE45GFLAiHQUgSvPCt1LNNcIKJEuzE79Pw/iSFXLUHEljoizT+htCLTPAqs+
ecw7El6WkjpWJS9qQ++790ulBq6tgBMrxQRRpzNZUDoClhMbUNS7eoszeteU5HjyOOOUm8rz61+P
JErwNefhNSuncwZiiXyJ3tsQyXt59WIIw+R+O35T/8/g7BAQtcpYVacEfMFGnqnjQ+VPujZKjndm
4nFrbZcIyfJNf4Mml0l4gn1+nqYU6KAwNU0XZ+HPzJzJBiWLXWY2C7UnDt5g73BVMcVJBwCLYgPs
sEZPwfDZ4/ieZtzGwXIpM9UyWS0UczwD3EdrDS9IGgALCHtwyAOMUDZlgijrr8dUtqOuOa7Tsrl7
euXBG9y0AXSJo6r8IL+al+IDTKDaiH1UramOs+DUM9yliFt1yStibrDj7bKVk+nL033yvVm4M4hv
fyi130DiCWjLGh6GbBLqb5dmrNPgyko63X0iSP5iNZ2lt4/DesbOyQMFndaMNFC8gdeAb6zrP0Bb
H64AF1qKIAubUa/gseQBd7cmY0oWrZJQCKBPEKp4QYeE4Wm7XKtyjuG3eVocFXt7V7pazvzgwGkg
cCVY7IPzF4Cw2eegarr/icUUlAbqWK0QWNqtS+QrMZw0hmT1UO3Q+XW+MPTcbLps+UH0E9FRJnPD
1OuQFTMn0KvvJdXx5O7hfV5YdXyB0aUvHscr+5a+yI3bb6SpEAa47DyleostXNvYLvjjZtzsTMs/
bKj+2lg8ha3aYC+Gy+STlOpWn8+m9P7hu5ZuDSZsuT6n4LUUk+Y5CcgGb1YvM111NrrPLxuF7hZe
oldRX6sOEPsM+SUB3mOnAa7Z11pr+ldDsw6fgd8knpNuoUHDih8xX8R6Y5sRHtExMsOFcHjJvr8F
PiEeUfadyO268JzV4PNfqRysBx/TFenss6pXQ7d7nKfEcit57AcnkxOdpjdMvPjhHIfZligYP3Vg
q0EQV+/ugEnsUnTIVARDGYiCUhSKgigqzWKG3tTT6qyqB30uv2bWi2iYZp5lzFRLvFh6mQs8fVD3
BaLZiD0ZYPNxCwJWqaIXf9TnLwMEBWgRnTV0nWTeeT6u9Clhtu2WF0ZrUeQXrrdsUIbVuxSIdcWi
BK2SOaa0ZczjCcsv3TbNf1ZQJpxwIbXmseW+tIgHB37zhX+kwaxlzPyNlclA2cQWyJxGosrxr9Xv
4pVw9kyNgpmSNFo+QAQVUvVNSNQaF1S4BUwhZ2uim9+9QeEgXGXq/GuqONjphezbj9cwgzLVbSl/
eahoX7GtvXJxdjUEZ/LozLQKi1Q9wwokTNsDDxFaF9AWidYC1bLBy4u4NVXqQLyvdN8fKDpfh5if
0RDxjf1FRlUazuVq8XmOh8PBTiGTN3JS2bKOKgo13B8M41fQFXN1977JgOlQ9V7wJOUPwlZzDChw
eGDo5GzfwK9GWlxbSuBhopCiYN0tRzFfmL0zlksgG/LxfPv06HvJ/RDxinANP6Xmhnc4LlXZ+gu7
l944WQiLcL+Zwv7FLsP0GLZuoVKkJux6eVrXwWN3wNUWoZ0AJToERfGT9V2hiI1avpyNk2D331rh
J8Aog9ntja6kDs0SlWEROnF/TksIj1HmHymJqxEs1bB24JsFN7iwty02fL1JQcaVeeeC0vpLDPBF
79xWeUaeFMAPvmB3epVpUk8P1TxGQIvv7Wac3sCpVmhhJxnUtDdfFWXkJRo1Gaqf44EnaeO0fntS
02ujJLEqePlgG6CrHItHL2DgmvOUpONlGJGypCdbn2Mq4XZgY0sVRR9UtLapox5pOoMao3hwnjdk
Cf/zl52e1Ikj/W8iR07nZrQbQGWQ8gkM5GeiOmLCQM7NFFSQFIbRnk25/TcmjKPp0i29Nc+FFEzb
cSI0LXKZa3cxYPqsZxNioE6t1RGqUEKDNFIVXFqpZxWQACo18VOB5x8Gy0umBOwa93FGyi5ASKzj
FaQq76h4Frake+ETlzJ8byH/KVUFdUfESIwASNi7ZwaMwA85FwrVK97gLFag+V7NHP59RzZOTNJ/
UREm3Q02o5bJkJSmH9k924Dxt7mrpIvSadDqwp00K2QamuoqWC/EjSSXMXWeb1joI5cEwMI7XENE
LLx7LuFFSPNiS41AlX4RmahvGxQ4TqFXlgr2JaqvMBWzwbpPig2JBk8lqQ8Iu9zNdqio35WPt3qs
y2khi1zqWd6pZt2jMA5IKkpZbu3AuTVVBqh9DfmoQV9W4ptrHaAxugR3YFHzDW1wd84ZHX0tcvcs
F548qoRJF2iSMrkz3spywoTzSThUwZWhpMSLdAM3pp6nHdZDlChfvqIEh1N42S0qLwh34Do0vO8k
o+3XzlkFM//ay/ABvFSvmuNUgEjo5zdQWpnoMTzl4QL6jWGQRFmVKG8Atib7TEgWV/WrD391tiC5
ZVmnNVjcutaycNNQ6WKJo+uQbrYvxdUjxw0GEZDHLhtWaWr5XeMNngU0a/IDSnAQiUn5IMwBZf72
YiZFyfqPfNOd01rdrmAXEm4E5eP9AIheAjZC3Y9vd3i24aRnCa+VnH2Zlqc/woGnj+krBd07ecO3
yTb4A6gity/GWvuLTkFfKTnYLtxyL0uUZvQWzPWycuR4W+T7jolTG1WKpVCC2dhMkevWxHNzGJyx
2rNdjYMf24Hsk6GxkoZul7XTBWnfZFZAyr9KYonlewREu7fxdIT23/ady+G+2ea6O/5d3GGQTpib
hhShq5pc3lxDGhTyi2LOqhrFw/OKcYEcYARzGfor7XR68h5vOKBDiukc8TgqQGTUkKnbTs6iMRPW
ByKhrKISg2JKBO30axnImnWjlOSDtBtnbgGDOU8j3Z6wTqWMSDllijZXMlxL8XczLtOIpxXB4zSz
B2rWkmgaVYX3Pr0c+ywY/2IbAajvv/8tppNbKLy5r6Qk+H/IT3EtwGc0iXssOXGIM4hrqVVJIz8k
juKio8NeqFQak8ZO/1DU0wxevD1qH9P/CAMUqIeh8YUXvBCYOQBs8+0IHhS9zJlNVHfcqQKm/Zqz
erP/DcuSRAsfAKvMq9AkOWYG9cfSDaKPlZZcPDUkEzXcYDugM5TyygprsmP6Uha69nT/yvw+kEGn
nj8inZY1pqeMXxIe9GXVLdszjOSxDucrlGJgYprBqqd8gzDlxV8t6fJsUGLwXJvOp4Wudevx2geD
x5ZEL3Ks2eklJw5aMkLzg/vrAQU6wbmLcwbsIrQ5rdOtSnJuBrt3zJcJr/5q8Q2Tb+IGUvhkBztL
Z0Q9wekqOqYl1GawYb8Sbvqa2BIRRRiMTBadYI0QrF1N/a2mhTsUplABmI056tkV9APrJR2BVJ0g
PJPOHqkhfTuwMw5O54zgOzayznw4xQujj3hyXvwYus0/YHpVrirp61o5TypUBDfQAJKxvYKvZkg/
VpFROT1yB4n4bxYSAAzbwe1FZvn/MBNU/lIYxphNVE8MjTo6QaJCyEv2XHB90M5vK3YGmGF58olZ
+3BwETWUDotERUMsYeluz2WElsJWIz0laHWNBSJR5lu1op1/61yHjI+649Uu/43OuxkS17nJLWW3
iYHhPzhqQB88YAK4RIuhCZr7ySCqllHjAUENOTcGAPnhdMN60zjfjR5q+GzIuMq0zIJLnqVeIWnB
Cmj8xYiN2XDk6xLLbC8P+ml/3O/qQXy/oGneKpN2ikDpAjkQTfbBeoYJfb0Bwl2y4JV6ssQO1vY6
Nt7tf9Vf9tCdTDKfqi8ZQlXq2TS3ZJl9iAUyrDtPdwIthmPFxhmTsr0K9Xkhpcy2/xLkxc9/5zed
YeqOVTBI5aki9VP1w2xaDRE+Oc1cuHr5EFNWTtNAPC2/sluWhih/tc6zZKmXoNT6mZv+IGvf613F
UYwrrWlkCze6xrMPXmaY/w5j6WaWf70FZfZrCKZJFOv2dwuRaJY1Oh3UWS0DwPmGT6HYoLXKOTBC
W+M1CkKaF2xiI2sdflOGOlWANaL2DwHzM65pfl13nArZJ6isGGDpC12+hvWTFjwYnX5gQ2GOBE5G
EjpoZCf9oKJjyDTKpR3PFC4wGBTGcdvgsDrWf6gstA1iWm9PT6JBYCw2RuR92Z+dCIsGXZ2NsUSN
uf+wN+o88S/Lu7U+zoKonSZMYec36Y9nM1X+toUKWb8G2kMbqwnnpEo1sD7TrD4LP1gn9vM3wHYj
y7W0G0phTq9uw7a+F/3NHqccUiRkF50kAEC1TyQrMvVy+KmXvRRZqZLu5aCVPHvbigO14VLjR226
JvNqlD4+VUyEnLjv9dK+Ojc3YoYYZV2NE6Pf/Z6ISkXtIO4R2tx1NK+Y2ykeevg2JgKyrIQK9jNB
lokx0wiAuLPa/AuTMCtG5+6Z3E/hRGqOfAl2UumoiBe4nehvsQ1LHI/k48Unq19gmsTlU8LPwzRz
38FV9TnXNeEkQBxDKC1I0RucQC8wC1BBRs+Qc+iG8mr2WO3MPplKthpYbY64Gi/D730OxPYcdUyv
Gc54WjHVdnf7dvrm72vWFNETO/FySKzY5oiHh4kSJTnGgEa5hTMcvRfyPoU/y8fegFSaiJc+3WZE
Ic7PzaKI1RIaF09jQOh1NcOhxGPr7EDxoQoY25bcrEWLlUlo2FIMVatWaBwf76A22xakW0Ez7LLA
xnZwIDX6iqIaDkRuhD+F0PP7fiiWnyQ9i8YxjPeCoq/Ed0PTuCgZKfnb+XSjjfXjL2zZ6ZFsRhTy
5mpKXBeEW+2Zh/3chBqQQPcjfNcPawIjJltfHuD/chcxXIpXvEPUxWJXpO1E7rMp4FIiGbjHSfgB
5XqAKSU0Z6QzV2r6K3BZG1vdiSAFTQmKm8MCblUyUdz8ZC0YlH/gnSB0sZriQ8ISLtNZ8hLwZjec
xixUBi6QONn5lwGr2uyzOiYZuOurPohLX28XlTMpin5Mpj6QUgGKV5al35dN12EY+ZhNPMY4w9Lz
tYI2uDtP5frDdP+rhtlNt3W1AWn+bidSwiFUSHsy+npLbhdeInoVhLycVp4IeavtU9eZsB4KFxXy
vt3jB1195fYscSAHIDKiz0gC7NiCB1PC+xrBxG5+ZezNxsIqO/5jL4SFoKKkyt6Vq55AquKcWx+w
q4WWmNwbdAx7BH0Mn5+ssH023RnALa27pB8NIWw7Z1m7GDRbxb6WKI1QYSJxYhxe0tYSBJ7b7frw
xpjLC2p3qyBAozy3Jd7OUY9uKybhGSKL0x3liWYyWi1cxcFCC1ijiwA2LCS07ph2plixBcIdUr7X
Tvee+HvyVgsOhRWEPqHLCkDBfG6HGkoPBNZdp63rh0OJ8komfn9GzbMiRkAj2ZDYfFL4FgijNa8o
Hj3wOxxZh0S1IMSbIZ1Lw8KuZ1OyOQxnSJQEJvKVtX14+xycT1FhwLhRwaAYo3INiS0rwYxxF8yb
ZQqiaLcW1joBJRk3/i+O+VYbd4C827pNEo85cJKRIRXStb4uOves3J2z7Xl0Cuw6ukd+xB7rOYUf
3IBz33m1RldKyrWO0L41zmN9HN+RUsde/z9tnEPVcomGNJE+KqtfIx3R46pyB7dRVNJ98CExm+pH
RWrfxbG9pRhEy2QO58F3NjVbPkzhLbgiQgvHYoyOSjMY7b78cfZM7a/FyHAMmJ7gGNKiPL3bM5Pp
WB5dtPWuZUOyMDzWcqYx1AzTIvFOSi4H8Kr5WfovCf1Li6zXIKB43nrDlWeVLMjQtlGAYNsv8XRo
bZ2msNJh+2gCTn0jhnmZfQFbuw6nGPjVW04+wiWf67RWKbY5orKSwCpGR+ITfTUiSBv8u3ZONvI1
dJKRkeqHpn4yLjfuJkoEYsw/YetkuuxDW9tidqdb5PdPL7VGtAstWewJKc6FXeMFMv7lUfh9J7MJ
lwsi9+wgstnjhRYJrkuV+uXufpYBReUXKKqfYW8ik80Q16ZLN5Wd0zx+1fBh9AfqR+plmn/ylNyG
m4LXzH3Bx7ZVYQentZazVep2rBYuTbaety1J61yobSA4va0SLVY2H+grdtDbzueTrdJTeVFZuyGF
fbw4fiVh/Wv13J74HYuk5yu8NzybV/kLGocGxXibjjce2nIOIEbsZIwQEdaFC6xsS9E6ZUJv4MlN
9QbK7EgVJc11RFFGg6W4aFa8RkHG3p8/IjpoQuyjw1MnNd3CJybGTRHkDZRiPn2RrYzfLzqSgXNm
m5T5KT8z8lb9McCMd6m5KSvMxGul7ZrmxBWvElkH9ZpAZghSYlp3MI7azvllIiOdjZ1TjOzaKA5i
ZUNaiEKtR9dFnO5NEiyWumG9koZWZe9gHQKOiz8RQ/fugVR61qC/D2C2jp1+jvvqsOIG6L1di3ri
icWIeEaaBwSMtTI4BEw+wM8S0Bg2s8sy1WjhbEvtAyHZGXczpFHxu9gFvAcyTmQ32RluJ4jjQUeM
weWTKIYmWnlwyAujEoJJP0fQmCntZxipYiTv3AkUubJmeYCvWMoH8S7uoDkDMV3eOcA1U+p6ejOv
1WAkuVUgkHLySJTNHVkQgRleoQUlBGbXeBUS6R0xcRpQJB2Pp5nCROu+98HTZB3ZISpQWHjHK6JH
34o5x4hUISmQjWZublTBiNOtdelFs+Ng6n0U/TAFx1SD22vY2W+YsYcPWnIRChfglRaC6lnCFe/j
lQXDiuZ/4+4mnKBJHP7nhpOxkt0x1bas/k+7WMdvFvuZWWT/l2Ai29NjCmcXpSOgC8FYlRLYoDwD
PGaekCERgBjllt/Wmi5njwGHsBoFUoBk0ztAd9wvk5/kvnE12SakH6Om5pSv8WdfZPnS5AHHM3FV
rlt/uhvLVTQEzDMox697HQbYsANUPWpZWWZP5WFFL+c6SErBW6shDuCMcPFDu7h13H+stfI4r0zw
iE982ZQJq+oo+AEKlcd+eWtgyZWpQXWKzQHK8JjGhTy1KJo+kIXPn9QaeeWDMmA9fPNgACnhy4A4
s7cNdiihcf84kSWSyzCpgB+6H4J4+bbArWQI2QOUGc6WdMb5gg89LjaXgfnzoIVAUnHZr+l3qku0
6D1FW9Ce7FMHIDwEgcliaTdaBw3x8VDq81NA5+wNY12Qg0ZvRYHEggGBEDv0O0VwWPdEZfabtMCY
P69NejLbZklAKrcqnKsHiVNurG53B8jRVd/L/WbYHFMnMkTemPMzXC130XaB+E7yBSC6t3ru0C4u
Y/+cXXtaQy/YlaSEXTiY3BVfvDm4kfJwL3uWVdxsWgTRcOnJQ8OxlpTXMOcnvxjK/MaYGZ5/H1I6
Ihr/1UUv61yb9JYGF9HK8JWu23bUtwgE0fkr1Xo6On45+LAkjJFNfCjpTLKkEJjNeC7lKGsavP2K
iE+FEDA6CLTLV/Pu8ISlonclqi3/cvizedv1V9BCTnYpKHrYf1JvKGfwUnRaTjH++ngJUrWrR0Fg
mhVT6xOg9XHLvrhKF2HgJ5wVFNQPLZprQVFaD+GvcElLXmFiq/EWJkN47b8C+fev8dnyGCpAICl2
YvbzbPQhnZGs/2HDZLei792zBPG0dRjl11B5JAgulsGO0c0+L3pM2+ja5eWdlSF79oyJwbnP7Y7Q
8EsBR9SETIaVtAMNmCv6Eh0dB2pIouD016qK5NV+sovYypDZT8U63fvwpiPm3ZR2DCFSbbQzgQ3J
VibSxfvsS5uc00Y9C0xJJLG5P7ndHCzL6KixtPpCRn11XqhFEEZH8BadSOWkchAIqSuLuTrlCrAw
VnbZbEn05AeaQjaeFsodaSuXF8aWxIYYuO1GPyTceNYShNppYWVd5tnaL709TxP5T1yZC3jb1K5i
nO/KtGOMmwqcRA9RSgcJWmK1nlMwF1+SBVU+bPy4E3wm+hJ0gaFtnd2k9UGoJYT1GYQZRK/axU2O
8pwONFb98dfAL+4ApiW5l3/0/EfYl8unKG0v7GvTZ/AtGThO6WIU+dL109CsCxwic0/3wIL0Ew41
lklsapzUIONQ2JYHt90fRNJuaAdf4ejNoGU2HzI6npPXt+cpCYnhCHLbSM039IFxDZNKszyo1nsW
P43cY0SbFotj87yKqKesR/r/luIQNuPxFGJ+Tf4fqHOI2sKmqP8wz2kpuYx6TiuDIihySfCICn92
Lo7/w25yXu3mQ7mfRAPVT11fyu4nj3NZtZXQssFUPBdBiYHq5u8hWFT6kUnwpOlJAlzBELqUqpjw
5sA+GQd2UEf6NNJz8rRldpk2Apcq/DvltsKtPzFgqZAm/wjeBPpdaKlLv9XAo60PmQZuw4U/3t2L
6pitX03BN8H1Pm/O8VRwYrLcYdi9vviremAl1SlOrwmUeA+qpBl1dadlUYTGfJ+fk+TyD/j0uUm9
bczXX9/R7h2bPctppREOFkmLWzGLG15PuCTtwfiPCfF3hAcheq7iMiNpmxfXfTwanLxXpu5XdfVd
iq+Qd44gtTygzEu7t9JUTTBOYzlkM/6QHJYMlUH6ypo6Za12LD7EhRosNlhfwkNnzD76lhfLTX1H
ry8YWfuLiOA2c71SGUVpQ9iAddeodJa6R6+JwrScNmAZX8RAifVT2pawjswPDmzqW9wk/TpjIxD6
TxGL5G8giKlijwIP+y5iVtO9lfPUjCBYA1pqjTwi/jSM1QbwUqnlVsvneqHywLMoT9yFemgpRvVe
QszI+GqmW9pDl5DNQIGTzCIKXUX4FyPqIDmwkaliviT64MKEIjEnp+cX+ZudgtoDuJYg4D+Epw4J
NXF4qMfdexe+Ro/r99BpSgJJdOnDPEaw1hTm0Qv5d+sAs/PhzaGSwobdrM2IMjQEXk4qxJXlo0jO
biW2WGQLGnLGDhRt8SdoDSZRTCUN/loz8wAznyw+J+P2jU3y3fdYd+KXKgVFUaQp34GSYp7O6FoO
aCx5Bvo9QBYmLsXQrB38790Kpy781mydD/8gs0UC4eSEuaWFRNXrAwAbPX14T5QX1KrjktERGKNd
Zbxk4+YLI2UWVxHgPf8MA/G1AHK40keDBewbXG2X+vhHmMosiwe49InuEtXq8O+dJfAuKYw6MuJw
ClFW+q8E5/avlQdtjmhFSljoHRGdsnMHTAs4ov5z6ogvYejU+kh+Ijqllf+X/tbOGB8uZ8e/M/CQ
rtf7K3i/FGD4NV3ckyHgOTjA8QCeKd3j5tT96J+TkGKNwzsVNPOoAnAGek7Klnw3cBcvtBI1inr1
GTgAqlwJpge6chS4hj6PGMhhb4NL6guyuqHaCuEoo1Lx+j2WFmqhXKnyqco2UjNzQJCYrunK0+LM
7nJW8DhGGBDRpvX8VfdN4UF09pwPP26rcLM1YZD/2FwTahScq1OZb9Xj8Pop7ONQP/tlXTtLHWbk
PartUWI6rxCZbUkLPwepXipWaxngEvP3Ypq1ZaOUBDnwi6SOOus0QQv+XCLMRxqk+fR/NJqZf/SC
6K+cIiBh1KORXpmZgXHaS4mvdsASOEVnDiNwZF4+FS62eAvRiF9BppmRg9Qdc5m3DahQeflGRNty
c5y9lZnfwnjT1CRII/L3bNutU1ox90xlCC2pmT/e4h3A+ths/UD7HT1KmaV8pCGpySe8lSfwsi6q
hFaASiSH+uasbT7mDh0P+sgp7uYoOrEcVlseVQ2vuN/vyPfVeFtE9WoRSeDm0tzEO2FSgnoQbvk2
7b6RvleP9RdQ2ZN/+5ylyB6iqfXCRl9u5FvxTQ31B+C1s/mFhOshG+180dUf8HDs7FPrP6UzGHGn
M3eIhXLBXj5NRBXsyfwvOcysrk8CI0o4yPK3kQqFiPr5ZULkJ1qch9Kv1bAabmIKhasF4sOGu7yt
1RJOlKgRGOSPQR9jMGA2DCdcmu3dlpWU/78GWvVlML+dZeGbfEn9KBxaBk0L35THGjAdAX/rSyrs
sutYlVure3HRRRTweQ70rbaRsL//oxSAJMuNTTjwwgBTh0wOf8w8xdPvLdSkWRqd/Lir9DvvsKtu
I0DQzXVYb0Yd8MyrNxQkhikKKslX++NjrQ9HUSrMV+VmCM5gXS5pbLrQQ/BytKXoVCyQSUx8cOEC
7xkZ7E4ZLmIQ+ZC/U6eu2NQx4PCMjxLtoENV7rVEkI2N9UEHm/AFfOuHhE+XL4p6Cr2vrwGnFpAf
Yhp2OctEEx5Q7lZP4MptZ5U7E2jJMozDSjizzCgYj28ixRWjna+tYGaRDW7vbm02YfXHaicj2dA9
cwVfEUDQDElkm0EBK4LO9NYv13DeAnoUEG/5sZVyhzDCIGS8jqdxIR+w34ZC7/IdGkP9BmbgJO6h
5wwn8LiUNOS+eDRt8E32sRjZ/cHn8BsORbFTwFcSavBQLEz4bkSHTjzWvZUhGtwDlLQflesTvPMG
/OMC6dCBFu4daVkPvXxMCnA3ddh6GhgakPutF2Dc/z9vo0Lco00cX3R3IlASR+wjlXDrfZUT2guI
8RaS+ble4uhnUqY/6bAUj6Koe4smJAV/L8VoMVqcxO4ldXGayT/3pyoYUHiE4c4mED1XygjAwOBL
K9GjvXa0eJS982Ty6XVP5hygMsEiAKkO33lLpJeZiVGUOJUaIaepiyhW+5v9mPw8qEWJxmOwlzcF
8OnXemd33SGKGFCI6SpmdwsHtyEheCtbPIpUmSQgBjlJoyXoC92RPElDbMfIj9k9QOQG1sCrIU7C
BhCjVzzOH0uxlJ70Bl03UCLcRvOKd3BX/bTn9a7ztYQjuNoVuhICmKECQ47o7ly3L3OzNC8Rz040
Cj15XC4oQvHojHX2OCacHbxol8noVFJDUQfPU9G2UrVSp+XN1hiex2rXCSl4j225tpObemRcrUBr
sBH/Fw58dokdRjjo2YJQlu+m7RxT8Ob+wXTqM9p6xOG+JfHjX1m+cwOI5eiEltX6SzryiPYx5TnL
PK2h16uay+1ceeLsiZGabRsy7okblIXK1X2YNRh/7fBjWZmUVjaZOsWsr5pkpJscwoHFArnD8AT7
jP/iHQgCSFiW/53ZX/51TEz0hNGzoOlWIpZ+wb6muKjgXXYB1SJHxtUeFudlLBxqH/NUVcKqx8S5
S+lMjw6v0AeaV+9hrOXfaIJWg5g6/tv90kGG9OmrMOgLn0k27+TmpDf68hFQSGeg27rN7lHryIvt
VZeIizZUbnAgLNECZBEhgN1UAGxhOAXE9BBAoJ5hYKP6/gMP/aJWP6Ctle3OedkrwJdVQ4eYsaOw
H8pXGL9y5ShNbXT40ckTtlpQSXWIEX8TxvkTrNeHsB0yA8uqiZwM0JAekKZ88u4A8ULgvNR1Uahh
mA1peXIi44Zg+ZoZkHmfKXOvNuwGeW6ioCIS3qClpj7kqSV5aFKNrGIQd/9Qex8fQGFYClFozXsZ
0fcEh0lced3fUDthWNZYevY4c84SdOpT4+CIECHMR7I9ocuLDa1y8x2W4R5gXCta/XQjtvIJ5WBU
O/gl6YtJEavwxTogd8HASHEThr4ITtLXDBmXAOt39rD5Edcs9ubqLcICEkTgLfQ+HDOiN12qqtPP
Cgs/EiJcen2YhhelQf4KGbkkY4F5DO0qQvNBAeHp9EIcyLU8ZxpLR75dtT4pSCnlmy/8gVrpAU2/
N5pkfavSBIQY3sOPD143n0EjaCUFi4CqRqo7PeHWue589kV2kAdEM8gMH+CTcE+v0Q9ilivx4EmK
h01Mw7rlbGu+kZlsL6hTY6V+8tplvSXGkXVwzVWbPOGNZgrwZm7bJdKm4fKbAJxph+5d2/mYAB5w
bYb3FDZhRDhZgQJB0CVjBXJPuXwAFFPG44KfYhQ+w9uUgysEVkUg2yKgLZsQfMjkethWANt3ple5
wo9T5kb94Wi2xcdTMocopZ+d2vaq3CaCYOaYj/GUyogZmd9tuESxNju8GTh2+0x1npZmy/WLB1p4
dMxwpXUrmGA6sx4j9wiJXXef7f57nffUJjeOhAUCQ9Rw/ZNuXVDBBTfFcvhn2ajGl+I7IW0IIuPX
ElYkJ5BQDffblp2Ff30AuVgnC+qCt57kO6rkkHUAHAE4gX9Q8G5wbLnU8A4iBZ/Bb4ilTHDNdVGT
dpvJb4wTUEmZwSEQv2lDrbDHt9z9vZ7KegDwX7FKE6cBXTxg+CsfuDXBTsROq9+7AUMC0+H9BD6p
nDqlB48bnZMnmTsmy6tAfLmKJYvJVpRPT/vAa1av2cse+w6EYZrs9F7vp+AvyacFXu28dGzGr0nL
+qEpQcB42LLxKCyk2FVI5fUf7aLwq6jBjc/clhqOefYF84Vl+p+7p+2xLpZ74RgXmHtyCTZXKGaU
Pc/uW7liUha+KZXbemXqb0Z4pSAT0XmN9hABtOW/2OvX/bwxt17ocpndw4MW2B4l2Y4m64Lkcoja
Org/1d4W00REswBTCbNeosT9LqC3iJhj/rEVrbjB+vyBbM/qLUgnK0uDrkCO9yv4QNPsnXGfNJbx
TfRDVP4UsVVHJnPBgQrBpSTp7Xy6KmTA4sxfDHIupmy4QL01EzMMNTj8rNxTJ28IIGMVZCSc+U2y
66MU5QgLgcf4PyhaII/lz+LnVd/VG/Ks1NvuQy+tBF9cyhTs9ShV0fZ5pA/MDTN/8JHXL0BWeg+F
s4xw/ZmXH3Hb5gfqwHJ2GNl2MlXsubyQGbEqMG0y+gX742QfgFNYNacqIQdVYAJAdObeual+MxBL
n5YdVC7PWvh8khh1tkhsAtDzaryQOyIrJaIfoYau6DU7FMaRy4uCEKNWLqybyLmo2fuiwX5zqQje
mazbqIfavLpFcoPdZrMhbdwqOtFkP+vfaSY3hEuiWjjeLuQBVMjKgRkfOZcT5DzV9clm4boWf0yr
YnOo3ss8IcVvth3qqjdvxhq/IyYGEjtlSof7NxNa9SB/yPI6flPAHhQLMKcQi3C9FDohQvKpfgbl
IexSWc+y9i1nygQmBh2BgQDOdGlDKkEvaeyzazfpXHjcz6mpwVrE/pm2tBBJIxbiGDmAWRG2jyIv
BYbODlyNgyUVu1EGaXLBG4JV997ZBuZA4LnYZb/xMZDU9twPHBpGaG8i43eH9riCTOq4cq7wHNgv
3sEulX1TP12dIcC8qlHU56iVWpCUQhHQ9hDmyFMKnowAX0MQHZ+14kYM/oO/h2zhiJEYBoTE0WCT
aXuYHTDaRdSp8pyseoPlBco4uwDF72fwnBCuHtN/Jw89jphk8pJQO6r66Pu21wXlbhGCGBPBv1Bv
fHNIzwZ2oLLYnhgrD5Ty8EmSM77uAfANlVVwe/8q+7UyYA077FYhuO7YtgIP2DG4zVkl9/KEA5/L
0YR4oZ7jcoeUqQH9wYLmCiVQjHHqEHwY+tt1WV8fu2HiDhflgp6BCb/b7qMXDClE0YmHwSY3Bmj0
yyEY4hfoDef9ZA+ORaMKINUTzqHGvWn09ZUT3YdeW9u5wEudqnW71c3hxDGtgwR2FAALIuQNRrmq
EZwEbyMCr9njcR9/CTD1ZM20Wh1vNwFPFeb0H3t9wr8lMdsxK047s1/2SgBrVDK4pr4YFIVI25qt
sWYJE0FkEUeP/FzucWiBga+RrSyD0Ea49s/Og3haUzz2GblnoF3AocJVnHuRP3nsx47FWcJgM/nT
BvEIzwGp8Ce/khy47zgoiN1OTG5iaHdRN3ohhGj4OTDIFFRzGRduWN3kE2OEV9eqOl2sUQW4FEJl
b1BDM5cYOuHzeRTNjhFopH61CfFqRMys1WhbJT9nZhwAevnDRgR5CktnnGJY0dBezKhHhEFOW6lW
SK0teqcSitrdD51EeITLwVQJp5wFqxq5SM07Rdkhl7PLv53o2lesX+QekeCWS/SJ89DQyXkRhyRu
LgVVtTYaIfer4Ra5dYr55ivxQ8IygeROhjiJZ6FYFND7QuOGB/64M+sbY3g+uDbVxxIHJTp52kBv
ARFAQS6o6LeNtGaU5syLZbWWzLQfr/Bv+v6zZ4A6nqiY3l5EGbKALfwsP0AdZlecBRJrjPSKAvB7
42fCoJBaUiERtXrQe3f4IGWeogKXbvewafghiuhaH15wCptLFmjcD9YFeHClqJSNwcHn7FzEgTCu
XaJSvahwHU0kXJ9caaL4g4pcPInF4qnDBucC2bypE6jAIdnOzY41rkVXnmYsjPtnKKtqoDDhvI+s
EXr4MdA4X1gejeCV6MLKbgIC4bfyRbscLV06xdOi7jF6aLoS/gWSONXUcrvWtHUe+WTaAU1H9FVi
q5pUnYmAJsxB5AZEPkXJe5+n0OIxKs452nwOOBq9VwMO+EcZS6/D+b1LendverKEFyHz3F617vrF
ZCgczU1mit7wu0qD4iju4dIqRCFc/iP24hYCjcGrETEN4hveZpQ/EHCoVnlJP0zvO34CORb/enDe
Lf7e0r9nXOufvzJMsxtjkn60uN8hpx/YZW0+0LM9Nx/ktJXsYN44TBBa6hTA0vN/Rxe2L+bMvGni
EnH0qKqTfrHmuYs9nl9zom8OftVu42FOaTwr9HbrLO2IhmCxJ8o+OnSzdF36aqJ/QcSJcn4kZeD8
MW/jTap5IlCaq4TdCin/GbXa+u/zTh+NixjtQfHFFBvGhWS790S/f1zI0qoQo9OGNMjLbxwhKj7A
XgBHl5dz/Dhuv8LQTiwC7Q+y8sZLabHnHFnOJ9PIAzZZCe+Mr498l9zPa+1R+x+UjOSo+Et05w5a
OtniVwMBmUgQm1m8yt0hjWzp9N10sBZoNYQ6kHsX2233d2Na133BbJ6XiESl968roM3IlZOnjPHo
tX53TD0OSjjNbJfbaMnIHRuYH9Bv9UKuTLxXlKVlXzT6rppS5g327LIXJsqF9ig3D51Uzc0L2POs
qszSGvdR/kN6qrXJ+8cslbJ9oPBtM+0+yXjk+RWrnD/EkqeRp3bqLArD/Y7BO2W6tw4rIUn6PrUj
2rhX+NPmWBZTEvLdQcm+k8Wr19ViWO9ktEJcqA044IqAHsL/Dh/r2FGTExVR9IEaUuG0XLD4Y6FJ
5vjmGHN0AS58VJjySy0mR70TS3e/cAp4JXgCknVqH+SnocPsofWMfzOCQo+G1/pALv1bSAbotbrj
xIuNSd0kPKluHuSk9iu1F9i2DExDe2c+PE//v2hqvzfkksXoqDb2vyjBNF71m2rREUKCaUCqZLrn
dqaNIfRRjt9BSc50zOVBZNIr7487yrBkywXJ7b57PzK1K9tgXDixQxDl5vLsbVUiYZEHY8GQZwtD
cNUSEFUluo8s8Xm2EydAzYZ7WKgUO/LEbZHsnRWIlNF1U9r0dA2bjn50xLzoSe+ffk3grmAdIa+G
xsLArbGW9I0JQWNF2wIYWidkrQWiLWOWGOAHxTbRSYTJpgqgRbQt38xo+KI6IyAYp347sLQ2V3Gr
PhOixZY97JwBSanixsuBBZOYMaZRP9IY52Yy3poJ7OwBM3e9y9SWOTry6+ndexneTgib1XxOdUNG
BsTi0AD09at9+VwJdxswFtXegxzTxEHicA1ONjbkNRpUCMwje2NJ+QEJnHAwuX9NISgxugJGjsOP
6ECWmAyoh19+EjgySGvm4wjzqOK0p+Z/ovAaboatOfpmEadOYkJ2dQbUdn2IZa0zgc6T9/S7k8oE
dftTIy7yxESwYoLyg1WGNoB3lHzZH8QTCJJYYYIWb78orlPU4mc6uRhr91INqGn7p81ZMFdj0zCB
6VKjxWzPSM7COxZ7a6i0A5X7m7U6s5lIgIw5MGmTyHz7Whr9HFIwV4eMhV21RoB4cBrkD+LVRyeL
ttYrA6uSF9IZh1QuPOGPDywZIL8hInlpm5dd1tPpibPIdsbGmWCZzEm8MUPIK9fyDA2wLCnUfCuI
pzMA7kSYC00GqKdhCbespkEDHuPJfRBBmCTWXx6djxR3rgb3WbfK91wVxnt1JDPOTTTifWxOEn56
fUIRDwdSWdhyACoO2NxG771cJHyFyphbGBioiNt1CQbwnlCDc0N2QcyU3TlnRg5q5SJbcVbJMoFi
VEiS7XHKvJppC86UrHXxLqEgK1fLvgGEOpa5qqZFtPvmA84t/x5RFE0DimPGnCNVr4hY9HibZImb
IIq6LCDi7P0K8gJuUY9OoMsyhXbUxibaUDZTjQiiAi8BNjkSFUuSQYCZtRX+79o61CW6aapXQml7
UWecSqg1VIJ+0KDXXiRpHXQ7zYQupsS8L3HGniRE+bdkZFhyrBDnfx8l54WQw+nrBJr6+m/2ZIxG
Ss7ZtDPcXDCmMDRjsjI9G35rWZuiYHy4M3wTkpj8+5NvYKwawv2EChyGWklgpMA0Px7yH6O5vDew
mo66jNFfrdIo3vVqq9lgvoNqZ0vbixgbWfUWgVz/QoYFZexZEr8vTsaIE46fuCXU/CkPwArH7KYO
Zb0nXf15c4gwoZ2RJYiqjdDCpA5mZbP9f8A0hYUG/JCBVrKMyhaYOcX2VUpicHLu2tHTP5yl77a7
8L16RuEua1t6kZswEcLj9yDT0V6iYECU3BQ1utSxaXYgBI71z7IqKMUVkiXCOLTBm5zO41eL4T+w
V1M9zjvQ2LOsLKdgODEg/7Ma7MiVZr7H01GonVnDpKQit+bKcBIveUeAgKFaVTAFIFXBeVotAVY3
lo6KTjD+U86mtsZovjKSSFrooE9wvdOB68dp/bTehRbHETD01LdLOlYfCUAaSl/reV5KAxm90L4Y
NC+lpcSavZu05oOArWdsRK3cnjXeNuelg9PveHDJyPvFp8I6Etj1IH8iuOP33KOBD6N9hD49/AtH
/KrKajPfJLHlCffLE0KY82kJ0SAMXjxDICzt86vdmcNGMtRkS7NGU2NXLXeYNG7R6LY21FVGd57U
sLUMiKxYPsN5J6s+99TAAgbrdNppKlZSbB/N051ukRBJod456JQqcdvaW/RxCvPb8bTX0j7Tm8Qf
wSEORkCERbEveAGCBBYhnhwATGvsWLaEUBsthV7DVHxh31/szY1gFBEXyByGqF2hzC3RVG7mir0Z
FaZaQQbIvBuS/xHDem47wfAfkdxV21qp1JlwzMSG7XcSQX1MWCAMT6HFgHTUMB5zgB8fBXoK4flX
T/tJeaz0/b5WmgUzwKn+ZzOO9ZeuLFZ/UkkAugey0BQXEZjnySGtz0Mc7FovKczTLXzZChb2Bkd8
I4HQ1yZT+bwYo8sDnu0KDM13srwzzSUWqrkG57L4EtXN1WVpLPPB5m/IWltMv4EvusNx8HUuvzIP
CR1c918QREF4+vy4odueim6BDmxsYn2oSoih4x6DvHSAMrlE4UYb37W9yZ2PUfDEtL1c/BxblD0R
0zr/lpt85LzvLtmRX9xLHMTtGtFZy5I1jSHpuwF03CBhnFawsiUeZHn5w9c9ZCg5M4ujjDlAj6Wy
QpdSLoyr63PR0wlSDVbHF8gK3yljgOhY+oxBnePPoWpXAP3ZR2hiRniJGRgl+Yey8e1Tll07lJo1
tN4PudSTNnVkpwOXatfm2izn9btNZ8l6dj231DOnHGAt7EJz8SBrvKtLV9Y7JVt1M+E5RpNHilTo
jYyaK5kErDCO5RXCUlinLQlAdBk1iXYKgspf3xCulS5TY8qWh/qM1B0kXRmusk10W2tSKf1Dd2pq
eStHGpeF6jdyEW8eNofr0L+aYr5opl6wEm3+KIA9xqc5r2wA4jM7wgyyVdXjesVObmaf6QHsFkFy
ZQIRPCJO4it8ZH56Ng9na7uYFx+1cl0CKUR6h88xgGr/HnejscSpTdmd60zNh9wG39/t8J2i/fZF
ysGWVy0FFuMJQELFtUgHxrwR3LxTnUZKMv8VAvrtuSQq650hT7bhIe5RFdU2Q3dRzlQ1fzU9CCeB
dKAOfhdNZLaR/DmBlkYtRHUxt0LVCQzeW9sveK1zbi+5zKCH/Vc2l6qw+ZamJAVW9cVO0zbP2EcS
9KSqNbNu0tTV8ZlT7fGdsPmPIzWIcig1upgoyxSke1kDcecY1+oB7wmGHLmY3CFjzWmxVJH1ddW+
MX5I6ilzXZvZVGDfESoVZGRqsq4mR+NZ2QGXUU7Hf+Ba/JevMCRlJqgwZWbPG1qLNsGGSCYdiS/8
euubVaLzNy1oqTTCQGPHB/u6OhrzISpVT69IHh9p2DbSeEo1BoONiTU79DoQ0fcBeTbF4b+AhOX2
Q3v/d1ndgVfqwrUOhaomqL+//k862Z5zvanPLamH9f8jnZhhKme2rROiuLpFlWQ6NCVURZed1Vyy
udW+hIcgDaPzNEu1vqaDQOW5ONrtckvS2e/Os8xQ3Hzb3M/ik7eNH7DptegWG6Obq9dwX1BcaP+J
+GkuFzJmqyrsC6Y/ZqSjJUBFKt1CgUk3aaxCHHifHnSWT7XeMaGYT5Wy6A6PyzGdnhqEez5JkBVS
FRjObETcJOmam9YTdHED59dzzwRDulNO8pjMnlASOpOkusThqYSe0kA8fQ3yry0/QOieOf9rkiCF
BYduHd3OnkvuoPrSzs7Rt3u6Q7t9UmP2Vve9hjPchcn0/P+lRXwaZtZEWojyyoVhIsJW2qVsjJ3I
STl3mRUqmZUY4PSGVP6WjscZWiFByQyws4uqCoj5BmE4kufMSgISZvUgu/cRz3LMu4dm1gJPQqRP
sxpaga2H3SwgCYCHAFnTGrfQFevugeGcOvTAvJAE6S2yUcOBltpiMMIKLptBPt0MKTRjTvxRCB9I
0TwwJ/dXns+T7hind85TgIUIL2boaykn+g3DPFBvwadBXNvjYF1otv6tpuHzx49xZ5NQ0haFID0P
c5KUiY49R/PMDnOPiCf/yS3XPEIabxQQR9rNFJ45zmJAdtVcWlz5/xzpnNvLWV9zCnc4fG4dL9zq
slIohRYb87stSBdgfAu4CdOnVlTrMKnv/ReoJhwHCkQCda7Fom9GFBHHSAbSAi1TlW7gbakSDPbw
R1TnRgPXAaJc/73sCl1ctE9qymCRPtzTv+VnLzXBr+QtcIYHd5YmrwAiSsdSznd+ytFSYDIrlGFo
GfPA1CBpWDBEl7AxQx2zszQ7gjb3S6NqcI/teiEdHA+w7asg+thgO+iPaX9FLbImwLXXTri2jExV
68CJ8fLUg6/Xp2eNVxqBO9bjKvtcaD88MWi3/VPmUFWUqYWswOjRpbrYaRA0IJPscrkTc6WLvXti
eAou9OO4USeaMNjqTdv5XdF+QCQyMWmQB0U6XpNqEmlvFNegAT5MFqECx7frm6E6ydNJ79F6uD/e
GnCevXU+7Xq+CZ2gp8jv8L0phz5LtPwTobjjV68kH4zPXuZD3MqTEKAUxRbRQ1fRJzd/0L3av2D2
gQN52pGktWEASeXXyubeeNkot7tyoZu4HxNpBrhH4w7zvycMlWAIC0ghCjcQ/3WhqBMJxyoYhMcr
vLM63v5BTxuOOYAwcl9fxaFUd55v7GsQwwOKb3x1OvJSHpypADVd80O96IJRQ1gcPECp2fc6ID2R
KHmKotsCgbBscqLSe6dw5MGkavVFdS9w+5JpYzqs9yjOJFA7xkqS1ZiuZELjuN4LTNjyFMD70jO+
mdB0zoy7dv85aPAdUfS56DQ6/VsB8P0YcFt7ObCrrJbFnZR4N54PqXaxWmzwtCFaWm+WC4Y8gtQp
JTxQarAA0P+OKGwjmNlxcnSI1RyanzGYdC58qRrQ2UyFrYOuY8nqJC06/LYzcioS5Ow0KACN1Ai6
OPCAwGWPx9APXz4zQzrIr8hct2xqUutH382VPlN4XVzXIgDmz2rqqaJXu3Mbm7rR+l/XGfXpVv1h
5jHKxtFx5AVJ7d8sLH/VQAWz1YDTSpWpfFiwr5JnIUY+zOf7/JguKqa3QK1Eoick/UlIxKiHawYb
dkr3G/tT8sziwHerlM2luceW3QTMbvPXcci6lUFPB4drzoGAftckoDMBxBMD0uCvYRNifR62AzQL
zwwc4CZbMWFfGKwH50Ln94QKXd2kANv/pHm1KVwHoTFVEzOlDZ840M3B0JG7xL1MYBmCmzmbtZ1j
Ga+BXZVaubj1NWhT1CXp1fft2rLMQTHrCtWq8Cz8ciZpbWNR8gNCf1zR1Avrwv1pcjgfbBxDTkwI
AUyz23g/ERSfXtoGlRKmmzKqDYr+eB/qM2jVv04160j+Dcg6R1DhZY1fEfLxpNTAQiry8qTiMVyW
zQtVkU3O7iRGi+RzCo3afkWfZpeKHiaKZgJBki3vLO3QywHSyQvTFJkMrqy7kxEjDodO1jyYzv/W
OY0MK251IuGTOLzHitC2otq4QPlzomp+FQoztWI22vBnIT5dOK57i+MxwdUyTuugM9D8Wd1dEZIL
9kJyP2xVsQaR2aC/N5ZKlm9YoE1CqGzPu/q9W6QtN+8ls5lRBx4cnOpgzzxotrXa14aziZD7V8TJ
OTmvP0VwBZ9/K1eyL+UN115qeeJFbQWnAOWfVBaltxLCVfcTPebTLU4iPb6prpUO4xq9r2PPrezV
WfY8qmjQDjCMS2z0rctKESH8lOfQlqNVrZUCV8ZGSSSfct5Q84GsqPIs+OBQYiL3xOJafGJBiJ2e
igeohrph/YZ3oWOcbPoMYgFamT31TS843iYtjpnhnSbZAngbMtY2auf3gsJUFd68SxsI/laZM7MI
tSuXlrC8rlDt3jSIOrfJQAWrJsEZ0+xweeDwsp1kGS276s4nHlPdJxEYSVWjDzPwu6/kmcmZSzAs
qjVhYzfMrtludS9p4nIsOb4OxZiKDQnO6NViFqm4GI8bm+YBvbqX9vfjmafD5uRf3l8nFStySc1U
uoObX31tRex9J3V8RNcvMEk9wfidSuh1lYV1vS8luHh1jONywWmrb5WNMGiUWPw/iVntgXgV5RDt
dL+MDQ9JlY9EcULFECV0+EQyW6yCOwvBehmi8hgjG3+8XUOI8acL72LIiRbEPcsOUMYIyyveEKVt
Ycnaqud8hpEelfBUxfmSfCAFdl69F2ZkjYqH44T05tKKyx4InbSE0cTWl+sIUszYuVDlxJMSaiEH
kNlfHzakBfe+UF8J0VS3e6yRUcgL+W+95nRegBs5UNwUHFaX6P1n7ZQ6up1aH5NxGHWYdicF4Ca/
DA+MiKGrT3NMGtwhR0OarN2zQOWKm55FJtcpWBShPtuzxTALe5OxNUe/kMbRgCvanu1QXqZAZnf7
tzgq7R7ceIW5VJTUn9wubR9FpmwTz8xrqvojRj1/yrKUhB020op+dsaq/VuXLZzWr/UKt9S1Zoow
F2TDv5Im92dXs4Grb/t6c0sv3MNkyOQjDydCQ0TuykLyqQtwDH3i7VouOrR3tMGWhEqqMecC1T4a
ZVBwSSixRWyuW8bJUMr6C1YfLCTAlz552LfklNhfrDuZbf6GPkRmzbyART2ub/BX0bGfOVRoNe0w
Oe6lXHxd0CA0N/jcXA6esQgrCXqKinnFoC0VtlVgk3p+7Q6NvPi7863f0tTkXBVg+Ta6LbnNO2+y
LnmuBDxLWDFFwODdhMJKIrlmXhHB6OfynIsYEtwd/ew8neiI6wmoyiz/OPJu45hqhS/ZC4q4AAaG
ixESUENzsVZiUbn+FIR9y2zIIH5K3oFZX7D6qfwZ99BE8DXoPOz/FLfMd5YfBysBLM+DMbqjAzzr
sAtRXjjpKPOTO8K/BKksl5K5PoYcoBH26OzgCBx7nUaNgTkMv6buG6S+gMmmH/arI+8D5vp/nBYb
sIUf4DA71/LhYEdPRmSX6D4vuHnSZQA03gIX6J+mbvBA2Ud1p9waRVOb+7QW11YjSUXXWhoLuHIF
Gx9B24Mjef/PDE6Ctg0/z1tPWZzYg8C7zkWdIzwOJI6ESpid+n2iA9aABAUcXK3JaqC3mejqim3Q
EvEMy/r23zilpxNCRnHd/srce6pvYK6r/fmrUOCg0hptVGogYCIb0K/P9PrCutFuCJo9PkzvfCEo
D3K8je6UabksM4nyJfbqzSesl7CJlJ+4l5u440+Nl/CHjxtwUdhIdiL8CV+qu6iHWJJVIZk2v4Xa
gVQKdcX2m8XmmKX95KXhe3XvuEAD+LA1Qepykj+VnZATVN+T7hDqvYLYnc/DNn1dr5xp0lJNTC7J
eF1aU1IgqilhG7HMedJ35U2XINtkmfAk/JHXvSyhorWL6C55+1/7FRWJk0SI6ORCSJ72EX4huaDu
hACLZwy+e4o/ESBw2fv8PdCqSO2pPaA6mbvjc6o4WwOJalxbKuwCRckPD55+yxXlJMoNmROWI85x
//DTEjJwTIeXqK2HBc1WL9W4I6CosZkoRWeVUBjDCFrjqX67XavPTlE9LCQT74JCcOu3p0yyfpgW
pwfcL6aKAFsNbWXcAmJ+AkUOHAspc5yDhEYd8kCkH8IKd24FRQkDfI6lfbiDE3MsbCq2uFKVAqEs
Hrol6p9IDS3vKms9zP8YXea6BHBxFq6UzQt4doKtYnIS8ACmLUdMtnfbqxaCzzAZAZ+eDe3HRUvX
WA2bJplX5J5QPlCjJ7pM7XJqXBeg0KAurgWZX19gev3lMl1S4YX5LbbO1xbP0/xqJdphq6aasJ1n
PfC32Nq0Mv/VIdDuAAqVYcIcJf2RTCcSAna2r+p0POIY9yc9y4Sh9TPu9TnmsHGj1cyYGfgyYYOK
IM8IPAEHrWvtZWpjVWcVLc1SF/uP9hoVNveix2zJAygnphooR0hJCsXOH67i4kB79rwMZy+o7LRR
G92UN2h5UVFRJDQPPGcq5xuxUxM7cRNIYrnXz3Q2sT8zcTEw84uaEqLGJ3IUXVCY/aGy6kvsJtDd
Zx9NX0KJO1/GBoEYErM0uKhLX+Thd2oYhb28QNG1VBy+T8z8mGVErEg50JCB23Xn9WYf8GBeDGfq
pCNDLieMnP3F380v8mWZP6zuWCswsLpnVDYQrVWLZOtCzp2xb7r3Eg85drjJW0RR0ebCURSdGmYb
cJha9l+KjEFRUu5hkotWNnmdVeUh5a3XTSzmmlTvBeetr2G6/ZdyNCnq4RjsJPlzoWGjKwlh7hMt
akf2tfYrjpVanHpIjqj/gS/xs1E/uhbh4kwzGVhFhgF/Fyh3Mh6xtr01rC4kpFChlhbWzcpf2Fci
2AEimOWPW38cvUuOtUeKtMKleCyxPwPh08ksYHK+EDQQB+AfjsT20nZaXMtLlESL/4umvh/Pwrm4
mGfrSqk0zfpv1s1AL29OX5y1oAIaXWcAj5KAWMG2jeJUlPJcGhOK6oczGo/U35viPQutkkd+ff7Q
Dl1BG/hrmzPkryeGoy7Pi7o8XzZX4IO7gm8Ze4w82eSP2gzVzH8em4vXZvZI6Hns6wnlVKBNabxi
8QUsfkVl3OlVRWjeQzrT9viw/Dzu+OUg+eIH5fWfUnBwtRSwqpqTXMVGYJu9Tu7WbuzYOci5kLGU
Abj85RGPHE/W7OsRj/IS3zOW0U7mYB1MISZD50PHF291H+5p8ujYBmwrpDZIKbYYjyYZTPl15Cpc
m9i3G1lY4c4Mi4JfqVZVb3vRb4nL1t9+oqxXxd4ZMrnbceIDnyZmq/kncLyomGlDR5u9YDwQXJBH
UOKY6ZVhEHxbIB7Gi6V+qKccd5ZsDsujsEMJkKilBGACDiGbNZVuleFTYUwWiVJPEaOReM0L00Uf
fPhH+iN5MJwx5VRtbxdrPK3bjlaMrfOA66uE07DbI9cEz0v+i6kDVqD1II3VjxUDKtOeN3/szCzl
082Ci4njWrhQBp8sD9ew8ufwp2JVxJJVNkSiTMy1qClXm0OVkFIP7sXSaD5lSCcT6gdBO1Rt4Zzj
+bo7wP8hy8q3i0M+EFc7lJDaue0McCeJHVRMpmOhcAKoX/L1Ws2inIiSuIDUZlEEl+3OhzPsG99g
851PGV5HBcpvcxOWc2sYdR1MKwn8C9FFQwC5NuNEvf+d5I8DHuuPNILLW/f8amsea7oCTp02qy5/
5u8HzDwf5cunwutyg77PRdzmhbwFbLfW/ZhQrU43rejAoFUk9Rc9fqw+SvcDtEXjjq1N6LzZVObD
VmMIibwGLbGJjatFsLMpbkx/zFJRi7T5IBnBqBvDPYrCH3OAbhMUgNBxtiWkD8MdBDOb+NVjeKDx
oj11VxO/vQRRKXVT6cLtl5uqzZD0ZNVuHTy673D5gdnulvUKIjLwCG5I0gy855hwIoRrdnIGo7UC
RmBy4XwDeDykuqZ9d9sDTPIs89D9sozCc22+0g6g0vv6WWyGcZn2uUKbaLAahPRyN7YPXapdT/mm
D4KBg1PWZU2AxvdFKKYLgnHc7+/R59POEkwwfqC5j/uG1d2Pyy7QGROw5go2UmP+Slet2q+dPfXy
+gGGzHVCrO0zG+WDISVVdQ+3qFB3mXQhVknxhiNMyUSCta2SQKa8J4HXVdJLXscWEdo5v45xI7uM
vKWOSO9pij7MlzRm6NuMmn9OZACRFtW4vF7Wi2iX14YXXOFoZOYEpcIBBwNw5CHZ3GxDRHg1SlQU
o3xQMv877bXOC+zmHtl97GwSFOWvPKDWT9EtUPhyv4zEE+hrl26BQ5fuTihFrb7QS1lIaHlIoB2d
pUt7Z4Pz9C0b0ANY1R6Th3HDqKleTztP3GmZld9hWV1bHbWOaq/OZxfTazp/l9LO2D6cgMV+a9x6
Cfn7yYNea3N8ibEIb6QsSl9K0WcYAnO1//EjECY2fmF0zu5ywYxIaqSixsdJU6hQXzFKBHwn7HtU
kyhDXHWhKtuSTfEciLvMDRb4JMv85xkj+aKG4Zm5TqaYuYbeUkHcCTwlnLHrCdndAcdZOkHkE8hP
gow6A12FM1yctLG3IS3zgWOnW958MYBuiVbLGdLCLIGuYtnJ2Wl1awgu4sueuvHhGegwn+m5YcV8
c1JOttFn4pG7fGX8g+n1gly2DlXrP1u4mfOTALeVxnb1nhedC/oCKnxeZEE1QDLW3xoVogAPMJuz
Fki2DL5KfqS1/erA2uzlhPIbQnY2oKNq9vwrshgSGJ5dFiJYQcFjvAjXvkNdLhc3/on/Q0i/oUwn
/TK6qcuKrwWE/bfsh9/JDbqqaIHfDj0aJbki2Coy9UH0RXFbIhwpKxVq77DckbcvSKeN15MWQXoq
wZRCKJNU7KJLE0yaC0cEhZhlI3YRjV0TQ8K31ohrFdwk9A/wngsDkx2ZpTG7I4ofyiIt47RrHml9
mQX2hhUA/17v3ZA8pCUMpe6Tn6CLiISUbPWhy0qPtKNJRI6R9rFE5AtGRFFAemCaMwX1tBdR5uAx
mlG18obTOBYvJMolk7o0MY8cbu1lKWCUnJbmYrSeKKzxvzQWHQSoqANctf0mXX1HaJ1l+jjfHOXp
1jzieNz+4KtzBI4ycWbkJmvxruqGVwe1kBC/SUGFn7UMHnCDgfI1X+hOxeX3I9CyA2ULMs4urJNh
VSNerVzuwstni+VyVqqE91J9JI6Ge73TANJhG3GooX1u5LumJr7ii79LxSjEvWCWlE0Qc5s9rSNy
awtQ+a48Nh3gHDW0ZkhRImc85FU/N7aLh9mk2fCVpm5e+GvPGsX8Zp+3p7UsMLd5h+ouHaGUEwnx
w6ilFYmBh6zFPQ27wnWFRCh8K764kvFaPIqMceP/TarqbO9/LHnpq0uhr85GFokv/CTc1LYpBVj/
dS6LPbvrGKYK0yPf7vJHfxmoqVKi11ljw3ZAcBkKBd7QNYYfxOCC99x8gvsvDc3rVa59JRAZUrEp
Kq3kWRhtzvqOlvLckZbs/IqSBB9/vwWhZgtT2ABXot4eQOQzSb6qZrA3Lh+UyB9vyyNxcy27An31
MVRYui6ef6fXf3cVs8v6jggGDosokBTqCKNeHFekZSerpA3prgRyTuzle0RI+b6XaZIedmp1/KT7
vIYuiCH5FOgWWpnuKz0HCsb3MbXNEelgY+NAxdCN/qOeiqT9gCrVPIjG+0SQBB2iVl6VR5kRCzw7
V/zTKGak1nLTRYQCWZNPEPCKFdkGEskaaGcYt5PjU8b+CgcRAJG6eU6uJzYFVCHmK8/OS1wr9RO4
H0km7IZnbHnIiRbwrhRh9ffnsNkVhB2ojxgEEjXnC+dAuYq5OsyFbR6rRUHGm6tGmjLydGtn6LZj
PEVwFAEEkpN8B11SSUvsFnDlB465X3U5W1UqrJFMvwKZZssmDegp/dg6wHQls/rdr5GxWADB2hFT
zRUgMmO84Mp/csNLlhyTCJihErruqH/HmHNvO8DmCyaYKL3cNlVTXhBG2klvwh2GdqT/ktzsEoH9
vNu7W90HgwE9I2Iumzduh++oknks1ZRXlq1/K0QTUwCp5Ceik5CU6cqJmp3SoZbdFHd6UPQas0aE
c0goeqDyKEkKkeXz0fQcyRDo7dvw85HjfmX2OR2i7wV5fJiL3DCnGmS6W89Z2f+2mDr4wx+MxgP+
p1fkcypNe3EXXBLfEV+U4qwvIRHXz/VlVHoiBowLqDEH65sPVLkuU+7J1W+nyW3bqDlDPtHaS/tH
w4zx5RE/If1AZFFcKeXlLIhTsldhWAZCjcTHIruCdT8oZ1Au9iqwzEv2FFSK9qCy8F7izYU7bYxg
lC18mfL8A1pZxZPeQa9JXMITLFOE1Yg9OzwHyoH7Ih0sZIciM487BdMyh7ek78BE58kKd9StCf47
X0tz7FrNqR7El7mOQ7i+NTUIwcH+aTiy4pSP/mkk1NWSROxtkBLp61AnNVJDen278HWEGtEFqvPq
/0NraTUKuUXvEKQHhcvJC+SIXjdpk2wrtuhZWmOTR00LPNbhEPlc9YQybMlg3Gm/lvb+BFIe1s8e
nhfLFK1M6HmOOSt4Iq+roN88Fx2NG9x9Zwc+7Ey9qwxof1k/HvsHX5b8yWd4+Mv1LCWhFsKCZu2i
v8SSls5/W0HJGp9MKZOJzzs4btS+a8sIDkrVphPF/BAeoTQIMz+glkWtsHx8nBvdVmD8ZtDb1Bse
biegKMEEVuMfiiBQihxNwWY/ofUNSRJF3/AfoDTZPp+3VincRSrQ4LD5Uqvn+42noJiOsSqQtsED
sfeBTMeNuBEp489HfByAK7dN8bT9caQu9yX1eKdmWOZA4uwjIgHmORdKuNXThYMurgJmIT+UnLZ+
cnrcmWL7oyiasIh0V/5LyAiK8N+tiT6OTDkKUnWN0J/KEmQSR3RJYAI7ufJbx68nfofPlywNKoNM
C6p/rPhfsF7pfNRDB59IjpG6BXLB/2CeO/UKojhgEtqyFjptJyLsvbbJcs4tfFd2D7S4pSP1sYTY
Nzm0zfLx7q9B2OU8mF4rs9Jj9oXt9dfyRDh+7fV0MIzzVJT3mhcnrHtFXWfi+NJNd7D7tA1JjQWl
4nKqJvItg9Y4Hh1Jbw6JKURL4m8kY0JwU1AVcVISkT5RrkFNNIM8qywidSRVF91r+qIsPCquMlc2
o0UrHl3v17gnClQTAqF6AcTOMSNLmLqGFwra/1G8aDyODIkncRHDu5zXcPTHIHVsXhMIsniQBCJK
opiMn0834fie5p3NDYqqHHGy350VnelzONf/GCGNRDG8VYobJDnHqDJJgF9I17WtuHIEhP2Qk74y
bnIfmEgqBz7pV4Ym4tcXtUejwJKEtflClsYICdWL9I5CQTT3uG0g4xSa8H8AyznXEnRx/rMZRSw9
k3Drl5bhMt5CQ5CGTuBFZ6EkRK4rjJnPlnRisjCq+4qgDD2lH/qRVqPkvAPlzjjKrVkthYOAK2Ce
4EICnisxHhCkA8zwLEnUbpxmfbdQrGghQ09dO+gOV9DzxlweEEUvxZTJpYFmuolSpkORExph0Uxv
gOug5+CueHlT/utKbI7oFWwYO7fwFyfFVmCgxNC5rTA3C+zZJBQ03wHvxfVUT49vi/ONTyNESMcw
9HdKLUcXP4LT4ZmQmZmKxgYYf/KgyZb1tqfgF8jBWNO0nPmEaBAzFzJzkE8TSF44MGyG5mlHnQq/
7cWirMYoM6+oupSJQa/OGz9S55yJz5mu8ePFZWbLIGg+u0TheP4f49y2/JXLvktTzdyVmgEXqn+2
mrI1YbatPqfeAsdGVZ7gF4YfJo15JQX0t94JXHginEYP7C0yZJTs5WPk6NIfV8B7et4VHpPNKTEx
8YIPfPRi5QL5QgBW3jftO2RhmT/Fh7DkJZg5slsvduh41kfmgogoCMudJ3VARB757RMqNGvkkjXW
l/mGS4ZWDnQIxmuZrJSPUI5o6GaVEX1ATLBGu9bYdLJso0V/94HM7Er3pd0TzLpsU1NolS1Snhyu
UV13WG4kZ6j+xubAz85D01wbihsDmD8plLAqx0la21EjKKWtl5Uz0dtFXitipe8lXlyBYUGKiQaY
UvBroI/9d9UsNO9EMaMC7Xst0b+RBhbVf8X0+Z1SCMI5yZmfe7C8+UFua9zug6taSpzW7W0vk/40
+Kfa2EKK7luvawf8wSK6hxSxH6eXqECy0yUqrh90ejnlfXEHmULDh+sYyN8ccDmwlN4VkpUoGz74
tH1w5LmHaFz3j288SLon29pcO4yOOSciYE189XTOX0tdphi8r7hcfC5zwsX1EALaXLW8U4PSkw4p
FbrdIwJKmRkSnh4mR3mhe1hSJKDA1NwF8oJMJKR+gO72QrmpSRCwkEUOdhmAVsMAL2+eylitamMW
ruINVRFMrKGDU5nW+rnfMbWnxRCL4ogGwY7sc7iEiaQgWmPmSy79OmtagOebyt3qsRp59FZ0Ddl5
QquNggbYiuIUJ1zasJMtJylTrd5F7Oja9fe9gzhOcOebjO2lNu9Y0Yky4SXsvelY88s0H3IBPt73
nZ/ZUU0CyaanC8NK08kApbcewLKt+VrxyVq95IwMsPfy85NvTrqOomyimGJd9uwOa9f+07XwqA1A
xtzd7bN9O8+IB0uETnMgxeuDR2S/C9sRwl4h+eYbb4jiWVxmnJU+WPmnl5QjT7GoNqR5BdUgao2E
qF1+IlkI+xdNl1C0ZPLT68VmttbpQ89ZN/e+I7aaMGrl0J6KL/3IFm63on0Bhq441sN7PhVwIJXg
Q7r39Aqn7OMyuIGZwh8stBVGXIxqg14OtjAVXClyaFlQFaK2tHWcCdkNgKDM7iXvfCGXy7cnKYt6
6mSRdEJxFTBFBZXo8G/+wJglyN4EgqMyfU9759SkwNzhjPtBW/K+zp4i5SFCHE1NM4tKKLlW1WXQ
zsOtUdfqwO83/xOFNrzOzl8uoKOS3hHQlwF2CKoXlOrtOebwTSy+CBLuRwQ+avYs85u69xXMlAKU
DVF1HoWeeOAI55Fqw98L7etSY2cMVLx8Hl5Xm1IxcHQtJXPTQgCm5iDZnZdme8uq7XRh9PZ+vdYz
5+iJpxjf4cI5BGLY3JLw9XUoxPX1dqhwELUFbvPuAu8OukR01ruxXe6RdgjljgAb389V0IO31pip
lVIwpkXossdGACtR3fmLiTJT7pkMf0L94k0VGhn/i4qMhxjBjXkrh4zm1+S6s91piHuSVEv/v7SD
FrOjEkodezhQM+DOtcgee6IZK6/4xWz+QD1FT2J/YooHrXXB+LKAyxKHkwqLpI5AAnsUDezvaKWD
sW9f+hU/FaAW4cJv5fHFzRYWAKmxC9Kbcx4h8ZEJ89V+yKrpqv6EvusSbPjt11g8e+NW9Vwcxcks
ZB4LjyfDiLOUE8Bom3XBdA0UouMrpiT18bq4p3PZeHdHBuvk2lYyTHeyIs09MdPluL08Q542hf6A
K+gdImDLzr/O0oLiyuR6tDwaxRutDERGFvIx+z02mnOQtnpNeSYBmkhhW0WqD8Ecw0VoXJGqcvuN
9bxsUqUrvG12/0dcD5vrXJw4DQ2a82awnMeNMl2EWar/TCB1pNQTI3HjFBXITuCbh1+tD0Z14rA7
AAgTFgbdOw7/V3bpmZCrFR4VusFyQT9gQYi4YO+3fdDO+9rWQne75xyhy/QrzxpCoRPZt0pE9Y0q
p3dNoKhA8WiLFKDaXiw3z1jC33qOdiAmtXeCB863iMqr4mgDPooJ6jGeYHuemf613PR86gkrxteU
ss9UUwCRmcLmb+HchQx8Eqh6RUF7uvTXRAlsZWtK5nD5VE4Kz3Llg2cZ16VTtOIJksa6eCZ33dyx
IzvpA9c/sYH0b5NTOcNcbpCHjmpmPQ2+GXWDP0ahkucjmCaVhModdspt8DZ9jHAM9TP+eLt79CN5
lbSpxPK1p6ycofv7ZYE4Ldc8WFeplPJitTavZYMKGzxRSMUcsPTpD2JA6f5C4jaliKkhMSJzwpDq
XKinUdwVx+xxkahcMIS/SOm4zPMPeoaLgA1EQFoGv8/eNrCWsf8Xgt7A88smJsMhtzofkCQIoQrM
3NlGaepKjvzvkoNMMZl+epcmuZVUR8cASQvdhbiExWCkJW/G8FMGcHxMXuL4LKKXubQd7yzvFiVu
SfXmXQNjGvRagnKONy437OPLtPCh/Ku/67dRkBOpiTXciIMgEa5Dae/fNgJyUTLKscGyvLUvsW+s
II8FcRrZVl3Eb10we4E7B35l0eiVr+ppA611zh01A2zfy88LVdubXPBe0YeqFQjX5F3WkfHhBkSS
BM+9vT2upPL7cECphkLt+KXEVcYzY9znvbPnve0CiHXitYxch2yTyqHd967+unqNyu8ijyYuQdqx
56Ntirg4dpU3wUi/un+aGDuMECESwVdHMtEEQimi7MX2cFKKEsG/ILBhKHrzQMwlrTOFAlvmXK2X
u/9qKqVXTBZQR+VgkDwi0E4pv2aJNePe3Rc/RXTssqnueqXZ1LeeybK6yHmE9YaFMqZmmh7EKkwF
0pFiFzosKAPvFAG//Cf1edY7nNEOpoXtfU7an2bzD70Xtp6nyZuQTs2NBtpUzk/EcTvqYx79mrHo
Do5UHlxM8gLj8PCAHozXTwN3WsE0dJG57tC60YBkVofIEA4eN3zhGE7pkXqnpDr+8XxAw4Hy+pvo
oFTUp5+4amJhayAh871l0qp7J4gIa3zitmr3tawAlsWIytRsDNw5akYtWbWIqZOpFkDMh6ISifAc
R9ASZq/cG8di3a2t0kfnSt9ePyHoLPQe+ICEx1umnFKi3i8DubqjImClCIrPRsueMsspHuvJkJyZ
Q74qnDHtc8+2c17LChmApq437SD2df1PEq393kFSWwVs8Odojxzqw7dgMhRKwmyH8CEQg1gn7OMQ
E8W+P2jAEM16vwxlrjbW3RC+UA9u/iRiOI4dZ6vEqDB9/dRFCWqauVijey/dRbZCh8bM/e5kPx6m
UeF6l3CCZ6eabQ8ExccqpF5daIwtIO306JxrfbNE0J75xwyb7ubGQDcBJlKYnBjTgDrTnw7/YSFz
EOPAa3VObO1qXxpuoY26NscJWp2HvKPHClGd8JUiwaplNG032/f6zDR6TpGmnkCgVxgl2oCarse7
a8WoAZDjISn1lvL9tdmEjX0a/5CuMzu570h0Gp3iIslM8wFZ3I2BA8wc+IWs6Bk8vcTa7Dzk6RaP
MAi4GnBG8SsMDfz8rAcCvAaDuMYqqfx6RqsriE/bQE53MqeihxH5jGMv+tyE53m5TgoU5hBZvs8C
RyA4KAknCHzkap6ynCxuUs7Jddc6ndfbmCx5GIwhZGe+uXgxpgZ4JWhNcCM+X+4Bczt2DRU6PbOm
RE195wV21RtlG30xik0BxmajRXe1d0YXLuOqMQFxI/80+DbBnikVJ0OmGtUVqfhnvB4LokaYaWiq
FMHHmbniIt3IPdQFCrD5pQsezBedzmTuMcEux+wKSLRli3XhPq28cnsesA7UzkeRnNqDfgzI88rg
et/OSsqk/DbTtZowxiGk+uNyAMQSay644eiNhjkLbMMU0ybBM7U0qfvMpd2O6jtpYQZGsEPHa0Hy
vYm6BMAG9sIqVX2Blp8fXr74Je6PlOIAC8QeVEv8Rmo68cq8Dch58272d+aJSaHY2kmtGuWdDU27
F3HyAoI9bJvkI7b9hKZU5zGfye1IaO/agxeVknSpxYv8EBFqo32kHUJAh3D4iENg28sRLWYz6hRd
k5YbKRcx0zlwtMZghdtwz5s1z8iKHTiwCDdbGyiXd9/2PfUoKt8NFy1OJ8EeIH1xRoUmmMCii3fx
C0O0GUkKv2nLjCIxsD4Ch1L8egWexQNLWJGhB4NiOUYiUS5yQV1tvXV7BStNb/4D04NJ2kiSCzro
P60cfMlVqoqUA8JM/rWt3zhw1rQy89qGisScGAnBCDxcBTVnRkE0Ug8R3vK+pERQXeDnbzbWfckW
Lwji5NhbeYD+C7hoBolk24Rq1ADV310blzhyvCEEoFfR+PDaYySL68j7xmvpSUX+2nlWLi2HQcoI
Mte97ndm5RPa/7BkUPUG41NOChAg3CloDff+ujB6/6pIQa+4BAO69fokg8uDCqcJ22T/Mqw4IXuD
cefb8PCOS/m32qNFKwkC9nY90wABVyBmooSnxck6hZNA330liL2oAI8I0ntr5C9aVgy8wMhnybyL
coILqxQSHUjAC3WF29XWCEQp3f7TaM0N8xAlLmGvFewYNSr5enQgS6HMCV3d4zEAXCeIL3Gwdx5A
8cry7tW90SFlhM/GWINCFbDrw31v0e3UAZMCkSQaMFS6EoRpw7fyYXgHcGAhQscctWhEOuzOmNgL
JbDcqcQ/K7zBiRkkCTA1vCzvRCsYYfVccPP8vvLdtL+M8GF4DNAM9nIltcC8F5mz0ReQS3TwrT+t
KDm+qWm4RHweKhUhJzp9MfRTlJ3Zh6vHh3zrLievqGStueVz6zqw0K8hHCQmqCZXFkes152TVyLu
JmKCvbpVoliJrS4kZAhRlwuOGqaiCeyRrE2DF02fFSCtm5RIXTmUOqOCNeNdLoJW6osxVwPN2xCx
Hx04R7ydQ6XmKuxO6nPBZ0K/+P95nwk4OMzpdLsQuIFnXMFIXqymaXQelGjUBOQZmWoKfDmgHkqG
ZBzzsKH6Pr2zuoXZnSL5XK2mGWw4ySc7YHgP2FKC4W4zlgc/C5Rbq+7bKBUeLA8/m3CAwzwuqnRI
4FjRJQ9hnLar75Qjmt2DwkbPPa1kN2WyN9W06d0PYIB3UD1Gg1i22knAoh2InAsHA59/qE9jV1h2
9SGoC1h87l0ItBvCeApXosJmUoDevp62N/0ndE6quQJjcZ7rKM2xovq20zTb1v5NoHuCSOqEhviQ
10sdXOUzoUlHu6MfjFeu+wQi5B7ZYMfQha18KjDSYzkNzu0/2hNy9J90Wmj7v7p03hfLxrjcUV0+
ZDC8gSV/1Y6lK1WZ7hsCeN4cqAmbOUHozdJObALBb9DT5oYxuww3+pG75gLp4k0XsHXkbAdd3CIG
euY+K5RSQAy3uJJhowslfWQNqzo1jmlCEycC+FYmJiR6F+CqiljdswUu8kkzJ14LFUeNPPIJRgMt
vwMLSu/REs45WFmxZy3nW+a/b5j813mnHJ6h40II4fKnxYCTkDZw57XdJf49kbmSfuVtnuRRT1oM
oszcfjsl0nKeV9vlVlddyQowOqCedrUCWBPnUag8r0gUdYBZrSp93VmH0aW+djd19Nng2nZ6KK1S
J222TGP/HEbv/TeY1mqSQBGAk2WgTH3ve5LABiszU0U9X90BByWFUe5ytOC5O1kkWO+SfrALORvo
EDcYCnwr1F8V/EOhgVKsz6Teeea2lGAa92ky/ZjWO0j72XWNwE1gpjvfu/BfZTkzlsIrX5Llbfwk
W4Jg/i45SK6NYVAZr7BBBIjutnYFZgyxL/gCAx9yFgi8dI1Z6G1eqhgdrKWSJf6isUSWzr6MoOJc
Wz9iAXGitIfr6aJ+h/gjmJ8d1q4K6IypTHqwm25PWCH1T5WkYDNm4kxQF+YBBEc7uWnR6MytCUP2
+dXaBHdRsWgQXI/P22rAO6WI9wpEiCYjrMktO98f6Eh9TIBKN2zihkcRlFngwmLtH2N01rdGxGTt
f5xgm6lfD0cWSREzcKuZW/TjZEFc+Lap+bi/q5/lhaCQM561+VstkhR+vxZMz5+4bu3wpQHX1/fF
ezAoJ761a7BL7ms1tRdJrMHA+1UkJMBIQ0uuWKTFeyFs++QEXv5C7AzC1tipvyOrvghQrFiK9t4g
BIaGSEUw9NiGVTYKg17vL0Ea94UW9YVZNvEGiIbJyYCNxpxb7elLn/2yNy4QLBMzr01xvGNqgYid
nguj8r+GD6g9uXbKjPM2DgopRVdn39CShGdwgZWl7mS39uSMOrKaB68Gzo/IJTJWMG6jf2kIRlja
yGcZa6CNatf/RmF6C6pbQW9nBcFX50jYbaX2LQWPQsa87QKWT8Ppc+Ghm+eUggc2X/1hI96ZH7s4
swcb+1ZaZVytAcp3B6qYg4I0v1SpWQN/tN4h5d7r3nHJdlhmxHs7H7s9Ascw5Ug6DM6yGSn3k/Ka
18i1fO6D92ReXW9o0Azw5fssvh2dAdArxxqPpHbyhUzd8YUS8xPOgn+eWdok+A6UrhG4UC+2R7Qr
LxE1dbChSyrB4IwtkKruG57/TH+pfx2T3IrTAhtCUW+m0guvN1yl6kCRRNLbJ3L5eDhzZx7M8q94
oSFSAi99JzRUdzejAA5Cl56QXN8h6k/MLtytehWUiyjIBDj2lbckbFgleeoSaCm5WmhRVIq1ltL1
hfSEo2m6Rrs3WnOoF7z2dw4KvkI47yrMnHYU1MsIbtmUUTcKa/dPAKecE4fB8cVLd8w1+FG2n/l7
NXJid7uBgYf5ckb0Lhv/NNpSeJcau7QTBpUhHFDBaTQa/IaIToHn4RBiJUZI09aBE3loSqBHupYT
+2TPTAr90rhavt/R8YbaaHkTiyVfgN9jgGwDU5KTnKf7+8XTeZ8yDHPVwjFv2HsGrS4JKcOcqbeX
t20u5AGtNiGzh9B4lZffthi08qZZ3uHplhQd+VEFqnXyjXp7jSstn81uy8GRhiNf9aCjZEv2qiFL
K396t8IS8L6YGckhhzOp0bhcqvm3oJOjscFXxQXQe9s5+oqtOI4oyrGsXfddQD7fyDmruGOToROe
nMVWk5wsMRI2oAYt4ye6gw7/0xiPxAvD+kbDjxFfg/V5Ok+WmhtdPN5QgRr9pXh+4LaP4EztnmeC
50yaVzKgIYwoRCniD5uuaeCqP3ZP/lYNlpo9ulQ7p5LuZW6g3kttgcRQ/N7AMhA4oXwtgHltnXMX
mSRw8HFBdq2Dr/W9O+JHBoKdhBDxtf2ipwBLfNXIFag5O8thD005ipEC5Rjqgm1hp3zKOHzQajsz
CYWBTF7CZ0SUFbmrsnIAR2cb/wcrNoJvLyprB6mzjLLrtUQdUHRr5LvPqGV3U9lhj6G5xo/DeCES
UfNVfQa3baahAaX4NhTxdWGRcWGiJbQFrQOd2lHoxBEim1c5miFBu+Od9PLIixYg9whJ9xJwl38z
q/1v7klTEqoPeH6vP3QPkG/CRjw/J2BC7KaVwai6gkAizj9B1ceAgz62t7/KdSwLVJXmNn4JQsib
+kSH9XB3/jKd8LvB0soooGlzqMTYXDyAeGiIYI33v+Pc/EMZZb9jEVlctvDexHqjGW4+cDs4Xlfv
fPZt3LtBk8v5nLAu9hEOrmlK7NRbPLoB9CdszJryOm8C+4PMQuuSL5MQ9vva/muCEyUaRImSbLbv
nhxYj4Dfp8cE4YR/sTKdmCXwYm8lJAdKqz48B9ll5jMDYD9HM8T8WpBwngp9GSwIrjiBz7ahJpAz
6i0cv4WtGXnMlcv+mPDWPDwFj7V9dDfaoMfGqvCk3eJPBCAce+MNTEq+3gMbqX0oi8gwWrIFssvf
JozPa7ynGWTRmNKJfounJHfSORPMFZZT//G+BHdMORzNQu+COQtYhCaWAEBaFB1GJqMRASPK00FL
Zw4rXQYLwNsMNRgETipFZrPepf1RjwCBVY7UXCLcbI8UY2jfVM2lyvv0w87mqWoE/OK16hFDnqv1
Vq2ti0lExqdIyb3KmdnnGIRtjO6yjl0si1Cpp5azdYKU09fi0mvfnlll5nWNmY9Fs7p3dOZmvb6x
aMTxB7lyrH3QqsYGq7RQvhn1HdRQi8RiaOJPH+usJq5RR9lFjOZr/GO+2CPYWtYWezZft8eL1Kqn
ELf4qfLPAK5AbQ5XYSdoXB7R4R8CFVDUWaxlOi1rVWHwlecFwx54hTmyzKS3ykrvAx66AQ/CyiVp
OPYKdxFZXZ16LJmvI7cBF1+MlPWEuC15OllW2JIfJYxrgY9PCpG2H0/wib0DUoC5nlAOI8yuW5Ra
FmTfbAmCtTCX4wZnyEXgg0Mg5s3jIClsY4q8++fHUiMb3snY+ZTN4EJVOwBKZ/E8I1qkpPaNN0Aj
53AelaaPY4/I5dACdPrzKOCyQLD+9U5VMHyW74jb04HwIbEZnT8UN3pNEYMnWHEG0xEfp0jd5+Ae
qxKeuIy/miRbnbEKqoBaJcbwWoWVRO8uFSRGvdTIjryl3DR611hzgyCeuo2rsD6U6OHWvkCGPkms
2dstr6Kp2gi39Lr9v4lwtc+Jir8rjFEGqSyEQTk9ba0eq7iUZccab34AWbZn5yZRnLy/2AaPvwae
PrNILSzZ469DRC7dPfbpttiYl3vpXTQq0ZnXFT+AnrWLMcrPXodsAoIy6rp69yYGgDeHgw67NO/Z
r3Ci682HH5lG7frabu7+Opxrrso=
`protect end_protected

