

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ej7EX7T6jodI3eeD0H7xP7NEyUg1taLKF1qpZ7e57tL0iU6rkTK0vgAE0UOu/qCCPgUCRFleMSr8
MejlkfKVxA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jjV2dzJX3n4L3HsNul5cDmWrVN+3MNoQlg111ncXDiug6c+Hp0AYDW96KLd1U6sLRz7QUnbnueaE
xF+B2vnLgBdPLCCDDfcWlmaB/J5jr+esdewqp4HS/vy37HsLlnK/FEFLOzJnAXzWtQyhAT/4QGLK
J30Zap//VWyOMWyxDzg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FWF3yHEVcnqhAkSUHTIcK8E/sEDnrqETjeI22zIZ2991OQLC87InFw6ExM8zuDjmHMeaDVhZNgEk
FOiHQQgqAiaDBSRrKIAnmeTWOUZg9GXbgGqP5gdtNc0HO1kk6Yip1QGxfbhRFwh3YpTsYnl42SZe
lwn+xr5JPt/+LzO3Ucy76PxPK+my9XGZy1z3eQNpZ5DPXLmZrEePKNE6iSZ2gdM6mps3ex840jBP
9HKbLlTih2X0RYcovpKU5Ee2H4f4JH0qesE24/5PPimwxsoEUCELdv4WhV6rnOo0NummHoq2Qiwb
ABs3V96fj+4Naip9DM3txQ0UuI/Fn6jM5HkG0A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tmwC4GWVR8MCeIowm/YZbGdijHlwWOF+IWQekrx3XWsOmCPuGxH2I5rGh/X2IzvoT41kcgt4ZlEp
hafGLnA0b8klMWRXXsc5z7v9ErTJr/tuDh1yutzKl/g/+7IIKtR9a/XXPxsb/HsXJTieMVqfGEk1
+D9EIqvLpdQvN6aNsvs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kViVCZwuwF5OvDBJOmZQL62U/uf5UrxeY+HEiUFWYn716G+pozUBiJYEnGflxxZLb2rwSpoW+kJu
v1O+hPcgXm7xcrQVH0H6WzIP+gkZcM+HALA+PMYyNmmYtuHaOILNZeCTvfu3PAFDi8HYx4PJWJWQ
OFmtcTxihVQQD+JdT+Pil++JGRoxGJJNnwClvJdJXf41fyHvCBC0BBG68nz+8s6lfzy0gNhNaM/R
3c+a1setSuKSAuqXS/QeCSWdaP43TIODiOXEbfcQam4akexjU3juk3GoTJK+24GmmAIbiwEo2RVo
YLpaRpIUYqkEUAusAtWFZlO3GITlrPo0lSa9BA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21632)
`protect data_block
wwkodWTK1cO9AV2AXlYpdYKtSKXHOl5np0qTboJyb/rQQNtI8w91OGnzHUw27XKrnj9I/VdGPTH9
mkXQyxCyO+3RJGNrD+3VwWyK0VNl0x/UrgB1IuGJrcNRsyMiHKOXy6GwhKxYnpR+ZNaL2P7cvad/
bQD8OBQ6HBNbGNeinEoJRx1I4a+Mn8bjaX3C5OKQc1zCPPBKIbkwU/JYRnwTbDRcoITBCVyuJETJ
Dddb7giqjcq9T/W1kAc+ijRKcVBk81gX8bv5hUhzRKozU8pDyabDRkzqr6tM9/YZLO4mS7SjhYio
AgUEBS+C1vglTTn1V3s/tFjfSKdLBGHHzDp4s79C/1UMpks1GKWvptL+XD32gmjcqLKEhX4dwzip
CqC/VSRMDZ9cGqXXBoXG+DwfqAj5A48TcyaIbtUApo5KkLxgtVMwLp8xPbvxuNvapBadNZ0e4XDp
uy1xyPW4ydVyDCYReztG4bDm4fqYmoPHTyK6Lq6mKPFc4IMsYz+mAghlLFeNdVQGIyGvAOQmqWv7
USzSpoAdL7yTZwBHE0DM8pjWpMmms+9TpDH3ei7d5gHR1Uhtc2DMgOj+ftxLjcfYq7NSCI0wnGGq
cYO2rHMzbXEdddJCX+3lDpT2nBwCfbXerj7DDMHpM/3gxpVaCnQ9JqgKWz3bF9PS75TKHXJDbvPB
IfyduW+awomW6iZhQf4ejRiz3hfmPlrjxlzZN2yH2j2dRLTwX0mFvYAlw23b7wZ3xVDmtRLgKt/W
Cy4shHpzhMSLBt6HddQjJuGTWA4cfMBVQAF1veClvf8oRGTIakosW1aWZ8tj3vWI+opI+as76Shk
9jLkmnXaxT4qmJ8ptqP8qf7V1QQps3RI4SmJzgPFRvFehHlRz1OVfx2FODl7bYU/7XxKLOg3RxXo
q3rcvivaXu/fGoJlX0SGQBjMgQNZqw+669Q3kiDAfBARKKbpiAi+cUi4GU+Choec69sG60RA90Bl
ILlLeCBnFxiXT+FWZuQrLRRvvzPS5oGBbpQW0W1UiU9JrF/xNpKsbL/PDZIuuT2Dm7BQXrVia87B
4v9fFUeg+d+8sgXQFnDO1A4Qzn5BJEaLWfOfcS26Dl7FRrk5+pT1p3cPyMCc4nkPrhsmsf6OMhTu
Yxi7mLoAHCMpOi8c6iYj5qM1Agu03mQ4BzG65DEyJdsaDP2bZiq+TEuyR5hTezLidFW8lVqMn0gf
urnzd16idEQMNn7HnEIRCTlcEQsOqwy3idfBODlkITfIitzZDUxXTO+Z0BNA/rbmCiLHwrn2kFZp
Ho4nkoZn4AyHIjM2Fh1Il2lPrTDNjj7YOSyvaciYRR4PqOSqcYWVS2Vh+JXxinE1ZrXv2p7NeSl/
0fCBG2mLj+5nBUYOoEZXFZ1hWxnc7uQGrGurlV10nzCiXduhtVmDQI6v3h7gs3XSzpJPllpDm+VS
0GZjW2I8r1+ALMrtmHJlNn+BeHZOHh0XMc5zSWKCPy5NCHRT3hIcj3SKTwoF9jw82EMW5vTsgDlm
BIXzUO9MaB2LQKUjUTq9OfIIjPcPVhzD/xqDqd2F3K7Cdww3I1zUonbCtMAnwDJ60k2Vkg3EtUNo
fyhj8UPCsUJRhN1W0cplrdMOjuKXCDRFBihaaWYJ0EIFgnMcC/eYm4508iMZtrJkW3SmxMHt8OKY
Au0vPNE+kpAYgph3JEjrWfQ/g0dffQNpwna5tbY1KLvjdOi6M5KDPpb3ZTCZMZ1KKn2RQwsMT8IT
r7wJzjehKnvMILmhfH8eG8AkhCIER9Sqa5D4OS9pU8C0zIZZ833VI8xmq1mnuzsWBzu8111zyEvf
Mv/oAjh+a/oVXV5fiiZTBHrKytJiPfj6gV9YKAMjb+PTlBvVYg0ZO06JyiLMr/eRjWoyHFzoFDmD
9Vb03Vl4s+fAW1IYFjP1i8BmfPytaGtd6BjQa6WaZXChDMzFHMG8/1HqVGN30VbFUlxcny8g5BOA
AEjYxrC6EgD84fzXuIyhmfUsObQNd4mmBCERkZOP/0due+mPYVpwyrVm73KPou56F07QOBlMdKkU
D2vlyK8rxrZZHbU8QDSa0wr+zz/e3eQj2zS+tM8EnYaoeIJiermR6A6vwliatFc6h6q0OY2rGJ37
uQRbeTjGGY9T1fMAxiSeaLnnc5Vr2SMDHoutGjKVLx76OJYY6xP+WXRjB0IBSZVuDg1pPByHaqGH
rcXmdbpTZioyj0H/9BjL28cU3z+3I9QY03TA1Gy8KOpXVWK/Lus4TZa08yXYG6IBxgPDWL7jVMcv
pqMQIgFYfMYFpRua1eydYgHXkG0kmIedIWk1A2296QmXSGNV9AEgIfqSFamfhk9WvwDyD6pvXlrq
2ptoN0Zix6sK378tyjCz83LlyA2/gkB3FMBE2ihFOf8GRG0Ia/T9CX2QN5dl99jZ8h9gLY2lUn/5
8Vr3nfXUl9dMXbq3V73yjmBNK98ZGOCH3XtfCsE++JPBUYnZVRWB1nHrvl3E0r6fRCY1ZD8lOJ6+
8QXeVQH9sHHvBi1smmMNeufSnxAAhShFOPvVjFzcrJ1el7v/OTAguSmN0qtmS3vsgwaTg3NJ5RYi
+Ymw62WbvGl4o5JJv9N0y/UJSIHdHK9lhSinTvoMp+Rrg3hDrp+9R+TYDWJf+ACx+ZwvFgO6Vc7I
BFbWgY7yadDPDcWBAYJGzwB5V9URVjxkX5IiEpFwiU88UloCNG9HtUDRmcvsztq8yeb3XWBO9odM
50LTnelfl46H8CvNgQLCM51TwHdmLfPc2AmDYIpf/xDbo7E8BHRN+nhXAFr5Mt2OVWGmvPOWLHSV
xNPwdbVxo4ETv3DFVyuRfCtmRpQKhGKm1qeOjHpJfgx+d4Tar3FWcUPdiGn+wvrO/xiZs11GF8Za
WTLsc5Yy4a044cSaNZfI04KqOATdVkMqdxISw6Yqh0MZ5xQyyXL99LeM4xSX32fR/xCf3e/n+KgZ
x6kW+qCxltRXcfuiyKpUXu1b4BFpV+FXuDd6NubJndX2Ds7rUOjGokkfNOOcbQu1r4dESmklQlHb
0bCSf9CmHuVeXtC4HRFdG4BKGXs1+ZufWZpmH1OQogIzRt/GL8mtZFZiM/nH6eGDKgzJjWA/eRzJ
RSzsh/aCuprtv9YMP67VjmObg/CC8rTGqxCCNAw+kRvEW5pgLPDqBrR/Lx0FFLtG9f6/M3wNrdWO
um8HwjUjhAiC11bhSrsyngRXRJ/CwCih5APYm59wKLvB8nSvSNB/xmnUfONTc58WLjhoPOnHiqpQ
6J2Oo4RjxxbCsKMQry4Na6CwmW1jwn4/8Y0W/dkQPY+LoofzTCZhzwxsdDjur1B/GT2zOFWsXfeN
43YEZadd4DzXUul/ScsU+KpDy5eUZzsf+smeDlGma1FZSRFqnRtFR17ciWVb3XP2n1rfnNNFS3ZI
PclYVk6MgPhGtcZ+M9sWd1yWYR1r+E6EwJCx3KwG1J/QfyDFXBoNIY0acyXjgVq4uexJcXRRQEND
ySlr8Q68WV5MWbvNU8lBB5jHfn+RboHTEKSWhza2c1jnjYNyCCEUX7JFhc9L0silqvcbQjiHdC9s
4IdgwtSrH/Yph4ibj/d3Q8YoM916/C33ytJ/db8ZgtKUR7O1O7o+U2R085if+AQlHUVhaDxiMmVa
JBl0NcLweKMVER5HArhmdRmR4beeUGPgq4GAMiM3Lzsx7DTs6unQuGOGeehdbtjGcnD1mLYiHYQ3
QFs4ZCnHPd+yAQkAnXgaAFpfLPfQF1cckVgzcVTXZSqe0W0SiUU9poOXNdb9+thUoUFnMUgmWCUd
TKZm8K30rLqvBPp9ue9U4t9xPbNnPMP2Zq4nsCpoy5Pu+FHxgydNm3VT6cuaX85SZ1jS8aym8KuB
xe4leRPC9i4509UW8nSDpKhYyldM5UCG6kmJ2tVtVMofBBUy8Mz+id4uPclN1Ozqur7YNr+Q6cvt
V4+MLWmAE0+kMDo92x4wYJB3IKTgU7L8f9KwHb8TxYgXuvD75N9Aon3ZA32KDGGhYEEGPsXtw4a4
rTb3D9O9bEVk1Skj4VH4rs1EK2oQj1uIZJ4ydXcOFSUbqSvHuHtiOCaUvr8vMJH1e+nePJOgT5w8
IugP8e3J6HQ6iJoEigJlRilgPmaXMjWIMbCM5ysF6XSKAXYs+0MTFycTrQBtvs+IPQE8VUm/Dyc5
JG5fPxkZgNEGj6dw+b/rvwPWuoTUr5dbLIh9GAG/+Vc60Bxq2LfPYCbiAtmae7/GCcLtDgqBmbBU
DGBeFidi5DlHl6707PW8pxzK8tSGZ7cE9+H+lZFvuUIlD5lMPlkEVfk7qBucmwIswEMidZCXLmZ1
nLfo744a79hdL3L+a0nEEnBBHbslqyjQWEG2pp9CeNDjT/qkE7pySqrKimsMDvMVcWOOpinR5hQ0
fBxj01PpFylPZVfHQ/AGGSxD7xjqyWzsmxfjXMTDlqU9qqg453/AppCGatbrSpEmC3NnJTAj8ZPD
Ras8oXqSMzdFbCu7OXFAXZ3A3OwiLnoPTfXysm5Zoous85TJ6RTI7vWiM0wRz/5QpFg3x0WCwQJ5
byqvH1W3OscqymrRM336H5CQGjwl+ZfI/8pGmEkttfhkXw2VNz+By/fwdhYvjBQH1EJKm3h7XEPI
hdqNvtL0n7rDsW9ca5k/y/creB2M1yemIsLtuQ0FExqFx/ovCEaQnfBAEr0BKAo5Wxp9cTQBs0BV
BCxMQDK93YjDuxhSN7FRqTX84mftnlj1TyOvUEHjovVQ3Qtv9qwzYK3KdUmMYXl7cJExcdCdauRW
K6K+89fHFT8zhvAW+mrPNyD7hVWTTNa+PElFMM/O5rTRCJgl/VJC683AKWlb0XbGyot2pqz/pf0N
b67WMQKTJ+oSzgqNAYN3faz0D//K8PMHeIiP7NelkFi4AdrwOLi3qVey5gkhTcSYmqorQU16X6qt
NkgIhM4rXcm0bn61f/OIjLFZmyBobb8w7heyRNF32B2tvjLXnqOtxtLskSCuK9p6/w2mrXqP5iVK
TK4gVacfXVIV1l9h56QDVmu8DB1FoyFiVnsIjwN1/unaYqGwCLR88df2GGkxqdL0NWgVPtdnHe7E
A7CBLmeSdQwTz3VoNm99YyIY7pP0HRTSGefC8FYDotO2cBA03DnY6jU9TEdSnkS/NaB2t9YnBhkj
i18qqZf+V9+jAoNZPgmBmpoBwWZH+i3WacA0aYOKuHxF/MQfvYi7w1wBC+sL/U2gpWP+uiekSasN
PEZqlXpSjiLGjKw0Q+eM/GP9BdnLukwckEMW1k2CRIPv23NAwgXphQWVHpu3NB/y8VQpKbPPlmCI
p7zlSyW2UJaglbAp0qrUwAeh6Qh587cByOddG0sLnHt+pg5qdcWaZhVTFDlRY6qCI4NXMn2XXBNc
Mb7CViKIp616CHs+xO96wI4x0NAUslqzyuZoBqPCfbUjo/oRvIr8TW2joCssSO2FilO1vCPEKguJ
BSH6d99uNuPwZ3XfzXdsUQAO5pIsc52lX640nrrqWw5FPlKpJwzCyPsqXgvRX2IBx3dpbTZcWSLW
gXy2xdNtLuV5t9ScxM6YI5ovsDi9lH7npSjpMlAHcucXWQ+4U+cxVBWPKuf6Z6l75kLtNwvZ/1Hn
OcJOifz/D8wfgvxr/Am3IwEJdUXuBoMPNu5FkVzJruuNZPDrrijaTGfTIK22LX5j7AT4XW30E38G
LaEgG+2w1MbYo5Hb/FRSZEXEsKEAhDw4lW1etOYxeaWveWiM1SHMmVjbEiRheneYFot1a6HNu8WL
vgsp5zMxAAQMZ8jEAODBjeEIft+xPQZi/gf/U1gjvGHQ2reBHw3Qi8PJlz30vprG5pQ3zqnB/S3+
WU818Fp1vFGkDsAaZOfLc0/I8OF7ZJaAhsf9363q97jpnTCDe3jzn3PIJlXmV+DSAFU2K+i4qNjo
au4h2GyPD5idTvBcjL9b2lk8RVhWLhjJwtV3Z3txfdMvTAfBDSltG5zXt+tfohjRPcLsRVvXNp7P
S59IXyuBeXvuD5M+nqKXgt/Q/7J3KGhiOTc55/X9wRLoZeZDV3mpRVOsKc6AE8V0RrHXwoNBp3nA
sdSQTf7SOLbgk3uoRgl6eOKlCm0cIYsevryE//99qzNr1e+bocruanzeT2zIWGlpCM/kZIsl4NLE
d7AmKxD+IaK1+1usHeMlDJRSrtT9MmhaHmdwomZNEhTO/auclZg5qEe0nH+D1hYEhbOt3clPGra7
ZEdt5HvDeWqe9/qYiqEbQFsUVxkYYI5chVLfrseru+h8x8+cs7bshWgN0u9UnBwfmdZ7sYI47dHr
xUSe0FWmsasJGckGeqqI7xAfDJittag3vHlqqw+zDspgmMxfNkyACrS3JX25uQF/Z2M+wbM8JWTZ
nexyYMcn5sPDuc0McOFf8CYtBG4A222M1GkOasav1vsTCTpc1byuh9RK/khYSojfryBzLdDB5qqh
QQcpUtHDWGRpyyBYaCeXSatEBUl+ZF7YH5gF8BjVpF4v08VdP81F7T6x7/iemizykS2tgckbP9Nk
wolf7TPBfQ4FkW5MZP/oFOxr7rJJavKq8BST/4xQyFz4sduexyLQJXBGtKhw2hEqBs+2cGNLGiCA
OUpnbWaERBA6nlSP0/2YYoFfg9bNLgCJ4S+YtVZSAXskdvT/R7qj9txC4Wvny77iz5qYzbVD0zMj
8Zi+H9nfLR31rVBd92VkedxeS2sDk6q1vnjAg2/JXLS8vOErARuBAxoCg0oToP16CF5Cqn2cAo9O
LFk+2KlFs7ZXG19oJDWKIkSv4xtKXSE5Xv594tV1dPN6AUiHa2nLQGlGO6qxrxgoYNRcGNT+s3rE
j7CTefMoUlTKF9DMnS9AmhQwlqiU236GijG4LquwQvLoPIOE1xahlXKqF6yUDKcv7f6oAC2qv1Fh
b1VG34rTkuwxGF5ZmkgFWeA7aW6jHhKGuzL9kdFCNyTeZlVy2UT6W/saRwwTRG1jYqVk3cjxIv8K
ORUwrCFFbBIITSYFo/c1vKB13AqKkIvOobMKJjhIj0A0JFB13v+7LH7Fpwlgq9rU6tGFVQnrlW4L
hX8NHYapnujgr9Dlhom+thqxZqf3NvxC+Luwaf87ZcLPOF/I0IJ6j3IWrlIal03w3Ye/nOMB851L
/Fn8U5kG0UAzJD4xvlQYboKKRunnEaqO8S78LIzK9xbZdINcwwLM7VykwssIX7ZNlhADs76QnmjR
4W15FORfYZEDO5Y2imZwkE3zKWP6hwP6dENDcN1HkVIXnZ7wTYFjrOrydJDaeDVfNeN0aFYz0g8r
enu/lD9RvBP2ZHca2RvgWL39CmI/mhXc86jGuSnI9SDBEeZw8kimtaTCwnUs5mtrxHGSdlioNrG8
eKRdPRGAyZcZqIO/Ym5ovbjLK9d1Aq8m7DBD8Z5zpiNcLLDtXxNJCIdp2n8OsLN08oelQ9yd+djo
dXkqY15Y/Q1M50+9y6L8mw6ZoV4Y06YL+yD8DtgWcI1Dqoq2cIVvy2o438L5+EBmn0w3RvH4gN9j
VoiosbwQQOuZOFKAQ9ZBdd/9Oj4Qk0qAUWfQ6ug3r6OmsIaois6joh3GAQrYdYsMtUCBUktpOCCI
XOypKqkca52yMsQ1TU3UjhjbxSFhYRhNGeztMm8cbOh0Nmn9qeyJPDXrYKmNfoMC7dH7yi4lPxqo
uWF+JvXOOfbL/yWBNEnXBMVA8ZogDPYE4ktW75ZoQxjYlUjSfsai81tHSYGj6g9JqZEeDHfsvcZy
7E9R0QJTsTTBlpXD+01MZ/1IE6X3SAPUK717oEiSBvxpyY5B+w2Vo++uaTKGrtwONQp3CUslJlxg
SV20VNpOSg2UCsdY6b/5cniqTcLHS85A9ErZYx5LJkS4w6LX2sOkKEBk9qW+6WBKKyqvPiAzdVTd
gbRR4P1zKk3uwBCz2qpwybjH6cn5g8tJlJrMQ+pc6S1z4EW+hujgx7ZGXf2HRk8NXiWIaGIMz+/n
+x2hxutw4CzECOX9RbdZv3bkRhU73J63yS7lz2LL1gvTg/jKnShhDfjjSlhLwkGtLh4ZmbeQe1GS
GCQI+lFg4sWUhaer6AjHYsxx0dNrmA9oWpsVlQBUScnPoHflunkvbhX5/XehMgkDRx01KEzs6Q2g
2J7N/W6RdrA6PsEal0orl2dW15hxz9uoJj3DKG2WRed/TPNFyJARBxUCvkfhJmI0iRi/QRSD7mh0
3/7IRdgFHzMucnBiGoGVPXaD0kDt0N7cTkSAZj/YXKMzLh5QoT9hmBiACzUkeUgt3hwr6ZYKR1e4
yT/Qsd7ujayZFuHWMM5oJZ5gC6oZZ13dh9uQibtLaJK1oE7lqCQ6zTrR7QHnrOpxiU/tsnYhHPVs
EKIWtj3NLtDN2D5WefDUFIMS1tIuJL6xLEciWa6IGpfyHfKMwiyhR+bFTAXwkJeLnbwbE+lbC5Zz
COGzmwSuNNLJYR4ISHi4Nr6+Y/d2vU2rPMzqjmAfCsmo+DJEheypPtKKLYESAd+lDcHzuSKhLmNX
BnlHL4Y7o+8w0JpxS3GlbM4jLqaQOdKsOmzOf5RP4JhPOYEGYypyvFnln6ie6c9g6eNKxB7FqWHJ
xTU7L4e3l254Q0YAlYmRBWqVjuhz+uxPcWvXfOizrx4FeI1DALwdbTkqPCKi9sGNYDywyF2XAVej
kN6/3UL6fijdYhuXzkhw6VeriR5ACCEhGB4HjSqzcAbXbuzeJlDX68iIhzhFESfkplMsFV8cdKe9
UHJU0+YTvygjZMO6r4K03c6VEoTSSm97lALUzlxOr/bToBLAJhJIGfXlqvUbKefCxdu/Xu60VaEj
+W8BO2XKu0aA395bxUtVotU0BYisyVs3GwdNgDBz/DIrN3oPJFRRRn6RwuV7z3f8SUfWqtwvrucg
KTYOiBAiH2PFL/aonbB368fB3lfBHFMohgNeQDl3vt08BK126qtHeCAhvDmBj6oDJChMMoDKHfuA
BY7BIcLf7usgAKTSEVa6EAV6di4M8kklk5B3g9YAJdHt4B/WQzkOotzD2ygMQjm0TwxiCFtLi/sp
pz8rd83cYB23BJfg9YGkTUrR3vQRoWkzyuissmH7jN4Lk9S83b6lmYMEFpH66F2wNMX/tx+3R2dO
G1b9GRQU5hbMiZMX9nYgPX+T0iAxR2ECWT/AcVokEj3Ha5zNKKuPiYUn+OXx2u2wBMRGNQ/AiH5x
UGqOiBHSJCSqUtvE2drw8GqzQBJuHhl+xu7o8cUpuyQPUOTjNrVAlD4tBeAAqO4iSXktLOZV5+ue
8PHcye0PW2XLiW5MfXJNwHFwWk/4XSp15vylDD0dJECd3K3tYC9MKA+3pNIxQdYkPyD76dtHBxmS
fbrhutsaIjFN4uWz/u4mOSfeoXH4fLEwW75r5g4xF5C7C6+eURS5A/gvj41eUxT3rd0Z6cMrAXdt
zyVKmPSzU6pVN4r/NXBQf6JBE6UuZEem2pifObOSe8NIDNaKTtWPOp6kSg1ogCmZcJ9nie+OADZe
044xe8MsqWcIfTWOdXMmzWdWmSeWkOkYHqb3h7KCxomVXLUq6oKsw2oJstIKJrsZ3CT8KMElLW0i
0qTcIa4MMqCzMjlEds1pltbwM+3iOaLLaUDxA1LfUb4ndT37VS0qS8aCxfeHE9KJdO/8LcxVa/Oa
T92x4HzRB7hqLNKes1cCx3pPLA1aYuDBvLdLBbfXKxE91Lgj+A1o4bYr0UByb/0E/a0yqGyvv321
XQ1p+IlUpNoqYWVjPBvL8DRxltIDaSkWBN3b5ajAbD2nRCNA0K0j1MufBHEKzdmlT45UO7OyXaQK
Sbj5QK3j9pWfofS3p4vYYDwpQspGTiOQZhT8WmXES+AgEsXJUx1X89GXjJjk1JkVtUvqi4JMV37w
1m0ZyPugHRKZxuEEzZjOnFtKeP3fvG2bu/22LLAz3t/C91TssSABZXKSlUQSrE7zR+7dUV7FocZE
1Hh25ByAF4CGU9pTxlT0nYhNRT8yHJ5v+YaFVw57XYG36KCGDMUy8KmNDyvB8dGPZmuRSQGt1NbS
2tu4tmARYnqQRIOrgg1RGuBpWMKusiP4EXwHAK9gyEXhiZJAbhmqRgNU+ixyu7cLPP3eEdmp6T9K
bb0EtdyvRtoD9Rl7P6AG5SZGsret48fcXAYPICynb/VS/8Rvd73GlFpT0g7M0WJkyjNZqt///GNJ
hGdIOlkv+QhDamWCRjbNRYRzw6BbMQWSBNFGnuTuV6kXqrbp0vPE1cAV5mfG4dXUp8kVu2ZO3o6h
csNwHvQbc2kJ5HmtVGXSRNGX59yGnh7gx6CRkJoS0Sqp0omBT+opaMZrhHjSzwErJHaK7MA30Szi
sJGa85s1p/a5Xg97Cts3NAUV/rLbPL9KApJ3Zq0UkpZN46HiDQaWFmWI6DR1aBrxfJIAnkqsI5Z0
gQ8MTSdV0hjw6XED7ITJqGl8vaw7gk0IqzmMN6XOu0kIulVf5VWBS4xrdZ1kU0u8gETdQFCLrwU9
Iue0onLKIB3z3MWS/lWi/a/CePUXDM4byxl4xg3DXamGW1DS/vq1kdNr1QOMpVvp5E2KOp6P5Yw6
aIUoDpJ0tW9x+qEIYaaasK/Pr3YOB0zricktskeRmWtwSOZpdfU6ZwGXBWlRnhs6U6xvLXEz4l3S
Ryy4ryNkytnC+pJbM35ywGAYYcgA+jvIyonJuDAKdHF7hL0ABK98Y7CTTqVRUOgA648ZGWZD2h1S
8jGgewEb2h8qAQ9HLiA4u8bDy1dT6C5xj1Vi4eQrQrfFD5Si1G/UcO7gYyXerkH6RFlDf2MkPqtJ
xQ67m5O4Cveaawz22glLNmJRNjc6VqeOETCF7of60DwJgCuUEFW3I+wcvdq4F0w2evznJ13LiHb3
wIO8Jc4RDdSOtYVL84FQSRJB3S0a3ZK+Rzix80Rao8RD3+rlyujmRBu/sVq4lSX2nrvdMMHhLJwG
rs15atFNA8wkyY8sAFq5zvT7JHSknPt03C2Xf5tR79JV7r8s8pxkrN4eW3sF/esM3l/hpxbKX9TO
Xjn7CyLjbCz7BSlOmC6B5uSA7YtAGE1aptsk/mFB4dUIJi7IT+5LNQ3tF3xuMRT2zaXEqth5HB9L
h6xmMy1OFKQSFiE5wVdtUw3XMq05B48+BVa9hdmVWp9m+9oQrQ1A+jx53TdVyddIdiFD7cTrrHAT
0ik3m/Q80CTWSKgdjpFi5xFkB2rnqen1W8Gp1nIR1C7UvQUiP1yBfw44hUV7nv1+8bmn39bat/Qy
IUui8ILlai5fh5cIMrBp45slLgNy/NZ4iFrrXhGqWP8aFeAb4vhW9kZUuzghDq0XFB0DfkzndO5X
LtCr6yEord4zrzfrfhk2Bswa2PPdAk3y1fvwMJ/TqT1eLDdZJcR2UFuHTvrDG167stcpV1L5kq+D
svBDU0B8YQxYLCWX+HikJufdHMcb83mQx8v21l3xHKlmTLX011TfQs6wRmy6t5mnlTi6Af993xeY
WG/2X6Ixg2YEIdADfdWwjQxYFfx9NqyAFBwpOlXX0djf7wg0tUuCzOp0DmtpGCNaGFfECDYqjAe0
X3c8S8D0ro4cANmwMM3sL1pBC21UyLbaA6WA0QaGDm4k7gbHvGNI0OW1f88c0QUt4npBGb/JfcFG
cUSQh0mi3sTwzukbSECBJBqpomC9gC+gawuElpjfFzspDSca5ZS0gubVsXAYIUuv1547EnQzOKd4
Blu+vSm9dxiEi0Ec4xsroiPTr16A2EYJz5bsKMneO+WqhPBkvWeMFHrG11sqejKGhhJUt2xxHGgz
jv7wbEOk9ngRRn1aeALCorKzx9SwNJ8hkxE2CaRFiRSEHwC5KvjmOXlYnlBg7dyb3TBCUmQNyYa4
nr6WpIPvsH9ZhYQO8j1lr93XhHkhisZxfTuBV0CSY6d2xtrSRNi+9jYxrol4//+yL86oqBxIgSeX
Z0loBdvMHSmLFS4f1opn8+hqBS/HlQ2RTHCkbJVQytbEBX2avfIqbXwqWshUyq5EK8+4/wqdCS2K
n634hM4RS8QRiSs5Dtzi1828UpxVHBINZTGWXbb2F3weKiHWc9Z0Wg/3tOqnYg3Qp9mgv3Vm8fWb
YGdw+/JwfPaXk07kz4LTltv9WMCcj2oh6lUAj/GpI8j58N777EM4PIhlHSTbO+MO7ZRbuaNUfxj2
g/z+Q8IjI+tTg+cOkSYOoRizzDMQm/jX1R9ykXrC52q7ICDrH4Y3VLU4VUlO9RU+4CLXz+NPyiRF
thsyGDLnst0cAPg5MClXP2gMWTuxI/H+4+ZwfNT58w92Sm2M/Ns4lqhfLJ+USmUDYtqxdUbSaGoQ
fqHUZXF7OwmVg2bj4qQMgYT2wD9DFR0FK82+nfWjQCbqF2AjM9KvXPCDf1VJRRjNnoIalFroXV2b
lxl2qnl0bhmi8++7lcyRubJyLISK1YXLqTOY9ObLGv6xAEvFiTLh4siGmcUdPSVBXKmoKx9UM7Oh
UPvieKlbe0g0e7G/Evl4cG9wG1pzkytUhqfpIIaDWoXd8Ldva+T97cgDnVM9cEru1V2bj8yTDkJ+
7o9E5fSaf5DcnGaPEwjFRH+amvzqmyt6Fg9KcvZ7cxH7mcrFjy+5pHxdKK9+eqxzhGbZJEqidK++
ZPCKOGZJp9lS4OeeJpNFW0xilHqFMmqxPzwEiGUz9Qi8ElUd67ygqpwulNLClNvTSpGz0JvsMqUt
V9+4tY8SRPQSN3a0PauB/RDQUUKV9zm6Z0uKkHdvrxo5iYn/CQXRkcW5gY3Ugq7SmYoOWY6itbz2
NEJEyFxQHUTdHAqi+ZeHknXX08HBNW/95saaMTBsBKMGBuTqXg8+cQi+BPIo8WZISAasNZ8OeZpi
c+8D0WRsvBYh59g404Ss+Hj2pNPsDJCaBiV6KwnRRPnqZOZD3xKST3ZVgiQDNaq+rZM5igHXtsQS
8aZ1yol7FOPIqltfGqMX+W6AcPUOoSM+hZZGiTwpQll+BftWblCr7W2AyPvgw9qUedd9VzW2q2GL
t7TIjR60iy3j0xK44coSrR2R7k9Ye/wlPvksZwqmaEh33k9U38m44pLVqG625E2GZpGpekTbWhHf
FpQKkPsDg687aWdtO/Q4r5AWoXq9hapkN57xsei8wXobLITW6NT0gBd/QwokIXopw+m0MAJwDU3B
/y4X6ASJDiCJvbG8LhOIS9qN+MfiV0eOxVKuTAmdHenBggpjYFeDEvg7LG50UKoOzW294Lh9hjbq
74hCCmRIBimkCp42Luy9xFWmyLMTEtASU47SPt2zupwUpbTOpv0dEEFETfLAUqly21ZqQg3XaZQ5
S3lIo1IANsP896GlPyisVaUyBv1bQ/R9aoedVI5jLORBI01+xvH83RWE73kPpHmsFWvbUMpF/dDC
wjZpcU+rdIyotvIW6eDsAvx+sf6wBsjTsbzLFz5QppWWZKJUDYxChAe1tKlZCIzBCJXfB/Tz1nJO
8J1fh7o66s7yG6TCltu7sY3ywaaPasynA45XVXQ1tqXw7/fwIUg32H/my+qY2HqGdcY6KquzwbmF
8mXHV1/8MVRVtW5lDPVWuyIdOZVSswXwS0vsSJmSNBXRGSIJdRJqcFGZNa2C1EnCWy+XYJD5HrWF
8oK6ou83ePdtyVIHhZD05u6NxOWxtPYwR2FS8zRuArR4z6afVJOictIfechjjjyF6baCikNtQ1/n
E1Q/SLtia9Fn+E6n5BaAIQlDYc3kg6IXZcEb2PqRilK02ev73Bxi/+UQqfQbcEKAZg6lg4r+G+4H
qlEBpDUg9V0eSaf3Re6s6kWs/Hevcciy6YA5SqIyYQGyuePX0slGiF3f1WfKkm/G1CKwiZnf4mqZ
Zfpx4khNYR+TaLo1NulOxKl4vyJwtfQM3lf2g1TJzbu8F7oQIsgMti3HgsLyzyzDg1/BdqT1LYeY
y5pGswpYwnlz20/zNOYywN5saCb0fix5HM6LFksjrO8INGO3+YTXZLPudncpD7B/GYZhLduKRJFa
gkBI61D82sHJHTnoAiQswLxW24fpKBbRHGCvhgugoKlVYjDuMCPb+mdOJZ1Q4sk5Pj7k2B8GVCIJ
1/J18yeUt/XqMlR3B0r2BVeIZI7Dnms0jNbUjvTgl1B5Af3srPbtM9Lu3Rvao7ciS2/zBohil1cZ
qENKSwUkDGmeOm3w/Fyc1qsLE9BtgfGo8t0sGvFc5ruMor7t/lNwEMGGIF8W6ooghV99AXqRo7gX
wQoF/sLrfl1TY5fFjbSE30LXW5shgCul/WdQIT80vresVROygb+oL0Oc1v0JX+HsFAlEdPZatouB
RDiY/P90rDNuHAOnxZjBKFG351/6N1kc8E0Re0fD0R6uKFkn4kKW31oqrb/aU/o5oa2w/c7QNBeh
NG36umooJUvNFMfqSaQFxfbhbeDhds7nxDOz4kTXVM2NqQkXjyTCsZ54MKHb7HKwcHVkiSnM/TEJ
St/ZEUjFmbqjLD51OCw0mwg3JbAJOdTAY9ZUJM+Xm3EeZny87n0zdnFdC9ZLztYztWlbMom0gc6b
ZVByd0mEd1lupjFJf+BypUBhEa0fxN53v02G4Qv5gH9riOyys5Nt4xEGYxfYcT5l2rpngEB1g1WN
GFg7mfm+MEmCdaNx4nQ9PPclR1BWzcPtF70dNa5nsUDRhV6kbUTHSPsL95t/VVnOLBBuxxVvIKf2
04uiu7YOHZgMzVRpjLCKa7YzMlmm18rsXvd9xlv/nPJ4UD9USXxLyUCJuNNzvz7kwrGc0SwKjYVJ
X3lA5KTDjNoY3J2EbiCh2w+x1jTjbNFFjKf+ScaRs7U+WL5F3NqqdI872MS8IEZSM3JkKRtertFN
cvwzE0D4O03m5YnPHDi7gYfExMjxSe/bj3EAwLJml5M6aZohk/9qHVzYVsLTpuC+XP9h28iPlGYi
EH2HD1jxUYeBB1ZzTM7KzKUFhVCVkcPsNNfqkJCri/qCIe93aUJ7N49yoU+Dj/mu+UVhmBODnhU3
QgbaVX5w8ASVzDCaf4G3CqXKZ/MRdTNUkulyxvNy5zVorJrj4HMpGB57agJIa2wWDkHDV2wgco6I
gJ2PbkFdYhahrnWZxVc3QmI0WG/GpL9JKlgmfQVn8C3kXfJCDLGvHxf//c/U6ytR94wJgfI3kOus
SzynYxpNuQKKMCI76xrRfk5jxF4I5DqF/W0XZ9om3FYxOfJwvYodirN6UIS2cufcoJhnDyJO7evV
nAXyGOM/9ehzAzw+fGzyu1eRfJgk9FUgiZ4kan5unCDGi1yh3aAhpgfZm9DqN+0L9wQR69Xqf8BP
SaYVMUz78pn1ZwD+zbNDDJdit1fFWsmEu7i6/J8NUwUfEJg7ldq63UbAik+dVcR+R4UyDSbDN12x
SguhoGrjuOM7iqhbt+akGppgoLYqP0pgde6O+OM1YdLDIkOo0PK8TWmseDWEFMdckL1McIoAceQP
TveXKR6uXzA1a8H+5bcPERdfP4zaIO2Dy7EGnviq4EXHTy2rG3xG3wQz9JoUPkaiospevyR2FR/S
f2WV4LfWIxYSsF0AH4TEwtecHDZoedgH6Z2kbWaMNwRna+TOPAJ1YiVSTYkQ65Z9CLsibB9piZVQ
oJoh9RI0qf9uiR+CUMrjFQgGx0tZwljrKuqsWX12vOtIa6t6CgNia1LfJhW1CD5no1tEgPUxOChv
F5acU28p/pD4XV0/r+FW/scj7AxvOQodojE90XxJi0uGP+56CEhU+TOX1VlGIeZZyRNICPeehAsO
1czaQNkON3m9aVhwZ8/TE+3u38q8okZYgnGtIRBnLn0eCEjyjeAz58hG+XvCX/Nv9Y+QM6vEuuE5
+w5VyFtpjbaHxLc/K7q0DMz67DQVZxUbMFU7k2oMw+IhkbkHOqdPQm1E6jNG+6DSzS+AKn9PJtG6
+rBdgQx9blfjfcAn7WszZFyABHkCr9Ptjz5yJ65ebin3oYI4U2QM9kBs2x/NAtRiXTiPCFtE92FV
WZrdeavblqmqTikd+NcfNJfz45nnPzjPKo1DKCPujp56a1L9LREGo1mlYQ59SmbgRTC5TDEjBos8
ZpSz46B0hFbXvN3Ux49LVY+hRhPlXJjvYKnmWjtaLPdgDWF9E0fdSdAmLMOzfC4z/apapfiS+18F
/0M7/yBXANLG444kSzAHU9eFE+N33AE1Br9E4LfSwKjTNVh5PUonv9cvQ4ymlkVZ3t/FF/Zzik/+
TzcbrMGVSYQLWERAaDx36vRb8weiSox8rb/QEPk3N5ebaBQ9UCA2aR3z9IP/377H5t7njGUe4kjj
SZ929M4mE2SP2eGSwtsT8yNiB57zAJcy77VE5183AHW7xboTBDuQdoos+q3Mkn/u1ffp3c0VGl73
XM5SytsSXKLe4is2/b+WtG9QBI1aTyicaG61GfBwaNXCsva3BCrCFMg22Gtu7pdcm4M5ehDoUeT3
QfJf3xMCoJn8nehbyqvWcXlMMPH5+gyHZcWWZ8mUkLYaaQjdom5Vk3XOhiO1toGmn8tZQZ2wpEan
R1/VprbrwwE3BSp6Ogi2JEgUsaHVIZkyaxSm1sxXH6U7tru1IYccQH/m3KLIBIccrHPFwKXCVP6a
kiVJdlaSyze8ldxYGoACA3PxbBq4VwJtD22naslHl+MNqDOPPyLF7njArw/EtfFmucgecd2sMOgM
gOVjiY/A7nrsrks/NIqIASaWS2km20Qx0pbVu4PSEbJ0hi5hX9wchuYaSfwUluBUg9BbLiF0c56C
JuP63cy3TJvXe2+z6x2hkqEtrndYMSpdSt+UGBY0m64gg9ZMPjVMY6oplyyZYqlfrRSeJl87M+o0
SLwsx+7bY5TrnE38kChxvsC9M0FnfwRkKn8sGBjHtqTqimI1anWjny/7AMPWaD4CGcI7zO72Kjrv
l/q4LsPzflI+xcn2EJsyaLosxeKxRMfZUEwPF6hLb8jN5H7LuObu2wjToF5ULvvQ95qQhmFY+jHu
Oh2ReUl02JG1h/lDeny5Gmy6l4LmZOEfUG/m5U1ZuZuGu4A6McMQ2u5tPWvycgC1mLwO4VnuNtas
/qJ1UivZFJFVJGkoi0emrJc4bpR4XJ/e7dkEXOq9XzuxKl/J2TCg4HbYhyCzzWRNRADrsSWRkGIA
TjZjwFL9hXYt6idg8MEa8iPtLuvXgX+O/oTW1xJxt91jW6HTI5dFaPbtoxDwMErCUIdfn3Mvr7aZ
dxo309yQwZwlZOAI8bU5S4LLg0NGry6F9uaWF6HxlLzBqaCHao+a2S5RaN4qi35IOXnUujlNKMr2
UIsTXdi9BFnna5uzM69JqvYXAqQ6/jBag3djih4lj8eXtDNgb6Rv1hXrMi+v6oRn+SdI9pDS1WYx
48du/md3qUZd16e7//N1VRRWpDuqIQ8Oy1kyyCTRJeriwctqaOSFs0b7IHVtF/cZVvg5fwLZoZ+v
lZa2WoBbO0Esnj909ofakRry9atUbQL6N2gm4yfuBxCJ2M+GwzHJIavZjHiSnYk9ThbXxioSI76B
gi6QYT9yHiTgvrZp5l5QKsWJ+8EjzDQLySkMW/baRPgYXrA22ipIAyqhHhKSjIAVCqURqMH37gT8
rE4W7ovL2GRycA8h/tVnEu6e4mmFa8Uq4SOqCFxNOsJoxktPok+yRycDluF7avD1KgtCEMjecvEu
Ou5O35ANsLwOl7jLopOYNZ0xr7n+HnKu+ILhSlWlaHUHvvHdfN3VM44HTfJlz/E2/mKiZCHGtngT
d1X33M6KKHVt4JhbOk5UHoQME5Wmds3jGbRozEHLfWuJFl1r9sqLz0423fNj2xGq84baYbzZxqS1
g/4KhWxwLMppt9/vrh909KgYu2d0czyl5lJ9BT32xI8eBmV1g5g5fAsyW7nsOT9mR+EwSY2OAvqQ
qTZqf6IYS+NudJgBMzbZhYEHF9ASCC9Ply72XsKtj+32D7U3FC66TeLHGbXev2Br5d+kmCGKNWkV
H0pdxy5gAkAs9PXH9GmzSCffVq+m48hXpEFgV+Jg6QhFFKCjvjSFoC4UCwfLlfO0hvlCJGYdd2hA
qdbWuFeoWW3C5fsEjf/u4tYlcKLnGj/FBQNDv1tHfgK8vIwz8XEp7TCzjr0eYrSroc3iDHsdbVTj
Qfe6k6pq32gHT+VithqN7Phdg0AWVSyiWvdv2Cl91m7pHYSm4Xf/3vI0qg1Cbzas8CNjfLivCXGm
umdple3APwGwQoSE8Wbyf2tutITKhvYyYmotjvkJBJhGCUkMDA5ejWXgVUOj/ddYO0tPKvEe5apC
z9oVETNtWs1dYMgYNoQ6jmBBVDN2m2vPf5/EkajJBH+ce8HAHD0Zpp1lYisevZXAxCsKj43kszwP
S/Ct3hUpQXQuTjwNoe8TfimrjbBM0JiedC2HBYp+a+49p7NBSjxmvjO1GtT+zJDJBkn7w8lNlwFp
cbvYHYUseEBoajXTcmd9VoAo+4yfrSFxg5RaU19JFQt25DqFRBBrzXL1S6z+4UmwlmN9ceiP1uDD
JOtNwXbW4amtv03YekgUckXz9wZb2MiNl0xLpbZivrhJFtRrj/9VLgVZVGzwSpyUBsF9nTEM2PBd
ljx7H1Qyle/TeqtsK7qz2Rg11t8tB+dR3Nt1jqBJRO9WvtuJZx+saeNrR13yNKkOOBdgP/u8ZF2a
nvuYqAO9pVzhlizAjJGAR/zWpgfdAo0aPnmGUBAGch6hdZuIh+qAPpdPNBmyoHc6VNTNVO2j8mIJ
EWlI+5ARpLVBZpYzf+Q13HvAHotR8s70N4M4yqxcDjltgSzFTZWQp/2F4fCAiQo15GTgh8Flv6vq
kh1h11OUVLV04uWrmFoDll4Sad1z15OMNvxXbZ9CkVPBS328MImMfNLrNPADfMUsI84Xhy8bSmBq
NE+/8PwnJxLBSF3in7sPzDP0VR5sCdDbmi9yGrM4jKkAwn3Q12eh/eUE2bZlW+cpBmyhMf8NoMeQ
hCoYaw275GdU2H59drRbJWvYIr9TII+bkD2TS3LYRYes0FOcJ7dHYC9R0aRYL/xgg2Oh5pAuVWUm
20mgPDDJGJOpB/L69cwPTR+l0hM+fbQMkuhs8VTr1rQhlTaMb4JZlzD6hRtElWqjTmYdS8GSUMyf
myaQUQX6BtpxDGw8dW42PXo2Ky/6n9X+p3jhpRXH+vamLYYcusol8TctIxJXUUWMhH70sTmIvKdT
HC8YlHjDgEztUqrs7a7ltp0tJPydDztDS5RAxfVJlA1Qv08FRY0UmDkjhRrgD27U9s1htbIQk1UQ
FQBNcnwT9FIjfJ7GSfY+hjEPVgxnvqjYO4S6xYF4uKM1QiGu6fsDj7U+3OcU1ZKYHDBZF5DceL8i
nVttitc/7Zi99s8ifEJDiOVEx2bt3rQ2xoYdm4oBkKSS1fUBCWil1eW3XBMAW0FV50xZBZMAYvju
diKpzaCCiZOUeZb96Tb4ZuSen+1hZFjWT7q1DgeWwiurvzviysztReI0j27v5n8woUJVvQcg+A5d
rA5LObG6cfbze0JH5HXjvfKYXepOwZs9WhdDd26CRFPOcu4IvURd2pqab94gdhLf+2v2AQrUBd7A
52rleqhPzmKPrGE0JNTDyQR6xTq3shOv00qThOLpbovh6NjyQ8LF1KR3eWasEORWW5fFZCDQvtSD
TTQje1BzN45eYTf7YzOXpmh+97irYe1xSQ8pT0FdQvLDTs1eO9o113qdj/e0S7CjxBEQ4vY8NSVc
wodeQ068VEh1RSFDAq4iuAg6eOZprNkgYavvEhUxihvvkJa+DhsQVJnyZ7Wi6/0Hz29JC3MjVC8a
8K5gnttcYmnl75Z+7y+BJ49wh2kBDi/brVaQrT2Vqe1LurZ9n1P3HqqeCygmGyPIVIbKWibEptE6
JI5Fe76v4HQeTccS4JdiScxS48YN3wtjWm96pzHgRDMwGAD9o3vNeET8iAvhKv2qu5bKe8XRVPt8
alUGlULMB6GriZRnbCcjzJKhC9VOA0Sf5GPWqhGRpUP62fkldwS8pMXFkUPh+tc6gkutesxAM57d
uS1wGcMb+5cbWrY/k4iuOz4GNzFQqeVaM1pDzvDNCzd7cHdseIyXWaZveXlYuS840abMAbUXGkoI
eoxnYnx6HbzcC/Pr+eAD7QsChn0QxoikMbVZpBlkUICodAjSpV+FLbGlcpUQhFmlRdaI7fRra2ZE
fUaiBiKI87PojYf4ZuvGbdMVyDqeBElQK6X1GVfcPgPuedVhe4wooGv/wGIYzWGz30z/Eiow5SNA
14hfBD5wbqV7gNRVFsvZCaPw5KAPw+qBUFUaOngXho/RQoZqBXTzyLo3UuSMev/5aDNTfSH1WHH3
syRtHOjXZMyAVY6GknkIB3e417iD38IaMu5eZk/xLvSd2Qg6iSlX4xRNODZWuzS0M5ePxR7l+X/9
s+qFitNAB1kumHWFb/giwMPECT76TzWrO7HPqAn7HlJkwUCECrHjmMVJtkpqs8U5kB26zvd2qO1N
ffZlybN2L5BP1pJTnoX7T10YMl2flVW+bPqL3T6Aj3+W+uQilzquh4uZfnZF83CUZBfOCkjbulPS
Gbkivw+6vbxhQJYHSPmujiMpJUksstkXzD5SGR6QGTxwY0aFctJkISbjKW6pocyBhIkHM5iJ0hj7
0xqaduMhOZxptaJj780OoXrFqeDcAYJOjU4zBI8dW/ByYG3YOx2eJpjHIP54usgu5p82er/HnNGv
JDUIv267a1U1SVZzmpFLCANSjZPMreGkTQiEuG7X6szbmqFHNPJyRiAIUVwX2eLm7VMB1ljzMU/1
XZE+/yIVXnPszo805/xBSXFgg8Ckv8CUo2Va1hZsKW7JL5+vtoflxspUCSbO304vWJny1Y4A41Pl
Fz7OUT8y9EM33ugwzYeUcolg+prObV5xt2ohc4NoteTsyq8HumLaz4/gVxEYKb20P386qshk3MyJ
kaT6X5eyJ4qeP/pSIX66d6thEku1wu+1cSEiq7/LSHVGpV2rkKgcWY//GK2vEk24kSOdU6pne4Sh
a/81Pu5zPg1jOPbMPinGtjeFtTTVf5sXjHLf/rh29Zs1jippkZHGQ8VkN7qyjo0pQ3TIYVdENqF+
wB7E1cS+xm2cuiCYByanmyxWCv+UBgp7vW0OTf+9BI9XSRBGLlPsdXNlJnuuuugi3p+2O9ZLxY02
gtuLtyVFO5+ssisan6gNTQjYmh735V3CVuLbQ4foi1Y4UOZnSOmTPwI6kGs7zMy5o414T0dgFqI4
hI+86eovA+LpdZXV4op6LeltpdLfp2LVHS7gx5Z0Mc4zK9P2wpqOInZgXC2tPfIqbj8ldAKyxhlF
g5lIc0jSvaa0+fuLT7UozWJ1NFFA/nK6IkzKnssH43fUSLabpG/uDRCdySYc0jcp3aOfaZ3Na7tn
5TMlw6sUq0optFI9gRVnoDgC6qkQRCYKwwuTjEEdEahM2bHjYQQxlvp0Xe0cEjOEaAT78W1NS58q
y4Dptrgs5tm1+5naa9KmrARCahUYw4jJljzZtLn4QISqvENbNKTk/ok2lXJyURraSh7+xU1gPHIG
Fa1lljOFQtqNYOX/za2vB929b06LzdcLuEFHzJpHn7fehj5uA7Vyx1CwCvJWHU/BNYeLaaelmXPD
LJADtC7MUu2Ij5v329BRj0Lak/EoUCRuuEPsGPSD0qBPaRM0mTDyHM2/tChI3Myuzswrmt5WGz10
XDx2SVLgfa7u5n5bwLaOAjbUtIXyAFBpCpeETTxRfVdIh0ZeTNgNPETWWopq3z7u1lXJppu6bWKl
gLBw3mAdufcrUHx/IiKidQsJXMzYQlS4tEschFBNg+wL1e8FIxO/gC58IDOYO1emLXQnLS3uXXH8
zrfsNxgj0xRXm23BjClY7dxhC9f/f9LbOG2KZusz+JOxXMU0ZyyCfbeu0gm8e6gHt5jcPUbpd6cD
qBdcdYbYEY9QZR8Aoa2HKLZqW1XgWBMWSNX1o7VW2PgyLcN8BWwFsdwL+Ph0T/xeEtAXwSFJ+CyU
dQgtbkSgfwrw1mIWkdKlu/kRA5ZzhYPCaxTs/dFww/1f9hXm3A2xYBBcP5YTjrIPz5TQgjD3cZyJ
82hhTIhsUb+cqsIR+WdvdqiHbBWvFDzsRrIDamdLoTlmYu/aOVrRxl6236lUCxNaXpjpYQgvtK+m
illbVtByxxNCYycSSKgBlDg15CfCahVGQRBZ/cxNPihZMeal9RkTMfh7cveoEzbXz/taJD09kuO/
6lPqfu1G5oGft00DZWkux7969AU3e7Cvs/0JUnFRAyhbW3NKGdwcvmAOhk/Y2TxKsWkDVHUcajiJ
vsKpd7KiYpdD13G8wl7F84vGa41VqrKdDbMccCxB+inNt5mvKBaKptAcfOwr0c0eAlKN7OfeOeiP
I0SCmBlgE4OCJZ8ziZ77lyFQJQqmzf4lkzBMp5aIBR+dR6cLYlpm9RSmHBNFokIgokJFZpAZT86N
UUqPBIy6/mUMn7Pds6hXTUzUVAmMFL4T6VjWinw/z14m7ihy2I4C9XwSjmDAOTwfs2sUZy5qQBx3
SrAdFH5KOJASG86uzjvpkpuy01/ks4Jaj8dORt2rkV7HmECijjb97RKFcP98RHYxKW19Z1Q1xsF/
f3wE1fEIa42VlqEnmh5Gq+4CAbq9TC0tGOZ/HfKWrOKiBJUBvPoZBAfixJ5GaugMv122RK2E2fUH
J/IiyLrADk4FptRMF15vtvt47+KriowyiVx22xEJP6Y+zjezv2V/MBTy1DA0Ka7muwSRyayXSF2n
aeod96HX76oUbSARzv6c836lhLKuit7qt/B8YQ8+DZTVq5+cfNEoT4lua1T7XwLChxDsq6tYwO1L
q4OED7TKv7mm0OOyaj71XmxBVdczuhi/mnmvoc+PO01ijUVlhLzh2dh2Y+E8KN57XOXhnhtj21mx
G4PJeiDEmzJhXvQ6ZEzSbFHWcFh+mfzOU4JNfkkEYk11FIgtSNMxgh4DaJluU9lLY9y8nN20D5Ec
L9pUzoV9ipTiGd/9gUq5JfPC+BmKXiBuZ+5/ct5Pjtm4m7HQaQKSvfdqI0Bl+7Da5qZlnfQ11rGS
/m1ZrFetx0s/Wn76vhsCAny/c10AFMs8VenUkZFrxuOjZVGm3IpY9gA5TAQH8gUuDIwunkhmo01D
iILBbMDU5esOmhhdf5aQUh8rHumxgWC+bYj1eLkJwb82ybe/35Epm84DWGecTG7ajcuXNii+vInk
ZYHE2TvIDOQBfe6JHWJBdJ82YvElM4gk9aZsZGBImO785YgZzZ+DtfyX/AkFIILy42edH+AMpMo1
f3zSQfAF2yAzqeod5yTqQR5S4/G6iJz6z6ERbe04C93d3po282lKD0zm9hGkZxK1+/A1B3x4xgh4
qEOgrv0SVTf85+rIRf2XowwT56hCuiZ35FXOfG0e1CIjuebzcpJoAk/bNo1MaNlI+alZvTFxQp/Q
o1MUu4Jk7L4rspLD7MqDXlJ9XvJGdXuet96KMwt57bjrH5Xe+RRoh1sOoQkxRP0G4kyi2ZwBWzMs
6RPtWfUN9X/Zid10/kPYF7o73ZPqz9A6HznDE23PP7zaKvqt/+2mbc8tla0YZ8zPwvvXu8YAewjL
gpL/9OCa7C2PXmUkLHyvU58iUBfgLibs/q5Tb+8A/Fs9dHMKiRWpF9TMT7+9mwqidnY0Vy0ICNl1
ymj+Gf4+2ClJxQGPAiG+70uCtXC1j2Dw4ZUiKIRVTD+v3NQ1GkZL3KdYmL9vtg8YKhQ6S2M2pJBC
OqDqi541AilYI9Jdm+i3OwT6uv7b3e3VthA+e6f8vlE/BaFnTlic8XnA4dINHg8Rt+aR/HRdpuf9
ydpBHRVMof2h5WVqDJRC4nCvnzBYB9n7OSHDctPK3VvJzDk5t5SJDEraX91v58ko+mxIhJML8MSz
7wLfK6eyEO074crVEXuzMvGlBL/mSlJQ7/NLS4N2hvJxaBtYi7H3+mip9ncofxVbtSIl9XSNcUat
sWlkOveuRbtv74IJSyP0LXaKs+uUbbHGQr7sD67JE4HiIgHqaw/GursF9kFNmFe8lrYpTUPgI1zs
cS7HnFcIoyTUAFWd7wTDkdwjlE6zqTJnEnjQcBBHh7G+RlZWJc1tCAWGanm0IyDhYXw9dCIMd3Lz
XYlI2vCqGn/LWmuEbDonjdT77Sc6eBhGL2pVeAlv4uct199h9aTUo9M45Eh2InG98tOxMm6+urG+
k2Gj/plR5rStF1vFPI2NWpqorbHINqmqUsH7/iz3WM0ctilvz6YcRf6RUrlG1NcAPjqh4hK+sJ99
J5pqaG0PtB+xbrlteCZh5WG/OjH6SYJZnmcj3pS/GzmgO2eVV3+/rNKmq++NUsGuWiA7SO8ATQTZ
12R5nYG2vA/xzVJq7h0NBwtgfzSHX7yeYnQZtmYBxXXED9eBYUOjj7KnFybz1DcY6a1nZ+pbNCSU
E7zohpKVgpIh15Zt8fBpP8WFHl8woq6td/FFGrxsi5dVujyGgs2VlXIGllt7yS8xsLYJ7WhSbc8W
U5X0qnyDHdt17DwgbXWVEy2SVMWzUHSwjybIk02zPN4Y7C9os+0Sf4t8/qADIxK8hfC7Taumg56X
60+XkNQMfe5CZgYVICOf1C0FwmDr1xi1aE7IrhRJ2yqxXEkwWq6atugJx87ogBbvgTmXxQJOaKKe
2xkYD464r/MW0eWN0dHzVyuB/sCfdSLsfz4LFUdhWOgqFuaZ/v/MaY8jBZDB6vFa0kpG4E+6TLus
E1QD2HAi5hC/yg3OYJhfa6OT/1giga1GmVu0AH+vHZZs6waxMJIS7YzBeExF/8ci/7zpeuXAU98s
q7OwU1GUu+FmdT37rCz2N5IhUcetRG0QHD/WmCO7oKPt+1qip5kpOq4fL3fdnRJstOg5eR0lAK/3
RWGGZpPUzvOfYReQc2cRIPM69zxtXr3o4cZnAwrxiwF8OC2PramW+akky8mM2PVkw5ydTxGyQnzI
OSh269LaUjJjPsbsQeXd173wr5KKowaTN6b5KTFezl/AVIlvBa/57lz2JS619/CbuzMahz6Rx4Fi
4Q8MQbhpyicadv5+UY1q8HLqGukKux1Cjju7Chhv0yF3Dra4HhFrHqQEYhrjEpy/1bbzrGWvLVuN
mQojd/4ODgS2W9dNYGcfGwPXfXHyfKWvSJshqzg8EuoulUgpGJ0pettt86elxBHmnBELMnAilDOp
6f9iLyF0sn/byirLOYNpQOP5XtjhwasXm1xZhqga9vK5HndXb24tyOuOKZWbPmeRJw+708P6hXld
mqAhw6I42zhwefRCYwqXGFfsLKEEB/LUhqTITPWra4wetEZFNgn0ALcha+hKYep2raf5OetNN/2j
50bdmeMp9BDyB9s/2Otkvz/AXzrQPi5ANJK3UbmKCnhNkC6cu29hTSn+wkzuMhgHWu3YveQ/G+IP
fEeOo/VqmaHFRucj648sFyxTvmSrDZj7CLqIyFfGxUt7TREJCWF5dOuAHKVJARP/AzHnY97xtshh
KPdvo7aN27k4xCdvwuKoHZGJb3zi3g8wToJKgVL/hGPNnZBPwNXy7s09gkAO4bASNZnNrElXTjN7
KAg6whPkjtL0teBvpyTzPzV56I6SKQ2OVT+xBC5HubnXfDmrWooDUoBdHK6ZbwOLVUbtRXtwoXlI
ONTvchYxMNYk7auqwY44JbKJ7PMHG19I4MSnLwIhMW2ZIb4xl4Xl9yr5unbFDchHyxP7mADK4z72
e+hpn4wXLm/gmfW6dhqXgQsWaqghhs2cf2KszBNgtuGQAK6U+CsCfX+NbSUD5ZZwAR9+24/yWCKu
YrwuxKIV59MZ+ke2yOyM/suKgt8C9KqPUoTFpVq0ttpnOS+u4sxLe8hCgF3iSDNWiN3C4QzWPb3p
twn7MCz0DkmHVkTLYyNDwdGLGMbmllQcIrlMX8sJfq54pmv/mFJV5Z1R70T/yPtruXlf7cCVLrQB
BHgBkTx/WV/NV+E7HcuZBnQMxp50mVozrxTuQW8wmP8BL9b5i5f9+mS+LUD1saPS5g9fVviQSXrJ
X51DCENKMLUDl0yADsPgCbKS3lQ+OakHytWXa8s525ShO8TGKnucDnLu0hqKLNdgQ714ZmMm9Zev
BWwE4H7cNFjp24wPDbMYhRx8GmWzz8Ula2yXzbCnrlMvKeD61d7FnYdrxOgLfBDujK3u3BNuziN/
18AnzEJ8OvNcAFFyB7bz1mjdNCF+SCFvAZ6My4LPeRZ7yET4ceMmaL5tZ9nEmsXR7WtMN042DVV8
v5ISzNvIeTP+LdB3ImBOi2h1q/2B9505HmAoTF7+txQp6tCmpd3tNvpX4RFxajNRgD//NH4KDV0N
pw56H8MqE44ySNVHZLjjt0vuRlnv9cLsws7/gXNwpPOIlQ/XG6KmkcBact4nMpVqsj2xMdl7PTZk
AGlLCUHQIgsPE8qfrS7H215NiviOwvarxnmJTUUoHuuipQvki3Pn3sRRWQI24sJRqiUI9/4xdxQy
0PxVUfhR73UPqO/tlJfXckNpVYeiungz+clBRegvvHTHm2xfeJ1sYFnVTFQI/j1M+Iqq53Z9i29p
SG/q9Gl/xXcLRlYs8mEVlALM0L5GfXi/VOaZlO/83uF6LmjqYwNaLgozEJr/0/Pk1wf6RmlSjCvk
7hI7k9hBTy1Z83tFcSDtorvFzckYEpgXRZa+ZNyW8kZ7x6nIw7EjAHwcUkqkM5afOYxOxqnVz1Sw
ZzanVz9oMdR8YEr6uXVOqhC+5NEzCUsuPd5U7IBFgtcCh0jRf+1IsED5wJIiUtGTa/AJRW1BrXoI
5jQ/K6dsJxI46GMiHDB6c3qyfTR4KzOr7B5J37e/noV6PGS1hMRKqNsBHuWKEN4nUIHTcqw6EWr8
9EH3vcDGXJz3pg5Ts2H2OqgRTcbZFH58Woeiuid+z8niDgQibhG0JOQGcrX739W7kwfJ2hx7Dl7M
U9JBCT1gNLkzqZD7hrfYrrpVdUAwCxN3LNc+5hB9MOkYsxYRz3151CYrUpHdcg0iWPtoAOKcBfyk
UQ4ixB73mgwbEkNeMhNC2Pt7ZoQs21rDCY4PC5oT/NTZqtKSaXZaUHQd4SIOkWmwQqNeOS5JIzt/
mzJeR21OGj/DXetaorpNEePeCLnpIDopuqeD1hsAUf6D3DeNbn7HoVN3v6083OsKWswrgWxniJNr
DEQoMYvWTACaczO1ZVJ57IrkbFVgk1XD+W4ydt2UXTxJvD5LFH/lqbTd/RNARgMbDUjUsAGqQhqU
KOYlZLCLbatxtwdHWeq8o/zypyl5XE6EpuFzR+3zd6Df+CzKZuhb6koajoteVo3ZnfTivb9RzAHx
gd7grekJdnX10qcUPzz4W0cNg6RuTocmlfkhKFp+Rl6mCLDwyhoN/6yTmuAL0+gf82VqxVvVNgC4
gBDNszu8pG2Yt233GovP3kOz7jDkY7FYTSBy7Lgj9RvkHGzTANdQXubNOQzaSXzfaMTo5u4e0efQ
9UwET/tzv6Nb9KW2V7bU0dPFxAGAp0IgU65XqqXCgngLJMKUJkMslRetmp3TvQjhusiovrwwhmu+
SIjSTdgJ0OJ45y8HAnpmP8fPablkX7fK83zKgcn0Ie5W3KliMQgA9Ikjw+MDA/q/hHpY38q6hfe+
KvEf0PQf2tODpZErcEAgenftMnPJOykZ6JS6mLyXaPhEY1kdDMg4vm0VIU5EWFEO6m8ufTqFu+OI
z51gIhHzO59EMs+5myi4taDEnMbL9feRCPmfxzQuWl8Qi25rCIbgqpjPVJE5xhbtoFUTyP9KVnIx
5KGRHVB1kg58AI/WuRvt9AqwAckjFl6DuXtN1/DzCS+yGInzjC1vOr5zHleUzEzUJX2RZePZfmqB
ELYTyzUCS2qcLy3bOPU6fVPjGLjrVhE575zGK+WGlriT0bBw8SEp8pTcA2hpQ2oB8JSNgsVeBarR
fKnQFLYZ0GDVvLgU2NCTMNIWPHiRdOqOYaGrPcBWDbfrBkwW/7O/hQD42JeZlkws4ETBwlYNIfKR
A6foWjVKXSGeU2iA12MAMuzm4RgUvL/KIU+XhEhRp3noWcDfuXPHiyv/CKShsAKoGfF3YiLu2MSz
wIVe+5MI9slsOW/3IFUSaS3L0vpl68m4owe2HR91P0/OcgYjtoSyfWzhhzfQxtMjbrQxcn4U1A9U
OQCU5ygofMAbIktgrnSXQf7VARgeXrJGH18mjk0BKEKG6zbdV9j1Oazp2botu9tRuKf1drBJIcVP
ju+6UjLsVEfsK6WxE/9oL/bb2Axej6ht2NPwnw0i8I92BD34xDZAL4Ww+LzfKeD+hVnUPXniHGUW
teGnwpIAR287vbDbh00CVK31ArWOigM/3UBgfEigGlOauCsqbTFVkwmb8yB1w0LgMg7PAyOpId7D
ofn2GYJ3gVi5p3kpOIz3Z/ZS/5GWAEow9AhAmtle8HGYB2Gx2mui/VN3ZwocfjlgztoLpwp5z3rb
yKHXuProuSkMKXuIBdOc/Pc6l3qAz8MOgmFW01Dz7QE1guxMMI6BO6iRXmJ6OEbdB6ArKamva5c3
4kIv3TjIWnU9snt6HvFTZsu9JlPpu86ka0SqjAS+6k99VMM2+eI4LroklnW3yOWOqL0zpLK94Wpz
4CrQMzd9B6TIyQ55FN5yvFcV4t2I4vp72UihxTjJmDgxCmhvfT2GTR+yby/MvYyu2jorzIIycB4c
8YEIUREmLEXAO70yC3zb9MGD+kEYimEknSw4FrNKjTewb/Rw1X6tVexPgOVy5NMmAwdEFpPc817i
lFnMIQYToSPZ++ml8CHz4diMsS8Cejiia160Xag0UyzDhUp4KwS6cFXpH3fEIShVnY5rKo+kyHQV
5NIuYcHq1g/WjZmN88L97ysJt5/vudDKtnW+jgI=
`protect end_protected

