

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KmBQFcd2QD+kNdok9pVSy+mGWrLkX1cfjcswOe7HQkAaL//+2eh9MyWA7iCeyf3d6lt9rsd77auE
ZHTB/Fk1dg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QEzlBt9msTE+rOcclHYmjKiZokGI/DjRL2yt3XgvDqGlPv64JOq2dg7pr5CbDR9qLFFLRNKC/Ave
HXTRb+K+eTpEPc7Ya4cYQ9g5+MXiwB7XQLPa/aEyjO3get5293ggZuzwkjZSHk+e9QqEk6Bt2c44
54ZWwitNxoUsEtZyS3w=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TL0QuMHUSOmzGzMiljwv7rv+fdjjk1oxddi/yntmPUYv8VtZjSw6bnlL4bf8+q0960/PHsqwyv81
+G8ArGsFjA3CQMteKmkfl/GKlw/jFc2hhJ+hJn1EdTZ431Cju17vFLrxGbmfF2JpG6uCGt3WAMGu
G1fJ/VcvUYAU7TOa1hY2/jyUGZ+kSwhGTZ/4ly4fqsmslNZ3EEbYgLpFAp/bY89KPhWWSJnAqVdS
qCq9OYjG5kABfXiZN18ABG0VS1eWRKOZaodlce+Y/gZM8YZj2dctmqg94KhruUweeysu3c48Ck1S
AaLBgWKSuYgiZzrylr7qBC5Dl8oBgOPR5lyerw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dhihncQPuJXJisBMfg6qt1V0/kVXNX+63Zw3PO0eub9NsIOp9vBY+EvdwHq1kfbkAnPnkJp5g5dj
8jo4ZZkQ4/P6qlTLOl2VSHJYjdrirUyAOSEdGt3l160J7/RiV1QcAcFzPoLRIkYo/SrPrmAgOSjD
13RD+L4ONrHTFwpLC+M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
p/aSq/rPYB4VskPGN3ZAnJ8z/CGp43GAjjH8Zzz77N5ByF29mwa2r5fYMj/F9VkgSkV8YsC9Tznw
lI4j6LMf9xzEX0HjWvWZ8pW4ITmEXtFV6uNX6FWbH1T9+SQOXk6jlchSOVmnkJTb28ykZodOoHXV
sHyYMhT/OBUCY+iWfh8BYWXEVyyUd5vsADHb3MkIuYdUTbUUFBhXMe9Efyrrd4jCrnlgHytJlFzc
HHZNJzS0lT/zBck+tKmXy9DwdLnPca6apjf9JkkmF7kUXw59bl0WfpuUVSCTVtnv4cgTqLL7Vr6F
wq7CBpoBFMhcwFp/IV8WLrlN0XiNXXNJSRga/A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5248)
`protect data_block
RkBvTSH8yfPz9hOEZxnt8QHEGBPqVeFyUxE6KVHzZ5KBCx9CNiKTpgiWbnegPpl1D8gH6gc6AbdL
CvaHoxa5XcrW3m6e57kHgGU3b/X4JJ3UULvSVjjU+USm1UCGg6JuewCkYoPbQ+vXkRp7xD5QaYL7
qKEDRq4qgL8P0NiLu7vArfPfqCUTj7Yly0wz/LJPMIFImKaT5CNhxHXavnvyfslSUrZcW52EYbrb
P+tnQJSM0y+F39/A2S/k7l6BUX3kENjFSia2N43auoxTigQqEU8g4bf6jAltGMAP2hn7qLMuFgk0
L6/mWZBGYaT1Edgfa9W/3tFL8yqVhVhuX76ndGeW73IcL0k0d5wi2O6sn87udI/j2pSkQZLIKQuV
+NKCwkcbaEpGWTo+2mCeWULbfgCvxV4Z62O9ePkrrsKeO4wHjwF9LlNicksiB6r2kd/XAq5q2evW
9qC7YcbSMpGPG4KIbFpHQxhTmLBl6TKe469HAskVqiEZYOOa+HTEgMUuCGiUh0KLh6N8c0zyKaol
rp8GkvDPXwslw6VS+UK63sTWEUmWMVLPQ9QgUyvGo310YqI9T7uMtLQDiMjJx8M4WWk0uO3jFXVs
evbBCrrPUZNMV/vjHX+Zr6Qi0VZ69Vfex1xNIBWRjcSw4apzNXP9xSo0E8b6AIcade1UhR9kALmn
lxqITmryV6MFGQgApzXruTRoUTvVsrfuMfTAdAtmDSJU07//DZ2bDclnZyEzmrUSAM9svKB/MQoJ
YiAHMAtdy4sAXURk3As4qwbFAUVtTqsBSs1m0z26p7SersfbaH168Jwqgm47Kh7+EXLTEh2hj8km
xAFaaOcaEXffDWJ2WtCq8Bvls0HYiQzuIp+fesiW1d0nkP4SyPXhPD3fLr1cYfiHefpTG9dTT/Sq
cEP8yJycGI9Y+vuvCUcbmyeF/GKW1r/CMTtGaE7XV9u38uDyBoGiThIhO/Qt5qorfjA8wJcSh1QT
DpwpM/Q2+OSMWbEcmiqG3JyKYidkUw8KMODHN3hs396XC6THGcYOBleI9lb45NbnsUp2bUEyy0cn
oSkjFLwJtT0jUv38k1nMBykF4dYX//BJMl6TwnbCVm4dB+SKLJzfm61m9S4yfX7Rc3YFgazV3tQU
ZvF3/6QOqVxb+YEje+Hil3QDF3QpnkrmVoyHp7zbzyDcqC62kHUpopYIaf+SIum5dz2aq8Kqyp54
ALM1WXgRmt8By/A0VLa9W0yISdKgQHpbdLXaFOw7qm43OzTRxEf1i8W/4X9ALr66mf8pkLliykUu
F64z8J9lE5pww4zQOMhfj8T2H8pJ5dT6Q6eV7TiiFDNRCYb5jF50PW4meMw/GNXlv8YMHmQxYCQ7
LCIKEpQP+XlskNpFMxMhUtFQ514zwc+p4I8fUoHc+hnJFWF4qGbI0Qa62hUV80+/kYRG04feNI+9
yIcUjPhOH5FIWuTVpqHpQrhjKEJdoVnuwOnDpBp1oKS9ZvSJY9sLTC6yEZwbISoH7wnAP6cXMvly
OhEpNJg6MWAdXJqkBlSTVfn+tqxrmrSgbFAYDnHddqvCQt+iln4OZ7BO95RyoOykNCQYAtuRjTtB
I2aD2EmKPOwPsLmYwTD+qruZRj1aV2uMAs6hLD3UifOMSk0Jtqvy96/exsA/Pe01bdc0+TzG8KVs
KSjV6vFJLbycwXgsPJfph8Ia6tbTuViZrXZskHKYJyMyh6QRaaErh8JXXnAGPCECig5e3a1XcapF
sBjDle82Rix4zdv6w0fBLtw9lzRvx3OTJ04Gbi2NaZgt7vfWcrYa1xz6krOyKfXnyC0yF8t7SAiv
avZmUliHHCF85bDsB3FXvtxJg+F7KQkTrT8b7nd55EVKorkXXGj9R1/Ov3SyGaKJc2/i2taXCDAg
Z1RZ86wfgBY2aEOo1LJIVTI8JE4fDhOhUk+9a7/4nsq3fTIb4qU3zL53IFBbgEE+f7Z0q+ASnN/O
UdvKdssB9v+t157BUpaPYUDCuGX+erRSYNeJ2WwpukfZxPKsXzoAV3479xgWCnWd5M6R0QFDXEK7
x50JsVx+VNcWmerQRi4BcqhbPfxkJOnYXW2hlKbgaJC/99vDylSdCm78+1TthW6fqYCgrgssljUs
9ZYtIhcBluVC96PCu2XACQfX6Uh2KsaJQ8BqOAsLkI6ZUqrE+jIZJ2aUiDBqs9SAuTUylAiP36h3
5EdBDPLGpDSZgrcnoNgEKo2Ea9zllltcr3D1Ekb67crkZpVLXTIi/XUHpP8QEAoscoDSkhg5bw3l
6NJSzjCTrjKoHucyk8yuXroaPWzTwZANSaPWUqdz6X0TvrvHSBnVdEg3Y7mRBAOy2sKk3TmtLdvM
eNxeLZSxVbJJdb5jdCDI3IO22c/2APwSVuNVQv3dHR3O/vjHxSbDj05fsSaDTd91Ef3YJSS+fJNq
jeJZdGwoNR7qvAzY3ZeCmcNjqZYQz87IrUzU1prLlhjLW3fea9EUTCkddEnEwi8X1hxtfnMcMDH/
iNBVSDydxOMvdNpLBFVSzZ0W1JystgiQtR8799yOezy7vTQH+WCNqFyDy0O4m+lr+erEwY2AAvTY
KIOm8dpKlpOkVp+vP6CZNtMWJewaE9b0vNn1utZkRJvZ3QKHnRD2t6yO/bJz3cg1WpmQNFpkQWv6
i5dXqznSqFGzbkLKFN6oEn60sDYrinBIUp2jcR3hQtelyi2kr2zdMDc9Gx3ks2iujdFSWyL4AdK8
iU965QfcIqfw5yxO/FHtUnyZSLD0+6BJdqAXoXG67GOot131PTurWm07DSdRCA8oH5cfRFUfZTfL
c0a2xuyHZ8fCZqoMimRxbENc0UfZbJf0fWWe4TSf/mTGy+LC/VO2DbsK9UlOy3H3qkzloJeQX2Bs
OWO4zo/26s+CTBU431jMWhdwz/rwPkZUK1WGsMYTWxCny6Tnl0aHeiiS9wNxKeU69/PjaLMCHvJv
2/rAmoaa+UV997rQzCleWbszo5+ZVGD0OKZaEgiYPZMV6tVNmNU3FncrWp2Bf7Q1v5sikJjbEgPZ
Xit/6iY8+S6kzmNJhdi46pXDagbURFyA2ly/NmvxzcLVXvnlMtYJXTU10Rzu1FexDaFVafDhEr5Z
pgANuZRNoAbRDkw4J3JrisR1F9VKWXYWHCzYfQrxZYd94wyFM2MtaqoY+MQt2xPQNJyyYrFk3VOG
CVghi1JvYpIny2zyzDeVAzfhczHqNhqvmcGz6eZcEvoXRSkN6V9U3ctD9cJMUdp5HFGJK+c9LyRK
wZEbxJjQ/CcCytQh8SzA1iDkI85grzCj9azf0HXVWcdG2axouqvrBGJnwhpaiWEN7kvndjDj1Kvc
vDNsZ/YROk9q9nevZI83KIlj2hZatzn1771h3qH/sXXmXVa/JgYQ8zHsH8S9Hk+EBLo8WcRlu20z
+uh0hHD63vkn4WkXYQ1xk2bqs77ps59+vcJxrDDptrMc23HHKUk/0Xh3oSKUn6dVKIQJfffVQRq2
zZGOK2rPToPoI8hUNVq67JtF8ZjWnNw5GJCHIdEO+JdIBwstoraI4QPXDj8QtI6PYOmSqc0Y1Xvk
sYtwXicBELZNzyZI8A01KGNFtDiH9SvdT8fl8kJBHTc+dZ2kA62UqlJpigyJoBdngwVP0wddGR67
XhyuTKioZ4GQCHndKykjHfPDe7Q2nzf4BddNK6RIMyLPazPgw07poVMq4geXH/kI8A70YJ+VoX7X
IQ1omBC9wrw1RPT9TbE+eWwwwBk6a0NmKGHgSV6yaL4qcqcp0CLkg4UfixbiySdGYSd1WpT5yelG
Itw069eHm0M38Bp4M6hjTpdyfBaK0qRhRIeLCA/xqO/Hl533piKUcjX/bM+xEMmJlLNAVM0Mcyys
NFSHK1iYgwh3ZPMtZalm0t+4mlFfm0sJJas6OzWQfhQBBBLqrZbp34rnMWbmpByDae9CIwa8OJV/
UxYZz55saxWU6f7IzShgjoMaReEjO9Ovj+Vf8nqiTZktIYrtKOrrK7alJWNlOoJJ6MHySTIIxYhn
YDv6S4SzbxWEH+ktJt889yxaKplh4/TWHzzWvboB9J/+SUFVGgPGk04xMWW1qozn9UJD9QtnZbmH
3lj5YUgAnqs1XGEMlTHGLyeNizgT904f4GUxH9x/04i73SVoeSVqFT5gTVMx/KlJyqL6Gw9+/RcI
5JYomV+3ujpmOsFrodP8aaMiTJLcVYNOkeWntMH/Obv1cZFbprJK3PKgWa/Grt7clcXcMSBUFTfh
7z5guZqZpGQbf3/jscG/zDtGKTmydZ6uCA0Y53zuxpE+yWluqKDox7LRVQVWoM3KuJex1XHQFLWH
7FR/LsVUo3+h/dG6cTnqbnmVt0+B2DPYoG0Xr7wEXiPa2I2wpvruLS5RuaidYVU6ar8nr6AiEGnO
E9irPl6DWV1zpss5SOQBAai7pWnlyOSfVMIz5bVOLKwRp0A2vUO7nLC22Sqo+NIs14fVgEgAVjKr
xSO5HZCePEjuX1FY28ZrCjRV9zSfY2qaY4tnoSLRX+2G5I8unD8db6cYw/1pjiI6FxWRu7v2/KO5
+xW67pjaAe4qfj7EPkH0ZERIlgxAavuw2+/r/8sVMJuKvK1GRt+Na+o8EtydQab5FTxRbL6woa/L
Zs0gTvBJlY5g4mkfmOTGZEOYI9Y3paamYQwSNZ4fMznDFH2T08r1DFuPMcqbDlp6IYcveDJj91LX
WqW6MJrtREkRK0G2Pm6X9yn9OMdKGQ1LQ2scEgVrz/THe5CMIqDC+C1+DC7/P+6LjT3HhgWLdHtY
2Dl8vWxJbsyojQbjTJ77gge9hGLdazfsiqscIRAYNj0DVTXMjiiQY4jSee6PNfXLRnCtlCRzu6Lh
xL5gUI0OisLxGMWex8YaVizgC9MmdG0Xkq4lslsWk3IFF552WbxefdgR3tkb7QqyPKB7HJBIIFUL
saBnyeeYf4Q4UwaRDjmKjs5cVPYe/6dQWe9VnIeHL2tKOzmLOcQHbrXkGhHoASjnEFCHS+e1Ov41
ed6Dm5g34aYq5RJFWDMLzBBC96XdYCVEjMPQNioArDrY4W7ds5OBCaZHusLL3h2hqpCIC/eOfhX5
0rhhzpOg2P/zlgqrsn8pM2wvXZbuvsDmp9+U59YSXzia8yChNd8XFrVgGnDFrdSW8b4qYdHwUqQO
BSW0aILGQKG8gDnLK1+WYRJDqgFueHac0Lh4vGTmywA4mririYun6Y3UayMQeETcdGPjtTlyyCcw
nn8nXqgcOaTBs3klNyyxfEetIJwcdwXwt48EGd/xnBuu7R7qJ34BLN59h4bwZognKiHQFfulkpdX
7MLZuxf/mozRj5d9myVghSc6Dpa/OBwI3xCxnrQI75WLKYNWsSSYf/M/fUqbG95poPt00Ne8dNaX
QyRAEbWdp2K1R+CROfWAZoqjXJhuZ+d7Af+UdecPceSwl+RCVIvq22ThDq1D7c+dbm++AriuVJbD
RH2hpMnLPVDM5wQWLVx2MjIkYigXHXiwtEbWBLkE7yhlbXD98L18C3QkaPueTADsQ8aUk0Xmirs5
+/ZuHOm/IQ7VzWVSESQQgpaEMXPBihYYTMFwS6ZxxgKJ3SicnkzMHYahcMEgsPUThlGagp++FTu0
0ksMAgznKkuMaMzID6ztZr0GRgvlw26c3AkjtlldH+CjJfijyJeCHUYUHzHW/Bcwwk+joMeX/iyA
LF1ePFweBe2+Dmef4y13vBsiBtm3EPmFchCZi6g3HdJfV6JwiEU0FJbuM9bM1rBn7Lzic2bU1pTp
MoxwhaidXMdZphraMOz7Pa2qUqULlhzxuJ+6XdW6vQpW/0UOq3tdUjaf4433JLyY1FSOWFKxLA+R
iFkJNK0ueAkpdarFQAg+gROCoL19Tt1aF5xartutIokQq0eyFmtO11qtQPbYrC9hZrn7/UEBtE8l
lGTqXOKD+Z1QPZL4kb6pWZIn4zvzvrH8FPYLZcQEZ9OBIJrULPB2z+4ukm0KeUOvUqqYdY3l+B4B
g6rQAkbcvGlPUIFzI6op2qy1QmituFDzufa+gw/9el9+l7ZFiNw2ylbgMFaEcI6I4KBWh/gO0zwy
vjOFCt0O02TNKmRenXSE6MPOv7PIcEryKPAHSRyPy/4+uSstfAqec9wmBeogdJ5py7KAk+6DFpr5
KWhOg3AYNR4oeg5FqU6ax4BlMcQW9lqlm7vCKlqs4A/ksFN04bo4aAm+IKQ6ZBsgJzLHRvZLkHdw
0BeYdvLU1Wec8xujsToMBPjHKtSh0WyOY24P5HCuoSXULaY3spzVpbt+Fw+vk0bxA+Pk2T9m5/J+
uizRpRLNdv6zI7lSqZkOLePfMyV53EB+4WO5cHbv0cEwaiRJdVFyKAbdr8tuzDYCBqZypmXrHtMh
uYpl9yFVzhoG/mg9tA/NEubb6K6XiJ7PpRfY6NXkM+pYgboz6aC+UcvIJi6Z2YeVSDn5aMPBHmJg
oumBWGW4CsraU5tgak8D4G4MZSpCxNEFHK//p7Cfq3Fqh2hIxKt9+X1tgcneWYYSnayqs0GTy4dP
PpXrLhIQq3fblxu+qiqfWFjNmE6/o0or1HjGDcvNNQVBQXV+3pExAnvy6z9fMDbSD+Pka29LJkO5
NowCQEikHnkvDb0gU6A9vwEvROPPZapox+9n95kqpV7dJWBLBNxUlBYZ7XqXvqpW1nh0RrvaOkBV
6WqdhqeJgoOeq1CNY4grco4yTtqN7RbUPhyOPGVjARnSzCJHJ6W6E86rY+Jhke9WOvK0w53TAQ90
KNHufUzqI0QP63hYkrN8QkO6McfhZyVrIf2hQh58CJ04mh5Vqu6cs3VhSRSsGdS9b4FId3SJS/iD
4QPoR2B2s2lQtz43c6lPib6EfK+O0qZtV7duZr7nGSuZqznAu7SPP5NpaOjV57W665zVdhFDesmN
hHu7mGh7ZZqSYi6ZgAei38b+Qex80Mm0pVEl8ytaDT8cMvfBesQJwOPD6U94wakoyHt81mKpTqiL
sOkyNQ==
`protect end_protected

