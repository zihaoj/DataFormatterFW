

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fAgj/3WSjBpge3uchVtDX1gnE6lYwU3Ik35plPnBc7INkwhXmFekzwlzr265C/YPIU3XVsqW2FoN
0CVd41WrBQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
RqUgBWoCMo7SQEfDigmkJ6lkcHYucDR4JCcVaoVSlarFEhuWTQt2MdfcInSgMRRIPd9nZY4whSoD
i/jJGZiDiMo+rw1ZCBCQazq4qIs0e1RmgmeDqeK/KYVr0UrfQzdfupZavc3oSEfQmohAallkX9Wb
rNDLho0zhfmvp8+jVq8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l9XLKMRG5MiOtEZOdvmpYo9l028C5HJHPZzqr+znaTnepyKu4SlmYY6FAIItu71b4jgSRH18MpW7
PMrNCCYACgViTcCHujVkz0P3kS3ywfhFIgTgXSySBIm6gWujS4+u5LtE7xX7qd2HBVjPXAuZ7LOd
8qat/wyJroJ38u/NlaTZczHQSLiNRzVQayotOoUjIEqXPJ1sKxkQ72mhbnSS/sVqCUbkQZgYYKnW
1Nxz1epBr3IVuOz9d+IgDovkv/nku2ALV9iOKAwIoy3uoZldkM0aOCML6bjO1fk7xtRqBrURihmG
b1/iCEqMyKTu3JnduGO3MxZUkVHAwMvKtTSz+g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
byrph5M1hEH2q5NW6bYhEW1dKKxfKFWeEICCVqEKT3K7lE9sudxZhlFKJwjCCt5fyBvUpOMpq4bd
z4d9dwPLdi4nW7QlVV+HOjnxSvXS43UhWGBYUFWKt7IMzIj61QHyy4e/M6XEWj8wWAQEezpHNokX
87dtN/K6sq9iQ4w2SnU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OnvxgjxKvHOLqSfnT3+LWNnahbfmZ1FCBzQnL7P/Zj1qp60s4ZHKPqV9VB74C/UVIgrf/mQ1u2HE
nTaj6wP5RybMtJOYL9J5oYZ9gBpoq2DUTgAFSjIiNmcoV7qw/yrpDuI1LgxYonyVxelJjGSbE25Z
Mrll5wufsGMyp7w4XBT3amK5c/KTWBUCNbOo766gLEqzviFbmUYGYIG44W1KA8kgStjNbUKnGvFZ
vAfmEZPIYIeZA4OjoDumPDJji3vJIPqXCdl9PvhqmyBPZ8vfCbXd40dyibAL65H52sZyzxYU04CU
r9atC5/E21lZQq6cBSeRhJcYGfiupwCe858lQQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 88208)
`protect data_block
EF1HB3xg/IxxVsh8Fu3LfYxlAQ6vD3VBrSvFK3+7Ox5pQuMIS72/x8VXuFd/MgUuFWEQJfvGBf9l
HrtWrL1FjXlaEkVaEJRWZElthnGA3acbx9BvXy1NNj4Vk8p9+tIhtIDu1XJWhPEJILueI6B0L2uk
MiLs/tDUo55htyIAYxLEmAaIeSXijMR+Us8U5NnhwYdVg3yTFQ6hFnndUCeK/+GwwluWUNgForeI
ZLHRdC85gi2PMxxzl/TkrmkL8/h/PPSC9HoBOqNy68TaRiGU4UJ0Q3Pr/0Om07kSvf4zZ26Od38J
RfFWMPUkKMp0MMJf4CM+jzdGMbEhBrW3gLGvr1JWwrgvdDB1Rq6WHH4vxgJfav5YxT9a0R+wMMLB
Z0LUTb5Xo4Vg5+n3YmcRTY6oJ09dMwberaw9TxL5bP5e+FM0n4T9wwLiQrUyfXO0QQ30VkcsBYp2
90lwwBTTk6Svs6yYBO9QX4gXRh8a4i9cC8o9pz6FZ9M/oqs31vmvYfINm47g2px9582rumF2/oJY
Fga8Q8zclWYYuHfB847E/DOBdy9g02W4v7hUURd19P+WaSJdhJ1GS/b7Uxi5R2yQ/Iw5pVvQJgh+
ZjIIHNAEDKFJL0f7m4gvS3dIMxH1lGJNZ8zGR8tuG87uj57Yx54SbISL6qyiY2MqmNkxy5S0yQ6N
LKK4i/4WyXJaDNp4TJO+2Wyx8L0EfMORPvgRHENzAXrzfMML2Cx5E/EdXfmIfxhwlZ/cJGWUuzUH
sOCowZr8kgZ2tN6hqDDXwnyBB0G3L0Z/ofw2DWJ/SixSR/7ZgmdvJjrXQNuJ1U+2FKiHeRNTMwN6
NHmcfRKVTnkLzwRZuL1osPym1lOIO6t4IuUk46Fn27SnD9jbzKGkr8CAXzqwc7TTqw+IX3rFOvow
5+jd13CRpzVzKIy2mxvs666w/sMwsMhROmE56dELaAE4IeYKqTKCNAikgJozdXix/3yKiIwPU61Q
4XmnJKcOzKy8n93PYKdV/TENDu3aSAZfIv64aj8xle3txMsTwic8G/s5Pc3zDW5EGrfp6yq5saZD
hE47JbiMKAsKw+voIiZxzT+/BQywaQMXGwZuLXn+XCWj6dLjDZkGf12nnOlR9qmtu08tE2UO9xV9
LQkKtxPOiajLC6NyP7Lp0Hrr0ikDcowE9wnprRRQQW2lTCcttbsEDZPiz9Xh0slBybL29/kJmdyO
qllFgcIyzkYgDB5Q/OyW2FkAwdpLpJzjnNpqIf6ExzS+/CY6mrUabhsyGO/VGhvWDL6Ueu5+xT48
7L26T7/dr7pHdqs5OwgQa2eRSC3UWAPWpFsGu7N6J9MjLZdeUaWUT2uwYRRNtc5cyWeEhcEqSoVA
/EVyw6PBdJd7GtbTpD6A3V+emVkal6mFqx7iLYCq7Jo/me9RcGhEKc/NgoOnLljmliOaEduymn+Z
FRsubRWB9ki3FTLV+OTEAouaXF9hWgq0ley4O00CCeXuA7odnl/mt0VRXrhMAtQalLpDer8qstzN
CEEg0ZH9Virte7aHkVFbAqPD/8sXCY2rxoGNGkH1YCuY4D/iaVDbrD2zPDmfiDyYic119rNWZ2ZP
szZpbA2hkDwM7QXXlqC50v61ojrP8oN4ejVKqkKO+ccqeriaS0Is7XMUU+Gd+GtUL86208KBpKNK
qtjAFSlJtG62S6jQIj9iAGutDNjbrGmF/afLu8RalD8rrJlMWgyxPrpJOZfFaXyPgpoG+MIBN3tL
EvPgsR7Xlj1uRBvp/I49NyJT9FFX4GsLuzFuxSkn2JGABhdf8g0hq+nQ3yFF1wqdFZj0lvb3sS3r
rEgn+BwnB9RWJqBABdtrxyE7OEdmv03xnmrD4kQiUEJfF3Odmf/nHD3HJ1rfoFdtjGLoGzVfs900
BBpUQeCx0hOLdymDWZyEKhYi/2vQNYtoMgIGGb0CIyzIdbtjfjrik1TWQwvQlbR3qeT3mJQxKIBV
/TKBH334KgICHFKJLkHpI/8efAKwb9ChFQmcNDnuJx3qAIQwSJuLEBMtbeSvPM45DPDYKma1x19D
gS4koCx/GQWj/EzsrMoUur+AwttMxeAOrTvZlOk048l9ii+hcNfkX+GIObXG+hddCSsPgcdHdcMC
DV5RIGaB16IdWayXI0Hpw1Jj1eGHJqFWfD7FFDHtctUB/LxyVsu7v5T+QpidXM3NlMl07W+M+4BZ
qHhrWBP9cMtVTuOycM5JFIvh5IvJCGFP67Z0fB9EpwB/mnlhiovlXfjwHw0HfVpDmIThN/p1vCF+
6M5FPgAgav7W352rLnFBfdDbO2Zvcx9q6NTbLzExItt2YdM3y/wCn2qPPXc3kfjyQcYUL+LKpr3H
/oa4k55Z1J+T36HWXQJYu1xvauNSAxJ+VK8lTZJTbt8GCwhVB3f4HEHlZ19XGOOcQc0+fEJ0JbWu
UVro76yhlLTd5qcWjiGliE4UA9bL9LYnbJUZVIsbg5JaPnAziYCtfeX8KLF5kQAscE96Kj1RH+kJ
u+U7n+kqlV2P+0A+tt0fvvdI50InzrBiSMoVdHSxOnFI0ZiC47CXeO/MCYTQSaBhjZHoG6rFfgyt
vjivau13drhJMtvMgz7V6AnL0kiCGJw9yx1ljC++NGZTWALRCT5UTeeLPD+GegA0YKtVBlRJQH2D
hspH27JO84ZpT3wgkrzHox4zLU/j6YD8nNjon1E8h9t3wpRDPQPbx4N12VA+Kc42UQlH2nNP5b+u
fIFgCYkxi4r2DBl4MklL5RURrkpsvCne40EIIYmzHVArTkvHPS0OJRijr7HRxVoU6XK60Oqo3arv
K1k8Gm5kiZk3uu/YYkTsEMKEicE/jQaKq40NS6w1JAwGFP27f0DVAH4aVgytA3VSwTf3lEZbvr6G
V+T8KmYqHybAGbLnnuQ4PsTFDtRWpu0BraKSl0CMfPig0k4ykU/4w8rlfLgiDMXsBgzrAr3kbpyH
Ng/KEDGU62mS5I0954jdsmkq6Uk6nqYM6rQW5nhPKwZnVJWk+4SDfL70FXexxXwUXvK2N2ts+lt+
0iV+yiqC6/A2R9FwhvSTUpkwKkbELpbtTFbvpGOaKYoJN2/oRsAI6UGDEbuYgonC2FPT+oTRQ0xz
XFraNPmWujJhc+TWBQYcWiyOnxL3RM/wFazpRMP5600OGnOKOGdK4ve5MnDaqu88JwEUvH2nUXAB
xsG4/GlrEgPbiQky9Zo8RU1GKNScYQK1C4SHmjHU7cws5RdBmtespJ0JohnF1psGjpLePK5k3uNK
YwJ3tEvXRm+/Bxrq3Ax/amfQ3REltuKxO1+9M4PzoDL40fhnsTtTItgUeh/EflzOWOnRJLcJjehM
e1KRdy/FeG7P3vrAKV+L1VCn+ZotMWCiyVE5SeanBySudL4gZKQjfh4EMjDHJa/ljDdm1thwMMXD
wjWmwRj2ZX2YT+49ZEWmH6mP9XprYZIq9Nf2pXiH0mRBsLYF8c+Mj9ulfKS8ZzLJmYHkK4scVUkI
he9NYqpJRb7upRezapjl4jMtoJ1xWJwkN9/Vf2KRapjNg0RrvFP9fuXLov94aWYuRrSfhcpXDisL
0VO7tIW0hIxAr4fVmfYKxc/yIoOzF4UpeG5gTg5Q/vSgwWrKl8xooL+t/9doKjq0rWhklzdbgCFw
cQOC80Yj6OLPhNgyEjlaeJ6THbm/A3vxK6uCvQMi/4WlGw6onWa2RNBhUU2HmunTEo9odXUHV3op
6/ohKRghqg3exlJZM0dyXMLns4jlL08toifP3tTflR9n32w1d2NG+dALAGyuvvVyrCtLWSugta3g
3bO/Fka/aCms9korn8XBsv9idIMMOVvHQNbIUPVApsd3PNfWj2mtlpqpVXmFV5koxFatVTdA6zI6
pjJwImsdot2qPbsmupxDxIpdXanZ7m+UkRLxtbicLicKR4nZWX3C8is8SVv1DHJKl2nxQIDWGmrK
bJa3n5fm8u8/tYNlVNr7pwD6TNGVeRQ4TrLtubEYgfp1YwaE0gh5prx05d/YMSeqkEn4LzHzXoTW
VS5qU9k6hcfZwmToB1igqD/pN2aOc3J9ULjDdUM1NKgYFkGBgc4lVkypd5I45wMonEEN2AAP6w/5
hkkHbgKOplvSUC0gkEsR4t29IKfxN7wcGIVqt3HJFENafVOPwjy+a6peawfa/ce6sZ6BymFTDz7g
DNh1tFZz+iNrxhRIoiaam1E+6c44wfhS08152t3d0Fc8y7Jk0OQE7ItRep8cLwzw4mK/788FKlMN
PV8FI7UgLi5t2NnPTaDhCsSBZ3mC8+Fb67+mCxtUGOjn1+WOkwk1+hyp/XcugDfquwZVVAfw0da8
aPqu2TiBZYuoazYXDoBvuh6fyXR+jjUx6jS4B3yEReqnR7vrA1S/nEttwz+E+DGsA3hc67x2DWDX
xVXRaPnPKSFBLy+qJ+dADHdV+IJZHbGi4e5AFVTYB3rwVuCpHslKJsD0O9YyI6SZd9JIrNEVbNdd
FW5l7xfHYk1fCb3JtoTvIO4kFQHnGXTzFbDmbrQcNRqX9SCPCTluyXRmE/r30y0YqPbQfFR3TrGL
Y1cwjMNAlOUOcqAQAuMVBRJJIUFaIM8c10w2SB0nwE1KhYX65bfm2APCv17w7M/cZMGf4XI4o417
4h5XcW2YqsDm0L7vLH9V3fjx16j1Rp7/NsAiMV7m/pMrDRv8dwGHsmmeIdyyc2O6PKCtIT0eW8HP
O0iITgYCoFvCo7Vn+SbAkw869xVYORvwdIXMls0ub9+55wm3RQEySgR4XSOwyneyRr4tkJ37LZ1c
xhUnzk4HuYaW/JT6oesnTdAU37VU0TOIVi+dCNEptcoDAmT7W3YerERL6voOOKJP+BypgR0pkgHB
I8O3YKllmAwDAwyvct/KGS0td8M3hGiBcPd6H4gRoAtwODMY5EMdHR0+utyBajRar6ywUzDbC0VI
MgytOj967/xZS2hCaehdQ7eO3kNzDJ+TxISoVS6MXtLze3c5aplQ92stugndOyEfBXIL6/4KN1Ym
Jbd/LPn/u7GmiXlkKJ4ZjRB6zicHxIgkHHjPpi8iZmDu9VErbXlXa3llsruN9AM2jr8VCIfyliJ9
Df1zpJjJXWX9vx13xB+Jt1roJTFBvQy0R+jR3+Dmc9xV8B7Y+NIQFaQiF3VekeWor/17b2lO2HbZ
ygj1jJ07YAIYu6Ij6EB/6cP2sZlUbdywRwY1l87JCNvg4uSTwt8riBo2xfX2gYvRYG10sCH7UW3X
gs/Jvf5pH1WmnqaUrPY04jw6A85j4G1xYTAp9W6wXysbfex/HONv9VVL1lXKU8RbM5gR0pJ7R0n4
8ehRitNXDL85Hx01Dg40Zy69tV3bmntrhjkX19QVMTHlSY/KvSycK0NzIdFjFModZWVOPRyHfX2X
wHPa17Ecfsp199ZcuR4nUQIh/ubmWs0WG6icGC/lDnTXRoqYNyKneQ0jocKSiMEMw5zRygtH4yeZ
AcNYOuj4PsTNmTAESkRV/gn/nAhHflNuhugNnIswRc1pU74Pl+xlofOmPBhEEELwTILJ0cXLymkX
6wdE1jJvdyNMJXkveWwX62nX6vxixYv9+0wSFQP6JR+YuUlZpch46GShMelKaPV0/TrlCHjA6lMR
ROf016MfIlxU5vznbPXSTCvpyV/1afe5wS8izhwBvavMlpExeOwps8XfRoJU77w+uU1XoJjNMSG6
kbpFA6YVUTJXSkF6Mew2Xt3eJ00DS/fXv3wJEJJnABtcKs5M6xzt0T1AB/vYyJLu24wTc9WhkZE+
JUbrnC5Px0PclIa2f++DNeQN3S/ivByoabGuITx+3IR2YsadClw+jvfpftxdeB9RhLryv4XXg+RS
1eVOufYgDQkvPft3cTzlff0pp91w0tz75zEr5D12XZJX5LBS0G75yQ2mEYj6W+cOGxd5Pwr0D8aW
xwHzB8stgmkwnw895j07YyCTol7MKNQJXhrFp9B7RKr6ihdneMLoBFg9/UMy1TuAuYgo/X6qKRw8
qZBxPKyR6kgmp09BvKVlbJDClmagCy1bJP+BMdHfXvjYw1e4DWLTinI/VnB81KwIW/S8x/aHhQkH
aS93VN/CPdDlQMDZvEOaQlPpy4Mz0kYUpdYpoYc2abF1tHhFDmquWNuLqqpg3W6blF840DThwf7E
XzBsPN0RMSWHDpuYsetzCjnhSsa27GyGSQKc2lUFlPMllf4BBzr97VBD1q2rA0PnVTQiiqgZ4ylu
dcWxGvvAO9DNwGeAlJKfQzvb2Lr7LauXFESSAail37n3u062EZ7OaMId+jdZWklqcoobuqc6T/+9
fD2LirpT57iu6xj2J06UmZrNKnwSgvB8ry548TM3eV+TiBqX4ix4x6kMLIx5ilu97A4XfpcXs+xR
urfZCHoRcFVSZgIXBD8nsaRZyBjO33g8hmzhlQo9FoInhOp/XEpHrej09LNYxBC0MxDsZ03cwow4
MRjwVWTrkqp05aeysC6jIh7s1vh+n7p1H5b8EHAfKhdfeK6QIGcTEaJiPOKek1gvWVIy2a2tignp
c47Q+yACmhsnb+scQ+Kdc+fjo5kFS8aT2Q7OHzdUEiB0iQ1ORoGG6XIjlvkVfniyYqy5QR6UIgcD
NxySIwpiTiLhPsqS/GBIWdGHQlQ/BfoKECZ+V9Ak0E+juReNTRc1hfzjGm1pIcXE7xqoGs2rfY1F
30K8dmcdtuC1XISPt86BbpqH4rhKAxdaWeo3eqHzLHu8zWpd0v3oxopFua7Ob7+6kToty5cTHN08
1NQR58gLGBdq9TdtAopdOj0gfrsnmbY9cjHQXtJIMotIw9Oz+FDcwPAqPWgPMnmt8BBwCq0c/vSG
U2Jm5I/kI4H6zsRr+nz1m/dJMvhZwik5yMSCWBq8Ajn+qDFGCHm4xevhGX0zXjYjmsLmAgLmQohM
ap2+fmGbxomEiX7hqbT+8XTakGCmQmgxKaUc4eHGDYBf0O6u+WWp65eaxIEKHV2ageTDZ6Om+it3
31Y0azxz+bmGopzrqfl5wtl1aHDCBaC5+tHBlR3qDDzAdcrRPiGgAB2AbCgcoCM7NwvhHk2QBqyM
gI35EIc+moFImLgXkEGp+SPiBxvpX9i4Y7txa4/F3IvJ8zCnj0ADeLew+W/Ih/6M3aD2g2XdoNYH
WLFh9C0mulSTbs7QojTwEGYDRyljJuU89Z7kVwiC3SB0bIKtcoQuApLAmvC+MN0F6Ugqc3lwPcwG
/4R0jLbkIwHvNebTJcgzsVUCe6VcSOB/grcvglJTw4JlKqFWWeU/lSfgWMdgJpYM73/g1RwVEM2j
FetYIzbdNHWBRwVfRsn4xPz87wSeuskD72zztqcVKwL+e9wYmblqjs8/nQnqZrRtOKWPHLZ12r4G
EzxH7w8BIeKBGdXp3aQ5tAvkhi4DKqmBWk/5zV8P+VO58Ri8zGLl+v/8VCCidDq4tksYgfKnKT5j
5lMTb8SJjpotkuL++oYE9BrAZdd9SbK+UBNROX7BV0ZbwyhqsjYUnvqU2BIc0vflbpYoXw0lSWrr
ZynQJhndTU/iUscYKyjB4z+r8MoQRZEdCMQlR8pWLtMQKTcSXXjiquzxoqMiQTSWCgwpDPDR0E0G
vFP9ntdigjCP1NrKC3K5WyLBr40gB65IHTATHhrRt0jtVo5NH+xVBODMt3MET4tkQA5odYfWAuZi
pIX0SVhHWDnQNxTzD4vYVushpwVW2pF0Eu2WSr0/P2S5PUvNinJhew6Dor06/MFb59+EQsab75y9
SFz2ZO/Ltry82hRe+Qd4BrQCTU4LVF5kxXjP0b/E9pVobQpNvUPl8bqf3gnzRUa+MZi63wn3eEl3
e0AEiuVzWOFrYbf9CbPaIMT4aZEg5qXpt7WBeoXlijrxZo3mXKplqzIepZRPeRsCPOJ8YMaZXwPO
6kElyTMjaYF/goHlKrDTlmDLKrTvdCfUGYy4DkSRQ1K4IpZv8H0C5X5KTbNMj0LAQhsyeTfTg7Qe
sVtHjRYrTT+QB2hAWer/vT4nwPQHgo2L2RFL8gicKyR7eZvc/tanMMcznlEUWYkfDDu7TGhzeo4T
h6yLSpldNmZOK7q0HW8hmkyJ9yy808wi4lR9K5FTF83TLSNoubwsE/vUczMVlW5psPH/A13e6DqO
vC2PMZ/feLgdxAhCjK0QeKpeVuWCl3xaNkL3FoaxIECHMIJMuxcykzSPyX66QeSqD5ClIu1jgd0J
A93tE0GL7l8eeckaWEdyD9ccCpT1KOvWrwG19jJs49ua97GMCXAQ+SICfDpC9erlKGNXD3NB1E0k
ZyLp9YmNK8PcMnihbtsUxv3Xqj8uKB21VBD8nvJqt1Po0c/rAiHUxOentR1aJvURrYYPEBVfyWuO
hNyBUuV5cU7ge4Dq6JLtEes8zOINTdFgJD4qxaYTQZZyluIJNeqqssIT+UsRQ5MoqFSp2pDUEmOi
VE2Ux5iDehTA+wGvTvOKxgKTywmQJtQozNHTTSaCtpXYHtVZELaVLs8Izmm2gJVfj8TzzADCxkS+
obDMuXJLFOI2Iao+ymocH8031isYBM4gZi+V+Hu8O7dAfPhH1Kx+jGAPiA9+GU8TC3oZilrOXhnm
5eE7p5ETRYB8gnfvrC3krdpnK5Fo1LdU+dmyKcgKKh1vS44efTKUM9pICLugKnY4WDTsuV7bOAdM
DpsTsTGKmKe/J/DKLMgjGAqYMoaC5YTAsn59OTbMlHFaC9jRaFwZij195RSkRGWlMZ+yxJx8JiTc
D2qz/wAF/Eog5lPaE5O0oTuSHO5Ch33ZdAUzQ9DicYmSEoppdfNssG8dnWQ+Ai95CYSflE4z955X
V5eaqTzWmsbr1NyCDN0LaldHjYH2pY332T5u8uyZYcp0Zo48kk1sZLWx4uh/bKDGUsZ8lYiNzTyz
aatPYKxH0v9TB9qThWuSkV+oOwAZ7hTIsw8hKzdgFpnjXogDI00F8C2Qc0xqDe6f9v12xHH14GmN
uqPjm97Rc1yuL1zPFFXC7sOrm+x6Qqer/ytHN+MPh7g8fyH//JG6ARh1DGMo0iCrqZgEkT40ngL9
gZqLsdcaWLuHLoUTdRh0c4i8fXv6G3IDjwvankl0nxMVMSdejKU9Ro+gf6lCNSWfhnXcuxO1B0zt
f2x1vBgOyLZkxFRpI99nhvj97F8PXZczil+PbAyCnzBtQaVACELCoFC6zbR1Vo6G+I/5CzaYtJQA
v0w3n2SwKzAUOy/zm6XHpEYx4i4G1P2M4VnJkVtoyV02jns15S0deuPhYAV9Ux4ikxPYXb2Fit7A
7qm1qVBlngIahnsSOTJxVOSazAIfu6NcdlhYrSqjyV0+Y4oaZSCP+8G29EEbn4153Zg+VWw+8zwr
J3/EAAijH58tvNM8gyrE+HIvPmtJ5U4Y4Rb6iogqatzFUUE9BFjCGolN5WfJv7s5TNPoooLwWyO9
LcpSQSKOZXi2DNHWRTOZmVpue+vRfp9e2TrhEZ5ZkW65MS8GBdGfx9dNFm7mlRxHCJk/F43unjPG
e2pZp7RIChMM1RAvqJyQZrNrfQYSy9rMsogCPBl6yiPEhbfK7sUi1uxxNS71kTj92GQLVIbyG4pN
IIsGXtjRzGDr7e/XE1OtQg9qxxQZIZkIA+ETk8bOQecT4pisKie6OvKDqzaC7iPQCrz0zDHjgwu7
t3KUzZe8aYOm/Vix+1GGE81k8PUgRT6G/UD08VJphp2oO7NOCdW5PTh0vEK6L48FwC+fsQ+lePR9
AyWfGo8RPQCgeK0W+5QV/H2S0mdjVbh+TmXUto887qjfXDf6savg6Rs7TtnzQBesQxqNU6LiZSTY
pxo6Y17WW+VBVF5MF72NXoG65LPd4J0miiJb/l4gDOgvZfW6AJ95njb7+Yi9O+GHVarM+4VoDxgC
hNl5TUbU6ojmaeA2PGwBr/PRxdqFuyOU4uhTCuGFkbkloyDF8XXLmMa3FvI+LwHISv9DcgKlqOSg
Au9TO8Aj382YAAV+9MhdQb2vlqwq07efFZlEJwjKrhD4VoltaCHdw+K8E4MpelznQzeBS23+ZACD
yaPxNqdqblP2juVewbWMNjAw2guPTSp1fKlWDmBx1Nh1kGq366mI+cDUKdecP/WcAPwcrY49vcyZ
OFelo0pr4rl1/7xA93yDneQr+7eM7d0oJdW8pAum8agU0R2IVOE6sjOAIIjC22sA5TilmNaII7aj
GEmch0y8jM99YBUJKQg+sPzrm9de0gbuCutRQPHozh/4NiniO+KmVNQ+UvpSf5QjJI25msXLmG5J
nLRg927Uzn8XkC1ldSExLaWwQCHqHjAbdKqN+qhsCZpBi6Fh8FzRuL5Rm57tfP951+mA/xAo9jIw
3/RyWpBBFmNyvpMwYzAth2i5H5UD2fUhE//XIy8E9rzGPO0UByVPL7OzISkQf+Km7ebcsL1A7ZQ4
EBV7JBA+oxOdyklCPxH2xr4uzsL+6nklgWRgir9OYR2wqf7dIcY0ZU1KVDHteghFLKVxx53F4rG3
eY4UpVrV74E8lz4sEicQRnYhS0klnDbH+XAG71l6DlmqKDQk8oD6Q9cj5DG6jgsm2vp2ggxpj/XM
qVZwDvgBNpFKXLtr23cUtLXoNzmL/N6eXah5yg8pJU7MR1lI29TUMcDpeo8WdjvN9kbLRu2C/GyX
+VA8ZJrkHHAtBplu2O/36OcBVSjUktqb2pzCrThR6aOVjKXI0LB3D5Sqi4oYXumJU+AwWLTV1/g9
7eK4Vxrn5S3s5HmWyw1jrP/Pyl4I4TiLbN4/Elas9W7kf0Dacs9wxFsfXsZ6Eu5ZUTE8CwwOhNFM
4Cf4hq0W/+WtVO9tqiKlVqMyuE8wa0cpN0nSBpo/kaDPaRjNUYcMiUQOhhzVx030yqCOX/JCWybs
vvwUsAQ+SFbGFEzDXKsGPsTnP2GabGh/OjxVqKOhfw5Gn9/1BOux4G4EoQOd9jbMbw+FFl9GkdGa
50IS0zIdtGSNd+EuA2u824fhzC5/1TaZMWjwArW4T3zZrOUZeb5IEPvxMKfRfQSN9nSZuUq1tqUI
j0YQ6QqX6TG2jvM4zKwGralIHOBehBqJiVzhaPkDPh0wKuYlRgzqP/RdGczzty51NZpa0Pm7xH1c
0w0s45zMQehxI42ZCZDxTU6FupjE8mwa+duINDukInE5PXhisoFQGhmBRih6VFj5vM8Vsaf29aVy
i00p0wGMbsvZvwisThC7HS/99G5N1TsyGUzRIBtIoqNiUWMuf9JAlJshrVkB1AUfHEQ0El/IO1YP
yKNICmReCtFNHsQBD9D10jf69M7c4hPxA4iyMysE7fbVilNbBSWuaGPzi4WQhbkZSvpVoqqcQNd4
WS0+YxMP2yfhjhQpqVIbuy1pHwAedv/IwEY7EhgAnHb+BtM8C6HGTRXLIc4Vs3zDfXmuyK2+aCqw
N875ut7zoHPWjq/wkAgK38SYBe+KA9wBGv4LY5dZqADgh8z2GqOQc1kdDFe//OqgC9ESOSlGSlLn
kxnAs4IyagGvWtNjEWagY8KWHvpORwFv9UTafAz5detTCjjRUElnnFH55IniFDPKNU9xoeQ9hyds
R04AZiUxaLsA6ZHPp3Ie2VQkhSNZJhJYeekgZLd/mvF+PrezcPARya3Zdhsr8fRi+nEiI0vNuMBs
xmNYGJTEWluAV9js7qmLhN8J7ZfxN6i2ZP6qY5hd0ruCt0C/hU7eavoZvnbSNW3S7P+nv5P0zE/3
IOz0Ollykk6XbcHXKcpAMCsCoyDZzoFM8Q8bayot5ZjIl02fVefkiVGobbfFYsD/jt5tDlqgUzSR
bE06cm2MS5POWYrxgRtTparaWYDOMKM0LPs3Ew0wsnLoEr27eMFdkx94a7JzFB2WFgWCgt1PSjwm
T4z4hLV/HzDHTa44NLwuugMnffhRUGKYpVvFn3v9ItATG0cvP2oVAxyu9BeJfUMsYo7pTajMHV2t
h7W8Gr0Gcsqv7M9ov1Pt+gtEn8boztPoPTKuZf1VZsVUxYIJ5pY1lcaLttde26HKVIuvbgIIBNGT
+AHtD74+SCCGRDQLzopMBkF+6GhkHE9K3kKdiy34A2fo2LX+P6HmGuVOqQAJFcq76JI2pZgodPq3
4/wZn1TsAkoIgUtPQViLoUeB1KoG4L4Y0VGcdtb4+m9qnKr/06yI1j9/nJOPeNTrbPy41y/BY2Zh
RpQOxNWGsLP89BoP1JaSbiFThL5YTGU1qwp3kvmhrvTpQpS6T4v5VYxQyTGeXSkssbUzDRk/LvBX
II5AwHln1IfV3PNyANIefXvkeZHRrZU/fyN8fziylWY76tuNOaIjFszVaV5vbLi0r2r3GPmgqen2
D3N+/QnRt73FjfDYPiBOOFwy2nyY0viVH6W7CplC2POxLKmslQHLEla7Oq4h3gtpbwUs6Ux3JGXD
gj5y/098mnB3N8iTagG3rmZmlJ+98V3XRPHepyTHHbU76RoklaSoWdfCrw2WOGeC58AHCvsYBrvZ
sRQu9cIpwjIMqpsb6Pp5CeafTL19qf2pTzLDfJ6/wRi+Pvgmq1Atlvd/kOxbFgTsPN4J8wpiHe8E
0yCFYFOzvF+t3HHT1lgPDu7efsZOwyRkTmyaF5OPx6P2eKZI1IwVr5F0nTTj65/EZvV6Edfy9qRo
t1lZr2iPimHoL8pPm5fasvKOgwYHCPi1hZN2OSQksXv6N8rXX3viKBUWR0SLEUtSLB999BJAnKUP
/c98kabR/ECmmwZ0wJ8m/nSFU3b0Tq6PAyBPFEM4ozBomZcOgGLMHgDLcDnQFWI6DNM5ykPWyj0s
38zGNYzUdkUzJx+ivxD4RVg89R6w8wZwFsir9Bl2rBUqYhLWKtMtBWCmRG81+Qg2H81TUwwmY8x7
hYv9GuK8vW9dH7y2Z3ZIf2wF4gq929aKXKEI+NJyAjEwFaAmt8jqWD7d+vns6e8YdoeCeIgvbzU5
c1F8T8P6bcQbogwNVMqsET7+EkdCdwUxUqf8eP8MalOck9deigmQDE5hHySauMLDmZZWrikvan/A
kvV3C8j8I39GWDgxjOIeYTF7/wmU6KxUmJ5xqDJiax4VijaQwfPGNi32LrenfMy45YBtBD21i4c8
q9J6ysi8WctuNCovsmTA4TaXq1f13CSq/+0bed0oSHLN62zC/VQOYy/mIN1m2zxDxCp2tE9GGi/0
5IbYoST9aBZm+QKfBHrZB3enfk5Wb1rSXoRGzQCHwEFYE+1wnm4e5BrhRxIyYYAI3PixE8VkCKa9
5R9viwI6/GOzuPlO4TctxMQMkcHfxNF6Ez1IkoQ11mEBLvw9A6Xt4PX5oNwA8JBVDRLlf3k6f0lp
behJS2dUtP0dz02WehR2Y6I399LdtED/H51sdpLYJzqiXvFXBGs/3glfZB4N65UYdDgmhdVNzGQA
wHC1Y92vyQlLop/gVSVtp4r9h7bzu7PgxeuVVy3Dg8GEcLk62C9H19/WrUxYVROB1i3RK7ZALXGU
38YMFYeLfpUeO/zFWdaeBNPu4IKcvswgzQXjKx//EzUCDWdcEdTgBvdORjInFyIClTmG4H3uUahO
Ma5SOWSG3dR5dApqPK9za6ywRx9ehSS7pBt+NMpaZTiMMJxACUJKRYt/+1Ma9VwqLVsGwk+GOJ0A
l6enupHU4T4iFwQ8r1kcXwIM3kgsN6367hrGaycpO0IT/wKg4dxUOu8ZI+4nDkGX7wB/dTLdlFjx
QKdoSygbEMVXfmwcR6Ue7jAas2AFZo+SOn55RyAr71ezv440FIBOPoRplpBU2kXueojhTTZG2RRT
6mHxApGSjLTjj2Axkygg4q3Oc3Vv0S5dME9kzjDSAORUUDbDaLQYSIWp0l+NvoIBv30Nd4KH6Jil
ng9TOedRwq3DmUnrVGKif8lxlWZIgPM/A+OkdHxG9lreFZfG7CcXfSiUzWLWKGwkPoYKX+9jtLvh
YPH1vyC5+t6GfhLunfKuV223w3MgbSYWaZkxes2kS2NAoaHmRv9RU3nw1IUVAQG1yspUtBuAjR19
hkyq5SEotCtDfx1KO0px1Lyux4+yFdQay0EcKlNLILCjJv8wneVt/quD6MNlQkPGqhNcOGsrWh7x
ScRTE3WjAG7ndje6hteG968n6VeGl/ZKYuSi7lO0WlTBiqjSxr8y06+ssduBRduheReY14sjhOEl
ejvSi/sCrgMXEaEC7wiDO8g4BT0HWhrtQQxtThwx/Og0oPbYR2tRvdmAoKFTKOv+TklLYjf8T4Vp
rTr03qr07QH03nYI2drYtMwBINW8bJ8eJxnhF9G7nuvoSjlqaM9ds28YTvMWSBzzwiiC5JUXHbz3
Yh2ASzChA4tJtz6ZCzz35UzT9D3H4eygf6OUyZHMxf4OeUlbOOaPqgIw0PsSHBZ++inSlMFbeSvg
TYevJKj38NF48Su7PPbMSRsU6DyBbt2DUtJMKo32V/BEcDoGKsyE4EiQoIIcsY2jTch5lenMXDoh
IUj7xsFQzluvmfZmFsAJdDkB/iPoDaz0zBoSClRhunV+HaBc+cfMCx4HenM/WYlRIUbNO/wAbDD9
6NkWAdBtoUUCMeMNmZFDLEZsJ2fAKyESbJU3+sip5YUpv2kl3sJzSmNHFHR8g0nD9gjWbxXibjFm
LslMVIijH4uS/NhcfGU/1WnN4GJuAxsrORW8UKgPlakkGgDWDGnMrkb12Z+zajHTXnNE5WqHpj0j
Jj7pExdUrFdzcQmMQGnaPVLEufJIdg7CUwAWgHLqLsQDOK4CHhtCaUkAu1HeGzdmRZWULAhutYNh
HzUCqWOcTo1FII8+GglSCxh0VOC9XkqyZ0VNO6YSfEsrN78a7n7y4Zd8q+7Vxey3TK9s1uf3s2tS
l9pD40WycWgQpnpHVCmlMb267+49jaije8wtRXdtyVrrVEJ/UNYrE6/kv+FRSfbJmZ18QAPtuKxv
q8cIygiGHkH8lYvYRWu3e6pcFKehX9UfOEjf8NwH1tK27f7iFaQZrB4oz0Eqkjza3F5pIuJzEoaL
i9lrwxDoFP9I7bd1gVliaXR2RGVzJSnDuJco/TMMYFm8o7Bu47rUMu267/ZwqXnEThrOD1AhrI0J
rvrXYPIGowaJg4a6j9gSQPsxLnHgbSM6a2SUrkgrMMmJdxWCRkGHgeGOn+Xkyt5RCd2WUTJ67T9R
bfg0D/K4t041uQ0jyAqQzDMxK2w5yuq1MOg602kWmlxLjQ7qGibLcgC6F90c+VyrE6Pg1rrfAWnX
19mjJD8wTNswdanFYL8JWmR+eGgF8vupqqFyIrB48gDFb8QPBTVdBcdNupLgsBRKl0H4tYE75l6A
l2T6mdBMdzj/FtlRyXOjREitt3X9QsJAh6C66Fe6WsW56ygZxrXLGZ6bnuSUYswOzK9FfPR5i+KL
0ik+pK7M7PR7rGbiGhxWjpnvBefl86ootQfNMqXJajjq89eTSNOg9hrA50MYTBYhX63/QsX5PnDq
1Rkpl2N/kjKU9uTVl5imL3gAsxyUW5LRLhoBkWtFv4/fZiv12JcqrX+wadMy2fPuLaPEJc1KCzX2
JFnVXIxEdh3fdBu4XFseo3tVe6ylJKApBZc27CM0g/A9VDQ8yK6c7x9DYZ3ls5p92/HVujLkI1wj
9aSYytCRkmUJ0ZHf6MFkvQ0rgochYzBGWKIPmSoeAb7pAEeTwIkRfHAtVLZm0sEvEEwhrwBIJxKX
cRMoV+M3Bn0gqGNp0+plhHzaTN4x6MFcSX0IOvBgMsZUTYyZxrcU1uVMsxQ4BYJMx4Ac+Qw5zA9Z
8bPxKJHIgMXNbecSGrC6TJRQnWSIhTMCYeKDBj/R+tJ5govl5vDuOS2qMHEsQ+UUyWlOKrIb/Wfh
CpKyqbnRX05exNBEn6kAgj74tr7/f6ZAz59skt4TvV37Q+n8VEvQ6VOltHPSuV4jhBj9jXGJLqQE
Str7CM8JEqCmyAKUJXOqSJhANOtXINV6uS+xlpay/xCBhZJO933MPKzXPEPc672ZGUpz9gy1uzAI
+InG3TyqStARbuO6Stv/dOfptnVzUqNNI6FKBD85QknWvPxkObGbBTt7u8zojZ22FzveBH/UfRmK
NyUt9MRVYkPIbXy7CVz2p7jkr0gTUfKp2MKjt8WLK5aNiMf0dqMI6KAcCX6NtJNeBy5gmgLl3Sc5
Srv7RDcJV9Mw131FamjwVtaPN+/kyrUgkKZ2Fp7w9uo7nqXqy1fipjPQ+pRYz9zX0HKbQx2H30rS
l2VRqsD/CKN+sUYww7jT37GH+/fyETUmKcGYKs+jPw4B7RzFfLubZvc4FSXiwm0Qi92VqU8VeaA+
OYXx84WTTZ6ObdoS6OgnUeT2V9AtTOsNohxNCJjJT1fB/xkMUi8GcKKc2MoT3gI3bwtpU9Xb5PfD
vAF2PkiV9ZuiKhiVfZxt44af3Fpt4IPVgcMaFgvMEdoY3Oa9OTxyQY60pERmqZAvjkzv5Qu9eaX/
uqIgcGG4Ik7sks34KltR4iYFEjv/0MjvD9mhpHAlJSXieAPCp6RzvcW5aGETLONaeaBklroxjpBl
xIU4mcj5jc7TSYAHqPL1Wa2y60HuBwMFosjpJkYeJleGDtea7H1hxYjIFu6tBlPGR5uNZgx+6MYK
6M9wN2IuwzezX39AM0KyAVM9Y0NQ8zXX8WvLTDjD2YOwBaunUBi38jafv8cxxV1fyol4ekdlmwma
J17WALRTklYFdVNALXx9x4TSf0KULFdgkQboAdH8U6K9cQCmCGWQuDwsU5izdsk9cUIObs2gZIPg
Q86pYMAI8qYm7ut50DFBdca7f0XsFFJpxVrNIdWqV1PwUPRUIaB0XNh/UfOq3ZWna1sZp6qZbQ4B
RfhVc3qwbeY0J1l/G095rqYObkGh8sw1RAb1gmVQujqBJg4XmF6aGDhLz8hKg9We6QTjg0yEhVWh
i6ijBIbGUc+TGbM8++m47GdlPExEWbnbS1OBBE5EE/OeLA63Ee+K2nLs+YO3KRJXkTPb0pu4cjsg
Bo3wxfPZUjVv85KkrzEYtMQYk1FRpTa44e/wA0HbZgvEGvadY8XkZtGb6R6LcN6+zYabLDBhcFad
98HDLIoyu8zi4cdnnCERGTucxU7zAqTaC/A0MttMVpnAbXU3GOl3gXZhfdSse6ZStK0ZlyGAQdBI
n4SJGLPuWJoep8oG7VuqpHDP6Ji2+wQraErlbvbaQqRSMfsX+ZJsz7X4ZuzfugIaYX/U/JoNAArx
aOY8vgRsQw1opEiIDpcFA3QuP0pqA9KpfLTbKuQlWo/XxCrrTrlO2+tggrwVLJLOvJ3XYD1AKxv8
8IxwzEOA6B7MFNIqZRIDE6RDBiyxLRKgEYdTMqLDpdn7wT2OB5RhV0yxqJgK86eEvgyJC87PjcRu
qjbjRH6MBnS5G31/KcREev3nx1yjOgXEyjRAG0jkBDzelLgQxdF80ObWB7tzHQ4trbFVdq/d0FpQ
IX9jCrFgk9OddlnRdOGQmZ0FFN+BcjrwnQzrkTiN6GZKz+GThqQFvhUVqbQu6Vp+KyrOO/w5TKK8
inIz/RcuO+Q3HcpPNx5rtztnX7o1T+iXW8iKBOva56yQvvqS/fP26mfj3zewmgxtZ1shPFXRdg+n
asL8qeZBjiJHyeQTkW59hAuBpw0UbTr6aik3ZCBhziXCUsTaK6g5HUSMNiso79SkRjv8DpwbK8u2
S+vQTo0Wey2vSr43Qg1ecKsF8zBWZr5C5q61g38Cc0INZv4fnVmHBEBTwxgWU+I3I/Air3BQfoH8
KUU3GlaNFN6Mo1b87ssARIoFfrDS5cjBkpvwg+dWInr+k2QpEw9jtIKkEhoo6RwyrUumDILz/gzk
LLvHF1/vSjMZUrtl2WB9LrhjGRpB9krrKSasZkR0MxFzbKhaWwA/XTGHZT7PalfFC2cjeUpmG3r5
PZmvjmS0JXPbkGnoDajnJZg9M+sDVIwkOaFsxgC+ABMrcIrdtajjwmrubWCoSs8ODZ2kJ4/4KSIK
ENI0Y+hqFjBu7jRqsK/DeXCBl6t30WbG4vpBNm+2RNl2Vi1SggjRNohF9Om3hwE8yrjv1Wan7ydC
FRWDr63NuRGGc4tjGgXpbYyjkkSih0Uw0+coReWpdyK8cNpLUN7OOBOGshv7xYC9c/uhm8yIDVU6
OCwXiW4uWK+wB1qKFQmh/5iTQsy15ilNS1zfCo2YdIRTgIyRjFGUjLg3xfCToUugqnw1hcSDWOJm
H2NMO0BBtUG77hB1YLqNFL31sdwd/A3yKHFDzOmQVkbTMJ27tvHXz9Ro/dNSxfSll5WXqoE39TGD
3K4VBPAi3fLtP7g3IAuzv+pCn9DLcfNwLYrAfvqlvINo0jvzvC2WgtcIVb2r/5Ho4dnM9O+LFOu4
obQRywfl1whT3pxjf/NrjZqtk3IGZMU0hWEY5OAErZHYPd9Ynhw1RQiIPOix3+rp0ni+53SMz55F
G8veG+EQ+hFagMdUzpvK6P5zR2illEKZZKW99d6vNWgEpdTrB4KGX5PfreapTo1X13iBWqavNtJp
9lbTx2cMrb/4PLQVak2QbWTkQZiOxRFFkzhIbSNUqQzzwivYP814hT7QemIoJP0FCxfNtKjZ41rw
PcPV1+axOPgqatIUNxQY76ghFDsfFJngd1CL4qKet34c8QKLirheQ0ISJkC8OeDKaRDX4vtc5Ovz
UE0gDZ8C90Zr2fDkZih3DPZwxwb60PV3trzokwWxHeZu4CLT+b1pyo+JZcHNRjSZBeaySOIFQCob
bBlF1Fkffc4xgN260RYwBuZM8l3jrnMPSnW03lYlRFvcOyaF3owByjsmIzl7bLrGyTY4i3tUv+V1
hxTwQ+BHOM1g6MmUVjo5wXKPjIOIvKdv/5VyVNf9XuQMEk8lsPHr4ekCJyeKpHBan3mHVQZ34xal
qbU86cpbUbAm73isyOxv2ISbGcvoWAahusjRN+Yro3q7ZQp/DsYWzmgc5ud3NuBGnEUJBzJck9Ya
nhjeoT3Q88TjMj73CzM4V0J/j6plKTjNodDW0EDRb9zvQrxSPrM1QKIqwN7OqjoqNQpHpG7yf7cr
fcys0mO9COLWe11Dd+uHdPHYapp5mljiArF4LzaDx4qvyKfTAOrG8n0SPp2k2gCNPwuHg/RMf0PG
L9zJ0UfXw9Afs/Usm1+G1Z/70kjORFZBpKl0yiXkwpa1BvzC/NrZLOI8rRFCoKOpdcHo3LXel518
3sep2jnDVbrhUxTUxjH1e8mBuWz2Puysky5BB97CPIRBJlIIXDrW7joqBHGPyCMLPzqglKOI6tgc
9eSYwHUrUF+VpvEgcXF+U9ipLPdZZ24z21/8sypGlp4oAo7gdPq+YRny/p7cmfW9wBLRCKKgekp2
Op1YnRFPOFEi+At0Qu34SsBlx1e4CcKwo2X7wjCjQsOWvdwv5Z0MnXMFOofaF+hVqP2OMEVqSXk/
ImSGxE4IthHhdeWznhMru8r5AnncvYSp13YCp2D1ew5W8vQ0WFs/3En18u7Zt5kjqFA5kW6U8zry
jyJTZO5hNFUPGBvfPMRnpfV9pYif74jRtvRuQYr4AlLKnnz2XzV0GTHcxMigoH80CVjHqhntpxNZ
5PQ/Atkbu6eJeY6YfjxsV4YIqgeZRZb3wx9FduztSNME+E2biHEMhMTaeg16s4ir4CmiXEVe7m5C
qaoV/arD6SCNJvbqjPjjpy1o/xO63+lvlcMy1ulyPyTcKS+GvL9uW2qKb4t88U4jVaN4kmEnMyoQ
qDJ0QRY95mUI1xxUkmcLKbZr9PfK3xV4xjSRNdcwAIqdES8C61CRB17CYQ8NvonxvD6lVdGfdOrW
yjqyKXZfiXb1hmBMqC54zjXPbhf1FW3yYLAC9vJqJm2yBwIIoqb7tHKTkYb/G3h1jxBiHseIItaI
DFSKh1OQb/0vd2z7plDJ7C2j9xMPBlMQyP5olftmx+4dN33+vH+p4dmxYiLIiUB8j4Co9+eprmBU
ARXmzjS9u7kE5yilpppSJyYB4+nZNkp/Ab2wAMSEOGGsBzeXpw4iZ4cJ8n07mr6SArSsZA+q7Pw3
PErt1jgsPSDfY4A+ictkz0NH75cQcbRgnvyIrfIxfaQAf6iqniEif7ECy/Qq2EBVRCW61dPe//C0
fExwytOLsjUN5MEDVhHesyT/tP4ElD3ciNsQMl9oZcn21TZ32jSSN1pODMrsWnV3/fmGScK33dmt
Zkc8CVUmFrcC6KQaTacdW5pdGCiEHi2saimNlcC/trH/qF1UANBgE3qywypNVd85ASZ5W61f2mSH
F7+qWkRqtYMOnpwz96Cg2IeT+7SCZtjwL1+aJIAllRrkZLOLfFqLyppyv7HnFl8HSTJNULPGOZyg
mqbRwPdwcJZQgfkvDVRGXbmgRG7hgu4FjPCcpEk3bReeoRSgoONDA+luVXTfF5STR30OIZsOcAnH
JEPUH2a/Bs+qjT8/Qfv22PUiWjKNRZ5eSu0C30dy+7WvYHgI/4a+4e+ZXt6DIP812SNse38C+BOr
8F6zqPGq5P+i+kRx2rR8YLRNqEfAFF+S0Jij5PeWy44mkzjGFHnT2NLGAKcUvbLNi25OZlrkvJD3
kAuOT6JD17vwV0cagZL0DseOFRj6dHgx0Btg/GyK7PTPhruo/TV5ZMTBAAWzoO57e/4bVtbLKm4s
MlDNwXbdgzlbo3LhqT/Ts+cpQbSfDRGCDVl5MypKITdAr2eDCgPAQBx/gcbC25kyJPJ6WKhqU0/3
AiDESwoaBYlGgCxPYVlAN2hanG1pBeNc0yMPd9KVKc2MLI5VyTG7wPW6MW0J/pGWTMr8ngfv0UZy
CkCpEzaW80+iZSw0lFt8IRG2IKjwHY4PQFHnLu73+FSB4QYOhZk+ZHUUcKduAWwLQ47MjUmBeZy+
SAUA0NTI7+dzyhabXlHKMyvERWmLYIxF6B840ENFuvg7qeXTT7vlC0GCCyxV7TB+o5Kj+LHJcF5k
R85FJNF9PXMimXlsAO3xnAcv2TU4ZlDIIEA7EiUyb7xpMZtqeT1q+pBdr4CeB2T/t3JaeJ4RmNVX
+s1bhRRA6Qa39daaJO/q4b5FYHcf3oPz7gICHz21gFJzvepC7babFtg8EBGDnvegVn2JayHO+Ey2
nqEPzCEfghZwdYc2Z96tN75A4cRVU4cwiD2ECYIjbqefXwHaQOtWUvuKmw69g3LdJyxw0rbu7elz
x1bro7Qp8Vy9IdH2+s+WCW5KzTmCTO3Rl9ZzylB1YNtNJ6KrByt3dZuf9sB+KR9pLhEivlBAFFhT
6J4nABEoLSr7rzsiRKkhGmjTYBTyCGy1sdvlpCBaLMUyCHXRrS0ZA+sFRVMLBHrV4R1OsVny5jsX
nSnqiTaGGkk4MinLhW1TQaAAE4YJLwGf6WQ5ZoD+XrVirVKY6d8mD6VeEsvVu2j3nVSOBxlwV0Ig
2ZfWCIR9Or7NVbTpaCR+Gj2/8P9kpX48FcYNeYW0EvlV2v6x+AwkpRUk+l1cEGqiyjIcswkdi2pI
n6b4TMMXmxKrupTyfCwaGFX/JaCFVN5ZhIdsitkMcKU1stTrHvVRHE/C1ZWnwE1Amdw1r88aUMiq
eW7whKjQfVQySERyzVitwLavs5sDE1rla44XwXIEqrRwyISl5NHhwi3GnJcmWKWyjNFa9pMB4vxk
TQn40h5VADXTPtNvj/RwNOs7xjEgGpr5RuxovAlO/+zu+eQWscE/Yua83Byo+RTz08ObqRMmn720
NzW2v/LBMmu/cOlCaYSwSBk5NEwU8Io1+fHBzppp1wFVu958dW862g38u1oH1pd/t/HuzLJvRHpF
U2fDbmECZw+V7GPHQfltSPfMTt3byk0FPgS9BXmXORH2OvwqJXpLWGv/J0zCE1BmPyPpunAkwuHL
LOoa9/vA/Tq36YXSCe+Gh+rLCU8mVCQwguXvvZQa3DMKLYguHGJKhRBagQmsBqSS2pzGO+ftA80S
DYHUB76aVK9fH5ULPNEvfpKJ6NWdtliWMEwEoUfOqTjKBrrVtttP7feB9/+LsYlbbN4iccXA4GKg
Wmh9Tk0SFXD64m3LPx+vUwK43A8DrEvM26IBUF9lPWURplJdby7Re5t8o+GB4ecdOT66xAW0kLcy
bbPMT5HpH7EeTRTHEdZzR7EN4TlxIq/w1k44RsNwJs8sC6BrKIBqnpq+r4MU7sEzfxslcKnUZ9GN
J4xd6ApxZ0naFLmgro6+DTOUjz8Q+dB73hvI1T0iSRotako/JQOODfzBZwZSPso5+shGcC2QACgz
ZpPe2EBVE4gaYSyfUW5tnktOpb6QDwq3OxbJEefMoHhoLwdZ2BXN9y4HB0ITsLi3tPRB5CvhmSjU
W5i6t7EEcdHTGgKodM3fXxn0C0OHPPZ86mBpESi9xUAvCLFvyDjPY6143bhr4pBM8z6blCv8KsUl
vuX1emd9WGIqSukfkKnTrfj35k6KK9dVqxIzdQiPI6iNF/O67fAg963bwTWaxmJy+0B1lO1//1+V
6mPPatVTyyGBsx5bQqgY+kjgYCdopGxmogEY6DZjQWBQ4HZttn0bIoipixieInzvRHbSf3HnSFcB
wGQ95p5ujUcHtvE6VJ1ql7mJ6eazn2W6cHXEjeC2DI6R2HvWTEFmliDRSCVhArCyEJtqLfxXi7v9
bcIqF07j45PcjdfrfTbwpsvFxNQV0QMxtb63XxE7o1RtlgofEog/eGvBxh6Ph5zX0FB8GldBAUr8
jBDeaO1tkECjPbt4WTI4zJJrBJotx3Fi8E2Zqv6l99H8C4T3up8jJusZCkFx0w33PQ2uIuHCkqtZ
2W7ogHIdAuc4qj9WJZkxtLtLDdvCcKnPb0sf0VHqhbCoDwVNZ6BijCMkla/yve+DUnlQiKWSheND
I4/0PMMFBIegQNebo9gdEKBiMtUjhVMdeLFHIlw5BB4BtFXoz8vwNPFhW8Kedltrc2SzEAp5qghy
iXgy5BXPkALpX5FAz4yAJoLk543yCnMsqLxlw8Ppu+gmoI6WC+jzXX1HObx/LDJ2Tbr7kRxV7Fts
GKgeh58H59huSM3pGSPicI47PyiJLptD1MHGoXaTIOpBGu5IGzP8Qp2sz4g1oV4nEE7hD1wMtYem
LUriiIjmX5PPoExhv7Wh8VbK8jCA2/48wjfSDo9Y1JBrGTK1H0DEaoR+7LTxlO362psLJjIS8tyL
L/P/NeJQtWg405UA30vsf4HtwM7/NzgUQVGIGQlqy7nhgSQS5MyRYwZfjPc7Gkix056Z4wcTgasc
KcOp7JGzIQGeMQI1oBRlIy2v297rXX4Q66z69dPTmGwG+WZVQ/sB6+W5gSMjROLE7TRzJmqe8AKp
GVbSGyukwkwkT71rXFB3y5YN3FlgZzphaNZ03MVi0LZIJ9T84Jgqm/b6h4PuG3RAfsC4H36rBM/B
ngluMrW+L/KYrkaIreC4+XburMQqAE1WI/X2l1Q8k5dDsK8BxeR/IUFJuzfQr6IjUDCDGm3rhydI
gYWwxKW6/CBQE8b3fTbdmcXmpLbXM8yt4gEXnhQHRZ2ekDBV4pK9BGZ8q1DTqTRhKpeatAalZ57f
8WIwN2tCZIkUUd/Q18XtUmdQNlOjWuYrsyZFWJsG0/DrUHZOrLUjSIKz8puWzL1XTlYKdukP8bts
1Xrk1g9YoV7T0T65rlUiiuNvU7T6GPYq18gSi52Y8zwZb/WzVo6fuQA5zdz83YWWVjz3RtpV1Z0p
mLXzjliIXNj9Ve0fkhwwaj/auVw6cSwABYbIF7tV1EM7X5TSivCKVrmfnsBQmVoSFPTM5/FWx1dD
HWx74k1HteVooZWz2YXiaKBBLK0baRajwhZcLSkADbDksMrhOPU+B2mJYaH/xHr6TnC1hpaY/jmE
c2SplErhaFyH70vOne9azqi756eZQlicKrZjGPMCNOpVRqK3Anm0iOQPjx+T+j+8MRAWoc7hB5FT
je8SHnLgo1vHuFMEFMzNct0PU9Udpcd9B0YQwliqqbqEUSQwl3WzsLe5Ghs4RajWDYeUtUbc6AX3
Z0LVNjeRY0Rf+Lmy+gq6Vz4ldxHHmfZg2zsOhrW5jzbuvphRg8CN3KSDCNL2EBACwnBDo6mErSCg
deMj79JTSMQjWxRDukz68cuyowICawO2FjAJisEXYL9g5luDVdJbf8olPYYFfF4EW+d804L64v/L
YsPu0mOBQfpBTMiq21fIDcZd4hN4qXdSa1MBETU2jGjmZkcmhy/MU4cbmxBqGeVfsScMakmG2g7v
f/IvmsYPh29qmDI8wTM+mxP1ULuKjxRyIthM8R0V1NbESF6ZZdvF/KEG10AoDYU6wiV75zNydwDm
WT8CA703NCyS0KSk0JUqbhO2X0zt+gSSN7HsfzlqapLIvPbgokGnPEr0TPMdSGEXQ+INFM8HIbxI
+vXO8i791b96E9ABlaKNBJu6M9Bi92aT1BmLirve6MGG1rleCm2+dm1onQWG8XlYZ/7f2S8qSIgv
DNrnmnKoAeOSx9zNLc8SW0GWoPkh3b7bKUkxCWN5omCgDeLAHf/y8f/4vnQOzVk3qiQv+OBitJjx
hb8WYw3pG6OjIGlIp2Iak9MDTpr3NzssaWkBShf0V/pvj1n3XCKqsAwyep0k9vaValDwOJ7jBh9F
hQXbBokFr7eWdw7KBFq+dvBNSXZdRfAEIujT+oNz6VLHHeBEJBoIL8UyW3R0foYcf6mkLAmvZXvm
gHYZWsAHOaGAH057arH6dzCpdbSsUo+ujEM8AmVxq0/632ZohoroZ+CI5cTokbXb+HSdWXwcB1v1
UA0ZFUt5dsSj1BFcwbnGWuU1M+fRo89LLs6gvX3W/eM0jzX9bmT2JVVabTePPFZCkBdXhxoZYP5Z
4fdf2XsdMqs1uU1QCaMP1iRyKKE3uIpJ/4RghqGDl8KtMPzGB635AeH8H93c1Xsc6K/uS08dF+ZY
boUUkpB0iNrXPoOIvchkQKMdVqqDYBd1D0AuNo9L14fm9q5jpupWAvSXQx8gBEifXCnF7Ws26cNn
4l9PUc2TaqbglC0Q6I9uYNOL5ApVJBPkXAMIQhd8dWe+h8lDva5PvCMvsVNCeky1mTXA2+XSWzwR
hAMiJogXtwnI/2MlI2kbYPjjbAAvEKJZ5XciLXPj+B5srKE2nJc3oBg3XRDR1w8MSSWNV6DLwe+4
VThPhMuK9K4zJ4BJ4Zgr+dkvGXwg5V7KaNYIZrDRAB/2ryZFraBvyv/H2ViUZSLDkYhvcUruRxME
79UFEiVc+ABMHPkzFNjH7w75Qm3ZLu4tmxDZBkOrgX9jkOGsiU6vqj4vFbpvATnLDMIH1nZkZ0Jd
1434m7rb3vLzR3ZCEFGrVN9kYEJP3bAHs6iEfY5LuMcH4roYqDzkmf8YjDy7Kaa7GgVFOsQzmS8X
lQKZ8plrGVqi3CDpwncIzC3iBDxS2vEjnVFKBSVCiXlYYLbQI4UgGV+PaLOV8rpSdh5JScDfcphp
m9pptciKcxgWDJ94Nr5xtIkctJ8iwld3V4vPSj1Ldrt/WMD1XC6r9O6Er8wr7CcLUhUxTJs+c5BV
0cQyd7l9FpRITuMJ5afZp2c9P5BtYVzUfJYOvn1PpG/G+TAAPNtgFQPzrujad4dWoTbbQ58JWbJD
JwVMAlAaTrks2E1NI73LngqRdBe4juLydWmC5jqxxzxGZh26FFKUJmL7m4nL2H5iixlgXa3jChRP
LeVm+NXTpChtCooLQoblA88RxAZQ85THkw/qanESpcl/jxWC8FsBYsgPLDDcooya/DqkimcgPxMK
vP8GMt3QC7978i8ATHF26yCGlxOI2KBZd+PZm20IhoW1fPsOMT16JxrXd1wN8Yb08V/NofZVUwq2
m7Jen5yZu0H7ms4BaQiJ5/PRZQzDIUey75wVLGePi1hYmSzW6AJKDU0ayuSq00AF/Line2KonWkL
4l50+7sJfIFwCMBA6gmOvjJbdd2RgNQUYTi3ow4jgz86qoH95tVmG1WCVksjKIOl262OKGOfTUfx
n8H6eYoaFbqWyrDFWAsWTKloPi2k7G4NuXsSInd35J5Dk29kbNYrqPEnI6Aof0+bcZqpqaOLlDDU
gQQG7Z/H8OspSE9Eqzjsno+jJ4Ur4rFP5Kjo6C9tKEaFgkKNYofx3e4LuoNpblDhB7pvdi1MWIYx
pKX7lI6yf1pn3B3EFwjZT90H4QRAr9uudo3oBVKty/KJC44xALYTtLEorpLjjvpiYkaRTXqHW0h3
fsU1vrt7pBlsOJbtVWgX2gzPLNMKNurw48FKRyivCtUcT+0tbxwbT5t27AYYGu7dDZQxLfenBtmQ
UlpuNf9s6zHq/+uttf1dpLSsmIF/YCh8H9y+oLwh+pftbzv3HWBdzZQYLuyv/wrwTdWxV/gLFEI8
zwkQt0vgh3nZ1vbzuIf1PUPnTyBkDJEcDpUEGzA4UhuoE/73FTl8Kv/I/QyxcGU+tzjhYoTqDw/b
ziNG4NpahoIAKbCIILDVhXIoNvxh4if8VefZDV+6zbkaR0K4Q2AAQza4ZTsumAa5i/ej9nVv4mxk
HK/aWKs2MW+kgePhk35vJz+O9hLOSKLYaZfvOlMBmim4O423PuvB096BnL9MucOQeQ3NJWgJVpZr
Mt3EGBQtsZ5ktSBbw4yxyzNmyn/1XO1lbLweL/RevBcgLEWfCpylvBfwDdMYDo5ojmlYjcMB7M4B
AITFS37Wmf9rN42pvluirWKkUqofQBljkdC0WN+sYh7OGdIrfQKEtK2xJscwjNUpwwkBc8l84PRo
4Jar4Y4+q47gDZgCN7FNmpRUZViBAVcrXOLBrRbeII4hYpdPnAftOdyfDOt+3p6uNbFQfa6NuP4G
YxrboMCkIrevWhvXCu/cnrMV+CP5cYTcr1ScbMw8qVw8AASt3/9mVXZQV56n1ytY6PSIwGlLh4hg
WLjHzPzRH6Kqs5EjOR/msn5IWbZvBlRrsOo5yZeAitffUs+CarUanlzEFcgs5RLsTHgGWGtIrW1y
q3fBpM98w1X/N8mrxm72oSHwErJoFVZ+7k0jugNJt6SH5v5PZUWOkTuJu7tAgp43Ktivm0TbUvWV
HqTMkhsymupImnH9C/xbPixKCRBzT6zyGLujjwpKRfS7zYm1rqZv/9k9CAMLhcYUdb4FfwGbpHYZ
edfXTFRPG1rPuLrteaYDBLR5pIY7w9poqpjlttDMb0Pr1byIAcijERAjPF2LXrGvBaVyv4Zj5vcB
q/LrPmve4ajn0jKdysxByy0z3i34BV/WXAr5P/9c+J+EdyZVKDTdMDU3t6GEOFRRj7rqw05r/hED
94IH7b6a+IPAlqQV24TyDGxOLGNdIB+j683fREkr6g9Gl+i8w54L1ZiJeMbhVOJAxULv3xDVunMu
VX3pRWdG7dA0hDa6M0svVFPsGSbjzVFcv0Sz1fzMWo25g0EcK7Dv9Z35IGE+lvg2KqXfot1n8CVq
fYl4pVy0YW759p+Ff5SfKogakJGiqqdvLOWeZVmkTkRYx+S8Ft40E3Kd4bRgpG0z407FK2UVyPLD
8Ou1hvrGaxGV5qVkG+YEfJU/+GASWDhT/nT76rYfyXAF4qyh/B6ZoPCSqF52nAJVzTEB4fV91nwB
SSr7DqPV3a6F1XEfFxIa+OpX1Bz3w+bGzu9IQ0bK4E5iqLQ8Xv86IRKTuKj7IuPi7UGtx/tU79Xy
zj3NJSCsSvIuNo8By6QoA2zcGdmQvMmKuOYMkbFl2hP7yppaIhJBdTmgmv4YwU2cVtJ18SeeZrM5
SknPKgh4r9DlqvSKipmklZy/Ky9oQ34Z+arV23SsdUEhqdSo/bNN+MiFOsIzMlGRWvSW0xqFSe1I
2AJliMF6+BgubLNc0EjYyJUdaLJrO/WdVbwKUJb8aoO8QXeerKGphsSMteh9t7GAXHP0rdZsE81O
ijrMX7WcO4y9jKNepgFBABNjC0UFNr8Tl2Js68q2Xr+pRZedbggF3Y0/LcmAanD5vr9tW7dM1/mN
Cgys6T05BvS2B4oSezwEpDWisz9SCpRxKb+/oni5LwQqhRNHJHZiCHBqrB4CcqWsPJ5rFY3dmmo2
L/wEs37Kk0mp+7zvV/h04XRG891ncbAQNautMA982wuI/0211Oc4x2OAiPrFExgGOAPWT3n6A9xf
lbP+WCTWsaFiQpdFdUREPqjcmWTjQV5k5NP1NcUbLGc4Sa4lNqsZ7jVV6e3UcRygoBMPr/51kvgo
H8HkiBgRuALvV23lZApJFk0zmBo1qDie8Q+67/BNDWcwFpS0IVGPdvErXxGVUEx0tLk2eLnxZ+OX
LHLuW8sZLmDSdx1T2hRmi1zn6JfkSICcRU0j3QKhWuEbS4QPLTCJ5jc4Olwnze4qfBHiBARCLt72
GXOA1cORQUskgBrYtHu9WSN0JwcJoZ4KEwRkpti0ot3A0+ghtm3mIB2+mCMP7gFQnwiiM8/qKR0Z
N3VSapvG2eFaLNw+vMM0G47EnV1KI3HZbdRQKlkxAmO/UaFzGlDCG6JgMZfZlukC2yf+7MQkktSG
pSdtzE7WmdB5Gm1R3Dsld7ze266UDeS1At0/PNeHoZzeHalmFsyJPkCtNxZtOaNFIPW/P7Qyp/Wv
wb3/E0BPkwn+jA6vOJEpfJlQgFhKKoi4R56kqKtHCwOazdFbqozM8Svek5Om0YY5YmwXTaiCdfIW
5DKpNo+JwjpEbxrQQu/TvZie4P4ssnmqLd02Yv16dqaWWES+GQVb5TcTsuEoQ0jgMrSWnECsBm0q
8VBPjB3ziXtbtfcT8KDXlFYl1BxhJ5yWy02EMho/D+luOntb7RQABAAwPEuxTDt8gLpB8ffWPL/o
g/QHfpGzC+F5VPF4lN6gJhU72ETEFk6cwC5T25kj5L8roHstMWLf+EE2dOR0yxpyu6luMO48o/B5
zxEPBpSdCSneiAtRwOjKRiCr6gKnLUnGSRU/ztd0mj7IaY13R6rmbcUCCEh/oJecS7EPjVwzN6xE
0MJcN+Bi1sPLeICvMNdVR/RYYTDtqsmdxSvcws0mUM11dYsIvk+Plnk1GGWRbWBlxFzfJsfvdfnd
UNYLpQaoPzhcqYimCL3m3cnrT6nk7GabQ51mn9RI5DCe+fyk7eux6ZCI3/0fvH9UE1MP13c6r7cA
SJCCS/46KUK0Pwu+DJA5sQm5fG1H9t6CsuA40u9HeTQSTN25jCnVMxchU8bez0cJF6forOPhW5Ra
TT7vfNsOawZpNsWNjV5X069VJZ9npqNmvig7Fb6FJ1LMgaKrTzGepgOpECdTrXweh+UTrBGhAlxR
I8J/T8bQ074hAjWj3FUO4ITyLZ7heXieInzOZYZ4ti6OciLr3NJDlYVzyVIdCwYE9UFCQTu5GSFY
7wGIcGx7ApjAcH+C/QVA1YYNKfxnWzzzm0j/l081aj780eW6vN8sy+esEqHh02aACJirBrl4GBm8
uMbcXY5qH3O0+63gdZ+iNvRXkM+qPrEd4I/iV+Xw7ev3/RAFxMIkRT5FhMPXTrCHvTMLrpWOel6p
NU4XCS3NhRibxxepaFjCKBvniUJ+s8i8ggcqep5cuP/Iw3HkgYVCCrwLP6wnClGo0Xt7LLZEVymM
kW3yR9764dg/gGCJpXTH3dVtA5x9eXff55lE/7sURgIazzVTfyoOytKxYySlxHLOoTrbtLKaJ4sJ
X5DIjhs9XMVo8YSF72p3DjOhip2Cx7pmRIslW8UZ3w7DWMChaOLn/fehT9kVJN/St/6prhumo4dz
MZq+YMjWzC2dntuwvsAUc6uR6Ahyt25i+73nCUIHk7u5S4p7UUdkZBZRzQQ4/FXagyGhUm1edVMk
fWF9bdHodoYNArbwTCAY2fa/iohjOpWfz97kIWH6f30ZAt0jRNRpkHAVvXnoCj3yRiyCLA+xxZqQ
6bdS6ReUrdtGvZtagi/KjCyNRD2lcSnmV9bV1vc1oSd/6JWvTupMK35j1a4+iloxcE7Kv16ZA7Ku
Qdp5pb1fei0PSODdvk8Ekwmwq2wMFvpPRNPBu1H5QjcLiJ1JoVSHWVsu16J5+WKX/8VwWE4Tn8xH
bQE0KvlzXPKHKb6kZ7+nFv7UWlrKx+S8VDpfgxKQOm8x1v0Z1NTilHOCvUqcv1qZvAsSFzFrrU1G
E0QZnsc+8JNvBsOQNPTI8fJsR2BVN6ae6GZBTs8oA0vuHPlzDg8SvRew+hAogVWqngHgeYZYaFfR
fi5AvqsTX8voq918obdheFWi/TsJBorZkl8aRCcuRdEPNU8lCKf9jRBYynXnn3ayUmEFt8shGOq5
EFErFddR/mH0eCyWZ2+FqUnNCXl7aJP6cN0hTwAYqGGxEq9GtP4IdhHuNPxLUp/F79z3rog8dQ8u
oxm/WbtF8I4tscqhAgbSyrIQnrD6ZJh6F0ZWdWUre9AOjxFq14o3IxUDKjn0Jbps3js1+Ts5Vxnr
3H9QogC01MVmYlkMV1+eCTsUCSZ+cP5PF9gQcFlPmAQB9+LnTgRdsfzwOkEzeRCyk9Wh/ly0LgYJ
r2PrqlBNLQum4j/HlP+8xfsjR3rqEH4aT3MeZMQ4PzD66IzSM1XFZh66GRdzR0CayHfdcC63bKQ2
kFyk3Ku2NzBvg9pinL8nU2Sf4YBVYO72nzwV+U1tImRLVKZIwgSRFhshKymbnC5tVbJxCO/qBVVV
211vV/NO7g4arK6mz3k8ZiqSIlZbocuSQ8Mxnrl/MznCY7MV3W2aiH0/6ZlQTahfLDIRa9HkOqcp
Ll4MOluLXndRVfOo1HosXrbXC0ehRUATt1njbzIH2tihBYpm7+G/sPmsGnoqLhiYOXXEr+Va4DM2
obZJekybKoqiaXj3efF0+kZnhve5+mc6QvR6xDtjJla2Ka3HPmtab0J82LZ8eHrT7WE6pjzGzjsm
NYxWtyONmqDX3cKyhuDyJBAgOk1mwXckRRf1bm3aLzzolJTzV5LUFfORU/zckbC5e2/p5StjJ9zg
4QGKiHsXdnjrC9jAYVQLQNUvGh+If9ryPvx1aCX8rvTmoEx4pzScxzUSjkQdrPT9GFnx50WGlsBF
kMhSvtsbldnkZelmHiKvCwcOG8UeDHMEfUZcFExuM85XrgeoOdCNgGURx1o342OOJHXcsEmlTcXF
J/Bu5ujbiZ3TGcUuVzUT733ImVDCgmVYjM6CIiD9++muLQOgFVEIeQEOrQm3+B9Gy2S+mX1PqyM4
+USKYuJjxUegEaPA0Pct7a88QvwsaS9n0qqDqrIyefaIyuRzet7IpfYm4c9h0WKE/wdPjF52fD+I
/aUqYSpVOwLHk9qjNPRJC776H3W+Q9VrEpW+qKbZCZyJZUHURJDZXSFwg0WC+SfJdc831WtkBfoy
H/WdM0ucy+5ocCzPRIbfvT4tiNlbYUR5foO4k1MNlbPHTxoKPNMB641oCpsAKAtwS+pfOIuPW/5N
0V69fUFuU+DSAmnbS9RcZ0O0TiRLURE19QVdGFAkih/WjrOoGIu58JJ599rrsNzYRUmfSKugW9wW
dVts1YGSEYCGvA08AdYUT2iw+yyWIc8a4/0j3ZOOQQshQZc3iulqwNVCn18GygrdwltOriWTNL+u
Q86phO81hLQUNLpFLoKX6HLXBYEgsUnoxs36jlDbukwu1NdUA7/usVXUd1W++eJ1PeI3J0iupfH7
eIABcTJJgeHXJKfaFhx8uHanpfYEyaRnMCmBPkV87M6+YmCuabFYda2XWkkzrFPUTUE8qO+w5yJW
MsyL/FPGC5QrC1UQXqeeTSXnjOm7q3srY620cSFadTs3qdXh08jMEzqSIxTbSLgPIOw3RcVuQPc5
7qAC/E7eNfY8yviJihf/h2t31btJhCkzUvisT2hBi6HE9j0wioJWOZypHU/XNcKHGapXPzp6hWkx
oIRHAebF7FjwT/IyeLlMEcWCfonQyKWLAbl18C/HKiylNgVa4dLaRnQ0UWqfwKwMr8uTlnMQTnGc
KUeuPq06J5V5Nruj/wyuCWaC4AIVtcAOCRCfqeyyV5ejCov3f0IBvqlFJHFP6TgODp9v/QJCVt/s
jtM5rh4KoEZTz8cvtqTo5bssGzzljeTfkue16furRgxYIYAs+kvJ93OV9naIXHEfzAg4WGmOfsKE
95JxGDS+gcZH8AlTxCYfFzwcoWwIDGpqTBh43B4KbJxR8WMyGLLM5xjNgGBo74As/y0XABYHtoJg
BYok4wy6AylJW1+/+Sv3Y0JrbGDbLDYazX+hETj6gofjB7IEansWeB8X44eySa15IFCi/xmVqDZa
tmYejh+Zj9Tu092yDdKBr43dWdW8pmErmg8M9fVTQgG/n8VCt7oBaYqwyXZHX/sf3n4ib2g8NV5m
0O/Odw4ubZHjWXDQAvzxNpI7YShfpfdSCXr4QvOqx3B8Sf96MaPCb57HPQXwF7u41LPEpKYFqHk7
OkkxRcrFHwLNAk83bsEfOIxf64Tw2mG7vKnxoywyyf2ZkwmsZz5T6vmo6l5OP0iNNGz4KVF4Htbq
GPmy9O++raWbZhG3WD7qVLZl06nXuYf6ZmaXnlffUf7FkIZgOzHkYpse/VooNdslG6RF9Rl74dK6
IrGnN9mtQAZO/Af1VjRdWsR2iymLVrZ3W9FCD5LvE6ZLnkmtFq0VsrShcbFACW1FlLqlNyG6MVTj
ofOGgZZ/POP0WBeI5/AyvolILJAbKWFj8qJcu8Q6kCo37NeJaMZFVqlKJAQqO8AkYIp/nOELIJrN
dINL9zjmOFuLxryRx1yU56/Nk1gKr3u1GTNcNaD7kuqMjhCG+PqYm0Nh35ogkNBdeQjomg995IJY
mVU+SZKpHLsmAjxJQy4Q57/DL+T2lg6cKP7VuGxij1h8Fzd4Gr6Got7afC4Z7jDbqvZVESmDiynt
miROwRDASxIgzIenfj1mFaTczGyvQ+AzIC0BzMuZFcXL2XGDojzLUjiRkxMDjeUoRQYvJNsOVQ67
lZRcsaQKATl20NabGOprgolaJTy+LcBiasUSoxUF8Bqj3P8UW3xgGr7miOPdrzJ7JzgEmRFyBPCr
AtYV5zt2irCR41GKdQLk7DXJqBoflGmJOhtEOc9NYkPYa+V9tUv/LTtznNSg0pc952FPrvhDEfeV
QCkI89xXye1ZqXhRSRkDJsrRqaLtRw0hEnt7KkmMprLPNb48I5WO9M7BT9de/ldhX5DXlj74OgYA
Jn7kLT/4IPo1Kim+C5LZe4W9othwI6bRUk2HkWnNqxos4duQYYvZyDcOHL6z5hdqql8sIcU4tDJb
OxYk3kqqVlEM/idw0zLYVfa5n3tY3zfn/8MK/oucgPJrFBxekxFilDot1mis4SXtKVEsFyhLZk1d
SAtUtj/gsLdf1dRIdB6ZzusmhNWgo2BOyvnlig2luYtIBUszV9j8uOVaeooXWQauVf23PfYvGIU8
mcaW9FbtFaOEWLJDu49W41HP9cCu+rHPvRAJzVOvLdTyQv9RApbPFjuI1cd9I2C5yO64fWoIoar2
he7gi1abGLijo3awkDHEF4YZVhXEHG3oV5J534XYF+g2BJPJC6ovmMlbaRWr1HfnyaYiJJarpUTt
4Iv2/3p12giejN82YRPipwxg9JMqPQ3yf/LaGc1axADm/+zCg0VN36qctbXgAATuPSgXRIiNj2Mv
LD5bm0w2hB/s1WJCi/10TCbb+DLSBfLjdaby4flhlT0gxeNOBqeDIF8fFw5TEUWGyEIDR4An56zG
z2hLg1cz0FvIglpo2PUvKz9HKGC/m27yvJit7sHbl3eq/23LmcN15M1QWk4cqetF6kK7OBQPM4bf
Bu8ZXgb7IMuYgT0I4YplUS8JNcrJdUetQ4LX0v6VatRGNoRT1EovvZP8LD9mosZQ1M4OkUtpuWg/
gAl2s8AQxUS6mcuj9Xd61LzXbAW5iGWT1oBSjy8nY9t80rtSiT8Ew7ocGpFGfVqFKKqcO0f9LDRm
TPwx2jBwEsjRNrSewlvMBeAb89QSwBr31/Z8PuA1ehP9J7OuD/LQr5EDR9qh4PZ+u7RgL1xmiTIr
vqIX9Dvvr1mzcHO5GK6DUV2Iql5PfstAO+QhqXZdqWIVoe0utHIShyZGUBy8BdX5iHGRq/yQ4hgY
wusOkUkdGaG7UEoU4qoYpdlTd6kSxQz+NEhdzfEqEiyyPbsHiy3pF5WelScSdNdf5XMNe9lO832K
PPkAP7PDYfDuqErNChSOAmmrgnEpUTbD+qFTL9skd7HQphxlRW+nqdWcFOXLbDLNHyaJvx+fa0Yv
Foi7jq7Ymo7HAjribhy9G/okQwFIKGFB6glb3BsJbHiAx4ZTZFc1JHU1ZA7/gi7tyu7unJNO39dp
h1hXmBV9PW9aMXe/TOr2b5tlBsQlJvxGT8h09DrG8xlnyYctzuC5OENOY96Ib/svKyxrrcJB2+qm
bYo4oy2iMjqibktnmg0hnRZIk+fOCVksH5VcbRHmdYTYDk8ZWIultVApVPVKTARwTN2uL02jutWd
xC4fcsFkQ3UwVkmgPfq7kd6qbLMetVxBXsy9/adsH0zjlPD0Mw+Uwt8+mosKpgEffP9bmgg9JBcK
q8fYvFY6NTF+yOgm2HpsBZYaPdRIl+VDHols51s3z5VRaUQxZ/fUpKE9qFHZgT9+Imiyq4EVjMVO
7fwYOM4BWrXQR3c/vG2oVqqRzS3YIH3ufVk5Dmn8wHXK2aXH9rAAB6H1DE+KS70M77UySRPRnUUR
7wremT/O4dOcSzA/2/7HB5vckcNX4YqUyC18Df6NS4mv8IBsyMn5xMSdBtXFt2Gtm+3Mf2jWtc5U
zx0zTLtI7/ur6lEEYDHfkx73iaNtXNgLjqBevyew8rHDaJPNyuXkweSU34PmV7/n5jCJeUo/vuMk
pJe3Oy/cHoV/t6P+FaV9rrpqqUJ1cEQz4qF5kw4cMD+DnJFw+oYJIKcffvcLa/JCAgot/1fmgODW
mLUDxRT1YBqNhgmSoVd4liHnk3YHlyL44qVFjLHknw8VPwcMe5l3eMxb/H03O6RU0xU64qiG7LbX
+j0/1GdwW3ZR5lI2leAbu0l/QngbrtVWuDL3Ix5jhl/0wy/Mxk+tP7nAFfe1tvTBpTaGl0OaWD92
OQbfRocWyvWS7NNk5TI4YMyMkiiEvkPt7rJnKZwYhnU6k/ibe1kNKsOwd4OR0hPe6W79g3un5uFc
+Js/WmwQ5PVTI3iCxBxfwIyPhWJeoWmr+PQTmVNgf76T7QkkPUmnZkgExmEcA9BBKvbRUrnIukCy
ytAYKHNQYrPKx0gNbC0ygehCr0nnkIvmRV/mdu1hbBTdZdyRqOv0qWwF736eXBhBS9cCqkClx4jM
4B5vdR5RgIDdnLQ4S/o3PNkatjXY3IF8FWauwbnADJWNzJAomds1VzZbS2uQbzR0v1z9/Y3ckhWK
V9sAXoEeLI5/GApwc+fn4x1PxNtDU9919ZSsFHYFr7RNicBWelYdHxh+XhUjA2vSUITAvwgJ/wXH
+uR/wRG3+AV0IHMfDHCGkRiDT/N4gyN/+YC3bea70I4UI57B9MV1pvkpTGAeEo8Sv1xRQ8NrjmkJ
VD4ItFqUlYPJe9vr2csF6BbNZ00uisJ9MCyhqTiEnjJQDZ1Vx1IH+7YQ0cSq+Qws5Ek0UTBpaGtg
wPCtBIYxlUyt63NgXor2svMuHKve0XGHvEXCyT7k+8tm1H2e/w2IDbTKmZR7Z6BP1GbNnUv8FI59
LH0riOrGtHI93Vr6y5XPlmnIPTN1E3ibNkN7hsjebnkKSEmbOwCy6VQthMm8tnI7xa/OG8DvGiKs
ewFidDKhw2v9rcJNqfioeVkwr0vRIzP3vjHvnXfJvA21eS7bwAG3Oh4ZkHVupHC0tveK/kzk6q7L
QDYN4ZFt+FRu/UgHKkRklcRpsY4cfyShRzyGbvm5sugajNLMDtBvw6BGQGyc7Beh9G1mjOaiHSBg
Q6Z5nJP3QmqyfqHSwghPhjdEBFTNyY8FptW1nWsfCS/4H0QMGqT0Ij9q28bfOPLxl6e2jrkTK4EU
XrdT1CcIGMUxudNHTsoLJz3UgHg0dHbyloJxK5Exf/yWlagyOnB4xE0irCQSVAy1KrqyGFhSpFqF
MxynHVbA9kReuu9FzLmSGNmUMKEa5FPpkICfO5BOR0tPi3pRcsMFoBDsCj4hzrfIqQz7adrXcUkc
T1pZeoZeKnf/DuWhy1gMxfKUThA56opYS5Pgggv7d6yUj7q5OIdwKkNZn9WEvXK0sN6gFJH2nYk+
S7FEK7LyIwVNMhAMiW6YICbG7KsTE61L7ZUdRzAHOSPfn/ujDdu9SIP4E1ZuxsPT6lQphGccNPFz
gFA87CKPPKtYyAg74Pc/bLAXsvbv68D+xVJ2s1/yxSq8JugxZpfo4jqbAVSc7CAgjVXtt9nvuInY
bGCXHPkds/HzAnXnK6x7GS2vfB8TIVeqG1ClCE2LBxKGxXG/KnqGtF9E9GVM/011BXTHYoptUvy2
2XK+5UjqmFcWx4NQ5BFDz7W14WJxcy4BAgE9bNUOJ6LzmWedzroir4HEe72BS/pC3b5LLB5wbmk4
cPMX861gy7dd12QPHBoLTFGjcXMoewcJizb8/82tE07Dp+WcI7HO6xd7EV4xEu14kfs40FNyFO4D
SMMnmdDKA/AzBIg3QV08wbVK6YSdnQJ4TqYLidoGfNJWeOdmvg/2wF50cVfwG1v5Ghp5W17Z0Vp/
JOct3VJqsIlV7bPOQrDqFHQLN94JMryGisw8SLEjQAXheY3sbaoafqkM5cmyPZZhYshaimIyLheW
Wd7umEN2WyvW1YUWp4GPL8Qlkh8KLkzMhpJ0rKfB8zgHpIA0w9SlzrsEA7/rOC7C5n0pMdf6Mb95
eJWJvrh3zcKOAvfXeV/2XZ9kyHGfPRJYp59AJ6h0Btn6aDneEXVF9cGWAl61/ScjU6ZEz10LMBYU
kCE4G2hyAB2aS2P3rfoRCNsbNTJZnjPoBF4/3sp8Jw9NqEkFWhOrXda83D16cNdnP1NWrOB8ecnk
GhxkDymgfZEF8Tk0v2WdHTpvzoqAm31joxQW9XA4aHQHNF7inTBl092KszSA1RuzdzEb0+0fmSUQ
BwgLCH1f7Ryy6piKHNAzRRIv92Ip6YaVzfDXW2s0dMvGjartsOFRL6M30Hloo1rvd11VigQ2jboB
YukRrHpQgr/fu2CB0GELp3mWxWTkGhO2WENK+G/5bqMCpHxDMRy7mRzX9R1NtKk0IG4DSn+xFqL3
xVW2dj6eFIo5qsqG1oSnkiGAtJmrIgzGZnqEltIW5t2n6QnHM9nvRsbhsFtk7cFZQyvkLvfn0f4A
azg7u/s8S+l04o1Wv0VUZJhkhFHwMb6mMmc6TK9IMV9utxdbhhZWa/zI6eFw6nPBugwcMBYxMe/0
qqko7DSsA0Y/UwL9UX/s6aVgT94X2nkluk/aiLMe26KEF3OotNqOBsuMfFA2NYl+hWXujB0jAtod
lmW7+PTooTWcpnfFV+CxbnEIwotJi84EMkl5IHkFKZzVFwTTm9ImF03FMlQurXRNKDG/84l/2MjB
CGCX79jkIxAZCRTSG1ZZKUqWU+hZsR4OP8C6mkAGJRIPcRvGxFwQS9jb9rPmonvFVyBhx0kErWNa
ty2kNg3bKkCxtiOKiI9FoxWQyy7PjBBwYKqLwhIvX1E9NwDkYFopXxdGVLs6tlE+nOvV2QHoyps1
+nCiB2khxc2lYPaivGkHDDrLRVhH277l418rzjKOzp3/v0ik4k4LHdDPtaONlKf3arCebXmxmwgb
6Rz3iRDKWiFe616VBvIP8Svkvoe6y1t1j6a3ubKvU2hZbmy5460FZ8ID9Lk9b/nz6X1RJgiGcixD
J7pdnVkK2p4sMmqMatE+qodYmYoAQW149IJmAvE1ZrFNqmkofYAFdT75ug3CI6u8J7oO0qG413pj
ezFQihNh/3oJ2sPFbcoDt/8JNRToUiB+H9ch0RxEfainXxtPVWs1cUl+j4GetX9KAjVOpG+MkZ26
+m1Orr8fEmTfS0lHcLgRfLmuRvhpJjwB12QoOB2NwRmmWZYYzZ4Mf3TkafoKYHvPJ7NlO6jHTiP4
wb9H+Gw7VpOLYTwU8XEzfk1iV0UG4woaS0HwOlOOSOd05B9APzLUOkcCyXweJB0yyF7OoMC5vjRj
v4LaecpRPwEo4Psae22VnPEaAXozv0hyWavDL4CdYoxSiK0dZvBb39/gR/+f1za4fX74L3CzzmM+
ou4qN705VTarU2HsdMabLxhrXwDEwnhDKT6qvDd2VpjMZp1R8VsMLPyRTYFhNoPkuGMe/6DUWIaP
eskK0AOempaaHot0W0CLuh7t2SzjVUOX5xMRbWQhggFrZvUxHIpEKuINdjkgFRnJtlFtNG3yeEr4
GHiel+7HMlwO3th88Rctkq88ExLz4Xd1f9dpNXNvemTvZqpEGAB+DoJ9JCh6BAWvDR628jOAJVrI
RqP/fNUigWXdyMrWP2sW/ciLSFa+DNM06+gDHozn4uHxT6bxE7LABE8c2XDUIkKL1uG6+6i0GVXt
wCBQ4RLR/4WoXvkSLyXxHX0pEhl2lTCskgvy10/IeXFoqJ1HuJSui1H12GVRlv0nX4c+5DXxFLBT
t6jaOmCPjX35/xigfooxg8Nq43W+C+edxguJ33b9Rosjp1pqyUuNdtJVp12sJLnAZwFylNLIwBcy
GO2M2WYERk4zUWexcGBOthH3R7tIx5NJibO6Tei5iFlNK4XGEPe7zVXzL4ejXP+p9lI0c/P21MUf
boINM+vdQSxhQMv5xZ/EKsay4Zn/nm++wMyxZ2pDKGQ71YnF51Hd5bFnLaJJPveKfvXMgPwcPqlo
nRRR07Z8K9yyE9MdzyMMlOJW5fpWkf+Oze7Xmpg+l+xPbEjlSx85SIhGZJAOefarWMdJcbPeq3Iu
hi4r3+jGuUgWY4egA3rLbutjvfJt8vqhDM7BljXxIQu+D1n0gTOLwSbbEdlOX+BZI07hxEuZiCpy
L9c0SV+SxmV5J3BZoL7du1N6GGyb8n9MN3W2alRa3OfUKVS/DfpxUSStmobf0JSce7vHiB01V99F
JVjXICD1Zy2VQbgJe47J4/BdM02EqqV87bdspP4syY2+5hP0kklgkubekNzQi/d2JA5eepe6vOep
5GR03B0mgvTWxuM880n7LhqzQ77Lw6Fmfojpz5gTrPQC1dH2MNaakNpXH4IMn1rb/VpBP6ncZWMv
vgx33BLyRrtc5dO2q4RJiIIddk0wNAW5pSf3DSIh6cbjrhU3g4nqnSYfuEAw0f30aXxmIuZ6FBiI
iWxYBzI1XnKNu23wQ4qgHTBN7388vwdzFA1fJ7gJdBut+JdfNb13802vwU6W8OWjhxm6XTFYXLe+
zae1tG2B7HwQTRx1Lro/NS2hn83FEtBRRwxGam+owwzOUBJq3d8ALsuwA5cDyq5OeyYTzvn/UIH7
hLyiErLSrF85ypiLPFSzCiultsbS1JsG1MKlfuCVX+Ncm/NOv7zK1CrZggoUIavsHbjJCwNgKK4h
0rzgDopCyrs6yCdDP2bYqwnEn+4/zqbGpcOYZBSDViYx3d3cQXUb5vx4evTUm8dJrmeTlX1FVPpB
C7OxHOLVRhOjMGWjreP6Y5NfSkUkmaZf/B50Nn8hJQRZSEywzFuSHC+vL4i6Ki5jcxf3XCwM043T
zqOOWP9MzqSlYpOhs/Sgg7wB0gGTakSxgTlqBJ7E32klnp1fCt6VvzziueSqXwOoVc3WB0WrwzQr
P3/TB7txtgjdTKwA8vp7fEENsACBLMmM+uYFkK06e0XdNTMkWoVy5H2d0pmZYbNwaIDZEY0Crfwc
v5WJ6LzpZaLm0CmjXGw3Y5WixVNhSf3GnOgHW4UludhHPZuo4YN5NxKC2LomQi5MQmJOGp5MK0ek
iJaPLV2LUaUq6KxtO0V0MePO3xmQM/a43Wd7xFRV2PsqyDgNwDUTZsRrswW4XWid1spJnGyTUsDt
sd9JKzl9w4gjHyS0qxy1X9JM1pUM7LKbWAyZYH4G3MgELJeFixrws7BScdC6JZlv0RTN3haN9AiR
x1a6gkh+WqUK2kPEJMtFOHP+P5EygHzxnElRlop3rrQ81ZlcE+vZJjxDZb7pgYehQbwph4fQySRf
1VUAGqOPwp8yHvFBMQAMJ9LOjyQBJFDTPLAnNpcs6PUfPWIcxQ6nU4m3KnihnyfJf8xSPbyEmofn
8EwnDfDGIFbX0x61vMBZHst5kApGBecN78RMzaQmHtanlNU++r8BnwiocME9cJE9R5gzKMC8pEDM
W95pLwhBaSOB/vQe58+KShU87srNdDJWygurRtD0u8c4l5grKaXYYHYuAQ5ah6hL6XkKVkvS877U
2iPQ6kwdWsIsBM8KPhMwSoWwCsdpobX8I1bjbpviFDE3iOxcN+5olJE7CScl6ZGbMw+KDzo5ud4E
5Vl5AubEowD7o+ATGe49RuYTM9DztzlUqzocPwp+LUVe5znbQ6/P3F3eigExuHj4ZCs3tDZ6Qk6S
fuow/TgU4OlWMCuyW8m0H0sE8HU/6aiXOnJ3Z7LdPMMPC7ucqVe4IckmhUlZ1hMkxlFbYVEUurQH
A3AXOraJbFwSiyHul/lQ7Ur+30wfjAzqJqytDUx6LkF1myFZcJKHR5OpMjlvuTAmtTOFvFRAgIC1
JF52nrEhuz9esFdGJSeElTEUgtdz5+IJOsyHaPlyZrB34ypg+IzzmR9sKO3XkLGBY8tAdS1iPKEF
qwqgBQjBXxntG0VoNqAgfb5qOgc7+v7xBhgGSZF0zeIW1v/wnsNZkan+/R3mV2wQKou9PITkumhx
SOQpBTb68ky2fscWiU01/R6Snq0G87fdBFtQr/d7zhRBPKmXT0E8218dpXPVtQGpul1dpOoo57Ib
Iut58LJb8kOJQOUKpMuddDMUElMyKjCSsHz6l0JxST60BZr+pOADmfwwOB8LF+Rf4g2ikaXitlGW
tKkw6ayRni3g8s1mI0aJL/zUdLBYRZHzDh9WFSNGVKHbloYW72P3vVDWp6fzUxOTw39yXpSXuSfh
C2s2uKtlBWi32DRYDY1K9XP5Xz+7Oq+hUGSZTpM9gorsqCc08nYm2Xa+7TIc5DhRGMFRMhqL0Xss
A4DJUDA0BYNHg5p7dzWG0IjGtb9rHDojzApU8D3sDhaH6jg0GRSDz34XVF6a1y0PP93CzEQu5+5U
TderGr9Abeq0qdm3eyOTKJVqX3tqX1KCREdB4f7+eMzoDgHeHbg+qKg6HGbB+KKNAoQTuUH4dGiA
lqXVCNCsLQ0jrojJgTqzQ745sKXJFKtBfmPjiV49RMrt4fzcJ8HOL2dNXbzxCwjxNOhUzOQnaNrU
LZ5zHYiCX2Vq1yJuMgjRYmIOlTnl4eH64VewziuygSa/JGN5mkdsy+3jStPzzsogcLYyXvMWzZA3
T3pikD1bZ90d1Ml0lqGnSFQzc0Dp43Hm21KPGVaF7ZI503QJy77T/Pk7HrAY0GlVEmaDGBdV/ISh
GTKmgDD4/sYWW9d5oyygbxw+uVYr/HEBSckbsAuEs+ANEabIYYuPegcrPeN/Ue8jvfDGpcGiGu3d
6zEZQQul/jAAdQx/IogCoq9kqGNuVp/I9aDyGt02pFXeE1juu5OWw20Vc/XAJLO26ECzoyN9vYij
a1aYVOaMw7ReA6waFtd4LL8TGBoson9mii4btG8yc+DwU/fGeovdH4IeCLEIiP6FwXhnyjTWBOqP
K0Uj9BlddWYE8J+qz90DpMU5fbmB2mRUSRs3oz37skKqdwbvK1G8Hr9GsEJW+9ww7cNIa+UpTB/J
UV+0MsT4iPOyz5JjGr0Slno6RHlWOMlwS5Pj2rWtikWq/PGs9v0jKfze5p6NgbUifVgAxyYPFlwd
e/npqu5K8McrOqhaVPaRacAE/6IGqoloi8FhYcGn/S2BH7iC6gzrXEMPIj+ir/heTwpFaU5SkAqN
pp4fdmLsBMGvM9XgAgssHWorsfB7KNRSeIyOwMOwgKs46aDU5xYhsbK6dXwrkNOxTjNjJDSQNW+E
rpALIiD4Vu7OAffTIEhz09tauzMhTRAOcZpcMkyHPuhgviSo7zrBjQawwZUedxRSk6PAmAJZMdf+
lF/C+0x3oGnETJotHryIW7/4t9VxA8LZiGihIVXIpbIfhmsqtrGw0axpLofa9as2YLPrJui15EkM
IwMDfV95nocnSb4KMT9dxPIw9/nu9n+4zqWR6i2nlUZieRAFesSfAbvmEeYoMfluRnYqyhYYS/XT
+KiqGHZxvZquWC6xwt5wqvmDr5tdvlejO4MEFN/QvCDhSUCOKwJctLX7ZIsAZVDzncErojow4BLu
xIrFMU8Bn97eCAtob+hk9Q2H7b8qcFb1n1L3/35Zlyp5PfALbNvSs/lwP1z0o6yHlmwWewVqGvC6
Y4QAcuKzzvIaUXsPx9S47SSsLW3vRhJRkxpCaOksO2ZXY1WW+Kmblcxx6cp+L3HdmqQ0VMBLjvMo
tz5E6IrqqokHaRzBsxdI2lqhT1mGvC11SMkkYaASFU6idVGrjdVEnPdbrFge0MON9Nn+Wj9LFPdy
RzttkPkPkNtRfpzrPKG/9bgEI8be661IH+SUqIAYQ84//dYOZB1P3dmbHdGCXRwhBDrpNnhl5PGE
4SPAgtXPWeval/cwX6b1sBbs6xun1oLfhe3VrPxRSfXS6GF5hPAGFZXovFXIKr0RJOM9A7zKCvVB
qTno4aWPRcNdiwTABL9LvzZLM3v8jHCZPPRo/fhbKosjAYOHH6s+r/MqP0EGW60ORFYgWv4ZVTPO
jGcrHwKEkRHpPhjGZZOWTWbqMms+NpYVtl4C0IHS9yBd3KSztSLk221nkhMmNBA0Z5MeMfvYstVf
L1Pmnoh4j/JwJFLniT0SmU39jJ8A1akVMCfmnpDpyCX1x4c1z1G+kdTKSJ5VlYwpVhMPWV4ktiSB
Ir42+Hz0/WeeVxDhfoZIB2oHmdTrJFcLcjhLwgPn+CQ3ETBvodxiouDwxZ6/AU/lg+WOMXlaYDTu
JEavdRP9ttztJ1eySbBg5ghPCGEaSxxic0GiQnbCiKkYrEsk1AU3T1wF9xMqwL3DIntSREEw/aRT
tD5ruz/usXKlwf/iLO6ylTYTxpflJPbHYcxvGlYk1pUDRIqqj1iXq126bTY58pGCT53kQMKxUVda
1s7jeoEKz8mKVv6yIsVcQN9Dx6ZXDvdwtezR5uRw6egx4ezTwcb4J+Vg4qdsbgbBw5CMCcZkxME0
op6A6zKnO53j3X/XQvKYYPNjAqOm+2ecfW7Rk8z6GUeH5V/viAoUCkrjxV66fo6Rtpji4xQSY43e
WveROx+Qu9ducoRF5ahXflXTrffu1KGWizmD8KQfkkXtWWO+Gd18dz1Z7Yh7WqJSUabg7Ywct+Pq
xZnBYMUBZLHSyK/xjfeo1C+EV6yJ5sS4Cn7EX9Rw3+p6defzpAP1+nHEN7Wa0qR+LvoPvrbt+m5w
tYVTUNofa/KaUr3BLhLPxApdYenETT0qbuvChAAyijzcp02ZmXPTC4lXzTGumFn8zyOtJMwJqcAQ
7SgtbR771QkVZuWu2Ks+BBPTfs+q4DSnrqNOZz4befRBKIY3Pwon3DghmmxEEQXIospH5OiUMfIT
51dsrHsUwldPoGJyJlXyfaZJUhj0XAygq94aU1es85CCx5Z3m2oIoLdCez4ZoxMU/7rRWLlwSsZn
lbay0u9lPa6QzCHd3jmyQ+YWLpl+wlkBMa0z706Kiajt4jbIfsgZCZ0VTItTMXNr5AldZNFL8twZ
7yILwT5TC3v5uNo8OomGCpgZ177HP7TM/02C+2JmKrLKCkfRB+sOWzI2077ztiXec0xp2p2Dge9N
Ly2mrhgKdEujJ1kk5C1Ql2u2dT7rsW3LMOkh2bT+u1p9gAt8xSG1W3aOCTufoztG9B6LwbKVQDGf
oioqLyXlRj9v8owjc/Yw6FRWCBkEkskCMJNWQmj7UC/6u/sPjTiyd5C4ltLpRPSoj5xRVq6+kYZC
Gr6wRDzw1pqRB56AnXjfcRAhLhCIfOuYXnaiwd4TExBEfmkRnBs9wy2jpp5UrD9LhuIwenCdFTc9
z+ca5qVvz9mtJJ/z5tke7/s9ab2p6eVQRLrz4Ktk4yhYiO1A72ib1JMF9S/HJlaeByTqn0rsI9ZI
DbGPYFMrtEBjH6m/JnGSLWoPVfJY74/yywHUYuDxDjbRDD/mWaRvUqxdqTUhFHoLaeQh/Is97I+2
vJgdgTaETQjY5Ixz9RDP+uzgams3x+j7FG5qFxBkXBerPfOcQoIevTp200u5wC3zXiyHSAaZHGBG
MfcreRkxhnQO1MMBUihCQT/pzYnbVz9HHCyyiXX/6yAY1L9QjdInS/B+Bx0iywKOc/FaRMCOQFQv
Gc4qOVy3+p6VpO/efc7Z/3obnXfQYWwal1gwtHTQyKAk3EM8WwK3FmF0fyHCMHkiFuTbZ7QvAqEd
BJaI188k3T8FRUS34KAZL2jCHXUt/lwyoHeFR6L7vVF6GK7meuQBe14K494QSiJMd0BT8lUvWZxG
5NZntpkmJ5px8vVYAk/1ER4HM5zheJ0Plpjte4UigOsxq2ZGKHe2d8grbhfUsuG4QnTUyBtNqLAG
GGJ+qtYjHJXnqa8YJFnNxiHoBtDIT0cFi+j6a96HKLpxRFa1WPL9sCRogbs77u4BrLVoIKl+L0ND
M2HCAfT19QwcW0HrJkpIjkw4Oz9uxjO6HFiPkKU1ccaN46rVJxeIkmJdyB4d9j11kQCffHe4xw6N
+7C0Y/ZH6AbMLIA5xEOifv7CDZT6vTaLmtesvKZrutG+U7r27A/5BLKxM/2qTfoxCyDWRoib3Gqz
H5VNXk+qt3fryWwbgWyMLEtNfy92bioiwNXFv+4XN9SDPqF6TAQpaMgguKPhsSk5bxYGZPW1IZ65
3v5PMdK5k0PxiG04ku7BA5WoKs51lVrQjK14BmcPI6G7/P+TWu8vHPMRYdBoi7eFS4WorY8zgRol
uJkQmKtr8kFUZ+07EWb4loc/1DB15SE3/In3Tpg58LZpJ5uuUeRNELIfP0jN8BFXI4JGNnJMOVsa
et+2rQmNswws56oFHFtr0vfBg5y+vHm7hgH4U9Uo+VogydUCSfZuphK6e46KvMOUdWxqAe+KO3Rc
dL3llqimTaYxEABMP3Q39xVBcMKpt8znqAJg+0uQSsSAJ+VgfFoZwuQBqKjDzKOvy7131orNuEKE
91b39FsrnDjJQ2/GV8q3ms1rag1gtHb5/MVuThzaARzbR2T4wh9nSlo+IRyKJ39J0T49bN+Pc+sq
VfwVa3NZ4hZxdE8FNfKpZ35ZLK3QDsV4y3LREmidnyRLQHR40Mj4X+XTsRnTEnT8oXnqgGoTEpZC
Z1BDn+tOBRaD4voy/cRJPVK9/uTgAOHqGK3/NBsKSXYPDSbxD71WSN07ach7nWuBjFcsQRe6Tzad
0uXvEEna+uM1wVy3OxletfUnwNBhdz7gWelgo5rrN1tPvXug2VrcJ1wTria9zXuSAOW6oBaXhvv4
dQkrbSR1hWT9iNU3EXLGl9W2Ga0wMEfr6A1G+mhjVhZp5ecBnZjbRd3PvB1DszyAPZp1gVSK3Fzp
iaES28EwLFUxs5EPbR8JYAfyBnAC6dYDRtz5j4Lljl7WLOLrxBZPb4H94aLQvUuePK740SzbLRZq
TOqP5zsDWDjx94+JAh9KNYcjddhS8hqoCUYXBjrNL5pnD2JoyFBlwiyLiPcYG+spRqmvHopb90M1
XoY3wicAssV20sgVfzOtQ82DV65MaHkTWJRcD64YIO6QVnaK6ABbK9Um2YhY9WX3r+p/X63xWh90
qsB2xs31Cp7h3nTLMTotWccOs+YZl/6p8NRJGGO7z8/ezEUC9UpFU7pD4JG5zcg1CPMWI9swGmv2
yw3PHO1FBrvylS/mSbdYR5lzDvsH0kxwx3tEc8LS5/r76Z+uHu6gUsAP0yPpBFDuC4FBwFS8fHcV
rFxMsMyEMPg815knkpSRboiCUW8b6mIfmnsT90e3FBj3WkaYNSdoTGVlH4poKx72QGBr1KsV12sB
QaM/iydPCIHzrVZ7dkGK3jz+yiAAasGoJrEHLeS2KmZ9ssI0rbGs87vfZmFLE8pe8xmJC66pT1ey
9F3b1KpU1B0R8mhd8u9CavyRInnK/xwApM1Dv8Zr8vTO+ld1RXvBDwsDKi2F8O2waAfjHWz6JR6Q
yFSArKzmxYmXbktKCM8mfV4gVDWN4rkgzzrbZPDOUjlSaZvEiTCynrAhNoMxHqPtmS/LEk6bQOBz
LHjmmJRuO8TOK80EgsACiRiBScaETzQIPv2obp4nIlDLN5mVlXaUo1XZTwMZJBPFLRQNj1tlcY8e
580Eh8pBFVCwu6lslPQFX6WI+jWzG+zmDrG6gfmMu+dP0Cqmiz24WdXmheOIXBeL8C5Xn21zhZBU
sgi4thcoDPa+GUSL8hTgDiKlGObl3qUyw05JU8qclZQMHjUifH7OZO0JQxI03j0bEpj8lZzhbwF8
73EDjSqErrwkCYfwpUKsT7CbGNgbxytu/RW4kgGoDiJyPJR0e9eqXN/YlgDK2oztW8n8xYbHcidG
t3lcnbPWBAkyq4Im4rC7Jw503w3/YS7m8035cZQGEltel1DCgJQ3DoKCCeETI5ISyRB+mCqVEHzI
A8R78uIIL0AJjD8eLIOuWJbi6xTI4JE1j6GjRponfuRVWCG3KwaQBpGjqakICGS3znEHTkdISi7r
73NAAUW0ARhqo4T0OB1UgH9UhtuA4R9lP2YyXTWDw2VegKcR4Hl+ClrsQchO4dzSnuH/0R5PqMfU
MvSQHXlR9T+a4fa3eSablzrZuH0Y1ZmxgM7kXrHLWcZRic9RMZc+tRO3i6bvoPifZtGiQObDaP7F
SJC9SFoktIyIi1cePGsbJg8SadquQbgoeaurEkLCWoJrMEIH1oUVbmjpCnBYhiDDcjDLo8XQ6g4Y
XFltQSdzuQ2QRrmeejc8hWJl7HaVDWKgVhYE8U0hNDrLvECb/VQW+aaeKnth94+STZx4PNXwIepy
lQsntgQ9oFnstmKVuxeihFw5+MrsmyVaRlSChe5eTXEKRlCKJo47rImB2ezuVFKQ9oMHp8lGLpJq
ET/s5o6nXUJvVlawzFNnhttvivLB82O+tHMPT+J/9AYZ+NJSdJ4CAJ9RZSathrJMR8FfsNOiWiXX
PpuEBrYsPSIQxK9Cpqo2afKwu2GxFPs0u2h4Wm2tCIk9qqszcnWpXwdUn5Rs1/fPFyPPRTvuwUR3
q6AxbUSQyG4bv33TqVOGgnYcpjGHfjjsMP2ilG8gendJNRNn5VkeEUPOw0EgEp/OrEsB5raB1JuM
ZhIWkr5leXdAqLPOPQdACOvNpgNkdOOrwFbn4Nk6Oc4t68n7IrVaVHAyj+HCYpXoZxp9qBhLI+Fc
zLRYbdrRwtInVlG5OnsIohnhR43NCf5v679aB16HJDoMBAMn3W4/Bs8T3/MDemjCjd5OUaCkjEXW
qUVx/RbdnCQQw49BReslUYtyBp4vzaNZgaZqZ2HN4hZdaLGNfnITuaLNx0aLZFgjxEV+aZGW16Am
podtRJZevx/SbLAXnkdH4Bj4b7ditfqnsgLuklB3uMBj63+0ioRk/FFwsW2Al4mNJapwkgkkA3Un
NteF0uYecaOvqErr6znRH11eRkEm/qFc8RBOdsf/RU6eJll0CjU49vgznzcZdmO+TnLZNw4+K3Vb
vsuy62EEQrFKai7HSdjkhTl0bmfXWeBoEJz797HpExDW++eCdx4K3sRqBKwZMWut2dv5UTOwxftz
PO9rM3KhT5rZaXU+4RwiV+RG73LRShbHvKVeKzZ8hGg/a3F5UDZkzZqzkJyrEqk7IhiufwlU+6XL
JyXuHT0DDGOW30W8z5kxKNWNNA8PC0sGNakiZ/I50UQW+oD0rB0SxDRebeyODMQFR52YhctyeXkR
Su9y2YHa8xQKtdZl1utdTAM+e4NocJNtcGCDo4dCM7MZZnDm44rW5uiLRedeZ8iFpFuk5HvumJbW
2Dytbc4aaja/1q4zryLfwFMePCuSjzAfdZFgLytCeU/nGvFLfpUoIQ1DVdTMJM/stAB7BqjCbzfA
ODgzZC0SABXcbGEp6v9+eAg/YSb3xPpxqhN4n+M8pEli058yt77rDgTuNtz5qTCefVQ/lkGWNkD/
sgry/YjLGp/MkHk/hCBXC5HBXwAgbtvFzfN7+brWnthWZW1XQBnEu/f9pj0dZ0WtbWDU1wT33VjK
2P0VdEZL8yOahzzsII5Rkt0yIjPRrCjahlY1qcvNAXOoLRSLi+IAAtx9fQhxugLdMpYcwNLV+9ic
v6zO+kd/qjVRbdgzGcqwrl5ZSzJH8JstLEA3Wq72abHq5SwC49p7MziTarkwY8u3WI+zApZlLrvK
AhFLnS2T4AtXr/vprqfexoadIWaMJvoNT86uadS061blNY468oVVHKgqAQ8sU92/1ff1iNLM/hXC
fyDqfOWgEB0l4RvaTCHOwbpXoNhgOhIkyH0n258oo0DV6NXzP23+KIoT4XqssqsRg36o/tnX8Y0X
zaFB8bQ1L7VXYrQbNRYEgZA3j2iXnFcPTUi3SSOGwRdBAuuK3eKUfYO4gvDnwfqXqcJDR+Tr7vA2
in4Tg+KUf+gjUrD9STDgjR8HGnpNaQYoFLzkLW+Tg6QvGCOzawT7432rt84SAT1GXzvTsqoQFq7I
hkfJsY3r9B2D/C1BvxCrsgnpOsRmnXTjg7rmo9iD+c/uC8Q1TLhNlf3BjGgy0Ut4AEjDCA1/ZNxx
g5W3PFa2jKOyWKbi4ll/kH9K44dzXizNfZTLj8JemJqxBtzqa2/pI8XvoeKtbjq45byHLJ+yhvV0
bVYkNb+oz7wCO2AZx48BX8LntDw42QL6OTrTkjBf6E6rQZSoGTZiCsOuq09OdA/W4PLzk3ze30gi
swfGpnRPSewK1DPcOcEbHVlheL4NMHrJ85lCFwr6OFCh9kiZDq7kGzjJfPHDS6GcfS1XBD3VlBnh
t4uvAQxzN1An3n9+gNcGf1rVSFyJpYsvF7zTr1KOL/sQHw003SqZ+w38j0ih/R4iG8jARht3ohjS
Etb/4mlqImPAqFNE3Z9I11he5y3kSFzYzCJE5wAfaOepMdCjjklViSZ4JF8IpQ2tKO41onHHztGJ
xuU6L+VKhT2ksLlEUodyBsu0raE7xYu/J1zBtBeXUMR0dmVOjCrsOx6P7POXKq0zcA+rULS7GB0a
5kBbwrV3UeJrE7kNUTU7k8qqPpyQvOKDqrUbFYgCMFzQ4mJa1RhboUuQGUvQsYQs/NAbR4013+r/
9T2LG8AwmO9NL7wM4kv/wTn7zteTwLZh5LrB6u5Ljzf0n35fPb7HVkiOXPa3sR7M4vybZf20Clw8
7xXpWy0QsNJMJpum9oSlVDwjpO6vNsTPZD3zm5KD7NKOxErcaRnJp2ARcbfoUmMy+gyI1bUvV3d7
D2Ww5AcWXKXDzU0WpoPYr9ynga3zkJ33WN8iZodboZx2KF2jAtstCANaH9FTJs30VszYCmASrsyy
VK+vonbyXIVwmlBw++cyiMKxfhj1bvvHs4P9H8TD7ZjsQjDzL1BHwQ81QYuLYfzthaQWiuP032Li
HNGxX158i7CK0/fm0smmCy/rTPE05Iq2pl5Q51HlV95sX3cOqWbcIztmBm22jsz3a2y/iTrI7bL7
Xe8kF6Ok2lrqAPQ2V/hGiEmIusNPqF+8djhNY2HolTT5qmvvxZpBvLKix2uTaRy4jXqDme5TZiGb
3DAK7bEpevcTo+cU3aug3Spc1cUvt0lxZ+FqAxcO6OdkRp85cdbym5STmhk7CYu9HdoLtVtrVTGP
J2WjyFBd198zTKfPmJnUD1wOyJtrAIwfQcMzjaAVWQ83YymWNm0kxLxD6iTDvlkvcTbLSuw3G4zv
Ec8WUt9j5u/5wc5M8rwy0eWauvUnrjeIksOh9C3kuz/iubGiXOvhtOvMRAfub0vbMwuivEcMITFs
M1buWILfMTTUsJiW4qtnH39S6F/ltcythFOwNroOzuHBl6vQIUVU+BXxjRHWDvB/da73HLQfsShk
BUDh4sMkiJeW0JYZzhVwQ3nyPns41orw6RbEQC/K6MsSW1izII3ALpylonoNOO3mqeq9ezC0xBdQ
iBmRoIrk++uEHnA6bX6uluvPvszN2BAXwll16l2Co5JvVpqgqFLF8M9L6FEEE0mq2mIlLJymhuE9
YwcUH3owqUW8oaWshjbVQhN3GzYoROh5OVMHlyLe76WDIsQ4MH29UVZNrBlFkIDyvzHrKQTpkpdp
qJPM/12miR9cj2t0gx9sOMMbpNw064BGfbAFlT0YKX8FcAv3kqeBZzaH/2ut/dwnnQe0SgdylC6b
mgdr+hRPmbY9z7aqAENEn/aTPEyOBqxWtFrcJBf9aS5Q/Iwh1S3h33ShGzLA/R3/kJGT0zYQxVju
OuV9a2NnYl6Jd5ttRH5soa1OHvkGjhn7rAgPdzZK2aMqEuBB/KZyMj6bPKyl38evefVpfQUoqt8C
8KepZbgJb9lqLGPKy/TAknEn3DFPrRr1JsBmx3BXCvP+h7W52r2/jHUZ00JaryeoWlSCyIImniK4
XUa4AxjFlHEPCEUXzfbGqPsIGdbKw2UqGQM1TaqH6BGq9HtPOzoW51C0VBKu2ksYl9I1xxD6fC6Q
NGfP+uR03Xw4cDFlHLzOmS2L5ArikKzuEnfvSPkdqhpPL5uYbjvfenvYMgTEznjx/AQczGXCNGVa
hX2A99nZLhLRxiy4IaEjXYN1XIPXApbk4Efo9K/Uj9uJqqSl1nROigpVBdGTzIPP3+uw/2j2gcye
f11RXNI1lAj+uxzVOksLBGgeBBUW1//IWdssWXzaDXAxKVxDMGnIkCd8ZHaOvXfUtXlVFUaA8rvw
JowHHYCyIm6VNfT/HS6V2oVHCuXCxagPtCuJZFVu5Bkw7t/TDKpFE0egf7puLSZT2ghX+BZqLfrP
hTqmXQ0hcGUiUIaArCIfqbY5bPGpZAilYbZna0E4iKtxABNiTJ67KRBs4SN40EpPpuo6/EOB3xjd
MfF/h5Xufa5HVRYM0XgeJbYDBp5tYR2jAIaVzueEhwbvWh9H0J2uwrUSC4YbjHgVXewRe2ImzGxS
8gH7lzKf5pZi6ZC0J6mXtZclERpzSPjOIGeohbFl1s257De1lecsmxYFZc+xtDCvcWVOZPMfxSLC
qKbGyG/Sjj9XiKZBl4ZYhm9oM3xrfxAZrVzz0Ec1Z3WjswNpqRCDe2od/83R4JzZpEI7sER50v39
++ypNV2VtgCXMQ8iZt18m7kPbHA5fKrKrFrH8yV1lDVYChT4GBuIy4P1IhviDvEPImCJmfEZ+v5K
fQlrmgcH4obvaEO2IL4BruB+K+8z04Tvas2xz1sJMcUI0cOvkbBgEoaMBDjb3j6cwO3oSWDVlRis
g/KAlDG5tqrBDE2ZBx8xO6ZoMzW3s49cF8E4z7k64i4bKA1kN2WT8WhpxgwSF8p76u12qi8oB0GF
F7w95TNMpeZuDlqksluTnP+s7DyZNUihUlcPxqm6ie400flaWyFNSNoa5t6snRvBpTuMIJeqA03v
yh9q7U6/rOcMsOReEO43McjB24powpN7G0TNg5sIVbg7MZFWkAhUB6Qv/F7z0E+3kH88DPxSvVkt
1XXQ0yBitPDOvG78cTSW5TOy/36NVaWq0rsu0oV6vpNNTPJpDY72GUSKDk0XYFD7IKTuhKSnclL6
5a3FYOeTVs+vvlSXT7ePb4HVCt6gA1+K8hPTUExjLOqGx/y5PNgPEcacyLIcpY8dH1zFDZDYROlJ
f2sUwhYeUNHPHBTrZowNmSvw6Bx/9JQWT4AX6ck2Qzn60u/g5c0Qd826vzrGQenudz2/ktMRUbcU
3Jvxq0surzwqjyDkH/NM01Ej1s3U46ex3RuhrR0/0n/wI6qK5LAI5tzvugGXWCnIGTh6CMBIDmY1
wPnhfZ15v7ZXRMGRvpfiESUUejttlQE5ReFsHRCajH+66Wi+jgo53O1Gv+FkYmimoYwntsQxY+y1
7/w8+6KBNrKfN02k6rHaKYqK9LC5avyJE02KJOrAK6tXrboaI0Xjdcyt+0VnGkz7IgYUV5RZZaGU
qsIBYl1WDJlsl9dgyPCM5yG5W7spJ1+C2r1vVwNYFnT4cbxIQSNkjLf9i1WS3yaxBZFpOHb3nAx/
r5T6IJkKHIg84fv+6EOmo8KCuPvZD/MjXL+r32Vb6S8pk8mXSoo1jwkPPZS/+Jx6B6rtNzVZOuLd
k4K5n3CykvuLdmDpNdfkCLKru6eYbqzTbcxGX+tATc09rHHDoEJxhK+eHBUdkRIgSwP8zMpG1wSJ
9Peg/Na04SIyHWsVwXPw8RSs0kGsAXQm9vKZ7rF15ap66JoYu/obcH7CEW6vL81XG/pn1hQGiWje
PKPek6VtsYyP5BKbmwwxmt/KXtzZlLsU56VJuq0s8PtuDlajtE3qW3YSC5OBl1fZisgTrqtfoXw4
9qkC26vuwFDYfWhQbSHMzsoPHodZ00Rodte0BaGpfanKzLSWhwrcB1IwwcyBIeCPPQ9i6dFJ9vRw
94SKyQtmkdkP9+iFfh9ywoViJjDPpIogKVjdaUkS36BFXhbxGsw/l13E4scdJyJftMMZExkXWAAq
ztmAr3teBuqdxFQGvRH2S1T6Gl7XJrRQb712JFyB7jyaELhv5WnaNCOgMRU6DQnabiGIFdUYGyup
zbM+CaxrqC19CRwLqUdZwiyB8RWRSs416Mq/+zEmW3OncduHpLmwKsICqMmBGMQf/qKHPbHmsO7V
CNPUdrTEm6nRZnwYtgUkPOg9tZssDL7ZIXSK3eCTqBOvPOnTV693qqHRMzdfORMgR5L68x1+bEpk
VsKdxzsKW/jK2lpB9qGgBpluhL1ODoB8y4zOKjSlOphUzMdrvx49m1k2hoUb40g3Eo2EBhXaAm84
Yq7MV9QYS3rGgKIB9y2PtcFWRBrpOlZXaXj7ZJIUXcAj3ls9i/iUz+BDbG2JhruMNvD0MgXTSeLs
KjhrlsVQrXIuodpEk/VdjTsTcKRaQ1qy4z5fVSk0HlF5X9RE4yQZB5deI2RLBYaFMEkI3090SszF
sjRDJJpciWZJeeYyETyl0He8lFla45dsL1ZzO82xAHC857IBJss6ubnURIdb9HDWqYbp7SWqL9Fn
q9GnsUGvDXvRQkmTQ+//ZwzQ2h5RwgC+n8LCSaHIRl3MVgXfbiMagxsgRTAIaDgf3hejYF384Wnm
mpeuw/yznPNtMj5s5gRRU0/Bx79Wy/wAIU9m6Ud9AnkRMUEQB2aGyth4ZnlwR7E08bTxZ9NjthgV
LGhOEFXz0lpdPdjcacLxX+IAX0j9c1Fzesde+b7rsITl0GHpVRt2FFONzLpUWvxeo28ApmxWfXfg
5jLttbYeSKPnkh/pNLHcrWtc+PTH0FGjJPXqtsWKjukiuWTcBEUBYfPEF6NGqLLyI4MMi7WQRTCr
L2HQ94wA1S6oYbfyeiXBqITboSeAnKAYPiN78UXYbbtcfo5dAJJy4dOj+Cqw2woFpfaLXZsrlXKm
XUfibS9MgW6h5zEiQSX+PleFQmtfFovlMgOXCEt31GiUCM6BjBZTNIGZDMCi6grrqITZRWsib6zS
qCH9C1tjvDewcQD0B3ogsjt1F8ujLL0yz8D2IFqaJMpc/gkt9aYdajBESuA/9Do/zkEhA4mCqBNm
QDIyHLkBXK/CCF/yVZW+3raI4ydRVcC3nmN/joOjevMBbdk56LeWrY3W9ercFPpAdvQ+6qlMmmKW
yG5CIT5wHCaNHFNpHRskpOI6EOB6W5AYm86GyCMqpKsYV+u91EFSxz7KBDyxrsgLlk+kYcvkj1Vj
UBW4/yA28qkUYFVnsyDx9TL06rlGhXPovIdFooQSV8pxXy/v7b2RWC77hWC9bMo8hD/Q7dNZN656
s8aixfR+l9G3wQcXYRtP2+0hQSnpXKtEMPrkTmZZbIstnNY4PzeME8xuO+mYxay3eiZSTPHWfK3p
3xl1VJu9CYgbHUIJXdyJP0rXS9YkIJV7yawhWIWXBI/ay3+lE0Z++pRQ+jTCfBdbKv+lGmLvqZav
NdaaXpyD0kl9WAcDuqsTxMYIKqoEBiH+QgXC6vgaptKCU+RZFMvFJKgfMfLUmlm4/hQ+9LvxZk7Z
QTF3/5waeAGqsy5+OEV0S/AMUApMdj/WcCL1CkY/CuaUV8Rba0GrHHZq9a3bU+TD3RZdA+VcoqVn
Ex8UCSZuWgNjwLFFS0CyYTOwsfIEIA+YLsZBjg+nXdRmoYLds4U/m2zL2clNKbrAuVB//wAjSGH3
1SSYDQOHmH7IZtP379xcxaiznc5ni075R1ifV7Yi6/fruBebtNIXaecZK3QL+f0v1zcKuJ0EuoHE
JNG5OpM41xghjxSR47OLGoigQzoppjNldl0T+3JN7DKEMSae8QtxNfwVk1IUgHgqKx6MJsHlJxMu
b16ULG3bVNuLO6Ajf2Ndey5FTQOf8fw7y8iPD/pzOaWBIiG2iysMG2sIwfEtOzhHeXLDnsocfTov
SH35J2wjI+vTd7AkKhbMqFYTdthuQBME0/1PS7hOlKDd9VepeuagAgWRbozqjV77efHwCoJIYXuk
r3HSHJ42QSCyw7zQ7SvrzmyHHmJiv9aKPIVr5ZMxloxQ1Yrl0LWckSvpkwt2q6k7xNScYBHQqWKT
h4DKZTcpF/hHAdMx8dE+NN9vt15+guGgz+5nBP1MVObtURM+j3pFh071oME9rmt7MohA8DJ89vNp
/qnBpGQaSOj0YUAFO3kPt9gSkaVGybKbbTefxFp0hwpJNd+KgyP15lFdrVfsWWFzsnyQv1usg4aF
2rg8cQr7c8yPMfIR/5GP1142O4Dgar33dNsNGLv51bEITaRQ83f+c01y5nrk4glBDfP59n9iKDml
uKTaUh4hTafS3AwMwn7Fv8mAtK6GtUmo7c0YV2IXlPA93fuMbWTMb8LHSpM9U9ddn6kxfYpYhgUI
EKN5hKFHJkvX9+xr1b24pCpBnaU8EW6n9+B7lwrwCz8jNUvsGbWsycLHUOc60aTOeBFwH5iHweNy
ry1G6gnKQDTMFsXNYoK0SSunWH+QBWF0LuUu78a3S3hec0fbRUsw3fOOFEij+ob0gU8fn+mqp1HJ
J4W/gmteVJ5DyGIdsOTh7rn/5X6nDe63Xrg9iHkfr8WeD0MeVostmfZHJXav0pnb7J+BEhkOrkWs
bGp8rv38Fav+sqELTqTFTwjJCU2RfCT3o43hrPLuimyADPSod7VvU0pPfbQhVXCSxgXXdY5N/EYl
SV+ue2rriJgtW1IMV02YnE9DCIbXKzCMh/kqrVUP/EedpIHqi6knHK9+C8cYQwC+LW5nOHj/t7WD
+oD2o4NEGFAOslx2vZOoWXVNCZtoiEQtziaLYEtH5yTy4qfTv1dUkZULbabn2ln4/uLH184YMLJC
QcIZdO7KulYm25tKCc6oRr8fZjZKM1f/2ZSvMf4SsJGDy7IuAR0ZKdVarDIbhVtWTHWb3iYFlBFo
jNT6J9oASOQBaZfFkGQP+E6c/sMIsbWjsV+bXwneq/Dq1ttEycHwHZ1TLTlPTMwZKkUWMIvfoVz9
a7BajEEpeuMhAz1iEjM/d+Kcxpx1sDH6Ifa3Y8b5o0a+11Yxa1IwUzQTzSHr+nUJSjgszanxR8FZ
fzBDDKtFhWHtLMnrh4enmn+KUOHr6aAxWiGZuASlO6CYrRT4RN1RTkOGoP6gOLEFehqxTjABXElQ
A5ZXcKMljjy6Rp4JaatKSbhtvqPcM4C5L8RlnYxjZmgSwkDaPXkJde14KQlwMT8fwigTQWdnxg6F
a9r/Mi7jpTCXyPS8cJiBi3bLvwjtQ+UGIk6aMIRsexR/QgAUbjQXy2B46MfgSNqoSj/GNjCYC8Bl
+AqRKE7NEaBS9EtWupQg9VdmTwvrmfFPaUPO3RvBiz+m41secOy+xqDnK/kKKlzelrgr6DlMhCNy
uooq3Libkd4zO44E1Big6FMlJ7WwF1kl8/Hm7bAJtHh+3BvppfLfNLfcDMbfMq5sbFXXkM6nfGEe
EzulTtbywkEiYHvLv1/+xUXvDHtZJbXMN7Q7yERRdXZ3XMKbqk2dLTXnR3O9cFD+7XiUEAiPNn5Q
iCqfvTSEP9l0yZldt2aDTZ3n5d+MVdpSOqky5SBUaRcVPWxuq0dUuPYC/QbD8CHy0fxPHZfNlhw/
GZl+66sp5l5hP62ogVZVcIsIRvyl/KfwsM/Atk0ZE2aulKCB5pe7SgpIxAsw2AGcvCRFaRUNlFo+
DIyyFiLWYUo5kpQsmyM8Zse5PRbG6j4dfWaGajdiSObPpreF2HEa5+kjOgvPHjmw+3j1D39MVvLO
YJ/QvMT2r2eGfEG1lu1Xu1KzG5N+E9FxeDTjXUNpW9xBOa7qiMT+FspjV2d/rwYrOe7h3BFMOnF0
zBJyKDY/IREyUZ4Hm6gENu3IHYXuYJQDSaNEbAzmByBPjCFf2SMHb01rl2KXWEchIUPASP2O0gf1
zvyDNOU8kuP7+f0T80F7hE2gXkWfirToIu9InqG/Wo4yumhCWJCQ0xvb15b8iTvGgAprqX8q/h+4
SS3Y0SF64Yyugm2i+kXpjmdeg5lxVmG/+SxelLWb4Y3N7TOb2BmqdzzehTGqEDXNtQQkbnQdEiqn
To+Cy4l9E0N2UON6sdWYjIW5/E/d6NsjnYIpKqnv+Frt2SQUE5VjkRV4PwDPyh1d8+KDx/+p7Tfq
BX/NGofATy0ZGaJVk3zxoJ+g+11l3rphQDdRubgWrdmL+m3MrkorOEkqjN3wZbEVeFzE7QlOEu6L
jweXADFzO7r0DLyfCcA3GrUxj1G8uFCowM2mLI2TX7elcx/0/6F7ZlVpVm43XSzHzvhK5Rxjcbpm
4BmwiWjuHYkuoieTJwm9MvFNcB+a7xALxGwWQAljylaMfk+B9dgF5gsKcx0Kg6OUHg9RqY2LNiSf
XGrJ+MqwINar+7fIWtu6SBzGSBxrpdlBBqsyafJtarPSufcqZFR5Ep5vQ5x5dtHXRemFNpJ2a2Z4
w9l9wc9UxVuCI/SNE4vu6XUHnBoUvm3VJ3RkH8G+P7l+Ce4xgUSSEFy/fr4UtOL5bBrcJPiV0zew
b5SKVpn8tLnFBOXZTz+RNz9vPep/VjkXUSBzHrsiq9jSnICHCPscvXvar2rYvDzL091qygVQj8P4
IE/R5WXoAwyYN01BbX/p9BJJJyhpR9p1Ne+1Rv//nnycUbMVwjee+x6cn0XB9XdoGQWBHmXoKSvk
Jd8y1BxN4PRCB8N4Gq9YP0lgP9gLkPKOTRfFFKTU0B85Y8Hfi4GmrQouTkuI57dwjdn67xpLrye/
/Wj//prIOJK098JxX0wGG5NOywcUZy/ogjINf/N2Rg2jqa9HKbSsdOKM8hNo99m/VwZG/PnwixnQ
+zSEYDhi1nzKiOam8zuBiwnR5cOemgHXsk3gzQc49nCcDxsFpdZUDUP1q16L1A8wJdn8JHhjrS3g
jZr+jF45zEAKgmyWBZ+NoyaAFu75jcKMQn11ItuV8MzYweGAiO0Szohnw6X5CA5fy+14IvAC1Pv0
vmzZ/P+4mbNbn1yc1nI52l54LtzhGnhdxQo+Z40IOrtn8qjq1OlL/xYDvArGkVG3cVRa7nadgROW
6Ymuu+Bkk8B6O3QLSemz8oc5XxRYcaF7H3IIGw3u0xWeVxcsknKH6dM18M+dc7sZJYXf0OM0qknM
FK/EU6x6dAlH+LMZmqIz1So6LKCh2XF/FLPknoP5rxn6UAh3oo0z9LuhIGOIyO0yUUjsCDSlIezc
zxcZyRg5N6OkPNUBOk+b9cOIRViJI03Fo9AZ6/hTY3RKmsmhqRFcgFdB/gosT5kUd5Y/D80rMW4i
msvH8xSfD9b9a6KEx+3WU6StrZRJttkzH3OlTnnezXiQw50T683SJivnlfJQJ1huxvFwgNXlKnFb
5FZMKZ3KZHE11YX060f6Be8G63e1hYfFc5qAzqCXygNc05npyAna1lR9GcbqU3TvLPXIGWcpctDu
Sui7mUhIx09DEzZ3Se6d/9QAqT4lflbd4lHYHjLgOQyRfeDW32F2tIZut4ew8v9SDJAKK6MlPSQw
CPkOyawvjjBUDhU2QJBH94/+ShdBqWoTbkpJbEXcAR59rvoL2oYN79H2ZjNH2rvGg4HSXDj0bXaz
3B5nf1NUzdQnuvASYdI55ig8h5N4hDrf0Momp0TFOowRHop1a6ktKzakze0TGH0Cy//avd42WUsN
g7fTdrWu1hKUT9fglXeAjgOENpwB6DzVGR/2J4TXzsPmpn2qvk8uAVZEFs+GJBxGV+D3ENCkX6M+
LYbX7hWVpXsA76nTlL7M45TbDsBzMws2AnmtiVRgqNlXfk14sJkOEuTc/lTo4vgjE6wQkzS+QZmO
bCJKfSVloVrqybmlfX3rONjKi0T85cPqdMlCmYM3TJiytbhcE9DkC4+3+gYah4qVJ92jpZGdRfDb
By8poTJ1EsXgAlCvGF0EZlFejlsw/bfQx0bnOZ9VfsyxpRpU54cP/sPRuk1CW0gRaGOTuaLYs3K6
DjQh71m8XpkNkygk7v7YHPpeT/aCeg6izDgwuIYc63vbOx0rj5ad66xKZOfV18ul4aS5pOtPLzgr
LplsEW5W4FYgd4j+/+3UG8CAJUMK91wAIYCdU+lEKLGDwvb5ktdWwisQUd69haXzq2UV4SKw08YY
1y4Dm60FRkj8E3t/3wEwR6WgtRXhuvnAZpkRWwzE1nutz81LgOrF7EL0bpUAZ5dlTffheoOaMgOA
q8jXxMqWjH+FLoLx/VIUILSdF4scJqBfCZNZBMpnzSWY+1KXwcY3jO+Dir/zjrtVmIUGY7mRUNvY
CH1frNFHZt70A+Q4X/OWYxvCYoAAabBzA4v85tMtEtMAUf4clHZyjbcVsdSiR6UQBNVNlSK/zJ3P
R0ruu5V1R7bdgR2PIBMylWb3h6z58Ci2aKdIBYOjT4aMS1UBr0DQRkJgkhWRvqPIwV9z4jMe1psc
aC0/TH242VlvprBKbVERF7sqmgyQpxeynt8np1ZMSUGZn27L6aSxb5+d7+n9i33nhsHrd0lPiOjq
oo9aTTuypOF8IDFvgzoT+vdOIYVHIQMw2LJuI13bu87nGTpLxz1O7tFT0Bcslq+kWmBt6fVR9v1r
QnHHm+wOwjv6XytNacXVf0dhfuaBSYa0FWLPnvbF8/6gkbWLq/85bS/oJtsnQqSJPq5qLKWf78Pn
Z6vz78wXx3k7NVwONa6i5R3Z1HG0n8BgpIFOy+eev+FsMXr+Ssf97qV7a5aLSgF+rkeh15GymEYY
HnUDeKmXJZkW/9eCeHgUMAFReUYrYHuwI2bx2oupF3DOWoVazjNyvFFV8owumc4A1q32NiI2SKQv
d7qGpzsYA644ceW3ojH/kApkdsjVeAACz8IfgMbbLdW9BSyKQ+ACnoKxxvJ/GUPOO/oqxi4aykEj
TowCpPG+EjaqoOKRAAeNg0AAs5BEtB9Ad9VoTa3dTlUxTh9/zKX+N8bTN8dWwN22iXgM3iz8hmg2
IdqgsCvcg2AKuVQJY2D4yrPgbx4tz9cRxF6Kep3MBEQuHgZGqVv3XrstwihFqemCVGXJniNwT5DL
eRq5p8GUhTefkqS4DRgKHJcbirQdRh/7v6wOg4XfJkI/Smg+blTxu9LoAV7uONAbwWiabCk5bSiY
77+rO1ZVXFXX1UV7gM7eZF6j3T7+wyIKGVby1MFfvM8x7MMeBEDQIx5Sv4gNaeYBJI2q1RLbfxFG
wIOCtCx/wLTMbTsPJfYtDsqJ6VGgoY0IXseS9vDZ7SNvU6jo70JwhfWV1YN/7Z0Q7nl7G/HYbvHf
1dxZ8yb4yrVzLOFrqcdB2stu84U7Mz/msflwk4xnfJRP84chzhc2eLcFBTW022HoqsurLmSjAxYG
8SmPLeSxd4P54DFMaeOIQNHyt249p0p4TUJ2uXjnNQf48pSLoHjPEWkJStKsKmclhJOVpIIaNssQ
hAPjO5Xwh1EEPjj94KEf2jRhIOm4SfmktKoQvxggAlTFEE72MYxPe/E7GnVAqlrGTt2bZ7aSpFBF
syQdd8/jc2kZ6v5hPJ0ECpMJvNIa38ggXF5fCOyKwIEFIhY/OTogiQ7QkJM5hkRUKueeFDsRpzhP
l1skPesAI7sjb+o8BdsiCTtUC29f/m1Kwat/KM6wg8eR563EjgpsdjDMWGFWM95c5cpw3iYzHLMn
bmBXUJf51F1etC9nehEMIvHsHbVxwZVVj16PPoWcuQ+S8gD0Ok9qZfJ0RYAeGe4Kdiw1aJGEZ8rx
NPqgay9T099leL22lIZ3vsGpC7tt2I0pVIZGtEy1Jzfg/3MvomfO9njjGj6LOuhBbAEc2aFkNaAV
KQxjRrlwnuyMwt1G1/LoDqqh3CMYExXF895kfHwNRVEFhtMLRNK/ruIwHRPa0M6J0bXtEF3/3O5W
Tp/vLPCN0TAhiqY4gwhu2N9+qHngmaYB/7g/Ojb7BL5JHtpI1mZr6Q/10T/GGkOOKbNaab700+9i
57ltsNSEayO/XpKZLbcaTRgpLXkJYdr6q6GrAkb+ZWsc3Y1PA+Xy0IKdl8HIg+xe/kxuCsyNa+Zp
hsyrjxvqC62IkcqcwQicMExW6KhU8188EL2zpTMWINbJVWA8SdiWqdP4aYEMFcgI7Bf1UDXl6Gkm
T5FGImTeBgpPSB66arIeCA5wEP0NpZQG4ut9zveAdFEeioIa7Le8ECvAer6yvhizRS8uSuqvkeXY
B4z38aPVc7uqp4nYYNgYcFS+OOeg99Er+yimJbSh0WxLmgIqb5cIPHQ4HgQwCPvRBf0SWi6kJ3hv
EJu1MSrzD31cynez4p6cf0P7tTzRjPRcKahBAU8fRqxtEP9jj5cbwNUulDhfEq4rWSYeoPlAilhG
Zr6lBX0Ve9BvXhkVc2iqOtHv+LvTGYJpESuQNauMhlJGSIOKadY4FjQ3iCerInTW9CsMM10s50U+
+29s+bTF57CdYqcpPcUWk97M0FG9NghPK0rwF1UFc6inz6DqmaFhljAgrukFUV9h2PlxGoTTdTrm
TlvRC9G/joSLPtzS7PQxZoETcY7gyO5+MHkjcKpvgk9F5EUFMq3x4TYG7kDlwdDdUzbOgZs1wEmU
J1z91ciwdQlVezImHEjiqg1YDbXoK/XUvupR5cB/lWJ0r1qKOQJAqO6mKagrAS7P6QrG/pAQuT1z
prppiJBjnh+pZpuvdjmTVvA4HbJVtmOHLMrPZpNiyGgAWdh7Rdv3OkLhm5X9/3gbBXZrNBVM6KLF
e8gIU/VBU1NfOupRo/FzCYLTfRjqPYLAaORnWTdTUPz9VtxJOGaGneiOs3HWIboLXN/9KUZs3Kwi
U2O+v6xcX0/Z29WbriMQpoSfxsq22IM5wOyz5iq584SscA0i3l6I0v6OyA4iLdWCtTYNiDHO01ka
+KpkYIOsoeIckJA2mC+N2zUudYVS3/i23w73OG9KaGwGWhVbK38XI+0e5os2Pyu8tkhN27kaRxwy
ylBTVZrQbNfte5H0U44dWQp+EXR5ogfu1aT216qZURRi+MqfTzQ0zwRXqYAUACHoYkb3okdeqbfL
PUjsBOAcJpb1jThHJYTP8r3gKvIkNU9b5Nr2pjUQjUKdyMjKmstPJjtiwxuw3hw5k9nY5JREDHnw
S6P/OHookBMjB/5XOIzGi9cbxw1HandRh5N/lt/Qy7HbNOe8xXIeGLteJ3Ehfi3hrEv5H4HJelMo
Ubf9cJ33MN0SWaB+LUngndEqArxm/ON6oLyTmVjLJtoSA7U/UO82DmN6UmmUJ7H6ZKQqW1jZDrIr
4AchvLyZfL/yy9OkKF3u4W54VjPlSUZ5UKW9VAJMIgJyBjt/HbVmhnSM6rzlV9yVWTjZtSJCxG4+
QqCbnrLJDZHzJxry+MMh4VocKiinVfEFSxubvRnmWfOsK7iplwqNlF3azCyNowET5OcnPNorsEpo
/14aj7/8Od0Zb+noXSpv/P4CgFyU0nQUX30BFiVpd8GOtnij1ebm5axPZWp1Auu6AasuzRxilAzj
iv5a8RkaLgXEDEGm/YsEGctLeE7N7E2BwBuyRgGcHbBbButNtzyvGwKNdrnvWC1yp/w+vU56fe4f
vtBOc3X4/BIjGEkIcmr9Ldo2hXEe+rW0A8W4QtazAwcr5PQEuOg1kS+DEp/EITPwAYD0useBbabA
ZQ5Mr1eljRksm9hQI7Js/c9Hy8dOih0mz5rACKwSLV5TP5DkvR5Z5Lidz9V5DniclIq0P5DP/qGY
DSU50noUzF73zHNeKDsRHJaLMKW4kUdjFknYPdNUKeSNmyf8MbxMF7i0e8sHMAkAyaGi5soYP8SI
0zeAzIwrIyd/T6e7IiJ1tSsiTK0OpwhsoJIjWQiPsl4y/xofsYSma1xn4p+ED95TxxWV1qb7ziKq
llA+W/ZoegkncrS3SxYsb/nuEAjX6eDyOnM5zYJmfAQM/w/Le2afmDAaG7u0ma2eOUsAaVtFX//r
3lPrJwqr5fd/EBALtTEn/3OKkM6+5C2Le+ZAspt6lt/xh3zsnBtitlGscNNi1SdUvIgK2+2C/TLb
b4NtQtyU3M+t1BWzeIRXivv9x/7qAGgWt6BaXkPh+6yreiShYZolPa3rpAZcRY2ah13tjO2tdF0E
LMgcqlbiP5Bp1bqfFpfkcGwWcgw/j2C+hdDExCPGVa4nytFBdQdfBDYM8mqadbWU9DwLg659P9Qw
+35GgwHPueBtdTprpV59EeTltGYXZ5EfR9G7ZeM/fF1BqPiy/4CZgS93S16DQSUFmCakGl+32OfY
yVlGHp+sOyGMc52uonUzRVzRh6g/V/7NNtM1J++CucM6mqai3qERA1AoR03Mw0IHbWCcUhFY80pg
U6Z2AklcfevCcBcLoezPGDcDFqup2cFCslyNwTY4MfdCaJM38LwCqyXdbLgxQXeT60ZjurwiXEHw
FRiuHqdeAIJlmMnB2UJO/Dj1o8wgKHeHwbDM8QyQpcuMgk9Td9pfSSDa/AToGOWdl7v4hr0S/auz
nTqYe4M77DKgWL/VFOSGzeRer6dcw8jHhO88H/+PuxQh6Dv26VGiSQzDl0/JiLq6aLTjcY8fEaWF
wyu3QAQa22vCXgUeJRvWBts8Ei70Fg+rChhAPYCJ0mEqVKfOu3i+gp6hH8+BKL7yHjxpxFzL4/DR
RoUwDjU2765TVOA25wNquxyNS4coHVYVKoYSye+Hd+dI+R8P+yoBsxEdZ0+r945w8HbFx2S/wJ/q
g/TCQHEgLxg0kUUCZH5iYNcw1s0DY3irMbvP9IdSmxT+KDPaQ55BPw6j4nYGwHzRfAtQTKKi8BEU
apoNta22mH/92iPJJmdZeXuRG/vq6LpC8TCqgYUcefvn51ov7UIlgFxqYhJzUPX1E09nNhGi0BlA
k9g70QwHuo2v0xLdWmZy1+U7vHd9rX/qiofKkLwQuGbegewTZyQxni51yrk7Ib/oEeV1D5eePZtF
cgCe3ZMb5V2uN47Mn3wmn+EfYaSb5MwFUT9XUkbwhSItXzc+Kxd8trcndGGR5NYRxi30hbtdrqGH
fBk9mmoU/uxXPITw9wDswIdy5Ee+ArZQAPsVJgGTgK8b0JuKZiRQTZ+v0lbTYh37x2+5EOQkca6e
SyevzXvfgbWqPU/HV9VTgEux3++k8bdKVXpFhSxieDxnQETIgK+WiiF6ksWiVIiYBTwaHeIPE6Nz
OK5BanKczqkCoxlOy8Il5tmEmvBISwOqEpikjSQC6mz1mmTEG/YekmeRo3zr8plgPONN9HNzT0Lj
UEpVCOXiFywRqZ6NeIEc7RILTGxgpAc9yf4VrV36T/ER4ZlDx3xkPmX8WXGPwMmgYO9YlhdlbMyv
gGxNw5zFQ85KEgUYsqMgskoucTwCxjY/b5ZSmvCoHCybngrOrKWVHVDh+HjjxLZRkfVyNdQ2CZKz
Ww1+BETOslSDQXjE+q1nn/8+Z3uI4HqSwwMnJInzJ69CWlNt8nIfgy/SgLa4yTqnb2ryLZKTQw6K
y601bdmkkPO7pSMPOatnDCXWvpciZxQ0zpD+JGLJUjanf8lPYucbPtZlt/hxysSb2ha0QKYVcSpO
3ofWRocT/xCYueLFsQq9kfsShv2X9/jwCGK2rYRagDpxLkK9SdZb/s4bxmdO4g+O9ifLp5SnDt8Q
VzYr5LRRJ3isz24eE6NWwAqgbvThsrfAr/k4MviMmAB0ojVHRw/Fnvcf/+fYY4oohiFUAj4chVDB
Cj+GP8qaJNUBm7tDVulhNp7qPSxakGXHMFd4B8uWe1/dp8csbVGqYGqsRYMBYx9wwW00OHM3P1ye
Fpb66YxcDQXm+bJvH2vgHtGVlHUqZCJs6+B/8fUd2RHwhYOICiDiMguKjraAbeYtfo94oODs0TZ8
fp5E3j5+J/WZAGnUbTO1FcnEUrJUibcnPZ/M8oetKXbaKGQKaBL8YUkcb+6+YgmVsdEwIf04zd5Q
0X/8zUATlttJUFdfh9lJBEGDycp7vK8Pr5kzT7XIvbbqMvTLmDqMmLiDr5o4TcI1WQS9ps6S3PqC
qdvVNs+TwU7SAEC7tKCMwW+57W2/h12ddtJlMilwqVFWe/63fGfIXxBDAqOMObebUHkVBfcuMwWf
/+rFNsazzhJC4zw81dP21Q1oV9A7v5MamtiyVLaOJnovWo3kVwsEvSbQl9tsvVsZ3RcVJVutsqvi
a60ihIEY7BTCQ/RpGJyzx1K+HAXBXAZh6Ze0FwWuFlozWaNIhWsGn07aTCS1+BM7wKOr63pZR5NE
wS2Ge0OaHR5vHXXEeGUgr3J8dkD90sP9KcLkPIqfov77uvaPlVB/bLRTb/2daycgC7gBpgyisdBh
xZtgjBak3SBhOS2O7bOn/GJdrA5ulMFfcE68Ri1CWlnXibf9yvfawrtRgpisYS41YNIjzbLnUW9g
J9eMJabeArpX9Yo5m0rd9ctbIhjgjIQhmNCxyDdlqhtW76OmpDDZw1CVGimaOs/FJY82/dmpMCub
23NE5cmY7GgIhhQVNViIut2Bw8houezQ0btCxNYdaLIDY1wImK/S+J2oFGCJdYgfFIwwXtmUSS9n
5AvzOkVdwi+/89RxedU1O+5fcMSWHrEwqymAxRsUtFM95OTS/A2j7LlO/AO5NQvi+PbIErED/Fgk
4EMfoMPGepgG5N3ryZkrvcyWAskhwNoFIzeMXmhPm3JGWV3RPtuiNNeO6PuzJylDVAkhLipfJyyP
a8HWptzVQvZ4VjRSkSC1MJtliefwsBNCLzbnX5nP8smEvQLfGl0HmelRQ8DhTxijsXy3QHrBOPp1
gObbPTcrMtdf0oE1BgvjLD55pXD1L1c3/wb1ET+opKN3pXgr4aFzGQv7aiyFp+4/an78vniQuzBv
3hGPxX/XRVHcjoXjVVI2oUFsehPFISP6o/nE+GFnEMmqcpO3zscjdFcwmesL5j3Ync1ntcZxU8iU
kkZXFq6QrFdEA1qcK9l8/WasDS57oXxqEECLcVXwzXIV7VJX0a+0TwJviJ1PSwNfC5BlOvGXRf5z
9aj5iq73TEXB/aho2KNNc4uqza4PVjIIssVJ4FwCaKakELdBwFjeUed9bD+7C1PhHOTV0OniVIJp
pNLLfUQnGwouhnztPh+gCdv6czqw8OjjiNJnro0iKa7OIbhXPpNe/MCdoahm/owN779kCWb4ULqC
RrKiTC4Ow34WdEw64OXoJqwstSDXoI87oOwTlBHqd3yQNFsmXzieMJoyVlta6sTjDCyuL9LCPTO8
nTpW9Z1+QBxOeTkZwMx7H916RBeZO4ynZQeq2IFNQLxJrHe0FQngTDDqkx94B0bM9oBfbgRgfibL
QS05iaOUCKAZ0N/wOh//eEs2EYuc975uIm0+d0/onbBjYUjeq03cQV/A2/hSLezPpagCYdtDgmk/
12PDn701PhFroRShtAlhiU9dzHPWBKIIcPIt1hLPJTibNJkQWFlMb4GzNdJpiVhw2aWZz8wRKKDB
EGVuENi6Dsab9iv0Cj8+pC5Icvgvr5xuI/0KfjgCqQfdNpp1nQI0lMpXITZEej92tDkCWJAJobj8
uiEeonlK4W/NwMN4+z6pBZb63EJ5XO7P/8G6Bg0kwWpiKdP5qNlPzdE5HUCasbBHzQCCKh9bcGFA
i8Ko5+7OznyUpo859SDQz4R+x9eEsZXiJ/n84Mw6+dbBSR9kDr+T36svPwjRdB+o8cfByiGxO2oq
v69hOI8qO4I+UCMpFB0EZYkLZci2HCHjP860Wm0Tc1BLez3YQ7029zNKZp5+Yi79HO0EMKHYIP0H
di+UBxx/SsYynkc0VAqpgUWCGCTYBXf9gSndXu3YgTfutB8EjWUk4JGTD+NvQwVJ5EUXlp3/959H
+3Bk8Ae4osD/SlDgObCxELDRGcoigjyjvDGsOmS9Qr/jfIkpAphaUEjFZMJtN5efirlLVF7UfCke
yvTkuz3Juzx0VtqR7t2r8Bd2zNNIcjfzmSw3JL0VVw6qUHlFhVp+jPgSJ2UielkAcsNi98UxTbDa
mlrsC2z07LaWMBpZzKilKKnTOVSM5mSglkgBSd7mrPV6GLdKHq9DF0Zw2N9j5aFJzBMWqMD9KE8/
UncRbscQUZmRCc952HIxHzEGjbDqMm3UMBCah3Hb0xPBx6KcKL7PVv7QXgBd09pu94pS5QJhd/G4
+eVKlO4YmIpdx+wkwZv0GAh3RgQQ6ai3bmDRDuuNb4Egk8XkpQZYHghOvAiTHIJzH7cXyBmQoD+o
X9GRZIc62bRp8LSwtq/HR4oEhSxyv6BeriC2J7zVb3flJoyc7Tlky2U79G6lXIAwpgQjNerUAbCA
qbMQ+zbQB1eBADcv3KaXEfv6o+vecjdjB0FRvMGnqpJg758dGJ6gaMEzUIz9Xry5a30DUeVAXCHZ
SZTruiW8rNCYb+V+yaRQTpeuvLCO9RG18PeHm0S6ThKUiMSKKz5Kva496quasThK6XeCPA5sbytz
ifjHHe9PSqfW832sRnfW3IZZuydC8bf5XcD/gN68Mf2Rdd6FXvvyB84x/gz2IAp2CV4zUSq4Kfkh
cBslgYsLjPyEyog+wonbsPbt1tfXZD+3NFR300hwmNCU0Bn7UbqDNYcZNHcfa5fCs9Mr46Yow2Ar
qSyXf33QYxhC5B3SsNbeYyxYYw2+eiZAdMRhBN0NapZoftan/0vLz8EBTIsvGIta4Jl/gAOQQkWA
cfmIkoQw3cH3B2h8XBqBqAtNlbHHiB3Vv0DEO8cV8cDExjWFivm/U3A7vwh96LaYjT4pV8bmZcMI
0LBZ4WbXYMRN+YgotfC1DQrMFDD8Zywt1RuV7ubXWaWC9eregJyfMrItdaUnM80xEEGBKP5bNdEd
KzuahrYfuMoCfoDfLPqKggfqcDan7s5CqXcGoLtNBcuxzZDFal/8s/MBMqCrHwUClCIA05RTxpAL
1/PyLimGzm7EHeje/9489D83S7nLix4IhcPnY2ue4phU0JA1OGe2hDo3BVKTgX3HypsNpFrYRjNv
BMR+nAQGMVPQ88rGtzhdtAP6Ahh8SCqR34DUmMWAkaTHBsXOo3dSOyndJZOhzxiauSEyF/guOwmX
aSpUjuexCMOuMbgMYt2Pq6hYbekx4YJmmbDEZtNi48qGe4uN8eQJzC/v2VoAR6x9vCnFHSHVMkE5
2l3DQZaL7fHKGCuEokuuYEVjjXyMHIUUArAzk5EhiDRqnJUdxOVFGeQYy99Fn/fEkBH5QW+3pAdW
wZMD+DDOrXSAm3dHmHpI6I9EasLA+h98oJl9nibAmhXv7JqMxne3FOfCPT0DdACKSkp5xpuwklX3
nP8CPhwnHY9/1EKpFYahOrQExPcSN9MvqeYo+5Srd3mi5LBTqYLj47y8ngZ0gZXP7Y+5RzjMs1fH
u37H1HrZVbSCiqnAdIgqLDEf8wAURGkBnaCnoa+32OZp2nijsJekbJeYrJmDaVT/wJamrSqf8QuC
MXJ5zrKQW+UXRggzHPP5TRAOZYhuvNXektCbraEhGArHpFFKH3PXX2YadwBaZdepBcXELjv3kSOO
yciZUNlfUZpU6O2GO4rQLdxtk4Eev9XHtqsrsmTtSJvoW9hq4kWKeflD651KYBq46YD/ABa5X2wu
AhmVHgYAVfK6uR8krrpVFqPurG/P9x2YP4oZ6QhjKhQcNt3m7ejJ0FkcvHY6/Z8bKvM/pDWq9Hh7
75zip2TPOp7JqcaZgcCj4934xuSLfHCHdnAodgkzzpNdlwFxB4CCF32NA2zfWFtfOYIp2Jud+fVY
bjoPF3TimDyvp5fQUQZy6F6kCn+BJkoqEt1+AZaEnjaJegkeyLfvPGmYORH3JMwD35ZLliMPkUKF
z3f7XRJ8ywLtDGNkT4QgVog0w1jX6UKKQVQ60rOHbu10zapvnIItdIFRJkBMn0vWC0k1Y9rGpNaE
AoLIL8M6SEV2uYkYSDK59a6iplxMQzedcA8b5I9R9eJIFthy3PAjdHl5NY0LxU5E3yyPHo4LmPpL
Req9HcnXAC2LquOY4gS8qL+NGvjxkllK1wk+T3KIq2g60KOKHOMz3WpOosXv2YLnk8Zn8ser8dhn
hwHxxr6m+I+0vR0wFuNeanHVU5PxpnMJw2/JoTXPQ3N+RxzowciKKmzSi4MOwVzzkTuY36XWMaUI
EiI0x+qdXjfIVoYXPZmH5Mmb90UzBqRHgzOr/CTLh5fpt6nHnFwLm45N88k6raICzZMieOf0iaA4
AdAdfdEcz4aFjOZ2GS5LWJjOuuZwS6Y7huSMEKPFOZvo6FwE7xkIklQyFIqqRIKJA7KOTD7FbSIb
M6p+xqoNkdwizU2eEM1NDOSUt95IdDw4SoNhgNWaMKhsAqfwjKko7zq19pGtQZeOXCgg+AwwvAIV
A5GLeFKPrP7YleNZlheI/VIxK3HDWDhG/f2ZZiBkXQGePrFa6++evF+PT+mG/8PBEfc6u8E86z4m
xUvKqzK7wUW4yf9BPbw6g5pstx2jmXAhz+eGikgZL30ECWKOf4e6nGzvC6xkTGF2Z09HSrmhIYIL
tT++wCP+OFP9Pohu/1/9i7cREPiJ+6ZjTj2D/gonfFXyHNEGpgWVxjuxvwAI7RVe8DYmc9ngk/ad
UA2V5VbuDXXAgbAs7G6xgI1suli8pE4MCshlelrfViskIYZW+0+jcuf4Mb8nDkM+CABxngrpXu+B
soxWSpZ050Rb9G8pvPeGFSUU3aHN130Q9tx5MArV8hZyPmE2ZcXzILapmhwd7nihDa1QeQV0yqYL
QIpVOh8bGN8y8BB2SzS0aeHGkjAxsqnD1jylxioP6FQuSuYPCaouXfsDj0mCBaB2s2bMCmHsQw6L
y3FJxEFNJZrLxXg9go6IcUnUp885itsVeK8DTtRoYdAMxHDRzHQmblsiv2hHuAC0HEIcp+zCgII1
ZDMK5La/dpFcc31dy98rfJ6VOuhGG686Ay3hJoJRb3LLTkLbWfWeE3fNMUrp6omVxqazS6FUasY0
WMUVAXKEZnudco3bOTsTdWXnd6qYmTOxHXG9J8F4jadU1KeZ9lKZ4eTMXQfalfD4B0gAEiH61uFg
UahWT8bi0kZOjgXgO19ChgWR4Yp8Oxxm7MovKQOT1bNk+Yzg3hrznHlTZav621dfP94a5tHwJxq5
+He/uRdeV9Erv141CiP0cU2hK9u2GXiKF1DXZbJH3IjS4ZzMDMCZ9RxaqZ+hvfEGY4BAtakmphda
Rwc+i8FfP2fed7oHPvvwTtZNeoDBEEqleRIaC40IGe7NlWkS/hJCgJq7dYozIEdKtjHun6tYpGOr
/0/KqvsVpHDyuPy5sW5c6YqLnett9LfO2fuV+MIeLgG4HFXXiVNOOF8dn8tZExqjmrkgL1y6Yiwd
D13ljODS84g2pjZHpgDolsdW5dGkiFzIrBIv1d3RbrqcRvh88aJ6ouF/jkNcKh/BOx4dfRK4Tlup
ppRQJKfFUwfaLMd4pRyvHhsyswgSR2T729cZt6ziEflm8snrbD8YaFNnWQgCAL0rXRACtyToszp4
7e7E1eFPXpfunOBsZdzCqwRP3OdqZ0Dke6WNn0f5P6whu0UsWO/AKLeZi51LAGAbB47ibzpWKRVk
2zRRu5tn/Oy0XQjranqGX7OIBmRC2bKv+O783cAZWxgDEPKg73JIQC0NzOOLhWRNqPi0er/aaOTl
ZAGJz2mdfWamtfraz9vj2z22GiYD7CUu4PeXcsbVnpejKG6RucUvkgbDK8rjXkzO7zmnabwBbGJq
1+Xj5nUozpmrgJ/spq7p1XXKcaEmpryDeHoLWdfbOnB8C7Pc1G+j367EzRmJPlyqhw0lSZL1kr8e
XtOJ4ULWEKR0eUuYv+xF3EkSkBT7kciinmUAyzFrpfsBt/iDiAime5Sh4LbEOM19i+J21kN8WrTs
8lkLajITOybwd2HjPaDQIPtyf+CpqVpDce+o+xaC9ZXW2BKRxIMS5Zmtk7484eUFgeQfdHjtTriZ
XnBWEHMjQLNSrSNBtAInL3ITVv8a0u67UBDE+XBYB5+MidRxAw8TLkQU4yaMRfXHWZTTpDns5YE0
Xl0yzj5dnkfrjv12gEoVUD0UbGuCFr8CAA6mkuhPEnXCCVXnsbUhvJjLnRiuhdJTuxNqkWx5BbH3
YC2XXNsWptFA4Xznh98HUjkUkCZn3cC8cilPI23dK3yh2C5V/VJVCLhFEq4CeafEHJTexHOoWEa4
/mvgDZnevMnBh89OktOLunWavvbK//uh4k7AHdn7JonKQu58cgrZcnj7e2gL6pK8n8VR3hSp1npV
hmY1m4SwZoOfKrIANoQgSfHY/Eysxje9Jszkgh4jX1J2mOfEXfyeJxSGXgrrzUxzntFUhyTcYgO8
gdJW6KMKgd10zXPW6C4jn2g601d4jrA9Pr18NJOTcNfmTtdgdqf96cYhdeCKchMnGBWJGMSXYIq6
sKtlbloJwFKBX6uelpQs4nAXkcMXW+qvIKe1+ZIzNm7QTG5QRjEnTf98vQ1N6qK/3KOzYTZpXboJ
zJa32sohgZH2Dg5VHCRDENdf36lwGZMN1GpH1Gdw5wmt759nWSLYtbFsCJSm+D8QbrRw4i8YzLzN
zyi6mJpqv4EB23udd7+Cg8Deh2n4eyaj73A8tyQKNDPzjcRkhD4iVi+8ppfTGlZjIG5FQOZfaz1u
n16UjNj2ig1ixpi8Yb1oYSKMNnmreiAEJ+RIEhMF/7yJc0D+ziumYGMd5ou/TP2h6R5axVeQ4S+d
e8Rj+D9Ef6zFh0Bg6oEzE6bzvURmoKOWKGxWJfv8liviRi1iscBTjFJvAISH6Zpxsx1nJ0kzZCbd
X87dqe1fi137QFYl2v51g2LoqlBlvQnZ20AwfReDwfc4nK4SaGMw3cP5KweJw19dOjMBXiyXyT7U
E+rMXJ3Jx7FN4ybgbGtkLCnXQDWtNNj9+6BJh0LJIITj4eGGvkqoczqeVIf1nOCmrk6j0VjQS0Em
5XNoC73WNRuZDTuOaB2FjAcYzz2ZC6laZ895fwt9susnCGxxhlM87mTRB4wbEpQKHGRWDjhFbunA
isu5iP5si94kyEmGE+OtclKp2+gdGrdkipxdVSPd50UXXV8a8ew/35DkceebIQhDDpt0rbv6OUXn
7mnUjp90fJFKnEF6F6BorkHwavfchONp7vzwq8TFBMnYUGkv1va62aLwLizuchjLY56tlYvpM332
V+WuQM2+b7k7gEnm+ODcSCK0raxNrR93jtjUhjY4gxDyc8df6Esx2XQRSDW4fK54pVAH6MNT4dfh
xK9u0Dfdo2hAKu3M0N6/lKYFF/kC2WKqhwPitifGp3X+J/inu8AgHT5F39JxXsW4BdLvdvgDAXeJ
5KHXI7hHRIOJPSN6HIf959YDdRgVMFkDQaPNKCPYQWtmG2hn8xHZrJCPWI7BAk8a5oWVHZb+jB2G
luuRrsiUxtNroysztdqWzApFyFF9STbbOseuFxO0r0e/4Oib/jnexwpkEPemreJiVZTGQQfubBCI
ETZqOlMpoa7yhTJHeOaGmFg04GwDCYG0SPDNr6xq9qaTj0+qsVLaHBVFK9r2j9/Y34qryIXAwUEp
2G5gZMxMKyHzgZJ6JcK44e5HVSc4tGtJ4Ma2pAxjTkk5LtSMC0UIobLykjvClt7OlundpO18L9Ag
F9WEJOhRoEalzEB0ZQPijgPFOZLNQayI456CmaiEfcZ6NBF4pkcHrRG5eyzxmq8GmrQxJMBG3GAR
1oYjkSVhEkMm+GnoH4YxZIe2YA1OrtL6I5scDfN5IZvM8mNVaboVhltUnz7XqB5O9nF6Zsu1R5R5
QJHQUFPev6+BnKizK37bn/C5FxDHTLxyN7jUTpLmCj5i/Bvm5iVr1inntLG6GI9Fqpys4RGFGhll
mTHJNCyZcTJYAxKeZKhvWImywgnti3CI5ZttQqraubSb+ndNrb4jG4JLaiaSlPoPV90fkIl8ANOL
ot2LNqiMYIRsg5KxpMfgL0cWzYf23Ru5KWDtZPr9vBzn8rkdsoKDj5W1AErVKjcSVe4B/nfukAw2
qma3IXUmmdv5K5wpX/YbJdIeGXWkcuJi92PQZbSdgIiyn4pKqqTj6pwntLzFdCPqIHQvbTjujwTZ
z5pBJcBDhwXn/YtRRvAaoNVdimRKzM1HvMB2wRXLVeVA+2avbZcNU1DslIdA0c8a78b2LZ+fqm/r
57Rm78JmwEzNmRvcCIR6dfE/zdV5XkaE9GqAtpobVxpRBneD1kdiOGQh8FLHCYlWX1KbQhZumHt4
sxvOPza8n5c+qmD1Ih0yoyKgAUlEHhjgLmQPAR3ADuQzIH/FAS5XmXied++eozWWKNav4iu+TDXk
cBpTpJDZELCYZRZFzDhD9ydG+qVDYt+gv47CI3jHOwsr/QDD4VNHM4FPIpBA7BEBJOF+8dbFnBzJ
5CJVvYiJfRMWwLGzmMZ1w3sOHs4yRSOCC3Kxv2DTR5lqRXLVCg96b99l82DMa55ZR18v5IAduLOR
OdmOpkYOtPfvVkJFnPwIwRgImyhsUxjyIvu4DIyMjpomaPlUbbiSnN86yBLpF9lMWIN01e7/pPLT
H/W3n2lmrNMhVuchaYtRYBsNHqecdz0mC5e6uJ1aWSFaiQmY49krgbl7buh10wacGXZ0RTE40QBM
HHCfrYrb7EonfF5PD5yOk6XWxO11dfJ640XYAXRYOQ3hqyJtl/R2Vy0EWUGg5z2vChSlpj9inFRJ
gDh5QDcugdyiVbz0ZDZgr4TTszGVo1I3yBG2C7lAvbq/eaFD4kxX7jwhpkFgPacn8fjNfK3YR0Hz
ysX98eB8q9v0JgPvkAA/6rCwzb5Q+7Xf1jJJmXz4gZtM9k6UstEMx33vIrDNQMUUGLeGfwAEuFWN
UfZ27DnqGOvisvrBSP11KBr5WIwknhyXb0+Du/6ODmN/Uyf8SDHVzemEHSaXgpH1oXT1xPyD/iTG
pXgJ0feKfBn1tHDSo8ePvvm5atawUxEo5T6FEhnBfS9YFRTI3uOA6LlybHOgKo+Dgvljt8FdZ65X
Ni2u0RtZx4OLfa6RhvkPkv34FEO4ifoEDRkW+KnoV+NtkRz85D3ZYw/rIuriwCbdutAOrZ3BkfIQ
4OviS6gVuTO8J+Pfby8oL3OBtk0CEvYI4KKBThBDUg56g1hGt+7XHGIz+e2AabYa8o2i+N3mZZxI
0QPInkzVHj+m+JKrhlSPlWp2QCBdp/ffXXokeDFyC7eoHsgM4YnTE8A3zQPuvgZL4q9IOCPpeY+t
87YzJDh2xCkz8EfYurhuhrQderofgFyB66C/5tC7LZWlIkbqaFNvcChmIX2Lb6hHlRGu+XJzhHIR
YouWr1Z3rQPRxfvIOYjHGM+JBWh/IaXVZm7a+Vdsy+uL3hijBKUT6XwpqQpj5kbCU484txQM4I2a
vVVs/sDuo5usDjPRso0IocwDlNJWa8RLIhEb9aw+uZxz50EaGRN9PiChLA3wrqd7Jo5WZpAP3nhW
2Uoso/KL1vE1EnXDOMCIcNcB6k8Jxac2V/KvVOkAjd73ZwrZ0J35+1n8bhHJ47W23ResbvLJLQc2
nvbT4uU0PMKHdmrjjpN79Bhb3QyqKlSTwOR/qyLvozw7l52xUIR/iXUbpIHQEZ2BXsgx8b4bh9WJ
jnq080IaTt0Q2UzhWdnmkV17zFVn+71kf10CUjke6cLvHLZPMbOEZms8ok6b8psRgxWE2485JOiP
vdUJHQjCbr4SBU49VmFzJxQN2VOyNaaeUOAB48DAe/xzjfU1mEn1isCEwiWi3tDH2UwtvONAfCVs
QQaRYMOJtGYTcE7gmWV3mA3O1WhSke5bSBRjYRdLdywhCOxzjsQYIbDKYPcnSGqIELLuglxfACmB
oL18FsZN65kEQKFXLWxLJMcC9ZVGowvxQpn4AaiKtyyQOJwLgDkFlR1GeLeSHrK5XtPv0iSLFWVW
jq5mhIeWhDt+oJx4a1ZbpqCXEHBEFPK/0Y3fQ2fbTgKW5pCa7qPePmJ+NoJK3YYez4xKXuPqXzeG
7Yv4MlkhYEtn65wbaF7lVPcF1NeNV93ckEIVfqEcjDADVKRVYXf8PaG3pBY1pqy7FBfqKHAbmupg
NwplPjGJTUeIXpf7rBl4nL44dqX0A4YiAHeviPRUFCrElCm/+s6nhvATPycytn/E74oiyN+r9uaE
LUZe6EchNfRn13YfE95hp/eXkoojueH1ZuyFLTrgaCrhJ/LXgMUNtAoK4ye1zw0nd/O1BtJgwDWu
ziNPxhmW5zVz2/EzSfHbaO2HfkKjatd+fq2SPGtOC4LjaHOWuVxbKu8iboAv1POo2eiCC6CtEFiE
EDC5CZ/kvNqmQ7izKTWWK36Z+hOkk+1TeHTrbJxb27fD6C/reH5B1uh2xEnOUmW5+jW1xWqdlxVA
sh4plpbHAZcd6AXOP9Tx74iE6FPfefH/T8JIOyW9mHOvTGosBONg0hE5G2csJ8B3l/vfBvFeqiGe
WKF4UBAwU4Deiqqtg6EgO8VNtWB6UtaYgeMdyLAjREaFFBAZ2B/0jxiiF8zkp75iVbc0hs2H9mH0
h8uFBaPh1VtKziIvqo5wrXV5j5R5q0XRlYr+8X/iHC8Kvz2Y3Z6VrXvdb18vm195aMGQrpgreVae
XxpMp1cjATa6WyKhEVxeNQ5hMguTA8s6PFoMaJKkpqpzH0qW/7fLYJenQvmnl7riVaaS/dbfW3of
WvFkir3RnXvCwab0aLKzJThaddl1bCbCXeim/Apji+3h2pkXlRcGk5bFYuTZeamlb5xlJNHCTg2C
6O7JNKpG3DDj3w5a1fnq+jszVUhTmJrNSZo/B7zsF/uInIKUpg/UdWxjBQRoWeo0RzBjHrLcq2Z+
MJbCWbTZMZU8aEVS2i4smwdJEYoUF5LxYIeQ0mcUlIpgBubIDzJQ0IOcgI5f15piDntWU+UxOYTl
LjlIMmjo8QdeBO23ETJDDlRMe2dFWHKM33qZXjUKFH7AVdpMhiQn0S9TlsmqU+HGPCHxz1CxMaMp
HBbVPvOBvMbGVljftWIbCev0Wfxu72MMM4ivQrKHiJxrJgUjUdjGbiVKpio6KsGFWBfroYRAs+Rk
zlSR/FyFn9+StZayNpQA/yJgVQIAm7/TAkt0emvv+yOP4KWvSaVa++LPKr0EicHG6rTFsRdVTXgG
Wqg0EPXAiWFx1Q6tnvdmAYQ2C4JYCvHSSqc2hMMpIusv1gYG/YAll6m6lYZPjSHu2wjaOmxEudMN
gWaiCqfwaSxEZdIBk6xd+oXdYm676BsEiBgf/+EY7ezSDcp9fmqocasf7NY8FG7BBTe4/5445DOR
AvxXJOs8OzD2rqjF4skwQxME/frUAidkar0dIu5mJC9jU8J7Y0NsuSPir0b89qCMh8Kb/lMwwTEp
CxpuUbScFbxpFc99ls9zTRS880o0Qd649he0GDeAxkJik2v85KV5PwIXsce3gMBkaDaxwSVkJE5d
Swz6gYJc0tndZh1YlCSYXN9yhIfeA5V31oDrlVZYP0J3pR39mOsnXV/8fq9EsLbBlUoF+Mus+/u4
MxRr6qEspHFJBvMupgKSQv0/FG0SlW9NPzvNXagX13dCaZPqevIHl9VdzvJEY62PwLpfl8eyEC/Q
33G7VfK1YRzfGB10qL7T144nnN3sF0h20XdKB09yIS8ZXNPlYha8/2LSVWV3x6ufUhzTAj0Ix81m
OB3ct/1TJNhVv5n2eSOa62gxgRviuBqvCIOyhHwsNBil8kSI3274gN+Zoyddk8n2G/vziAJekejU
2OeM/pp+Sm6cwQTCWCXFdlKvURA+F4AIju+UVGMmvYrpCAcNUUxMRvZypsPdgwfLO6xuBF6cYjtg
trhniNkIcgsU8plGZKJoufCyCUYSJ4r9dF4TtQxXZlFldFVv5ItghdikF3dP/T9dxSg1ES1wgdO/
TOK2a8eC+iUVRomJNNCPMw7nuROTes0Z9NKbey3Z4FNINI5H3bknqcXUpYVL57BVMfaEAvARX85R
DF/h1Bwra38EzjahgV1vK6cZSoFLuhgtftINiVPH3jXI3vml6Kqzy8CgyJnEM0I/r3IBWwuKbffL
DjTbc/1+WYXNY1I7qXLvvMr3G5CMo/15eNfUU8DWoxFuOdQ19PJcNMzIYNDHhjVTXeSucmgAmbY1
rFWH8RXyQmPUAGd/ghLQ+JCvy/Ly95fT0HID8ebeth3rGO85fhE2Ha4Dhnskd7J8o6XgA7eFaKwv
Br0lZ/eIQW7xEM1+43nJJEQxKYrO68DumjG8auKSmQ7FmWZ7d5f1UTcz2QvNcBrH2wzVccsQviFH
0OkW/1felbiIkUEs7IODCAGN5nOoqhD2z8AfbPl+DpxGKwNQ1RlNJiDXdPYxVerJhRjQAtIFPKa7
1YUcL1K81m4He+5CL3fJA6KZIumwoVycAcHbAzdf3dTtSaqBz7QVZ3XAziSKX+lEih/ZyfeGXPpG
Ip2maArJXP0Bl9U9lRIl+uK9ran3VW7DeQ57CvrQAMNLO0IXfxhfM8EUKh3Zm4tTjYp32sYHejmJ
sdiEfPeVtii8w2K0XoAbuTDIVjUmpxmd1tZ00FNrNVQQPwOzjQEeHXEsBBg1NuoMlUrNbSNg8qHN
tmr+CQH5UBzoKcvH4W6+ypQQ04jzkqFOOAgMRJhfzkbtbFrX5uPgkBRPfrwhDBf/ZGJbcQwsclQ6
yIiQOG3fXAmWYTxQQJYV1kAzfahRVm3IWcTHV4gVeJ0CZQjdh3XyHJxpoBBiuNECwWpZFhqH8tbU
9uc7OwgBvemjrSX+n8c9WS64ypyx6YtIn4zP+eKSH6Ga9GoR7OBLTvq469PPmCIAxoTt9iLOsJyP
930eB5o2YZ0zpn8JVGfGiISSbN2/K782JBM+liv+NIuoIrwzbQ1d0MQQ1+qAV2xy4BnCaeIiVnES
qRuw6jGKthqhDBpTGBbCmOuSKmymatfCSA+yNmP6KKOFzQdctenc5Hpw/AX/NjV6Pj//bm9JvrUx
lhjTvxWzYnvzx9EmgVghMcsGHpW8SrsJJjVLKbpfIK/j+HjZOeK+pSa9XI+s+5KeqYzc6+uVyuKP
LVTNnwKuYopfgJvT0aX1N9Pob88R+CFUrQgumKI3uAZCQlssPcgdmkZqQy++iQo7AZUFkAXWwbVs
DYjaVd4xnPPqpSoe6DEoz3OJ77iwzYY7coazyjK/8I8oZR7AIYeBOyzQ7bZA+rmYBUbdISWedTWF
YmV2/2eGRXARw2el2vFPKjyOI2Wp4IFY+tFQilZ+jaClgoyiB8lA90Qfn/tKGoIigFlHlmQFzIpq
UQlpr5XgYys3F27cHbA68Rw8e1tGOQrVhvKlffTE2S0KgUwsiB5JgENmyI0sztTgIKBXa01eOD/2
h7IU7wIq3xZHsnm8eINR+K5qco4L3AuZY+qSlhAbW4sw7F3Y+8KXKQXf2dgttaFRRnEClhsGt+ut
53dXioKAiFvVFsW7VlUt3tMGQizgBTv+5YMXc+dbpe2aSuBQRcZrUsvlxhNUX1etIWgVLPEU4Xd1
M0QQ9RCA4+QOF6ca75qCR9ZRmaLwdSdibI/fWONu/KBvlSHNj16MAVMVweHdVRavbYdMhuOgzHnw
i9EC+zyqBm/9wBPHwc7nSqa1SmnYFBeor5eDN24DGbaauVoVCVy76wU6/vk9BQ0j6ZgqzzTrv9ET
xCxXkNV1P9RsnPhL0vO303CZZHXjsKu7zbwDYuhLgDwPnqPcyUkLhtQVQimNylxqbSXUk+9eslvk
Tj6JrKjYoFKIJhkM5965FKrDDhw7ai4WnJG1SdWIQKVTDDMy8QbtiLSk+D8TKvTLACMJSjSelW1Q
wosP40dSggYWa8ibJpQLBQy5nLQ3Mg8j7LogcSU6JK/POei7Jt+xlBKsa0nwN8Vl6xqzI3EIo+mE
6qUerkLBL4ZTAZIGuRAkDY2LvQt4vK061L48VeJLs6ZifAohdAc6XVOBYr2/RpHapKQvBG5uMCXN
klFBzg+yQLIMVdZM7QXTqmHSbPFolovNs7FG7WEKekEOMX7+P8JzgzU9krIhn14JJVUonyXobFe2
iLW1xwsrCAQ8h2YnJ5QyuWAjKxfzL9ayKS6sdT0z7mQLMIix1LSiUAhtgz/QfFRvcKCjIZf9WQAB
/cHdKPEpwwRYUu6L6Xu10gkMHFnyEeKPG3TVZmDVRHVJEOA4F2ZRX4lE36+LBm3+ud5CC+b4Rgus
iTVI3RkAEdtLmm90FrQuC6FJQg445Sk87mhoiE13Z2vGueUgQCe/OEvfmOGBwnFLwIwtLCafQIcw
t76zlT0bIuqhNyAT4/D4kvljfSJoVf8068IAEeZkchtKLC8G+/685+P8yd6wE98i7n+UVpXvQR7f
lfVT/Rn4blkhZtF2Qe7WwB+Azh9ZAWI2q/zBseYjXVx7mw1D3ztZ11IbQ/90BkU9jbt9EvODfIGR
mxofx7jAvVn1I8Yg/SXiidyS3D45C2tx+IOcVaD5K7hNtgfPccsXqgj/sITmXLSvpAp/OfL3wBMw
PwuTJS02Fa2eXHupq+ngGt34rmMElUjarjYUNdWQrCv6qYno242LGf7RrJ1BHayGMY+XthYy0ctM
I/GQ1DQDB3X7sT9QnZcXZtj6Fkyd0JOP2Q3zCvdW10Ku3y/eYD7tMdbMJUGb/Bh93a0AaLM+uyEQ
uAa0mwe+lcJEgBTxWqsuUowbsR0eEidg0NhLomEZxg435BQW3FHLs79lHgnbgv0QeKSMMetEPdU9
w4F/G+eBFwwGGnureXjYE949wWhGIIP52haPulu6XRBvzjU1Ho/qkXjrrl19vZkL1+TdMmUQ3OIp
UR4kFJzZW+RWJTizTTLSWGwcwNMvAf2cSpharfJoA/VpPAnAnCnZ6L/dACq6aKeZtCFVGWqT0kbm
ldP9on4uVB05wBILMP8cthTAgX1aYrR/3lFcGp5O2LkwfJwu5tAjpcLKndFai2p3U4jLKTivYEDw
WJV1uiDuX05RIGH5wHISxuTFwJfKdoX88Jip+syQJdpbw3tS+VUKwd/F9sDBXz1nhxKpDuO76zOy
OqwS1pRNdWaooiuKdIBzDbTcof9SnH7CHxc2fX3HnM1sOQH8QyuoM2TpV4Oyg68F/HX80XzO/5HQ
WGxkfZmK38MYgbG98xKhn2ZOxFZvJpG1cGi77Phnst1w5/GCd+gLxyuL/Xj1UqAce64ESIFtpj+P
/Gr1uI/Na3M5yYAwbLVB0RF3ekqCYMkQtDBI1VE34Zf4tU/08Gr3RsgxIqEAUCwmeWqyuEIy/R0N
lvNydtKBQSDRtBCXR/zVWlR50mroeLo5enCIc5WMs4EZh9z5YHIPDeVfDjcfx2E/t+QUQaSGUgbG
c+6x/SWe+NEwr4kBS+anKGHGAWRKaFdIsgT7F1csTbFOfoeSdFQJbhMraXxL5Etwo3Zh3MOnt7QF
w0350kLOIJNVqEUPaMRVWwwOu8BMwdGqfuoKKsNu/9iI62wkfAWIn1WJKmBShZu0A3+hUa9/b1py
RmKKwRpOOhXYrt9Vb0FBP5Y7cyw+zsNS3hRMNgFVqzZVKf28dCmjOTqH1vw8MK89HgpuA+t01M5c
hHVSv4dOKDEXgYJByDuCKWqd7cQjtwPURo4n5xim8apFpn2h5Tp8jDvxiSFGhKAZITeKT8dARt+n
IkFGzdpJ79IBiHblRnb8yIJspfS8VmlI9JuuGFcB5Oe9svkoQDm7dWRvDF9noZcUcniU1X2Hy3NA
UEuL9F/DLJieG02zkE5xqGsR62mWXwv7u+QhfKY+p9sN8uYzne5GTs1/+E4D5N0gJHkdQuobCgDf
AJkA8HFYV/HgA7Co+wr+Bmb0mIgoTHw9XQLiIAFCifYHuOcSbzBIfbfAmZfpUusWDKC+plKup3QW
uPwlYv9Mgs7/6j5j6PP6wjiwtWlJxsMJH3oyRhEcR9zFJk233vrx8vjpgy6az2nftMz1eaLCHGo+
JT7Lg64tthpeGYjSzwRWszAWU33hAXNHJ9j+n3rbtUoXaSIwfiqI0TfPeTG7lnmSsC8cj+Njyusn
Gb0qpwxQm1goLMI/wotv/zzS4v+GFmcDZrsFzJRbwNjrlT31dApNXLbb0NC+LfliNdHE83LDeJbE
HeyOS4Zhv+uHGQWcTIexTcwH69wWt9kZXZbUf8KZ7EnqSIvehgRY+Cx5O4Ri3V0eB4M2AJPw/Dky
BiVos3IwjEtU+lqbEokbu6LNoejxgblLISNLUNeK1l9H3yBFZJEXVQHl9DsaJMdenEGUTPHdTjn2
Aj8hXRDLxp5WkrU+iOWPPDqePVpInG9LbEV/nw+GsLq309Oj2ZPxIcPJjhdJHUA+Tgiu5rYKTsdV
DuBrRgg7hSuIfAWJIxSGVKp0xn+RIsd0oBgTViZSzM1MxSKZDvwfzjE+0Txt5r4TWu9SDnjYPc+1
KOAXltCEQmyf/4t7xqQvQovJwYgVVyNTnpw35Sfx9Vw6uBQH/cKv4RqrIZGrBccopQg5r0NgzjxG
HZrb2THV7aqWmBmGYKlr+KXnkxUAxmq785AoqeybYuQWPI+bzBkP6WufstQfXkdCiI+xQu0bUScy
ayqUvBjHr4vVX3quvGHxCWlGA3Zkarmb7g/rHTSepkR+JczgLZLU80rXfsTRlSB1IgKbG+/E7xez
LZOHdtSMlomPg3GLgkwjJbNicGPHiDZV1eCkpYsb0aHbDZUfOdXE4hWHWshrlWI1TekuHRKRJxLN
YYabBqul1I2cGF2NHmV986VakRDRiqeibW5Io3s8EE+S4bN3NmKaRuGHhQh3uckVUgs56ZXKio+/
1Cn/iJWR1tLvDcwzKFs4IIEllgumqV5h6j/gbAodwLA1Uc6BwYjKtUTkYYh/Ym5Nvc/JVritHi1s
yBS7+kw69BWAuzq6+vVX3IGbNWghPbvfnDv8R+PHQ0cduFIjzV24Hp4+q1DUqUVc6SrjYJTeBzZI
OnVWqHjlv7p5EhLT/XY93ujmsp+uIXn8mYykDBOkdx68Jf9hOgovMksQJdI0cIqiJdUglVk/gzur
YoyZplzblH+2MvQCUMwzfhB8nFsgSPbJxTa4Iox+pKo6W0BhpXo1/66FRWnZOjfCO2tV+OhrlgeB
t/25xyiE7kc2oot3sDAMYEupDF4/zR3TxyX2ibGWHg8hf+v6pINdA0db2eHpp2JxdVTQLGNnvKSx
tDTRTburU+EdgBGpxt2E3ckP/qf2KiYtHFEdsH4YsN2sWA95U0LBN7+DufSMmR5HwLvz7hPeXSqi
7XeGKxFJFxcHa+VFrd3aAREDRn8Cg5GXV0XT5BXABlU/Z8xVnQVlSgH2/fvxptxDA0A6JPCi0eNp
7EvOMJyiNIO2RMT4+uOnMSgk+bnKRhGkVwVcRIvv6dmPOIg4UkZ8GxPFSyBD2w4Mc90ZF/sofZnC
k+m9IKgzLcmytYEnefPprXGnwA3ZL6BUbggkPaV6uNTsM2TkBccvFHRu1n/chOT72Q9vCK497YD/
dpjL7EOzxpHQA/9tl3UVIG2lSnyRzNVLT3/vY+A4AAsIKF0WXiIiwSswVrSpx8ocNApFSCKeGGLa
a8nX2EDUdNYvfju1vbuPPqFkhE4JEOclmHu2swD1lPxVNz6lfVN+fehp3fDxhteqKhxJN8+gK3PT
9mlXkTdFrRLjgZrKtZsTuiju071SvHPR0W8A1GH2P5/L9Sa++bolAWGkCP6X9CrHT3UImDarBH9s
oKGnzNSuCBTWKovU8EeorHjnRHChB2UqKtPO0WCvDwzbAS20+wLyE0bHXx6W05RrNICrxYWIcfga
0NHd/POlr31k4Sq5zHYdtXCqqCC+UumPT3gJ6RIsNAfCc8N7eWF5U5rg1pVxLkHhBfw/ccHFLjKD
zGFp6NxpnALMPSImX3Sqz+cX3G0AmXRO8BNYCUKntmIlXvKy8B3hC/PbBjBalZUa6rpXOzgQYn8f
IO9TC+GlPX3WS9cLEDuN8Bo1osThQ8Aa5OIHFkRmLMO/xA9XxEO8bGCaDEHY5qFOIU8keNdpiFy/
4dSZkWS5kHPGNTmoTcgX/thw3ODY9Y6Apwj3CYx9ts1dp1xY3MqJWO3GF/HKL7luyTnTgvduOYuE
tQem22SSZEtv5oDCpA5cXRK5p1TFSyLh8xDeePVCQo9lcIl1JGwDYgIng/6Oq6BSJ3mM3a/aQE9s
rkFGl6Xp3SMJHbhO/lgm2vz5f4r41LovqNcDgr5vRWGvFJNN6AxpJAECOSW/jOvBmzJpLU52W7nP
B3YtPZE1+C426OF1KFOcDzbkRyoDr05SX9P7muHHFW0hgsmf61M0EiG/a22zfyLHe+vxU5R8p90X
XXyRLVEAgzfwBFnY/X1bCdLzIKocRA4sGE+r6NE+CzhuxcGHAPnccDTPFJeXdAkIhMl2fd3R2VnB
njZj6MNKj5VXAvPzOohuBtk/SHbEHx5qZOnsYTQSaxrBrl68xsufCZ+HgaD/0QoQH05aQAv0bCYh
4LS68Zdv/wtmu+Je0OaTw2cNwGprj8smclhoX6V/9QXLtdymmoXJQC+f+hyJx57l++viTSqYT0G5
XqSX/mplVNDf2zt57/z6PH8zwWIn4Z+7tW7ET/wuPasci9TDRDTnPzKVgd+jeyK4iNX98NJZUxAy
3RM45NbhxkPCzYN/v0N4dwK+W6rnTJ5LPVxE3SB0dEeCxF5br0ySkqYxGi6pw3LrlS8FGxsGlEmP
4M6vkfEG5YYsp49N2Jii+ha31OkGy9xvv47/+Rr2rRQGOo2uka/ovvWs0wZwE7aBe7fv16ERydSA
jNhxqSyzrgXLM1CcwkfTwgeDximM7ueFoFknAUadUJUB24+Xmromh+eIlJpAaKeS9Xf/1YayrLhC
aVbYNtoEU8uEAJWb/qkIGC96ZYaMF543aMQdiD73WoyY1BXRWtZ0Gh/sPwi+zhCFMRQ7iSZHjlAc
lSFy/KUNcQE2ij+XAL55sI/S1SHTXeDOPI787TT3sQLHc1e6S+S1slXgDhd8X62K0HglDcUVHpXs
VE/BkrXaOg0ZfQsw+g3jF8Tde4mgGtUOYO7I1rh85HhRlQFv2XgHFPR5RWbvIFqQa3AqhzN1Zx0E
Jj24thPFqwnwmYv0oXkwb2VuDNK6o0KRC+xJzz1r9w7knIeCLvloPtWRo05OGbf0Wb9vdr8nLnNW
NQcU0y4DnaHKHzcs92kC3tiO+bN7ChnrNIB6wZef62bFB4bZubMty4RpWlMc5s92cKZ9ObK+pBcX
+tnl7cAjzKAVj0k8Z/IJXY+VNPkEz1+vTQsoh7hL6PsGb+YCUD0QpR07Igl+tEF6Q5L5CRiwD/hi
QVtLkLsjsnRHdnbHjg7V68BNYY//ao66MiBKu7I6pc544NGRo0MPg+aRSd5QAxaPtJ53A8gQBCgu
9mfRnIqqSxJtx7YNgD187BAiaBUGc9ojf4NtMYnjG72eAEV7SH6cy44DZ9K3knl8sEcA5Ie6dXiv
vo2HRl8B6rpyRu0Fj5dPRPk/WQ5mqEtne72YnWCV2lshwD63ME1Iha5YxYoIG94yjnc/mc1M80wb
2wgE7ZnNx0uFsjJIxZ+9t68UUNwGFequ/dwSRw1sbn2Wv8OvuZbV3H5LW/WoUXKS1373Aq0M7NpK
56EOv5XMpbTu100lsyS9G5KiTgOxlUNXH+5/pUvB16DEclu5eht/KRjQlapfYGT810rFt+bkGoP2
xJXuj/+DmecK3r5xUcjzT2ijQ4HdLmPMGyHrfRU3aTwQYNJib4o0t9pfPZJBI+7GPHsEyjNtw19O
AqKxxqbAAt1t1DxbKCVh+BHdPjEZ41GsIN9eNQLl5ZAU9ItXqX8xENSNTyUyc7lGG+iQCPLMwQjy
WFSvrJEQydid+Se6l3oHZCwvLcNSzWFm6QVk0V56z12WVKC2AtBSaIWX6VA+G9Nk3ODTu3p9JRcf
CPTvBM0qxOHykxKcyQ27vRM7LVv188L3OM103D773xkuPaOh1fovh6MXxthJ+bTPGrv7ZCqBGcZT
dDJOSlcnUbyD2ekp3KtFR93bR9UfpYGcwXmx/MRVNTv470NnK9eDUeVPRwICsugvgWdJdZ6liIL8
MoSll3/T/xdz79VaJkPOrADyJnU4ki3SyhfW14GiRuoxhtJWMLYiqPMJKWh9E+9vWmAPXl+f+wOC
nUC0mbbUnsID2A6sZ/zNDHGp/N47xQ77s6noD1A6rIvCdmqo3344vTxK0Q2RBtiGD8KI09XsCHey
2G8/HMNo/l3EiAkBRb7rAQEpz68r4juMlc2DN2ktxVNBQa9quheE8R28Ud1u3O+ZjSU4D/RjjNvH
RrarSS07kX2Hal0fpG4ZtxzHpEjq55AxiJVtP1+1c6KyG7v0E8vsY6J91CGDD7A63r37oVeTunaW
X0aU4rRliFgp2pSKoxnIOPDg+1SuSUFllBvyL3lLjKh5vSXkq4edyM6Wae2DRqAOWuHZx1hl5hDk
zMEFevSHTjazU0CnRYMVDje2aOnrOdI+Wzh3LLcebmYyEh/QcGmwam1JrZSE5nH45VPXekKkE6EW
7F9V8j4HSvZpfMC7DyoN5kxVf0aWOGB6DFB3YJv6bhtci1kQLXjOocfeDyCtCLB4jV23GCGSH9Bn
zt47D6Xla0tn/jYSQfqQXpT7c8q6bRgOhCi3qh2wWsEEwNiSKd1tX8AlV9f9vPUMR+3PmfEhkgh8
grIIFJLw2WaxuWxt4Kc3+j/WDKPPrhiV+sTAwErs6u+DmW8rs5HSclzgmG+WtGFWPralfIouNDdc
o1lNadRSs0+uOajZbL9muOgQ/085A24EmRWwwZzvQ1CIbu8UUWY1Wtjc1NWc7twwoZa7pyaF5Lih
EyHuPYdjAOYUtcqJBDwXiAW4aHe6CReFlgUGr3IyHY6mNh/+CFkaZVs+zvqA4lwQMBokBL+piarr
UV0wphBChkutwWsrcgoN7MH8hPL/St9s2rFtiPIr5es0fF6Re715UKih5N4bJszCOJYzSUE11jhR
0+mvoifMfDEa/x4uN1wXx0Wm53RxpjN38oCk6YPz+kXpo18Ulo0ior2dhR6wqdHEGeImWo53X14A
xxKTYVjG+2N/wMmUj84Xk+bBh1+/0Bq9Q4YT3OlPvUF2LC0wSOWc1Vw1xddxx6Uf9rgKNxjMpXb8
F/AigPgMIsSE3ZlKgD9n+5HzpWEglH67eGzgDOcdhq0yiU5K0MfSinsivbd69kz3OkQOLbGuKwSH
NV9hlMjPSApeQnAC/ZPSksBb8AMlz3irIRDSkZn1UtZNNfA/zUXjOhv3QuDzplJOiJP+j8dYzbKk
o5Y92nZR8lxlghpY9/b0jKFruKtoa8oTkjEm4RVTTAgiStJoM4WlxjitQZhRpNdcD/VA5vEDxBdo
3FfugH+boE6k4QYBsjD8ET5j16fmeY0hvJoZqSAbiOiCxjuaZz7fQeNs9C1dT3Z7Pqj5yv7766PT
VhurC2hGNSNUMHN6jzM0s/tz6sLEM5CNIcKXOHJDJcGQMYAYqUeqGrWKS6oEmWuFmFBAQeMX6QKj
ZsqW/LOYnwtOkkj3l4xpwXt7liP4YdJMfwZvGVms1vw01gTnPmmo84DFFBLwoW+A+l993Cs+BlPv
AcnsL/ypnD6u0lqX/h6mUGh+vdKxx/ZDeJgNWTwnSJmbH0LBpPdEfnF6Tk6qxLbMWZIPTOTSqnTJ
DIprLThaqVphZz3TuvlSeTwQIgtdBXrdqhojv7J9B1X9PoVrE+4cw00AGvGvkc02Nnen9PUeNAfk
PnIGS2zQ+/uTQIhN1oKdrKCdo6szqZJ/uT0YOWc/Ji/1FC8jUlo9khZuIR9Z8iZSrZ9niyY/7l1m
6RmUDjvegl5aWEf3JD7F07bpHsd7GSO09r8ZduvGFzfEyw3b1wT9g6UZaTaYw+/LvBoYOODznj6y
dmKOeWoKBa7ejs1q2/9o2S1bKzMUcKuJ2yhsbNN8gpV1Ih0cB9EnMIxXB8eB6vfRP7q+mnOFxq3B
vXI9UroMHD3cUT1lxYF7DfAbmG21EZKHLrZykB8FHVYIr7CKVDq/xDMPULOwFkOWmUkbs8oRkZhD
bPvhBQXXaa4iMxbdBfmSBKI4slaf2B7ATIRWuRINLujQT10iH7ZJUp6oIv5cTEa4BZNX2qbeIKbC
550xtCFd9Auygx2Lk3PfcROZEcOWk0wWOSDbNlZNn+q16NggYzE0IA0e8HqfwcMCZRjjQEHvq83Y
zoIWZnid6PCZyljLUe9T68klxTce3pXmNvkb7fQ2YC/gFHJczNTOR+aSEZ899cjAZcr+9Q0RwAbr
WydSiyV062V9ram8PnglzVxUbDI8qhb+U0Z9QjDoP4cT9o13VgK0UMKdr6DSTR4ZGziZiEGMk+VO
OE+ZRySk0C/D2TDVyxRCPYf5GGLummaNwkJ2/6WvHuaOczYoXdVybIiu4gy3DDUDgaEX8ZmEAGaA
RNpHfIMAiIVfDzCMpslVv2mMWI/xJsqeI2GEAwmvNn1GSk/kOa31+ZwgfvkoHFvRHQJxPBkHRYB0
yoqKbYhntxxl8kQyh6WMVPf6WsJT+z3eKAcaZQ/8ygjKnR95nBZbdhjTVab64nguy41iFu8/IXNV
e5s1HvbNAfDp0uMqyENK0cy9WrA5zPWajdmX8Ckjjd3pJZNoXII68GWo7Ku0+oblljHbmwVeNkQ2
3EfyiEIBIgOm1aqMzXJcCUhWmi8HrNCeiDD4uCbHtMrlpZMstkqbEyRw4HSgumYheSmPjw1nKogM
6ArnOo3No8oFnY7wrosqaXkWZ3xubpfMZltQgQstax7zkJlq7YyxWUBF933nzatHoY/ZOxg3Wby6
l2DxsoTS7x4S455Tbf6zm4Uq3vy5KOWwOwf+UUEdeqhxB2b3b4KBMn2QPoXglbRB+cdxfr0P0EXq
oJlbZrmlar7DT8agO9vh+fQNcoSKwl62JEcH4hwc0y+CmQug4rDYpbjFbdGoksgTFPnzYSGOi4CZ
p39nbNtQHBCicsQtAJFT5TCVYLAiHrPR1mz/Q5fllbTQOz0eysW1eNgauFWJN4Sf+ZU1OJMZV97E
0622yv+S1iPRpwpA8unyDA/cmlyVlSMgOTC/FCbPMN9m6D43dk2xLpbJk6Yfp7dQx7TNuDi7p1/e
oOWN1IYOOML4qEN0hvJuBXDs81SzkSoFyK8TctGW0YMpyD2xyKp0zgiBepxf+YZutbc1BbRrxNFb
Z7tuyg3pHsror6U/hy4ERfLmgzlDBvqhTxi/9n07GSLZg+PGT7NJsLMi0w++2acf8QXzBjlMIab+
qLQtaxb8U8JkDyLTwGYDN0Ma0ntGKmNaY1YVOLK5HT/UVitgWnVKkB08JpkFTdNXV4Ra/8ITlSI5
uaMJauEjxfbyssap/BcfNgTYKtxpEp9HLM1N9Z4CYwqC1+0D3G9Hlq6Qxv7Eo2cOWALu/lXjlvdy
sigmHpFKD03RkvXfpM+D6CBHocLKWYyPwtVIwq62IZZb7yspxaTYvIQJq9zOcZG9u5tuogz8nbVO
htFIeOHzgVC0UREvLcmt+X62MYZAUsRplxEdEusLCjzoAxdmls7/7FXaA/l7MVfUTSs8Cu1AU1oL
CVAhENaVvUWSIHXeOFqqXKlKFccHwKhFUZMAh/jGN5oOqx/iUHkshYkbZZ/yhR+nBy9j9sbC3/bS
NqFSZ+rc3r5nY2qIUg3/BETVKUOivOmByWJTFCSu5s2ijLlHMlD0ZlHFuJu4JExHhHxKyr3rjsbj
tAIfW7BxKqjKWvXn0X8o6epX/pEICOmRpABF3PPWlDUR/4czib/F1zGdbEe/kVviGLQpxYoWSRt+
DfjMR399TuaTFnWsqgxXmakPVs4HVeubVGNeqCGxkBtEV7x/F6zTNriPXzcMh5HLslGjCNfeTsL2
2sAzxZsR2XRxqIUmQgg1TrluulROtO/3vybIEksbNzV5nQsNcPnRbXMNRXeW8hKEqhFaGb8TcKlJ
Lcbpfk3oD9a/q/A316jW3pFUbGQeRQm9CSBiv1kN4K8nRkDx5OeNsaXVNeMIJYx/DHlc62Ci1xVt
HfnzXBzG6O9KjkwxneWf6CQJK18YwvYMIMRdSuJYdjO8nP5LlWPN0wfRedE1DtLyL9eiyEMQrUPn
6mLqUpi/annXzyL0TsPo6sBAQSKg4Ab7VBJOX1bUjbz1mEaMEzEEA9K7vhGYUMXvA+tjRPl8ldVF
E0TWm4r6Zp+p5J2hqqP9ebqExC6H5AZGNSYFgrwWdujRdWbudsBd8+cBIU4udkn2QBhf8Zl9iCg4
bviLCLGrPGGSbGQLCMTzXvOQh+cR/Sb2D+oLjGNQbcuEb++QMcNOfwKAnTsVjZeR4VFrOP6VeA3k
nz0Q5vOJ0P55lGjJIeWvusPhyDG52PEK1FBzFMk6+iEe0ykIglDzVjTLeRrQgmChQN6YCFM2ZkbJ
/aDY0ShaGxeiR0oBjOLtaZMxw0cGBByqRiNQhCGhE5RGsSUkjRMA8z7jTgcD08Kh7GMnAXRsWU45
mABhf0dVFE8QGB2Y4uQ4KqQPhFlcQa8EtRcqclWv5k+udEXzfE9XOzPU7LXF77JXYKWpyD7ByFoW
vaOSOkPE79/d/cAD6wpKmTuy1XAvuO2iDXtTIRYAvPtlgUl8K9sUSU3iqUpRoihrbW49aBctHaN7
SXlEYAJH6oPWjdajC2sV1f1voalNYvyhibfDFn2Nxdn/bgiMAPNGhlzhYaUDhXFhTmgLKFgM+siT
vrEtUtRBZCBdHJ7HWVp/jPNvklkbwn9Qpixm1LELyOn/miL/M2HJ+aiLLR23fadlNnmmnAHWyzba
wFZf6B7R/FChS0CdqC3c+igY7OxnPDXKbeeUOMvRQtrAL7gtRjjUIORTb+0zDL01ssfQZmUfUsLy
6IMWGFC4oARERMwIOah/I0U4csxrg9IxPXZiMIRsTz13ANp7CyHdhege4LJB2NZWIh81m0KGNj3x
tvI9RrSE2hOynPoTIySxA/63PKRYjUaJrxgzmjbxzDRkr3oobqWZbUaIZT1MFirBeiZty0Mdj4nD
+IJ6bd8ZYTEdmnr5tPr/6bqv7rk3/2Zr4nJ0Ge64Xs88DJtBvNJumhb4RPzKthx9nJAsEMxRIX/c
NuaJPwRlCLlowDiNnRPZ8FWAdnyUfYuteg3YhVykXDLZTzB7USa1uKSTM45dfq+DRdSZfocLNBLy
azsPBBrdsrLlBTiE7Mu/lwZvbzzNBwnI539vy3Nrxf5lWhyWeyGu7y977CvLkBBwstlAii4pR/YN
GjK/U9NCR4ANik1ai1DDRLewaUoePOqkOBk1ydv7Y0AcbjVaSACVMCANirsfiiEujcjM75K6dorQ
e9+3KLMrN2jESr3JvjTvJPyXRw41eMWq+C3JuY4EaU27CcHe6cZwg30tLDHoAQj2inElzJuPmbOi
Vk7uS/HhVeETFVSehh0U0G4ah/39t+uw7mqrNTHxy8Idfb+KKz6j5AaoI9Zdrnvd0yv/OgAjsxQ1
gSh+HSYbrsRIRt6iYq10q2Ql2vtWZhViXjqM5DBYMQhe95I7wervHJ/xtxwSdUKQ3T+bbWkNnUIN
AcrU/tchwVSxzE1v2gQ8cvzHZLaBX4QjgOLRQ4e55dJEGBUrG8Xeem0/CGa8Z4Wem3fVYT2Cd3M/
JgkDFWHTvPUny2URBMmO2GjB0CTD2+IZGYn7jKSkdoYs5E23BzHAg3l37ARKx/uZwEQiJc5qd4KN
GTqyP9Wny3ttpZf37ay66uFy0iU5DFGQrpKOkX7VjGKqAIdJ9qd67Ep4Dm/vB4S0wFBpzOyOmUvY
17Gqr5ocAL7P2FOVU3NF9rpUd7tVNmhGDJU6Nt7VXI3rjD5btsFGskw6UuEyQ96YEx5wLRWMIrdE
0msYLtR3iSzyTUCvWTqZvhhKfJLvZYwMeTvQBiqTji6CN3/C2f74a3UP4cFW9yjxKkChRo34OgCr
KKS58bmquVGavkyoEfs+WRTI3Or7TZY1X8nBeZTrTBJBdDjCsOUmoDZ2Lz0uDcQBaxQPtR1CFWU0
dEFVfn5m1ud20KxzfgJZ87Oyf1mJ8ur5i2VdyXTTQQHmKlYxSVKe7hlFKdJwjaw7UfeJEYV2OH6j
IeKXe3BTmJ7qATavEpw337E4+7fshBfLolo+DVE+Js39jHJjqibckxyhqHDF5CqZmfZv/pu/7Blt
+Aa9wlS5mbOhf5ucfFplMZHruRqdOCV6GQeZO8kTpkvcETlL77cUGALVntscraUESuatpTaliA5T
wmAwapkNBwmlp7JyVs0P54QcQ0c2NuqeNK+L/qByNgc45ABiUFxb6sZHfQHqUnd3XUBUz37Gags7
Vy7gDmfqkQsD4bVGa9ewWmsH6fioxdQBKq1KFwTorrFJx4AKH9n642lauqZ9aZE2TU22HQTcj366
9MgkyXlo50YxlgRfVat/8S5dlJ/UUU82gw6Xi3ckr5E1AaEomW8m7nqozthbpAF1/H20xRdO0353
CcXXO3+6xSeKmXTQ36sagHBzO/Z1e0yhoY+24S3c3CGD3kFiZwW6NMkCsmTjpEDMTuC+AQoV0j6x
S9w1S/I625FBgXnllEZKIgDyw9nKxy6f3B2ZBphswzNMvurrSo99Cf5A9TPZne1b9Fj8LRyjO2A+
CMftU7eNMQfKR0zK30IJ2m9Sed/FlSJzpgAoO1EaYfr4UsMNLT2DVlcB3dv3o+nFOW28d3Mgt0oR
2bQH6zAPSjx1QOmMohT5fx+oqE9QUA2ZsX3ZvBSwaSeBQksbIF758rS90E3UwmuOcbcB3MA7s6w3
KGm7iV1ipOOdQmoCCRRdWDjPdJ/t56OudyBtxsHUF6gg11I5+KV/QVxsW2Q9Z371IcyXLqUB2vlS
stAIhHPGb4qJDxiWJUYv6JapJQwlt+1Y8cZeBeoCkK3HdckEmebKnAV0J1dL3A9A9AU8fwlAv0Tm
wNiXCiCPnpFhdNiOGKpkk/24DrLkheupXC4b5r/H3W4Nr1vwDs62Vsxc7sFKdJ72OLFIybAOw/7Z
EoBcnEGyRkPcfgeT6pX3JwNjvCrXIKVkZ5eDPn/AOx1IhbaAqoGleeJD3u8DPN4fweHturdi9STX
vzGnwkAmLI5OwN/x0QvtBnHylhfGcIPnft70yNTLB8U/KxucxHWMt2Lycp7V1MwoVlizY21/9bga
FwsNy7R0+4XW91HDkHtkoOfDaO86VmudIhDYqzOdRxZ/6ZETcZg0OKhH7EhaJfgw6DXIJuwn2Iyj
jhU3EPId1fRK8cXG2YU1vM1ELl4hRbDlq1pb4irPblxd9qKM4zXnYByeEuQ08PNJb7bL0frcbCLl
OuvHVrncR8Pr00Z7eePmZ44Ya0vH7MjEw+uCGEyiQgYfH/7C+F8zbEulcg5WMFW9xk3F8mlep7dO
OSlsN5nbjZyD1oxuPbxcgBega2/0zrMUOsOT4lmHRua1/Sc5fg9Gr6/rBnOKBmtX1R2mnoG1ErmC
BFe2/CeYPG7HpI3EbqJpwjpCAiFWJ6ra9q1MDHCNtEnofxqgezFQhLak877qvzs+kUDfYcob+en6
eGC3/LpgMRreiISohXxYSWgLwqRPUDDah/BORtY6MD9BzfBlLbdeSrtpvj23I5y/nAEWjbBR1iE3
ZHg9Ag51VVHwaLwJVQUnoKyB4RyLkC+dsPDW6T4W97AXvsbIKxwwHGCNG9jT9zgY5VtZq7xAoVeB
2ZFcgNFFqFDOmlgOQ+03LYyjiOWbsfaBN4dOI0EXxHUC2n1wqUXV2+stKQTJdStguQM79v+Z5wt3
kYm10M2joj+2tCiMqkZv1KLlyAr8lZ5mh3Ow2/tdYAMkmzpcbY8aJGaiGqudn4T32jTMwJDQXH10
UfiNZ5urZiUHkeLevbcai4Outb5PhJn7vKgXnMzFkzMo+nPHuR1F8PqZnNeXjdlJlcfNDb/2/cfh
jiXHLKe/IAUSbWKAUM+7fYL/QovtqDW+5F7+KjKbOCC5Zd9AxmrCdVFSlM/BdUd/oUtrHNT4ZzGr
2DzRP8Un1gdaUipfdO52IwDO4UNB7pB7HvkCMXg18Q6saCRC6YrrdmoTDt2uJFdhSbzptKfol++n
FIxaN/h+tX7M6rLI3oOzCjsOLZzchwXEWoDzi0qVKJmZpSl326FM6jS91UynkaUkF2W/NiUUQIkR
DsyUECfBsDEhYHTTjC3sU5gBvd7qnAH426hsD9HeAn9mHClqJTBOaqSbxVcO7Elv1u2WVsGTztSf
9JbpXKnIBkJyaPDC19TVdxTLXZ0VuFIO7by2qBKO+LP6g+4doMiIJgf/rnN7cYhP7FrLFHnvWqO2
yQU6+KzIJg6z/J0fSjd6rgsVUtysHdCvQ+pCSyaHOYulJxkTBmwyxblxysQuXAf9Ya9ne29E5Gl4
B9Xx+FdN+BzV/NOXHJpkeI4wRnmNWHfHr9DJV0HrHQX0xcfLl+WWOD/z5vI6pwr7HdsCQHdQWcfn
/dXWzAeczAMFOJln0gwN7DyH8Tq0ZL63/7QrQlKghSrBzIRg8PM8KXChqDSIOvaOduISlNgU7bw4
VhTPL2UHSgSdhu2XvjgAGaNwcXCcRwg2W57vcOKLeRfRoTi95t1dxZK69I8PWNb7Q7E40Mw++4ZJ
Gg/IM80IqT4+HYsT99DVRC2ldJjxj5VbV8DFl1EUxYh3SSbt9N9mgrEjmrN6dmjJmGwNAorsObia
llnPFpmID7k8k0A+KMzvoxBEWrtCOdiLRTqYT1STW7eez/Rop89GkvQkgVE2Z7FXL4YP6hy+S3RK
1RxYHl3ZWLj0zmXm1wTzcyTVltTgPCxH/g1CwVzXZK5fwk7UZB2y+pYhaxHuABt3+eL3WHmzt7QO
uzwGtCclZQd/T26xtVhinhvTq6bQA+H57fRfnxwWKgX6qz/dK+vKt7MGfMAdl8O0J+76rl3HAv8f
dr1G1XrYPYwQGPWY+7zFxdnUI1TjfBwZYOLMLTRk0tn9M9f141qJIwZnIk/B7SFGPvcAWpcIeayK
GuyO4R9yCtpC6r6q8OJ3mfV1md5J3K+SlgEJH6KgKl3KS4LJzJPkOHzrKAE2s9mY/qai9i5/4xvd
1CCCfws5EERmwmgZ37g536QXfG8Z09rV2cxkqVFI6DWZ5gYu/Wk8JjsQXlKULZO9mledYYxR7MPT
vuri4uRha3GfXF1dr3Y289QbN6Nq6dHk/gl6n+t0pVchkjF74ErF3g6qZJ5opwLkiGEwgF31bfP6
KbbwAAsxev1LzJ0jSmqleAHL8ctDirEFYWBaod7/Q4z0HmqBPhWEO1FZXOzI2/1CXFi2g2N3vzf/
ujJbu4LEEVawndLVupRSdPH1mt/HE5Wrr1QGla2hR8iRSz9uCsNPFflZZOpmWdW7XA0hUogDpTT/
MAgLcabZ8TNKfOReYlnB/VKVzEABDGnVpnI/O4v74H6xlSfviP/IFQx5ZgLiPR6IRRkcS7mWFN0A
nZXvURI7Ft90LST97DOLFOHvpYVHJStoLnZAMG6beaLO0t6tGI2JSquZZoL7QI7ewjKPF+NcF2H8
CRved2SAQgGKNAp8djchhhf/LF6JPoR0iBk749JnDBSI3ajhaJHrhkY7hSJJ4fiU3CuMtv3ccHV0
7JdbYzig6HDAEoCb5bDCLmppU/Txf0tbLBEsqPYIo9P8TqoS6mGz3I/KuwpExG3FFXQ8a2Oeg3wG
N0vOaiwzBzbdC3p/dNjG5hUBnB35oSrrxpO18/6RFNYORtx/2ax2+oKWg1ae2mgD1MDb3H0F3obQ
VW6NA2HyeLURIzQMlM4txevZdcZJV1EEugcm8bzmKHvvxYu3TNgPs/ty8kOTbm3MeZRYNbV2ubTo
uUYltCHLkA4AhSTkU/ikD3zDmwx1/ZYpX1AvJd90OhGASSnFk49P1pakNF0domRH1VrElfa1c3Cn
VxLtbEPN5SGBkf4RMlMcDw3XuWT4MsVf8KSkHaMF5ZERwmaEI8Gn1Qq0QW1Nu7vKjw1Z/KpI4SDL
KkDc3bE/hJpW1MN9ZMPwJY/b5L7l60H9xoZ19thB7Q+e8BUeORTqJ1MnML+SZ8nSnYp+pdbW+SZk
iX/H2ZtatBX51OK4NpUcFxfJDDQpLi3QWpsLE14TXgunaQECF2VI1hISjSE8l9ZoC4op6XDrqZi9
pnJtNHU1RzZA3ajdZlTm0f4eIUb+8EhnIXCGLHB3GR+ZP2RKMlgJZc22NKVOFKv5Eq12DqoPaoQh
KVmPN8FxyME+SI1oiU7xpUX6j3WlbVgcuYmNCriR8mAc2cMLU2oS8ADhOyA9wr2j+49znYNA1lec
0kidOwOl/9kM7cnRgFO1fB2vSfUgp8e27dUDpdnoKQfTvo3X4QFaADTioMvaX0PHBnW93t4yZFfE
6h7a/nR3zzPfJLK+5iG4E6ioeoNqvXIquMwIi3LrdpffMV0N/pA1i+F7NiXnNjcNQUr3t7NXDy3w
A3vbd9IXaNnz8zuILBFDSqecp/Fep/p5xcEGtpf9ePH8kaIEwdnu6xZZXKvMThdHF41xNdY5y37P
EltefpeuuNbr1zVvNi+VpBEd+OiXVbYrUW+MkNHci0bcJoyLkM5INM2ARvTVd+Cy/MVSNfUUO4p+
Yyz+Ie2ZrUmMPxWBxPdOptgskQWFZBzwm+buj7EbHARqQO4xAZbAXKDrX3LOZ0F5QtW+zq0RZXAh
qIkRHC7sz38S9QvJXPdI0ReScxpgyMvh5K+iOEgaXxHTgJBECowxooCJBvpqsdkEqD/0SMXJ78V5
9mDUCQsOD1ghk7uUIkGblEAeqgumRLoGz4rRviKnS2LroZd8nXVNVpyKy0IK12wUJuvDM51ri/DK
dw0OiFR4y8yr3Lt6oYSEdE/AS83GwW98P3v+HFQEiQPTz58Jd9hamOw2qOxWX5eO1+EgMkW5dYps
dLwOVJf8Rvrgps7ym8zxJ0Sct+t1YtjEpDcbkSnNu5Wn5cvl6bvKwlVvc/C8Gp8y5au31V28yTcX
AnCEE4sugQK/weW22T9IpDOBPgd16XP+dy0CtlrhyrJJ5W8hFY60euY5VFZ6nRA4PQpzZSMEFMie
KMxkb1QQ5SVzNhI+DQSIGi+3qcN4v69dBDgE1WYzhxki89PXc1ty+BjUbw4XYHkeZGG4X0FYUAYB
er6L/80ql9uR8RtRmwT4iXwyYVKhStm7v8gCX9b+RmVeit1R8WlTFfzs2sXhxzTWtfRgzjX5z9wM
pEECQ+yQa8iuIk8o7Qj5XSGHqFWN3JyPd/uVrRC84o1RhTBH4dhNxw3nEB4T6an7cnWXwe3s5V0R
jaU9QN5FinCo42ULJjQQRIfS6gMz79LVnp1G6FPmOgVhyfC4d1DmrPPX3SGSgH36mVX4KQQsfQEe
UtnkoiBb/TprMtOAvyDfk5Vp+mO+UCCCmbRFm9eOGx/0kFdxSsOLUfVZu6ho/dQBYZxbCl0krHg6
TUCvQbT8rCO+I/nbYYRYnIDrkmN6Hfagsys4gowTqSVRgFol08rvZq53YU6aynvNjlZ1+d+PNncE
3wcB/lXn9GcCu4pUti21WT3nHH62HbmN3GcSrs4l4rqQ1LLwfeKb02n7H9WlbSWZpgSFznOjKgRP
rdt3UxtrV3c1CIRpinka3Cc3v859qmnG2iLABkHSLPo1jLTpKfK+vUMfz4zMtaI1k9gkICKYPco1
pxFHOMKKLl0AYaNbJ9E2xMbnr6es27BvZPNFKyNcWqUJmmhah5YwNtTgjLIEmvszOvolUZYyQjl2
WBIvIrOnF21+eNM+0tFfdJTo5ExwReJafPpCKQ9BM+JqqtStl/ZB8SGwBr2w8AZJVv4n48d2X8Kf
COM4cwh2PTAL57E9DW9wztNhNlU7QPUjwCYwdrI3mAcqJdJeXnaoA7qYZl41jYcmwOI/0AycgEpt
CRDG3wNJSPwi/w/bUmPPgNFDR4nUfdv9RNphxQlkftOYqllnLmXH9YlwWQywc0zeCfRzEJUn9aGO
VNXBoCOT6RBaZb0COiX3zCCT8BJPEGahmWcmgJ0Ya8v03SoEV/9s7hhE0iG1JQwaxEPE3u54C10V
U04pnodTnmpMDzyYVmf59iRBPeN8DsucGvPSe1+E2L0pQ4ShkbmadphZFfti9dGwTKLIcG5gquFQ
f+cXwcs6EFxalS7OM8zqRyeadUVboT8Am7j3CHCEsF3VNTq/Z5WF1MiNxVNovqCu71/SAeOLD/sz
uI/Dg8qD/u02Jns0nYdXhrpQ+zXBAYtftMvLobIKcQykHVwkQFP5SzG5XyRieLbWekAlMzTHybYp
luCGos6mvfHDtY5xjeiFd6jg2h9xbM00+FMEQwWW5ZjOv+dVssBNOLVe/EJkFH/xpuTWvbCr59Xk
L9HZP9C+iVKtSwqZempHyAZpW9qki66Oeup8xMXEyeRcjZTg55g9hCS6Tg9niNN0wvB4H1ooRGjO
nbMtfg6H3teLyCnvJUIMhaSTuhfgv2f2BboCY4ohZBjjxeddEHDXe4wMOSEQ3t0+Z7RDpuK3wuMR
K8SDVcmLKnxJbHjwQ8t9nMB+HSZ6Oz56cki1hyYRTBtjagQN+gRUIrqOBdwenQEe6odK3jchSos8
IZIWR7N1M6EmnR3F0cO922QxxGuRp/mDvbeOYD95LnaH0wtY+JmU1P5fzRumrb2fo4QtTvlsO1pA
EDbXHy5PxG1Mdar1P1xP+hfvzQC5iU8olwg8weCKFCGy6Sg71Ae/o7CZ2Bt2MEBHNuj5Y96N/9iv
0JsisepRivUgK+8wq7I7OBGCnamb6jTkc9bfKHxaqGwXAHe5CqHrJHbINOhmVeWq04mYdu4F5DTt
CQWLhsdD5uv39aJ+aUm8gTKRp2+zmCShde9mQPhjs9PP+6rzGszUJa8+Zv4kQJbsZ5hN4M9Qq6+6
s+7iAlHy21AFX0lAhWCLrVQyb34ZTrlcmh0xZKt3slrgbcpVZYlNCfMo+OHkTksiMU7MIu33SQS/
oryyybX+ga5+AtF0KoOUXDDQUHiHVqO+vIxg1Yy0EQ0R0EKn8F/Um53+MH2m8Fs/znt+Lx6Pr4Qr
ua/JUPSWF3GkSjpVIPePncptL0yMXxMF1CKtkox2DD1sF/SU5d5UMw+fE9Rn9JwRpMAZh7gjQAt8
aoqbemXquxtN24vAH6ObE0VOMj0kbxjX4tpRBzQbYKU2tRWXLxtKBvkaaa7Y2s8HQIZ2ZrWTI6Kx
DjJjJmB/RYH+wChDM1axi5KkIziYdheDUICNM1HGHOABo4AUGB1C3OPv47qJwFlyMNqghl9ZBVlF
F0WrB+UNIBWe6KjfmYd/slwufBno6OiHjlpEj5N3emChbCtzXfLWd4PAcWIo3Akfic1M+RXgMs2B
3tDvCHyccQXVOdo9ULQuHUNg0pecHJ6PXmCMi7MCaWC4DGgFkab4HMeMNdvVv8tb+kLAm2fHptpj
NZItX7pm1Z++jmrwtrgAWKEMTbnriO5X2JOqy/R887BCvyLJ7H9rkcNd1h6+SOEmdZuGcQMRU+YI
VAV1Qy9f6NOStVcoJ+pLYqrRUQKrxPkotlGzZyJyC95U3d82S7lW1dxpdWtLPhGc/j2pOzUzxdoh
Jj60EMSnn5+svyEP0270hOIqPw/1riI+pkts+OheUVFEB6l1it2/cTNTEo+GWW2BO21Lym7VcfGF
jlsR2EI/I4rdm6wazfVx5uVUtZ966kggBcn32uXuR5tOTUTXtRpfCDc+KnyNE/3XomQUqBDATCpl
XrQiaSx+800YX10SNrNhN87cSbIf/iZLZc7IFFYafMha4eeEDcPmW4LQbfeJYcilCWAUPP3OkTSp
FkIuNqBhcPSBLRFyPN+KOg/6+YTuGbe1/NxKK+LlfPhneD9paIH/oqsJ91vQAYeG+9xkgJ0yH5e+
vn5j0QVZk4tQ8bnTwtSNGeU37W126Y9MHpF/OKhVAFpicD4zAHs1AWS1tzOquvtGdcmC2pI0Y5Le
xvm/9LeYjwbmdARXimt5J9x42n+4XgrWEIVKseUMJnPk90u7IULU0cJvFJzE2Q5IFwe68A2ouzJk
iscRU+gUUxNZNYGxxeLLKCxzLZNqCsFMHgdHbvxoh0K0tuK0io8oLLE58K0GQhBZF0Y39olD2wkH
NGcdKQ1YUHpzIREOKvV8JGKJ30hmIgA/fl9igQFiM/h28VIu4q4EtXVcgefXp5i++Go5IMUVEkJR
Me5lY5QE185/V7aTGYqtTGZZF78eY+nE9kImkhUriJRAg5LfnjeovVL+UUlcuuC6dyc22jpKarFl
dkjtxNzv/3ks8erXMdc5C0SvV7o4lqTWrFaeE/2TKBw+AF9ChVJw1+V7hP5KNUXGPqiWeML18MkH
TYWW1Qj3TvybBKxe38bWldTNw4VtTBVRCNQFpJczaDeKZ0cOsZoU9M8ty0+zaZKeEuqptxBtmXvm
bMc2tmGgxVp0FE3HJF8zRDnHLvcG7MG3c53Iwb415V3e9my/+hRdSyM4E+3gEQuAeci+D4ird0mQ
Qidwpx5qLBzvG5YensLoTMPkZOvG3YYCE6hb5QCx2MY4F+/CqP30f9A131khaLHmNk0dmprXFYJ/
i4kMiCu/4yUyQnTX1TudqYPA75kt0HWBxlAs9nqArmNob3nzNoLsFjaJX5yNPJI3z2c08xoyI11T
w1g+ImxYMhLK+v0t2QYiDRsckcXzjTcYb5/F8Z0VukZe+k7SQ/amiQh59eKHsKLqoanbf4z4zcNX
xZnV/o/udpUlXY4CJwq+g4NRdCXbsrKIpkMFH1E3UkJxGela03ze3b5rEvC8y6dEXPicG9itSTDI
9JGlO6b7e+ZGkjsNJZJdRsNzc1dxj9UX49jCciP506sYnXytkZGxDDc5mpKse8QHpjs1rjlRBXNO
VcXi0v5fEzed492E5ZVXM3xrF0a5tE4me10oEhfMGbd2cOpmRCU6TU3cmBR5clzSDNumGagJ6d7W
P1Ivceb+vQKWN49L00v4NMyNVHgpPViMp+VhblQ51PekomBuV0NKn3YzNtMIDMC0tdj7ZrXrrmAM
udMXx/Ui7i3U/9f1JqR/+i+ihwmSHnuAPoXuYdvkNy1yARctD2L2oA9nC2MDvW4ZZ3sFTvD9bje6
nQY9/+raJYBRl0DT/hcBrNWxzx9U29JmE5vIK8CmsQUQi3JLnrkj5wF5JcC/ICT8n+SNE4LGKTqa
B/KpgEFGKJ89qeV0jEO1pkw/HgJ+8FvdIuteafK+xwrseTxJ7BS7pAwFtuiQOK0U7p0Q+ARk8Xx6
UaqJbFI+bAdtl5AsoaN37AOKM31qCvcNnyb0ejaaj+2yShOT4So2RAvFoNNM1VFWVjUxqP2bMx5V
xYJ1AN7lClNLzzOLOfkNo3P7JWVgPea+xi1DHvVoI5z4mP5RElHym94InitgzvLuM5GnFAJwUWBn
9GgtXbWh0j93hw8wyXdk+Mo8TihqHpVjk6AsqXoes3e6MGF/Fk6RF0C+x48HVqk3hCpofz4UqbFL
MKO8pgghLQSYC1Me7sugs2k+wKkU3f51nCwQkD6xsj8+E8kLB5rD+MuWeUw4BdAkHZkrXhYsGYPA
qcJt9v66nP5zlvksHaMd7N9pFA8sOom4F1OFaE6RdHh/daxxTSykjKT0IAvmlH/VZtBmVgDa5L4L
4fz/AZM+XTwk5DW6cVga8sUxqAHSF5lCZQJSZsWLsqeq9QpaRUSAXJEDBrenmiuSsQMRDMorR0MJ
w05lRMSo5spNGzQUEHiy63MkoVXqMXlt9VdAWMlw7zSIvykQ//xiskL0Z74noJzyzB/2yV//Ezzl
Cs2U1ywTyJ8ykWhXjvH13n02JhjLJkah2IBbLYC6vLD0+WNDZnPjFow5G5luURsF3h7wX/kjfSGX
Guc2eyzv6/lfw4kAaG5458WCoyNaBfZeISLgvlOhaq5PjVJpJZJnezjs1GLZ4sSwPVTIuErQcseT
IZD053OTWpbfFl6FCWSJFmifx3TXdvWM7393cSH9Irqjo+Di+8Kgw+8hP9EuRUzxV/EBoxMCIYtB
hrQjl2EcugTDeZU2Bkv8hcFyofMOtX4ugpyUSVVu4nYAPFfqnTnRJJp2R+w5EFVa0uApdjPOSI1m
IGOIMP0JxjMVIlu1Zz2RmNhTsLiZJLlz94l8JDw9Jy/qgFtgtv1oco7YM2K4YtkyM+MBdbqLN84z
iC3e3/oVzqHVTzukt9l82umGJG2D3sudjCA+dmojDZ0Q/uQa5zRPMCDrLKTWlzliBKD0+GhNX6Rd
UQ4MT0Zesq3zuPMlC3CJ68yxtds/BFU0bBNbH3aqlvhSwWLokbYe8IIVVLLz236ura0Ra60GEWow
/IoMjdKbJgVhH4qkAv8FgF36KFajwd+l8EE6iymmG2GYOhLY1yaD5wFNaUYHMhq+4c+pBd1plxpt
3IwoXUfZB7YUQctTHlEcClnE+0fXTBbqdQkBO6Gz2+Htgj/fx5LPm96uQ+k5yGiHycYENOiHCyiR
WrpFxIN2REtHUHMS8Vg8zyeoPFO2w/V60anAy8ZBGUNLq3s0UwQa4oi8cQ9AB+zDMrg6OvOZ2IHz
ZbXH/ucgkU0rBkUy3CcveifHWCgwTbFcHQ5W+At9SsOVaXEjNYeyhdyGDiQOGq6Q1B44SVLLafyV
M0eEaS1xOzA5Udcg7klvO80NXCla1f9FwxPFo4q5fV6TBItFYrH3XItdGMIgvSsQB+a9F/JbWpYv
Bls48wcUcWP8mgTP/V0YoB+CsLOQETTVoO8OjLjNWp2P9bQU4TeC/eoOOGRIaO0q+KgHBQPIWtr3
RPKEklZbheDZugyEeBQHsu/+x89sClIJagxdhcyed5ZkG4Ngv6pLE7/xO5jMl4FWPam6v2IKe9Jm
T6DkUMeCNPu/rTWCOgN5b5pqJPhK9PxorTba1kTXAS4ZWs6kq5GnxZk7f+M0Yf4ktWNKT7zE03yF
lCb6NzehgoAg+AueqC9V1QwlmAcietQ7jbFvVdazXeXRuiRifMC0h6zjUkxRaxobzlqn5zL7Tp9z
hqMZvWvnphnc17vxYRFCNz3I1PWe5MaD42Nv6Lm8iuYViss5y+UQSJ3HLSid2UwO0aYM0t6+2Lzf
shiLQI3KRDiQ8n8qHmOOavTWp7T16SBWfU+YTYqhFmYSChGdjibbrbhAE741hyF3QXVkiXrlYXZ7
r73YsUNgKJ2L+97ED0ZvPseU58bDk8t1ZqodcN5CRWl+Z6cjK2yl9zxd4923Y2rKxiutnp1Ravx+
xHfnm9JQd4feBaBmgCufLOyxP0W4VpT6bzyTRGutfj0jU14pVwjFOSRuo9DLLGGkGxmmtdM5wMrH
ExuT9tn8BF/RLlLjB2zCrH6t7NP4JHN4zhwrNR82MXwRJB6ZnrQdbe2jCbCwWqEMDpw+mlB1s3V0
8EFaN29xc9c45rUYe+WvQLrv2jtxnhBHNOGgh2sPGU0GaqyeGuroIgR07hu3TZzTCaNQcoDj5IEn
nosVMduo+5Uag7QN4y3N9tWdeEZn7HA7FyU+g5w+de9Y/Tb2VjLtWF+KQHsoT/vxZybSYb5xhVY6
tCyoEqnSQ2HbAWgUptSSxGXFkiYs+mj+Y0srUcFskdsON7DNbtKAye+PEqalf5wpwVbXosX8z7ZA
KBQlT7uhDFxRFuV17GV2lEcfjCZ6he5UHMqhgXlJVG+N28zOWXXQ0FDeq0IsZV4GTO+5kD7Td4ZY
Gj4fpuglUsVZyRzTgZ+kclo4or9s+r0AxfxNMQ9uJeUaH5vlgSyvWztW+OIc8jK0Oc0sKQ6XaaCV
xLqNkNGIThCV89RlUv+ooR36fm+nAn8BzVupSRx0q2kODvoDJigV8UZhKMDmoJW/i4ewqV30OlFx
IElDgR7t/0IGYHKg+eL3xrv6SXxoBJVrDeRW5ZTCbwvtzFRONiAN2yZV5BX+nfNKMbcLTuYKn4QD
E4ZW2c4tyGKmM67B8fSHJju1kZJwv38KkstTJi/Ir3RDQWLcBRsJi+z9ee3HapEl1yzZ7n445CVX
cfwPY+o72sOEJGJ2brKKlxpBthEtz5uYv3/8Gjv9Csp4BASkDcKnvpZrLA7xzGNLiHlLx//Lq1Br
xGWJtTP1cGBSeLefITnCWKaV4OhOnrS3buXTxQXADUdZHOJ7iQpNhrfCiM0LQV2QWBUaGiXG/dgf
dOa0N/6oKlHnfgumNJyQtQ6FdspCRQ9QDdVkutnvabxBh3yoroOppRlcFgiEU9e9Ctav8XIrOiUP
h2NMesKXx1qW2/vG/HkAk8ElUm0MQCnkBwAQcxtBPHc3V9OXVcE4wBENsM1PMvYlF9StRRk7cqZI
8xWDa35Kft4D901qoGYHz9bT10BCfx9rDcAWOh2Q0PtInzmpxC8sE5Xlu0zpfDn8/rtfKjNgw4i7
Y5AqKB2smnMwX7TXFUaavmNpSO3rpcoz9Xw/cw8ydedkPZ5jgMVwC+ujeVEyev+Yr75ULZFWQxl6
urOB1bLbp12h87xM1eGde1PCwxuwy/mHI3uwyvUudaO/M0O8Yu88mqi+kC3HzAxlsZC23/nKh9yP
1NLZXvHlg35pki+Sl+V6cFGRWw+X8MdLYqBdcaFJGvxOoQkGzLr2queLGcoNgxqtnDf7OdE9fQtb
MOYlGcHJEeIbEtIcd4LSKhv9T0hTKLOoaSRfzV19jMiNeysyHWT+iULAVCqIZdW5OihzDz3+2TAV
npHZlDv8WfkO0FnPW+MaBvj3H1gtGfceptAq7EPRvN+KusAWvWfanEl+UavVJEK7o+a8KY/SKG6u
WX/iNH83MyMnY26sOBzwmHnBecl3u9V3XnMp1NvU5lJgOhp9sVbIByNQSqj4gEAjUd76EiWlFwT4
R6+xLqPU48Fge+BnxzDRDi9m8hsY27Din/kFUSQ0p2knE45TJ9CtYVHBtGM8CwC748R7SjUur9+3
Tz0Z+eKMKXprywKW7kbr3EYrhHKxYTP4x3aitGaYswzh36UoPfe+WIAEOUUPXGKCWgKYC3b/ZDNI
msJy5qaF6iQ+1/NkbowDEvF9kE5s8Hw4LJbrAOuUYUwU0WYbbQ+L2T1IFWugUl0SmXr1pN44fxlr
MD9TqbcQ2x9qOcaCf8luMjnua/hKrboUcanVrv4LkxPsTavgz3rh59A/KpqdKXpcec4CFOQ7FO5v
OrB+nXCUlxuLVWDtT0FqZAcVrYhThdCgdJ3uIbPFLS9GzrPk8iwgoumKB0dwSeEdJ6e+2DLG2bsp
4Nm5IG4BGBXXILODugjxTVEmQjHClgdkDKD7sLaQyAvWSDuGRD68rJBgs93ZivLcxOMNcdJJet/E
qfwVK7+TNhNQkrMHUpEeMN53ENlgZvKoqS83rRDx16lvN9fhUh1PcDORKVf07mS+efrhucOe4Zhz
jZnthuG5DM3Q+djzZQH5HalKjK5HxoFNiFtTZSjw2qqlaF8s+soHoI/zIDY6YqqnbBzR3rmcSgPZ
Auulw3pmmMF/HI6pAtWbPPmV+ZKV8b1UdAiuM9E6m4Iu0OcfytSuWAAjLxkPaLzlzr27rQrVgRbK
lQC3R7F13WdJYAC0hH4kzgZ8tpeIM+pnuC1Gc99s+Y6Fl2bUrrPzvyb2FpPixinih2Vb82HsCJMo
Kf54TLIZ5zi5mxwhQ+tq9I0aXm9TWDAsPhcxbILDmNYoVj00m76lBWBIVuBQNh6HNIsDG2bPfVSR
gB7OsValZzR2MHUN4rimIjiF7pdpfPCv3dzWb/AZ9e8wCW8Rv2RP2xMouLUe8ChgCfOemZrz7K/8
seaCmHGAT0fzLC5rcnJzBbChcVq7G6h+JGiSB+0pM/O7vYHljdmvV0USVfBghcEJxe4eB1OEqpZG
IxUtYkgvwpEogvmIULSxtSTBPd7OshFNVGAgyDf05uA5VaivC+JM5uE7IRJzexx6mimbC6G+tf9E
/7eSVk8TZsUpSN59a8FFa18Zd9DLrE88HYlsnwlS8phou11hDiz7+mOPR612P+0835hjakFIBjL9
BJ97EcOXzzfhGPrbemBGwRemsGirNQdZiiWbDKvKJPZUyRkI+PnCOtLpnjnQJHR4BIj3gxsXzPdg
Ff8/ZdgDRi2oFbhty5fawGj/trbe4eZR5hy/B7lWjqWBmwn+Z/b2Elvj8ADJfpnMphoU9ZtW2i3Q
lbPoxUTfXb9xFBQY+dxRWDs3s4POAYm1NnrqY2/VftUxseEgCpbwhOF0oZoZ5rfyG7Z8y0aoXMsJ
gTSFelMqqlQY93dZkW7v/uqEcXQKvcupPpWjTu30mjDCednJmCcQEHv++5yzJe9rEfebt75aGrQm
RZUTe6eCb17Q5Yh5UyfGSRoom5C8C1J6qLVKm8hCiEDE4EA6wrFeYfArgyCGhBgRalY79vs/CHEv
Lfz2bdad0jJeM5dbgZaWIaYuD1gM8OAfCNLLzhKU7MxHP5kRZzWNVQJP0l+jEt27XFGMHiLuRf+k
P3KNFJ9Guxz8Nisqobx9+7zUZUs5VaWEwDrWa0EpT3DU+Df7IAVFUvkjKWjhXAi/KE5tskiW2XY8
23CmtgKb/P3ZYRW0LwoD8ah8WUWco4GnlACC7aJl6TGANYE/5h/yPykWwUO8xyUMWkusO2SOfW1O
Ja4uT5pPnqCJ66FSaDXn/pZkvLal4QI5W2eC04YGag/KUnihp1RjK/8R17mNpkpf38AuV5EchUHD
8j7x8Y2fZBjh1U9+5n2p5etjoTFOpgjTv342u79SH0L7IEoG58ZUjsyICZ2tntxyPALnJtnwrRCM
YqliI2mbZGayuQfD3XX/DaRDZOf6UJoJNGgMwtMut1RcYpAhW4QdpGAx19bEsNNrXog/tiyhScZZ
L8v2LILdm/Rr6CGrL8u8GTtjE9345VPPBhJ56CrJ9GO2Y+OEB9WcEQ+HQ1Cte3mxRwN3fqvz2fTz
c6MvoK2qy/pvQXye/KXZpz3RqRCucRXx6zeJfluS4n4ut5t5yBxFxmt791FQXE3U3ZdFX/hZAmk0
ywnQF3gh8G1McqEntFkXIQsbplCQDEdKtDvbKNMwT0UXtVjxLv1bHsPDrMG3f/Zu1Je8RrlotITI
dwWvGUHY7Kh3guBOAc8adkck9V18Z42GIqOXZKGppPLRijs2ChfBOeStd8VlmpgQTYxvUACBv009
MpGhu+HMFXoWbfw0Qd9rUJdkV2Ilbrg5LmE1qaHbNVm+a7HiJf4TLG4bpObhgR/aLeIfSwB0BELI
y3vN03mf/cmO7cfavgHnDZ26bMy/cS1NYPrWaDL2DnnbAb8wBbHWuyUZ7E6q+qHnS5ITDXCUhLsh
uPi6leNAhEQerSZLiJySUrNl3XqnVp9Iyo12nD6OiGnqVKY7aN2gkPVEA+Y6EIFbfBCBEL8ljm6T
tmcF/DZFWbzIQrUW628tgGlHYqw+IuCpvlAhScgQMc9CWLfB3sYhTyOkx+RQlb8LohW5JzFTGs9s
4mlVMn8u8/AMV/6hfWWl/PiMtT8Ob0dZh6jNbBUWYTLJIi17ouds1L1mroztr4KHZMmH+FtxAN8f
d8yXgsgae6fgIxGQOgoaedOmswdVFErrJ+A+Xm8Tt1v6XHMi5pn/M/zMaR+gacniGhNR4vkj9M17
d/7jXlBOiEe4cDu7NYh3OBQvd/QRDFnw2mdIFclDNpQzgjOh9lPyzJnZCNABuW2hDjqpLfk0HsF4
p/53A4OKcoWAxn3iCLTGRdyHw65nwqx8jVBcTV+aBcg9UmWgHRfkN0Q97VPbm0cu+Ta/u0psFx/F
RC+Qb/mKPpQCtCj/GUIieuIMGOcfN3oL85a3G8+c9qG+d+uvm+U6T+Dz3x1r9Ib+Izt1urT7QyJJ
lLkpgjUUbBpAx3h2dSHO0b8upqMtUJn8da75lm63S8O3YyiALwI5yOaZmSicyY27nrg3gEqNs/Zc
SnCMk/ki9Jl1V+NmKQRHkZ2yVa2kBuRUQgavdk76Q2fQg2HGf98jO/6zp0Zg1sWz2/LvQSBHRVM/
3N25zWryCTI8rO/XVtMkK6Eh/AbS1L0pcO+zNyuhge80gj5nYW0BL9V3Z4QVl5JJ7O2lCpi+6/4E
5rr5CylvUc5nGd1AXVz2gAXeD23KhwMTrzvY1+jUDelsS5PUh172e0wmpiGwsJfFsTeGiNbCQkI0
0F2wnvnPHv8oxtb+GbrKSKrSwel2hfAEV4rkG+gjwuDglv2ivi4Ja7RnLPxaR/IXHynoSfKobTbo
0bQlyp6ydlc6E+WlPT+g6fi7WI31ps1quM2qdmqecTT85peWW3JWXRkfG3Wl9TO9wKUkdJiSODin
u1pLO2VZyeMpoMnIJNsRZrQgbDHJ/Kb4czJ8oGIT7S1kAJ+H3o0X2Lv62nxxPeeGFgks2EYniPsj
97RlLp9iYT8qd0njVxF2Xc72JAT7u41OPN2w1LiGNgFP5n4cJHv6fH9yFtnHADWx47tNtCVxx2q6
Gu1dPwJ7yMklE8dhiyrnZ94U9bccg1TPy/tG8HegM7esW1WcZ3RaFtL2ger8lM9RnZydN9IG495z
VaR6fsoKf5I2jFDG0WP/la83fLRV+Jywh7oaxBC9OvhbS2v7lQJERZGI4qx6pKizxB5hEZBpMo7Y
+NzdNc4rM+AevzEPj1FGShdK7v0UeRQv07AthCHDnoA3BUBw457PfJtfDNwMRXVwXtJSqz5c7OFt
JOLte8Glrp7oFskE4RtQt700EKb/Zmk2ELmm1b0GY/7MhmrhoolWQQi6G3dK03Ojv6pUA4jm4Fst
GQClpS67/aHRHwjLqkdW6gN8FFeEUHk1U/U27zgDtvii0wmCByUK0aZpoV4xkVYx7x/awiBVGCtz
on6CB+TWwl/6atkyS8g6VnhBkQLslPqy1jt4o5m0qD0XY2Gc6hyvpnfXuJ2V4sQqncv/bWLnEg3J
NEfoDtqtgAn2VoJDymMFy9Q9e7XdFqknlTsbtStI/CoegP2OguF0V+DxxI9HbgNyup5zJX2KV2VJ
Um043SyU0V43WfqWdf8wxFBrhtbvO4denmioS9t38L8rlQOQCRtTW6osESBZpcMEVKrYe1lCO2Q0
sP9aaU8Q04UbmckEdQZ3naynOhzJCZXL2LEGacpzhv4GQBmb2pO9JDRudlY+XqWcVe+oyHH0tnz9
Xfp3LeLwcQZYt3jPqpx10i/tRuRFQhY5DFhVGkuc2cmOefhoJdm14iXSQ2j0HgcjrZmK7E1YjJ0o
N2CsFP/xhLdvP0rEDuhm1zgCy3HrOQRfilNTnEY2hVylsOSUJi0GSqbx0Ab1NFAGt3tzFRmbuiad
vCOwRXj9jiJmI8aNt97OpLCnFOw6KMLRlg/pJzWTlbrUA8JQftnPUAzfqXDkXR+XcQpHLZwHyGLy
GOrGH5MfurPUuoT6adQqgxAMpUk9r4Eyl34GLmiHbZEU7XIb45GuPtd1ciEbVmakf8aBkRE1R7mh
CFTUtGFxMAxBCQa5TzW9mrK6OoYBJXc6X/MpNJY6o3OugzsBDvAB0A4I0dUkwqQdjmwONhk6Q9gl
I7JgTLQmKFxEvjoFnk/YGxqp8aDOcnDjFszVzGtauGA9Rf5X87L9FNPkziZDraw57NjcdW8VirdC
jqRID6ff/yfwD33ptc/9ZHI4Pt+fkKCP8P2/QKomk3Gtap8aIhAAUY/vxYmWSs4cU6uLW6t5pnoT
7E4F7tS7yIfyL5cKM1KHfE6Y9AdX/YBR9wGms1JARIhfo7DvEegwVtIZf5BM5Jy3DXTfWAyaftYD
6U0mas0O3XIXXgEvMLvSLbXDjn7kPQJzjcfI3m5gaUDbnc02emHqMPQt8rzwZsAHXAO2dLS4md72
mcZJBGd6zaH+8SRmQELYhp2JF7b+QOVp5EDkThDTLvxYW03/MYYggiJowjpzFAxhZJwrH7OUWtcE
DYhPM7F7KQjc2yqBKio4xGBqti4dD5uf8Gj7exuA+ilPln+iMgjlkTjWs7u9USoNvNxsaaSQtmtg
esOzfuwv+aKVdn3iteySJNUiki6m+/qmZ5hxRyTOXL62y1wjcV3uHrID79tNv0BQzGK0jQHPhQ/H
LbzseuDWEqbc2VPZdSppe0L8ifBmJVBH73RevGC7FtCD/bZAO7E676h2ls/mh5rQqMC08BPKQrs4
9C+EEfJqHE0i4EwY3o1XZihSqxBJZh0/+fgVTcgV7fzpACoNSfEDHjetB0uNE4/tzTjqj5nENC/S
Ck2lY7482r0zAB3mHwUvLUgvJxe9syukFHQ63rmon9TnR91zelUOOShg3Rm6PbiVvPNPjNjEUwWj
q6/02fq57dFYZ36JM7oBp2vchlluwnFXFIgogWz8+C39REA0SoYemm0HM29ga4eryK46KDtVbjyH
A2QbzCQOa1eyny6RK5NE+NQ0nPBRgs9TzrHTeRVUUljRkPm03Ces5FhrQBXVjmfHbdWEiefkF8fy
TAsslobiGtqNMXdjmrXpgPuXKpZHIoXtS9M7uRTmbHEJBtfi+QgAIV8M272okeDnYHPj6+dUkszK
dPWvO1xLGLNOs6DRr0lh7D+CF8zLEdRFCSt0KocoZpgFfCksddFYmvkKXLGD7wIlaWr3xJ354YnP
hwIviP4Ds0Gf4zqbS4UjbM8SLIcyDMErNJ362aAUEeacrXPcopIGrc5QZGhMg0iYfV8kgPC1CE56
+taujK/aDcaYZPzmVNa3Akzm0S5fLPxPQ0ztzw3MpwICuH/FCVKeJBRpxcIYW4hU2v3MX4xi+8Gm
dOIvQ3MqSEtYoPxQGkvKQ83f3GIue8j1xiTo5g3nYsIPMzCJx6S4N8ct77Q6pD0Kycnmy0hsL2Ep
WDtAwSWTBA/x5HHKqroNU+YfwXeEk3FphvnYhaGUJ5p71a2N8Te3k/2w6gpOd0wLA2NJIFfEpWp7
HyrvhKFoAVBlj2kepQigVZEtqImuqzozmRKTRGGjX+CPTEgSmTYfGntHxXumKrNtMzPF/3YNf0cC
Vcn+rPxEHI1RIuia6wy/n0Xjr84JsSpjgeutSvlEADZWOXUmUIMaY8/FzMn+2b4jMd3/TLDT/Uek
Z2hKuAYhaTfQexC15Jy9f03qCinJJRAT+k6tvE7+VYfXjpidZjxblpfX8Bfr/IFGxyfbFqaZl7ye
AKd1qKz5MwZAWsWdF7iivo/Oz2xaEp6MtTPqPZHgPVca/LLYiM7i9Xwb9IydRKWncoX2ClagSY80
uy3IkDJpdk9MNeYSJl5cTvEpTYcwGlOvnQaaoezgvsfzxn96HHZiSPs4u5Wwhu+599v3Ah7ChaS2
e1+C7/mGF3zuJS1J4IcIkZik4XIopRX5eG4Tg/Tv6kquvYOtSGa4xs4Aq0TEjX9ER9shQJrTDVG2
uZg7SM3Qs0jd/Lt6/FW73mwAAH6c2v3pFL0g/FQQqfiO3b2cY0DCqZdiP4szQIQbi8e/adilqRMn
+Gknqim2dmtuLFGVi1GDFLwkTWQnObdOojXCvJCPDAfmJKza4WJQY6LOqFLsjFIPiIHf/KxTHRUB
3ZutBVvVpgkgk191yuhM64/47BRBZBeDzvPh/yiFkaSVY5M+Ne1yLbiw0v+faa10ocCFuSPq9CoJ
lsIqMce31qCBn231chRPI6ThuaKUPmjwGM7vNhl308dh7Secm1nkosoOx/hqNh+oQoQ8GRjWzyrc
ZSazi/G9p4TAzCAfKBYlW5QDCtjVBvubviMGwMrjIzQAXnlQAiTUWRfDUpj7D5yrwf8OYvBmtWaJ
nC+xtL/yZhOlS+gtOv3rpyD6wuDIMNgNxj/WD9DtGXbfZlRxqmLj2qNLmcQcGSFRWaIIysp7JGM/
YqVfuwBfpq7HN2MP93BHfIm/9cvPtEc018Cl0QStugk8Fe2PfkCG9JJFli0tbKo2b4J4PmBXSJVn
C/L6Z3oS6tWE2qqbOuvrhxXv/OX3/Fn824O9AZFshUQamtvUo+kdpLkWYHamWLffJALwc7DTW/H7
5smxTo9mEPnjPLpukWv8W8dySjf9m1w7CSK9VecOgJRkvHi/WEBU3DuNUk7+l6E3KYeXxroE79WS
dqVwzmzxRfSsWPj6TCWLqeus6w5CzdBIdlfxVYQSq6Mk3p+PgiX3YocKNncmA0NI6Z8/AqA/3Rxp
XyTycdu3VGxT0QMarZ/8mtW5pLPVaQKd6weQ2aV/I2Gqw2QdoTCR+KYGRor6r5B6sU7Dw6B+B3Pp
YKRF93o50VJugfSfVW6tlmVMkHpJ6izz+gQy/4u9EltAMT05UAdD/a2WnouQojT+cQefkW3OaRfM
gktyAWuYi89YUWofxWu2qTPV4lEOnLwztbEoqtH486kUQgmYW9PYWCVSlurY4FWL9dl1fTrBCp/q
u/77fG3hpTsMSBj40udwNY8MRWtcbMpzdwY0R0BKVmy4Zrv7lJJcvMPGwCe89TPWbHHTJC9njG0X
vmSSkSHcSnrujV+6Jec57hYoJqqNuPe9Qwl5jimEvpvCH3KKMOYvxWCh1yOZ6+qrU1PTuYqaA7Ql
BarcpbJ0v376e58xhkWfFbUNDNX0oPSsAjkgeBjf1csEeKaLhUZQJ69jnw7lyiSy7ehYTDlbYAjH
ozRY/c5IXcq0IodZT94U4ZiYpFUVltJhXmUNxtaMCC9XbW7mLRWm6QW1ssz/PySP9zo1RUmfkWLM
z8aA6RmURezpRT12cpA6S6smEc92v83vJxSWkP8x6TZDpjIw3NyZVItGiKRjOjTYhPlFaos/Q/u7
kK5pwvVhk7GpWe66pwI6WZn7bmNETRJC6olmASiqeNMzkPFbbxDWNuC7PUbt33bf0EFesY+Xv+xQ
Gjr9yn2QA/lhIveN5GbxY4hBKe6G+G4cdjo/uicsRvofYeAIvvJ4mk8ju/Uks3hnapY6kRBS4fIw
ilr0Ie320QlI3wThYAs8svmgggJT9intLIAkTd6FDqL7LD2VvkLRCG5BXrZHoWnrnhsEzuMJFEVW
gC7gdpiqIi9KXj+h0/c8cwQwkEUL0iz5jLzrCHc6nQSHYUiB26m9d9CLjIfjrWjyXNs6eQvdera4
axvhhD0puQTzLnkhz9s9UABXDqjhl0dQvkdSoOidnyaTG4datwhKsuNQ3/gYLxIl7SEBE52p8tDe
vHr4kLm2+vrzQ/Ft+x9eddIgaxPvVkIYxdVjxNUMuh/OZ6B1oMCBUqmAHKUYXYPHhrC9XhUSzHoH
scwKkrdxxmtCEuCAj/gNbdcXIBmtZsbMpp7NY8dnClQHkKhqU7Pbh/gVPfvD/8oJN9u/S54UZhzF
kj6uXrLPEzghxcVDmHpE9iTj+WaXrw6hKvtJ9ST4CAEcHuBn5zITwtrlFQdfHsuSgaANPYFyoIqf
bNdC7vZmE1g3OmSPGY291VXoY9chgPa4vmOSe9WwRP7b4h+XgHyRkMojqVA+2pUxvMJaO9eHV1HW
N5h2FFLarCeOMNwU4ljJcUz7vSIft7Ego8AePHab4sVas4z8CC8DNe6vVbIFmXe+WRt8Y9kGIhhT
LYTMWVHvutBGT4irfcTj8a5dBhwFfc7kb1hjyvOSILMhzbsjqNwjJ4WWU7F+ceD/mErwM/Rf+Iyh
im4UQwV9lVTzeaNKYoX3GPb6t+9v/vpaNeBpy1RcKn9rx84q3lbBDH7x90nOfeah8y4GXKK/sYs6
ctxiC1jyUfQAk4L4vKanSAYTYFxI7nJqXCS/YjakcjSPcmI/1WEdFZ/UHoBwTtc+EyEcP9en7LsG
bNE/rmnvhSgCp1upKQmEmgk6WxbRznLQ35LRuVNoVfcLJ8RPPPLCynyWOHo04HgQjH02T1RTVksB
G6erg1YtUq70vUpibREVNl2m2Bf/DtiMbBlEpdFzl3ImpD5JUifE3wCGRSuS97zxUOOFUJjjSjOJ
m+8s/OuCdQ+1Psztt7/9PYr+Bf9YPm7F8adjzscKyY3tWfbC+pZe6wwrZH4COnDffDj2qOtl/bor
gRPOHBWnKwQFt3Y475hObOZSMEAVkCB2LRzAfEjrOkfKtok6KraMR7aiZXExf4UekcelQsJegUbx
IEtO5EEX3C9CD9+IouxNRUF0JLyCEuNgeCqRFBv/310QP2EXQ2o3T4mIjP7mXv3ukA7hJpVf/b+r
K5ckpeHGpKJ8IJeDKAdJ5yJqUDF4Gs8CBZIavziB0dpGrCSD++OoZvzjnFWO+Nxhhei6IRVoLjfB
fYP0VkU6tsxIiRoH3JsgSrxQ2DYAUU9oxC+ka1N7Yzx3quHEEmFHG+cG211vrBAw+n+dY5RW77KQ
+Df9QXPenbYPRS1vkURRbyqNK/s5R/FgD4EP2XWy/JeiN3pl9/6EvzUtSNrOPSvuT3Q1J7As8pDk
jmUxQp9+9fKDA3nDBX3D4AAWjPcc7aL0pk3I8hqt50+CDvqrGnCrP8u0FpKi+FRWTxltl4FVLM8B
8j8q9nlIi8gKU/KopEY4pWCq6St9/ye4zz3+2jgNhSoDqVeJvf7XBTOyMriYkxvf8FHS/AWW4DO4
ftX5Zf2xsVBcxvLEawVjiLuyHahLNzn8VeBXlxt8Qeo3rDg+ve38IJH/0OHfGl6By5DAHTrrdD7b
+jb3bJpYtgvyfd9qu++hC1skWUmbYTcXVD06WLqJMYpQDWGdgTsV/vXpL0BbSR19zacihhJM+WP3
z3lXakLMBuVohU0BLXsnCw2jnbNXwdZH/tYDRi0vgX8pkmPpifYstRRE0wjXsuwwaBnxlA0YhQFt
szSI0b8E7orbmrx22l/fJCU0Zd1gVlybbZ0k5hBEf81zSORkQ6NvOxArsiRc7o6Qo0kMMKYifKSc
gLuztCjmrnqz0dLvrcJOsGk6HN3E9GkSMqlQOv/I26TGy5sO0ig0KeWeV73obd+5pDuFtf0SjFd+
I0kMcc2fvd4X3QsJ5Qs2oVylCzJZyA2nDMNT4xkIyuC9kpeJe/9OwmsIrFfhd8mxCw8pmE/MisQm
ivY6NxgA2bAHL/YRBqOQEa4YA/Yolqz6VUEkz03tTOvaX6Z+eCafX7cMVEknJ8URz/pAr5/2Etgt
dH+1v+dxjk0daOwSec3pMIlb9cEWJs+qaTP4QM12EMzY+fEtkzC4OCFIAsm80FFAWZKRKUHUKGbi
jZ268Chrf2a8cltd3gpcs/vOy2VhArYH7P5YHuFXaQ6j889s4hTXg7pGhVkPVpoaAx71QqdrY+bT
LItnP7QQeBoDlamXUu+Oq0DT8jXmZIf4XLb9Mg1/Iq0hAV9hTaDYMCYotTcPvCpaBLJ8K60EJooV
16Gd2Wc+4XtGvs8CN8TQg8SqlG+6FJX8Y5kjZaWUraH839zvM9xrsFf76TH94KW8uI/eP/fd5MjP
qy6XOGdfyzjesJR/JVJSI7R/Jqh7qhPLbjkV2fjLWQ+pzL0mx8AsEpkTIqo6nPHdJD+HwPbWYz3O
LcvNFBV8FuaDKlPJN49NSBO3fmf1CU4bWJwnAtqmaNYJD0dlM3vAajN/hGVve+PtRpVqGuXZsv+G
2QDX8fKaiTmn4wT0u8Pu52a6OKPgynopMvGSq/tiko+l3e9Wn4v0ZkFkDO0YT/1QCW38nhS2vPBn
gcIpu/jmQZInKp0pe9RQLpuwUZ2PrJrROgz/OLaTIA9kWa4spslB3Fga7w5ZmOjEAuFY+5tblEti
ek+4xAC0gW6CgPK/dQzZ6Yu2H9gJjb4+li1pucLeD/8MsgN1Nl9EucGVQy9hHl8ecUGhvdY3Vwgg
PVgfqq7j1QxwkGklUgFpRthA6yeGdYf1xmZbSqUoIWd0+DXaKx+wJCmJuajrcUeH1fGFqlqKK0Ah
OtVlRsR5pb4hvS5JbUm3UPPopMp9lyhvpTZr0iMWeZ8oo7o4VDSsPJQHgM/N3Soo2mAA0bFLHXj/
ROwxSH260ldAY5uGnZbxyx7w+X50If6mnwlDyX558kjeAOOUpsPFUrfBve+eXz3iI1CtXot6miyW
cwkNyNDF9VFJUWc+2XrL5uYG6GaZtIiW5pohITHmWVIN+ESjdrNxrITsy3keMcXISH3/UDC+x2ca
1zRaL4whV8BtG0rIGL9jJqKdq43SugKHMLUfobsUPXU7D9R7GJjBN7MpoX16HgUdLWIJUO7FE+VH
+YUthQHs8UUD44wmExuReGCHEuLmRLltY8clL6C/Vb8RMV+0R8jmec/7FauqvQM5M908+RfsDxox
NpAufrrP5MfQuZhIO80JP4pTpnwfdFyxYDkYz71OtX5jPOF8aR8hf6qzNbHrp5jyx9YQqPZiFC91
n4+yoFCVDVhK8nTdudzwKqvrg8owvS3j5kCNbr8nERCGjmifPhMcFN4N6EfIj+3aAYdSuZySrZ9v
6vuWTHw9WpmLaODyBAaiVcMFJgBmoxo3bWUoN++V/9GRGFTuLPHI6sInA+/2iDLAxKp4WjnsuoK3
BL2c9/fELNXAjeXDAkjf6LuPKtEnq9nTFPflxnt40PQHM1DHDwz1TjCbeSM4eS8naKIXEJt/hSsd
JrqbjQu00qzUKp5No53wJdYn8ysSYpVyVVjw18l2ReMs44srb1PErScC9vAIj3DX4/lYXPbgpx4q
FHYyt18bic3eenF4lWHaHTN/x49CjDcrzzxOK/mCGkvVZsn4gQ16EhyzV76A79rg/12XgVKZKZ87
83D8MPPRfo4M1NBhHvO1/4gBF91FVSTojDSKsTC7PxDhxXCFeVsfwvbQiMEU+lU4FDexuelzuIeJ
o3rZS3G91eQsZkV8/3035D5IQK/+xTDhJJ0YoQmNmyk1uoAJNA7WePiX2U4uu75BTySeR5u/WBqF
8jjyFWHjrVl2O5nyMwmfF7w0TQGZMw7B1oRUJTWC+YfZOnonbjUfNwbkUkTWaCfQ1A6aqJprWZec
1i2FTo5MU6UKoG3PJJwm6DXIMI38kiUuzWYCMJq91zr+QI/1jGxWuygFCTdDpZJdRusjKgDEJ2cv
GvKqM9l21GSq2eY/1JoOml4B1DT1KSjH9sZ8ZQhHr6ggqaqKB7F9jByroRQvmq3lZXH6XJFh6mcd
hx3vpoPdEFxUV5G6dYTHJaZwqCf64l77Te1z4xczW7/RjaK/OE1rts9jLG7R0BX+pno+2RymLZzi
+SSbC1+VXFfWeV0YEIfSn/Bya+CMJ+o3sYlp9yW4JNaDupRuvdX8YJnF8pwsQ5Lg8IPRrl4RFs05
Zjgo3J53AeE35k+Rp1f0Q66y/Oa+YYrqHEmzhqfrMTvwjPaTTo9HOLRghIXLw/QDSJlFkDiXxA4I
FHamxBuO4OG++PBCTvxGkoDuyM4vS8QpNYeqQ5gM0LBkbGD5x1A5VD+SQm5dWduiuoU43EJ/VJRm
/mMQU9G53RE/Yc9jQ+zzYmFQCJlVAW4pM9xn9ndmPlcRG92kirtUQdW9mBSe1TRgjKy6hdx2H2b9
LvZv4gRh9dxUre4WgBrZZsUP6PjhsgNCOJNjRsRVxTmA137Eziad1Q8q/EneocBl0OV0JAP+RRwV
O8FXgSLkBRLYXR902HXbV02emofLrGhhkvkkz7XKyrgBQ4kAJR+t04xiQnwwbpv6UVwwTrQYOX4v
7oFsST9k1K/O6Gi+McJ/WqLKvdoqkwErtiss++TnnrYPQIJw+B9HpSkwuzBe0kaqLyM+lbO4Zxxp
q9mU2L5FTGcgmdihpTGCVEP50jeTv7aIsbQJmjIbBnxsFrHVaQxABOhS/gj1zFbZg3m45nG/+5JU
wLHbeMoesXjg7dcuwvUTayejHnQGkm0ns9kqEFe4mxyCnEDbBnQid3M/rep+7Zkhs1AC20mh8lyc
kJVjjlw31WQC/1A6PwytSaKKqluC96sAGLwtsC1qiz7WKtb3p8DHtEASLbdl3Vg3CO8uSH0NmJPV
wuTSquL2dLur+YGtkUb5nUIcVPF7NfHY4t9rZYKXOj3NaQJGvPjnv+UDYMCkUIhSE5IM3U5KYUHs
ycWTJ2QRhnLmvZCT9JCpRQdRqqJo+JLGQp35vnDu9I0Rl3CeQS8fcdiurgnT9ordLyGbfxknwPqh
zC0u+WlHu4UqY+Lgy3wPGI+TKw2vqomXr6vzmP23T0TDiPHqrm84LCRKkk08hMuKce6SCP+0NbMk
KsBIU6lym8t/tHhQLrV3DsOc3HleQRMvrR0zHbBOPfuxuMG5ohC0YpyzVTVoQubOW/QF4v9zrU+5
GWjQ6hHDBs+Hg6ivi38XW8C+wysCXwF41tKn3PdrpwZya19CPSQDASXh4yME4pZKcFygqP0D2te8
Iw3lAZzU1zBQTJ3MWl/7tHJUm1daWAwPlOw7X1WnxdNB7BXykpYH7xNDmWXlVuV7fdfgmAPLP+DU
subh6VoIY1pT0WA2ly2YCHrpdpqCu2+yvMlm6Fc/R4A7WCVsohep8IuOKXzpXQEplLob2KuccHi5
PTWJ9/h8eeo+iNDPkpBjcPJWK6G63i9Lt1OiCpwlryPtjFGertl+XbWXJT6pcRiMo/PIFt0Y0gfI
fbI/8pwYNdSisJvvHu26XYtMlx5YdhwEJ0UzN2CO4eIlo7809fdYRNHgThFw22+CH2xNGlnRmRHV
JlzaSO2Ndj5oFywMPMh++Mox2V6Pmr8kyvIVjb/p87EgctAylT3Td92ElpwXptmHBGdi9360G9MR
pq4qOIIwG5ff3X8PdlpqUiwGqFlFwOeG0sYxbs8UekPsBAJPqkodz8WVhWAFDaQUzq25SHzKtLtf
jzui1Q4p1wTvYJ2k7Xmf5mMgA7PLy2vR/UGeJoThqzChMHJmyJwbC1hjKDkOaDB5I2ghOsVyQbR8
AQC0s+v7FPZHpEIWLP/EbsyNsLPVErSDTgHGeMjfTKdIsCG/OvJHNOz8+/rS2rdBMJf1pIwVt27W
tKtVcqzyOaclkxqsmTvzQEf3fuNiQ7khATP1ZGGpFratUmWj6pGDKTb/GHpKr/Yv53JoRvU73kDA
kryPDQTlW7ecXtLUzFuhrHbslZz7AJ0F6TmZXaHUy8nlryKvJJkYKUnCVjCf2x5vk+b72ALnGUJw
RyxuOtp/2tqeh6Pwpwo/4XtPAXOLLzMdrhwkG0USTPMpbynfoqpliMTxEO3eA3/iHn8xxUeIGqJx
4VNafcRuN1xXXMsnqljYx97hSMMTwyX2N4hl0hM3cQ/zVePp9bsAgzZGeAPdwqQsYfi9a6Zp1iTu
sD0y2sKVeo5FOagQSFMGs5p/5OiaJmKVJGxhQ8Hxb/klAY3ZJSO46dClmKEWFYq6HU3EXbdqdtNt
51Rbmz0UpTSsEP06Yn+6EKw8lXfKPdwCIVZN6N1ekpylgSE1NYymU3wV2d9URwejU43p79JgpOK7
Oksgci4uVOtcipteyQvKsuYHbZ7XjJJTlEdm7iUJ2/hsunTrn9+01ceUyptpRI8QM3PVU4CjJIV4
WSwjASFaZyk9bm7hEU8WOa18Wo+IhKsp53OSbNI=
`protect end_protected

