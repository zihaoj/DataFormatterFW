

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NXzbaqUbNopmRfuMl2HVT12kVWF2tapquWjA4XXIer8mi7ffCBnM7/NgFFiRNY3D2ryOG1Dct2dh
JpGD6YkBUw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hJtxAVssqqD+RGS64FGKHB0v+3PAzXPHwEqp73Yn3r+APiiq47f4Y30aTfVyU4q8KqIbivyZDgpI
INLoER/EdfKNKBRUCTLlZhYV4TFnipTNqHukfXO7fjMCxJWcAVhslfIqZMgchQ2jOgdjMPO8+ZS1
P/T6fOvCQuXBJUKPses=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rhdi3KcoP6AQydprYX6tjeWukpgDvF3B3GnijBS5iRt8y0JAyD/AtZKU7ELOfIy6zVHMKDwQnqR6
mfjIpeposjciWLOFJGvsZSdRr4REeXeRaL5ze6jFecFYr91/O52/k2GfitfFSDJrO7SseBFcgPJp
2uvHMErTv26sBO1UfM7Wd/Zb1XFFlNTX8matERVj0c0IFEb1gnFzu7EmFuPHCBEh88/YgzkXVbVZ
L7HA1KqWF+j0UtjnF0ule0XO2lL0RpPTGsCA53lsiCJ6zIyLtcs+YR46eFktLjPztjnIMBvUqk6n
O6GE/hBzFg9RLriyO+m38T67kmZW2I+9q/iJBA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J5zNxEoSPyQl2zDMrzPFTS3TdI1dTyIkSwcMyjgYCkJjzWXb/0B0ErwYjIDCRGLofR5O667y6lO6
hAruYy/x2xlf/RmIJP+8QR+mrsqyqTxvbCduvJ36gHrqAeRLcwhwUtn8KyeY/Ycn4vAiOBcGGWa4
UqvnluDmwMYM7/gMNVY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hkLyXHJhnwLBmJTFNR1wAOeuvKaAoxsu2JDlKAiil8QxNGEywbDolJyBlta+GtylyaaIDJYeU3IG
VHcCiVhVZjrJGpTEJ+ESvyo4i4XdytMiogaBpWNMrV8E9ddUNJLuzk+39DRkllAHcBnxSzIbZxOv
VyIAYpO6W3jM5ohjRWNmVXxi7DMP9g4BLHOcMspFDxJv+h5UiBIqcjEo9PO1N1FDY6z61/YFc/+C
5yvReJ/a29i+ryL0wRC/eQNnbceVccNPkhvXSstkZRFA2/e5qs6OUiEq+AQ17kAco3VtieF7PC6S
ftWFCui3wy2Z3aCxQMOpsEcE7qfn+R2zxkFyVA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6704)
`protect data_block
aUwQ3NdmwFcb5ahwwOGtDtIBHvtqLFjmk0SwKldWVjFcoqatE1oY5ob8IzkaEQyygbzT3nzDn7pp
394VSz3IUVpJLCLc3wPtQDKNWvpTbwgtUnW8gnfCn9eHoplMurcEclQDdZoZJjhIoEdT9pLGQXrF
owlfJSo6Qq+4E4lKh8ce0GeP2J4k79UJw6RIiIHLpF0Nlwp9jknH0odWS3JXlw7he3/TDBCxrd84
n5J96ARh9SdzF0sRkd+HBRWA/LyYDGKib3gwZTiwzeeI+gQsJ1tmGK6jwzGa4KBEztiJNAXs84hF
EFTLts3i0Z5r9ERyPjl+NJ/kDhRb9wyz7uECa6Lbc4FY26kvfIYUdR7tZtBqIwh3AloA4wNvPzVv
z0TMA3LRrKVtOLhdic3Pxo3kNHEV+qrKDBEiyobh++U7l9k66LLZZz27MVA3asGWvzd+tkLIMp8s
0UCoDxIKHE7KoQRMOHQzn+Bj8ShRXGS6mm69s3lLMFqAUc1E8kxPdYG9Q3G4qiPyCi28AHTr6EqV
BhqWdasPM0NEelWENUOM3lrMd0jDCCDHyE/IGS4TgCl8EUhrLx6EzG/ANs1HXliigzxDD3/H056G
OdLSHzns0Z64T6jtEfSzwMRxn3IGwpHoCnLc1buca+wmFgyquXaEs2Lk+LzncLEbjxawC2EI3SD5
mHoE3YmuTuCpSrkOwp3Lv9riHEz7TXi/Im4W61+u3gwpsbVakqpiNywBZ3NGgliz2Utjk6vwtp2N
/GXnWIdNwuwynN6gJ6h5PVva43pFH+8YrGukC1bop10vz0Iey+4n4pgDHKOSPA73f08LyKoz5EsL
6PkpwPVtRygYjwqAZ+UsE9qokNeI+0QtzK9GqIfx591QFdKEK3+M6nSDPGK+bT23Ud40hhF1ekqD
kH5bRSZMqO5VzQO8IY5Fm2qU+DQcp+598vf70Upsq2kORZ8nUR1/QOm8uk9Loz4mhsQIaJQxStR0
2fwl1qUNLnVdSirSf/7Hb0zNL/XFDw02ljZi5582Zzqli/x1APWk+bS0mdJIAwmt3oVGgIiIhp18
VouhAM8pxqvHSjzkExkFJDiEzAxTvaMhk8W5WUhmALGhle5Uv/+y+vVIDKPQ2dcr2K+ht9QNljzg
XQT+1qvpww2rIlWEDqJGL5NUD7CxVjZtz+QeYNAXPnIKNGV1WO0GKpfvdX//TC5qnkhcp/C79CeB
jtP53UYVnTCCTWd+lOrxm/oxDpmo64WzbQlK+FCLPYuUYPwFb8c3DFr8UNMk0WuO0pJ8RxQ+5suN
1DvgbVgqkMRv9/90ULsyzTHWF2p5N1riuyBoHpPSsrocfK+IrxuVwOruMjq1330+xbSMJt6jDMP0
DhG54nfQJkQ/Y1rtRQQV01t9HCMHg0AEiUFQdBS3fg5P/GObbiho8V73ckB2zm7o2sM0s5IUUDeN
19SiIC8sYfYOhbpoZvcoZNmu9F+BVrqcIPa40CaC+7RVwtyjxSpHN1Z7mNudMqq80tv01wOyQeVX
iUPNkGInMUcMpKvhoiFTtcRkg9UF3HH162IOalHHYXc/arNZaYT4Av5DlH63H7P5gWbUTRLlOV2l
f1d7Jolymg8XtiWXJC37AHcr5oF9WnSRh1DVGMdXxRBFpmQ1OpXUpUbMd5hjAmPOpx4c264zKdAg
RuH02WSX2pGMjexzgjhiDM+KhvV0nGHWyXtAY6TPByfLH350lgzbF3k4sGo/7PHM4XPv+VpJNXc8
DQPV+Y081QfY7B+dK1U1oe/do4eN5PRsslTUqZmjFHwB31adMc2xBI9Bn6ulrUZb170nAAoMVz0A
RFJDOw3mEpexqMHMk5ztOyvSIBN6lGrB7KLwX3HROwsmLlAp6GS1qvR8CbAy/V78epX4lj9yloXV
8af8foD83pji4LpH8D+U5fDKIz1BlRpRyYOshf3vz7Gx6/01tijtUkXwRVWHpy+brsSIncsShXAq
dJEE1x+1pDbyP7VXHhJseKagFhFPvmdEZwpA3hRe/op6/hjOypz/E0SBARwZVosK4nBYKFWux6s3
0Rl3dQlB/6083DL9W8LskogEkghqQHw+Q95nQwhrfpo9UXOs9asSkZSscnVfKVvdbyCZwRq4mWpD
s7UI6vFX98fT5ksCxcYw/XqX5rLBTSZGDaaOqBRIrNMSlShuCMs33idEKNymUNID/fPJyiJ6Uaww
ry92slHwvAg4CgGGUsSJBmfd8hjppqTfHIRPFD4/PMtF3V54fQj2OWCJ/HqqtF2vlylTRGKa6TdX
DFaXGeriOuUlAHEtPOMjCcr+P7kdeDSTGpgJeQZ4a6x/otxWVdKS37vRtFQJSuEnQtKEmSpbP+YF
kRGUmsKG47Wd2aWjAeJBHurYOAAftxGikM89hcV7SJ7Px6ryFcGPyK4g3LIvpSoF67T2CISCCaLT
CHbA2a3Jo+07B9qwrW5PB/+TEJMGDCnsgpLNSCV/uVUvPOSrqnC9la9BTTZIYbKCAnrtV7rJOm8Q
YcFc4BGSLQt+vcCJeHwE/Xgij0S9A+YWGLitI6uQXXqG5l96c5I6l7S9WI3UjffD19TbnFRf5ZGy
4DhZeIKP+wXSaaZcXF6SBdA9FrBJf6B9HXwRjbuOIGrdVp/U/JJYg1q/wEP51qto3GoXhkOi93bC
KHri29PIDMsGAg/tOz3P5inkV06vji7ShGHHlVF2OlT2eyRFFWDDOYYK6h52G8XItrTO/+YqoXRb
DiDcCWBc5JeBKxi1ZI3n5NvAZ90+K4lZtT1DOPebSSUHLVc4j+ueK8qZT8caNW6F1b68Ycu6AP+w
x1dj6ymKx/upsoGhia7zApxS44rWxKocXKJfocT4aQohiukFbRkI2ZV0M7+SbLkUalqzP7j8Qxdu
43UcoI5NASqY9uPaVHYZslQaevOCt82iq7GrDIyO+oD4eNikF17551yfNffzeFQhmmD8jPzE93ZM
BuPal/zPm5aaRfMIFhGfULCEU2NEyYeEqdexi1ZLVEiSIoJjlZdluS9DuMNPrJ60XQXBdrOOD3hT
ABna4TM5FHhj8oMxMaD26o3GCetSfiHQJFb/lsrpw9prkVquGZJUoM8fl/rF9ZXQxFKnRfSpGOLE
jasWtQeKo0zBS0xTYIotJyIPMDl+AV5a2II23OQ9wYzzjiy2aVuWUD0q9mqEW6wKWd8UXhSL5++p
HGmttOwSA8gogyisN2WJrhs1EHkP5R2CkEUYlnH4N0WNbuMfxmV3gpVT6BcCi9m0th/Sopue57vf
mesj8gO4IueeqWHpHZvS2GNcix8w8qR1eFCNrbWwcKE+YAnuTHxh+Wg+ofZcAdBsg/0Fv6X7BwdO
x0pDFp53EexvI84Sh/IQNEZfgEgreu6K/iXaneYEk6h8KyYUUXtV/KN6fwRjU7jMxgNnqRu8emcR
JQr1j27skbz9+oCYcj6VkDL+SkkkYkBPHqe+/CHC8nuUaB5dZeknsZBTtCewA0iFJZUo7g7MYGTw
VKTyQsasMqGprvephSROhWK3kyhQL8CMV46mrQpf5mAk22lx91SGoYOxVHGRd3bN1JXCWlce+GLW
CgvZRNrxRyVgrZXFosO8RoqFoCSmK4V2jvqRxxBF3phBVJ18Ws1Uszv1OxNyBpzIYuXS54inuYK2
iKAOXRUnr6YQtNRQ5IiPYI/ErYaLLf1NjmkCsWgBYWuQbwp69t1dCBlZyCcuysGosjeTrvFaaoY0
nJLlolqhmGZfmwHaHjsCD3EXY4AuzDPjg0vQZNacV/xQ9X7XVVmeqpgu0gmQVBtwl7SSBaJXuSvj
COgdbca8S71/33avMav8hvB2GQMdcZlPH1UqOfpJ1VaPSkF9C9VcoiAC9OpARCgt8J69GEeH0f99
cPZe18tUJlXqFLLOhv/K7Sup7Y5/GEFYXWEW/kS+Lt4qJisbsT4bMiOwfK1kW6U6OWNHaO21JDi9
FvNd1hhgy0pa1KdeyLdK3eKFrkokhhWBqhjl7pT8kUsBQTcRQHlOm/4GjwADPk5xs6OO/Qdt3J5w
SImcrr/xFI42tjtDD897mRLJ1BzjBkPgUj9GIUBVyDrwOF5tJyetHY1j78dlZK7xx79NwKnVuVxr
8vkVLtj3i105Loul+ADuGLOmYZexADyxvXGB12Zyco35t5VrxNBrqYBrF3QxK3RqvACtSXQCadZz
0GN5CjH/4WNJcQYNK1HLBsEdIoBpBAw61bsihNfqZ8y35fsn2SEGZzCPJ6t7Vg5o7VcmVjpBaXZB
qPodR8gAqCewpLn9opfzsdQYooskt3yoHRW0qLZ/0dalvxMtHlBT+vXXO6cgLYrAFyBvbAplmr0D
R4Cj//vL8Mv4BjGcXzBR3spPiwSLhR+ho8YfcmU/v4qpfKKQOhcEwaQQArEbRMycFB7oKtyVfOg4
OqEarDNM3fRlFDZoXj0hJE0cKnT3IGFks64B5CDQ13zHKeTdDzWNT4SOdNB48gAFuvWafXTaNHQG
X09Josr0E3w8lv1yYadEUTz0KbQcuXKCGu1HsJ7BdVR1gz9wTjS9gOi609NnvWbZT83i7joOeuB9
Sixg6c+71P3VCiaGW6jImf9t4Y/W+ONGXUrETEeMwFPcRzppdQX4eFLsNzpmgZdGw09F9vDMm1pb
5O1BZ1FnSNscNE27Ltmo7m5cHObEBGEZhRxywEod63qWiHu0OwZ+PyrWwGP51MGbh9F1APkBHfM/
xoT8jrKE6EpMV0g6N4RMqgKkw60Gq/34C2UH0+fc4vYZGiGuImU2Mtp+TvHcxCZKjlxO4rVFALC8
qLeo1ATa8YuaWuz22861ZruynX5MuNYb/3D+joIyTJnfpN+vKF0xJaZWiF0xMW0Xjt+2e49lQ5Cq
hUX5AzgfMLWNOLevVlCNfw5VLJ8PhMcHlF8TjiDmsmPYp+oEzSEJw434x0m0Tp03sYjVVvl3zJTA
2tqrwGRGk63pndwYR5ncwOaq1chaO6qO6yt61k4aMQMd14+s11S5g371yZBlvFLvYRDqpbdI4TG9
QiOQI/nXY6sTD/SP7g9+pySEcg5pzlZzEy4RlfI7YnUHYO4y7eFO8xnv0oOwfIJ6sKT+/me1tRcs
AGy5TAHgjJTDlh4bOT0rNZ96LQaqvhx9s/Jke5cLFxMzkJdQ0TnwLQjxiZYbpMRIj7sScN1SdDzt
Uc0yWApJFklOxBfoXL6L7V9uzkZsHqVbC4v4ytBe5zNvHV18GctWVO+6l31a7E4ocoAHUtW50RX0
pURBGgo/zU3k0ZpDakHFix9QOTIj+k1unVipn8fktbWuKCYSli3rLUegFMo+nlrVU91rrkhqfb9K
NTDdfCMfFE1eLBERKAbCSAlyAVYDTeNSsFf6qEj0aimNwH+r+qH6fsk3dc1W0rCRDK9SmgtAGsxH
DCBNEVtHIIN99VFv3acXw/g9VEWMhbyULBy2HdMCHh9eHzH2nSXxPSphD6lteyjOb11ZqfVH2gpu
bkMYCZPDd5ZAE8GgKgbkk/krVK0QdHF1uiFG4uhZtsPkJwDO7bFx/WRXcyHXAGBQGqVbz1vbgxiX
IPWszGiV4CdykkDMuESA2gCJzy052QmQOiEfTdWSOwzgB7Okm5Rl0bHVSaVWHlllN1BjvNY3ej1s
eGKiDRB0Atbo/VC3ESrlfYSe6B6X3juH+15m5upg6/Y/o0Y94S1UYGztJVl30WfwXZjZNKFYpyOA
zVmjekH2xhEro/DCoJp4k4XYupiR8Yu6zGNNNCx3aJQbumLnEIJSckuNTGixH0iPSYLSk/BbZm3G
Rn6ZWCnVxmN9NQKMfJOEBt0iy/oxZZajtfyKWmTukbtU+FUzLR95Kd35cNhYOh+/iJDVsg+2WKOO
fCV/oQdKXqNIjLJuO3l478kxSWzIYZ3RTce3sYb9tosdaoKmxgSObiiGEyosF81Xog70k+/rstsR
6Y6NL/PxdutnHSyx1xDgu9JRoUG/feLhpVpUpzpsNJBEOFQo+6c+QhGL4/TxnIwaksJlqBY05SDj
c1wMyVjtohqSQIf/Bix+OBnWKYAX/1nWFv0XS2sXTt5Pnz73FO8XVtdgRzBzI5mOL5pPExJpwqG+
afwTAjxUJd3oe4V4lO7PJDpT67ECgR1REZBfSnA58tnveqJlYGpirVp/UuEIsfg96IB48kFHV3Ch
1y4YVdw9h2O3Gyv20E4NwmI/VkP2ZEyBWciOn3ZjlFQogl2QwHgs73MCpBqJ3+G9S/iPtNDcFLPd
qWEj5Y7Gi+SSROtSEMQu7XK0V+nQ/VdvmDrirY4RA9QKBflzSKPG1tHDTPzAA3VTA4TLGq41KsrT
NA1qhYEjMec8NvpB4EXtlbhJfCd02vHIVvg3YTS6l3ewWktCI8hoT+yMFM+bAG0JlqOZTn/1DYuG
VFCcmCEPlNcFsWNdLrj8uPB/h3jW2RPLjUfKGfinynNKKgrbOO6VQC/Lr4e4DjjNkHQ1L9ukCAhx
7KLuDuRHM6HtMGTBCHyih34tsj00IONBXBbX6pDgYhlCyrmTWwJZmCwaWRuNMjFj6dMX5/9pIIGz
pE/K8kvzfJNJWIaVISkg/3QlylTf3RtqXgKx+XABDtoHCstlve4g4tLabAqrqt0DRfMxoJHZ3EPl
q3+cI5wc4Kj3EoKUZHYru7fxFxCiPFPadt2bG7AHZdsYmCTADZ44bKZ8HqbKztjDVUShcNHhxOqw
t1SDE/aOmBhaPY0kbXm90vXX4CXIkMoBryVahKEsWiUkdDqDXHgaee5SrFzOuwlWT46IWlezF5aQ
mlQaieid5SmilhBxOMYuKWQILpS9EZ/mEjmlPPda7aOOJMeMGFUe3Ja8ybWG3011aTtizcku3GqE
zuRMtmEjsThENEWBnYXjoqMu2xtuoNDHGLNQUaxj77pgXPUd/5u3SOdzwvFbkGU1M3DqhFGwVJ3e
jXzUUwEbB7K+eRZWFihnF9D7y6oy0BkJt8qyNTCoeIbnuYxeNJJEOK442pve/IEgnS3UFiWP8k48
SX4/6bGXQLOcaushvQYfYllU9yc/yGfPd/yV5DRmRFfxxE84fD3DYHwg4oBjcyyUsV27X0j8i8hW
Ad8QvfQh8MItpAW1oDiaJuegMTEQ0PMdiJ/obAoHCHUQhmjnNJbyC9G1yAj1pCyWc9X6qg1/TjK3
zidf3PB8IV06kFtQo2DmB0uA23KLqnpuy+ypUIMyxQIkX9QBCUrilT9x5AkQrwkx90nSbBSTDH0s
TH4OZyRH/i6fnqizWHdUVHBMgitqtfb8Q4um0V4tNcwya6ZMXo1Fj+GHugnGQd356Wc5xOW/3CpF
iB/yOVn1rjbr8odRgXRRa9WR3cVn65X22eUTtfVYaJUK2up5YZfJogsLPMzPtbdQu2sUDWxymDTO
7Uqa2YZURLgH/bt2rmXJpv/F3MJWgXa92+oYa/7EyYhI7cHfF3ffyM/mHfOEWzVO0nvV4Xe4EEwA
scLL+wYVLi/YIDJx5ZHCDc1jaUQbs3Bz6KUYVHKBNEY+00JV7hegmMRAPCx95HR/ybrSwSFA5P7V
H4N2mDEdfNYO3C5A0UOOLjSVcKLq44x7rCPJ6D/v8T8f0/HKcNOREATyxza/8iSEG+v/d58jl0wC
rrQqqB3s0ubYssBfOgs4xE47/Ck6aOABig8zQ/5hoVXvByicpAGGHDgGXUPLf79/HIwN8UgcG0Bh
G/uuXGcqR+Gnv7z3xjiXB0O4YUnJKl7eWjl574kbRjL8OlcoTLHMDSHULNBp4jcePTHnFLTILZ/Z
fa0eVaLmn141C8yLrcmdd9a8MR9BPc3QgPgYMFN8UXdhaFnjapJDtUsDf/uUabqAnRM9RNcTT6ix
QN9avZ7J9l/M5CnHjzle+NyrPnsMzfXsIH0WEyfYez/1kNOLVJHdmGA8ITfg2sKadVbvzJj9xitp
Eaq4ylF+nkUBPyJniDrNtPYB9nnhEf3PK43MSFTKJmFiOj+01rShGDwjLYQE2shkFMktgT0/QNWZ
nVPzO9K3LMk4aUde9Rudsmu5lnWVTlMRJLuxrCC+5heW75ldIgo+NtDV8m1Hwe1LCo39ZWbkiF0P
Nng8L3fDrjlAhbwEPQR+urL+lbCMhajTKOTxWfUudGoThnTU7vyp2u+AbnncEto4YJxT9rM/0RYo
Qf03tFAj0su2RFwjSYiRhenbf8i9lZxUAmVPcAvvofQJQktK8EK46VbUEHOiNsQEO2AkSwH79FL1
JNXc+EZJoOWYbfTPfr1Jg1aQQOjdm1c5zNLeuwUhKnQF33/LPd5RqHA8cSLAV81CHH8LSu/I6ges
Lf4R3WjYdw7dqwEI20A4ufFvk1ubVtx3niq34fQJOV0kTWZMhojg+TOWkoaYqWj3g5kHsKipPPwp
GTmjXYNz9aqGK9dFzYSx44B8NoLlRKTDGiOYH/Lk+ha6HF1A1+WnNIsk6hTsyBhmAAO5YjyDwYYo
Ruhh/BKDLh+1b9QsteOIz5fN+g2WBYjO58lOh4z71NoOx+ob8AQ/3MGUJG7X6Rk8httWItX8tLTh
WcwH7J0M2KoCkoxOOAZytwMk8zD80XHSJ2VNIf040/1h4Vl6QT826/QYTyALnQss5XGg9gmtIUdj
SIQI/K77a0SvR793MyMkOzR9rjn8NTnTl2n/lX+XnYFnlLI92zBEkSy+7bni5FiO4xGw5m6mHfiE
MMpl24wAeSsG76Wdixj8V53/LnPz+J81TJiG/CfBmLtzHn3mRaRxpu0GWUmdt2SFx/YhB5RzMmYS
GKjPXur72RB8BxWQk5AJHiLEc0WR1mxpOK75yb0TpchVpQXyetYkP4v8q6Y9k6GWQaz40hvswfI/
fF+bWhz2A6neKHylqe3r3TO6e7Ti2ZLXFhSs1SidIkfDSH99Ry3b9PHmJ2ERB8m3fjt02guMQsBV
gX1SST+DhTMiXXj8/qSk79qafxseEMAw1drVPoHvDDOky5s=
`protect end_protected

