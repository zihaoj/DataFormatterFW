

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AQtwTyGLz0NMO7LyR9Lhuv2cA/4y5ZLMBit+QBleYFW8IhTeXqKPD4aSeseNMhUuoCyqQPHKXbmX
LeVqKxvarw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hGVhv3AqeDsw7H+uancFjD279XefBZ3mwEBxW5pFk8a3sVNt7IAIfyXMtmp6XBWsae0N+Ci3/npB
3SasZ2GaBZBVMxZwKr7R+ZnX6uwtyrN2AJndaqNaMftiUp9xtV76bCQ9uH42U+M2x7hR4dtD0fvB
LYvzs92V+0bNZbbueyA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Rwsa6WOnTwbkSOakIUUGDzVbehno+eVI6KtkIdY5kK8lPoN8q0Kbk8vzYaFYPqtx24HeGf2fCrmL
UEBJpMMEdeDUWeTdVGVDGgJQqfSETdgcbKy251IhCrCQqWqIbqijbXpSb31jgoi6iOsGmyPpR2m6
gAug5BKSALEa3o/asLI95p58SZhkaUpFyJnRspVoLL7h+r+QTO86y/MjL1M2HHbiMVbK85YFLHSo
hReZLGxbL6QQS1znPiQyyVy1PkLupBaKBDXojs4pIX8/CiwzGsFTCtFrmYLQ0UqfaMo1P+9NS07F
kOR3KwphHArLEZjIth7K0OygkOWzpexPymT/LQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GFpv4P68gj6yK06WrGFskDzgRibsxHI5jWrB5NNgR5jAhsQi6zUtxk9D39KKYeNXJovsaANReMqt
hhf/9kQFTUB17gOOYbYVuZ5Jw0U+jkdJ3RB0GtDnyrRDOZ5DC6YyDUkB2r6PLs+CT20zanhxcEtl
sQKOEnL6phaWOedi7es=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c6+3pMI4bZ2mi2A6Ycj7+UeOiarlb+GAsf/fjV00iWC1qCUggxIKRxP+eJ3z6XT4BZPrG1RsEhpx
pNg3X+Fuqp0RwnM/yLWB2Ltk447QmP19vCUIvCHgqjPtI7kt0WbjsDqel6aoZNnpmEL/7gd6/3NS
nhA3XQ5QMumSsq/7bmoNg9hBobg7U7jlCr+9ZUf82X7MkdUEYGN/bzCmelYTt68FJ8ZlCW3h4ve+
YiX/yE5WOCAsimsuL0TKSZhntBGdjxuGpkF0yYXDh6gl9KfRWWkqdZXIh2qUMADKH/9YGGslBS9G
GFME+3dogZLUU37G226tsYdPFlDiwh9fU/p8oQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14368)
`protect data_block
ndbh0QJbQR5DRd4rlOC4xajWsTbjmiYXrdtsTFl8IahhsGd4bKxPzkHNTGYQQjGqJ/9WmLcEQYYt
7haWsjLCA6qqvapS6/ONK+eTyFfNGOnwXeZZDQe/AGDTkxKDlkG0Dmc3Hje0BLptHoUu39aR9vh4
MOruo+C0++ph8D2x6qdk20FRPY3SZe/k+2oa2/4fC4wMeN8soGxPOmVrYPBKUwh9pcOCrE9kR2WY
oXDA82geyA4AVWs7UlY9CMGNLmyvOWA4tE30m5yxqWJ3LJxqiHanDiFY6G/6n0H4EwvJ6CX7t/O0
DqfnGZKqhh07CjfdmpwYJeazdd3C9y0E1qr18nXQ1TRsEvIQNdVQylCN4cWYwwZ2iHw/MPhNddZ3
ZJvxAclJSzP9Bqx+vNlOBpU/gCrp0pll04ifUm91tDcZc9KTo76ThVTLmugo3xf6ykIMUoFQGm4b
JBE0o4BVS98+XqaJMB0D5zSZxTXXD7Vq55YbUNyMbGoPcW950bEvtQHamSdbKlQjNGK7JmY5nkox
hiyqYWB1qUpRnKuAQ6b5+G6OPJtwp5t4KVj+FethEh6ORYGJfu7nzwqUlR+St5TvbUgU1dRzpwFc
yj2cO7M6A5slx3GZcq8nEGyZ3FZMV960fuszecTzFHAEqckcVbO1/Qm+w1l+c/8xU9uWIwMGB4lU
z9ct93KMZeZ5GwFrE9EVwdcZSR/C31VF67qVj3NBGS6w1F0omcQYkO+A+8sZImsYNVASYci301RR
Le6TQmFFVYOMxFDQ5f+Nkp7HqZZen2A2yYS5jad9lgY2A2arcDouGKnClW3Xqh27Zcw2ReMupXfQ
8iijThTSq1QXSIml6L4Xf4brT2AEQVlXhHTWBGWtPq9u81vM79zQJA29LWCSZ/qwa1Vq7bmhbGJ8
ce2aDLk81uaY1qvUeOkcuNUtfLsowhGdR6ypjSS3qlRzCBxkexEmyBODARYabcUCm1xm8YVxu3bx
rk299YFBkY83k29l0rgVFqGpc70nb3EgDgbSug0pztcgrG9OGORkwF3nUpUAPSSoG4qenNYSCj/x
N5d0uV6hWw5hU7izkJHDAXRLZrpd5RuefTk2Ym4iHX0BLXiPsSWjADiyyOYI7lYfjx8lbzofnB2S
srypC/8fi8Q4JxD2ivh+NxKTJI2mnOWHascfhdTS1IDmbdmBSG/IvkLgqclIb/JDd+PMYvZff2P2
fPKvbiFqspfZL4BdFyXX8qq+e18V5kDMtqko8XW0hfUSa+TMzsy3mga3q8JOMGTuHlwLWckx9+PH
vwKwrPYa+oTP0DdnSd4XsVNH+ytb0KbYE1fLcc9BgbBlhkLwrH33qrXEXWuqp/kb1ry8UAgXdcAT
0MDfR4hHoc92lbF73RYJNV76bnoPgLlgOC+icA4Nuwo0WYZXNJ0H/a71bo1n0PKzDJkLS5FkcR3k
ySmHwoYNaI/r3lJ7aHn0wq2fQKc1jHTewv7Ydu8s2PPOGrYtZ6nwM6kHIQUzSKee/bGHKYYLC8C1
q0IUNkBGErGouhNBSo63iONZCNg7K98/qqlmhKI/dGw/QXN+sCaf6nQoaOAFsY2Q4G/ToBW06eKf
v3II9zVo+sJ/65jcr8XQNwima4zUuzmMsbKTS5Z6Vmlr9V1xNk+opsTI1b8Ku0IXzE06VDzyU6Lz
MvbIN3bffmaV+994OcZonla6pk57qM2Zp1QjDW6/fYcP/rlT303oELWp1LOZ3l9234Nxzwim9ths
d3O7zi6sqr4Dx/yFwZPpVxeTlgeniyloZVjIWKWYjX2sUtH80M4FgvpgTgFOehUK9y/GQKenvv41
9ye89IEjRzWg1+UkyGRA3cN0MdDpaPRLsk8Oe/nXIRSUClzCfdG8KqjLNGCEthgtXvkg8NimOL1/
duixwYjD2vwv9A6ZmivfEL4JEY9OKgXZZc+rqXMwCI5z8V/b3N9jlK98J4pztsjsNSvjRw1q6AtY
jKtEXlirdOl77g6AuoN7Sc+AVham+S/ozgtAyg9hdggXV2RgAdVpZEnZr5DAh/Lx1ZnPtQS0sUye
VRIzatAB6M9ks6gg64XiIPFYIMiL9TgZL/AaDDm7vkzjfjlWf3kgo632vSRn36GSNdw8BelwYOhA
zaeqU5riMhuJNQzOTE3gxUawNsWfXHE/j+Udi2KcXTzyL07wGA7Qb2CN4IlEKeg/pbuG3KaFooJU
5Ac2LnDv/4S0mCVG3n+d7EOPfogHBGfHN0v6AmhyzuqvflLJ+ILw6xLS9RHOHKW2EX60KxWHxN8z
PftaSoJBQpSSDSVWeok0sAkZpgM2EXGMCysHTvzj6TN8VEqD4DviefInkbsZBBEyLmrebpQ+5YST
541O4DHxh91S7bIrsBPSrbH2QMSHcAk/cB9axUa88UsG6prlKyjduAjkDOeJgpDdon0IK4UHwEaR
5GzocNdpbuQguUyiFMZ6HR9YLFT3nVHJh8wv615ry6IKhfOKzLpqZk3bLM68N6cV5vCFxzf/cEor
5671cyOg5XSpbzTEomv5rllMbXhIclcpQxWk00DDPGJ+N72y0Kid5Yg8SDqsWV4JayerRhXmJlcg
YxdUeeoq4DBEyd2fiJg+kzOr7YBjE/MgXlV2UMdFxLBPGE6zmwSsmbu0mFlVx4VyMYzelSuzAXm/
e3G4JRlWPc+5CLzxVesyqsg2N/pS3jfBfK/42FBwc4mWs1/MTdDHKnx/ZvR9oX+BxuboblT9ofHL
dtSv+24D7uYmRvp/lq/CHjgbo7pLFRX+bN6kjh7AXvS/IJZHZd98JcDztQUXsIj5WRhpP+aIIv0a
Ph5StL/xWk0xi6ypycBvRDgboZtWRKPtZLG4SGUJ6ZSe+F/SVBeIDpiExQ4Mft+0h6wmtimmh+PB
lPzCEm2n8yq2z0Be9mTv/zZ97Xl5R5wmovoVl9dEiHS7DVVcAgeZJTygmWj3lKv7gGTQPplY9Bxn
8FhvmL9lL2kvG57W29qX9gPXs7T4cqlj+lusl8hfjfw68zx6/utWLWJdiq/1kK8OzjsfbxdxhswK
6IHzS+egClq1vrKLfwoZahMB5jiaJeETzUkrmzRAfr6OimCYAAO/AbXJKAhBixy/SwHncbed0QR+
gynHYDlKGEM51BnLUHd4JqxklaeJUtabtfAzyU+WQ//4UOHGNMR7v67dOBLsk8Pkck1x/Zw+aFMM
mPdIiOmwxP7w0QFxfvyy2oEWVsuFuPPFpMUxVWe4Q6vj5/5eqn9ToUbw+RNACzeW3hmMhyj4qAeT
z6Q4sY5/AAsJeFb52qE6oBc5026CgL/cxMCf8l1sGMN80zt0ld5fDcbEG51Ihhih0HZ4yDhggsmd
WQ0QYI6ohNrPKYH8Yg+ju7G3O5g2IfzSbcAUtQ1Bwm3+wiyon0/ffFwMmBOYgljHxayXIcdsDagL
xzY8X+LZizhILRoRbcofRA9KPdzJwnttoV+aWJCyekRdZbyucrGPMhZ9HnlufEnnniOe4nEeOCxp
wg0POMXGbtG7Hzi50/2u8qkW4wY1XG4kfD7LdxJreTm8STMH08CyLXbVgNlG70JkfxMrTwYo5/TT
KfHyx7l/8b/TQSWurx4DHozRhDMHEh235noxb/kBrJP/n1dcOfSTB2JJ543OYjQLufrxFv0qTP+0
O2o5WVfbNJ43djFTwoX4q+NSEVo4YKfUkzAH1MgrX0DOkM+ZqDoH1XWxJFoPzXXXbYMP2G2yakyG
1QBklQl7clDF/xWVH27J/CDLR6iYQSveBM6fzui3Mh5QC0raSUWn5eLHuDCCvNr65ozUqbwpBWlE
kVRAOSlIU6RHN7wm0vMLLtRdk2AtwM7yhjz6JIrtP6hb4hhMK5yDPW0gAU9TKWvukikfLLrcGb8q
X5wtbcss9fHVwv3obRwj4icCCFFTusO4dVQ+IPwBna+iPANrE9P3huOrrnZ8iGGbWmefu1q7bFl/
YjayIYCjrz7hpcoWucok9hGT9WPW9KPA7ZTiUHgKooAFtMICd5xP/AmLhATXGZHt/F1jtmOnjsDJ
J2NxWi42/5NcKT0a08eU5nsYMC2YtlSiqN1cMVqY7daA+W8E/9ofJxNOJs0CoO3WzuMpI21bl+Hf
SKi5OVLyvnIiA2l4Rcga9xCIA7hTRZnflmbNtnd0rygWHN+urjliVDzsaD+qitkwHlzkhEaTgvr9
rBWXSvMHDvut8vvJneNeQJgfJ6nxGW4an953yDcvDV4vUK9KknIORaYLDbD2nqUVnNuZplxWJ3gE
ugTPtGrswHnfqjHnwbjo3WkUx5G166StW0pmELSdlfZNV6Sa/POhAAWlwinfL9h+kHPXMasRwdw9
vnPaK1EhotMchumgmapXSvOS8UUrOs5eqTv2f2G0xA1Ln0dfZbDL3MCYruLQFmNmefVBYm8kPZMN
RbvlKEk/8rMiDx5DZJEceIBxgLyB4pq29e/PRde+U4SRCeu6gft+UROzbvvISNl9vS3MxNKP1ylw
p84GcOa38Gj+0oWO4ExZQ6OV0SFtVbKOvYlJSWLRk+bYHwZ3uWgg4njw7UcveDI8HKTyGR+Lip0I
IzFMK7Vs5ItTGwjoDh0FA9jczFUZ8oaPbkTpmn6BhFDqOEal6VanXTlr18B1XgAQT8B0k2S8vGhn
ws6ZFDfAgu1O5DXpnInnWvXBa819GV6/tQI0FHAKtufdbKhf3/XdTFGs6eWG4YYlo9btR8Jv3u/e
8/KYuKvcPexHgKreEvxwUMtyYYyShsl2oK9Cie1PP2t80mbrn/AHZSxJVsJMSQtC7vlsPxZqqYvj
MPbXS79ZHUM+0+85JIomm72FrFEEnFdS1Ctj959LvXtc7inQylkhQAcjFM0g5/28WMtIwrnRqh0E
0P798YPLw141eIeJ99i+S7PMyrAjviyX+//wyyJFF7gO+M5glmBLqwxXyisXbEv5NRg3KWGNRrY7
9O6263qvXd9jg0nsTkNpJAOk7vubVH3yCd6CHQiS2m5oUx00SXu8pnw+6EJ/hHQojkUF7RmdS0aW
0RA7Ifn8Co36snarCpl7DrO4aJSYMLzHu3/cflwCEngnhyLRoWdZJ899uro9XEKLeLImbpRSzOgW
MXVEXbCWZ4nQMBjCXlov5ULetFbYwLF+qNFVNj0q+oWqLAYZQR/Lt/tvNtv6EAJ2SJF6LknvBilZ
x4koH2ehDcoHxwInU6KugjZPju2w+3qM9rBmqHDVvY07bPDREeSAbeHlSPfdBtiiRrKCzZVL342F
plIJP4Qr7jQVKq/XNy3hkuK/c4rRUHHQzt1KLT6mQr+IF/BAe9vro9ac8BJ/tvzIRi5TVrmB9R2B
8TgQZeJGb1btD+GsXHgMGfk2sfGrp8HkY0VSzsETMi8hropEUB+Id+VnrQ0dpFnwKW7j16oIG2od
niLGkI6ST5woxzqKkZiUYlzf0UkInKyHId9NQgh5xeUX52lpYRakXkgePchbYjS4YzYRXj4lhiEC
V4M3aCHTI28zC7YP8GetXUb1FZosTN9mYzdyIcYFW/ws/wJs9hqQRxr9ieR/9tYK2h+rehUoJjks
qicQg0sitEbotbNJl4s08hDcSbF/hrKZE7HzwosLbYqFLAYFy6y0WPT9QB+WSYbjuq3Vj3NW6yJz
UNKYuCT69vW57L393fyGqV3yt6ifmS07jC6MKfaT1JnsAIH99JXsei3+Xrc1ySY2oRBSlA+XgzEx
Nqa40lXjC7JWnhUqMJ0CbeJKjpUljoX2ecSZocdloSymC8CINukTK17x8I/RbsDgvXVbn5Huyag3
71DRohEDhLLamuAO8EsfF737lzsyafHPOYMO2SC9jBRtDPgHp+b3wJRsCBRxPvIHwsNJ1GJAA0ht
mSw4MzMgAM7J8yyn+VQuDWCPg1cdsYI66umeDoNepLqKehPy+G/BY/AvtF+npLlQTt7MK09wcctE
8Mlv4Bs2JhLWSBIvPqwCM3b2TEzDB4mOFhgB+fmnYKgmfqUOTtH5XQSnPJRSNbjADz3Sk0/VQ/lD
RYHpkOyoTvjyAiXJB7KP0WK3OsOcGhOcWiecdU++vHmAdhtm4nTha5qO6iTCack6fd9+e6U98V7E
hD7n8D/UissBtewA4X5PL6rwn9UulO0b2wbHsXptBJVkiCjdimXcmw9obKUTdom+aTT08OH/7MTa
sqqiCJcH6EMNenwIGm5ZhhhRFhcBRg04wupQ7vSLbAQKXrbeU/8tWMuynxFZbAkSM9mpWlG+SjaS
rEM0wpaOjF9LPGL5b2dWte1kVv4Hlc6H7n1uLR5Ln6qLaZUYnxrAFsw4SWOhCx04FAXyTBWbDY+p
AAYj1chlJHGDJa+lT4bdVVYSULqpUnYpTztRB0Liz/KfKpyJk97/dimAW2gATwXz69P2xdXVI4WN
r+DlrhRs2YKGsIiPE27DT1ZoGyDFG5+aDGqTeUGBGvWtL7kk39REyQ7CwbXV9BouW79Do9WDQgw+
9izR7llPAiCZ3wuyqjIvvCdbTleZ/R21CBde7CwU2GJF8QLRSqSfP86cXmGTf7NLc2YH3yjUNJsf
LhSJ2lOWL4+ZaSsIrNTtsxtqTuRo8vhdkG1lz1dRjBv2jCxKHdTcWvzCp4c/6NAWoamOVaaQXm3g
ITFEfhR+7krzuObadlV9lTc4O2/KRozrGbYwuEonIVz1YymTbxiOB8IcMKf6AJnjR6E/x/DCgLIH
C+ZcP8oGCjHsUwyo9A+7OzOCaNJeR7axlzhnEk5wERD6cM3QMYC0CzF1WewQKb9zGXrMxS/uORyV
LC+Vy7iA1SOLSmV7Gab98qn5lpxYF6n8fykZl4N/GTChXi2g1T5R1FqCIyeqSLjLtGuJMHsk5t/W
0dPRoZxKNsrcvfYllE1gVG36ePY5wGmu0QfJVLtSiOmnCmzMXMzX3ZccrpQJ7cC3EXhnWq5ptUpW
vwRk12XetqnKABHW1LUWmykvNkzZDZV3fakjEeeJvNqyBtz4WsqMVWD2JnYR9nyq4zCEFvE2Tx4m
Af1VrwGQj2XSgUNuBtUg+8/1J1guM7AyieJQzOiMRNnayH/VzmJGxH8Vr35sjbfaPVzDybP0I5tW
g3oYO0fl7jiPFy6FH5bBeDwIUcZ1UUlSLGOTscYi1X6374GrdYpPYoC9G1fNjDwOamLUa8f4XX79
XFMUV2j92K6bXe1iN1b2Ht7myW0jes4sdviGhtz9oYmdv4Q0NUklx6WaUmB9EfMAJw4qB2+36tV2
VxQioIaG9sWtohlflVdNt49kdc/sasAzRWOevK5NbMHL+EKd1FzBvrM+pi57UsoOwLRQfESHFPoy
FwnLfPePCSs07WDrHcEaZpotwRmjMExg3tpsm4BbpJIHXaadaR2jmZ1w5md5rGXmh7a5rZB3MNdU
H/WmXRZgld5FKQsQcZRchcd+PsbWdk8QpsdRLTqWYcJMeomsniTshFsimLFHH01soMUsH6+cOFPP
0T+8xQNiS1wwgt7NuQXHEENjZettxSCYzbkvnXpY6QBs1TvA1/qzYr0W+7w+8P5ncVtHg8ynOwzz
J5tWEjyi4+Q1p6yauhYZl4kafnr5e7Iu2ZjTLnmHzKYpe3tR9OSqs5s8+39Hplv4sd87ayYoHio9
qFf7AzHrxagBqNirFDaHYO9J4lFx59ovEdj4oPa0y1t7+246gl1gGjXIRBqRYNvCV5LZ4wgWYC1y
SeHs1cB1bF+KW/mZL+WAA7OlLkhleSMzwb8TBGGX2JEJxPFJhXCQmdu3xzasGIeiweXnDetLDg7S
YUPLg3agR6qPwN8b/Th9OfZDc3JnsZnVIGYrikSAVsFsctp4qlmaedeyppqiBoB3KMVWMhWeAh++
aplLWojszMbOCLMfdjZvehaUwH1N+rU3KWwLU3N+VJheaXdwyF6uew7ZYYsaeVtlltshRfmI6dzd
CJujwe5WTeCj/cpFA1AX14PEHEEDkZiFzEhVpPeKP/bYl+oOlBDD9znd7lQBc7r8qo3oiymMzTGr
3PneiYpvoXXt4qa6tIMuY9MmqwsZ9bnuW4nlOl3lvpSRtjYxu0kV2htz7361jz+kJ42MtbtzzW08
zLcTIFFBbX26EExbTHeJoQemB2lpx6kOlCv1JB1KTUZz7veNbbsKe9qlNwR0ZP17fd8K9tMZpYmT
PmNH9WgnYEMHyqEtBNH8t6AmtuyDMW06WS1CwtzGo1BlZis8KHMCena5K4GGJREn+k3sH95jLksa
xU4Edzp4PtveRJ0HYbogKfxRuGWq8JrMlS1e7Grj1l0WK5X4xENPGsQ1CBQukl/aGxEw/dN6K6po
iABmZS1lMLLQhKRelwZNG8wi8UrY3xTCqk8ARk1CkLKqWloVSj555B3DuSGjDhvbetmg/m7YXQM6
ni7PTtC8qic6CeG0aky941nr3vibu4fkNQIy723jAgND4qN5boJk+/mOLiN0FV4ckqNLX8ppg18z
5Gy/YgSx8M/CWUOr5a81TbYsO1EWUcFQ9TZogMm0Tkj+iQrrpO/WvILlKfInRvRDbm8NjMfcTmCZ
UKsSrUC7JqDQfD22DOK7UjlHTyt0+T46I0OpvrTokr2WRwN1L8WFRizDxEbW5I0QQ8AKM3Zia1z/
9Ke5I7G5EEtbJyV9W2HTge7biwpYFk0UJlCTHoL8WRayDE02JYo4AY5P11LXzyyknS9UP93pD2th
eCGEM8IZ3fx3KHWqym/oVo3XDweALSc2RdVVraEAyi6hj+DQBrfjFF948lXwyUqqVQL+k2B95BPz
5MkwdbFL5zUdIATdLoLFJbdqoAtIIrpz8KEW3JFfPCoZRi3liba0MKAkD9NsZmNhe9c8RKciETG5
xwlKvRU4WJ0XMCPTxjdKJ4qXPi1ZZhGiAbdMU1U/ezFfRxFI2aRNvP/Zjbh7DW0bCzUc2nj5Zrwd
530FAwSfvKQYnFO2RoX8c/J5qukNDx99xIRe+qTl5ZmiUMpquWzbri0UMJdrazsHrFz7OHWyQgHj
XaVW/HMn/jbEXIDBGvKmgOgTwOF2st5GGLllytDBBtO2YTLMrqNy2tgfkk55aHONVIm5KIdKziBv
s6e2sOJxQVof16Xo78qA2MhwPEEJC/s2q6iq989DNqppKtiYmaCr34HCdtU3uk7QZcoApwadPwpQ
j7bsXmzsRz0R5SWD/6YCmljHKdi5TR+2UNzdk9hXiJb6H/bcmYR/oLxpuaUsE9eJ0IYWvhl/9PRp
qSfs4t/HuTitmUwTmwCLjpc8L+TS3MSgdpdljpwqPCzE0Lgbrh0TAe/wrWt3ugSUqWZMfpfUVaJT
N6ueF9GoRyGw1hXhyTlLFH7u45s7irBAfsh28+SKDNgJjYU7ULZTaa1ra5JWqWLScLJwxsOFBQc7
zalWaoNOh8IxsKtyHb9n/0kVhi856JOdZpPb0EzWiaXbh1+Jzle0gO2eYuItlFPyu5KeRTzVzkZ2
XeDWScwoPRcgHUntbJZzZDSFyshzU6zNJPAiiwfwbM+3EDqaJNEHLwRiG+AvklfIDkwL0s1tQXmn
H63oqsJKwIIO/R/19f9cYRmBHvxd4hHAalzT/0nLZQWqjVITgd8U56BGYZ9eOtQHFPYo1IEKIK5l
5Ns+nOIg8lvaEoFNGbPqOTHVjE7J6gBHDA1axL5MfggtFR2HaGnY00GlkTt54QFj+6/lUL4FOxs5
1audTjVICkjR8hJf8bPJXJkThF8gVFIXjLEksF5/NBO2mwTlSvmvbK8dlojg6E5lZPTIHJRNAODn
S2mMLzceyB3r89H39sXJVWegXt+48Dt4odlVbvQ9eoiGGcx5LRC20pJkFWeqfEvHe/w+JQn2kmqy
ZVeZ1bd+lydY+1iPUNNRfJ5eKeTBgSP9YI7dNw86zlIpktGhn7Yv+p+cSrv1Vtu5AjC8HX6u88br
6eWntZhMEmYX7lksZvEZai9DC6YoNzD8hQsoj7bGX6ERBBhW9KRAmZPl5gqojyah9E7pzlNgoCB2
6afdB8IIxCeK12AfI/tpi6YsiYxnnKjwUcgwoUgBU+bhf5gmW6RRGt6z1Wr/PbFO9V++1XVpKa9w
Q9EGgw0DOQ93JPiAR+BygqLHKYZ0Ah87RxzRXScugdxwo6oX6XAY78kXtPz30ohHE7BmCHze6zHy
sfYdKnHJ79Avk6oYjWuJNh8wI0hZ3WEHaqvz5BewDmyXUt0B3ZCdFWVm/G8awgMdIKqdLEkuvXyI
5KcQcPbeT/iTTXdlmI9okEDsOFM+kSve1HRGK6oF6KnKaBL1zV3CVJ0nylfhEq7JLAd5NqIKFOUM
aJci05My3oUAfnWy5PWgP2wJ3/Vqlvy3jzSWSgnqlQa4X324h8M8PNpFjyVZNLV4noTMpcAxoCQ0
IMKRTkDv167JMa6tR1mWbd2+gNgFJAWeMBNGt4RjgRi65YMURnP2KYh79vmr1P0Zi1sS9BEeMKiI
YSUdFtnrtHJmB6MRmflSwVjISEL5JtGrAOLegvN8zjU+FssrRsglv/UWB9cUMRuTPTD2PDi30MzR
6MWqKYL7OwDIqTkEQkVNl5OSluQ0aPc8p5JGb2CM/I5Iddewn+wB/yRR3C54r8kMVtEbl5dugMrU
2BLUlDzj+aKbL9dwyQ0hZjKNXot+Bm6iAIw47CJpZ5RwdXQmLYeJwldHFHObPgUbhHw7hZYa1VzC
SqWTazNOg4kww+ivaHEloS+byla3sZnxPP5lZSIpdHsamPBL75kQXf4jqugZiejDoh8kcAJi2JRy
LRiTNcdkUq+X9DHklwehPylCPV8GK71HmaWc32K4eF99BynKuHKlGB3hGgA/8CKpHYLC+H77r9oE
UjHknPjM1uxaRgH/XsnMIp0SmBovr7dJ6JZLeqLC8yUGzIvT9C0HVEmrdEpVvE95FJKU1htR7Q9D
GxaWBTceu5t8VHpNngxwtJXlMmNzdS0khEhLFAeHLLBW6AhyIwx4Ya4mr5fARHTBjxVxjToPhgTc
obfVJCmPuctO36sgrxaU0n0KS+jzs8Q9XCPlVgReBMj4yUPNtCvzGzT31ig5bLmrTg8jLcRgiHUd
FCVgyHcZaothLMsZVikNMxFE8Po1qCEepsFzq1kzWr5PRfQADBjN3XaInd0NHMOZ0Ea1fuhmF1TI
DL+y/OH5eHLy9eVOnV18xMqHKighoAzGaHq2Vqr5yoZg1W8ekmZLLsGTaGqLz9kFVIv7H/XmKf/e
BWHe7emESaYui85iH6j3XlkJryaLwJqo7dcN+Qt1lq649cwd95LWJCWHwV3UubHEpSv/u+Ei1Nro
/B+DImOukSe26XxQiWiAxwfR4z+PKdh3sdb3Vhuuh9YcGz1MBvDZk8TID2W6aX0h1P4aRb5OEJsQ
GbRIqB49CGxmhMtF4E3zYyaMi+d8LtEK2pVZxeLwsnMd70sIPB5kRC8WgkWdqZguOEsVyL/JpfKv
vcm1YnNrHGP0sGbpBF5V5kbF6WLlGlaNKl7aCOYkUduaOZIvz3VSqP1Oj951u3QSkB0the/r+VJM
HA8KgrMDdU2p2jCfWqHcIsNQs4GB8pYRnsvBGFfDXiRFETQAQwLHbITf8L+Er4/Eub7ELAfDYDWw
TBsqhDbD+06H8lCcvpIQQHH8FtE3+ZF3CNp0aAoUeIj/2CNQ1BYfTbxhDNqwfyauWyuNL3JLtJMT
ckZsvtQT9pQtInGnS2Bsyalxm7HhwuFA6vfYxh2+CqLlHSQXfz9uGLT0FnBi/1v99EnipPEZM73R
RSqOSb4AVoOmHRfH7daGTyAa5x1Qo5FA1elDfQ1xnffrRqoKBM119eoEoqv1wEfuBO8IFwBRKMyl
s/92SjF6mytfkKtM0iRNxtj3bXs/szHuiK8HZhvNBucQxjPyralsDuZuveMkPRx8qlZIK5qpk31u
jY64XWfeDXP71l1RRG5xj6TzSpvDNH3/tbTCL9tVCIidhC8SwHpgg65ZN5T6z6Tlli6qFDgLopwY
gMjUSK2aGiT3/B4e51pBerIbmcl4JD9U8n499ORASfD+xR9Aku2LU3DWW3pZxdWdXClDNHA+m31z
KSSWb+aMXvEdCUlKhq1JBVhHaN8dDToKBtKvkqt72IKBZ2h3LEHcJxwkcupDf8T20cTxw0EzO7oo
vs2nnT/OI0j5eqFOfid6Qqblceobtr5t/Lgd5U7OVMYNyfmpIN4HDeXtx/SuSk65IJXJiKjFMlMf
QUEpuGYj7roaVlN3St4ZU8Yt62q1Qbt+TJEtTO6TQqJ9xgMOmSPvOGH/u9HsyMHZ3kwJ4MPGp70f
xxf7bB0gOvTee4GuP1tCZ/b26hx4lYkLVonq7h+YuV4EPDMCzq6+5616WMzGBUgjt9cexGds2zD8
uQw24NVC68Jt+dHG+hCN9fbp0ZiSYP9xsZpIiqT5j1I92aIdEEBcRFeprwfaFVk2b4Aeauob4aZ+
x+Z6FGaNl/vadzQJxAXvAjWCXX87J5ELDMPuAxpkR0HnqNQpbqv3VHi7spN05yKfZoKYB13jZCjM
TZPMAPkLWA16W4qtxKaHVK09uo92heqx5EUlvNnYmL3H7NGO0uH9AY2mxvyyueoYN9FE9u4uIipa
PWxbBfPQwD5UC8wUuBZj977rWKtbfPIDE+RC9jdrqNrkhtJFiJ3YQiCN0BQ3ZK7720P2Efan3x4z
9bsKArvHFXg2eMSgHhJ19Ax01lDqrEFR5c4vZGp+ZPsuASP/G4JsxBlMIoTLLZ4MBQLfiJd8Iq+C
SMsti3cIWSQvisPsfE+ErG8HcwJYm/hanbQA69tZBqXHpeue1z+d6OgQcQBYQt0O7ScX8LgVM/pA
MNhKTxf8B1cB34fSymhGwZ6qNx7FXYbTG9pW2HwXdFP8x3xCMaH1B0DvNznbBIiIsIrxxAVGIthJ
tosFf3VrBk7LfVt+TmVbi9yBhl66BEk1AWjsFB8I72M3by1CvIMa8iOK6Zc98UdnID3FKGD+v5go
SUzdZJ/dt+4QVVaEl55+mspKjemSTcAMGloOCD9xHZjNjnfHRmGsgemq8dkk0FrrI6tubM0f+ZTO
iGclKYp/gyP+PojQstIfOrrY8bNJjYTAS5VcClxo5iqUsBAYXZ/DzEfqePyHkQ7WZmY3nKyIK1hy
Ljw5OF1umAt8ZrcKy6PwbKjc4A+oYGYxCuAKKlcdw/D5jOJTbtxzpPAYskj++m/Axs+LPcufUR7U
0eA9xW8Ey75hamZnQoTYkImfVPj4aZ+p/v68kFs/zysK9EKHTvMtNJ0uvY7Wt3tCRR2RM4QbHXNa
6Q7o6Qivb20jwCb5co8d7SdkwzRXDGjR98TzIZK85kLW1DiiVYzGScqAfoHyzWHhy9F45Wuw4v7t
U/snw5/NuZ/dnXjkGeFk+IPHYYHRmxQhvxUtVApyienjwLmsZ9qN7n4bD4O7Y8RSFzsmv1HSf8rV
Ep1e1hiUUajut2h3RcUPQwC71j2s6D8mFcW7m96hK1RmkMH92Z/dcoiu+gGHcJ5mW+Et2LBV3tjz
C7iI9j4QyUfYhdNgjsJ2gBFq2rRBM9nOzLKWdsn2Qu1PZ4vpojfrqOIooVAYT+G42EDxXyPwjxXP
ogenFqXp6DhGXDh+Oj574UVUsPL6mo+UrWDlElauMELzJcWw2VLsl6BQeQzVCZu16m9fqATNTR33
j+zP8r61cQwYrQ4V+gAOYE58FUZzQV752PcyUqmatgAzSOE7QFJTv1A0VZD2k1arpBW199GoxsyQ
oXJFmYvkEV/GVI5HMQDytLyCpV3vtCQLHaY91jmwIlMa6r7fj/ofdrpBZpt3gqFpdGW2bSJ76LCl
5nqu6ZzjiGAaDalnYMnF63Eq8/DZr4+YqPckVkesV4MfJiMxb+pySDIkgbEU6qoRzBctQ5CBraR1
BoVJe59RblWoGTc36GzqJOWW24PtilDCQzUoPIhwTIw5Du0V1LFO4fqYRKHRwEKz6pXNKB2Qqszn
JDu7FTXJMz9curhDr0RS/oVzks5cSXs/XyhZpsF4tOocFPvm6kOgK701Ju7GfmbfSuLSetPgZwFf
gXSAfMLWzs6VWeK52jhFMef3s+iymQRw0RGgGmwDzI0z5xFXaaaaaK/tHMYxJC77gdCy7X6eojKv
WchyC6hviqqRCzdEeZdx+/XSEBC102c2z6JEj2yP6uYEW07Ex1/Wf7zGx3GYKure6TrcMN7b2Px3
6DDlq2YtoeVYEgdRoS+yS7+Pp2G0AicGZzdlUlowU6dM8n1WtGi5cOxbw50lFfxBKacH5zYqHkzc
Ix+9aKPdojZi1OQxU5cFZ1A/nVe6O1bWgX0fjQbeJN9+su8wG1Y3r601/9adh9yu829Hm8SSWOB9
QUQpzmqIwGDSWok0bQYOaIf6HkYLxATseHJXc08uFfL0ixsfvV8Tv4ebl9dAmNcT41Ox02gYZe05
Mi5wBOowDW1xAvBFJkVPp6KeHuMAYX1Po0DKbim3fkJoGTaaV767q5SZMAoQvGA2l8oItYeL8U/w
xvM+V/uuOztSE6QzwwER701yGKWXRn8xhJLauv37YqDjxrzvlvXuuYYa+FVMM52nSzG7b+5KaNQt
/YHJ6RgsOcXpy9SkvZp3jE+VdEZURWE6LxKQPXvookNNpNzdL0TAHkVuyhO0cx0pxiyDd/ZFIqL9
8rg7MjWdWV1WrImW7FbxVZSdVg0q++yKxswHTRDCHmfg7PmyWEZ1C4CKsSZo5V33zFt8NjmM1ACy
oISk8McJmCjtl6vc0c5o8glr+QbHyom5cYsLrxX4Mv+9sIJSLNNbOt2CkyK2ejshhC5b3Zo87rxY
QBtJprqiTn29pJfxnVbw6lt6wBoACVOcGrRBB1vA9M5pqp1oW3xfws5FZv9WN41F34h/AcO4Q5nX
XreV/Jd8sO0OxLjSc0WAzZxIqRk1wRd5a0YaaHaCl8CFeFvwy14mpaGGps78vdUVp6nhUR9+ZpN1
XwVIf3utVWhgv0vBPgkoYP+Xu1WZ4deOnfjMgE6anQg9HCJIAz737H7BtbAhyFB2DUYPkV+efuGl
pDkBeIlMFb0N3csQvFxeDcJvAh0CUBWm/8r/4SUU40Mc0KnXPEYW4DSYf3Kcm+9xNgAUo2l8aihw
tM6f7lh7vF08vkKcNegXZOkQezl5ODb7huPNY9EQ5GohV9Y1nT80GGptR77wQu48ogHm1EuI/yOW
kEyUZGSwxfy5dhNMrI6xKFO8G754Jc4x9V9vwG37OkuiXyo2TWwqzrh1aYwaxgkyzhM9hWGTnkbp
FmHPlx3Zl9gBo91/C/Ep4WergV88g96wykAqybl69OZNyAjI0pomk5Vz8CpQWcqXQdIMS6yK6tra
Tdu+yS8myJoX56gdaSN2Yt/RZ+ppu0gJqwa+PZ7ZeNoUAPwCUhJoQ2h3XEfL8Yl9G3EoUgov1Wga
6IBEeyBK8DuWEDZNEiF4TO8GYhEyxfD4avY4zpUyXH7cERRyOEaRuW+Tnoi8rKJ1p4KXbzgSzKy5
beHvZZxo5DLBFqKG8y6/8p49cxp1g/5f/7QcGavHQYrVyL4AGhOvbXp/q8LM9Nbj3PaDEwvuQlbS
3I1rY8GKlJuSYLsY2K/NS4qC9c+z8Il7BWk/CPS2NMt8u21JfbK0Yf+D8Va1kdfkoOyvjiSXpkJM
5VKceRN+LiMGCk72BtsrWFA7iiNTuBqq7vsvTP0NKfuSky2wOYFEzQv/MpbJX4YrgQrWT6oa37sP
efOAzm25UgJ6EBiWXlCqDjjEg5Hshearx9vhEZl5/DXUsYvKSdL3hRuVMDKq2gQAyttQB+yFzHR2
OV3Zqcgyl9umMatAR0rLPMNiSoF/tXHcAqT0dUlz299B5EE0ijnK060zDa8nC4IpsgAnM7x9PwwR
szjXfu/FZq3LrVUoCMhVKEoSSWPE0L6a3AHBfwTUTLJBuJIaBVpuyovA3qizGU4MZMqfUSoYax1o
z90f7bxPj3epwpbBO1OYIRSG/wWYz8ZXuRsjtVip+5PPCmyEAg91uyCLZC/FRqJ2BVc1st3z1QAH
/l7MNdvTFok/G85N0XtuLMX062B2nD4UZ74pjACjQld2HoL76YYdGV8hOC43MSj2E9a8Gp90tBPl
+De17nIawUF2osxtpnn7X4nnVPyz1VNXLNDnMckbuSuv+6wibTTB+FA5c/c7RBq8GNEV7Km28L+Y
Q1j85yeVCsL9jfkZy7ty+5TMu+cUbr1iRV1ApzFCN/fjHi7mPJKf9ddEz9kdV94iqb6YReeBw077
tRPFgU304Sh+JdAxf89g2+HtxuR+lqnZkuOez1sQcgYoDkA9qp0tbsNWl2I2HvlHxc8SHMgzrdrY
3ecNpddNIiRHp+yVRs2ZJA+iFjRF16lg9KGkq+TkBUdna1/QVjie1ycisHhMnqt0ud9A4YEOrIYG
K2GtuLgRM2ZmnHVTYbnMZr6icRnVgklbRu/+r4dlMGs02zNXYxEobExKjqLOkC9YcuwvrPaUvR6c
02jnbT1vM9iCqFBkHV+m8Bn57KMwEsqjQ3v2IRf/JemoMkmVuHKrZng6Xqa+lf425mWtONeAtzPt
ny2zuOqev2KWo/B9keFqz9Wpzw1k9FffnDuE+jfDkLZ2q42otW4mxQ8zWJ5WqSYXPETfagvJ17I5
qbcR8pcb0Vp0rfuv+nWqIdCMU0lWzMESU8EvMS+mhnR+6kheabOEfjXH9Wljt8KRJ0d1u0k/wJiq
4IjEIYgEAGv0V+3i2dCbVhLsOqatmiWPKtyRtVAPT/davLSfIOmVGOjn5nO1VzpFaVO/Rk16L79Y
bRewBqhOQQV6DJcFKEtQvBBpr+TT3T+TaYxij5+WfWlc2exZRUrD838LherAX9NWG6bGOAUOsEiq
ghWCQ/HHHK+R4Jj0zt/wdngi7+9XIPEyaVFEnqjx2XNf6dh6AgZa176tIrjtl5ou21+rzplHvNfY
6gnpofnxIWTRa8C4S2ROFsN9jtPvTQBdYujkED/Z+CoxYZoKEZK0iZbrZOGLS0mJdyYogFd9DqSC
AQJXhFmxUFq3Xnlc3UVTYv183wTWQkZAtprhrt8yYzFhrmDsgsmLXIDp/1UY7A95zjHiKTH/0kjh
K3BZd7hYhEFyYXtpWURoI1kE49LCoNA69BqurN9ZdVGkoDg0X14TQch2Ry2hj17EgOXaRx422FPT
YBBDn2NX+0Txf2BnhTF5qCvZVPO0znAzGRAGRcPeG5Sj8O9I38v/cfoL3cNHLApl5ZSml24RikCw
yD/8zKouhIdK/7VDjmpyAI+yfI82wTS0vfeLAjT1jxgCWpWHSlguy1xcD7UyxnpFrk8YZtPItJ6T
IsxPIKEzfMC1R85s/Y7LczsyL5M9QeJF154JkaHegx+NhPrai127VBhKt4YaYVuIfNkc+AWBUbn5
5bjxzsUSDUVA+0jm5t87pcFwdyYRrD5u/2xT2GN7qxEJyMEO7nHdO+3wKFdF+I663qIvm4mtnYpw
LsWJYIwgVseS0cW3yIZQAcEwSWUbiEp2zUFobMSywWmPe2EqB74ssk3/Pxf3Wvkq84KUK8UIOVnD
LSBt7hMwppV86tBHNwH0HU0I2cxyTzwZ/Kx3d+HN5EhdAPtfi93p1otUivsxAMWxqhv/rVvA1N0/
H9c/eWMRUQLb4hxDoGE/tN5ZEen5HIIUEmRNxxK+4iBEp/SuUB4fofuS+4n84+4kADyGUWYSla2C
tnKVb6H1bcgAl/qbzuve+NFLPipAYE+qloH4KHOMtkBNv6I+/Z9tx93dAYtfRK7XjLe2ImFF3fVs
/ZPj548KB1HksWSh4Z/KHJ1g7E6aZkjtkJA4UV39Y6sQZ4jzY/8+57UxKtQwu2nTL90gS6YnalnW
EXp9hlR689LpZb/wcA3qcQqVgKIAMJFmC1D4AHP8EeF3RTelYSFi9ghWS1yiw96EPEn/SwwtPs7N
02c1ortqB5t/n4cLRq5ZroemUGrDFTvby1gDo5IriPnoIh8AzUzngCP5w7vU6xDQcvvnV+8fVSwW
xfc6x2Ub6re0O0racyqiO7XMLwjgoLu1cIgzA+f4a7RFobgfSj6OuNx6ygcR4e/CvNrwVfl1UmTc
4f5Eob6+hokpYqnqLW8LUSXYp/zQpa+d3d5ip7OY0+dPw8BmNqFBzJRpuKEneHjNUQJxirUY8zFq
rvsl6rvdmwj3ylBPhEDqFeq7Cl5pCpVfN2CkFHeeMi+Ok+S52naWnzghfwhFnfHR4Umc8qe7zwQf
JT2t+cMTWHCBmpMhWbfqULCrNIWS+0SCpI/+YONHW+DB4eqSw3hh0E2QoN8DvZw8SSB5UbeC/N4l
05VI1AYZmifpKk9eai2eYWhDqbmfmj8SH8PACb5yWEAAsWIwcEWs0D0qQcKz4QfxDD9qby+RiTmB
odhIwYUY9PRJLTSRlzU8zGpGpuhPnGWCTo+cZfLZV7TgxtGGSScP1i1ORr2B9ph6QKgSgPmA3uqQ
aqEbVKAexSYp82YGNTHajRyi/dz8nvdD9Fv9f1NQ/1+OutApzy7CKbSxtn5MQ6iYkW8IjivBLaDq
CxstKcN1U9uqGbIFKeHy9zjiDUUQFWCktgg2jV2rHHtATWayZ8+hwMqJArpe3eKAfSLCUMgPSeBJ
jxwtL+2hxkmgMe8kl4xhRYAb5s35OGDRELLDvC/espRKKR4Gha+jLxexzLG/L+wZjMETAGU7I8SH
RvkjW+cMYltXvRebRJq/loJzghHmo8tUbLUdcdFT4+2EcJ4DIdTAfx+EeFYi0xfpODign5pIYvmo
ZLDy1jQPU50DTwj8X2o+LPbcw8XFJdrAuXRsr5H4v1dJVG1AzG5Fw6nH7kr5yEUIIVH6X+1rjr4N
0I9VRyCnKYvZQyf5dOIyX8djbIGdROMAShBg5MNCISgEWyhRGgb8/admXcAaQphWAQiijwDxyThw
eXTn5Zk3PtFxnL8kBFl6g4rfx6yTl7HBlkz/11CysmPhWwfQqIg8zT4K1NKWIZrs1k+MkTdHl3hi
k8eS5MlZpYkeWgfNNc5lcDJ6vMzSKT5G/yXGRJhIJT24G+Q67vXtcvSMN30RI0/WD4jh9oToJ29m
fbcogNOUAY7daF6Ywbrhe84deTGDNJEFcCalD9AGeQ5hhb73XzWYS2fEYfrGmK2GKF/eY51OzLTy
S100WUxjlW7TsZy4WwLpJB72Wgh+3XKkBDxDpMMXF9hmvnppOD18yI5BwhZBUW8qMEbAivN5c8fT
qg0Dww==
`protect end_protected

