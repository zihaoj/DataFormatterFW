

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GW7UNomknr5Dw6Tz3R5svbJyGexHUbbDbEMITb5vMnh20lFU2WL990S/aYPAkkqJUjJPpL8S/093
yhlfAz2oXA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VPJm0bZrrF2NVzuq7ao8MAK7FE4zNvrufu4waB+nXHPnU/t9wPsgu2I3ct/Bnh28+FN0cZR8TcWt
v4yqKihHeubq51JvQnSQBnzZnY/j4llNeta6yt/tyW8P1UQHd14W5LYJ3uilMxX+2FO+TBWdKAi4
WI9G7LbpVaiaSKjRrUQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QNxRzsRZZgR1gVuYo8+jKDYfKZfPisAg2DlTO+UtWSAU6Gzbvs6mMigOMdL9ZZV4UfsUw/2OJ5u+
S6Lfun4dcwsruwbxOy8picXmvBLUdLYm7bTLF0yS+A35sQViez7eTBeV/chDoMNsz5/KAmkP4uqa
UAwzHT/cuZCBNeVbv1n2bDA+5kMv5nCwcNJSACh254NPEvFdKf09AAIVWgsdVg33SRRzbYw85Zro
NUT2D1AiQIWC+D3eAIAGqV7MziU0hGf8yxoqZj28QBwS+/TDOZ5a96Uztx5lJuLm18w0vX0/3kFG
Ghl2uPWKnbELkf1REm3OzaVlFBuQaXkp4PEe+w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
j2GHCjMR7MSOEtk5/r/rouI+9tnO8tdJq5hVs55zjHiR2VpvNE4+EjcJr2mtVGWSh6GfYvEZ+lZ3
vnBz9lyo7eZUusIT6lSmCUVtb0bFg7Bu11ryq3Tr3LmAtKneid3NWKmkMaz1DXj3bq6CXcFApWmw
KzjnrK1p9eZ2B3zHumg=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kZyUDnN0bfuuqPptXshBDr81sWyb5cUW5RO54b8h2tJ586CW5VQQuS5U7tJxrVQsvTcWZuK3Ya+0
QfNJ+DcLZh4XQ5+Wjf+Q2uN+BwNpFDeojZKk0scqeFl5VTi93s4R6PDOeqscbqcxc/bHv28DahuH
F8iiTjmdq9hMc9MfxKVqzkyq5oYrXP5lx45V9Lh26i5lGS2NNXQMEcUEK2ioY6FbrOmg9jQHo3hr
aYsaMjn1BLy+9BIi5FRRfius91lUpBj93hqbxyHinQVQ0JRsXS3YiYqJWCyYWIko1b9NdOOBejVk
YlVQ2U+XhedNe/rfBgIVU9bOajnmSiSa7KbYrw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3664)
`protect data_block
UEdY07DzHl7GGwxljHZajresxHvgPg3IvugN2Vb1QufR0UBhXZ3iBtwbZhQXFQ0eexpVdq4IYVrD
J18VrjWIeKIkFB5HfJXxh1hshso1YubifIkVYrGzfgp0KMeNVx4kzpyS9WnmiEHRskGEm68w/xPc
6PGPfjnAFyiQjm32JPYXWxQhX/FBEh9Z6sGpEHgMiUEoQvc+YfS0IBNC9PWbQ9SC/tH6C+cUZAzz
TOGgep4Wnbt80x5sXvgTGQdV2SZBMgb7xXXyI2bdbEbGOLCXD1f5Bnng7gqGHSIMgV1TnVRMeuRM
3QhRARE+MalDf2SQ5ki+VyXLQ7g0va8V3bv9aPFOJDeUX12npOaZSKd2rQuMXobnqPkx1G7pxs2m
1TRW8x3KarMbTEbXhq3qEuAT47mcIX7xEnf4gTuZPXhXxNJwPILm1yoZpTuijmh1AvBJXxwC4PHb
jPNLQX9tSz3oVY0KuLP7cTDh+MGmROPcn9ZTVlPoEN57ut4m5lurrID0Ra5gIGKo/fr79u5EbbqF
QdBonHbkw7eHWqFhEc8WrsWd5gLSPDa5nYyyChhU1cKZLC/SY+crjpY/DcJPGSwidWH6EVpoDWPV
8OoJeLMUsTY8GRxxu1aATIXWlFuu4UQrOagT/0hoCtnrzdgZI5aDWLNE1Xa+k8M1mDLfnzoBbAJQ
AT7hCgP4awJ8M9mVCAMU4HlrAzgdhCxTS1v2RHr+nXhCjFixXcYnYa/123bd3ab5/X5RrwoixLug
2H0B7uZBi+RWAig0rNDMWddZdHJ4pJ2f/rgbrEJ2YoXYxWFa1QA2Pu8Aubz+Vf342VN9g5AXoTZz
Vciu7jVnmzcqac7HHLbNx6pkjYaYTiXVtdKvKN1RrLaTGdHgOjFRfwY0rJ5DqeGzY1BiX+/P2nvF
lW6wJ8pRlmShpt1BAbKjs0yHxwRS66KiKyuptG+As29iR/mBxTQqVvuL2wZWqMWkd3HR6ydFI8yX
NUkIoPYQ73/pNQSUSJWtd9mk98+vDBbuNhHgPInOD+5nNH723s46xu6wZZkRGUi52IsZcf5WWlYS
WmAz68MTalX1TlM0i4rhcBLH82L7poRoh5ddkmKF9SIMJnA6/qea/UUh7iN6woVObtNwqJQovrnV
HWOeGCqlPmIj3qgLgHMwn7c2hf0OjBx1B61Q/iEk3Bhyu9h3A8Ih6UeUtZHnp4zMyDd0/K/plbu6
8H+0nIN86d8nijZYBk7Td390qwcyRj+uWj83KAk5AwQdGlud9cWGSj9fIu5Ug78zJddsTJtaN+2e
J754ZzOBrnWqAtpbJMZqRbc22VIBb2v6+R4VFh9W9RxeTw4/Hc7DN7euCVmDPZMPnPIz3q3YyOYb
tDT6+aK1cq+iAfgtxoi533awcN5vD1PZBlzgX22mgI5Uzbn84Kq2ewKVMER4cW8bjuvhUTVvCkKc
aGsA7geBBS0yKC5+UJiriqEqP9eMAo2ASLhgID624U3ymBgiubzilx6IEvWDJnrDtEIf3OuUVOgl
sR4GsIpAsEKD25B4p/mCyuwMy9xBqAbuW7fXcodiuUVV0vqRglsRq5uKfOjoCDfHgzukqFFa1CXw
BSPRi+UTUxDjj4jSCAVB01VsUkRZls0fMYIEejomHQ6Y98D0tSbNh8DTsBwdKjVMNBviq1pPVEjq
eqTW3tYa/aKPwMnxH4U+FfYR3EuGSFY1N2bel7KjWREvrNOGv1rTA6mURP6cNC0cArII/ISdZLzu
fjtd0HTf3tp+T2tMOtreuag8is79BetZ9WzWOazoUg41l1E+vay1iT4Ht41OOk9b0WAnw720H4sX
uk10q+vSaDq1xj6Nnn6kl/t5wEdr089j0SEz48Z/J4pUFVnDR1mhkAvuONrNLGp8XVePF51MFbBx
iZGJtvUPFkx/02SPbSZ6JKh+73Cd+UomVT0EswGGm+1wAFLXSyO+qI/mmJ0FGerjla5+yRCkJ7xu
myvH5epkRcRq6bQdDrgMSQbjsUl8zO9yJEmBncIiLPVVVi9hQUJ0QCXNBwIc2AoH1g3F0KJtNgs7
ULAXPdJyIj+5J58F+fv0uwOH5hglXQwPafAzt4U9ODb2qzZV+E/EetuJweHG78U9G16AFGFeKiX3
fnJe2SvqU5ftS+eSBSQL54HHBSTjT6GJCFZ3r3aM4GE/xX+PgwqTpp2OEgwPSOs8SeMkkq81bCDD
bnAQD+d5gySInSOfqjfC3xpzsfwxBsZvLR4b+5DXKBgXuH3XuCtTWBdx3Ob06oZfbwU97BoVu7I+
wySYL1m91VwLvxd/cdFt0qTgwtlBdVTuFPaX5yfAlD9JFYY/sARQPkN9C1HzbwFxrfA6wrF91hFS
IZzHm4tAzSsUrcv6UuaalCADD8xLnBRnrNUTYTfLIDJGSDXpZ+bqxWkr6/USyV46MMmuQybhDpKd
JpNy3gqY5LjmTEtoy8SU/st4y4UlV/gBZLS1ieRLJCWwRYqYZCbr4mrZm9z1yjxilwceY0k49yu6
PVcKd637Oh2RklElk9nsxotWceicBzEde6pBQP4Gl4dJ6cjyH7Tz47dUgsA6rxPU5D2I8BfkFq6p
/i7OpDtgX9JPNoG9fcq88gUrrjavm+jdr6IY9J0EnCNf4xB9kE0LZ7K1LIMtIIrQpQyCwZrAuzul
9jHHbgrC3EupNreUnLRh+srj+gzcsUqsv7lNLteUZ/F+NeLdrCC5PPGgCJLjf6ACuNapjh4qDSkI
5ozzvkxSM8vfPE8Q1OxRKc6Bw1rtq22Cms/nZuvtOpMuGiNNkRg2/3pDlsx4My+WWf+wGhu/BUVb
ksrgRO+9jZgavJSRdMgthPDR47iFe8DmQ7G9BHk1D6CSW/3dKqajwfDWEdtLKKUdc+Ugh3MLqU3J
66vUrEZcGd4cxMIPCMCqLS++yFiLfL/MhKfxvk3KI7ZLm6EoX5XNftyjZiBKbKRwZJSmEQQPcUnZ
ePvLLcgv+XvCPWKEE2nOMeA9RjfUVgU7sNtt4+tdkRZ9bINjlo5bfOoOH41XBAZ0Xp3Aj5IIwYPd
0GodsE+bku9TCGq8vRlrPNnV2pf4xUNYO+BaxuY2E1+CameLtFB/2rf+ltbCgWQzr2BbSO4El23D
p0XNLf8uwVepHSH92VCVYVs37qzrheExJ+D7GRqHFfYzdkEFK17kEJaJ4mL4XwDSJ2uDsCVoJ0Ok
eAHVJi9pkDyYdMRTAD9NMqZXJDRGM+mz+7q6iWLcTYhNxang0eyp86iFq52ttQPMIIAbqXqAeWxH
udbS9DRmeLWvXFA9XAawSxJlsUSd/L50xZOI+a/QRGtmyAOQzYoTXiXq7lbQLa0iaAsTBLtBAqq5
Lfb35nCYvXEX+vc6+NSDq/ksy1cOKx4c9P6zvkTLDcP4QsmoWlQDsJg9HDdbC8T8q4MOP2tDDZ10
KWzxARe+aKCwyOyei6SaaDQHvcbIIuBKih7bn13VwliP50YWCjP57cR1hZ8v2inMxhVytJCzrfyy
ufZYwSB1yDzWAAC+zKeI//Uo9UnoJqpcLVue8mcZ5RYY/AaKa7SfIP9RBdJ0frvHHHxffHzPuKuy
W/qqee9NNk7Jt2x+IMjHUJr3vhzlwKApudJ89G7cqOKdEZ8sRBURDT0W+pUfscX+6OJQ2vt5aVzW
C2hLFkInImRCtCD3fBRWPguw+MWZy3Jy6WEf/pibVdeEeBa9qcQS2tpEsatuCuCqe/Gdk6Oiz3UU
Uk589YSqCKExa2BprGQK3bKNkaLO9NkcQoNuaQm2pPc5usRqEBQgcyC5ysJGm42NTMoKd+IhppVg
4AuaJFdONfG3bHys6Vt/iGk2Xy8hgtFNWHGfdcuZNGVNKhqGqnFTd1PFIXzHW4TUmkTLPJSoBdSG
X8i9b7oqeU3Xh+iBbq1Dn7u7rWug2BRMM8ZRUqOJZUGVPV645mWjSVrX3x8x48dBH83OHaCYztxk
DjkuooNW3rgH0ykaagjD+aTc8vGiT7rXTd+Ws57noy76xdH9Db+rQaU+tJ90I6yhtERD2BH0Iuuh
f3t5Qg9mNC3DH9JWXiHyZIBa0hqKTOXF1YUdC+zkN+l+INkfzfv/5w9zNxolIoiHwRTJFFHuVMux
41CyKcMVbKtUkzetLym0j1w0eYlLEf/NTZxqAFArHrgfFo26gemx0UqIzt6MtA2cj0HP1VmbUQWb
8wSibIgihSqRUOKEs9GpMm7HjDbXn/KPAVlG7xrO6wXfS1lSFYc81YpCKzLnngJaSgswG1Ovuqae
Xcu0EpioPArarKSANmw2Re9OP6bPNzTEz258NrLFo7cugXNTqYhnNnI/0ILH/iDdLYXXTuh2Yjvb
t/HPR45ypWxXdaVwVXw5yX8BuNBjwAB7yLvw0PCCNa/SodII5nO+BJ1FmKAlibvdwh/BDed2vJZI
E4wZJ6hIKwJCVBF6Nno2fiBYVYc9u2aLmShW/LTbozRCnef6v5AwOQK3SUQ6GypDUzlMBMvA8pxs
vcCfwAgrjSpSDTufNtIpgiIXoXiSkdQdYcjAPi9Lut/8dxbPMX5AdRToi8P64K0r9N+9GaVjUvyl
YNXkblVCgu8u2jhvPpqCslxyPJNNSy6NANYSqYS+rYDVe8nZsr4Pt38ElA6M2xt5ZUU7TXEG4E2u
+uf9D1eVM13J5Wg7XCKxUJfSKRPagGqQLDyF7EfjHngGHSBadYp9U93/EQatkbll8SB65+kF6aw6
1k9rsf/LCrjBRr/6hKxDEK2Rero9iRf4N09us0oBGERlf7oBGvKlfNiSeNh5EopPgFmD3Qqj3GX0
fepRydithbEeMi0XV5ELGXApts7f6WQWmTUiFR9bzzvkxGyDZJ99gmLD156AsL8gC+0WfBHnncl2
q1ekPFIH5xCQjY5yoUolpg==
`protect end_protected

