

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UG3jcx/PuaQu13KCRTkQ+xPvYDp3rT1vW297NGdT9K/urk3UFCpDApQ5LvNuVtk5A5kvEo5KkwDj
MOxFTebTqQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ps3S5pPkqVtode2oMxRgCxvnQZjEhHn6NFyuCKyy8TlWzlVhMiFYaxk034aYwfAZglveNAFp8rES
o5uVicjMbfBKNdz/kz5Gz/sJGj8dVtdAg/2pPaX+f7J7h/laI03wwpR2b2dDmAE40eRp7ULeEX/i
wjg5pV3NAMcC+mH8s5E=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VtWNnrUKkU/06DY2HIDBNX3jYmptyB2QYwRWn7WjCK0szHZbBQwhRd76u6uOnSdCzOZNosVH3d5+
gIJpuepx5Zit17hoCHQgCwCrP7Z9eDIqn5vONswMT630wEZSXifPherkwtr5CCKoG2Fy0QD+HfXh
WPzQZhm73YxcYEqudSMwm39kVlGe3Qw+5Sbt6R+0zQDQ9t1OPCrU58h1mjx8G20tUtCWv9x0owSF
g9A2Qnj7sGSqoL+JgtdCCZwKy/RDxcAk50c7xbgdlkLJkVDwGfD8y/kU/sjlRwsW1TeLa0qoqrw7
vMmVrFEEliPiIS+9n9a+qY94B/1lsCZ/l/UclQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BDAAmOSYJ09o6amcdQ7JQ+7VeJWei+GHMSXyjkrrEnbfYxY5NZ8VgXFeRGqiynyTEDr9VMF98Asu
JYDN95VwMAO6X6ID775tX/tdt6ol6sKDT8C2YXcC2vlr95iyQheD6bGpgcZ9qI6rDr79UhyM3QzF
iOZBuYSiLlP9RPMbaX8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aVgxDTLn0rR52Th3vaMDtAgpbIwpXBjHzKELwGi1V/6MYtCNDRFtQW0itNrr1RzTwY7E6HB5PMzu
UgWs7PhgAF6y4enQ6pHaP9bZWIpnLIU6MPazBrYn0LAmJrGKFCOQ+063nyrWXJE20wj1Ntp6LVhb
Qs3/C65i537WsJiIkjrfVqFD3zf6f0mHC3QC61+wSpmBNH8R1rsDrFFx9Alf3TuknSvWhYCq7gPb
d/Yxht4yTaKxMWXfSzE34zg1ZCTJAoqWVSdsulDZeBKLVCi29ZxR3yrliMDBPbRed2KwkVF8Ayx2
oSo2UCHd4ymI95ZXf6n5SdqWaYNZH9D0EBivRw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7456)
`protect data_block
Qk8yBj9CXiXmzg2ysfzCVc69Ea1EzELI+HSKLobZBdqqCFgA3xZbG5uyyhqy8eNXmEhKdDt1cOk2
3W9McewrCPcv2AyuLqw1N8xjUB2Gl1E+6zEHGEPIuoUbhzbUr7NDlXjEy3ZEWQBMrW1JzG9eydHW
l7I9r6RcuHfUxmIx6jlmaHOowUbBnJZDGaxzLAgyT7+dE/r0iQhPLWtkU+t7QvQOlkA73E8VxZAm
qoHnT25dSKJY4HDpt5q9RFiRbzkufPuQYJUBX/wEU/sxcXkpuFM1lqQ5dr1pfBWCJuWAVnw/FT4k
R8lv9heT65F/fojaepSfNgOuLJDuIGXFE+/b0Ddn254ssOHdKBOpWFr8/FWU/nQWSiH+QXb7ZRtL
1UZsFebfwlRE2cHnS66G7D4JzjQn9T7kH/BmuLYORqdfVLjHrAoKw6C2odMY/CZ5r6uX72cdboAT
l5veMIIdjF8oRusVvvyMGS9AugdNAnon9N9p9ArWqcVJtS3k7rJYenl0rmM1cfNDwfxpdwzc/Qx9
p5WFZ0nwEniMXogAGyDF8AexxsshaXx+7Il7ur4P/+m2FpgFDO+yCVyPTs8b06WZPDWZSuKm6Ha0
FKl1W0+daOFFHBmsBPiXhR3PdAri1YSaP4p7IoH57Atn5EoZijxQbTlcHxiyFYzNbEU8uTFjmyUb
y8NmqT0eZzziGiQoDG7nXsNWrE1xp+YGZioMOCKY5711SJOyvBTKLz588ohTv/tZ/ZrA/WoWL//k
RmNvc9MtdBqxzc4iEKiI0hDesSkLbdRVQyG5zG6c/kjNCAmcmnoqnq7EfrsPAjJeL0s774ZnMWrH
IxFv5bo9URAvSk9gVNjC3aTMQPS1oGEbjMQZ1gEbKrbQ80V29ZzY0FDsRYZ87tFisV2/HeZ2CxLK
FqS88ILgFGUPZ6Vq+l/MOx1jO+KbuAI9rXFwTvk4CAglrIh1tZ7n9jb1WwnTko3GysOMYv4N8dEO
jWMORv92ZgArtsA8pPL60fUWAcDWYP/GpFXEJBxQtawp0icgfXS5ixrlARQEaQJVI+4xJ8k0/J2S
++b4Kk8NxKTmZOOXjnVteTPcBCKXoZsjSpIQKCmEvImOFoox5tpyjNALNJtd0Tb4qvxcjNX0HES+
phgTOeEXgPXeOVAehy/uTdKzoADtF8/759qdtj8U2+B0s7B58ySSKQmOTO8EdlKKurniSW59+/eM
TH5mtS1Rxx35/tGzLyDwBUlpUNI8hD99EcVjpwsmD/Gh3xm68+kqUXuLSg4q8VTSvf9tvnA/bsum
H5gDbBCERQomyNtXnkOUZlJEls5brLXlfl/5pUOOjJ/D23lIuPrvpYK+quvaARBpg4y/NDzDdwYf
M1Lz9XfX0T9vj7b7Z8varrHY6uC3zKkD9a3W2Gf3MnasjJa45mwcpSncvJ0vsfQeEWQards2C9Tv
h1AHCakzI4iDnuWvrbhZjLrqJ3rIreFqE/kJ94q2fmrCOGpPJbw61+0sY2fx1E2Z18jsbT3jYs0z
ORnXO0yN3D3Qg6qKx8FN2IdRcPdzQPIwDxAya3HRkfbTxizEBVMKAPXJoAQGVC7hpjHIBwoYWvJA
JMvZuu72+HfmXYF9JSTJTsn08nHxMvgLctQqiLQrxMxu2WCyA84XvM1Rln3qMiabPWst3TocGecs
XmbHVJ+/OvBeRz2kzSUgMloITD+lmdIrroAlyAf/wiJKw73sqc5xHjuVuwa4IKzksmiewUCXX6qM
4KNKzv8nVvjPb+blAdNTypU5ZXY2PxFkq4t9wyvf6MjFvFJkkd1rTHJfbwqKmxgdhf0B2D+Fuq94
QWsF9n+tHHcH5yg5DQXwpwjOMIUdPNAwnLRBA/Y5k7fBcQnsppPpOGwI4iY116KJvH5KKXm5pLrz
ntZv1i1961sOskFWhYNaAGbCuNYSGrOhux6fLwI4Yfpqb8oXVYymrXLSWzGaRVjqKOzjDcXbvYWz
MYU800ifAb+7tr9iSEwgd5TPAoRQBRk14hFGao7uqHdeUyv4G8Z6IaXw5FRTqHX9b+55dbZTVk3j
LRFz/3REsfzRVmYr//6QYvMTdN+Kg/oFwBqYGN9IrGHMPGlvGJ6+ZklcnsC9Qz73+K9vskQlGR4A
O0TM66QiSywOZAHdLaJ2pU7WK3et45q9U/RbNwZb0uxWFfinsuwSdaY+PZ4eYh7Uu1rIXIPQsvCa
WihmkSmLTk0SRkWyoWS7B5zsJbZGiTsobUUaD861jW7qG78kSgDWrPZvMOwrSxO0atMI7M606Lul
X3fmwpeepvlo0UPMA53jGLYIzK93vvbmxSSBtZV7XG+Sh/scAHD0GKjFe/PBs2Vi6JFNr3GZ2fE0
xS1QTDsriokSMOvQa6+/BhHaB5GoaC6QUCwGX3N5/D8P9Kc73Jzy41W2KbpVcnEwaWATIfVQkDjk
lpdr/HmuSVMFDNW6xxD/wtFLXCo80nQ6y+IMoYD5hq+UEqMnv0byUm5Yz60wIAczRzPZ5WbXwL7M
XVp3XF67cSIySB4ApKW/E4cKepTj+Z0MpQuS1Ws7Th//sivggKmIiwkyck1eOiD4qSymGZ93D68/
E0TK0UkSNdZ0rDLrHds8aDfyI3rT6tLAb91Pes9tBn3mh/tjsSwwWBjF4O9BvXj2vz2QN6QBe4ss
urviG9hgUS3F1dqfamWTpS9gNT4L3DvDi3cm/7BRTI0qTpjq4QZMaAbMD6AIV2VqV4AxT1Be9zjE
qevUl1/rewl3etGltKQZmyuFQwzbLyLM1xQxi/03i2SqxbZGeWs25mjerKyv8khqwzlm4565EzVk
MAV0c3ZYPXVTjO9qTIT3HwwM1GBzeDLV4zhouzJN3RYXPPui9hJEyvF9XMUUQwF8bH5wOFvSzmu2
bX/VLb7JIlm95izWUWAUE5m4yEJcSeulFLPXjGJ3IycpjzEqJOepiRa5xSIAGYx6sGctO5XNRR0o
/v34IMDSPjjdMDg0hE1eagd4CtuNYKTcnJ1zMeLX4XJt5ABAG+QPRshFt60z8tvbfEhEUy7peGI/
PLMvSjjH+70RwRj4t6JYHcOcGPuHWoHFGWqa6tI7YM+NPjRNGtVynVyJ9qMEkrVtPgxDLj3VvOh+
hXt1oW4G2/NKbBdG0OqFSiCXjLRlrtG2J1LDKHKQ94sBbdBOr2k3rk6tMPkWGDLsMlsVL5Z/ZweY
A7QKAqLoJarUue1xJm7xV9pfNwzZc2JsHVt30EoH7Yj6IClxq0BgxWUJlqMmgJDCAvDGJagNmj4+
1g5LsS/LP4tsTqMCN17LAzvbfqzMHNoRlfBCGO3leZRU9ljpBemSgy/WTmoP3FfrUa2hKQccBZrd
PH+lcrlJ92blhKXfrwUZQrNqv6pfS3GiMcfAnBj3u5tbMi/Pg2lDyoiJ9hnvrvgjW1uxRcfzc0zM
MaDlOzv8dbDxNtzDQmAp0cq5r2iArthj7iGksfg35gI+zX3gUhmerbOQB5AOrteSNHJGZu1eVchu
w49vcE0Qfk64Sr2R8vkszwsDLXpZ9KqlouDgvzGSaiX35fbTMbKNwxqUkA3ijFscA1BQA75vZ9tS
8L10YmT3aKfVQZmJ06oUzQBzN2i26UMDubCHfbkNfEjQDG3p/mDCRo2s2yDPBU059bNKz+2bR4aB
lqtsirwjekl7bbiveaeD22h2cSCb1JsA+yC1gTgiyH+SzBO7cz5pZicwBVklaBNkRs2DB2Thc+5Q
Qzp4qE9oJALrJrB6F1EbB0lmAYjCp+01Xx4KXPIN7l3mJSKMDCqocW9TNc9EIfLGXCFgzOXS/5vh
Jg7qsltLnTOtbH+M8np1o4JpWL0kfB2roYSeI5PiqjonER3Lwtz9c7G+4ldXjiWLJqdzw2isDQcD
2Z2x6BH69HFU/P65t7UFDDtyKlxTE8cOy2Sg0KP5TV9jhxc7K+Dtyz/hf9wyNANz0oKkyWMfR47U
Yx2y/i72fwn5Z/Jf20CYvHGMhLWZxMStorElEEzDiCAKBkgXUsxNrEgp+K2vWlOFCjSqi/eJhZVG
WdrJ/zJ9vZR94/t8vQTaPb3Rl778JYozV+8GHXK6zyIUVWQpfZL7keljtKZ/BK+F0EhbfuyAHkFa
DfdsbvWaKVyBLw5fef/7v929HJee3nS+ZYxj57tGu/ZXlELkz9Ou6D4eWrbTq5bvgMMgNQUfhFFn
vP8ZiURgnSbE3FVXJpHLox8oZUJeIVKVy3kUDPOqO9upJE+n37t4p5fDak8x5EpQScJ4agfraeC1
iaJe+t4sKFcPtvhFr1T0T/9cW44rfAKGhizKpq6jsbEqN/30He2uGHrVooC9jQmzLrj5H0+ideqd
W4AsWDNbOyLvBm6Yz93U1rSO2hQ/VW5bHoReeFsB9Zy7Zhq0j2ND+fZhfCtmm9O0C5FGSIrXG9h4
P8BsOPzwkWN+8PbLAMp2sT6NsVzXYgjfEwUBaDMf95tCZ2oGe/LYQ1wUfwijl7fmgnTOtFV8ydRx
NmBz+awo7Bk2JFPcjgzvOXZdTb5P5UehUgKzUPXVuMaa5aq6YgDVBkH0vhZ611NzFlnTCPA1e94N
HEGwMN0c4m39lqMqGrwneCGtoK9q1/ghtwnAPm41c6gM+gvuDaukz6FKjRY5KjMZP6U4EYJ5a1Q3
DAkC9SMh+ejj9L+rbWTAaTVIyDvrTAzWM8FFQqWwNoOZ3moc1gLKap8gDTGun61ymwf5qP0qhQ6U
pcj0FwpjJJXpVZE5m7U82+mOspmj7XC9yuEE6rBR0MgtQDmNOoaoHRA+xiLyMvH43CcdVNclUjOP
YNSnLTj+848xYQdl12+0RGf44Bb4bn3xi0iHrDWmd7mm6ueTJDcIGfcLom83gDe26hTon5TgnBxK
5KNil8KE3R+MNN9Tl5qiE4TsWQ14H6W3Yu4hoBrMCm5HZkDeTT9ME5ttgL1GvGByUfpMoazfZdxb
j6dFsdqvm/VUgTekxfknFN5ytLHnTn6pqfAehEUbrn6vryDm213LPDOe8O+q2booPjxCJcqaGSpT
LimLdFBGPSiTp7vqb1P3su2c9Dq3TpfA6PF0bVH9zFie2/Bay2Mody+fALnNKsZfm3Ojr56douWG
ubuPaDT9iTap9egKlDkz96G+KKZEWrD2ac2xGD+xU2jvsS0xi34v8jPvhXuuHVQDWvuoWIBFpkX0
rl7Ts9olSGjBT3hHv30aGCWuE+nD0dKLXUpBh2I4I9vXrm6CvWbtYupm20WDGz3RzMl64vRwVuV5
ukFVBTfkoPoMNujwWpeJIHgwOzc+GzEPIRL6Tg7UK2qRwsNz1fpk86dpAqYuY23DKfu+8JuGCJ5s
s2zvMuAJU01Sbqa77b4BC7v+SDiRdhuWcvzsTjNiDixQJhn4+jDksxKYRaF2gqcOsQuS/DhMDR/L
QEWEecqxGwtwiALOUeoAHQct8LkZus5neLvviIG3PuOuqkgruZzlG2sXJT7+DTm+fYQKM+v210yK
pa2IT09ZuyNdi44Id6sHukAl0eZIr//FOu1ph6higjqH7SciqFpRiLNrF9TqMZOL27WyVyF4Hahb
qKYvS+VKgWmMN+He829/ApL3lEM48Clg7eOzWsVQ7t7xk5kZNDeqv9X/usbSXb3UUGFsd1CvSJ8I
VtlQ3mrqC/fOvpcnqOzPrmMyBIEVDCyuZFiqNsZdxPsGZm9ajbXoYssfJeEUTbmxh4snA9fXWmjM
mLAeYQB4vtvMP8Ap//ntfytuaA2rwUfNmOsuF6Ci+u+lRp1N6WWN97s8e3sfRqu3zNLsAnj1maiU
a5OhvLG2m0+FTnSboVTvE5Zg9TQxuDg4D0XUaAEcLdnqaVvYrO1pM+Zf6dGUllk9H9jD5uJzC/Nr
XQ61evSHX7d2/JsRLb2S3y8R9T6jF4+Mjeh49LGnd2SkfifczWqZ9Pl0DEp7Nbn7WCuvD/9ekBiV
ekGgHX1xEtXljdEE7bp5IO8t7ouhO7n/0XZpuTceZ+voGTKSX6rA93QncSv9jSoFVWj/Sln4uvT1
LbYKiEx/BUYD+jxfYNJaYqBKhJNQbtVHocPKAYtxkSkh8kSCFGGzPfkfMxm5eP5pLv14EIz+u160
i7Rk3mOwGHEIniYTYFbBjKwRpP4ZGcFCmz2xg1R0IkdGZmhuJyVb2fy21XapVUx+Aqvq+Tl4a37s
BUkty4JGFMbI3BWJtf2+SpBE/yLqcIybV90IFf46kUEROEGvTnOySR5W3EDH22+uLiuQYufKFtSg
f9RuX4OROpxGiwDbk/8XjgYzNNVkRz7Pu6qpCaCpGjq4llQOmYI0jCoIdfoQV9VFkVG+RcgZvyJW
fAafsyq9oOIQCmSQrdtjez3C3x8N7Y7QXijQD8aFMvmlHAH8LJhYZaL84cfMoYA+3Si330qN7Rdz
haozQ/H98Ci8FLp1uHr0qN70gVOGDH4tzyPZ+qj6VTrnZbZb2nFUmNh/aFsOT4YqW8UsqNddLea7
45zbPXXvQrGTJyw1puPzINaQ82R4chfBV1+4bMAIPafbgWRMUtf2tjbI4Bl9FOpMxDHjHp2Z5Hj6
78OYR7/XMHix1mA4q50YFxv21SFXrF9l8QqVhIKHbno7WfK+f/kX4zqpyfdvKP78V7fWiAkVUl6n
QtBRaAZ48EHkDaMEDH8xf6RgKW5sHkDVT6BB8SFJLfTWZdYZdWAZFJ2ZHT0TIM4yX/1fzMftYrzj
11g0blvQpMhY8+CVCoBYCpHHl8TQy+/nNHWMu0Aso0R3qtr05VXyi3QiwLaxgNz5xbFztfo/vFQI
KgVaLcthA/W2bSgjmvdSh4b3oal7WKq0tGC6M5jCMFngKGc/Nl9a01/a9Ia+2bu+A6S1eNUIamen
FcoyOOF4UB7zw0r9ZR70f/hdivBylSbRQKu9H0iH/LIAVQ5Ev/u/D0S9K2V5LFxmE+jOrsmsYFEb
70+Ve5dY9sEt01v0iXphZUPg5+W3GIptzE3XC/cl1xjxhP6J6GCosuPSECgNO4ngw/1J14pCjeyT
QQEbdzG9EpNiuUSLahlmYSnVmr0jq4wksTXMnaQ40xhT73dnnskIi9lYdsXU0Gl9mZMbS9KqGAXv
Rz1XYavneN2GopAGbWU0q1SqRRFfGXpM2QI5aBXRvZdNSEXLoC8biagL0Imk9J4QfGSr33OlrbsN
gf/fpmbE6UzAvLe2bHJZGXL3KyhicwkX6JEFK2nWLfCQC294ZvUtJDcbv/547Z1DVS3oY5Iv2i0J
gjJNUXA8fYS4UISZpg0fiK2f28H+ZWDU1YGKCsvzQjkNDjA/QgpCPFtcieDUj6Dot5kREfrEyuvn
HY6GeVWv8RyclmJJCdIQ4bBR2eAYjhkNNwgedF8hrO/2+JpPEHNMVcroEsF2zUUodYmQ4rKX4S/W
m32tA+i+9j02zHAVFT4xDOYV/Fts86OACq0zTYWM6a2CjiP2C49JrPkwtRciQju7JUZq3BNfBnhe
gpPHrK9ghWVDOF7gqrc1BM8iPiRE7NuTdlzlIm6sEAFkrw4nR9Mu8/Som6PaOHLziT1tw21ZCP4k
4JF2mv9qtMBzktx9bDl3SaTHY7xLpdMjVkK805j0xS8FA2MIaIrhvUuJug7QV3SODgmzkIxZxr/F
NVxYS5NCjXP2VWYf5Xsgv2QIpYodcFlSxwBHHMaKcoMDn0HnfE8ufRvNsMxcewhC7xIABNoMYTWG
4PM9btbkZUyU5ePZoJLl7XNMUN+OO3NEgLPRipf+QtepnxynSfoLgPGWqGQc7vkF1FldNJNK03uT
ZPbPPVTul9cHzIhlsvnr4EDCSqEu2Hs8U4X9kLJJDXKbrn6I/2TDCXp6Sn4IuMgfhzRe/GidQp19
GJbJosNoH214BSz2M0MzBnS+FPvC8S6yegUlVlsE//8vMTWlRfyAEt1rSlEfUjzH/sshl0TbTFW1
MEKLX9D7ZYoEe01eyPBmMBQNzuWfjDkezCHt9m6JRk+MmKgGLCiq74GZuNZmLkc4t/SxyB9F5pYK
68klyqG3jcaUbmZ3VF2yd2224Iyx9SegnTTF+EP67ebur2H1bgWN00V6SgVO9kHm+c/ZNpwYL8Hw
yQ+5zKi7vX8ZJOZx9/oYgWDP3Myg5l1I//gFGzG8z2PyVw5T7SmMQV06aViMzXLzIccVNQG0efIB
qk06iSAXrmp00NZimYA8EVJwukZOuyEG4lujG9rLZhm9n+yPyicX3vBUE2Q3ZW1a99mBp0cd5pu5
o1evF6u5GkuB0xhQeh4afY0huPpFuLCyXXbbWe7fROKUydO3Nq6SxZ6FzhvvFBksNJ4hnq8vs7Yz
Xt4cqdSUMpmH3GQiLU5XsqS5fcuzWKRc0rgP6OKdQfk9l3IA/k75UXWKNwCCUVFvWxyATlevrDXT
bbkD6Nn7bChCoRW6H2u2gP3Fg/SzqdVsLEHP3id1WJBqPMfPdHfvmgV1es2eRsBBc5Xz43b1TWj0
furnV97RiKoTT2GHh+P1Q68xv2tGn48RP+G9tEQKjVUtTSoT6AVHJyuH4lvIB3jt3xU8Via+fH+1
SP1EGp2uH68cA7SaPlzpVHWMfTUTytoiBzZmKjakEpVmu5qXzfdnqcpHt1OM4iq040mfScJkm00Z
lElKQb7AcSKIlDyXCKWYFzrzmnU4/x1jemGdxBkwW6tWCcCwM0Zc/3mI8V4utzeG8uhVbbS3B9EM
+UmG0UwFV14AhRytrQIr6B4MsVFmxRBTDRWNU/g2OBdvoSr9Ev1ZCGtAEO4Opx2N6tU8nX0n1Gc+
n9gtfFEdNgFt7mlWdB7UYJeQsYIZJfKsIHgDP3iywp12Wq17s7HC3YJ+TFhyDnsoJ196hPhn65AO
OrVIjxCadahuxPhNIfhQANRvipsW5TCsvNK8hQIySdEVhXI1IkNPvPhj1OUzSj9t55AkwjN0Orc6
GWuZQ6nSeJYwdD6ghGckfTJfV3WLKOeaB1/XGDfOKbJG8M259bHSl51L6Ka16QyYf7JptR37sSYj
t51YJqlhevbdkkWM+b3p1RuyrFd3P/GHOee8Xq2F0dHZhy3pb/pN1ankjfr/9kY7aG6Oj0oaPC2O
Cfp0lrT66sLnSbhGD10kY3Ub77LCRiaUl1KMVpsDXadVVVeRRcNr21PEjdpZtsyUnRMujH+xyxsP
ZVM+//Mk7QFD4mF+F7FBLRjszkwJte92g/7FMpZb64TT8F2hIbz7Ds6sH4DkJl/03KW3GaXWNFZN
5PikjF744D8VwlPyByDj3JvyccZpsBfpDdBnWaYGFpc2manNa4gHEAxs6Gk3OvWVKoaW9uxeQWQf
/JY4Eac/JoONpImo505N1UUIaE2Tz5qi3K9yDBz10WhPBzHY0axMYDvhj3DSLF74vDakFa9noS5i
RjuCTNnsxHYQFC2xi7xhaErmBfjYWV1IvgRLdFm5L8AjKNftIVtWHcq/GDlTSO6DiKA6iNHNCUZ4
c28UaYSoNXtYSm1iYrtYgQapzHujsZRUgkrMR4YUaeDL8fzWoIWXWLVcs3v7zqsfXYiT6H81WcWw
E5ZtH8ktNmYjqP7eArRNdVJh7LT4Ne3NmgH8EZt1dmI2oKqyyD8DBMD+WuPHEqejPfXkM+H+Mbh/
HRYbUXdP0+aBWULWjmBI1LXX85oT9P1Xg9LGBVzH04trIX40xBXimziwM1jEzY2SdXUEHQQTpSg/
ioXhvc8Po8DW1TH0kuta8GquJksq8Xf0JNSBCNff7ghuD6PKLFE/AX/9KPqbfxRoRnLoOZMVQ9ek
7c3maLALOTo62AJKdL1qnrNlKm65ys1Fs2yijapOWVMXFSdZfzFVb8lfRbDX3L6sVrsObzDLVIsV
ob386bmd+1Eqo0G9gk/TS8268UbmEaksofweNitYv+ylpSDoY/YomSQW3nhfyUbiEt3ISKZj5+g8
eLyghhgFf0gtg2kxBqPNvyPzCbW8ipH9cgop+v1xtZlILpHY/k6/Z6DGw+/BEA==
`protect end_protected

