-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.2
--  \   \         Application : 7 Series FPGAs Transceivers Wizard
--  /   /         Filename : gt6_rtm34l_multi_gt.vhd
-- /___/   /\     
-- \   \  /  \ 
--  \___\/\___\
--
--
-- Module gt6_rtm34l_multi_gt (a Multi GT Wrapper)
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***************************** Entity Declaration ****************************

entity gt6_rtm34l_multi_gt is
generic
(

    -- Simulation attributes
    EXAMPLE_SIMULATION             : integer  := 0;      -- Set to 1 for simulation
    WRAPPER_SIM_GTRESET_SPEEDUP    : string   := "FALSE" -- Set to "TRUE" to speed up sim reset
);
port
(
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y0)
    --____________________________CHANNEL PORTS________________________________
 GT0_RXPMARESETDONE_OUT  : out  std_logic;
 GT0_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt0_cpllfbclklost_out                   : out  std_logic;
    gt0_cplllock_out                        : out  std_logic;
    gt0_cplllockdetclk_in                   : in   std_logic;
    gt0_cpllrefclklost_out                  : out  std_logic;
    gt0_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt0_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxbyteisaligned_out                 : out  std_logic;
    gt0_rxmcommaalignen_in                  : in   std_logic;
    gt0_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxdfeagchold_in                     : in   std_logic;
    gt0_rxdfelfhold_in                      : in   std_logic;
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt0_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt0_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt0_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT1  (X0Y1)
    --____________________________CHANNEL PORTS________________________________
 GT1_RXPMARESETDONE_OUT  : out  std_logic;
 GT1_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt1_cpllfbclklost_out                   : out  std_logic;
    gt1_cplllock_out                        : out  std_logic;
    gt1_cplllockdetclk_in                   : in   std_logic;
    gt1_cpllrefclklost_out                  : out  std_logic;
    gt1_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt1_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpclk_in                           : in   std_logic;
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxbyteisaligned_out                 : out  std_logic;
    gt1_rxmcommaalignen_in                  : in   std_logic;
    gt1_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxdfeagchold_in                     : in   std_logic;
    gt1_rxdfelfhold_in                      : in   std_logic;
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt1_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt1_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt1_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT2  (X0Y2)
    --____________________________CHANNEL PORTS________________________________
 GT2_RXPMARESETDONE_OUT  : out  std_logic;
 GT2_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt2_cpllfbclklost_out                   : out  std_logic;
    gt2_cplllock_out                        : out  std_logic;
    gt2_cplllockdetclk_in                   : in   std_logic;
    gt2_cpllrefclklost_out                  : out  std_logic;
    gt2_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt2_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpclk_in                           : in   std_logic;
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxbyteisaligned_out                 : out  std_logic;
    gt2_rxmcommaalignen_in                  : in   std_logic;
    gt2_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxdfeagchold_in                     : in   std_logic;
    gt2_rxdfelfhold_in                      : in   std_logic;
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt2_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt2_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt2_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT3  (X0Y3)
    --____________________________CHANNEL PORTS________________________________
 GT3_RXPMARESETDONE_OUT  : out  std_logic;
 GT3_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt3_cpllfbclklost_out                   : out  std_logic;
    gt3_cplllock_out                        : out  std_logic;
    gt3_cplllockdetclk_in                   : in   std_logic;
    gt3_cpllrefclklost_out                  : out  std_logic;
    gt3_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt3_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpclk_in                           : in   std_logic;
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxbyteisaligned_out                 : out  std_logic;
    gt3_rxmcommaalignen_in                  : in   std_logic;
    gt3_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxdfeagchold_in                     : in   std_logic;
    gt3_rxdfelfhold_in                      : in   std_logic;
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt3_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt3_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt3_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT4  (X0Y4)
    --____________________________CHANNEL PORTS________________________________
 GT4_RXPMARESETDONE_OUT  : out  std_logic;
 GT4_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt4_cpllfbclklost_out                   : out  std_logic;
    gt4_cplllock_out                        : out  std_logic;
    gt4_cplllockdetclk_in                   : in   std_logic;
    gt4_cpllrefclklost_out                  : out  std_logic;
    gt4_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt4_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt4_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt4_drpclk_in                           : in   std_logic;
    gt4_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt4_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt4_drpen_in                            : in   std_logic;
    gt4_drprdy_out                          : out  std_logic;
    gt4_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt4_eyescanreset_in                     : in   std_logic;
    gt4_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt4_eyescandataerror_out                : out  std_logic;
    gt4_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt4_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt4_rxusrclk_in                         : in   std_logic;
    gt4_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt4_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt4_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt4_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt4_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt4_rxbyteisaligned_out                 : out  std_logic;
    gt4_rxmcommaalignen_in                  : in   std_logic;
    gt4_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt4_rxdfeagchold_in                     : in   std_logic;
    gt4_rxdfelfhold_in                      : in   std_logic;
    gt4_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt4_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt4_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt4_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt4_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt4_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt4_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt4_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt4_gttxreset_in                        : in   std_logic;
    gt4_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt4_txusrclk_in                         : in   std_logic;
    gt4_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt4_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt4_gthtxn_out                          : out  std_logic;
    gt4_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt4_txoutclk_out                        : out  std_logic;
    gt4_txoutclkfabric_out                  : out  std_logic;
    gt4_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt4_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt4_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt4_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT5  (X0Y5)
    --____________________________CHANNEL PORTS________________________________
 GT5_RXPMARESETDONE_OUT  : out  std_logic;
 GT5_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt5_cpllfbclklost_out                   : out  std_logic;
    gt5_cplllock_out                        : out  std_logic;
    gt5_cplllockdetclk_in                   : in   std_logic;
    gt5_cpllrefclklost_out                  : out  std_logic;
    gt5_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt5_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt5_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt5_drpclk_in                           : in   std_logic;
    gt5_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt5_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt5_drpen_in                            : in   std_logic;
    gt5_drprdy_out                          : out  std_logic;
    gt5_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt5_eyescanreset_in                     : in   std_logic;
    gt5_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt5_eyescandataerror_out                : out  std_logic;
    gt5_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt5_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt5_rxusrclk_in                         : in   std_logic;
    gt5_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt5_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt5_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt5_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt5_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt5_rxbyteisaligned_out                 : out  std_logic;
    gt5_rxmcommaalignen_in                  : in   std_logic;
    gt5_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt5_rxdfeagchold_in                     : in   std_logic;
    gt5_rxdfelfhold_in                      : in   std_logic;
    gt5_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt5_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt5_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt5_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt5_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt5_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt5_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt5_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt5_gttxreset_in                        : in   std_logic;
    gt5_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt5_txusrclk_in                         : in   std_logic;
    gt5_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt5_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt5_gthtxn_out                          : out  std_logic;
    gt5_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt5_txoutclk_out                        : out  std_logic;
    gt5_txoutclkfabric_out                  : out  std_logic;
    gt5_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt5_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt5_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt5_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT6  (X0Y6)
    --____________________________CHANNEL PORTS________________________________
 GT6_RXPMARESETDONE_OUT  : out  std_logic;
 GT6_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt6_cpllfbclklost_out                   : out  std_logic;
    gt6_cplllock_out                        : out  std_logic;
    gt6_cplllockdetclk_in                   : in   std_logic;
    gt6_cpllrefclklost_out                  : out  std_logic;
    gt6_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt6_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt6_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt6_drpclk_in                           : in   std_logic;
    gt6_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt6_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt6_drpen_in                            : in   std_logic;
    gt6_drprdy_out                          : out  std_logic;
    gt6_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt6_eyescanreset_in                     : in   std_logic;
    gt6_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt6_eyescandataerror_out                : out  std_logic;
    gt6_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt6_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt6_rxusrclk_in                         : in   std_logic;
    gt6_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt6_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt6_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt6_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt6_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt6_rxbyteisaligned_out                 : out  std_logic;
    gt6_rxmcommaalignen_in                  : in   std_logic;
    gt6_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt6_rxdfeagchold_in                     : in   std_logic;
    gt6_rxdfelfhold_in                      : in   std_logic;
    gt6_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt6_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt6_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt6_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt6_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt6_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt6_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt6_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt6_gttxreset_in                        : in   std_logic;
    gt6_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt6_txusrclk_in                         : in   std_logic;
    gt6_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt6_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt6_gthtxn_out                          : out  std_logic;
    gt6_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt6_txoutclk_out                        : out  std_logic;
    gt6_txoutclkfabric_out                  : out  std_logic;
    gt6_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt6_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt6_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt6_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT7  (X0Y7)
    --____________________________CHANNEL PORTS________________________________
 GT7_RXPMARESETDONE_OUT  : out  std_logic;
 GT7_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt7_cpllfbclklost_out                   : out  std_logic;
    gt7_cplllock_out                        : out  std_logic;
    gt7_cplllockdetclk_in                   : in   std_logic;
    gt7_cpllrefclklost_out                  : out  std_logic;
    gt7_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt7_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt7_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt7_drpclk_in                           : in   std_logic;
    gt7_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt7_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt7_drpen_in                            : in   std_logic;
    gt7_drprdy_out                          : out  std_logic;
    gt7_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt7_eyescanreset_in                     : in   std_logic;
    gt7_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt7_eyescandataerror_out                : out  std_logic;
    gt7_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt7_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt7_rxusrclk_in                         : in   std_logic;
    gt7_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt7_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt7_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt7_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt7_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt7_rxbyteisaligned_out                 : out  std_logic;
    gt7_rxmcommaalignen_in                  : in   std_logic;
    gt7_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt7_rxdfeagchold_in                     : in   std_logic;
    gt7_rxdfelfhold_in                      : in   std_logic;
    gt7_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt7_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt7_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt7_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt7_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt7_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt7_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt7_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt7_gttxreset_in                        : in   std_logic;
    gt7_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt7_txusrclk_in                         : in   std_logic;
    gt7_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt7_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt7_gthtxn_out                          : out  std_logic;
    gt7_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt7_txoutclk_out                        : out  std_logic;
    gt7_txoutclkfabric_out                  : out  std_logic;
    gt7_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt7_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt7_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt7_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT8  (X0Y8)
    --____________________________CHANNEL PORTS________________________________
 GT8_RXPMARESETDONE_OUT  : out  std_logic;
 GT8_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt8_cpllfbclklost_out                   : out  std_logic;
    gt8_cplllock_out                        : out  std_logic;
    gt8_cplllockdetclk_in                   : in   std_logic;
    gt8_cpllrefclklost_out                  : out  std_logic;
    gt8_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt8_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt8_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt8_drpclk_in                           : in   std_logic;
    gt8_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt8_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt8_drpen_in                            : in   std_logic;
    gt8_drprdy_out                          : out  std_logic;
    gt8_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt8_eyescanreset_in                     : in   std_logic;
    gt8_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt8_eyescandataerror_out                : out  std_logic;
    gt8_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt8_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt8_rxusrclk_in                         : in   std_logic;
    gt8_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt8_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt8_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt8_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt8_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt8_rxbyteisaligned_out                 : out  std_logic;
    gt8_rxmcommaalignen_in                  : in   std_logic;
    gt8_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt8_rxdfeagchold_in                     : in   std_logic;
    gt8_rxdfelfhold_in                      : in   std_logic;
    gt8_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt8_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt8_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt8_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt8_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt8_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt8_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt8_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt8_gttxreset_in                        : in   std_logic;
    gt8_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt8_txusrclk_in                         : in   std_logic;
    gt8_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt8_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt8_gthtxn_out                          : out  std_logic;
    gt8_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt8_txoutclk_out                        : out  std_logic;
    gt8_txoutclkfabric_out                  : out  std_logic;
    gt8_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt8_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt8_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt8_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT9  (X0Y9)
    --____________________________CHANNEL PORTS________________________________
 GT9_RXPMARESETDONE_OUT  : out  std_logic;
 GT9_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt9_cpllfbclklost_out                   : out  std_logic;
    gt9_cplllock_out                        : out  std_logic;
    gt9_cplllockdetclk_in                   : in   std_logic;
    gt9_cpllrefclklost_out                  : out  std_logic;
    gt9_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt9_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt9_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt9_drpclk_in                           : in   std_logic;
    gt9_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt9_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt9_drpen_in                            : in   std_logic;
    gt9_drprdy_out                          : out  std_logic;
    gt9_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt9_eyescanreset_in                     : in   std_logic;
    gt9_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt9_eyescandataerror_out                : out  std_logic;
    gt9_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt9_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt9_rxusrclk_in                         : in   std_logic;
    gt9_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt9_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt9_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt9_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt9_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt9_rxbyteisaligned_out                 : out  std_logic;
    gt9_rxmcommaalignen_in                  : in   std_logic;
    gt9_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt9_rxdfeagchold_in                     : in   std_logic;
    gt9_rxdfelfhold_in                      : in   std_logic;
    gt9_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt9_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt9_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt9_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt9_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt9_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt9_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt9_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt9_gttxreset_in                        : in   std_logic;
    gt9_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt9_txusrclk_in                         : in   std_logic;
    gt9_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt9_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt9_gthtxn_out                          : out  std_logic;
    gt9_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt9_txoutclk_out                        : out  std_logic;
    gt9_txoutclkfabric_out                  : out  std_logic;
    gt9_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt9_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt9_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt9_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT10  (X0Y10)
    --____________________________CHANNEL PORTS________________________________
 GT10_RXPMARESETDONE_OUT  : out  std_logic;
 GT10_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt10_cpllfbclklost_out                  : out  std_logic;
    gt10_cplllock_out                       : out  std_logic;
    gt10_cplllockdetclk_in                  : in   std_logic;
    gt10_cpllrefclklost_out                 : out  std_logic;
    gt10_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt10_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt10_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt10_drpclk_in                          : in   std_logic;
    gt10_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt10_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt10_drpen_in                           : in   std_logic;
    gt10_drprdy_out                         : out  std_logic;
    gt10_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt10_eyescanreset_in                    : in   std_logic;
    gt10_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt10_eyescandataerror_out               : out  std_logic;
    gt10_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt10_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt10_rxusrclk_in                        : in   std_logic;
    gt10_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt10_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt10_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt10_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt10_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt10_rxbyteisaligned_out                : out  std_logic;
    gt10_rxmcommaalignen_in                 : in   std_logic;
    gt10_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt10_rxdfeagchold_in                    : in   std_logic;
    gt10_rxdfelfhold_in                     : in   std_logic;
    gt10_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt10_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt10_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt10_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt10_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt10_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt10_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt10_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt10_gttxreset_in                       : in   std_logic;
    gt10_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt10_txusrclk_in                        : in   std_logic;
    gt10_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt10_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt10_gthtxn_out                         : out  std_logic;
    gt10_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt10_txoutclk_out                       : out  std_logic;
    gt10_txoutclkfabric_out                 : out  std_logic;
    gt10_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt10_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt10_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt10_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT11  (X0Y11)
    --____________________________CHANNEL PORTS________________________________
 GT11_RXPMARESETDONE_OUT  : out  std_logic;
 GT11_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt11_cpllfbclklost_out                  : out  std_logic;
    gt11_cplllock_out                       : out  std_logic;
    gt11_cplllockdetclk_in                  : in   std_logic;
    gt11_cpllrefclklost_out                 : out  std_logic;
    gt11_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt11_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt11_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt11_drpclk_in                          : in   std_logic;
    gt11_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt11_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt11_drpen_in                           : in   std_logic;
    gt11_drprdy_out                         : out  std_logic;
    gt11_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt11_eyescanreset_in                    : in   std_logic;
    gt11_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt11_eyescandataerror_out               : out  std_logic;
    gt11_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt11_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt11_rxusrclk_in                        : in   std_logic;
    gt11_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt11_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt11_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt11_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt11_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt11_rxbyteisaligned_out                : out  std_logic;
    gt11_rxmcommaalignen_in                 : in   std_logic;
    gt11_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt11_rxdfeagchold_in                    : in   std_logic;
    gt11_rxdfelfhold_in                     : in   std_logic;
    gt11_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt11_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt11_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt11_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt11_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt11_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt11_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt11_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt11_gttxreset_in                       : in   std_logic;
    gt11_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt11_txusrclk_in                        : in   std_logic;
    gt11_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt11_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt11_gthtxn_out                         : out  std_logic;
    gt11_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt11_txoutclk_out                       : out  std_logic;
    gt11_txoutclkfabric_out                 : out  std_logic;
    gt11_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt11_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt11_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt11_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT12  (X0Y12)
    --____________________________CHANNEL PORTS________________________________
 GT12_RXPMARESETDONE_OUT  : out  std_logic;
 GT12_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt12_cpllfbclklost_out                  : out  std_logic;
    gt12_cplllock_out                       : out  std_logic;
    gt12_cplllockdetclk_in                  : in   std_logic;
    gt12_cpllrefclklost_out                 : out  std_logic;
    gt12_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt12_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt12_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt12_drpclk_in                          : in   std_logic;
    gt12_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt12_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt12_drpen_in                           : in   std_logic;
    gt12_drprdy_out                         : out  std_logic;
    gt12_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt12_eyescanreset_in                    : in   std_logic;
    gt12_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt12_eyescandataerror_out               : out  std_logic;
    gt12_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt12_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt12_rxusrclk_in                        : in   std_logic;
    gt12_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt12_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt12_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt12_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt12_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt12_rxbyteisaligned_out                : out  std_logic;
    gt12_rxmcommaalignen_in                 : in   std_logic;
    gt12_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt12_rxdfeagchold_in                    : in   std_logic;
    gt12_rxdfelfhold_in                     : in   std_logic;
    gt12_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt12_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt12_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt12_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt12_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt12_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt12_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt12_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt12_gttxreset_in                       : in   std_logic;
    gt12_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt12_txusrclk_in                        : in   std_logic;
    gt12_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt12_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt12_gthtxn_out                         : out  std_logic;
    gt12_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt12_txoutclk_out                       : out  std_logic;
    gt12_txoutclkfabric_out                 : out  std_logic;
    gt12_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt12_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt12_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt12_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT13  (X0Y13)
    --____________________________CHANNEL PORTS________________________________
 GT13_RXPMARESETDONE_OUT  : out  std_logic;
 GT13_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt13_cpllfbclklost_out                  : out  std_logic;
    gt13_cplllock_out                       : out  std_logic;
    gt13_cplllockdetclk_in                  : in   std_logic;
    gt13_cpllrefclklost_out                 : out  std_logic;
    gt13_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt13_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt13_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt13_drpclk_in                          : in   std_logic;
    gt13_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt13_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt13_drpen_in                           : in   std_logic;
    gt13_drprdy_out                         : out  std_logic;
    gt13_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt13_eyescanreset_in                    : in   std_logic;
    gt13_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt13_eyescandataerror_out               : out  std_logic;
    gt13_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt13_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt13_rxusrclk_in                        : in   std_logic;
    gt13_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt13_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt13_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt13_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt13_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt13_rxbyteisaligned_out                : out  std_logic;
    gt13_rxmcommaalignen_in                 : in   std_logic;
    gt13_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt13_rxdfeagchold_in                    : in   std_logic;
    gt13_rxdfelfhold_in                     : in   std_logic;
    gt13_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt13_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt13_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt13_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt13_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt13_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt13_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt13_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt13_gttxreset_in                       : in   std_logic;
    gt13_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt13_txusrclk_in                        : in   std_logic;
    gt13_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt13_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt13_gthtxn_out                         : out  std_logic;
    gt13_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt13_txoutclk_out                       : out  std_logic;
    gt13_txoutclkfabric_out                 : out  std_logic;
    gt13_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt13_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt13_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt13_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT14  (X0Y14)
    --____________________________CHANNEL PORTS________________________________
 GT14_RXPMARESETDONE_OUT  : out  std_logic;
 GT14_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt14_cpllfbclklost_out                  : out  std_logic;
    gt14_cplllock_out                       : out  std_logic;
    gt14_cplllockdetclk_in                  : in   std_logic;
    gt14_cpllrefclklost_out                 : out  std_logic;
    gt14_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt14_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt14_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt14_drpclk_in                          : in   std_logic;
    gt14_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt14_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt14_drpen_in                           : in   std_logic;
    gt14_drprdy_out                         : out  std_logic;
    gt14_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt14_eyescanreset_in                    : in   std_logic;
    gt14_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt14_eyescandataerror_out               : out  std_logic;
    gt14_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt14_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt14_rxusrclk_in                        : in   std_logic;
    gt14_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt14_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt14_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt14_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt14_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt14_rxbyteisaligned_out                : out  std_logic;
    gt14_rxmcommaalignen_in                 : in   std_logic;
    gt14_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt14_rxdfeagchold_in                    : in   std_logic;
    gt14_rxdfelfhold_in                     : in   std_logic;
    gt14_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt14_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt14_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt14_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt14_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt14_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt14_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt14_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt14_gttxreset_in                       : in   std_logic;
    gt14_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt14_txusrclk_in                        : in   std_logic;
    gt14_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt14_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt14_gthtxn_out                         : out  std_logic;
    gt14_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt14_txoutclk_out                       : out  std_logic;
    gt14_txoutclkfabric_out                 : out  std_logic;
    gt14_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt14_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt14_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt14_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT15  (X0Y15)
    --____________________________CHANNEL PORTS________________________________
 GT15_RXPMARESETDONE_OUT  : out  std_logic;
 GT15_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt15_cpllfbclklost_out                  : out  std_logic;
    gt15_cplllock_out                       : out  std_logic;
    gt15_cplllockdetclk_in                  : in   std_logic;
    gt15_cpllrefclklost_out                 : out  std_logic;
    gt15_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt15_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt15_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt15_drpclk_in                          : in   std_logic;
    gt15_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt15_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt15_drpen_in                           : in   std_logic;
    gt15_drprdy_out                         : out  std_logic;
    gt15_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt15_eyescanreset_in                    : in   std_logic;
    gt15_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt15_eyescandataerror_out               : out  std_logic;
    gt15_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt15_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt15_rxusrclk_in                        : in   std_logic;
    gt15_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt15_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt15_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt15_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt15_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt15_rxbyteisaligned_out                : out  std_logic;
    gt15_rxmcommaalignen_in                 : in   std_logic;
    gt15_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt15_rxdfeagchold_in                    : in   std_logic;
    gt15_rxdfelfhold_in                     : in   std_logic;
    gt15_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt15_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt15_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt15_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt15_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt15_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt15_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt15_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt15_gttxreset_in                       : in   std_logic;
    gt15_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt15_txusrclk_in                        : in   std_logic;
    gt15_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt15_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt15_gthtxn_out                         : out  std_logic;
    gt15_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt15_txoutclk_out                       : out  std_logic;
    gt15_txoutclkfabric_out                 : out  std_logic;
    gt15_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt15_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt15_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt15_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT16  (X0Y16)
    --____________________________CHANNEL PORTS________________________________
 GT16_RXPMARESETDONE_OUT  : out  std_logic;
 GT16_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt16_cpllfbclklost_out                  : out  std_logic;
    gt16_cplllock_out                       : out  std_logic;
    gt16_cplllockdetclk_in                  : in   std_logic;
    gt16_cpllrefclklost_out                 : out  std_logic;
    gt16_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt16_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt16_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt16_drpclk_in                          : in   std_logic;
    gt16_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt16_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt16_drpen_in                           : in   std_logic;
    gt16_drprdy_out                         : out  std_logic;
    gt16_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt16_eyescanreset_in                    : in   std_logic;
    gt16_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt16_eyescandataerror_out               : out  std_logic;
    gt16_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt16_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt16_rxusrclk_in                        : in   std_logic;
    gt16_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt16_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt16_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt16_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt16_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt16_rxbyteisaligned_out                : out  std_logic;
    gt16_rxmcommaalignen_in                 : in   std_logic;
    gt16_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt16_rxdfeagchold_in                    : in   std_logic;
    gt16_rxdfelfhold_in                     : in   std_logic;
    gt16_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt16_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt16_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt16_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt16_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt16_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt16_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt16_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt16_gttxreset_in                       : in   std_logic;
    gt16_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt16_txusrclk_in                        : in   std_logic;
    gt16_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt16_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt16_gthtxn_out                         : out  std_logic;
    gt16_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt16_txoutclk_out                       : out  std_logic;
    gt16_txoutclkfabric_out                 : out  std_logic;
    gt16_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt16_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt16_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt16_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT17  (X0Y17)
    --____________________________CHANNEL PORTS________________________________
 GT17_RXPMARESETDONE_OUT  : out  std_logic;
 GT17_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt17_cpllfbclklost_out                  : out  std_logic;
    gt17_cplllock_out                       : out  std_logic;
    gt17_cplllockdetclk_in                  : in   std_logic;
    gt17_cpllrefclklost_out                 : out  std_logic;
    gt17_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt17_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt17_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt17_drpclk_in                          : in   std_logic;
    gt17_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt17_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt17_drpen_in                           : in   std_logic;
    gt17_drprdy_out                         : out  std_logic;
    gt17_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt17_eyescanreset_in                    : in   std_logic;
    gt17_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt17_eyescandataerror_out               : out  std_logic;
    gt17_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt17_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt17_rxusrclk_in                        : in   std_logic;
    gt17_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt17_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt17_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt17_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt17_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt17_rxbyteisaligned_out                : out  std_logic;
    gt17_rxmcommaalignen_in                 : in   std_logic;
    gt17_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt17_rxdfeagchold_in                    : in   std_logic;
    gt17_rxdfelfhold_in                     : in   std_logic;
    gt17_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt17_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt17_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt17_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt17_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt17_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt17_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt17_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt17_gttxreset_in                       : in   std_logic;
    gt17_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt17_txusrclk_in                        : in   std_logic;
    gt17_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt17_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt17_gthtxn_out                         : out  std_logic;
    gt17_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt17_txoutclk_out                       : out  std_logic;
    gt17_txoutclkfabric_out                 : out  std_logic;
    gt17_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt17_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt17_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt17_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT18  (X0Y18)
    --____________________________CHANNEL PORTS________________________________
 GT18_RXPMARESETDONE_OUT  : out  std_logic;
 GT18_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt18_cpllfbclklost_out                  : out  std_logic;
    gt18_cplllock_out                       : out  std_logic;
    gt18_cplllockdetclk_in                  : in   std_logic;
    gt18_cpllrefclklost_out                 : out  std_logic;
    gt18_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt18_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt18_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt18_drpclk_in                          : in   std_logic;
    gt18_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt18_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt18_drpen_in                           : in   std_logic;
    gt18_drprdy_out                         : out  std_logic;
    gt18_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt18_eyescanreset_in                    : in   std_logic;
    gt18_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt18_eyescandataerror_out               : out  std_logic;
    gt18_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt18_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt18_rxusrclk_in                        : in   std_logic;
    gt18_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt18_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt18_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt18_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt18_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt18_rxbyteisaligned_out                : out  std_logic;
    gt18_rxmcommaalignen_in                 : in   std_logic;
    gt18_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt18_rxdfeagchold_in                    : in   std_logic;
    gt18_rxdfelfhold_in                     : in   std_logic;
    gt18_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt18_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt18_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt18_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt18_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt18_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt18_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt18_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt18_gttxreset_in                       : in   std_logic;
    gt18_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt18_txusrclk_in                        : in   std_logic;
    gt18_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt18_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt18_gthtxn_out                         : out  std_logic;
    gt18_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt18_txoutclk_out                       : out  std_logic;
    gt18_txoutclkfabric_out                 : out  std_logic;
    gt18_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt18_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt18_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt18_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT19  (X0Y19)
    --____________________________CHANNEL PORTS________________________________
 GT19_RXPMARESETDONE_OUT  : out  std_logic;
 GT19_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt19_cpllfbclklost_out                  : out  std_logic;
    gt19_cplllock_out                       : out  std_logic;
    gt19_cplllockdetclk_in                  : in   std_logic;
    gt19_cpllrefclklost_out                 : out  std_logic;
    gt19_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt19_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt19_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt19_drpclk_in                          : in   std_logic;
    gt19_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt19_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt19_drpen_in                           : in   std_logic;
    gt19_drprdy_out                         : out  std_logic;
    gt19_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt19_eyescanreset_in                    : in   std_logic;
    gt19_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt19_eyescandataerror_out               : out  std_logic;
    gt19_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt19_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt19_rxusrclk_in                        : in   std_logic;
    gt19_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt19_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt19_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt19_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt19_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt19_rxbyteisaligned_out                : out  std_logic;
    gt19_rxmcommaalignen_in                 : in   std_logic;
    gt19_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt19_rxdfeagchold_in                    : in   std_logic;
    gt19_rxdfelfhold_in                     : in   std_logic;
    gt19_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt19_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt19_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt19_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt19_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt19_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt19_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt19_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt19_gttxreset_in                       : in   std_logic;
    gt19_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt19_txusrclk_in                        : in   std_logic;
    gt19_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt19_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt19_gthtxn_out                         : out  std_logic;
    gt19_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt19_txoutclk_out                       : out  std_logic;
    gt19_txoutclkfabric_out                 : out  std_logic;
    gt19_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt19_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt19_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt19_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT20  (X0Y20)
    --____________________________CHANNEL PORTS________________________________
 GT20_RXPMARESETDONE_OUT  : out  std_logic;
 GT20_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt20_cpllfbclklost_out                  : out  std_logic;
    gt20_cplllock_out                       : out  std_logic;
    gt20_cplllockdetclk_in                  : in   std_logic;
    gt20_cpllrefclklost_out                 : out  std_logic;
    gt20_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt20_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt20_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt20_drpclk_in                          : in   std_logic;
    gt20_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt20_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt20_drpen_in                           : in   std_logic;
    gt20_drprdy_out                         : out  std_logic;
    gt20_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt20_eyescanreset_in                    : in   std_logic;
    gt20_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt20_eyescandataerror_out               : out  std_logic;
    gt20_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt20_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt20_rxusrclk_in                        : in   std_logic;
    gt20_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt20_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt20_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt20_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt20_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt20_rxbyteisaligned_out                : out  std_logic;
    gt20_rxmcommaalignen_in                 : in   std_logic;
    gt20_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt20_rxdfeagchold_in                    : in   std_logic;
    gt20_rxdfelfhold_in                     : in   std_logic;
    gt20_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt20_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt20_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt20_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt20_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt20_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt20_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt20_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt20_gttxreset_in                       : in   std_logic;
    gt20_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt20_txusrclk_in                        : in   std_logic;
    gt20_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt20_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt20_gthtxn_out                         : out  std_logic;
    gt20_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt20_txoutclk_out                       : out  std_logic;
    gt20_txoutclkfabric_out                 : out  std_logic;
    gt20_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt20_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt20_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt20_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT21  (X0Y21)
    --____________________________CHANNEL PORTS________________________________
 GT21_RXPMARESETDONE_OUT  : out  std_logic;
 GT21_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt21_cpllfbclklost_out                  : out  std_logic;
    gt21_cplllock_out                       : out  std_logic;
    gt21_cplllockdetclk_in                  : in   std_logic;
    gt21_cpllrefclklost_out                 : out  std_logic;
    gt21_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt21_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt21_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt21_drpclk_in                          : in   std_logic;
    gt21_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt21_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt21_drpen_in                           : in   std_logic;
    gt21_drprdy_out                         : out  std_logic;
    gt21_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt21_eyescanreset_in                    : in   std_logic;
    gt21_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt21_eyescandataerror_out               : out  std_logic;
    gt21_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt21_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt21_rxusrclk_in                        : in   std_logic;
    gt21_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt21_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt21_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt21_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt21_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt21_rxbyteisaligned_out                : out  std_logic;
    gt21_rxmcommaalignen_in                 : in   std_logic;
    gt21_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt21_rxdfeagchold_in                    : in   std_logic;
    gt21_rxdfelfhold_in                     : in   std_logic;
    gt21_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt21_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt21_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt21_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt21_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt21_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt21_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt21_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt21_gttxreset_in                       : in   std_logic;
    gt21_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt21_txusrclk_in                        : in   std_logic;
    gt21_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt21_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt21_gthtxn_out                         : out  std_logic;
    gt21_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt21_txoutclk_out                       : out  std_logic;
    gt21_txoutclkfabric_out                 : out  std_logic;
    gt21_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt21_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt21_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt21_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT22  (X0Y22)
    --____________________________CHANNEL PORTS________________________________
 GT22_RXPMARESETDONE_OUT  : out  std_logic;
 GT22_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt22_cpllfbclklost_out                  : out  std_logic;
    gt22_cplllock_out                       : out  std_logic;
    gt22_cplllockdetclk_in                  : in   std_logic;
    gt22_cpllrefclklost_out                 : out  std_logic;
    gt22_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt22_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt22_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt22_drpclk_in                          : in   std_logic;
    gt22_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt22_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt22_drpen_in                           : in   std_logic;
    gt22_drprdy_out                         : out  std_logic;
    gt22_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt22_eyescanreset_in                    : in   std_logic;
    gt22_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt22_eyescandataerror_out               : out  std_logic;
    gt22_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt22_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt22_rxusrclk_in                        : in   std_logic;
    gt22_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt22_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt22_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt22_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt22_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt22_rxbyteisaligned_out                : out  std_logic;
    gt22_rxmcommaalignen_in                 : in   std_logic;
    gt22_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt22_rxdfeagchold_in                    : in   std_logic;
    gt22_rxdfelfhold_in                     : in   std_logic;
    gt22_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt22_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt22_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt22_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt22_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt22_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt22_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt22_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt22_gttxreset_in                       : in   std_logic;
    gt22_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt22_txusrclk_in                        : in   std_logic;
    gt22_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt22_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt22_gthtxn_out                         : out  std_logic;
    gt22_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt22_txoutclk_out                       : out  std_logic;
    gt22_txoutclkfabric_out                 : out  std_logic;
    gt22_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt22_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt22_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt22_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT23  (X0Y23)
    --____________________________CHANNEL PORTS________________________________
 GT23_RXPMARESETDONE_OUT  : out  std_logic;
 GT23_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt23_cpllfbclklost_out                  : out  std_logic;
    gt23_cplllock_out                       : out  std_logic;
    gt23_cplllockdetclk_in                  : in   std_logic;
    gt23_cpllrefclklost_out                 : out  std_logic;
    gt23_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt23_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt23_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt23_drpclk_in                          : in   std_logic;
    gt23_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt23_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt23_drpen_in                           : in   std_logic;
    gt23_drprdy_out                         : out  std_logic;
    gt23_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt23_eyescanreset_in                    : in   std_logic;
    gt23_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt23_eyescandataerror_out               : out  std_logic;
    gt23_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt23_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt23_rxusrclk_in                        : in   std_logic;
    gt23_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt23_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt23_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt23_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt23_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt23_rxbyteisaligned_out                : out  std_logic;
    gt23_rxmcommaalignen_in                 : in   std_logic;
    gt23_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt23_rxdfeagchold_in                    : in   std_logic;
    gt23_rxdfelfhold_in                     : in   std_logic;
    gt23_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt23_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt23_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt23_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt23_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt23_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt23_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt23_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt23_gttxreset_in                       : in   std_logic;
    gt23_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt23_txusrclk_in                        : in   std_logic;
    gt23_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt23_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt23_gthtxn_out                         : out  std_logic;
    gt23_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt23_txoutclk_out                       : out  std_logic;
    gt23_txoutclkfabric_out                 : out  std_logic;
    gt23_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt23_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt23_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt23_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT24  (X0Y24)
    --____________________________CHANNEL PORTS________________________________
 GT24_RXPMARESETDONE_OUT  : out  std_logic;
 GT24_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt24_cpllfbclklost_out                  : out  std_logic;
    gt24_cplllock_out                       : out  std_logic;
    gt24_cplllockdetclk_in                  : in   std_logic;
    gt24_cpllrefclklost_out                 : out  std_logic;
    gt24_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt24_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt24_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt24_drpclk_in                          : in   std_logic;
    gt24_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt24_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt24_drpen_in                           : in   std_logic;
    gt24_drprdy_out                         : out  std_logic;
    gt24_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt24_eyescanreset_in                    : in   std_logic;
    gt24_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt24_eyescandataerror_out               : out  std_logic;
    gt24_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt24_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt24_rxusrclk_in                        : in   std_logic;
    gt24_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt24_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt24_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt24_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt24_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt24_rxbyteisaligned_out                : out  std_logic;
    gt24_rxmcommaalignen_in                 : in   std_logic;
    gt24_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt24_rxdfeagchold_in                    : in   std_logic;
    gt24_rxdfelfhold_in                     : in   std_logic;
    gt24_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt24_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt24_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt24_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt24_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt24_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt24_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt24_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt24_gttxreset_in                       : in   std_logic;
    gt24_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt24_txusrclk_in                        : in   std_logic;
    gt24_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt24_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt24_gthtxn_out                         : out  std_logic;
    gt24_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt24_txoutclk_out                       : out  std_logic;
    gt24_txoutclkfabric_out                 : out  std_logic;
    gt24_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt24_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt24_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt24_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT25  (X0Y25)
    --____________________________CHANNEL PORTS________________________________
 GT25_RXPMARESETDONE_OUT  : out  std_logic;
 GT25_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt25_cpllfbclklost_out                  : out  std_logic;
    gt25_cplllock_out                       : out  std_logic;
    gt25_cplllockdetclk_in                  : in   std_logic;
    gt25_cpllrefclklost_out                 : out  std_logic;
    gt25_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt25_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt25_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt25_drpclk_in                          : in   std_logic;
    gt25_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt25_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt25_drpen_in                           : in   std_logic;
    gt25_drprdy_out                         : out  std_logic;
    gt25_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt25_eyescanreset_in                    : in   std_logic;
    gt25_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt25_eyescandataerror_out               : out  std_logic;
    gt25_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt25_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt25_rxusrclk_in                        : in   std_logic;
    gt25_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt25_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt25_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt25_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt25_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt25_rxbyteisaligned_out                : out  std_logic;
    gt25_rxmcommaalignen_in                 : in   std_logic;
    gt25_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt25_rxdfeagchold_in                    : in   std_logic;
    gt25_rxdfelfhold_in                     : in   std_logic;
    gt25_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt25_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt25_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt25_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt25_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt25_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt25_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt25_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt25_gttxreset_in                       : in   std_logic;
    gt25_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt25_txusrclk_in                        : in   std_logic;
    gt25_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt25_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt25_gthtxn_out                         : out  std_logic;
    gt25_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt25_txoutclk_out                       : out  std_logic;
    gt25_txoutclkfabric_out                 : out  std_logic;
    gt25_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt25_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt25_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt25_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT26  (X0Y26)
    --____________________________CHANNEL PORTS________________________________
 GT26_RXPMARESETDONE_OUT  : out  std_logic;
 GT26_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt26_cpllfbclklost_out                  : out  std_logic;
    gt26_cplllock_out                       : out  std_logic;
    gt26_cplllockdetclk_in                  : in   std_logic;
    gt26_cpllrefclklost_out                 : out  std_logic;
    gt26_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt26_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt26_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt26_drpclk_in                          : in   std_logic;
    gt26_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt26_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt26_drpen_in                           : in   std_logic;
    gt26_drprdy_out                         : out  std_logic;
    gt26_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt26_eyescanreset_in                    : in   std_logic;
    gt26_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt26_eyescandataerror_out               : out  std_logic;
    gt26_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt26_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt26_rxusrclk_in                        : in   std_logic;
    gt26_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt26_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt26_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt26_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt26_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt26_rxbyteisaligned_out                : out  std_logic;
    gt26_rxmcommaalignen_in                 : in   std_logic;
    gt26_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt26_rxdfeagchold_in                    : in   std_logic;
    gt26_rxdfelfhold_in                     : in   std_logic;
    gt26_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt26_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt26_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt26_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt26_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt26_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt26_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt26_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt26_gttxreset_in                       : in   std_logic;
    gt26_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt26_txusrclk_in                        : in   std_logic;
    gt26_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt26_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt26_gthtxn_out                         : out  std_logic;
    gt26_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt26_txoutclk_out                       : out  std_logic;
    gt26_txoutclkfabric_out                 : out  std_logic;
    gt26_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt26_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt26_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt26_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT27  (X0Y27)
    --____________________________CHANNEL PORTS________________________________
 GT27_RXPMARESETDONE_OUT  : out  std_logic;
 GT27_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt27_cpllfbclklost_out                  : out  std_logic;
    gt27_cplllock_out                       : out  std_logic;
    gt27_cplllockdetclk_in                  : in   std_logic;
    gt27_cpllrefclklost_out                 : out  std_logic;
    gt27_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt27_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt27_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt27_drpclk_in                          : in   std_logic;
    gt27_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt27_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt27_drpen_in                           : in   std_logic;
    gt27_drprdy_out                         : out  std_logic;
    gt27_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt27_eyescanreset_in                    : in   std_logic;
    gt27_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt27_eyescandataerror_out               : out  std_logic;
    gt27_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt27_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt27_rxusrclk_in                        : in   std_logic;
    gt27_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt27_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt27_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt27_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt27_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt27_rxbyteisaligned_out                : out  std_logic;
    gt27_rxmcommaalignen_in                 : in   std_logic;
    gt27_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt27_rxdfeagchold_in                    : in   std_logic;
    gt27_rxdfelfhold_in                     : in   std_logic;
    gt27_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt27_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt27_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt27_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt27_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt27_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt27_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt27_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt27_gttxreset_in                       : in   std_logic;
    gt27_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt27_txusrclk_in                        : in   std_logic;
    gt27_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt27_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt27_gthtxn_out                         : out  std_logic;
    gt27_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt27_txoutclk_out                       : out  std_logic;
    gt27_txoutclkfabric_out                 : out  std_logic;
    gt27_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt27_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt27_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt27_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT28  (X0Y28)
    --____________________________CHANNEL PORTS________________________________
 GT28_RXPMARESETDONE_OUT  : out  std_logic;
 GT28_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt28_cpllfbclklost_out                  : out  std_logic;
    gt28_cplllock_out                       : out  std_logic;
    gt28_cplllockdetclk_in                  : in   std_logic;
    gt28_cpllrefclklost_out                 : out  std_logic;
    gt28_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt28_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt28_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt28_drpclk_in                          : in   std_logic;
    gt28_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt28_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt28_drpen_in                           : in   std_logic;
    gt28_drprdy_out                         : out  std_logic;
    gt28_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt28_eyescanreset_in                    : in   std_logic;
    gt28_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt28_eyescandataerror_out               : out  std_logic;
    gt28_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt28_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt28_rxusrclk_in                        : in   std_logic;
    gt28_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt28_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt28_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt28_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt28_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt28_rxbyteisaligned_out                : out  std_logic;
    gt28_rxmcommaalignen_in                 : in   std_logic;
    gt28_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt28_rxdfeagchold_in                    : in   std_logic;
    gt28_rxdfelfhold_in                     : in   std_logic;
    gt28_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt28_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt28_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt28_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt28_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt28_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt28_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt28_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt28_gttxreset_in                       : in   std_logic;
    gt28_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt28_txusrclk_in                        : in   std_logic;
    gt28_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt28_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt28_gthtxn_out                         : out  std_logic;
    gt28_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt28_txoutclk_out                       : out  std_logic;
    gt28_txoutclkfabric_out                 : out  std_logic;
    gt28_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt28_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt28_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt28_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT29  (X0Y29)
    --____________________________CHANNEL PORTS________________________________
 GT29_RXPMARESETDONE_OUT  : out  std_logic;
 GT29_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt29_cpllfbclklost_out                  : out  std_logic;
    gt29_cplllock_out                       : out  std_logic;
    gt29_cplllockdetclk_in                  : in   std_logic;
    gt29_cpllrefclklost_out                 : out  std_logic;
    gt29_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt29_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt29_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt29_drpclk_in                          : in   std_logic;
    gt29_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt29_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt29_drpen_in                           : in   std_logic;
    gt29_drprdy_out                         : out  std_logic;
    gt29_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt29_eyescanreset_in                    : in   std_logic;
    gt29_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt29_eyescandataerror_out               : out  std_logic;
    gt29_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt29_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt29_rxusrclk_in                        : in   std_logic;
    gt29_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt29_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt29_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt29_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt29_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt29_rxbyteisaligned_out                : out  std_logic;
    gt29_rxmcommaalignen_in                 : in   std_logic;
    gt29_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt29_rxdfeagchold_in                    : in   std_logic;
    gt29_rxdfelfhold_in                     : in   std_logic;
    gt29_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt29_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt29_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt29_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt29_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt29_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt29_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt29_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt29_gttxreset_in                       : in   std_logic;
    gt29_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt29_txusrclk_in                        : in   std_logic;
    gt29_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt29_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt29_gthtxn_out                         : out  std_logic;
    gt29_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt29_txoutclk_out                       : out  std_logic;
    gt29_txoutclkfabric_out                 : out  std_logic;
    gt29_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt29_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt29_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt29_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT30  (X0Y30)
    --____________________________CHANNEL PORTS________________________________
 GT30_RXPMARESETDONE_OUT  : out  std_logic;
 GT30_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt30_cpllfbclklost_out                  : out  std_logic;
    gt30_cplllock_out                       : out  std_logic;
    gt30_cplllockdetclk_in                  : in   std_logic;
    gt30_cpllrefclklost_out                 : out  std_logic;
    gt30_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt30_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt30_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt30_drpclk_in                          : in   std_logic;
    gt30_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt30_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt30_drpen_in                           : in   std_logic;
    gt30_drprdy_out                         : out  std_logic;
    gt30_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt30_eyescanreset_in                    : in   std_logic;
    gt30_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt30_eyescandataerror_out               : out  std_logic;
    gt30_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt30_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt30_rxusrclk_in                        : in   std_logic;
    gt30_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt30_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt30_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt30_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt30_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt30_rxbyteisaligned_out                : out  std_logic;
    gt30_rxmcommaalignen_in                 : in   std_logic;
    gt30_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt30_rxdfeagchold_in                    : in   std_logic;
    gt30_rxdfelfhold_in                     : in   std_logic;
    gt30_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt30_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt30_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt30_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt30_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt30_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt30_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt30_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt30_gttxreset_in                       : in   std_logic;
    gt30_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt30_txusrclk_in                        : in   std_logic;
    gt30_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt30_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt30_gthtxn_out                         : out  std_logic;
    gt30_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt30_txoutclk_out                       : out  std_logic;
    gt30_txoutclkfabric_out                 : out  std_logic;
    gt30_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt30_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt30_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt30_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT31  (X0Y31)
    --____________________________CHANNEL PORTS________________________________
 GT31_RXPMARESETDONE_OUT  : out  std_logic;
 GT31_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt31_cpllfbclklost_out                  : out  std_logic;
    gt31_cplllock_out                       : out  std_logic;
    gt31_cplllockdetclk_in                  : in   std_logic;
    gt31_cpllrefclklost_out                 : out  std_logic;
    gt31_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt31_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt31_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt31_drpclk_in                          : in   std_logic;
    gt31_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt31_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt31_drpen_in                           : in   std_logic;
    gt31_drprdy_out                         : out  std_logic;
    gt31_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt31_eyescanreset_in                    : in   std_logic;
    gt31_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt31_eyescandataerror_out               : out  std_logic;
    gt31_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt31_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt31_rxusrclk_in                        : in   std_logic;
    gt31_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt31_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt31_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt31_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt31_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt31_rxbyteisaligned_out                : out  std_logic;
    gt31_rxmcommaalignen_in                 : in   std_logic;
    gt31_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt31_rxdfeagchold_in                    : in   std_logic;
    gt31_rxdfelfhold_in                     : in   std_logic;
    gt31_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt31_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt31_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt31_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt31_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt31_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt31_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt31_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt31_gttxreset_in                       : in   std_logic;
    gt31_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt31_txusrclk_in                        : in   std_logic;
    gt31_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt31_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt31_gthtxn_out                         : out  std_logic;
    gt31_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt31_txoutclk_out                       : out  std_logic;
    gt31_txoutclkfabric_out                 : out  std_logic;
    gt31_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt31_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt31_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt31_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT32  (X0Y32)
    --____________________________CHANNEL PORTS________________________________
 GT32_RXPMARESETDONE_OUT  : out  std_logic;
 GT32_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt32_cpllfbclklost_out                  : out  std_logic;
    gt32_cplllock_out                       : out  std_logic;
    gt32_cplllockdetclk_in                  : in   std_logic;
    gt32_cpllrefclklost_out                 : out  std_logic;
    gt32_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt32_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt32_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt32_drpclk_in                          : in   std_logic;
    gt32_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt32_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt32_drpen_in                           : in   std_logic;
    gt32_drprdy_out                         : out  std_logic;
    gt32_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt32_eyescanreset_in                    : in   std_logic;
    gt32_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt32_eyescandataerror_out               : out  std_logic;
    gt32_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt32_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt32_rxusrclk_in                        : in   std_logic;
    gt32_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt32_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt32_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt32_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt32_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt32_rxbyteisaligned_out                : out  std_logic;
    gt32_rxmcommaalignen_in                 : in   std_logic;
    gt32_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt32_rxdfeagchold_in                    : in   std_logic;
    gt32_rxdfelfhold_in                     : in   std_logic;
    gt32_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt32_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt32_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt32_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt32_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt32_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt32_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt32_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt32_gttxreset_in                       : in   std_logic;
    gt32_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt32_txusrclk_in                        : in   std_logic;
    gt32_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt32_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt32_gthtxn_out                         : out  std_logic;
    gt32_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt32_txoutclk_out                       : out  std_logic;
    gt32_txoutclkfabric_out                 : out  std_logic;
    gt32_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt32_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt32_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt32_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT33  (X0Y33)
    --____________________________CHANNEL PORTS________________________________
 GT33_RXPMARESETDONE_OUT  : out  std_logic;
 GT33_TXPMARESETDONE_OUT  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    gt33_cpllfbclklost_out                  : out  std_logic;
    gt33_cplllock_out                       : out  std_logic;
    gt33_cplllockdetclk_in                  : in   std_logic;
    gt33_cpllrefclklost_out                 : out  std_logic;
    gt33_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt33_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt33_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt33_drpclk_in                          : in   std_logic;
    gt33_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt33_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt33_drpen_in                           : in   std_logic;
    gt33_drprdy_out                         : out  std_logic;
    gt33_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt33_eyescanreset_in                    : in   std_logic;
    gt33_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt33_eyescandataerror_out               : out  std_logic;
    gt33_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt33_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt33_rxusrclk_in                        : in   std_logic;
    gt33_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt33_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt33_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt33_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt33_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt33_rxbyteisaligned_out                : out  std_logic;
    gt33_rxmcommaalignen_in                 : in   std_logic;
    gt33_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt33_rxdfeagchold_in                    : in   std_logic;
    gt33_rxdfelfhold_in                     : in   std_logic;
    gt33_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt33_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt33_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt33_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt33_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt33_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt33_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt33_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt33_gttxreset_in                       : in   std_logic;
    gt33_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt33_txusrclk_in                        : in   std_logic;
    gt33_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt33_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt33_gthtxn_out                         : out  std_logic;
    gt33_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt33_txoutclk_out                       : out  std_logic;
    gt33_txoutclkfabric_out                 : out  std_logic;
    gt33_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt33_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt33_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt33_txcharisk_in                       : in   std_logic_vector(3 downto 0);


    --____________________________COMMON PORTS________________________________
     GT0_QPLLOUTCLK_IN : in std_logic;
     GT0_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT1_QPLLOUTCLK_IN : in std_logic;
     GT1_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT2_QPLLOUTCLK_IN : in std_logic;
     GT2_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT3_QPLLOUTCLK_IN : in std_logic;
     GT3_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT4_QPLLOUTCLK_IN : in std_logic;
     GT4_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT5_QPLLOUTCLK_IN : in std_logic;
     GT5_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT6_QPLLOUTCLK_IN : in std_logic;
     GT6_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT7_QPLLOUTCLK_IN : in std_logic;
     GT7_QPLLOUTREFCLK_IN  : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT8_QPLLOUTCLK_IN : in std_logic;
     GT8_QPLLOUTREFCLK_IN  : in std_logic

);


end gt6_rtm34l_multi_gt;
    
architecture RTL of gt6_rtm34l_multi_gt is
    attribute DowngradeIPIdentifiedWarnings: string;
    attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

    attribute CORE_GENERATION_INFO : string;
    attribute CORE_GENERATION_INFO of RTL : architecture is "gt6_rtm34l_multi_gt,gtwizard_v3_2,{protocol_file=Start_from_scratch}";


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--***************************** Signal Declarations *****************************

    -- ground and tied_to_vcc_i signals
signal  tied_to_ground_i                :   std_logic;
signal  tied_to_ground_vec_i            :   std_logic_vector(63 downto 0);
signal  tied_to_vcc_i                   :   std_logic;
signal   gt0_qplloutclk_i         :   std_logic;
signal   gt0_qplloutrefclk_i      :   std_logic;
signal   gt1_qplloutclk_i         :   std_logic;
signal   gt1_qplloutrefclk_i      :   std_logic;
signal   gt2_qplloutclk_i         :   std_logic;
signal   gt2_qplloutrefclk_i      :   std_logic;
signal   gt3_qplloutclk_i         :   std_logic;
signal   gt3_qplloutrefclk_i      :   std_logic;
signal   gt4_qplloutclk_i         :   std_logic;
signal   gt4_qplloutrefclk_i      :   std_logic;
signal   gt5_qplloutclk_i         :   std_logic;
signal   gt5_qplloutrefclk_i      :   std_logic;
signal   gt6_qplloutclk_i         :   std_logic;
signal   gt6_qplloutrefclk_i      :   std_logic;
signal   gt7_qplloutclk_i         :   std_logic;
signal   gt7_qplloutrefclk_i      :   std_logic;
signal   gt8_qplloutclk_i         :   std_logic;
signal   gt8_qplloutrefclk_i      :   std_logic;

signal  gt0_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt0_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt1_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt1_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt2_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt2_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt3_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt3_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt4_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt4_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt5_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt5_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt6_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt6_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt7_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt7_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt8_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt8_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt9_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt9_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt10_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt10_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt11_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt11_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt12_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt12_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt13_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt13_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt14_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt14_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt15_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt15_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt16_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt16_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt17_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt17_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt18_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt18_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt19_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt19_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt20_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt20_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt21_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt21_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt22_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt22_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt23_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt23_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt24_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt24_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt25_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt25_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt26_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt26_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt27_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt27_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt28_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt28_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt29_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt29_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt30_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt30_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt31_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt31_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt32_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt32_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
signal  gt33_mgtrefclktx_i           :   std_logic_vector(1 downto 0);
signal  gt33_mgtrefclkrx_i           :   std_logic_vector(1 downto 0);
 

signal   gt0_qpllclk_i            :   std_logic;
signal   gt0_qpllrefclk_i         :   std_logic;
signal   gt1_qpllclk_i            :   std_logic;
signal   gt1_qpllrefclk_i         :   std_logic;
signal   gt2_qpllclk_i            :   std_logic;
signal   gt2_qpllrefclk_i         :   std_logic;
signal   gt3_qpllclk_i            :   std_logic;
signal   gt3_qpllrefclk_i         :   std_logic;
signal   gt4_qpllclk_i            :   std_logic;
signal   gt4_qpllrefclk_i         :   std_logic;
signal   gt5_qpllclk_i            :   std_logic;
signal   gt5_qpllrefclk_i         :   std_logic;
signal   gt6_qpllclk_i            :   std_logic;
signal   gt6_qpllrefclk_i         :   std_logic;
signal   gt7_qpllclk_i            :   std_logic;
signal   gt7_qpllrefclk_i         :   std_logic;
signal   gt8_qpllclk_i            :   std_logic;
signal   gt8_qpllrefclk_i         :   std_logic;
signal   gt9_qpllclk_i            :   std_logic;
signal   gt9_qpllrefclk_i         :   std_logic;
signal   gt10_qpllclk_i            :   std_logic;
signal   gt10_qpllrefclk_i         :   std_logic;
signal   gt11_qpllclk_i            :   std_logic;
signal   gt11_qpllrefclk_i         :   std_logic;
signal   gt12_qpllclk_i            :   std_logic;
signal   gt12_qpllrefclk_i         :   std_logic;
signal   gt13_qpllclk_i            :   std_logic;
signal   gt13_qpllrefclk_i         :   std_logic;
signal   gt14_qpllclk_i            :   std_logic;
signal   gt14_qpllrefclk_i         :   std_logic;
signal   gt15_qpllclk_i            :   std_logic;
signal   gt15_qpllrefclk_i         :   std_logic;
signal   gt16_qpllclk_i            :   std_logic;
signal   gt16_qpllrefclk_i         :   std_logic;
signal   gt17_qpllclk_i            :   std_logic;
signal   gt17_qpllrefclk_i         :   std_logic;
signal   gt18_qpllclk_i            :   std_logic;
signal   gt18_qpllrefclk_i         :   std_logic;
signal   gt19_qpllclk_i            :   std_logic;
signal   gt19_qpllrefclk_i         :   std_logic;
signal   gt20_qpllclk_i            :   std_logic;
signal   gt20_qpllrefclk_i         :   std_logic;
signal   gt21_qpllclk_i            :   std_logic;
signal   gt21_qpllrefclk_i         :   std_logic;
signal   gt22_qpllclk_i            :   std_logic;
signal   gt22_qpllrefclk_i         :   std_logic;
signal   gt23_qpllclk_i            :   std_logic;
signal   gt23_qpllrefclk_i         :   std_logic;
signal   gt24_qpllclk_i            :   std_logic;
signal   gt24_qpllrefclk_i         :   std_logic;
signal   gt25_qpllclk_i            :   std_logic;
signal   gt25_qpllrefclk_i         :   std_logic;
signal   gt26_qpllclk_i            :   std_logic;
signal   gt26_qpllrefclk_i         :   std_logic;
signal   gt27_qpllclk_i            :   std_logic;
signal   gt27_qpllrefclk_i         :   std_logic;
signal   gt28_qpllclk_i            :   std_logic;
signal   gt28_qpllrefclk_i         :   std_logic;
signal   gt29_qpllclk_i            :   std_logic;
signal   gt29_qpllrefclk_i         :   std_logic;
signal   gt30_qpllclk_i            :   std_logic;
signal   gt30_qpllrefclk_i         :   std_logic;
signal   gt31_qpllclk_i            :   std_logic;
signal   gt31_qpllrefclk_i         :   std_logic;
signal   gt32_qpllclk_i            :   std_logic;
signal   gt32_qpllrefclk_i         :   std_logic;
signal   gt33_qpllclk_i            :   std_logic;
signal   gt33_qpllrefclk_i         :   std_logic;


--*************************** Component Declarations **************************
component gt6_rtm34l_GT
generic
(
    -- Simulation attributes
    GT_SIM_GTRESET_SPEEDUP    : string := "FALSE";
    EXAMPLE_SIMULATION        : integer  := 0;   
    TXSYNC_OVRD_IN            : bit    := '0';
    TXSYNC_MULTILANE_IN       : bit    := '0'     
);
port 
(   
 RXPMARESETDONE  : out  std_logic;
 TXPMARESETDONE  : out  std_logic;
    --------------------------------- CPLL Ports -------------------------------
    cpllfbclklost_out                       : out  std_logic;
    cplllock_out                            : out  std_logic;
    cplllockdetclk_in                       : in   std_logic;
    cpllrefclklost_out                      : out  std_logic;
    cpllreset_in                            : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gtrefclk0_in                            : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    drpaddr_in                              : in   std_logic_vector(8 downto 0);
    drpclk_in                               : in   std_logic;
    drpdi_in                                : in   std_logic_vector(15 downto 0);
    drpdo_out                               : out  std_logic_vector(15 downto 0);
    drpen_in                                : in   std_logic;
    drprdy_out                              : out  std_logic;
    drpwe_in                                : in   std_logic;
    ------------------------------- Clocking Ports -----------------------------
    qpllclk_in                              : in   std_logic;
    qpllrefclk_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    eyescanreset_in                         : in   std_logic;
    rxuserrdy_in                            : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    eyescandataerror_out                    : out  std_logic;
    eyescantrigger_in                       : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    dmonitorout_out                         : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    rxusrclk_in                             : in   std_logic;
    rxusrclk2_in                            : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    rxdata_out                              : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    rxdisperr_out                           : out  std_logic_vector(3 downto 0);
    rxnotintable_out                        : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gthrxn_in                               : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    rxbyteisaligned_out                     : out  std_logic;
    rxmcommaalignen_in                      : in   std_logic;
    rxpcommaalignen_in                      : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    rxdfeagchold_in                         : in   std_logic;
    rxdfelfhold_in                          : in   std_logic;
    rxmonitorout_out                        : out  std_logic_vector(6 downto 0);
    rxmonitorsel_in                         : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    rxoutclk_out                            : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gtrxreset_in                            : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    rxpolarity_in                           : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    rxcharisk_out                           : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gthrxp_in                               : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    rxresetdone_out                         : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gttxreset_in                            : in   std_logic;
    txuserrdy_in                            : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    txusrclk_in                             : in   std_logic;
    txusrclk2_in                            : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    txdata_in                               : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gthtxn_out                              : out  std_logic;
    gthtxp_out                              : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    txoutclk_out                            : out  std_logic;
    txoutclkfabric_out                      : out  std_logic;
    txoutclkpcs_out                         : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    txresetdone_out                         : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    txpolarity_in                           : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    txcharisk_in                            : in   std_logic_vector(3 downto 0)


);
end component;


--********************************* Main Body of Code**************************

begin                       

    tied_to_ground_i                    <= '0';
    tied_to_ground_vec_i(63 downto 0)   <= (others => '0');
    tied_to_vcc_i                       <= '1';
    gt0_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt0_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 
    gt1_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt1_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 
    gt2_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt2_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 
    gt3_qpllclk_i    <= GT0_QPLLOUTCLK_IN;  
    gt3_qpllrefclk_i <= GT0_QPLLOUTREFCLK_IN; 
    gt4_qpllclk_i    <= GT1_QPLLOUTCLK_IN;  
    gt4_qpllrefclk_i <= GT1_QPLLOUTREFCLK_IN; 
    gt5_qpllclk_i    <= GT1_QPLLOUTCLK_IN;  
    gt5_qpllrefclk_i <= GT1_QPLLOUTREFCLK_IN; 
    gt6_qpllclk_i    <= GT1_QPLLOUTCLK_IN;  
    gt6_qpllrefclk_i <= GT1_QPLLOUTREFCLK_IN; 
    gt7_qpllclk_i    <= GT1_QPLLOUTCLK_IN;  
    gt7_qpllrefclk_i <= GT1_QPLLOUTREFCLK_IN; 
    gt8_qpllclk_i    <= GT2_QPLLOUTCLK_IN;  
    gt8_qpllrefclk_i <= GT2_QPLLOUTREFCLK_IN; 
    gt9_qpllclk_i    <= GT2_QPLLOUTCLK_IN;  
    gt9_qpllrefclk_i <= GT2_QPLLOUTREFCLK_IN; 
    gt10_qpllclk_i    <= GT2_QPLLOUTCLK_IN;  
    gt10_qpllrefclk_i <= GT2_QPLLOUTREFCLK_IN; 
    gt11_qpllclk_i    <= GT2_QPLLOUTCLK_IN;  
    gt11_qpllrefclk_i <= GT2_QPLLOUTREFCLK_IN; 
    gt12_qpllclk_i    <= GT3_QPLLOUTCLK_IN;  
    gt12_qpllrefclk_i <= GT3_QPLLOUTREFCLK_IN; 
    gt13_qpllclk_i    <= GT3_QPLLOUTCLK_IN;  
    gt13_qpllrefclk_i <= GT3_QPLLOUTREFCLK_IN; 
    gt14_qpllclk_i    <= GT3_QPLLOUTCLK_IN;  
    gt14_qpllrefclk_i <= GT3_QPLLOUTREFCLK_IN; 
    gt15_qpllclk_i    <= GT3_QPLLOUTCLK_IN;  
    gt15_qpllrefclk_i <= GT3_QPLLOUTREFCLK_IN; 
    gt16_qpllclk_i    <= GT4_QPLLOUTCLK_IN;  
    gt16_qpllrefclk_i <= GT4_QPLLOUTREFCLK_IN; 
    gt17_qpllclk_i    <= GT4_QPLLOUTCLK_IN;  
    gt17_qpllrefclk_i <= GT4_QPLLOUTREFCLK_IN; 
    gt18_qpllclk_i    <= GT4_QPLLOUTCLK_IN;  
    gt18_qpllrefclk_i <= GT4_QPLLOUTREFCLK_IN; 
    gt19_qpllclk_i    <= GT4_QPLLOUTCLK_IN;  
    gt19_qpllrefclk_i <= GT4_QPLLOUTREFCLK_IN; 
    gt20_qpllclk_i    <= GT5_QPLLOUTCLK_IN;  
    gt20_qpllrefclk_i <= GT5_QPLLOUTREFCLK_IN; 
    gt21_qpllclk_i    <= GT5_QPLLOUTCLK_IN;  
    gt21_qpllrefclk_i <= GT5_QPLLOUTREFCLK_IN; 
    gt22_qpllclk_i    <= GT5_QPLLOUTCLK_IN;  
    gt22_qpllrefclk_i <= GT5_QPLLOUTREFCLK_IN; 
    gt23_qpllclk_i    <= GT5_QPLLOUTCLK_IN;  
    gt23_qpllrefclk_i <= GT5_QPLLOUTREFCLK_IN; 
    gt24_qpllclk_i    <= GT6_QPLLOUTCLK_IN;  
    gt24_qpllrefclk_i <= GT6_QPLLOUTREFCLK_IN; 
    gt25_qpllclk_i    <= GT6_QPLLOUTCLK_IN;  
    gt25_qpllrefclk_i <= GT6_QPLLOUTREFCLK_IN; 
    gt26_qpllclk_i    <= GT6_QPLLOUTCLK_IN;  
    gt26_qpllrefclk_i <= GT6_QPLLOUTREFCLK_IN; 
    gt27_qpllclk_i    <= GT6_QPLLOUTCLK_IN;  
    gt27_qpllrefclk_i <= GT6_QPLLOUTREFCLK_IN; 
    gt28_qpllclk_i    <= GT7_QPLLOUTCLK_IN;  
    gt28_qpllrefclk_i <= GT7_QPLLOUTREFCLK_IN; 
    gt29_qpllclk_i    <= GT7_QPLLOUTCLK_IN;  
    gt29_qpllrefclk_i <= GT7_QPLLOUTREFCLK_IN; 
    gt30_qpllclk_i    <= GT7_QPLLOUTCLK_IN;  
    gt30_qpllrefclk_i <= GT7_QPLLOUTREFCLK_IN; 
    gt31_qpllclk_i    <= GT7_QPLLOUTCLK_IN;  
    gt31_qpllrefclk_i <= GT7_QPLLOUTREFCLK_IN; 
    gt32_qpllclk_i    <= GT8_QPLLOUTCLK_IN;  
    gt32_qpllrefclk_i <= GT8_QPLLOUTREFCLK_IN; 
    gt33_qpllclk_i    <= GT8_QPLLOUTCLK_IN;  
    gt33_qpllrefclk_i <= GT8_QPLLOUTREFCLK_IN; 


    --------------------------- GT Instances  -------------------------------   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X0Y0)
gt0_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT0_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT0_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt0_cpllfbclklost_out,
        cplllock_out                    =>      gt0_cplllock_out,
        cplllockdetclk_in               =>      gt0_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt0_cpllrefclklost_out,
        cpllreset_in                    =>      gt0_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt0_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt0_drpaddr_in,
        drpclk_in                       =>      gt0_drpclk_in,
        drpdi_in                        =>      gt0_drpdi_in,
        drpdo_out                       =>      gt0_drpdo_out,
        drpen_in                        =>      gt0_drpen_in,
        drprdy_out                      =>      gt0_drprdy_out,
        drpwe_in                        =>      gt0_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt0_qpllclk_i,
        qpllrefclk_in                   =>      gt0_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt0_eyescanreset_in,
        rxuserrdy_in                    =>      gt0_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt0_eyescandataerror_out,
        eyescantrigger_in               =>      gt0_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt0_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt0_rxusrclk_in,
        rxusrclk2_in                    =>      gt0_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt0_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt0_rxdisperr_out,
        rxnotintable_out                =>      gt0_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt0_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt0_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt0_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt0_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt0_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt0_rxdfelfhold_in,
        rxmonitorout_out                =>      gt0_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt0_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt0_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt0_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt0_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt0_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt0_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt0_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt0_gttxreset_in,
        txuserrdy_in                    =>      gt0_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt0_txusrclk_in,
        txusrclk2_in                    =>      gt0_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt0_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt0_gthtxn_out,
        gthtxp_out                      =>      gt0_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt0_txoutclk_out,
        txoutclkfabric_out              =>      gt0_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt0_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt0_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt0_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt0_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT1  (X0Y1)
gt1_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT1_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT1_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt1_cpllfbclklost_out,
        cplllock_out                    =>      gt1_cplllock_out,
        cplllockdetclk_in               =>      gt1_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt1_cpllrefclklost_out,
        cpllreset_in                    =>      gt1_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt1_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt1_drpaddr_in,
        drpclk_in                       =>      gt1_drpclk_in,
        drpdi_in                        =>      gt1_drpdi_in,
        drpdo_out                       =>      gt1_drpdo_out,
        drpen_in                        =>      gt1_drpen_in,
        drprdy_out                      =>      gt1_drprdy_out,
        drpwe_in                        =>      gt1_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt1_qpllclk_i,
        qpllrefclk_in                   =>      gt1_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt1_eyescanreset_in,
        rxuserrdy_in                    =>      gt1_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt1_eyescandataerror_out,
        eyescantrigger_in               =>      gt1_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt1_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt1_rxusrclk_in,
        rxusrclk2_in                    =>      gt1_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt1_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt1_rxdisperr_out,
        rxnotintable_out                =>      gt1_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt1_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt1_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt1_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt1_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt1_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt1_rxdfelfhold_in,
        rxmonitorout_out                =>      gt1_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt1_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt1_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt1_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt1_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt1_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt1_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt1_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt1_gttxreset_in,
        txuserrdy_in                    =>      gt1_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt1_txusrclk_in,
        txusrclk2_in                    =>      gt1_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt1_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt1_gthtxn_out,
        gthtxp_out                      =>      gt1_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt1_txoutclk_out,
        txoutclkfabric_out              =>      gt1_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt1_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt1_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt1_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt1_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT2  (X0Y2)
gt2_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT2_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT2_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt2_cpllfbclklost_out,
        cplllock_out                    =>      gt2_cplllock_out,
        cplllockdetclk_in               =>      gt2_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt2_cpllrefclklost_out,
        cpllreset_in                    =>      gt2_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt2_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt2_drpaddr_in,
        drpclk_in                       =>      gt2_drpclk_in,
        drpdi_in                        =>      gt2_drpdi_in,
        drpdo_out                       =>      gt2_drpdo_out,
        drpen_in                        =>      gt2_drpen_in,
        drprdy_out                      =>      gt2_drprdy_out,
        drpwe_in                        =>      gt2_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt2_qpllclk_i,
        qpllrefclk_in                   =>      gt2_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt2_eyescanreset_in,
        rxuserrdy_in                    =>      gt2_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt2_eyescandataerror_out,
        eyescantrigger_in               =>      gt2_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt2_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt2_rxusrclk_in,
        rxusrclk2_in                    =>      gt2_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt2_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt2_rxdisperr_out,
        rxnotintable_out                =>      gt2_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt2_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt2_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt2_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt2_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt2_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt2_rxdfelfhold_in,
        rxmonitorout_out                =>      gt2_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt2_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt2_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt2_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt2_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt2_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt2_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt2_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt2_gttxreset_in,
        txuserrdy_in                    =>      gt2_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt2_txusrclk_in,
        txusrclk2_in                    =>      gt2_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt2_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt2_gthtxn_out,
        gthtxp_out                      =>      gt2_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt2_txoutclk_out,
        txoutclkfabric_out              =>      gt2_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt2_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt2_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt2_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt2_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT3  (X0Y3)
gt3_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT3_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT3_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt3_cpllfbclklost_out,
        cplllock_out                    =>      gt3_cplllock_out,
        cplllockdetclk_in               =>      gt3_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt3_cpllrefclklost_out,
        cpllreset_in                    =>      gt3_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt3_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt3_drpaddr_in,
        drpclk_in                       =>      gt3_drpclk_in,
        drpdi_in                        =>      gt3_drpdi_in,
        drpdo_out                       =>      gt3_drpdo_out,
        drpen_in                        =>      gt3_drpen_in,
        drprdy_out                      =>      gt3_drprdy_out,
        drpwe_in                        =>      gt3_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt3_qpllclk_i,
        qpllrefclk_in                   =>      gt3_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt3_eyescanreset_in,
        rxuserrdy_in                    =>      gt3_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt3_eyescandataerror_out,
        eyescantrigger_in               =>      gt3_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt3_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt3_rxusrclk_in,
        rxusrclk2_in                    =>      gt3_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt3_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt3_rxdisperr_out,
        rxnotintable_out                =>      gt3_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt3_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt3_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt3_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt3_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt3_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt3_rxdfelfhold_in,
        rxmonitorout_out                =>      gt3_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt3_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt3_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt3_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt3_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt3_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt3_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt3_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt3_gttxreset_in,
        txuserrdy_in                    =>      gt3_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt3_txusrclk_in,
        txusrclk2_in                    =>      gt3_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt3_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt3_gthtxn_out,
        gthtxp_out                      =>      gt3_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt3_txoutclk_out,
        txoutclkfabric_out              =>      gt3_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt3_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt3_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt3_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt3_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT4  (X0Y4)
gt4_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT4_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT4_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt4_cpllfbclklost_out,
        cplllock_out                    =>      gt4_cplllock_out,
        cplllockdetclk_in               =>      gt4_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt4_cpllrefclklost_out,
        cpllreset_in                    =>      gt4_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt4_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt4_drpaddr_in,
        drpclk_in                       =>      gt4_drpclk_in,
        drpdi_in                        =>      gt4_drpdi_in,
        drpdo_out                       =>      gt4_drpdo_out,
        drpen_in                        =>      gt4_drpen_in,
        drprdy_out                      =>      gt4_drprdy_out,
        drpwe_in                        =>      gt4_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt4_qpllclk_i,
        qpllrefclk_in                   =>      gt4_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt4_eyescanreset_in,
        rxuserrdy_in                    =>      gt4_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt4_eyescandataerror_out,
        eyescantrigger_in               =>      gt4_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt4_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt4_rxusrclk_in,
        rxusrclk2_in                    =>      gt4_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt4_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt4_rxdisperr_out,
        rxnotintable_out                =>      gt4_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt4_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt4_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt4_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt4_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt4_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt4_rxdfelfhold_in,
        rxmonitorout_out                =>      gt4_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt4_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt4_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt4_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt4_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt4_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt4_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt4_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt4_gttxreset_in,
        txuserrdy_in                    =>      gt4_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt4_txusrclk_in,
        txusrclk2_in                    =>      gt4_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt4_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt4_gthtxn_out,
        gthtxp_out                      =>      gt4_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt4_txoutclk_out,
        txoutclkfabric_out              =>      gt4_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt4_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt4_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt4_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt4_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT5  (X0Y5)
gt5_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT5_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT5_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt5_cpllfbclklost_out,
        cplllock_out                    =>      gt5_cplllock_out,
        cplllockdetclk_in               =>      gt5_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt5_cpllrefclklost_out,
        cpllreset_in                    =>      gt5_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt5_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt5_drpaddr_in,
        drpclk_in                       =>      gt5_drpclk_in,
        drpdi_in                        =>      gt5_drpdi_in,
        drpdo_out                       =>      gt5_drpdo_out,
        drpen_in                        =>      gt5_drpen_in,
        drprdy_out                      =>      gt5_drprdy_out,
        drpwe_in                        =>      gt5_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt5_qpllclk_i,
        qpllrefclk_in                   =>      gt5_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt5_eyescanreset_in,
        rxuserrdy_in                    =>      gt5_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt5_eyescandataerror_out,
        eyescantrigger_in               =>      gt5_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt5_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt5_rxusrclk_in,
        rxusrclk2_in                    =>      gt5_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt5_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt5_rxdisperr_out,
        rxnotintable_out                =>      gt5_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt5_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt5_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt5_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt5_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt5_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt5_rxdfelfhold_in,
        rxmonitorout_out                =>      gt5_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt5_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt5_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt5_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt5_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt5_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt5_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt5_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt5_gttxreset_in,
        txuserrdy_in                    =>      gt5_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt5_txusrclk_in,
        txusrclk2_in                    =>      gt5_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt5_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt5_gthtxn_out,
        gthtxp_out                      =>      gt5_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt5_txoutclk_out,
        txoutclkfabric_out              =>      gt5_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt5_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt5_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt5_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt5_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT6  (X0Y6)
gt6_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT6_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT6_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt6_cpllfbclklost_out,
        cplllock_out                    =>      gt6_cplllock_out,
        cplllockdetclk_in               =>      gt6_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt6_cpllrefclklost_out,
        cpllreset_in                    =>      gt6_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt6_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt6_drpaddr_in,
        drpclk_in                       =>      gt6_drpclk_in,
        drpdi_in                        =>      gt6_drpdi_in,
        drpdo_out                       =>      gt6_drpdo_out,
        drpen_in                        =>      gt6_drpen_in,
        drprdy_out                      =>      gt6_drprdy_out,
        drpwe_in                        =>      gt6_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt6_qpllclk_i,
        qpllrefclk_in                   =>      gt6_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt6_eyescanreset_in,
        rxuserrdy_in                    =>      gt6_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt6_eyescandataerror_out,
        eyescantrigger_in               =>      gt6_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt6_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt6_rxusrclk_in,
        rxusrclk2_in                    =>      gt6_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt6_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt6_rxdisperr_out,
        rxnotintable_out                =>      gt6_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt6_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt6_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt6_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt6_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt6_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt6_rxdfelfhold_in,
        rxmonitorout_out                =>      gt6_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt6_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt6_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt6_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt6_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt6_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt6_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt6_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt6_gttxreset_in,
        txuserrdy_in                    =>      gt6_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt6_txusrclk_in,
        txusrclk2_in                    =>      gt6_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt6_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt6_gthtxn_out,
        gthtxp_out                      =>      gt6_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt6_txoutclk_out,
        txoutclkfabric_out              =>      gt6_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt6_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt6_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt6_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt6_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT7  (X0Y7)
gt7_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT7_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT7_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt7_cpllfbclklost_out,
        cplllock_out                    =>      gt7_cplllock_out,
        cplllockdetclk_in               =>      gt7_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt7_cpllrefclklost_out,
        cpllreset_in                    =>      gt7_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt7_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt7_drpaddr_in,
        drpclk_in                       =>      gt7_drpclk_in,
        drpdi_in                        =>      gt7_drpdi_in,
        drpdo_out                       =>      gt7_drpdo_out,
        drpen_in                        =>      gt7_drpen_in,
        drprdy_out                      =>      gt7_drprdy_out,
        drpwe_in                        =>      gt7_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt7_qpllclk_i,
        qpllrefclk_in                   =>      gt7_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt7_eyescanreset_in,
        rxuserrdy_in                    =>      gt7_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt7_eyescandataerror_out,
        eyescantrigger_in               =>      gt7_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt7_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt7_rxusrclk_in,
        rxusrclk2_in                    =>      gt7_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt7_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt7_rxdisperr_out,
        rxnotintable_out                =>      gt7_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt7_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt7_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt7_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt7_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt7_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt7_rxdfelfhold_in,
        rxmonitorout_out                =>      gt7_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt7_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt7_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt7_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt7_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt7_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt7_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt7_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt7_gttxreset_in,
        txuserrdy_in                    =>      gt7_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt7_txusrclk_in,
        txusrclk2_in                    =>      gt7_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt7_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt7_gthtxn_out,
        gthtxp_out                      =>      gt7_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt7_txoutclk_out,
        txoutclkfabric_out              =>      gt7_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt7_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt7_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt7_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt7_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT8  (X0Y8)
gt8_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT8_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT8_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt8_cpllfbclklost_out,
        cplllock_out                    =>      gt8_cplllock_out,
        cplllockdetclk_in               =>      gt8_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt8_cpllrefclklost_out,
        cpllreset_in                    =>      gt8_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt8_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt8_drpaddr_in,
        drpclk_in                       =>      gt8_drpclk_in,
        drpdi_in                        =>      gt8_drpdi_in,
        drpdo_out                       =>      gt8_drpdo_out,
        drpen_in                        =>      gt8_drpen_in,
        drprdy_out                      =>      gt8_drprdy_out,
        drpwe_in                        =>      gt8_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt8_qpllclk_i,
        qpllrefclk_in                   =>      gt8_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt8_eyescanreset_in,
        rxuserrdy_in                    =>      gt8_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt8_eyescandataerror_out,
        eyescantrigger_in               =>      gt8_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt8_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt8_rxusrclk_in,
        rxusrclk2_in                    =>      gt8_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt8_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt8_rxdisperr_out,
        rxnotintable_out                =>      gt8_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt8_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt8_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt8_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt8_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt8_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt8_rxdfelfhold_in,
        rxmonitorout_out                =>      gt8_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt8_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt8_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt8_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt8_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt8_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt8_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt8_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt8_gttxreset_in,
        txuserrdy_in                    =>      gt8_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt8_txusrclk_in,
        txusrclk2_in                    =>      gt8_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt8_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt8_gthtxn_out,
        gthtxp_out                      =>      gt8_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt8_txoutclk_out,
        txoutclkfabric_out              =>      gt8_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt8_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt8_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt8_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt8_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT9  (X0Y9)
gt9_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT9_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT9_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt9_cpllfbclklost_out,
        cplllock_out                    =>      gt9_cplllock_out,
        cplllockdetclk_in               =>      gt9_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt9_cpllrefclklost_out,
        cpllreset_in                    =>      gt9_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt9_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt9_drpaddr_in,
        drpclk_in                       =>      gt9_drpclk_in,
        drpdi_in                        =>      gt9_drpdi_in,
        drpdo_out                       =>      gt9_drpdo_out,
        drpen_in                        =>      gt9_drpen_in,
        drprdy_out                      =>      gt9_drprdy_out,
        drpwe_in                        =>      gt9_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt9_qpllclk_i,
        qpllrefclk_in                   =>      gt9_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt9_eyescanreset_in,
        rxuserrdy_in                    =>      gt9_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt9_eyescandataerror_out,
        eyescantrigger_in               =>      gt9_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt9_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt9_rxusrclk_in,
        rxusrclk2_in                    =>      gt9_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt9_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt9_rxdisperr_out,
        rxnotintable_out                =>      gt9_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt9_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt9_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt9_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt9_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt9_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt9_rxdfelfhold_in,
        rxmonitorout_out                =>      gt9_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt9_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt9_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt9_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt9_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt9_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt9_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt9_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt9_gttxreset_in,
        txuserrdy_in                    =>      gt9_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt9_txusrclk_in,
        txusrclk2_in                    =>      gt9_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt9_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt9_gthtxn_out,
        gthtxp_out                      =>      gt9_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt9_txoutclk_out,
        txoutclkfabric_out              =>      gt9_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt9_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt9_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt9_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt9_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT10  (X0Y10)
gt10_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT10_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT10_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt10_cpllfbclklost_out,
        cplllock_out                    =>      gt10_cplllock_out,
        cplllockdetclk_in               =>      gt10_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt10_cpllrefclklost_out,
        cpllreset_in                    =>      gt10_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt10_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt10_drpaddr_in,
        drpclk_in                       =>      gt10_drpclk_in,
        drpdi_in                        =>      gt10_drpdi_in,
        drpdo_out                       =>      gt10_drpdo_out,
        drpen_in                        =>      gt10_drpen_in,
        drprdy_out                      =>      gt10_drprdy_out,
        drpwe_in                        =>      gt10_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt10_qpllclk_i,
        qpllrefclk_in                   =>      gt10_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt10_eyescanreset_in,
        rxuserrdy_in                    =>      gt10_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt10_eyescandataerror_out,
        eyescantrigger_in               =>      gt10_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt10_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt10_rxusrclk_in,
        rxusrclk2_in                    =>      gt10_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt10_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt10_rxdisperr_out,
        rxnotintable_out                =>      gt10_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt10_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt10_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt10_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt10_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt10_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt10_rxdfelfhold_in,
        rxmonitorout_out                =>      gt10_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt10_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt10_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt10_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt10_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt10_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt10_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt10_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt10_gttxreset_in,
        txuserrdy_in                    =>      gt10_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt10_txusrclk_in,
        txusrclk2_in                    =>      gt10_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt10_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt10_gthtxn_out,
        gthtxp_out                      =>      gt10_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt10_txoutclk_out,
        txoutclkfabric_out              =>      gt10_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt10_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt10_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt10_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt10_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT11  (X0Y11)
gt11_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT11_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT11_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt11_cpllfbclklost_out,
        cplllock_out                    =>      gt11_cplllock_out,
        cplllockdetclk_in               =>      gt11_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt11_cpllrefclklost_out,
        cpllreset_in                    =>      gt11_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt11_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt11_drpaddr_in,
        drpclk_in                       =>      gt11_drpclk_in,
        drpdi_in                        =>      gt11_drpdi_in,
        drpdo_out                       =>      gt11_drpdo_out,
        drpen_in                        =>      gt11_drpen_in,
        drprdy_out                      =>      gt11_drprdy_out,
        drpwe_in                        =>      gt11_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt11_qpllclk_i,
        qpllrefclk_in                   =>      gt11_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt11_eyescanreset_in,
        rxuserrdy_in                    =>      gt11_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt11_eyescandataerror_out,
        eyescantrigger_in               =>      gt11_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt11_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt11_rxusrclk_in,
        rxusrclk2_in                    =>      gt11_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt11_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt11_rxdisperr_out,
        rxnotintable_out                =>      gt11_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt11_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt11_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt11_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt11_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt11_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt11_rxdfelfhold_in,
        rxmonitorout_out                =>      gt11_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt11_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt11_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt11_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt11_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt11_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt11_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt11_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt11_gttxreset_in,
        txuserrdy_in                    =>      gt11_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt11_txusrclk_in,
        txusrclk2_in                    =>      gt11_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt11_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt11_gthtxn_out,
        gthtxp_out                      =>      gt11_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt11_txoutclk_out,
        txoutclkfabric_out              =>      gt11_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt11_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt11_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt11_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt11_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT12  (X0Y12)
gt12_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT12_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT12_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt12_cpllfbclklost_out,
        cplllock_out                    =>      gt12_cplllock_out,
        cplllockdetclk_in               =>      gt12_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt12_cpllrefclklost_out,
        cpllreset_in                    =>      gt12_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt12_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt12_drpaddr_in,
        drpclk_in                       =>      gt12_drpclk_in,
        drpdi_in                        =>      gt12_drpdi_in,
        drpdo_out                       =>      gt12_drpdo_out,
        drpen_in                        =>      gt12_drpen_in,
        drprdy_out                      =>      gt12_drprdy_out,
        drpwe_in                        =>      gt12_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt12_qpllclk_i,
        qpllrefclk_in                   =>      gt12_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt12_eyescanreset_in,
        rxuserrdy_in                    =>      gt12_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt12_eyescandataerror_out,
        eyescantrigger_in               =>      gt12_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt12_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt12_rxusrclk_in,
        rxusrclk2_in                    =>      gt12_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt12_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt12_rxdisperr_out,
        rxnotintable_out                =>      gt12_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt12_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt12_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt12_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt12_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt12_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt12_rxdfelfhold_in,
        rxmonitorout_out                =>      gt12_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt12_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt12_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt12_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt12_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt12_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt12_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt12_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt12_gttxreset_in,
        txuserrdy_in                    =>      gt12_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt12_txusrclk_in,
        txusrclk2_in                    =>      gt12_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt12_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt12_gthtxn_out,
        gthtxp_out                      =>      gt12_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt12_txoutclk_out,
        txoutclkfabric_out              =>      gt12_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt12_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt12_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt12_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt12_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT13  (X0Y13)
gt13_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT13_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT13_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt13_cpllfbclklost_out,
        cplllock_out                    =>      gt13_cplllock_out,
        cplllockdetclk_in               =>      gt13_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt13_cpllrefclklost_out,
        cpllreset_in                    =>      gt13_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt13_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt13_drpaddr_in,
        drpclk_in                       =>      gt13_drpclk_in,
        drpdi_in                        =>      gt13_drpdi_in,
        drpdo_out                       =>      gt13_drpdo_out,
        drpen_in                        =>      gt13_drpen_in,
        drprdy_out                      =>      gt13_drprdy_out,
        drpwe_in                        =>      gt13_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt13_qpllclk_i,
        qpllrefclk_in                   =>      gt13_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt13_eyescanreset_in,
        rxuserrdy_in                    =>      gt13_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt13_eyescandataerror_out,
        eyescantrigger_in               =>      gt13_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt13_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt13_rxusrclk_in,
        rxusrclk2_in                    =>      gt13_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt13_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt13_rxdisperr_out,
        rxnotintable_out                =>      gt13_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt13_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt13_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt13_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt13_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt13_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt13_rxdfelfhold_in,
        rxmonitorout_out                =>      gt13_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt13_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt13_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt13_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt13_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt13_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt13_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt13_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt13_gttxreset_in,
        txuserrdy_in                    =>      gt13_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt13_txusrclk_in,
        txusrclk2_in                    =>      gt13_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt13_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt13_gthtxn_out,
        gthtxp_out                      =>      gt13_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt13_txoutclk_out,
        txoutclkfabric_out              =>      gt13_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt13_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt13_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt13_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt13_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT14  (X0Y14)
gt14_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT14_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT14_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt14_cpllfbclklost_out,
        cplllock_out                    =>      gt14_cplllock_out,
        cplllockdetclk_in               =>      gt14_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt14_cpllrefclklost_out,
        cpllreset_in                    =>      gt14_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt14_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt14_drpaddr_in,
        drpclk_in                       =>      gt14_drpclk_in,
        drpdi_in                        =>      gt14_drpdi_in,
        drpdo_out                       =>      gt14_drpdo_out,
        drpen_in                        =>      gt14_drpen_in,
        drprdy_out                      =>      gt14_drprdy_out,
        drpwe_in                        =>      gt14_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt14_qpllclk_i,
        qpllrefclk_in                   =>      gt14_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt14_eyescanreset_in,
        rxuserrdy_in                    =>      gt14_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt14_eyescandataerror_out,
        eyescantrigger_in               =>      gt14_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt14_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt14_rxusrclk_in,
        rxusrclk2_in                    =>      gt14_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt14_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt14_rxdisperr_out,
        rxnotintable_out                =>      gt14_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt14_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt14_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt14_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt14_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt14_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt14_rxdfelfhold_in,
        rxmonitorout_out                =>      gt14_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt14_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt14_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt14_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt14_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt14_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt14_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt14_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt14_gttxreset_in,
        txuserrdy_in                    =>      gt14_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt14_txusrclk_in,
        txusrclk2_in                    =>      gt14_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt14_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt14_gthtxn_out,
        gthtxp_out                      =>      gt14_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt14_txoutclk_out,
        txoutclkfabric_out              =>      gt14_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt14_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt14_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt14_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt14_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT15  (X0Y15)
gt15_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT15_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT15_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt15_cpllfbclklost_out,
        cplllock_out                    =>      gt15_cplllock_out,
        cplllockdetclk_in               =>      gt15_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt15_cpllrefclklost_out,
        cpllreset_in                    =>      gt15_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt15_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt15_drpaddr_in,
        drpclk_in                       =>      gt15_drpclk_in,
        drpdi_in                        =>      gt15_drpdi_in,
        drpdo_out                       =>      gt15_drpdo_out,
        drpen_in                        =>      gt15_drpen_in,
        drprdy_out                      =>      gt15_drprdy_out,
        drpwe_in                        =>      gt15_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt15_qpllclk_i,
        qpllrefclk_in                   =>      gt15_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt15_eyescanreset_in,
        rxuserrdy_in                    =>      gt15_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt15_eyescandataerror_out,
        eyescantrigger_in               =>      gt15_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt15_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt15_rxusrclk_in,
        rxusrclk2_in                    =>      gt15_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt15_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt15_rxdisperr_out,
        rxnotintable_out                =>      gt15_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt15_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt15_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt15_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt15_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt15_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt15_rxdfelfhold_in,
        rxmonitorout_out                =>      gt15_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt15_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt15_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt15_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt15_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt15_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt15_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt15_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt15_gttxreset_in,
        txuserrdy_in                    =>      gt15_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt15_txusrclk_in,
        txusrclk2_in                    =>      gt15_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt15_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt15_gthtxn_out,
        gthtxp_out                      =>      gt15_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt15_txoutclk_out,
        txoutclkfabric_out              =>      gt15_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt15_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt15_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt15_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt15_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT16  (X0Y16)
gt16_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT16_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT16_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt16_cpllfbclklost_out,
        cplllock_out                    =>      gt16_cplllock_out,
        cplllockdetclk_in               =>      gt16_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt16_cpllrefclklost_out,
        cpllreset_in                    =>      gt16_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt16_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt16_drpaddr_in,
        drpclk_in                       =>      gt16_drpclk_in,
        drpdi_in                        =>      gt16_drpdi_in,
        drpdo_out                       =>      gt16_drpdo_out,
        drpen_in                        =>      gt16_drpen_in,
        drprdy_out                      =>      gt16_drprdy_out,
        drpwe_in                        =>      gt16_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt16_qpllclk_i,
        qpllrefclk_in                   =>      gt16_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt16_eyescanreset_in,
        rxuserrdy_in                    =>      gt16_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt16_eyescandataerror_out,
        eyescantrigger_in               =>      gt16_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt16_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt16_rxusrclk_in,
        rxusrclk2_in                    =>      gt16_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt16_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt16_rxdisperr_out,
        rxnotintable_out                =>      gt16_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt16_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt16_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt16_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt16_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt16_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt16_rxdfelfhold_in,
        rxmonitorout_out                =>      gt16_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt16_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt16_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt16_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt16_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt16_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt16_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt16_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt16_gttxreset_in,
        txuserrdy_in                    =>      gt16_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt16_txusrclk_in,
        txusrclk2_in                    =>      gt16_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt16_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt16_gthtxn_out,
        gthtxp_out                      =>      gt16_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt16_txoutclk_out,
        txoutclkfabric_out              =>      gt16_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt16_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt16_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt16_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt16_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT17  (X0Y17)
gt17_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT17_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT17_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt17_cpllfbclklost_out,
        cplllock_out                    =>      gt17_cplllock_out,
        cplllockdetclk_in               =>      gt17_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt17_cpllrefclklost_out,
        cpllreset_in                    =>      gt17_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt17_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt17_drpaddr_in,
        drpclk_in                       =>      gt17_drpclk_in,
        drpdi_in                        =>      gt17_drpdi_in,
        drpdo_out                       =>      gt17_drpdo_out,
        drpen_in                        =>      gt17_drpen_in,
        drprdy_out                      =>      gt17_drprdy_out,
        drpwe_in                        =>      gt17_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt17_qpllclk_i,
        qpllrefclk_in                   =>      gt17_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt17_eyescanreset_in,
        rxuserrdy_in                    =>      gt17_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt17_eyescandataerror_out,
        eyescantrigger_in               =>      gt17_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt17_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt17_rxusrclk_in,
        rxusrclk2_in                    =>      gt17_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt17_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt17_rxdisperr_out,
        rxnotintable_out                =>      gt17_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt17_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt17_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt17_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt17_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt17_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt17_rxdfelfhold_in,
        rxmonitorout_out                =>      gt17_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt17_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt17_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt17_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt17_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt17_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt17_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt17_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt17_gttxreset_in,
        txuserrdy_in                    =>      gt17_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt17_txusrclk_in,
        txusrclk2_in                    =>      gt17_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt17_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt17_gthtxn_out,
        gthtxp_out                      =>      gt17_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt17_txoutclk_out,
        txoutclkfabric_out              =>      gt17_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt17_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt17_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt17_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt17_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT18  (X0Y18)
gt18_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT18_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT18_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt18_cpllfbclklost_out,
        cplllock_out                    =>      gt18_cplllock_out,
        cplllockdetclk_in               =>      gt18_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt18_cpllrefclklost_out,
        cpllreset_in                    =>      gt18_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt18_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt18_drpaddr_in,
        drpclk_in                       =>      gt18_drpclk_in,
        drpdi_in                        =>      gt18_drpdi_in,
        drpdo_out                       =>      gt18_drpdo_out,
        drpen_in                        =>      gt18_drpen_in,
        drprdy_out                      =>      gt18_drprdy_out,
        drpwe_in                        =>      gt18_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt18_qpllclk_i,
        qpllrefclk_in                   =>      gt18_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt18_eyescanreset_in,
        rxuserrdy_in                    =>      gt18_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt18_eyescandataerror_out,
        eyescantrigger_in               =>      gt18_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt18_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt18_rxusrclk_in,
        rxusrclk2_in                    =>      gt18_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt18_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt18_rxdisperr_out,
        rxnotintable_out                =>      gt18_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt18_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt18_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt18_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt18_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt18_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt18_rxdfelfhold_in,
        rxmonitorout_out                =>      gt18_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt18_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt18_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt18_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt18_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt18_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt18_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt18_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt18_gttxreset_in,
        txuserrdy_in                    =>      gt18_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt18_txusrclk_in,
        txusrclk2_in                    =>      gt18_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt18_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt18_gthtxn_out,
        gthtxp_out                      =>      gt18_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt18_txoutclk_out,
        txoutclkfabric_out              =>      gt18_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt18_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt18_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt18_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt18_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT19  (X0Y19)
gt19_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT19_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT19_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt19_cpllfbclklost_out,
        cplllock_out                    =>      gt19_cplllock_out,
        cplllockdetclk_in               =>      gt19_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt19_cpllrefclklost_out,
        cpllreset_in                    =>      gt19_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt19_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt19_drpaddr_in,
        drpclk_in                       =>      gt19_drpclk_in,
        drpdi_in                        =>      gt19_drpdi_in,
        drpdo_out                       =>      gt19_drpdo_out,
        drpen_in                        =>      gt19_drpen_in,
        drprdy_out                      =>      gt19_drprdy_out,
        drpwe_in                        =>      gt19_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt19_qpllclk_i,
        qpllrefclk_in                   =>      gt19_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt19_eyescanreset_in,
        rxuserrdy_in                    =>      gt19_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt19_eyescandataerror_out,
        eyescantrigger_in               =>      gt19_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt19_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt19_rxusrclk_in,
        rxusrclk2_in                    =>      gt19_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt19_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt19_rxdisperr_out,
        rxnotintable_out                =>      gt19_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt19_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt19_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt19_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt19_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt19_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt19_rxdfelfhold_in,
        rxmonitorout_out                =>      gt19_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt19_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt19_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt19_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt19_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt19_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt19_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt19_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt19_gttxreset_in,
        txuserrdy_in                    =>      gt19_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt19_txusrclk_in,
        txusrclk2_in                    =>      gt19_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt19_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt19_gthtxn_out,
        gthtxp_out                      =>      gt19_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt19_txoutclk_out,
        txoutclkfabric_out              =>      gt19_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt19_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt19_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt19_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt19_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT20  (X0Y20)
gt20_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT20_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT20_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt20_cpllfbclklost_out,
        cplllock_out                    =>      gt20_cplllock_out,
        cplllockdetclk_in               =>      gt20_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt20_cpllrefclklost_out,
        cpllreset_in                    =>      gt20_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt20_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt20_drpaddr_in,
        drpclk_in                       =>      gt20_drpclk_in,
        drpdi_in                        =>      gt20_drpdi_in,
        drpdo_out                       =>      gt20_drpdo_out,
        drpen_in                        =>      gt20_drpen_in,
        drprdy_out                      =>      gt20_drprdy_out,
        drpwe_in                        =>      gt20_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt20_qpllclk_i,
        qpllrefclk_in                   =>      gt20_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt20_eyescanreset_in,
        rxuserrdy_in                    =>      gt20_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt20_eyescandataerror_out,
        eyescantrigger_in               =>      gt20_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt20_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt20_rxusrclk_in,
        rxusrclk2_in                    =>      gt20_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt20_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt20_rxdisperr_out,
        rxnotintable_out                =>      gt20_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt20_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt20_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt20_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt20_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt20_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt20_rxdfelfhold_in,
        rxmonitorout_out                =>      gt20_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt20_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt20_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt20_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt20_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt20_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt20_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt20_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt20_gttxreset_in,
        txuserrdy_in                    =>      gt20_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt20_txusrclk_in,
        txusrclk2_in                    =>      gt20_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt20_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt20_gthtxn_out,
        gthtxp_out                      =>      gt20_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt20_txoutclk_out,
        txoutclkfabric_out              =>      gt20_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt20_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt20_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt20_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt20_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT21  (X0Y21)
gt21_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT21_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT21_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt21_cpllfbclklost_out,
        cplllock_out                    =>      gt21_cplllock_out,
        cplllockdetclk_in               =>      gt21_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt21_cpllrefclklost_out,
        cpllreset_in                    =>      gt21_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt21_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt21_drpaddr_in,
        drpclk_in                       =>      gt21_drpclk_in,
        drpdi_in                        =>      gt21_drpdi_in,
        drpdo_out                       =>      gt21_drpdo_out,
        drpen_in                        =>      gt21_drpen_in,
        drprdy_out                      =>      gt21_drprdy_out,
        drpwe_in                        =>      gt21_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt21_qpllclk_i,
        qpllrefclk_in                   =>      gt21_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt21_eyescanreset_in,
        rxuserrdy_in                    =>      gt21_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt21_eyescandataerror_out,
        eyescantrigger_in               =>      gt21_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt21_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt21_rxusrclk_in,
        rxusrclk2_in                    =>      gt21_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt21_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt21_rxdisperr_out,
        rxnotintable_out                =>      gt21_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt21_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt21_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt21_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt21_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt21_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt21_rxdfelfhold_in,
        rxmonitorout_out                =>      gt21_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt21_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt21_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt21_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt21_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt21_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt21_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt21_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt21_gttxreset_in,
        txuserrdy_in                    =>      gt21_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt21_txusrclk_in,
        txusrclk2_in                    =>      gt21_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt21_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt21_gthtxn_out,
        gthtxp_out                      =>      gt21_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt21_txoutclk_out,
        txoutclkfabric_out              =>      gt21_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt21_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt21_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt21_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt21_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT22  (X0Y22)
gt22_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT22_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT22_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt22_cpllfbclklost_out,
        cplllock_out                    =>      gt22_cplllock_out,
        cplllockdetclk_in               =>      gt22_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt22_cpllrefclklost_out,
        cpllreset_in                    =>      gt22_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt22_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt22_drpaddr_in,
        drpclk_in                       =>      gt22_drpclk_in,
        drpdi_in                        =>      gt22_drpdi_in,
        drpdo_out                       =>      gt22_drpdo_out,
        drpen_in                        =>      gt22_drpen_in,
        drprdy_out                      =>      gt22_drprdy_out,
        drpwe_in                        =>      gt22_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt22_qpllclk_i,
        qpllrefclk_in                   =>      gt22_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt22_eyescanreset_in,
        rxuserrdy_in                    =>      gt22_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt22_eyescandataerror_out,
        eyescantrigger_in               =>      gt22_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt22_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt22_rxusrclk_in,
        rxusrclk2_in                    =>      gt22_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt22_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt22_rxdisperr_out,
        rxnotintable_out                =>      gt22_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt22_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt22_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt22_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt22_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt22_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt22_rxdfelfhold_in,
        rxmonitorout_out                =>      gt22_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt22_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt22_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt22_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt22_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt22_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt22_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt22_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt22_gttxreset_in,
        txuserrdy_in                    =>      gt22_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt22_txusrclk_in,
        txusrclk2_in                    =>      gt22_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt22_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt22_gthtxn_out,
        gthtxp_out                      =>      gt22_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt22_txoutclk_out,
        txoutclkfabric_out              =>      gt22_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt22_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt22_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt22_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt22_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT23  (X0Y23)
gt23_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT23_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT23_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt23_cpllfbclklost_out,
        cplllock_out                    =>      gt23_cplllock_out,
        cplllockdetclk_in               =>      gt23_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt23_cpllrefclklost_out,
        cpllreset_in                    =>      gt23_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt23_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt23_drpaddr_in,
        drpclk_in                       =>      gt23_drpclk_in,
        drpdi_in                        =>      gt23_drpdi_in,
        drpdo_out                       =>      gt23_drpdo_out,
        drpen_in                        =>      gt23_drpen_in,
        drprdy_out                      =>      gt23_drprdy_out,
        drpwe_in                        =>      gt23_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt23_qpllclk_i,
        qpllrefclk_in                   =>      gt23_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt23_eyescanreset_in,
        rxuserrdy_in                    =>      gt23_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt23_eyescandataerror_out,
        eyescantrigger_in               =>      gt23_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt23_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt23_rxusrclk_in,
        rxusrclk2_in                    =>      gt23_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt23_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt23_rxdisperr_out,
        rxnotintable_out                =>      gt23_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt23_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt23_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt23_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt23_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt23_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt23_rxdfelfhold_in,
        rxmonitorout_out                =>      gt23_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt23_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt23_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt23_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt23_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt23_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt23_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt23_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt23_gttxreset_in,
        txuserrdy_in                    =>      gt23_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt23_txusrclk_in,
        txusrclk2_in                    =>      gt23_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt23_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt23_gthtxn_out,
        gthtxp_out                      =>      gt23_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt23_txoutclk_out,
        txoutclkfabric_out              =>      gt23_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt23_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt23_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt23_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt23_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT24  (X0Y24)
gt24_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT24_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT24_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt24_cpllfbclklost_out,
        cplllock_out                    =>      gt24_cplllock_out,
        cplllockdetclk_in               =>      gt24_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt24_cpllrefclklost_out,
        cpllreset_in                    =>      gt24_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt24_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt24_drpaddr_in,
        drpclk_in                       =>      gt24_drpclk_in,
        drpdi_in                        =>      gt24_drpdi_in,
        drpdo_out                       =>      gt24_drpdo_out,
        drpen_in                        =>      gt24_drpen_in,
        drprdy_out                      =>      gt24_drprdy_out,
        drpwe_in                        =>      gt24_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt24_qpllclk_i,
        qpllrefclk_in                   =>      gt24_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt24_eyescanreset_in,
        rxuserrdy_in                    =>      gt24_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt24_eyescandataerror_out,
        eyescantrigger_in               =>      gt24_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt24_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt24_rxusrclk_in,
        rxusrclk2_in                    =>      gt24_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt24_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt24_rxdisperr_out,
        rxnotintable_out                =>      gt24_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt24_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt24_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt24_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt24_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt24_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt24_rxdfelfhold_in,
        rxmonitorout_out                =>      gt24_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt24_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt24_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt24_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt24_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt24_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt24_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt24_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt24_gttxreset_in,
        txuserrdy_in                    =>      gt24_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt24_txusrclk_in,
        txusrclk2_in                    =>      gt24_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt24_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt24_gthtxn_out,
        gthtxp_out                      =>      gt24_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt24_txoutclk_out,
        txoutclkfabric_out              =>      gt24_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt24_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt24_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt24_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt24_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT25  (X0Y25)
gt25_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT25_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT25_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt25_cpllfbclklost_out,
        cplllock_out                    =>      gt25_cplllock_out,
        cplllockdetclk_in               =>      gt25_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt25_cpllrefclklost_out,
        cpllreset_in                    =>      gt25_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt25_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt25_drpaddr_in,
        drpclk_in                       =>      gt25_drpclk_in,
        drpdi_in                        =>      gt25_drpdi_in,
        drpdo_out                       =>      gt25_drpdo_out,
        drpen_in                        =>      gt25_drpen_in,
        drprdy_out                      =>      gt25_drprdy_out,
        drpwe_in                        =>      gt25_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt25_qpllclk_i,
        qpllrefclk_in                   =>      gt25_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt25_eyescanreset_in,
        rxuserrdy_in                    =>      gt25_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt25_eyescandataerror_out,
        eyescantrigger_in               =>      gt25_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt25_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt25_rxusrclk_in,
        rxusrclk2_in                    =>      gt25_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt25_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt25_rxdisperr_out,
        rxnotintable_out                =>      gt25_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt25_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt25_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt25_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt25_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt25_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt25_rxdfelfhold_in,
        rxmonitorout_out                =>      gt25_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt25_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt25_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt25_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt25_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt25_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt25_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt25_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt25_gttxreset_in,
        txuserrdy_in                    =>      gt25_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt25_txusrclk_in,
        txusrclk2_in                    =>      gt25_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt25_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt25_gthtxn_out,
        gthtxp_out                      =>      gt25_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt25_txoutclk_out,
        txoutclkfabric_out              =>      gt25_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt25_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt25_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt25_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt25_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT26  (X0Y26)
gt26_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT26_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT26_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt26_cpllfbclklost_out,
        cplllock_out                    =>      gt26_cplllock_out,
        cplllockdetclk_in               =>      gt26_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt26_cpllrefclklost_out,
        cpllreset_in                    =>      gt26_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt26_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt26_drpaddr_in,
        drpclk_in                       =>      gt26_drpclk_in,
        drpdi_in                        =>      gt26_drpdi_in,
        drpdo_out                       =>      gt26_drpdo_out,
        drpen_in                        =>      gt26_drpen_in,
        drprdy_out                      =>      gt26_drprdy_out,
        drpwe_in                        =>      gt26_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt26_qpllclk_i,
        qpllrefclk_in                   =>      gt26_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt26_eyescanreset_in,
        rxuserrdy_in                    =>      gt26_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt26_eyescandataerror_out,
        eyescantrigger_in               =>      gt26_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt26_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt26_rxusrclk_in,
        rxusrclk2_in                    =>      gt26_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt26_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt26_rxdisperr_out,
        rxnotintable_out                =>      gt26_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt26_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt26_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt26_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt26_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt26_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt26_rxdfelfhold_in,
        rxmonitorout_out                =>      gt26_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt26_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt26_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt26_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt26_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt26_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt26_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt26_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt26_gttxreset_in,
        txuserrdy_in                    =>      gt26_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt26_txusrclk_in,
        txusrclk2_in                    =>      gt26_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt26_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt26_gthtxn_out,
        gthtxp_out                      =>      gt26_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt26_txoutclk_out,
        txoutclkfabric_out              =>      gt26_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt26_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt26_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt26_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt26_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT27  (X0Y27)
gt27_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT27_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT27_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt27_cpllfbclklost_out,
        cplllock_out                    =>      gt27_cplllock_out,
        cplllockdetclk_in               =>      gt27_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt27_cpllrefclklost_out,
        cpllreset_in                    =>      gt27_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt27_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt27_drpaddr_in,
        drpclk_in                       =>      gt27_drpclk_in,
        drpdi_in                        =>      gt27_drpdi_in,
        drpdo_out                       =>      gt27_drpdo_out,
        drpen_in                        =>      gt27_drpen_in,
        drprdy_out                      =>      gt27_drprdy_out,
        drpwe_in                        =>      gt27_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt27_qpllclk_i,
        qpllrefclk_in                   =>      gt27_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt27_eyescanreset_in,
        rxuserrdy_in                    =>      gt27_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt27_eyescandataerror_out,
        eyescantrigger_in               =>      gt27_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt27_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt27_rxusrclk_in,
        rxusrclk2_in                    =>      gt27_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt27_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt27_rxdisperr_out,
        rxnotintable_out                =>      gt27_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt27_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt27_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt27_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt27_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt27_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt27_rxdfelfhold_in,
        rxmonitorout_out                =>      gt27_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt27_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt27_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt27_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt27_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt27_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt27_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt27_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt27_gttxreset_in,
        txuserrdy_in                    =>      gt27_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt27_txusrclk_in,
        txusrclk2_in                    =>      gt27_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt27_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt27_gthtxn_out,
        gthtxp_out                      =>      gt27_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt27_txoutclk_out,
        txoutclkfabric_out              =>      gt27_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt27_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt27_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt27_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt27_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT28  (X0Y28)
gt28_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT28_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT28_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt28_cpllfbclklost_out,
        cplllock_out                    =>      gt28_cplllock_out,
        cplllockdetclk_in               =>      gt28_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt28_cpllrefclklost_out,
        cpllreset_in                    =>      gt28_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt28_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt28_drpaddr_in,
        drpclk_in                       =>      gt28_drpclk_in,
        drpdi_in                        =>      gt28_drpdi_in,
        drpdo_out                       =>      gt28_drpdo_out,
        drpen_in                        =>      gt28_drpen_in,
        drprdy_out                      =>      gt28_drprdy_out,
        drpwe_in                        =>      gt28_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt28_qpllclk_i,
        qpllrefclk_in                   =>      gt28_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt28_eyescanreset_in,
        rxuserrdy_in                    =>      gt28_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt28_eyescandataerror_out,
        eyescantrigger_in               =>      gt28_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt28_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt28_rxusrclk_in,
        rxusrclk2_in                    =>      gt28_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt28_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt28_rxdisperr_out,
        rxnotintable_out                =>      gt28_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt28_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt28_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt28_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt28_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt28_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt28_rxdfelfhold_in,
        rxmonitorout_out                =>      gt28_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt28_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt28_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt28_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt28_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt28_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt28_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt28_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt28_gttxreset_in,
        txuserrdy_in                    =>      gt28_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt28_txusrclk_in,
        txusrclk2_in                    =>      gt28_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt28_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt28_gthtxn_out,
        gthtxp_out                      =>      gt28_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt28_txoutclk_out,
        txoutclkfabric_out              =>      gt28_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt28_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt28_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt28_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt28_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT29  (X0Y29)
gt29_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT29_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT29_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt29_cpllfbclklost_out,
        cplllock_out                    =>      gt29_cplllock_out,
        cplllockdetclk_in               =>      gt29_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt29_cpllrefclklost_out,
        cpllreset_in                    =>      gt29_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt29_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt29_drpaddr_in,
        drpclk_in                       =>      gt29_drpclk_in,
        drpdi_in                        =>      gt29_drpdi_in,
        drpdo_out                       =>      gt29_drpdo_out,
        drpen_in                        =>      gt29_drpen_in,
        drprdy_out                      =>      gt29_drprdy_out,
        drpwe_in                        =>      gt29_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt29_qpllclk_i,
        qpllrefclk_in                   =>      gt29_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt29_eyescanreset_in,
        rxuserrdy_in                    =>      gt29_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt29_eyescandataerror_out,
        eyescantrigger_in               =>      gt29_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt29_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt29_rxusrclk_in,
        rxusrclk2_in                    =>      gt29_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt29_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt29_rxdisperr_out,
        rxnotintable_out                =>      gt29_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt29_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt29_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt29_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt29_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt29_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt29_rxdfelfhold_in,
        rxmonitorout_out                =>      gt29_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt29_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt29_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt29_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt29_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt29_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt29_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt29_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt29_gttxreset_in,
        txuserrdy_in                    =>      gt29_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt29_txusrclk_in,
        txusrclk2_in                    =>      gt29_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt29_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt29_gthtxn_out,
        gthtxp_out                      =>      gt29_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt29_txoutclk_out,
        txoutclkfabric_out              =>      gt29_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt29_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt29_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt29_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt29_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT30  (X0Y30)
gt30_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT30_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT30_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt30_cpllfbclklost_out,
        cplllock_out                    =>      gt30_cplllock_out,
        cplllockdetclk_in               =>      gt30_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt30_cpllrefclklost_out,
        cpllreset_in                    =>      gt30_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt30_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt30_drpaddr_in,
        drpclk_in                       =>      gt30_drpclk_in,
        drpdi_in                        =>      gt30_drpdi_in,
        drpdo_out                       =>      gt30_drpdo_out,
        drpen_in                        =>      gt30_drpen_in,
        drprdy_out                      =>      gt30_drprdy_out,
        drpwe_in                        =>      gt30_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt30_qpllclk_i,
        qpllrefclk_in                   =>      gt30_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt30_eyescanreset_in,
        rxuserrdy_in                    =>      gt30_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt30_eyescandataerror_out,
        eyescantrigger_in               =>      gt30_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt30_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt30_rxusrclk_in,
        rxusrclk2_in                    =>      gt30_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt30_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt30_rxdisperr_out,
        rxnotintable_out                =>      gt30_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt30_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt30_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt30_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt30_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt30_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt30_rxdfelfhold_in,
        rxmonitorout_out                =>      gt30_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt30_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt30_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt30_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt30_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt30_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt30_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt30_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt30_gttxreset_in,
        txuserrdy_in                    =>      gt30_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt30_txusrclk_in,
        txusrclk2_in                    =>      gt30_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt30_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt30_gthtxn_out,
        gthtxp_out                      =>      gt30_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt30_txoutclk_out,
        txoutclkfabric_out              =>      gt30_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt30_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt30_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt30_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt30_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT31  (X0Y31)
gt31_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT31_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT31_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt31_cpllfbclklost_out,
        cplllock_out                    =>      gt31_cplllock_out,
        cplllockdetclk_in               =>      gt31_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt31_cpllrefclklost_out,
        cpllreset_in                    =>      gt31_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt31_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt31_drpaddr_in,
        drpclk_in                       =>      gt31_drpclk_in,
        drpdi_in                        =>      gt31_drpdi_in,
        drpdo_out                       =>      gt31_drpdo_out,
        drpen_in                        =>      gt31_drpen_in,
        drprdy_out                      =>      gt31_drprdy_out,
        drpwe_in                        =>      gt31_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt31_qpllclk_i,
        qpllrefclk_in                   =>      gt31_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt31_eyescanreset_in,
        rxuserrdy_in                    =>      gt31_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt31_eyescandataerror_out,
        eyescantrigger_in               =>      gt31_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt31_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt31_rxusrclk_in,
        rxusrclk2_in                    =>      gt31_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt31_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt31_rxdisperr_out,
        rxnotintable_out                =>      gt31_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt31_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt31_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt31_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt31_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt31_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt31_rxdfelfhold_in,
        rxmonitorout_out                =>      gt31_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt31_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt31_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt31_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt31_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt31_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt31_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt31_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt31_gttxreset_in,
        txuserrdy_in                    =>      gt31_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt31_txusrclk_in,
        txusrclk2_in                    =>      gt31_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt31_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt31_gthtxn_out,
        gthtxp_out                      =>      gt31_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt31_txoutclk_out,
        txoutclkfabric_out              =>      gt31_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt31_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt31_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt31_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt31_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT32  (X0Y32)
gt32_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT32_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT32_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt32_cpllfbclklost_out,
        cplllock_out                    =>      gt32_cplllock_out,
        cplllockdetclk_in               =>      gt32_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt32_cpllrefclklost_out,
        cpllreset_in                    =>      gt32_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt32_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt32_drpaddr_in,
        drpclk_in                       =>      gt32_drpclk_in,
        drpdi_in                        =>      gt32_drpdi_in,
        drpdo_out                       =>      gt32_drpdo_out,
        drpen_in                        =>      gt32_drpen_in,
        drprdy_out                      =>      gt32_drprdy_out,
        drpwe_in                        =>      gt32_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt32_qpllclk_i,
        qpllrefclk_in                   =>      gt32_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt32_eyescanreset_in,
        rxuserrdy_in                    =>      gt32_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt32_eyescandataerror_out,
        eyescantrigger_in               =>      gt32_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt32_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt32_rxusrclk_in,
        rxusrclk2_in                    =>      gt32_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt32_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt32_rxdisperr_out,
        rxnotintable_out                =>      gt32_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt32_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt32_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt32_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt32_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt32_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt32_rxdfelfhold_in,
        rxmonitorout_out                =>      gt32_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt32_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt32_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt32_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt32_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt32_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt32_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt32_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt32_gttxreset_in,
        txuserrdy_in                    =>      gt32_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt32_txusrclk_in,
        txusrclk2_in                    =>      gt32_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt32_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt32_gthtxn_out,
        gthtxp_out                      =>      gt32_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt32_txoutclk_out,
        txoutclkfabric_out              =>      gt32_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt32_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt32_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt32_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt32_txcharisk_in

    );

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT33  (X0Y33)
gt33_gt6_rtm34l_i : gt6_rtm34l_GT
    generic map
    (
        -- Simulation attributes
        GT_SIM_GTRESET_SPEEDUP => WRAPPER_SIM_GTRESET_SPEEDUP,
        EXAMPLE_SIMULATION     => EXAMPLE_SIMULATION,
        TXSYNC_OVRD_IN         => ('0'),
        TXSYNC_MULTILANE_IN    => ('0')
    )
    port map
    (
        RXPMARESETDONE                  =>      GT33_RXPMARESETDONE_OUT,
        TXPMARESETDONE                  =>      GT33_TXPMARESETDONE_OUT,

        --------------------------------- CPLL Ports -------------------------------
        cpllfbclklost_out               =>      gt33_cpllfbclklost_out,
        cplllock_out                    =>      gt33_cplllock_out,
        cplllockdetclk_in               =>      gt33_cplllockdetclk_in,
        cpllrefclklost_out              =>      gt33_cpllrefclklost_out,
        cpllreset_in                    =>      gt33_cpllreset_in,
        -------------------------- Channel - Clocking Ports ------------------------
        gtrefclk0_in                    =>      gt33_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        drpaddr_in                      =>      gt33_drpaddr_in,
        drpclk_in                       =>      gt33_drpclk_in,
        drpdi_in                        =>      gt33_drpdi_in,
        drpdo_out                       =>      gt33_drpdo_out,
        drpen_in                        =>      gt33_drpen_in,
        drprdy_out                      =>      gt33_drprdy_out,
        drpwe_in                        =>      gt33_drpwe_in,
        ------------------------------- Clocking Ports -----------------------------
        qpllclk_in                      =>      gt33_qpllclk_i,
        qpllrefclk_in                   =>      gt33_qpllrefclk_i,
        --------------------- RX Initialization and Reset Ports --------------------
        eyescanreset_in                 =>      gt33_eyescanreset_in,
        rxuserrdy_in                    =>      gt33_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        eyescandataerror_out            =>      gt33_eyescandataerror_out,
        eyescantrigger_in               =>      gt33_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        dmonitorout_out                 =>      gt33_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        rxusrclk_in                     =>      gt33_rxusrclk_in,
        rxusrclk2_in                    =>      gt33_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        rxdata_out                      =>      gt33_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        rxdisperr_out                   =>      gt33_rxdisperr_out,
        rxnotintable_out                =>      gt33_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gthrxn_in                       =>      gt33_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        rxbyteisaligned_out             =>      gt33_rxbyteisaligned_out,
        rxmcommaalignen_in              =>      gt33_rxmcommaalignen_in,
        rxpcommaalignen_in              =>      gt33_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        rxdfeagchold_in                 =>      gt33_rxdfeagchold_in,
        rxdfelfhold_in                  =>      gt33_rxdfelfhold_in,
        rxmonitorout_out                =>      gt33_rxmonitorout_out,
        rxmonitorsel_in                 =>      gt33_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        rxoutclk_out                    =>      gt33_rxoutclk_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gtrxreset_in                    =>      gt33_gtrxreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        rxpolarity_in                   =>      gt33_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        rxcharisk_out                   =>      gt33_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gthrxp_in                       =>      gt33_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        rxresetdone_out                 =>      gt33_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gttxreset_in                    =>      gt33_gttxreset_in,
        txuserrdy_in                    =>      gt33_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        txusrclk_in                     =>      gt33_txusrclk_in,
        txusrclk2_in                    =>      gt33_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        txdata_in                       =>      gt33_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gthtxn_out                      =>      gt33_gthtxn_out,
        gthtxp_out                      =>      gt33_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        txoutclk_out                    =>      gt33_txoutclk_out,
        txoutclkfabric_out              =>      gt33_txoutclkfabric_out,
        txoutclkpcs_out                 =>      gt33_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        txresetdone_out                 =>      gt33_txresetdone_out,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        txpolarity_in                   =>      gt33_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        txcharisk_in                    =>      gt33_txcharisk_in

    );


end RTL;
     
