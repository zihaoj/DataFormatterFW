

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QSlXH1KsKzDhMmuFBHpGFltPOGW6N2Nj/hR6wdz3GuFzdUyI73737RJtFqsiK4qgZqEY1tQue/c7
7H1YdFBcwQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FYqAcQ5nDnAP8qgwssOu6X5Y1/tiiXvg67DbVwa5HxrUahAjGi2tTl98n1DzLh4Z1jxHUstq4Fbg
WQwhIvMrEqvhtpOvBtRnrcAk82rkwIaBx5US08XKiCa9vkoMVNxZuZtwZTtrIM+9XUCO0ktmmPud
c08nxWNTQfg9hJ/b0n4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FjiSfv1bqWDMy6VzwRiW8VvhyS1saopqgAtovzmwm1cnei1d+AIzCwmR9dq2SjjBdQO2Fp/7L1vz
+UDC6Hoxv2bAr80IPb3OeByMC4PCaxWv6ZvnvQQKNeRbJdTihM1tavIitoWKGZHZUe3DQJyA2v06
DQBrSANGgEtOTUnt6tMy4dXMEIIZEWL0kL4IHy3WpDDif3d22xjAhFs3IscnUHqBynUrRy/VqA6q
fa49+QHq5sbAxHk9++bIP/bIIHvPtMMX56sVlDpZrRHJAWD4z/9ywl6NKvyZUuCmr/P6fA7rvBdo
3DCKxw2xp7ADQDsIjc/btZm2gugsXr+Bt1MuhQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o6DITVWwmnuy4+wsTemDOhT5TgoR8pvcv095fm91DzJt4bH/tISw1sAoTZUIM4aoMdidZbT81xNb
h8WqldC4ZdyVwZala5GRygNAuoUM9B25klGvzObmlNOGDchRuXoY/yDOhdp9O1k/bSOw3XvsPf22
UUOtzKeU1tEUNA0HCnE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ry4z6bB+eq7IVp32fBmDwE9VOaQNhDItOKWcz1tcafjSatrrqNfC4PuY2PxtPAHpJ0jSdYmLGeaa
ocEUIIyQk+UdRAga/cqX5xIJlWUXMzktat/PIvNXSPjouFsR6BX+J/XivrHLzzWuH1LTc663x/qA
xmTkreXa4QocIiBH5YAXHcEYhMVsqPcpKo9F1lW/othnEKkEdidP1RoHkyQCgpHJB37JJkg1ZLjM
yJ0ZKiZMCJs/lb20ZF2q0O1KJ5ElRH5GBzmYI3bc75ny9+iL5cF3G7M61s1CZwZqf2r8NKJAfQve
1o0xRTHtV5COmn7+rD6TMFnsY1hIs6XkKg3/XQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5008)
`protect data_block
y90rGt0re7CItT6XiUJnaSJd2MCt6ZoCnH23xR5W9Dq7YX1yblf/Q2xM4RhdJ0Sz7c3rUXvJ7gKG
LiEpJ6L5GqhpbK5zgAAP3nqP3EZKvDPq6/34O7brQHpZSLiPCyB2+eJvAJ2nhQInIWktvRUPJbdj
wKN/93HQssyOtSQFiN/ueotO1QISjjMnW+q2UXCd8GNmtSODNmwtLkW6kEKzus+SQLvokkBP5YTf
amq0AuSghbMhLeUOE3Qta71KRMVPp8DHdv9k4Qoy7LWjFYyu/6FbhwGh6Rcl3hTJ4hFRMIp1pBiL
sgyvbO3/AhiX4jynyAF4wI1TPLV1zERpF90WOjLk5tPgmmWj4H1JBQ561VEADIK5+zlMoPCwnaoZ
lZane9yGgjLUuvMZaV/RYJhrvlzJXOH92Fl/0XlXyEubIqbGsxov2gQ7MIDhpOa10k3YfK0eGD5w
zx14KTmWXYtNSy0fDQm5GmUAtrtZbn/9ji/E75bPxpLPv+pta6tyFs58ztfTh7qONHx9ovL1qBzx
wP/6S4RD0s4yWb0C4X0rqdWGtlK9hRwvYvTnICgEvfDn27VOIMLMsbz/uuoXn0+lXMXV+ImzLXy+
Ft2xl3SaAUxlzW8kJxGxG0EZMdO49rgWdXK2VOZa8ZTeUhWN4qu/oPX//zlJp5dmHSWnL7RsvAx1
DA1a3nC0MFh2JawbMLEGMyxPBF9cjbdkZkADzBDhUG5GhpTFUXnqrUh6bRPciV8n63SsxVvqF7rH
Os09dxbc+OxSJftdQWIoo7F0YjHdPr7C4XdoQGuaSLnm3crIfjjp4Wm02o6Z041FFNbiXbBdkzG3
vEM+788BFKPzL5cKWflnma1zNq+ZSo6iH8kcG0iqQAaX2/YSZxwrXzDuj+2VRErxjtJe4joa4U8W
aBFrDHpZmrFkpnnRX7xw9r4m4pfPNwO08tVCoqo2r6C4nFv30UbyBtoh3DxUnlLWjdsuClB7mALx
SNRNInrR8SxAWIlQdFkvYGyfsV1zeRYuIYuYtCF2/ZkZ2bk0F+uurHKO38XT79oPPCa+sc8V2hBG
fAcnm9uFBzFrnZuhhNuA3oEs1E8Y0yzaAES0dEqodRYFuhGd5GOcdPswvFk5LdoLY5jQl7yRc4FH
5nkR4OnLLphZKmU9/e8dioRnFqrkJ1sPVM5lyhMLIj+OQyZuBQbXU1BUFjUC/3BkC7UmV7t6ETm6
+SjulSntEBUggPkpCEINw69uobOrmdfZVkLxydGtIpd2eHNuNHYlIPGEOJXV7Qg9mZJA3+3MUtY/
p91Do6hrYWoZ4bNrxsgKbDbuoZR4yk7lU9jfuw56CODNrlPuxyOHGw3jXdKr27/ImbGsWr0zbI1X
o62gj811Q2PSPp3PYqotHZ8wOmDcNmyJd0TiiYkMJBD61ZsCbJib3E7zgUuOPWBGkgW7vTiKhTc2
/e2ZFa3Z9AB5HVDkcJdpyi0Q/nItRlXShHyDIEULj1ZzrBtCJ6hm0KhX0x850sIQyes05+lK9hpl
Suf8wUcKPj79XJF37KmZjlIgmexraryl0PkD83FIvaCGytvOzl8dfe6oC4IjgY9WlI1aI6SLBcdm
wEh1CaQocnNNLykI/8G/uMlYsP6dhnlSCAPZZdLvoUFkmmp/VtX34qO5GtXR4OVPsEaqw/XM7aMP
KAsDJEIGWehd/gmeEbO0li8cgP6biUIUtvdu1nk3u2QqEG5u4f46cz9oalStbcut8WGP+ae/jQAA
JCaDkrknqKlyiNNEand01FE/tFv2SSDXthsvGd3OZMiiweWFN6LCHcZYRja5mLd/bRy4G/gTmSPq
ddSMBarwQS5XA6ijz4+ZnQ2ve2Ab6e5uc6B+aiR6KmHUxAY+SIaf0YuVIMunuq1EgZ4W9XoaegGv
8ys9AJde1JXAnpeeM/4qMfAJ78wWgbbbCDfRy13cRC2t6rW2d0wSlFY0hBPLHCrSSu6G4EkVlIaE
jyqlQWKZdl5jVpxMngbCuZ0CcOYtPVUNh5NJ8XzMWvzK2/jysWaI674LDpARR74IbAKKnk75q5Bs
tejSl/Z+Ea2tqA4+Ql7ZjQXVXNhQBuAm7Vdw/qfH7HzDDa4r0IIRYyOhkuo6ujCPOz0IlYe9Flgn
M+AvDiVWLA4Pxj4/raKWQ3sOEJzs7qpxomcuVkhcSbWIa2KQj8adM2EQVvoCIIIpzQZ4FF2x+bSa
Ugq1N416MgoK21if/RBysTkczQQOA9pMQewZb8LUn6bezqQr8Nvnq78z29JJORhGbzebzIk7+Zrm
DQEPl6iO2+Az2NUBnCMlsxmTgIQvhE0p/p/gvt8wAGofFEuj7Zyz938ciopJEeQFr/YzAWRwV/Oq
0AfeIMhVXpKMmXwuD4oP4apDx3kXWcb6sUksGgMExLOLn7sF/I1icwd2L6yRI82cVfCh5VJtxG+m
tawE8b8bpKeNXxWBnf6ZGmtd8vxQYBvnNmhMyf3I7hmsYbS7tr4zyoudkFZP5s5OHvp9lq+Ampce
21sjm5HPABmvOvFfRhcm8PoiDJuMY6Cy7JwP6eHqaRlg3TiLjYU4pg6cf0zFzH5o5fXq1B8bqOEj
3DIoyAU3dgoxBkgsxEtFajb6k5uEADeHTPh1bqOG03PAKd+DDxC/2AW8zioe1hr0eX4BhiWihAEb
lOqEBtLjBCGZjp/TcINmtZ3Ln2TAhufaok/5bGcswCLdT/nBoUSlOk5n/qDZJ7yeKI7vCWPsXvlf
rsYPpmSTBqcuuW1rBTpdpBpTqPNpIGBRQhF8hAKdzv8UHkV1U1gKJwWzbfFMigAhjCSa45U2bOlp
HYhMm2xTuhkW1B/WsWlySE3E/G8h0NCSAJtz17f/OYTpEVFcLWzlzO24vEWO+SvKEf+PBik7/6GL
RCY9VhV5i25q8ALMY1jZ64ZHYXPYN1+0B0gxJQLFXObT6YMV2po3hINvAJRKa+D2uDVfHYtcHQ6y
7HAQqZ74MoWDDy4Iv9yti3KxhwjE7jc4DrG7m2DVHSxQlVEmGYzELpegDEkrsorLcPYYPPtheqKZ
SrdVO2wSgpo2KKvgPnQaR1SeKlCpsVPIP2UCaBX9qVbLycbdo2ObBVTffWVo/L/nEsJgkoURe/Ez
jhyk/4efAFZbQNdZWUfFSB24EtIgBza7xFugA2yqRTEyKINcQr22WVA+gUDqQsQ0fbMwI2y5/JJz
sIpl6Z182geYvH/ia2PQc0rrzNU7Vamr/eJtsvPIcPZmgPZEBnA2gSK6NMT7hMFQxXc+COFwXQSl
IjbgOLFpskpzB7VxRTBgejDaXloxErFXbXB6iW6lzgEvAc3UC/ofT8bbHuO3zuqPtsQSpBD9di5E
SoPsNVzemGYHW07f5F+x51orpt7JFH3TdRA9YKi6IsAHeU4SMyXyqny5OTmD4D4QuH2L70Gug8KP
EfgZTLVpqIspO0lHgPUoka3QOkJdLfae/9JA0F4yoSSCVizy+GgYnlOzxT2T3zn4BHyElRmWYXpp
H9Y/bMuLtDogyIEXDpakEgPK4X/cN8fpz2mqVFPoQ9KzDV2n4C7vezTVpL51+Q9OYhDsJzdNHoCD
1dZHVvlbcIlImte7nlB1GlvLlOtNrrig2iEdkRSXxWe12gL+uZn3beTXJKyLL2XVWktyiLQpT2ZS
acdY+hBDKPTbKI3lnGmkbqkZ0vNzljwVeqzu2DYFowo+JlUOObab9WRJybC1PPKZw+jTqdJSvgJl
kkfzZ0C0KtGzMuEmUtwLVfxcg6qqRVvrF/Ij966TDgS7Fl8kKu79n11MIRwEqFWa/uBSFcEzoyKP
zcm2MqMTNmZ+0jlUXg40F4MASpuL0mysYVF6UskJpv0U/1pjDV1TTbzNBmQie59Rm7PMtO9lr0uo
y2I7exjxWz7awqv0SygQ9M9233J8UONkCWI4+XsqZA+b/A/C90ezuqLMsxd13sZwEnp/1EHcVd3x
B+T+1DXLzCg1G/qN87L2eDpEmmlXoibVWHmJEmq7CetdeclLA1qjZIK3aJmp13MHW7SLS/6t4duD
b1kaEYyxVgDSWQiStGfQaSEr34HXdZO3pQBG7UoX2f1546ol0SQBwpy5gj/z3t+HgpEu9Ug1H7y1
q9rtIEk9tStOP0ZNGF1YneXk90zEoZWstEBPh7hsnw8RZKr+yBhatYoIIbwR1IMXY+cQAYitatMH
XF9SRjNYfDeSLUsar3TVModh4uc1V72v+/T2hN3eIndQui0HxE02LQuvhOmtsKQ29160Gew73hn1
Hhm+7IF4ujIANzahdOxSADMVfDAUY+zyiJnxBonl/UMeMlnELLvT/Uuz9tzyFVsYwPuJAGs6Pf8n
0UodvR1f79G40TNyHPu+X1tkYJNoBNu3u4XgnbaAVejyUl86SovR9Fv5/25NJzgluG84E9gY0cuo
x/SXtG36QfhP7UJvTTD6eyPyHDla0V8jO/jveyaRUZwFNDVVFTjxVePsXeGugJsfI42JlrqeVQPk
VhoMShWmiJbMALlLVSWYf/yeNjACg9PgCvqaKQ8/ziSjWnB0LXD1AkMGfsxvpmaZ/sfuRF5PvTc+
VEhv888mwNaqxAnNDPAFD9eb49bDXEuQb08EzHkWx+YCet8BZHUBhtMnIwfrD9lbxQe//elT5E7W
BpBrOY9PMYMNVJk4RPuODGr+aWuqaOrX/jiXWKqbOjkPTkCVUDaNk001K/gLyEw/IFg288OSXBFk
qhuNaEB52p2K7d5PMUKbhKz6rGGiGeKx3YTa02kdpVl3116/YTD+S1G4JWe9ivw+vq1Lid7b1gnK
KrT+zWFL9a8xBx3neb4Xhc9ZcctOYZvvt9YsYy0ALpqOG0T8RdMbAbI/85EN7cLdHCRMoLMud/x8
sEyLAV4v504JEJ5uUPomBnlTEbsNN7kCf1lxG2KjzE0fUEF/ZR7Q0pl342yVhQ+R9ZESZ9T3HfM/
geeXPA9z5iWp+VgU+R/xko/O/WDJ5AmayxpfN0PpK7q5X8blmPOVO3hikenT56nqXIsNvUYYytjh
iCEZYs8uetZLfwFaA/1t5JQKuonoH+sgK7hKxTSFh5ql3dYb1qcna8rB5BnhZz9RawBdblTbxf7/
9q8WY1jwRup/nfSoSkQo8zFNIO2jeuPvhYL+t4X7caCOCwQTNGgQQA/zDmRbgwRncMA6I/hzynSs
gy/QgutsYGFm/Si5q9pnfmnZV49J7uFXdWp7essFo6eo/2kF8rvPxe7SqcXxnUyxt2cnhoam5YrP
MFpA3GLGPZ5rqwlfapwbHkTS2NiCUvh92na3m/4mt1P/xYhRFsWhqnTesa6bzUPe/wBl1ty9Rfwf
nrRolcTjDOT+FwzhjUXIluQvcYzvULSF+BqfCer3C6d8wQoEyv5MVt17FUEb3buw8e6LLEYjVehQ
Lmpy3y5wtBJfzuXMku3Y9U9kKMesNKJKEZvdAccVVg3Os+/CFJeRUOsD1RJhsMmaqWWX1JQMopr5
k5dYouL3lApAY62VmAFsfojqYppF2CCqa/ialbPwW/wCFAlBY9feJ4xOGyCg6RSR4YAunO6inM6z
SwWZdi/Nn7AqtMYSUeH/rv2tmX/LD4CGXeZ/+YdAgAPr9ei/EfG6XTfVwnvwbyRtDz5A0eV2hbBW
KWnysAnFeHTDKlppraBfHBugHN7wLwu+U/K8x/Js/zyp7OQjx3M3IAu7axakQcPJMUcqAdKBw0v6
tPMGtZrkQ+aDgHSvdx0bK2HaHv0tDtYQP2kF0uOThTbA5ANmMbAOOxvHmCTWrAT1DFD93E5BieF9
dXT3Oi7Uch/WpBMVAgnr3yJRAvQRPUZ+ckyGAXkmzPn5oOmD0xBLTnqWPE5Vt784ijHMiCF5iom9
dWoOQR1ZHoTU7hOeEQ2erXxjUmtI1W6B7cbSBa/eASM9UsdGGNd1cjZSRJZcMgJIIds0wE9vmpip
P+KTLCVSALl6mrr1HNCAS/LVAjyGXKYRqrrNi3fjxzXCBFJ7+8e0neVdSyoZYkc9tcZraYv/oM/O
PZV4jubWQyjvtriDba7RoMZtvVcF5+pxd7DOZx8F3ZfGa8rfs+Ezx8VA+dXvFIOjImBZsgQxd//W
xbbmIwuFLGLuNdkcv5+3QIkc955t6SCPx3gwOAJ7idakT7yg18oERqQ6DPcCDTcbEjjy52d9tn4P
+ISXLDVpmXIaA0o0Y476jtV4R4QM+/FfIrbpptHAtTKpnTNVllLGGNoW0/kXhGccoShL6OJVFPzY
gkZepZ2BLlf168ofiLqRXCn1kM3RV3RELNz5dNAWbWRWNszwe7uh3F6bc0YciqO7eJ+GD0AbO179
e9x42P0zL0MgeP/qtj0lvyRdaPmSeypNDd3TyOGC1aUzDN81cpNQ+/TcCXYF9RIqcTtc4LSVjrjS
7GUUjt/jYFUN7KdqfK36/17wgGZ5j1pNtgn1ghYIUXoC/hot68YJ3ssYH8M2B2fZJjIUbKZXw/wz
i8h9GBR/5gA5JTjSqC5jrL0uhiwswc6/1f7mbDkE+/VIvMgGF9Q2vM3qsLZyF3OpMpLE40917OTU
5Pi9xK0aLGbR4MPnaGvv4o+CMMNzm0l5X+pB/gjdW9950BSBxrPCioNatBBIIstQxu0wjqP1SHRR
4H9pMtBGMhZhj6uSw8fgKAIR8UnJ8rjHnmu6zVbJ7XWocd2+E+Xx6ibLkN2y34LS0Q==
`protect end_protected

