

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
rKWwB0sGGUajpurVPwhHzgsZATzg6CI2fy5teGZgwWn6RJSxvVrm7X6KC1NlYW5YtUDp2ese/Vrm
bw3OqIV60Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BRuqFpGYGOGwcHOC9ByqxsqWUs+0okjDxEXI9LjsXxEyuWJLFUE7YYzNDASAihgXdiZINIm5es9z
yyLJWg7azDkuzQk8G9FmmXCb4GMcSNpaTGa1FVepRSL9Yvq1uMN0rfkU8OoTCb0JTco3mn42K2KI
S1jw6CGiZKnXjxgHNBU=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
X3xfyzvjrmPkaI9JdFIRWVWKvQVaKvW3xkPmxmWB+Bg2oVsfAsBqh2i46hM/Bcj4vTlgRohMAtTw
mZrr7U78E4bYF8iEtFKLdIJEd7hVOOlmDwsFBDzxg0k47kX9A3ruJ30LrjKdxboHAuMIaT/XR/sU
upe6flMZr8VBlv8re7jyziDyWZOLqFpjufskTfv4OQj1KszofT4kUnArUhuQ6UVlh5i6v/pQEzIn
QBP9XWEv/eQfQZl33K/QbbRAZIttPtuWp1T04bWkTuCPPKG+pDFGGGHJZvQDtAaxZSkHqZAvfqlI
CAW2rOiYEadE7tUwZCBmG03wqqm+cZJmCFoaew==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AUXv88ADQriH8V/F9F2bxLErHxhqOWkmnlCs9b253d+OgRvIOLCtaWRA9DjnqkOKIf1wnvs/R6pY
dJJExfXVZOjD4nIH7uFh77R1TOSQouJzgmqD+K5HYb0maU6PAGIafeBzcUv5XN4HOOPvm67+oI2c
ikEGUjjanBNxts7eGBk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UZCooc8nZi2nNWJ83Gcm6qAONngeeaBUnqNHZdi1nOU1iRX6MguqeK1oMSUjP/9bRjlw7Tp3sNmB
PWJn2GGi3l8Qe6b7auDrjGMr0IkAvVTyrVlPQlMaseSN4e4IeWhVyNWjm//n/TOKlr4NMKKu7xlw
UYk+ejL3Bl9bd8/cGgsVR5ZkQQavRAFBo8L2IT7ML5f1IYG78bF0KQzrmL9GYFMnToP9B7kVR7Du
Yb7rcfK2Zazdh5MpYg9XUjLic80aZcb4+8dYBu7XgEp/Ar3GApiNMnYJUmVK0q0n9Er1Tqahdfht
jdB1SKLd/YF5uaRclGtmIoZjAK3M+1SEWOps9w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12224)
`protect data_block
GuzdIvroURUQ8GInfYB+EofOwlQUPYcIBR/tcCGDvEWjqP7NxLKY1DNQFsEuQYuhNdg4eXvtkz1O
0kZb8TIvHb4MciPKsnK1f8jyN6PG7Eevc79EVK1efEeQ2B1XQhtlpCxl6HBvRJIyNSGQvgrKQ5W2
pUa6abRkK0o1nNnwhRB0qpPAIIyaRIwAXrMc5dFzzsVpacu6APHUhg3qY63pxg1au61Qw6GPmHkb
1G5ReKHvvzZ6qR/aTGpvVU4JV8U+UfbUfgshD8BTq1OBVtlJr8fBVdBoFcMR0JgBcgdbqZ8EBCMr
s4GYmmP4rDj1bXF+fzTjIrE2ucBZ1x+K/p4/0r/kkg2P1DXU8TnDGUj77bOGh6r/BbA8X9n9bOxA
m4WmzzfWKZJme9wImWiwZaGg1N17tWEGIv2mcSRnnFJCiyu6KOSNoa9d/ji5WVKG/vXwv6PsMuvZ
cW3x7X+FhacaNaJ1j1efncEwZ7GbIHTXQAIr87gt73dVcZLTUaKprD8ZsExRiw9ysVZvpNlkRFgT
/+l8wMxVKlPbhDGtFpgbauhj4QNYY1DO4RRgyD76fuOXNsmz/QfbnMINMhU7s/4/69pfvdKW3xZH
aW4JtoR4csTzvDYcn63yFybj7+QgpOIPFNvYh7DprtZBKbyT0cxoyr2uyD4YQC+t5eyLtKkjOqQY
BliRGogiTtVxPpzqiUKCBQLKGSwXg2tVAU9lOLbmBFxN7/TK9oIFtIg0iGw+iG4e+Ol1x8ETO80s
k4TpKfoPjPLWbDPxJWIhLN6TKOZeJec43+8NZ9s9L8U0XYAuEx8tSOLr3G1HMgPxd3BkVEmvdJRA
z9Cy0q4FpE0DOJcdkM/wgH8ZYFwNNxLtuzSgusYGPTE/EA6lWeFyyOsENyA/nIDxu5WS3AeGpWYO
ED82dX+KrHl9kEtXFraggKLddTaBqcAKxNRrNmUzzxTI6Fk/ACc1ZnurOadLlgNe4X1UgkEQJig2
a+gAW38L1hxFjnd3zlcMuvjwibrcibY6qLfcGtLx6eehBhK+2xDZ6jypKUc1o39E9+dBSh5I8q7F
FUlp1YZvRUVOPYF6eFrHxlXVNUXttuzFA1WHrFi7wTIigYNuMrkn0rrw6/nkA2fQUo7/JObih+cJ
EDXa19Nzueygh+x1EKNtL0QM94BaH+QdXMhAzmCfFp9GC8ZMvKea8B75pJxMzlLsmeoGUHjx84vj
ei2M6xivsoPB2waYTC8MmfonxUSNpRVsHiz4J6mJPS5T9YcNpxIfoLWRLl753XQ0g5tcHXkBDjXW
PtsYD4lvYtB7ZZS9v0lTezDfu2OWZPkjciZRhqfUvWaR2cQ7ydZjhVap38+gBSqZDGhoDqVtGRs2
+kaVAe98ejr98Z35nVjJVI7wJsCHGmIZXO3nzYtTRaivwS8K7TGK0dSRtB4fynug4/I2B2RqB5H3
UmTNxZ+pOcvvHpXaQZOrbFGQxCtSpXRfV+DZRDOW9nvBXPwglYMqOTU3k0NAR1LrMifiryD8VbPg
j0CIjQHVYlt1GS5J+ZDADh3kpdir3i8ktr7qtM5BRbtB0nhnh1glIZECykbm9bq98dR5mknWwAOA
2zuoW1koH5Nxu2AxBaXsm/NvyrHhzrE8ucJvhAdVYSD96aC/F8qFQV0h6zbIPc4QCDQpetDryYCM
F/EJO67mzj1HuzCITRlijphJ8/N5q4U5JbsJG20mhqTVN9AmBGPYbidOMrH7OXyKhe26yqpiHyef
Rup5rRbYbDbqdyO8WtOUXioH8Bv31QPBKu6TGOCxu/+L82mKUz3S4SUoOxDL7sNfyQTvCGAxMPJe
NJAyPQXZ+cWjo5TsigHmhzhAQEcQL6mYYdbSOIgjFb/8oxS28GB+RW7qAmy+2PN2AhgZ8K1zBk5g
7ccUkgkDFQF0QNTsr3P6XFwbVDi9iyFbKTGXcVIjoxuczl2DuPszZS2PI0+4GO2PLNi4OC7yIK9Y
k8p2DtkI+nm34mcQ89AO6iULjDtkecrCN3G2XxJUEiyNS3HIvjKK7sSE6b4rmSnNLECwn0FNxOyq
yh7rrPJPYN1+S7/1q+ALUymOJ3gbkNg/u/02mlDK7RwfpcJ2DcAa83H1xFCCeyRWs5gCydXri7t7
xpMgDIdq03D4t2L9+QjnKuUdJstjvi65kdC0zewAu8Tv7Z4d5HKYmwae/1JnbyIQw1INO2PtDzLs
cOJsxxUE9zNNEkBausj/r+Gao/IjOZqMBdLpfRD+Bv9yADgxapcRf201BmykaH9WzHMNHgVxJbMw
gDSEKnplHon71ze9aarHjbLz++S/VXox7EUDuY0KKnKSbhLD5PZDs9Scabsz5UIdUuQouvuGOLK4
lNbnAytnCW4UADf4csoiA7TXM7NjI2B5E/xxvlns3VRbSB1LZ288bXIncC52EVTybkufPruprm0+
hbgdJHBMK65BD9qqqAHm+Qvr2K75RGtLXSMXwgdTlTLWi4GKB+z/tXqHvbGYGSkwsRUjj5h4pVCy
nku0Xvlvpan5//Zg3q+TXezvtab57WkyMbVSpi6EK5pBMGMUv6bqn3IvrQCRUj1JhHH1O64DFj7j
Cx8BEItx+YPGSNufsdRu51nXe1SwBQi30/dFWcjm8sIzFRpCVqZo7cd1PXOPMWvlKdc5Q8FEEi3n
7KRWlNn2Z1/6nyJFZ/q1AW6AezxY8N0foEfHBCmXNlX6gVBUYjyQUG2sGIFWrsvpDQOJ0orOc6zm
nvAPvCEfnT//CtY6BBdN2AlXhxUUBGM67N2ubHkgvn4MK2Q6LRd5JaxgYtKHOf682Hfy5JYVyAjd
tI/4N5ygdyK9oZYrw1vJ1gVjw/K0R/+MSfDByKPW+yBKqaHbVQ+jBhzR8n1ENvI+/GiU9WCi9LS1
7MKShM1wPrOzTg8FJk0rgg5iPAy/nxx8oSfeHctCJA2SGTV/S1RFbMZdfGkIZQbKA41TJCVEValc
ZR0/OCGNqHQzOHgMHbwCURvPssbKymx7i+oFFv5SiGbJETD81IpvFJJzuUxq9pOc7ZEU/aLinHrY
z3XZsOPSeDWHrH9MJ6TsdxbDadwHeicNnaSE5xEUcMLFnxv2irtttGYyqaU5JwP4zoTVtqMHgmZg
Yamly9Simo920ajKOAt14YWzjjeyuU98lyXqYQQvcsMbcNntf7sHM6H8FRdZYup/xxLeRxafKM3N
KDqniU3tOkozbp0qnwuFRGM4tx0y4lXdHgT/+K3LYbacVtsF+98NCm7ZHUeKNheRkRsNFnTqPgJ5
vsu2Aw2+0A8wEdK9kwpfMwdAHLaDP4ZszIJNeLZyzKI78/6uSbKSKQVPlltWP0ejfnKsXKph1jLA
iiT0+VI8EZBETq1GAg7zRz3iQs0+yxO452R9P4BGLcbChwf3hw2ogqWtfkEgahbjdACMrQE6+IFc
5yLHpyLi8IkZN5gnZDxqlDPRMoNEQVpOHaHKXpFa3uakx19xLUCdX+5hgTFSMMjSW2/sjuwF7hc7
J91l5ettqInICRyYWHEU9kU8S/QbUMXuDE51WcR2ZqFbXAq+WJ0OXTo8UVrpV9TW1kbFrFsxWhit
y/EK0+f6ywq5QpWbZM5NTCebd/nU0YMG1wU1hqFpbNMdRJmBQ2CGz3KbsazSFtEPIq+S/92N5KpB
k5k9B0Tt4nRr/cqafNfGrBnF07m5poFJuJ9sAI350O6KdqmQiL3BAorsG6Mbgg2vcV8bXNpDulKx
YlxjaQLxz2nVdJRsLlfZ2XMOTOFcITeaVOfDVXkxebObIU4WywEJ/dz64mhKWBoDy59Z226Ztx37
eCDkQg7E9EiYshtw8rhqCEWvIksuhAPp21f9ogJL0akArxoTRW+5zgVejWZtDwaVLd4JqfdmDUe0
blROxbn7QvfL+7TPvhav9xs3kBztZj9vt4sGBH+HxNrbWrCnSLqW3AsmQlFawOFtiqMcObKRn1ep
BHDPg+X0X+DGswK6eEB5gDctF2/Yi9mIAS00yNRqa8pELYQ0WSZ2MxRxL83ucK3D7jA3fnHWYuxq
1BOxX36g4JV7+ESXPtxB4SV9ZhpZkKTB+62vMx85ZF72aGnq5HMrKgCOZmsGSB78YI3PlMEsZr+u
byd1UNbpjRMO8iGuCiPxxCtW0wpZse+30ki3ks3EJaZzzOQy75T2QvuvhV3PZEZkUEjZkxv5Vz4h
ado8oNu+NmIs9fvIYRvYkpyF9juQscntgx5W64IfMZN652tFZTPM4yZFt0U5ZR0qOgENQPcrl78+
RdGWsRcfnj9zcK+8ag3mRwpemP7GC9dRh7SiL6xgz0Z91x0cK3IuKy73oZFfJiUaT5sfbg76/i7h
syj46dN8zH51NXmMqPg4CX57J0QHLEcp2Ueq2fJiOBLizkh6jbpooCrnWzTwtGeGRwgA383X0dfk
7GyF6j6RsByS5gLv4EiTukTNrPpPgr0U1ngft99AYyBG+ixfYsFkM/U2o5ps701VeKH7aCiGOUBr
MZlM6l76nVbXxv0etxBkrZ5u+HQVzd+nuKFmOARFp08Iz1NQap0cSrBPdfifjnr98Ey7WrrGP3KJ
FmakrtXf3lx+z1Y4CXN2kLJN8N6ySX0cuc94uLBnFO/ayrPAF6+/ZzmKiwtdB+nEl4NI8kIombCi
CR1RuyLdHHDv4MitDm7v78TFfAP9TMQkhQ5axnT6wlShTpKD92JYpfS2a4HFToXASQjtur1J9XMx
Lc8JgyTvRZSZy/Lad2bWC7jkm/OC+cYomZ0eW4TVoDT11RS9whAytwT7LSX5O2F1wD7obv0P5V5o
PAHtOhvYrsc/beAqVtdk7XWy4u84P83QC8g4GgAl12eNAxcL+ZMbipaFnykBDT/qPE1Xb79nw9rc
X/NFyTW0nanbWORldTNTu6BzIhDyXzxvf23QMFs6zAeZuAH0djFTe+CLeR+zEu0obcR3yU6g2mcS
SV3plQeHYunxH/oph41wuw3/5ACADDMoBi2SCiaUhUJML/iXV4m2xI6r2sm7ZqyX4p58uzWLPeLx
JRXJL5bJTT2lKj6d2DRfMGsBz4RLcWn46yMP4XW/HqS77OVSm4CCUH3OTwh3Mahdn57yyD4PY7Xo
LJHXg2fPd3tLZrUa4ZsqKouZjgKLvbBfQ80eAPn+601ykW5bphjJAlgrYu7YtmkA4ZzYISCrXIoY
H0wYeYYqcx7P+h4tGYBeiVqtG/g7I8eu/whbMHWkoCZR1fALzGw6mvY4C1KRR29xH0cuubiMCH8A
Q2HfgxnFYpMS0rv5YxF1g+0MOslhAGR+jZ3A4qgNEBS1R3vUwTvdDkGAdI/ohyG4/2yepdjcByaF
JREop6fPF4+GkZF9KMSTXUd6Lq0sRriSNAwtankf94Eh0jFmhTlCitGFYBo0upcEYz9pZYgjK+pH
gcJokwNQCzdKjtXpegRuhl6m7M5zdZn9VCyFqUCPIBcV0yKS+RVw5+gTIZNc7Mwvf9axrn9/7pMC
Q20AhflGgpU0bPq+MeVS1ZU8SAzIM01f3t35TircVqDDMyxkRGH61BJ/nOsyOWvV6Hhow90TwjXz
6Pd/B9g5vg+Y+nxLIZ8cqEezeBn4vSPUfu8AfRq0FehpJUbE8cq8qVyiPTQoBzem4OibE8Hp0+4b
ErsxxV/R4i/6b/poxZDNG+RKbW0pknlzzfV+g106FqSHOudcjqdfUVK2yXE8Mob5zx7vrv76hXuy
6TMQ2yOk1pxSZ36iHkCPqsEmL4nc3ogCZCs3gMRhBqgYGk2M1CbBu6I2IOLV5UN6MfmBYtQAOzgh
oY/GZYF2eEXnFQ4/1H4skt5F1bIIsjp/Ev0ZV202wYXxsDZyJpRSFfv/mpiEYsFkOsHd5v1EZL9I
yoxrxKA+7HmEqWL2RoR+6UQR52mLLyDxQMr8lyyoZAszUJiU4TBpHWOkOUhViX5++aOfKLtK/QwT
Nnd2i0NW/fjbUIbJvETb/4j6Xr9/mI33WNh7NmoQ6LVDeRSyO3nr2xm2Y2oIjNzktqwpv7AvGC1T
HifSLoCrTmE8ReU7ncTe3saOommrAZjefY8TvLjjyFdBQoMKmncmk3kn6LQNHHnvZ5Pj8Z/FEHe2
x+2FHqS2EYR3QE9lMMWW06G0a94wvo7ABurnXks2wzE/cL2wkKW2gHWRIxEk/7jXI8dKQnWe+fXZ
AgyDIjPz/50Act/ggJNDdygSJXHsYZeXP0y4b15bhbComgDYctpCaisA+tAxgBDfarLPXAjUPOm/
tOQqx47aarcV/8Jon2qfrehHKvQrkfkbTiXljFplDBDm6zVyfvLVFK4zaJgiMI5ziQvOU9iYqvaP
3aFjZ/DBq7O9CKEhjyrOYXUoSXTVtU1BxECYBfQFZ02cuVO4NPLwZISFJvXt2x20hubS57Q57g39
P31xBC8ndf6OxDJt0C6xgd62M6VeiKkOihjc4ROR+Jtfnd2Bd2pwogw8XdbrOXngmMfsC28V0u/o
PgR72kxWTbHPlstRLDxQnHI7CGok9eku45/Ho7C6cax0WQ2Wc6SnfWjLaz4dtQ4GexlnUAvaPFTE
bGl0Xy4NjS3ZUPXcLXJ+/EAONThjQ74BL5cgyfpJwRISDpzEKQ3jfAdCRImxK168D1TjHxLZxrVf
eZoWavVC6F0YOlVZzoT0vhS3Jog8EY3X1cw/dyr6r2R2vdQA5knUsEcRa7dAhtN8u+qaQgPljez8
D0KOxldkXG0jIAW3Vv8D11utKDr+rzsDJ6xPcK0L6M6slbxgmAZjL6ob2nd0ud/eECO+EXTwCrTN
RFPxEYkTuk+mU+x1aOFeFUqmJ5VqWAoXA/2oFW+DxxyrB2Kq7tylwWqKD2VnTUyLsyaUPsmpCkmC
Mgmpn2yxLTn4Uf/wGePfm4d2xcI6k6TOxentwEgMO80O3ACbA9KBXlvdwof1ry3cxSDFflNCxG5v
pqZFx597+UYIU5/S6xVyjSyuXBCRRLlZh5RbPbk70Ti9qJp2LgAshq4CYGQ0R9XCIRBdfiyrVbdY
DfRqwCeRVxLyxS8RZp1onUf712+BWz9wl7FS7LhLqXeBqigHb7WrqHVvIqJlL1vodUvkDpDfQH4+
9qEmHOsQqavbcYcilhBE6zMEHAS7a/7lI9hlTzBA72uv+S0dxyXe/yW0BuRXXCkW0tgiss3uwz3+
VT6f1Zk6fGSCmaEtK4fi8xQtJEslxd7gNa56D+8N7ChPMr8SzzqimMHMWfWYuo8E1Npu4bcGEWK5
5t0crpTT50iVC7Z68WSuoQ+8PmkX7biNva4gXyW4F6hpv6nqtraHDLq07jXImk8KXndxtILUnAD1
rC5o4jM7VBYHf9YYK4YWqdx6z1F+Ms3RG/GpiCdNXfcHWOyDPkR6BCZk4u7a7aaHvWv+wHONbIja
9TeqFLbyoFsuasqXA9YPaqBSCukZiaOsl9RZu3VlhCmnWgkYB5dTrVXJh7YFAAAG/5Z7+rcfQpdP
Beczo9LWGS/vGDTD9vbUHDfllsHokpIwThRM+EYt1tRhDMJ6rny+aaGMIy5dvzP7o4p2R/6iUUkg
klNXRy2kkIAvZPretcuDmMSrn1P0P1EngZyZyWjwOPUkU6tMnc7bI8wa4bAHIKmWAEOfHs24FJys
YsjfFdvMRuuciJFIvlvmS3r4WkzYrvQaN3qIECuG/+c99r+LbS+o7ttOJ1Z2+EmvwDpikuuFpsot
cPJY8LTX4v7XDmYud4U8XXMTKsawEtNR+JHWeeHMU9SCSEDU2cmLeYKRMudiFrsI9vm5+Ia7as+G
u4quPzkbu9kGBXUcVqHDO3EnZcLIrlqb4Vq8wHzPkAKR9RB4x3BakA0BKaQf5TB+HcPQ8QHZuIa0
vU5uU4pLjJIYR4GsevZEPLB7ACR19VlsdA+His7n6XTKGiGHhEr0IvEc9NjkdproGXWGagb7TbfO
Otc9y9x3XpnksTa5q5WOO/82VIp+iptMucqxrLY2aB+HJc/ytAv/mtFHckak1wHGAjQXJQXjzLQw
Kd+6QY+n9DbLy6YHWXC9VzlQTtd1RVmKpAP5mERa4etrzhHzordFGvjAbsMRCF4CQ9t1D9HvHEF8
38jq3+a4WmZVtRVLMNxcUuPkwi2/E18vQM5+KvhGN+jwdJ75E3Hs2bPgiSJlyNPsX/wDeetAU4M6
cojZBkfgOFo0qxl0tHa52W+6BnmOYI47R5Sfc2ERqn2bgb4js4RMIQibkllaUEUKZjKBG4zBnkHn
xyOc8sTiXN7kD7n9hy+fx2a+U8qs3C6zVqv8SokU5yXo8wPl5snuc6WALs0/Bo6tpt6D1ZSdY4E0
gcrhebk3N5jrVE4ST5aVmzO/2E79T+Ne3dtBhVfF0suNBFngSWBvDVvi8rMltyGdBch0b92wKPzB
w4Qup7RYwArtrLYLBWfuWa2M+4VUzCJQLZQnxIc54HjR8IFNEa556RhEDAU7UyG2FlBBUY1evUCj
jHa3qxQ8xpdQJauJLnELFsIp+01EiFdccU5jMu4VD3Ua18Pd+uz34CbIofQ0zcmYCAE+9ll6NJxG
2n1NSx8F9qq4/E9JxjTBHagBnGwCSGibzvM/gAl0Z50XFcZ3YOQQobG80Q/hLrw3n1q1x890ADyF
CyT2zBsLu3WeG9kHkTgIEcciW8JWP1B4zq9uXdGuXOuuMl2pCx65qC8F5DvYlvVt2pXHwohF39Bn
d3EyxdbUxSoDopOUHNzQaMPaLoa9KsdHcu8Fqp3MsJA2u3j1x41u1de8bccFCuABV4uNYN2iUIM8
spgt0gWhbVigbeWod2I4lzuXABtYxcIk6qJXnxGpdmOiwrfbReNxPsTJmMTrYwRbc6HfCzXoi4zs
IgdKfJlDlB1Dkluy/i4b+oYJZ/LhoODt7KfeQirbAskbIA3ldW3XGXvSMX7G2BjwqtuQHjRHRT3k
KD5i7r6xEPKCGb9rupevcVv5V28RU9m7wyYP62EZN5mpiNLYkk9Fb/Tf/plFOrUS1+kwLF+s/mEw
x5vqUh9L0PrNZ8lIDWWBA+K9QG1FYUC8QlHj3mP2+LUs+cNWoOACWJcYiZbQLZCmx212aTty9TSh
EV1s2gib70kQ+TArsGvlqFFLp1cLvyjv+9maqtfXAdZgJYKqnZ3JuXjaLmPs8DC51fHU3y0kddII
sNr5h2f4fasfUJPlv2e3Y04UbU6g28xbVE39irzumlt4VUARGNSvdVc3jcHvhXkjTxQleyP5+SdM
1ttDmh+FwJ/8v1P3YPEejSvSGH2JFzM4yuVh1BVLDcYMjFjBUBlIAmdnyy4OJvS2rR6q5CLHJcEC
hgpZJRklq9aI1K01UFldD54HrtUgebT++3UGUaIExK6ksdXR1lqFqLXhYWsaZwCAc7MWOEhmAq8v
s5bRDGV4yTQCRoGYM71BYyMrl0hm5vQE6IR9oriA2QYDeYkuAB2f/mvdyggK1s1OKOxrZ4T+kq5H
KopjoRpgtIgTEHbrAIGDZuZ415cfehDSbK2pd7OqXDlVEq01I6u3wnYwmN+kytJfxKGMl2brw29D
z24P3jB3gk/MihdjjRFMy4xvTkALsLB+eQoeWJoE2KLU/9/M9AVZytvVS30WX2s9dSBIiTBkuf6Y
XECnOQSgb52ScaSJ8dcvoQYx5Go4fRfUoSobtR+Pz0KmEQR5SBKOtrHJP9kzoBX4y1jeyv4aBgb9
3iZhMZMZ6hGtXsW4ojs9G6FRWNPd6l1dNe4O+OOGiI5JwUTnfvkyY6iSPgKQfTe5St01lyCBMwyi
GmgdkqeLz2KL1wsLwyEdm1BjTxt+KBkp/0JRp0JJty97J8zGyE1Ilo0N82/xA3B9ucPxy6GzSVTj
Qcy9DaXgrCyb4GUH05UnrzywEfdBjCm006fnyJNAqGn+TpXCHAn5V4ZhntHjnwqS54xsyunToTdo
muQ1a5GjXWm9kzAXKll5L40BaKOzwIVl2FwHraYJthuIygGCf+YH+YxutQAhCEbGotP0BFvLL2p1
uOwAwX2AXuxgmfenmJfkD1SHLCmlg65oNAbn+9Fxaow9RX1bXQY/tgH4Hu46wNVFaCq5+BJiNb6j
akmlAwBxuwyWjvkAGsJx32WqdXHFamG2vxFEAgZUoziYEk9Pjg1uqux+qQ6vod/6l7QMuy9RBBIm
xH1J8UNpeWfuDCl4n6dvnQeaTqB8HuD5J1voo1OpWI/JopDznBqgpwg7Eh9zyooqUJ39Vo7unAMT
rCtCDTkwQWH3e2DvMIRjkzeePA6SCI8LyhV1YZiIJY+emfFu7lxs/nPtNdDDwT5fNX64IH5c6LKN
PzuD/UyqrkJPF98c8SQ08bK2WjcVqp0hnicE7xfZAxSgwUFRjZ9HUPzwwMVd7iQb7ij2uVyyaO5Z
PK4czNnTH5kOAvdM60Lul7xiHMQ9O5go4ZkOim/E3ju6Z+ezA/4sERSYEBNrFH9+a9mD0D0JS48X
0MZgnAfcnJ9nqMIfRtVzixtZClNwvBY8qq6K6WB2ohr/PgAbjvc70rg0TJ8RfqqGP0t5dQ0Dg/hQ
8ATnXrlJBXx1E1YfkE2lquiPl5mkXvHq67PYH6jEf7fSCxOSaVEZAiTAZa8OXfbmnbesuwLms5YM
J74E6IxsuqEVKJdSEEQFgXF7s8RqK42ZvEHW3oEWP8sX+46hE9uiymuoptdFAS0GD7iebw58cAZT
p+3hpxrvxgyjZSr4L3ZGDJisDr4eO4iUJ6kpkpY4lAsSVMvsyKUbgRVJL+PjLfVHKIgi8a/VV75j
hSwTTdbw8C/FEjiyuflozpjii8C5630GrNmZjiaMQrEPWgckVP/iK20fvFmVB5JpOs7FSyAactUM
7xUZe7L6RHSkcR3KYRt0ofUb096Nsg79f9RBA1r4rNeeEO1qN6Kdg+KUlubeIgXh2CLzW+9qvJKw
WrOapuJuTGCf3pbmqYIFCN2SF2iwyaEG9QcoGkVCcYTjeXYE6k8mMfsCDSKXdEcMQz1kb5YFyC/7
l5q3nvGRautxqbDSQ3lA28Qj9RC1e2JnkNxjpMXjksppoAmvf1/95bzqDFw7e5kDs0H/MRfBsesp
LR6Rd5pxfWyd3NglX0KheLbWxaX98PQLPYAwtPDR1gQJUv5FjCeKkchkglRh1BIW5Rhg0Uh6tcFv
fn8h+NR5xKVUWcMoGlA5EBgGNDJQecPeNuQJZlpFzhTBpcux2dPEh4XN69AIoRCDa9CgG81LAaHB
XujnTSDXFgfjfeA7kkeiV4pr752tiCvjsBgZdPSf+s61Vr+xQaXhmAfMlQCcYXxBVXzQzWbWlnFE
2jJAVhi2OFO2BQ/3QeR69amW3rRXwY2ckW2AvR9oFZ7WlVK4agAU/5Ui7qdSLKyFhrPWZAA4QF+e
HZbvlu0slOPr34vs09qmysKjpL+qwW2poU2OK2ybE1ZAxSro2v2z9tVxacSfBaKckL+HldqTI7Qo
mr63aUMnYAhJgvHnVflmQD7mKOwI5lxC9IlRo2fnIahj8ObEZe1m5NzpYouASC46hMpuL2kX34/V
rJAaUsxXamuRaHduQ01jtFO2IQb7wnlw3Trhvjzhfz7hNRRpnJ4JsN5BPFQvCx3BbeJ4ecVMXfgm
ImCukua2cicYrPNKf9PVNRDTNAov38V3GxpzqbtTFwGHeLx1YMqJIBJ6eIBQJ6wH0TblYjWUE5qg
bDpsWQLGip4ecbCRkeuQRKI/g3dlLNefmes1YqkcXigoGMgA7FUM3GtJ5ISd4MrLncDMUJwJPO60
5y/UO4NthmcEq82looJWOOr/OIzR3jxhgYSLMC9CADC/vYbix5R5FA3gFJA4kkAE6890AADHKQ1w
LXIFxNEJoPD9mJKkwAeWxWUYsDB21pRPo1BrOCyboRV7+vF6PapDRcPj/Szvv7CnIzCK1O4iPJJH
Evss2pTfVdKLadr3bgKYUbvn+O4YJyE7d4WtAe57lf5c2847BXH8+DhdWuSaKH3OE0jZ3cFZSRJT
K+yxam1jql8uzX6S8H22BoKpZRfxkAsoeYCGje1snSCpzcEu6mdtaXd3jMAwVmhbmwnSzcxhp7Es
q4kVQFSaUdM2r2JEY5ISu1Ycrk3ZjR6Ni2jlU2nf0G+YgG+Ry9Dqg7dr1rXjt0JkGbsE8IA6vBHL
1rqJAcHgMeDpagE+lZQEiTNQy7WwK6tiNVeM5isPTEi98Ht8XKaABFKKwhu/BoO08RcZCZydO25p
kVWArAx30mFCvrffkJg8JRI0mbfQLvawk4LWARG39PB4D38gVilf1y17kxhHWOplm41JNWzYiEJl
pODqHXmquucl9gYmeVTbcUM01TSG+l9EAZzgnCuvB9E8rbEYSde9szwTqCsSfQhBf53kV5jqUIzg
8Wn7Z3Z9NhTPOePdq2/NQNOdgvEeYuAwHtIBY/Q0jdZfO5n7FJpNYr7G70BHCzBIvEnTxLZHjeL0
4QeVZUAZv0+yj9sGRDbohan+gR/P7iO5cMfnSKJ12+gskGiuMGefwTDtKLOTO6+3vol+XZHsgK1o
3EIctZ/KLoHJjpABnKp+/TFJxD9f5000Yl3OwbT3hokyJ6eLKuQYL4M1ZZVwnRTuBc9+ReD26PoJ
fKPT3itQz581En9xvx43jfMKqcdjwlYNcoIQQz2/IsUvRcYM2jXuHQvcNohEEwpqvXPYI+8r5Z4I
18udeodnirY2Ob/T0a5OimNCC8WHJXHi8tqVkz1zHqTA7c3Gzjz4vVV8wPda1eOEt3DwNSSF6ePO
zbiujdNkOXbEbMnUcMpnlgmV5umx2pRg6mlsQeLSC38M6T69UenvJPUGC9F00+zildK7FMD8Nbya
C5TB1hXvmBQOsiypLnVDOL/RvV1xjxR2nHhhu/kMRuG8KsAVjAREUy5wRO+rket0P83buI8kqQq5
VtcNZOY4FO6pRu/paAnBMuh6XVgbs24RIWRIMENQMCgEVw5VXzr2YID00iBZfuncEvqdYZsmGYbr
qOUTB9PsqRgDzE4Y0Ce7ToMH2PvmI8GnBZJAfaiSF0Y0n9k8MblfxheirDV8/NR5jqJXACGueCLt
1JRfTzbWlaJ9Uz3IMrnAGXVmyFs5zTUkO6U4NiZQRKrP7eoDjUd1FDbtOpSfxyiM+VvKmRjp/Fuh
NkgdDf0jt2ujN0/cQoUiKoyBip6LKXdRHeMs0rknZRZb9PyX862mPbn9aQv5uTrGvnR/CdTvV3d9
t1uoNHFgZbW2S1BmefgBQARhte9Z7tZ3T7zFOEeDDGLZl45yslB66pA7mmq4WsrqPisE4sQM/tMr
59YNf0uVgDucM9NwtH5dTcyem1MaHqFiqCHC2PD3i5FUIbalfzL03n7EY97zTMBqFgZ+M6hCIMZ3
zNADnDx1jGfM1QNfS2/S1VGJR7AhvdqPVQBU9GiCuzEvQ2xB49eMeGFXxkmI+psHLTSr7zckC6RZ
QBuNAw2mBogqDuoE26iYx2czySoN9UjNnmbL9WlobGBER7XuDKaEHNQy+Im7aBv5SUZ1jJTN/cO1
MxmLSam2cPEuMPdkClkV6Im8g9K1OldWmWkpMLUf+7+rapLOwrdTyQIek8ak16rawsD191bFnPa/
//g3Bznofizm7XBXlDxf2k4hPl71aX1wHBG3K56nWkX4RRhLAcyNVyujWhGaYSXN+sET1GQbq9f0
EwlGxm1G5q6+8FLcukiasrNJA+PMpSyzy4maF7SsC0024/YimB1TfptDojlWpp42sviTpPkn7N7G
HsKOU9HfdhKUCqo3f2h/7NeQ17pOtU5bl/GUs2+z4GsVm8z1ZvG5nGmprmUWNaE+FDmBRqF8mNrM
IYSzV28Xnxu1yncgH1eArvlujB7/EXYVAcVx/VODUj0HoIAR2vaRUsyny/SAtwREH+xo8PDv67bv
gb2D1350gMq/7qeRvNKiqOVjshugBVtehcsD/CRERmXWce2T0IIxOtOM62hPjZX6/iGD/NAZSd56
PiW8gQdec6HrBcQpfYUXAUuB9EwSc/G5cC2n3b0kSRV3hWy4Nbc5Jb9upFCpnhLoji85yWIRpHqr
ly/sUqQbIcgxbZdmeW2Xg6sfrJaYT2lbKgqtObZ2URIEptreXwlaHmCEm7qZ4T2JKRUDX+56jjaK
dYFYlXzvqOqU8zrhd0WMuoU3WUku23/6H4vB7CynZyN8f+WCqfDliy6V4qtyOM7CvWIONkatJGBb
wnmghu62xZavC1dnL2FRxltFeHkbAFyyophS25UR+5N1/REJ+Mn0SyebU6KztoXFyBT5yetvOodI
vabPQVjepleC3dXEjBE5Gp2b5V8U3DEZ6hpvgSgAbKmEpyZ5xQHVz/YeJ8RV1VZJlTl1GxGohhOC
XVNsdj55K3RVAdcd/913V+D6SW5nnui3pm+9WT6j6aUBtgUtrxxoi88pdNPz59sxB2oDOzBrCaD5
JygyWrtnJwuI4ENdy88EgeUOnmoSa3iveNu7yZgxW9fsF1CZE3GVwALL1icjgsKbAi5EZnjoQZtp
rnOS2RXrfpkOaAXtE8NyajOIz2UP/ULasHKab5wjpqj1NpRv/q+aKkcC0BcY2pzsGFCFA6KRegUZ
Ixpfb9J2QJpt4Wl+4PhjEprVWs4iHkFLljRGXWn2H2jqTKanNHiGE1s+r8NSP7VMaC1EVfTH0FG2
mTKQXOMBgRa2B+S15qWjFQc/uFy00Yn9KrP2tGXlzPhgQwLSSg3YnVOAii9PPyg2AkpscG8tvSpK
is2PMZl3+p5C5xizwPRARVfONmJGMK/h63ozzqHqREpeHr+fWGvN7EVWY0qmPjbLie7TIolvhL7b
U/CCWSVXRhAAT4OGxjyYXZVeuNojdCTvVZVvVqABZ3m8teTPzdFw0gL0jRHJ4FIhT5I5n250jyhu
9R67saKh6i4tz3GuxQalKrS79DZh87TQ6ettDKgnI2+4pwq4Nhk4+LqNeXvwP7Q6QFOGlLMjawvm
lD4JB3E/PdrJMmXUHcamtBzPa0HLntvv7VdhUQ6wgrQObTdKh3nFoww6zEbl2uoGyXBT6XfgvSCV
g9/+/k7KhKdFjCEdvkDTy/3RX8Owqd0wEVyi2uHGQJ6UsAMlllyF8zn65eN7IyWdYx9kFqI4Q57I
SKf8Lo/TD4cDSlk/xnDMnLSZa2UlLphkOQzJDdO7SxJtAr3CpjJGNijgJGB43arKJylAvM1aCu/s
9XBFEibvrM5fr0HLEX5qckp2RArnRw8dCi5QtuvM/1eOvAofeF2aKA0YZRxzRzH6hqVajdpiearH
IO//oNBSJGF38tRhuCiyNKsqX18SHIb+R6zOxNlZ/IY85gsovahoGTI7aA7y3uQN1jqaeG8Y4EBp
1sN9o5vsIwLVfNK9A8N84pJZwc8FSaDCbm/LJ25aJU3VoNWz8UucfCOlbZc+aDNOW+tS0rr5WA6t
DOSCCw8+p5SZk9NoG/vZEwoaV4hK1tmhyGhMiCXo8fykbE0BM52IwB9mCjH7ffyX/iKFbVnI8otq
lHyIMQQUDuW6OcQGpYBI+aQVfYPH7dGMtkQDcFYOOyy66raPlNpniRwSXTYauxQFv8EZlFfG3crh
YS2GLt7RydwgJAwcLCNnH5Ik5YYEfrwTKLLkPDqjLNbJhh4f/MFvOOQmdqaO0oEezf/QzH79d9zc
Y8OBVZg4IUCVTwwS6KoocTnNjbiukURdGsd3P0h+ojLQ8s0FKQokMTxyDvdMCl6Wk99M5MUxrtTS
DRaFLbarMToBYHqt9bbKPfLuHPZbAnEfLXNNRhkwxc27HGeW0bwMJj3o8kFadwycNdNi+kubnf0I
J7rbOmEmIdWfxA/vBxaLu7LXFrFMMaM5w5nowkIxM/UKT21yGY1XeaS1FmH1VEo0P+rbxI4MyCEq
holJB/pNezINBvOzQIjyg+rgbxDfYyY9WbBXbc8j+ksEEYdDlXrReRUx+68FEmw5BMMayaKvYBCc
I4zLyFRuvkCkoiMNnMk+C8B/UJkuc7lzskzIgF+q6uWspzYPBZf86m0t3mFIVPUJjIrwdy0kCkhZ
Gr3YoPDHNnJqr1Vh2bOCKUrD8p+poLlVHjlnw7zPaWETyG91Tjb143NqkBS/CMwEdt7EqiE5ViHH
/ImOqC99Lpb/TZ0fKU9uj8QLkIQId2vVI/8D6lIM+GdaOhhEHrloo7Uj+nU6pY7rjR958r4jc/Gq
dVvdK3+ks2YvO5z50jf4R4zlUYqLXBFUnP3Bq/LrxbiMPqdws/eXLhVm3zEiMjAAvf+59TH5N/IZ
hYOsXciE6oJH+0kh6LjlUJUr1tH+VMI1C8Gh5e2SsCnZn9UuK/kmqH02PtrCxOzyQkahDCjvs2nN
aoyTS864txG+jSLdFfQge/+cxq9ONGjedEo=
`protect end_protected

