

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EQHbbfOVL6gqfpeCpoISbj+lHfKr4vlNCL18x6H0v0zQdPY/b8eADbNrvmvYjVcc0Tn1YlW6/oif
3vs3Nzg6iQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TWVAd3vZuakptUOe4SlR4HP/Qprg7tREK5KZyHcWZuI4prRJIyFeZ5KFTat8JfgFJYjNQZxQtMFi
t43U35kto+eyadS8hUd1lp14BAHOO/DBasc9vph2b2xCcxsMbIBLtNXOsOlLVqylmByUyppDFqds
sQ82BR+a4komiBeOV50=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
i3hdWV2Btkks5l8OpwnLTliwlr13EwxZaIAf1Y3tcSPZhDz6yEu7xxedJ5lV/LyBvH1uukK8zPLs
Mvzj9izn0HqDESKEPRrajf2E3LHbg36g3K/SAL+uZLuYDo8Rjg4qPZr60qGzcDINBVBiaBBVYaJZ
sinW9hN5toHGqKP3wZsxfdpWBzkFWOf+kDKWRV1ONKUusqD7q9a5/mIpC2pHr2Pn64xHKavTHN/y
IFfznTRSXKoPv8gqv4yllwaZtBPAFZakeoeMwcrBd+xjmTk0tnsXJzsi2qtIvWjU7Xa6vS0b1A+d
jq5ObM9OSnauk4yDCMPAepQm18CwRl+18wG39A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gZj9Iqx36t2MoKbloLaYjl9TNovjvifcJBpm50Bj49eEXTMMiSI47gg+XZa+IefOjgwy8N9yGSWs
up8fFGQd2XZBecmqIdgel7DtmTzveHJd1eWih2agQJJ/CKKN2wAHWVkuxo1sN+dFg5l/gEyjlOzc
xD4WVTcJCSefjXIZXh8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
d2ddZOSCnJp4objvLe64SilUiXTFDb90g73z8MBtePMbmoXnX5glCMa0KIQtm+CKbPk5DYnsMEkd
pbn2YC8EcqcJL/knJy/CgD3l9RTZtMeyH3koJIHeZuccfhbpx1iaQTf7tMFx81NrKmtv/1tphcBk
HM7xXoVr0wlE3XF51G96cxwGAvygKRbI97JtiWystSamKboZRyeAzZpl2Zo0rKOl+/tAIJCz+zp3
i90v3e9UQcn/BzNGJrJPt/Hfu3SdUtg/KjGA1q5Ud1nAOI8lq8jolI5fslaEEC37Qw2gUc2w36Wd
z7d5uWrm5mb3oJWstXofS6QSqCJBQlGpl5mLeA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 132448)
`protect data_block
zxs0UI0EGRDUsU7yP7kefF80C3dijPYSX0qkMrveBt+qCrQ0P5BEa6sMdOK29W2cuIetCmQuk9iH
Huh8URKNiJFwcxK20Plt0q9T8c/Wlz/pIZEFF1zgcD0OKqj8mmS27iHYfVoEAzYsSeM6Upv4bw3c
FXliKOmFbGyycN+4nfqAdmcW65XvZZDNj7va5Biw2nFxJyh/ghsD1cG2vL3cAgx/atUmIfyVJse9
GCv3ZNNH5DVO/a9Ci6i5qz63vpKVBfCq7ydcwA4fgHnlfFZWdnTupl3WHON3a5qvpOVOkOaXDnum
T97qoqhxvlDNPEkwkFF+3yWfPvGwv6/XXnBLxfJl0CnaSxFlpRT6rGD32Io8tiTVfqVqpyLWB/62
cwrjhsE5dWa+dzloM2viX7S9MBPTYurdzjMrK6JIryKBWboVKpNlyvwYQ4rf5LdJFieBhKyVIUH7
PIVliXKiowJI37OS4K/D6ImzYueq0odOMbGydZexF+1NqW0gbz1/399pHaiUDxw4ZFWZGx3w2aOn
5wsYeO3/pPcwWQ/uQ6bZmacJSiAqEtj62HHD7YbwXC0h0LYSxtlxCQmUtkxT16GeDZPlvfOphBab
9jBlp+Ah4evnxwI8NyX9q6a2rR1u2XquJJR0h3DDswDgH6F26gOxLK52qwjdqkSYxSgStheCvLPq
wNULsXjIHSMrGpnOL2s6hqao5NI6hgtv5uhoeq3LuSJ8iuWKrLzD6FxvJNb6dbBBVZSf7KBMBasQ
/ls2Uh8345wJwKZDIqDpzUNBSV2DRRJFEaNN756rjtDPTjoYe312W74ouhte6h/31P1Idl1ZI6NM
lncCAwsrdNw6WkUeqPwuyqFux1CzsddfxWM6L34N6I815oamgVBCfHi76L1o4vNp4Mapy9JEYHj6
rtxa87m7O2UPkZ7hmbQbE/EQ7QW1clLAgQOs2vSPF3Jx4lCpR5rEOhlX1q7DK2zK704w82lrsxjB
2cz2bY4QrY1ABlDgUGNGpHj0vvpaQKuEbfePg0wUyq+O2gQBM3dFTeqTNR8eSDcv//SN6S/6ZQnU
Zt29TQdhxsu52dlpzqMDsKLwUn7zGqzQIJufo/WZ3Pu1kO2oL8qQmiv7/+AHBXt6MuHnXctNG3jb
WkpmLWaVMuHEosSx2WMCH26ErvTtsfjBqM5OcJjHA7Jxqv5fdleb+7lfurlL1zjR2VEUWXDu03Yz
Vsb+k2bS5lcrQDcy93+eAvV+okoaZoDWTjzbACuFlvfsumpVrfNgef+/gGyPQIw6uDTexR22E/+c
je5AT/+xDBXMq1f8ceiKTgzNDkRykqMmy35GWOXxjiEY96vXaYTsa8kg/JBoY8NhCJ72MB5pKZ0h
Gb6T8DTW9sadWQRTLmdt6UWh0EbbzmmSg3nZBXMDIe755+c0H4rSuRm7HaiEM1F9y9QgUqNE/g3F
bjYq46lneYHGiCTXcnOTWf4gwZR5ZFKVIFvS4zdAVd0JFGQVcfRsTsTHwgMzOlAwmvBX2zwXT27W
RfGRzoHPFaQAdhMEm2kWL7HnF2clYFeQW8F6Ti0CGiWMAUFH6grpn8wIxv+dXzACtuw9043brNRv
bpz1E1O/iGkJMndmnJgm0ZCe8Nw3WIDekdJZ67IrITCrI5dUGxA7ZbhpYsQGt9fFq5ZvH9AJTTtW
j3oCQmmPSiAxQQrSjkV4qwCFnLb/PlnnfaUOucc71yNNMLQYFCZXDt8hURJSttbB2E749tzT+sw+
L5woOmYDVR7pgI9mZSMjHjtctg0qhTXonnafOAp9dMJK5X+bOgKK3Q47gQDmmhKdp52Yz0hRszdF
rT9TkvbDtVro/Oz4jKx3/khoVz3qgRLMnxOaeSmFAG89E+fXULwT3Ar+hVnWWBVsgi52svax6qGb
fzs0XwRu+DHr1ZOywCIJWaGRtWjFignX+sFGQZwlhYGHN6qkdFC+DWlYpfGzvkDYRH5+YXo85eKr
HGrFyweZAcx1JkZvNqP3FR6Ifw7tnfMW5L4d1gCQhkfqr3vukkqxqbVt/ZDjg4WlSiTl0NrlQsv3
y4eHTglefFzuu7IyNUheWtVidoMmzM/fg97kbQCz++f2AmCTj/pohoiWO62sc+xDydAojOnrF2bt
iRi45rU05NLRNe6dOwc5r9SlRhyJn/QS4DTX/jZbXIsv2xpFtZNXsV44ujcdaxqBfYLG1adU5dyp
YCG1ssCVPEzn1xZbWflK23NHc8X3wb0ocp/C9kujTfLFip2Nct0X+Szc/zm3ntBEKdJEj29Ok/bp
a0Qat2L7lcS/5KHBkdl1UwkTlvftaan72JzuTHGovP2u2XlDX/Y6i1MY/4z+FDDdQBqO1Nw54hYs
TL022dGRVV0Ut87Z1HUsR0FOKxt4NO+EXPSYEU6RlVIjONTyps0Xi6+AY8Udfxwsgsz2nmndSr7j
ySZo24Le2Wph1Lfyk4u7o8LjUZuUYLdqlPL9ApMnKNamfNCP/HYjuXMNdTbMhFmIcFFStSTjMg04
ALTqufw4nAN/p+NixtcwaVyeGNPR1Vogpx8lRVKw2hnUNcQH162QAhNqQHrqRIj2IqLHWsV2ASTP
o5ljfAopZXzh07NgU1o6E2jEeo2WADdZhCnjpoIvsDo69FzXi+QH3HJorkEP01/rqGHCsiYDWtjf
pxRgVn9K80MxEt5rYBhDhV054pB+9eSqw10H/9rUmBaW/A786z3UEa19i9R6twhn3DKXpNXjOZkd
7gw8tWMd5vzSaMXbho61LnIPozz+LYgT19u7DOxoX9mS8voZTS4HaJ9f/D3eI7+vvqGUtoUlmrQF
SJuhM4FlGpSWZwz7xyvpAHXSCf34EW0aqwmRwatTKBwPRcpAe0KvcqP5P70Hm/2iUGRnY4fFrga9
7BTEW6bvZYTw2C9wJ+7AcSt1FkvxUx2+4q9zHJ1BTsqm6AEn5xKf4o0ABFJaJVXxgL8OMbd0JBXV
1BIOVOCuN0NDvNTaslw1UybamaK6AM2PkOWmDhrdMF7gTkN/n8iZ3diQ+ys4zP53u6ReaNtEF2V+
lr+Bu5Ew/zTm1UwGMiv8hwMJuW3iZbey48shCTRX7DWv3T2XU69yRqAxcjZ8e8p1VyeOu32FLWcM
ioXiC8LS/TN9GIZ9zuHXAu8ckmfSllA8hTRL2AHM9uz3QJlk2vAFcwprPzoUM28ku0gUygcrhykJ
AP0I9j6Py9/KOksyOJ5BPZv1e+em5KKnFNzMp/Cj2sBr3wZ7ZABsa72Wq5BT/ORvza82/M6VrMGj
mOKHhrmRhWoNiT8fx3rJ2Tkv2BXbk9aAXPPpx4iXsB31qcYzzENWZPxe5CmoiKipY1wLyowsCqOi
tqEzuHnO9CEFMEr2TyJHJzQZegPTjFNLPgTyAj6Phn1sKTNJerK95KzOwQ96Y1gL5wvjemqFqazU
ynblkU3BTQ8QexGUx77I95hfWg5v6TYukYAPVufd46yiBC7SoZkppufTVmihiOOBfz6qAgNOdIft
YsQ6OXLdI368ve0T9wXy97A0YdzRRJp/QM4EKNlN2Grbf5spC7Y2hNpLfdGN4xFMa1x9GX/ICWKp
siUOWIecIc/uhtUB7ehGDJpGatGORP4NMMVjmJSzuuOKzg8EqFh2XA2/GfThbWybHIqMyj0XCB0P
ekXI5F4TBOR9/27SOjnR1hhdCAmNKC9JUj6oSYCL1wHvjir8pgr3pu9N48klpAxrrAz5lIWqheRm
owEDmh4REiINDt1VnB/equTCMInRD06JpaXRK2/Ocp7qmvJbM7KuzxPbsNIlk2cGL0VHRBp8meDQ
iMN4YryocZJtpAdV8c2a/PzqyxG3AVZvkemhRFZUJu8KbKeMdsVT2r9K5CydocB3/5waxXNzCXy2
iydJemQQzcQtlLuP0UwWxDj7H4DmeaSYMEFe3026Q/bcWJT6KAKYqhs+SaNguHJ8xWxjloAWC66n
HhM+Co7USuHLdhNnf60HQghKcnWoqZloJ7dgglvSpri8pvbEX/l+Lr1y1Cwxx/BVEweBAIUo/i45
2yXpov9d3LcqKvx46HVUOVG+VuCmWBApSSP7tBNhHG3uMrbqjRS6rZaw0ouL48Euk+gHUwe/WMEV
LFuXMHKVxfyZz1Koi4BbUUl/KsTLEJwDWnfQlpB0tnxis4q5zLaqoPAE6fnvxhf4eh1rF6AfzuVh
xTnUlliY7flf2ls6AXxB0NIku319zDeFNooulJ1/oZRSZjJzwT37fbNduU1/aR9XGuTTc7aaW0/R
fhmyonsIL/UAIMAFl9Bg6vJ8mLb1G+yufH81tph5rF+oHzV2tRh1ggTeJL5Pndq0qC9knwFILaNQ
lBBZt/MNwLm1vIkxjafLtbkQdpmY+3ET8xBIpib2e16IMQGjlR2oyu0oc55fG277mX4QRSODAFV1
i2s7Km8PTMtUR7YOHSPCEKeSJYN9gqwCdyXfhSZewe4Xw+KaE0rImBhJkKyOX3bInnQe9TJIdvQm
zsSH4Xy7c/xiy7dzEMK5uFMiF0Rg6SXSLUnuCR/RaSoAimL8vrdL73/cGwKYfYQqX5fdL8EoYAI/
FtyuNqH/8g/xYxdwGiijcYkn852ldFj97ZDVYQ9NNEVe8zTHhx9zKIyfEr52N9CWu0lBmPFWSZor
gGHkwv6XGEDbUbzFVyKcZ6/ZYWx00/lXFBQ3rB3r3Gx7YCJniURp4pBFbFUOJcvCaK0+nPzyB5jo
pB7w2UPvh+NbJgwtXPNLCwV+dKoSZa058Ys7nRJYVT5ZONtslFEfE/LKlXvepouOUbX1WV1Nfhux
bK/AZU4qaM89hD1SZk74Hd9Qy+BU4ch10ZZOfcePOQMRrRwzHBdjRhAQ9nXIooXZcmOpFOhXvRbu
yKYmht4E9vulLA+Fco8Yy3aHy7tsvtilthxeeUKzDlf8FMtbBInGfuANV9Xkhv3gzOIUQftlafcD
ggSOK1jNsto3b0OTA/XCvjbpXp47GS0CnMryvlDLLSrIg155DIJFLjePtreGEl+pu5jntS12+G2Y
vadm1EqZ9AN63WdUrYMgTn/pehqKJhsH/88FSuEGWN9LU+U9uNPCRqLyzu+XgP6qPBE3PjT0UpB/
okhlR7ohKegVzHh8oYK365v6bLyAiBaS2quF1v0RckiwtkMaH3/qMOtu7IW3Ra3G46pJLcr9xkA0
z+6b+mIHNu7K6QpntHZREdZSMPkKt40IJ747vhhRb7U51Wt5G0/QAbg3X9I4F26AQJcC7jxJqZC5
th6GhYZ9BwAF9G1WB4gfq+ukh7owfm2eNg/+3UCziaZQN3+RRRL2gJwtmm0NaFGgrNStT3rnTjGR
YtLXEvARhPwGA8nURK5SB3h7KGiRSpvoyagP2YvIpfyzsq744wQOjs2JPyTlFJRuc05MbK857hT3
xt8eAbNSo+m8atqrm5GAE8yeB7ABHepFZ498FroHJfdpSaPaD2PXdaKu4mCxVXKge5KXJS1rnH15
q4fq0/mb5PtXEqBa9wJIvqg+DukMsOAliGMl2aKX0xgM+xT625fOPhVvwJ/p+3PLGtxmYIldkwtu
EtXNX+dRHv0NyoVsoKXlsWuQu95sKVteKef1Wy0yc+7JZJ2C5LiRWsA5ZmpGxj0JT7aKZe6/4Xz7
9ZWzwv2M4l4ZFCe6D9jBdvlWuXSuHPo7Rv2nHojvimLE5zRfsZKSZLHElMnDFoaScz5eUM3drEij
2Ub3lgwRQAtxKwR4znbFDz+1LX5ONyj6yCqUiC4o+QVtbg2lTkn1KSp1ha7KmFrc6CrEnool4qKX
2LQfvFjkv0RNduEUvZcMb8sEPSovsd5fzwZnkR/pDC78LfpBMuOyAkJzbDWbQ/uL7Dj4G3ThGD5b
nhUlAb3C152in+sO+wbjMGB2sAUSc1IQA0ST5tgi2tuSiPgoRYMSXMgcJCaN9D/FZxTuMLCy48R6
F60IwEuBp2kfi/+2n6cnZe9YKG516w1isepr1GoXw80q/NTaHCkj9ewQkEkmJuhGImL0dUwzJhgA
q2xxUBLl+Tvg9eF/VccJjLOo8BYJbvXmFonvLsOeuq8Y8lWJnu9N2eCl/MnNadjXI36tkDn0SsFk
8rxV0bxoWMKIpFW0EfG48x1/3P5I/DovZjzjkapu6DRm+Jk+x/EnhsDzYRkfiq8O7tdv+2DXHP6j
UAC+Fbz7ApvVNRyGMVZ4iQY8K/WK3Vesxuov1UXnq22vCiA6q9RK5UW+73hR6+Tlm2tmZUUvOfjj
zbCijbIVUa+5OWOifQgFKeW7Hrmk/kKkZdWWkCSgB2V1cwW4Y/TV2VZLfLcyMnA1j5OTNA4Ydian
vCrgwUsfB4ISbM3nYh7dSrqDzBK+Bcl8KeyL7P1JIsM8k8AEcVcpFlVSbFYSX0betNxT4THDDqGk
nsm4C8WpsddTL/x/Dvuow+OLYpdUuO7HJuCqsLTmOPX01hPn1fdRQjejLocEStFVxhyrn9jQD4Y0
UmRUdexGiqwnxH0KhqM61ns9Egz9saOetxlEZh2GHuAL/HaH7XpptcHjfyZLUfnbS1vAWKEB2QUF
AhEHHkitNnlmbAMs4SNlEQONWpvwERQsJCMioVwKR4K30kEhk0bRfepVjNHmGz0PVazqjJp37ORG
GWmHhhBWfxdQ+z8PtS64xwznCCYz7CFqpl6aRloqcpJQZFSBpnSH2j+30os+PhhQxSvQSkR0jpet
FStml+rs6mRxTB7JkmnNy7/FOG8kFSg1K3Rl1yWBmOvHJ4cwBBkKqfP/PQepAOPg9r0PosO5LrI+
V+ekh5yVeg7Fmj5vvXA6uK+abpAs7u3y7hy1Y4FazH3m0W789CuElZAfHnfiH1Vp9RJTlQvF6Amh
/e76M+7SC/MmLEYW7YlszoBnYuz5PMlUNz1htJKfOSMJCvI+TJZvRfX5vjzSOlxl233+ROvuhYlz
VdPIUlj4ay8l3GUp7Fs16iPBlHjDXvGEEz5eUItEzsSqxoRUBwcPbAa6H+Au0C1xHarSg22y6UnF
p2XVZnVAByjBzyXGrRT9Ij3kJYQunrcvizx6AIDRgxf55DzZtBSBeVmfW9oTAyax4g1aP3R5QT2Q
3z0XdiZQCIebx91gPjG8yvk06ICCo7z6Fryl4Wu8xgERue2AGQH2vEe9M9zg8pgbPqeNiEEL3DX4
P0YGQrEWCBqoClm30RjxDylQMqq3u1WKi3C7ZDetEOd4XqcDeatKZBwUyL0Z1puFXID2LTSs8cdo
poZbbaL5QKSDAbnUP1ehUZTR5j9SfIyXBGw1zNKOK90y1FHuA+QAcEqBbNnlx5JKKDzpH8SyY1Ff
sRqKHiWX4v9buqjmZxPtujfHMLc18Mb6TmSLfoJZf/rnuhtVJY4j9d12JHM3hYqIE0zveE1L1XLm
FxbdacMSSQdN+xrsIc6hsDMvbBJO3+X5nRc6mw9EOkSK89woz0Zw94vVUvE9WxClNhovBW2P9aIh
IYjjaI25+RMTrYBntVHWRRYF4vk9LCPtGsU+1Zin1cEnHAsDR6Immnl5LmFIaapWDAKzRpzfJL1C
gyGdFYaYkyndH5eg060NsOJnlHt0uEtAVcbBdQ6N92U1wmhYqKAuo15YOlfCwDFjLpGF6yZ7SJUo
xorOBidFsuIB/DZwrc2g+aRphjAbvrDu+QbU/NunjVRLDtGZAB7MYhXUtoQmePxM14IkSZEBffKw
o0zm+DPyonhs97MeOAeN8lpP21eqFBevTMSdhiVjBHzFmuF6bBlGO5ra7OiHf9skFIgUH0zRXkP7
wR9fGeOeGzWYK2Ds3pYAYpCcqTrG+PHA2zfCEPeS6Z9MRfKH/7pmrfaHHdPHxEMY2/GodOA86DZf
Ct4efGPtfJb29fystA1yUwIDzaWcELRTwCRfWvWaDjgJse1J//3lLXJcIHbzw04XRllFkpYy3naA
2OpRgNSslESVQp35luWJVOa4XmdCNVNOGdtJLMkoyNbdLkNYjsOfyJtMlJ6ez8yShDv6N4hGzw4V
nm3ljRdRZj3Yuhs9jQciVUm7Mt0RxpOqCe9TLPO5i3DkLdT+e1ImzJX4whe003yMdO9vov/k6XlU
QLnuwMju5KmO8I9OgxJERwd1NzmAaCYvWQJp3JdncKI4CDMW4cfPvvFlFYREws90GZt8tSaChV6i
UFtzImaEEFA043YA3GObPbooRMJ3Tg5hMYqu0YagwSNF80OVqFj9nFz83p6Hu3fOoZkwoWzG5Bvz
tgyIhDgqP+s6eJjmyLJ5oROG1xa9ETWYELs/pCDrRGq5LFR3XmA9Fw52Bltbe0qKL5C8SuMpXbAY
rX29zQgPCRidxc29c2iWSunOk4IqGPBobfO4Q52pQyIWqnJkhAFFNbJ5z18Qw0IbYo9dBM5pw2Xd
xpWqg5niMys2g/mBwyoYZUOYvaEBSwHwzAS446BX9HUvgcwTSaxkvPVWNam0r2dPbG5unUydZIwh
UZWssgyIFvNB41FGU9iNQWHoh0V7UMkqfjtWsTnB8hRoD0GHp+uu6pXpqXoe588UQ5sT1diZco4R
3BCDRJ6UQ0zA1ichEOSwcAcAdTUMjvjxLJp5NFyi5J6d6QdgOtkJrudgLg3LJPBkYeYrGfz3BUjE
00NMRtnNDzW3wy9jdv1bhiDLnDroH/cupyrjEGb5FI8UoLeLAg4lIvStd1FYbPAASyAwf79q0VcR
lJORbmXJWuxqGXqIrXsOk8DFolUfau9OP06bT5hdl5xI6MJzIr6P3YBs3R30Q9m+Vv/0B88Tb3bZ
xSxULMXtevw8v+BKTSh+Qv84DF4+QGhuxweVJyHWnYsit/mGo1k24T8BkiitX6hShMh5sO7rkTmF
oB9LmypsVgDA3shwHx95lSOjy0Em1GRZXUl2OeUyTho+CwwldZYPZbVWvucnvP7Kw3ADIaV6LNLl
YcxQRXQ4ABFjRlZtFd1Dd5NFEPQdHRx+aKobzrY9Dc/BRFEkKSQqjtqJbzShCkXBKevjJmB9NBWL
3aRWf1JDJB1L4n2LHknXjBq8vKzMI/dUoISo5kyv/8MHfjjn0du6ZPmbQxnH2pjYxAYxzwpItIFM
kgoi1xC3cxKfcnE5go1/O2cks6A3qdEIWvXP1RA4NuvT3PjjRaRTBR3wPUBO9HsmT/tzIvRPuiXF
plwdieEnADL9x+gcNkZbLs0Mp6CMn83LVVXOFrhBlSBYjazH3as1r5q47zCe3CXJWXXV47Amu1HF
Mnn893KAw62MloiVvNfzE/NW9dXXAVIrN3gxOE7eEvrEJjG0xIRGnXByPWACS9JUmhn2uz686E1T
01Ek7SySXZVV8MieFA8CHeL5Qfh4ZyQDln/rryVw6Ysq4XBz154fA4kOhpv1QsKCoo48hbqGbQGk
VLOV7ecOA6b+qO/r+ZucASO8A1XkSXTtYlgEzFHkv533rC4nP3TZ4HWuBKcFpGlUH3eLwSZfW3pR
SLCleStB4JcEzl/VHJt+gknNvipcBa2cS9/huqYHuw08fDVvf0uKeUhOfSvd2BoYgGnDIAjTFjZT
/yjIHyrRbsauube8FDf01XNF8gYJcClcXLrWp+PR4IDBQ44OAKUF7PGd3yT6bV4K8N75fQVAsVor
Uaj5mOymP2ZC/7/IEXf/InHPOlaFkct6o/a0L7BhJe3fcLK+zurDg2vOEz+FvsKG5rhb7dGA6jF9
2YzsZeiYJBhx4OZTF+9PtFEFIlD5rmXaAAeqoRay2z91OPTOwFF9qwsBJ5etW70y51YM3DS1/dcy
wcUTguO5IisJIS0J90UbPaezZh9rI5y1yQLqg7Xhbih+Uhit6CV0/oyom8yfb7COjl/ZVuq1uKty
P/C+xotQm5LietN8FOsTBLLm/Q5ZeigSn+Zd/pOC0bIZdeLyMaD4mTUlAc+FqGSbqdlBcCt0V9KF
xiLhwvripICnXsff6+dkM77jTs4iGICxz674vU6hU/YlBDNJPbx8lQduOSD0gNDRANy//LWt9Rln
sFr0U1yEuF5BRC2M60FBPYTOlCPn4rmy8qDPnQZCoimWgAG1rNnALxSt/vFgLOXVzcygsDtqnl2Z
hmdCubSHk+EQvPESmRLP1sDWFA7m4cR/j1zcCDJjQJs8w4Ko+YOnrPIZRymmjYTnIk9QJhvRM3Im
H4jr99SELUSpmq8rIUzQol9XyxX7ewSJ5GlWe/4cJ0DKA1a8wl+QdjefcbHsRTizugH4TVngO0Lc
A8LLRmWuvRTN40d+Qo3PyA4p5ydwG9tr+o0TGvDn70zd53POVIP+ivRNdK571/2puGb91Fc1IRH/
Bug1n0g4p7B8RwaWTcaU+tdcNd9QHhNaN29Wbay7NOnbWvqlU2d/T2DZmCFqTNb/po3uM7VJDtAn
I6Hzl2+HD3MEIXPpOfHEhoeUww5y7+DvPqsbZR+zoEJ9W+/P8FIa2vnME3PC/BIzCgih3kuWYmDx
rnLvykGj+GNo1F+18ur1qPA087bWutHD5Xikg4aukw7J5SYUjrlQRQzM6kl3IJ8v8+W5urxt5DGr
9GV3HORgjs0i1se941zXOoCQFML0R6P/t3cEzTWBnx83GoRekJXHs8qfeFi5Qs+hgvYbovKeD4Ji
t/G62SBa2Tfv1jgsCBIditprqI99eW/HkQULhFqgSGfc2CgTapUEPxC4aNRukUQrPXT/UMU0njO5
oukxwQM1oEXtQJxRYDo5M6xGucYnFFA2fOCtCo2KiNTnlAbMu3fYh3PXeYACZ0VZxxY+6ptg4zB7
4CySD9Hn0dZTMZTuwqHN6mQSHA7aBAfZHcUyMCH2JCfBjMzIl7UxffxbM/3zMdJD6PYzl9Ne4QO3
fQNKTQRIy4ECt+f1CGJUWJELcu11jxqF/vJVOb8YJ/8Mx5kyNthfAT4a9L63P39C/MPZPi5zp2QP
5sYRIvnuncR2nZXh1qePBBYWOR+ArLeaMmSzbhH49PpTCYvbiW5x3IaGdvdxynpBpfAyFPuU1ggR
4V++hGZEaepV/glmo9R0s42cnFyacES6w1+fLHAscGts/t6afJlo1+dqVRwY+ap2ydh3HLZC+Vp7
NMbOt+u7MRnk2c2mzwGXduY9NzRjF5klHWGvLTwQyjtuejWqiirGDDoiH3YxppbphzjEa/eOSZqZ
uy6eiXenmGqWGtNXRAy8Oqm+XgZFop0tsXP7nl98g3hIcLL7UUophPu1jGHJqyLCtvEc1USrGq7G
vTdSfsSXJ/56KYpznh99xYCIZIwvt1W8NZ1vO7f7JfgCMSpNPO34ZnPPehxT6upD9IemegWYusF9
tbOrZMav+w6A7fuVg10pxiXc9reXE16YiMACvnuuaxpnF8bmpsNhgWpGAakSODdjACrVM93YfQ7r
NuNf/W8zXcVGqzhS28RDy34nT67/X/Jvap5tXzg0MU+n1qIyvakstT/5cJhLFztQn6htAjwx1mA+
FbMf1dPSxaoy1F6zXWOiAQL6KDtb9wH3HkaQC01gd3Tnb3hC91JHbqc1faScVrJYD2x865XwzsUX
cXyM5stHwlcu0d1Wf97t52AEMGQNgCLwgzhw/LunUtV1RDU1WAX+BsczpRY6/ZPuDewoBU/YfwL5
Yi42xKQ9xFl7NTK8P6aGiZEUnGJpAbY3cVTEEVDv/sBfgGTgS3LmpMTTEacH8QG231jl1p8kavqK
UQ+lil6igIIdPMZOX5i0N0/t9YNaz65mRDJPh4VGl/JVi05aga4Q0I18mF0PU5yoh222UaylG9PF
qZCFVSb02YDGNgllTfdCiHkAqQg/wG4cVOoOme1uP2T14Ss1XNAsUiCJIuztXHWomYOAZk/fRTmu
ddNsKihu1owlplGYLt3ARvLme9K9CLS+OevXjoaG1tzfuU3cekTceksSEuvVsXAi/NfH0LS9uHQb
KnrgSmDT3CM9+SXQT8mTu+y+9a7Ys7zk6/xBi8mr6iLzRO3znWEpEsciCvz7kL+LP8dGSrOYFBod
OmYHtJQMzrQd83l2vvEfN9jR4Fo79PCby2PFNmKNpjwmj/MOixh16NxTDTOTzmxVK8T8SYd/+nyU
fWi0QrSE3dnkFbwXNGuGiDXRg7MDzjvLdXVDXd5YwvEwrr6DSow2T3exS++9UVa55b6jK/d32Ih9
rLszezDyiYD6UpPTS0gs/TusQ6PO4wIPDJrB8txkkZ3NbTitTeZDpPOiEhJ4zy3nUIossSAEromm
5bUIytguluiEYCR95ni/aFz1/QLJxnYlgCaYLsTBmJyfdiJtCZ249Lmf1gOVYK5kTmjBDw6QcCiU
u+xbnBh0p3WIq+edyFnPWoHL8MRK+LFKnr4xbVfMmYnENSw8Av+vUYiXvUOZreUrrLw1UlcWNIT1
txFT4a70m41rkk2sOjiaDMlf9+uFJ/wwA7k6J7EAJyeyBktXkvAPHMNiuSmH8RtgSZC5SaBQ7TB5
WKUu5sc3Xj5/ueiVl2KO7B0PKanc7oIZzEs0vBI7zD7jyr6dOOL6uEIU44fiRvVLxycVvRfCSgWh
tV4F/vG+4VehohVTZd0NfGD6E2Io+/QeiEib7rkDymOuhbHGJAaGP7ioGEdTWea5ltkRP4yePYHp
tm5lYQ1LKglH0aWOLzRpRxp80R9+wreTGqm1rXQIHQIJhUXIv9qRVfE+6CESw9DSHCKwC/N4jfUk
J2dYrK49bmfVm9FNUwA2FMX+VbhkHapuEibG2/zADH0cJ7sVGuzbkhBw4xXm15CKiLNdiXdHlkQu
PfQ2fmsIzTCVvSwjfdkOU7PVSE1mjs7iWosWHFwpu6MqgvqPWky+JBY0LwFu4L2xQSrfWJgRkGgu
xyJaqUHgWFnjQDj3UojgFZaUhLb8oExeo1p4ZbT0A41Dq1gTVuqm+StOZkGVJPboQm33D7BFvoa9
gKqF/FN/oRaOGNv8Q1EWu6FVc4wk2NDvsgiNO32IjUMCaJz4gBIExkqosuBD9W4m4JpQf9KxjnsN
iDW7L6eDHBqelZUS7LH2ix4iGXWkMoYNoqMfKJDBv4l/A8WQB6HZ47y9Yy7fs0JPyf0xpWhVB1A+
A8+iexjAy28Dt4h44O5xL/R5CKpeMHyB62pugtgJiRnESNhlQs8P9LVYpza4KsqByaDnWzrVYoDu
nubm/k0mwD0eXA7upNTffuyPAvpjniti9EC3a83a4LuP+a7pWn1U3GjKmin7CtVvrE11C4ADhuw5
mNMcyKSLzAc3ul0HdrCw4LvcgprfoHIQiUELvCLztXmlHV7ZZ5Fjy+yDcQRHnhDW1ZVXkNbIEnFl
K83I7STWW+CEbZSiS2WQpxy9dfBezZ+wQaMSu3b0+TkQm6Euu8cdOON2w1eQEmiYPQOcE3oAU/jD
eILc58yN1T66sWkaNqErPMVzD/bVrSlfmsyHoCnFYMH9k/E44ic7ThrJPP/EpELJFlXBgLfOpxDZ
et8QxYIInJKhHvUkLXhIhZ6CZSNMwd16wa5IIk08Wo6iFAFWbQMl6gKJa15elv6AzdMydfTe39g1
lxEg7f2usnJin6tOTjJP60KgZSss2w/6jyLiNVEemCrXqfBwdPDvmhpNxLO2V0oc0quA4Jhu9ffH
nuaezq8bcjxnVtppFdRpLOg/g+TOdrh2qSjfhVAQkNVdLAM7nJjnV2v5pCafHzk9H4ct3Tn+a8Sv
qupTu2pbm7g5oH2XyHyDV/QlYEd3KWzgx4hF3N8aBBWMsmJdiMvCGOhffxOhFoum5JezLyX+FzlO
U4y6YzdbiEzklq0BX4xkqV3uqj16i0lNjWlwDwVmVuo39SO0XdrvZGNmNzBfAa2G+OunDJqds0hV
QkXiJkG0wosmL/BkpXtXqYYnSxuWlCqe9tWWfyegQZMARsK9YRn80OkeuaxCxLo6XHz6DEJtP4jK
RCfWiuhE/oum4eKUlV+NlymMfi6fXy5ksmsa3xmkhZwWe/ydt1FQbMZJv1BbST+WbZ7Vny9C5NdM
Eydqym9++vjLukM0cGv/IUnhc/6HbU8VTQYNxKqlKLCtI3MqYFeWn/ha6twdd2oqwWziiQjbxcN/
qT44silM3atWllqYYMHP3/S9uAkBUu4DdXn3Msr//kysE4d21N3W3bElTnyMLwdX/drCdQKpNYgb
zLV6wKP7OKJlOzouo4BFe+kvph/Ul0SN4rp10rWOVM2u6dspi/iZTe+QEr0/FTJAZkSG43kYNrho
ADIbEwAPad9uHUtpxEEuLABLHAHAfAbN9K78G0PRxcSnIyp6Z3JOKaPAnC4qDMM/XfVpo7qecBRq
33PTLm8kk8MavHrLWLYhViYCeHMPemDEAsgUesR0oOYDQKWZmzz8iDb9jksqQwX5wkUM8znNGqB2
i0fIkJQWbNRDV5X9d5TX+YN0Rd44LsQvM6AcuDtzfigMYS1sCDFroR2kQyrX/pZQaJ275wu884KT
r+XdzriqDiMxJ8N7dFd1mkYiVqFPjEbUa+2E4lGGCiNFqwr3rCyrLkhCqJkSXROUSkqu5bJTdmbv
qT04St7NPmFOjltXap3nBzYXsO/fvTyvQ6XpwnRFofrG7KzRU79nhBm6MBYIu9CfQBdMvApJPno3
NhhBtpFOqPssl9v928xoWRCtN+pnFmIoLXFh1MgPcYntD+ClQ/YqLrst8ngtS7S63WwhV2RfrfC4
i4/LC8BefAZR439B8oK4LmYzg/W5YEO+KEpU6TBgdBNFcE2Xj6W9O3dp8+ouU/tcaPsSiT0JN7s/
GX2SMVTMcVIC/fxMzmE4+MuI46X8GIVoMY7WnmJmdSi4ppmzD437wRnjDgrATXm7UAGBPexWuN4F
3MFpG3FgXRkkg1duTT5YlcV7ltzd7Ap579kE0G0FGqJxFt2WX4gmLfn/DX+jquYrPknETwFaVV4+
8FlBRBo0QgJzBqsWfN/FQnDTXnTjrXzuWxw4MfqQPtoSgeaxgOpL9ytj0oXmrW603Vq8NGKCDUIK
XHSHXqL1AgMY1NrbAXRS234NH0IeUU622qI6WYC9l954jxWCFAdbxPC24vB5LlzrmFX/Hh0KJGLs
rLHy05gzslBT0Z89LnLoCGtGTZ4V9KvKRyfEW3ls0LxmX/Y7UQEsky8/PozRdvwcPHCXWyOaK/ir
WRUCbc+E5bt0A8UrXDYmQD356Q0x/Xa7pShajTs+549C5v4Pk+qQXHE7xMJqHw2qw7qlmt4LaSGW
aMr3vbqIEhnQWNUsIqj8ETKDasp0GR1k0+nslRHo8A/TfEm6niyHpLjkd0OfJIvln1nF4GV0cs/b
/Q91oS4I7XnVeUGcyM1GoPv+g9JQde/W28xoKWf76zluQNeVvjoU1acRSvSoMGlfvo7xGe5vZ+WH
6VoS3+GBIgjiz1sGgzeflwDUUjrEHtfsXE84z03hZp1wUSqlZI4XAgPA0GRu0wgkPyCGz4dar796
8yp6hFXFpqlJbCVYqIppS5NW4pOz2KtsmrQPn+6ZAphpDVIZobEo0W8cW4dqnBOLVX6F7xVdNaeX
u9Nycb88Y7ZiJh1v3lX6GLwIW3/kCki7PO+CHBQAa41e7X2tExAkPXIUPVHxbOrxfdavJRyYU2NY
xB+/5NSUSUUvXfXh9S1H1KSt5I7ejAtmFWzQndJTqtta93QZhLSobhJd0NCGBZUHIvFsFFxP8Efo
/l1J/C0lnLCZjWFr4iZJwKbuRFnA5UktNRVoHtXLoZMsx38q1ur9rR5XiEWyLEgf2eKeXSMGzs6Q
v2n1E/JmWyCefRgvl7dN1LV7PxJZY8U5AhTW/Gvu4uac7EfPkI7dQLMZ1Clr4uciagMee1Qys4Yr
3OrBgouJJWY+y2Vfv5nd33gUtCR68DOKAEgRiUCCsMWlda/rRAW45TQ/W65oSvV7xMttNVjSzEsL
t2ApuIRExLYfhEdEF7ouPuC9g2OZN/4+fA5+Z8bI4DMWpCoCYIRjpjP95+WyTM8aoCBA7vpKEwFJ
zgQ7U9u4hh8A8jLjD99uE1zIbTqK9HW0agM+RIe3/sxAeg7v04qEbE4W4csGlNuH0FLRNl0C55O5
sK4Td4doLx2SuOpq2Zrdm4EbcAthw2HIqz3t91hrB6MNP8SfWDrS1Cw16Wy4MW5x+1hwj0btkmr3
7Mdr6x8RC6XBtSZrKH2i2R9h5epgbpVDS1b2Tz5syUlDesxovp2wz87ZDwIK0B5LeaAbx0EMlvx8
qVFVbmeAtGrCTOsgHtekAL8jte9xBEShOmqAVzHEnXyLNQHIX94gLx2xlg9iPb8w4Tl0414rZwEs
BO2gO26VjL3pzlHo2ax3MDN9c8zhhaspNJGk/T87q9rwLddLMB9Y/PR/rTjZr+Pc0yJaCrwJ1vb9
WS2Nhj77PwKoZp0jPJO4qaYOIWli96TNxAKmjm4zuJzyGwcrHWut86yvxhj6jEi5BYmuTl0GpTZr
+Z4KavM7sJUrNlsmSHUQlEp2LQT7ksxYIjGAtI3i+JI72HF1E/o6Npxo9Xfsq67dN6i2tAX/F8Dm
kAFxlaa15beD2yJmo1RBYPJV9s2yt3a43o5OC667jEZHN92BLlskf67RUo2M9mFo5l2FMpuF79Ov
JbG+Lasxzindj+WXNOlbTCQ+LcS8+wXfTvzzUFkAGSYh8ZwbjFrsOkphGKVDk/h+sQvKFKw2pLFW
C6gJLa1LCB4uprTnWqKKC8BnPDUpB9+62YDa6t+JyF4P7wTKLPvTuWBOej7vNSvVYoluukolTHaz
seflsqdcYDeUJFYhmQuU+hVNpLQ+o6Gwl6So13yR+9yUCqX3T/J2SMQ3B6O99Qk8qWDC+QpI6rk6
HHvZjFUeAbK8lGgc2AU35IZLDT5GiiC3PRUKCRFzMNlTRrSGLNMtOcy+Q3LiuI7TrUv1qkEXDKlk
9P3p6UZMxmJjaB313ry41h273Hs5H/Gs+wGrm+BaC2cfjPNHPHZ0sqPYb6H6fQOjoDkMDL9TXS70
b9Scukh/rEc+xHHIBF9DNxtPVRXF2qGVZihu/05adjqj/Qf3PFKJtFxaoNdCXQZHVXcbrmWH0Zb9
OYf8q01cohdAz2f/GqMraTkst2suoKyURADfXIVaoNrfM/yO0sf+cxk6n8QsN1ZbqNWXfk9ICTwV
nvI0G6pCoNgT3/WXIZYfUgbOgcaZoGEXzVrJXc3MljfaynME1B5G9FaCHraUwoqKXtzVSW004HqB
ff7yXW4f6wByyYL3e9U1y5eykEMkjwaNhA3sIeEE+9z1lfVelaeIty7BeIoefcA93TwPhnqAoF1M
CUMV3t17AtfZMyOYy3AaR96WK+7jhc/DeGIrdVzyof7G92vA4VwF1KqMu9OfnsU62r0wv2n+dy8X
b8rvhCrabRhQgXe1RTjp8lBlDPkVOkAXY+rJGROsPqp0iNPe2ZMSEPWNNDtr4jEUIG/mTDb63vKR
mu5TnWtLdG1bXY3rVHwyv4HfzestAuKKEVDCjXiQeOvEX3lghS9qN/PSpysS7LlBIBlMQ5ii0R4g
lSE2EuAJdT/kTghuGvkezb2qVXHEMhdVgF+3TIi0FBCaUPyeVR0j0SF/w8cvOyOiphrK22DkUg8s
pSsUz/JGZmAWCdKLFS8rcyj4GrvP22Il0ewXv3GqWsG+gLVT2e4y+LHDL0VcVc/eayXmUS6JBFLH
UylVMaJ039MTs4KfnK1/cNm3PB2zmxOJlWqLVkQ4iMiM33D/3EhVM/d2J1XkrnDib3SOQwe8iYkZ
/2gNBqCA+QmQGWlCFQ9g3XdKTfcZj99QNwnqWN8MEYncz+RdGtaweZfXjZ7FTDYbsvpZNOsxv2gg
G7ZRXmCS1Yuol9uDI6Cxux3tqQCi4E+bL6OmEsWCbxCO5ixuwpgYNzOm6cdxIOHnIPHsRihj108o
7mpem5zfoP5T5Lu5XTmYiZwf9SvI9zwT+mKYL9zEXib7nhr3SD17AZDTOT+92xMiP/uh7vRT2Vtc
/S3WX/gkZdigk8CvfXHaYBN5ENb6N2xllqrAY8i19X3FHH5eoj4PQ/w+umneg12dVTSVo1IBzF7P
rqlKiwikHftO4NaiVyGa5IUj11p8kiDVWF4OBdNT2wB22R3XFQLxYiazyHT0SUy55+t/oikrNEBe
NUapAUhugXI4EiGpMQUaa80uGL1W/gGYZd/M02lb6p2GKSaLXAJQ3E18amvtrE0EpMbw231sKDtd
RPCeJevUT1a3Xlx1VNpbkO9LK2MJqCzmj94ArOgFE0UASLUE+R5eq4lx2s241H6lv5c0ZFuacmrE
DuQDaHV2w6NMq71ld+p4+4rMIhfIaFCtnP7xGYlLHPDObNQA8rimR/U/EeuHPorb41++RVbUlvMr
uvrOOVia4lXe4fxOLcqGzO3Qgeih7iXx/Xvni82bIjEKh4/TM95q8zQ0liMTa29gSFcyB9P5WPj+
qW18QlU7uIAnBnmG/wY58zvobS+gglBNAnnn2Pa0Vra8mpv+Asokw8Y1p0TZYTV8CyC3RvMHIQaH
NPGntraJNeiRv4FlUia6cegqZ7JKxyRufEteUwPijkbkNJqzrC6uwqyGhhQBDmq06PoCESF1VbyY
6NnDNntFZMqBQQPSmzYbWz71KhIcVrO511DVlz/Qezlkoy79QaD9YuGqyJ3HMopQGnCX5HGuij+R
FTMNTjO2QLkjzAnFhJ2dGvZWYF4dChJbxJshMkXSIFL4plqtL222nJPLeBJr5Voyzwqj+QHw8Y31
i7Ofky3XamAn8NDLzQA9RdgVuq9t4UQFqG7ZstzuOR/sEx8ozFDa3HDLkrs77ZUhYj7NfNO4Efnj
RGxK15TO/ypAdxNw6g++H4oNKa2NtNdevLhtGWOAA3ALH3EhrrARmUhHOMHFT98k2pcgAeHFcFKE
q7eekzsYGxbvUMqptnyA5UpqSDkB7loLhtFbIpsVKYu1n/8NfEFW3dNHkmtvSW3jJy8qpo8cMjc0
i4XzYGoco1XoZ9mKWl/2oqH/iETk+5j5VQA3tZGxUcf4JrzBin22H2vF3BKyWzJbaCk4KZqRdR1r
C9JSGfQg87vBy90XDIxwXLrT9LKAXiHSo3WhljHoqll3Kk8Y82LjIjw+JuMgttcKxq6CtDUp3Mnp
NSUX79cMQHigdY4Bq0Q4F7pk55Y52of8iy68LYdSVm7F2KKJtChrSThx8yrOQGmxmi9aHa5SEpDd
C4M2+r9I9B6GJZCWyHevKzdpdOcQobh4U/ycOxWjhlFWuUWVyA28xVE7WMH+Snmi+/xq6hoAAdrR
gfv4Ly907N2nOOFzmlBxTDC23yGFe+MDsDqh7/uFx+V0lHrlWAtfWSo7RYoJeUBHx/B0+DlVcugG
0EmCt3id0rhT0iqha9PReKA1nzD/zHpHXL10LDoww9XLwI+3PaoEVrRvQRkTvBwlJgIuO4UVF0w8
W4AG2GmOag2474rJRig/yIvmRdRrs9X09MlKdrFyq/coETC+rDsLgC3/uL6b2ZK5oHccditNII+Q
FZGCWil9v8wtIrYUehbJLJgWhxIMtL6MEFWDXWRaJKaz6tyo2I2VCCN4fy35J9mAoqzs4kT+Q+0q
DjkjOeSVTwMiK9ivL0fL35OzpfesCc7UQTB0zCuY7NnkmmbnFWnPkgBGETbWFO+7E10EdPDYzQPm
I7JOORIQgiFdOYUFHjvhT5Nf2eRrjh2OJCrEbkw/iAePtzIp+v7lbrNN1Pw4MtL+Xi58ITQTeWPj
mISH9ydc6diGwKXr88Bc6fQ6CIU8wiMzqFYhPUb1tMG70h635GkOx7emqbo+8jAomGR84h1n9FMR
BCFIPxNVMgJeg33ziuNsE762VVuVCTHIrfTgnUmzg+1dBKJ7IPovPI+/9hUpgqbpuh1WHaKgg+7n
2UrBKANcPxtmx3Pv+36FR3+eScGIx1+lzUcUkGs7vvsvDeutplOxHnubfpArr4bsqW26SZhSlynl
oq31P9kw9eXIoo+M0qUdv/eICF636aujH/q6yNEo/oCOqFhIgwHajOAAU+JYDIbPKftAJ6r0iaMG
0BY8E53xHSZMGoCuvzWPUuN+tonPqfh+PxpvqFoAmuJl3snBNYG3IKZ1cqhGulkySuXkzSupZQI+
9vwf1GHWB068JLMjPvPioksM6zFTynZxwjuVsWJC9JmNktIzGTHrH5s5p7Y86aak7E97z2UOU52K
JIP6jouRB7M9FDroLGh7Dwc7TPiyDaRev3JY2rwcQPT9aXEOEEWyYUx62JmchZIuvfM3BMr7IEdw
iGRrolVmwqp5onyuE5w7BD4o9G8frQklDQ6JrjXNYlgADVa6HovgXFEfxN/gwRia5U8vhRWSsYax
CAPLrhN1vihuN7iGTgv036QVw6v5TDYgCnLR1yji/w8HnrhFyca6DoDGxzMdoSU4bMEmkRxWHyb+
EVhL7a412kHQ6Us/9hOYrHOdsqub+zb+3bVS225VMqn26N8jLoBtNX8vRnClB2HlNrONa1L7ISlV
epx1XJLf7PQgC/dKXWjkbDlgprZtInich23IazmWjVRWzaki3FZJdB+LyFdJh0z7kLPTs7LBu2wy
QWHggwhgQoYMATWaTVSsIbSiz6RoK94JYikM9lXF4kEW5UeolVuXTYtqUiNZHvIQ+oDeXJ6KbUeL
fgu491Oy0d3hcZHzkpQgPK0WMKiOiMwGP3RnTT9c9UYpWTT/PjbPaKZLwGxP+piOQ2QZweC4+0+e
G2GXZc3TugmwZi5MBAQTpLAZQo3zqRmFZu+ZoveZzmLJEiKnlJxc1+8GLcPxOCS1IdqjcRo2hkQE
Y24zxeNPWDHniJEwqMWAWAtLui2Vz5SGZ5lFuugwEhdzWnzpN2EMzTBgnPRkS3tci1IDsbnXNDhR
B6wlGXs98l769aKaRKromVubFug+54vVKjSiuc9AtQ+fDwzmaCLp4O5NjuRwQHYfZ+2NaT0o4y+I
tDVcySWiN1YQ3CgH27WVf3FawEvq2bUOgqYERWbGVBEFIZSOnmHZJK05JaMYB18512d8JvBOyYQM
fjK7o0dOoh9dqyRNMRyNTTH8JKtjmBMeWcPrLyrkdc+kAW+mzTIft6AN6uReINZs3GktYT4XEQ2R
X3day71FjcgKb2kWL3x2H5GotsSrou6thPs9XLh99TMzE4Da718q/RSLcupWcoilrUoN/NaA/VKz
LBejHO5GDDMIHjF1HG7PLa/K7aJtgF3tlPjjliHkB/3J2QvLe23RC2YDNkNFtEzOtOtm784UZ58B
zPaun8hdB0QjKl+bN6yUMX6cO6J4DqV/uaMq1OSEm3aW87+5/EOtBDD5bzQuKb4P/5g+8A28/U61
aSX853YQW2BGsQJ6mjMP02KQvbq3/qV05FtQAYoolEsUqsA9RYka9z10ZN5za/kVxSAlKN35rQ0I
XtDEC0eXC3Udtab8jvli+m0GWxLWMI8sZ1ufIMD6zI2y9TguCwWT7wbI+MuUEnvNZpTIQYk8T4js
5mEGvGSQThw9t29dLPjJd/27NJcROattL0e90CvY5LpXNYM0Y4xDlL7NOCd2ek2bVHbA4PwNWFUk
BSMfHz0ovUJKaZw8os2UWJzTWCcm/sRQ1uYdCBQi0O5PX5058GbG+2pQYkk/pXgmwHHwcHuxwIhU
4+IyFDH4w16Yyd0+RDZVekiGKqPpM3+KiTx3ImoPBBfCI3jgJsrIXPeOH4GxClR46EXBxr62kjFf
1fp9/GGeDF0cAK5XwX6pAJbwf9zUJxL58ApJBviovlmrb0DiocMLaeleqkOtPSseyrMibJeHGQhT
GjeX1r5xuP21AEdhlioog6xPPXS6njUcuvjzjnPeVQS1aVK7YHQ8wkkXUwiEHX2KSyuF8TYQIqJX
pQHHSR5v1z+sacv395z9mg9rA5YP3G5VjpxERuUmfoRIIT3+SW0q78CtAkB18pBxqhR+Lq8cRxTv
Sw/yf2IJSH+hmujFAl1WDqiXlPByYRet1HTYyVekdHF1bpw8JQP3Qp17ymVvduXUcsrEq60pP16n
dTIgs5JsKREY9KZKidRBxGp97qxEJhsgxh+3GyHDGRzze9erikKFRJR6ws/cO/eQ01SZwaHCJ9VZ
vlVmxuw7ke+GXc6plHjnuvglMKEh3ABNjgqDrbGY0KJ4kXdPZrtgtAL4xRRfpY/Z+hABfTKDUhM1
G8ud0mzhHI3XdUXbB4QybjhtwZAYtzgW8AkIu+hQagJLeg2hrXbopFjMv3jtaGSQgKuihubqlU5n
u74VQ1+xh27dz5cKIB8Hj3fsjZ587BC6cn6Gby0vWFQ4x4A8jPTD2HqN+s1GqENArQuLOlJ6DIel
23dD7MS+aGSUocrpiuTnAxwFGFENO2qLVdHwfnfKjumYzMMgr86+q5m73GkiiC+/Etg6rJTMm0X5
USiLM4JAdc8OOBpL/DgbRBm0l7QwSw7fUvP3/Fh4XhWsZXyx8FDsob4YoMNUX5m3ZzLDwb/+n353
RHJ/VQbBDbrgrZi/sfvsebz2DiihG9Py1SuZduTr+zeXKYSit5pFC4VJ1eKRk7iDvvAC/RkEs/yF
01FfJY0u7ut95x5i3XVBlGlTT7hRVY0lBdkzeP5dWetdhy57T6B6ZYSZiAEOmQU3RSaV7haAdiHG
rdyVUKMum9h1qJb8SXSuBMUXxWKyqmQ24buX5F+LtrxYkvn9Yxyf0VtjUvsz7fwSdIT6pgNcpp/M
pFnTFHxJ3FB1yiw4gkslPZ4ke658k3EQhuyV3yYg43y85GUzapwcDHoqoBB1h76Kx7Gy7M1KFXgv
oBSuQme8m1XKZcQrTvaxdR4tfDU1JAmdWLU0/tC9p9GTiS7/jMzhxFWTc1KJ1GxMYLm1APgnLUeK
+3/o39GrZTOwmRYw6QORLsNOhLqutqhx7236134EpLn5W529DUyoNK3jLxg7EevlAlHAXJ6aUGae
JrBkx6tyn+0wv7Nd4eW9/e85S3gE5ISXVU3PwzMdM+CHaiRWxbz5fOqq+gYFrUlIU+84vxOAlkff
UaT32ibdsPCcePRqKY34ynMskrqseHQblTLdvx47KDOsB4A391naW37FJMp/wt1AKwCKqEyxZIk/
x8BwFtNyTSLuL721bYudebisXpSdFG1JpwvNk2P/58yjAo0duTwyAsAJaohtjmQNgmoLeHrnC2xC
0XZow6Ni2/CcZs4nsd93MQfPOKXpLF+VAnScA5SC0mNoNLQtznhcQqLwR9Qcz+WP8N2ck9QcP0O4
cRd30fjPOCoadr0035g5PBNW3beVMdPom6MC0VIV5gko6oHPSYNj5Yn7dtPP/CErtQUyYTf4j/lK
4b17JBePDTaH/K9BYtayC0TfyJpBEd19hQGG1r5EqunOSmoJw/URFVqISityCNoec92L1uq+naQD
aiqbJ0Ie5h3i0YTbZljO2dnIuKTMTl7MICqBcuX5WC5pLDV0iyx61KK0/0PuL6rILiMI3ntEnuAx
NFezzn9NPGhW69JI6Wj7MYSlGa3YS5rS2ZqqV7dS0HvUktTpvcjGDD4c34RqLYgG+SamDc5FybBD
YmN9g6wOwe2NsvoVKcIStxktg8HFXwH73hyGly2MNnuJNlmCH7+xHFbYsfPXmCqomDYaRn0NBdjR
aux2eLj4PlTvXxS6QTbWPzoOoqdIRH2XOT3FPamz3OYCm9BA8GvxfbGDpvQvw+M1vaR6PLwFKoRg
3+BLWVE6nUeMBaPVoAo6Wrdj4DJeff8GRvreXcA9Eh0S3mQkkNGdFqIUH+UuqsdBzYR8QiPi28bP
J2uAG8XYCmBocdal665twniUJhNon5RC92e0730e5k4jKERWIBatQ2tzpGCOBijni5wU/qmKL1Zu
G73IYnyak0XTiITkQUQssmCLJIS/h7zOQ8v0T4hiOqEdpyWI61q5Jy6dKNahGoEk4jMRhhIYMoLw
pTKguWGRTwPCn3DgtAEx5/RbSTDr+K/qMFfe1G4e1SQ8uCFG7H+gYzHOyHY4PPPVJRU21RjkHvt9
rhoHMTxyWbtQndev3c+pmBjLiYNwm/K6zZBlP6t/PKQuqFrjK3GCSM2R0fMUVTj22PA4i6HRbPCT
XNBZWKnqQ33sC14nahx/w9JWPOTtsGXXS2KLGv/woZRXYPlwdPYv/ZSDFCOxLuJXEk+b9ddPCZeU
HAB+u3kOwbTCStm+TwzFfYdjVETBjG4VPYDPkLh10XX8pf/aCiuRR/WbLgFB8EVZCc+U+dRPNE+g
b+Tnv11sHeyjvDNOwHpWyMHy+yAlvoDYdzgKAAuS53U7XB7TpD2QC/xc0fD0m1Gt0nJw5QZiybLy
MKs/V+VA4Qd8nsNe9qv2FTYatajOvQgKlXLM3eig7UNPqqHsenzQOCNper1lOhBXnJQWaas8c3oW
N6kr1WG30GojaGPpNXeE5iUhP1sKplB7r6Y39Lr2O2xwuGtaopbem8T61ENF6zUmFYWS3uPz98+9
BQnsPvl5kxTSPBQmBCtTRy4tc4QvhypNgRqzdNheYD+Ir/YFwdPrFJRuD8FSr02grHKT2ps4H6CV
Sl1M9cxSsgs3b/HjUw6tTseF1xDQcNOk14a0rJ19UMFKNIbDDKg5zYAEuDErrm77ZDxpyC7wLfEQ
g3VrSBJC6wmHPx3fE+kZ3ccWMVr9gDUSMl4TT9Zoddt8/De8rxSiNUGQWygg2cVFxtrk4kcE/bxP
/VISZMIzUDCGHjCo/ZMf1bmjH1r+b2SEg1OdXerNj4bPGDrNa2Ma9iN4Cdm5bnoAOYN3c5I3v8db
jw3pRzeYDlLHEG5tbU9meMd3uD/ZBwkiIb55q+UtdaumwDYmikd3D6EPrcOwDwM6wUiEzaoHHMvd
moRFtJdQl6aoEmypyi/lTrN6JfwhBE2kwhxQ54JcUcrEDe4wipOCnd+4Hvh6nitz6E6COUV9DIyG
qL5+eehMAtd+LyrjOeN7Xx7JNgj7M4oktdDcR6AFYWlxdnFZ4WWCI29zqqz+r24FrozyBvqGOY7h
iVTXpWfXlMXadXFO2Og46YyEjGfKQ8OmrwKNTRQOEd5qmYr5RHrWXAEo06ouNUmUTkZczEKF61gD
bZtRPS7+jvpaz6XwH5aZp3hISLMNrK44gmEcWGB1J3mXpCVbc6yw17IxoTfRNNLy9shoH3WRGsf6
lXPkwwgp0nfDldgLMWHdgccioIldS3SL7/oNuO4+bG5FS0oOvh8vJJq7oji0SiVfm7uIbPbSCBms
oNaeaPMsp2EfiuN8XZ/lvCxp9+hmmc3JEUHgdirtTgpcRbs9rOf1TjUWSSAF961D+SDmx67zcPCr
MF7RvomHQNz97pt8292jk7m1TYCgRMWiUMGB4MqWuobfCX0a8V7JpqDmfHW/AlXM9G/B8AN7ortM
qLJe+tr0Cl/jJvPMzNgUcsY4+gU6BjG8BzbCip/qI75msTFqZgBXXII22ALpJRJVHzjrzzE1PsFP
XBPbdOUgdxZs57hNxtb3t40lwhlRBR/OP468wlJWkG6+dylATaS3P6oOiy+EPSHPYCNHURu9JIl3
10E+4f9OiYe9JpOlFYJtYgXjJw+l8tTbPZhdca/wZtV9GWd+NO5tdkqhmdJT9ohNpt1pCDbha54Y
8kRAnUYK/BKgU5o6Gz2LJFmO/Dn8O5Ph7H4arwAoVvSV9e/XulSYgPASzT+GxPGxHzWOKKkwTh3I
WMdGbuBDzO/a0W77QL7x/HzV6wMrWp0DLAO1hkBK+ZirfZ8fD2O9+jfUC1RqK86Gp7/YAZ0nLBdO
xc+X3ITIISYju6fUkmSBevLwOPHPmFq2KT5T3iDDRnCbgiqSEad6jMQJsvfwZ2dxWM9LD8mP0U+D
LvrLAvfs2enlsed8c7nABMLjMXsPp0+v3XpvwUeonxi3GEVd2pMPipjiMbjFeVCZTr0gcUqPKnkQ
fHyS3CipRRw5GUCJf6LOS7GTAVkF+vXtnpK8TVOhQd5JqHvBN3rkDsDLiHxCLroud7Z6eXJ916a7
5yoot621hseJeXopUlwFUKqS2IzacVc2tzRowpfiUP6pVn3XpSXksGjcxN8fBLpFkV4YObWAGb7k
xwxXfKgndqcJu36533SVKUoKE/LpMCVuDI+FxtHW1JjdUcIfOvEhYoJFJlmypVcJJkW9TSfjgr9c
NTGXcMR1wIQCHw556IX58PnErr5ItPN/Pq8R8lUZHgkahVfw7rJosDmYCNbGL4D7aP9XH/cNj1ew
TSuU/4j4+TO74+esgPGJDLDxa3PUYRzFsj1n3EFgqibOAP3MYGAEmCX/0Lpwwq1Uexj+/JfUXXVx
4Pc3JF5FbgLZUB+aArhkghdnJCouFGveHyd6+Noy1M/DftAeAkmIdZdY/D/lecxe/bXrugttvn+b
rTs3c6Aco64JdRRE3//Ft7yBmX+D8Jk1J2hl/CNjPmE7ZbD7ZF8boUeTcoo7Ge+/n5vrc9JVP/hM
zCFBIEM0zO95sI39d1wdFYQpRdx8a8WUxFYL4KlK+W4f65MdOnaeK73+sxUNP5ndegKRSBXtSE9r
wEcfd1P/3yn9xl+q9Km2tR9O166xbdH8FKUeviLqUQioTYiGwJCdeptnr2QlKS26bGf1Mmfi6ShN
sL90YI29J38HleNz7tmxdewAPr8YZNC5erRx9KppBZ8uyVdnkJwnIOT3fK04AzOYOAlk06WgI+E9
1MOIutRWtTbKsm1k5qvmjaboHqxcMOczyJhahIQnBle24Cdamqi4fR3lGP9d2EhaPmlKLTkvxARp
LnHK01oOe/6O/ahnBD8FwfFH7BzBLv/JywLrPUi4bl3nRc6oDUV8QFIrKFyBt79s6J3KIa6cS6Q5
ErqFlQNCZaxBO4m7MVAmr/C/VUQfDPPTxN/oUrigUP04nesuKL7ho1LT+R9V6GZ9GOtzn1JUOZpZ
v/KbPW6Pe62MZhh5xDa+dmdMRbLwGDzbCSkQVNzfQSPNR8/dM34tbI7cFHblACOfSF0xjcq0MjgR
SWkaV1qL3Qv7aBOtXK15gDyP/Q8zfEKWW+WdttsXVqHUIlv7WouKBK7/hq1FIAhoPwO3tDwQWI0/
3ZO1LT1gmZlubOt/tCTMWhCoR7/RkGKc8+evFQPvjdQjymtMg09Sg8q+IyE88CMrPPk0J3sOhRXc
MOJIAGYiiIBdzFzEv3226u8p/gTWfZpEURPEiOSvrBUKZhWYOK7oYN0QJ1ZtYVsmWNoS/C5snrWD
T/G1vUFy/BatW1y3gqYotRCV6e1N3Uyqz18aDM7ngCB5JkqU5mPRdl5CNC6Tb71NeXK3Xkb0+6aW
jK/eUhXFTDyKxwY4wb/eK90xo7M6lSZR1gOSm35bRa+qWQqjuq6KkqZpEbZYu80Ay8KKcFmW3nlv
YYgpnm3QM72k+FjHmdzpiLA4iZVIvrzJ9w23xvXtDBDfTxliDAdEU+OTPmEZBSIFDlqDaXGXs1xZ
sY540lMxhXGQUHmI/aMPs5a8t1bbrmZy6Yty/LOTlLcYjNIJxlZjqCn9w8a7AmzevZLKSEwBg7vc
u46pnfy8ggwvV3s/MWBv3vxPvaXUmOimnsn78I/2Is7PLVVM1468lQMWUrxwLXVRWN3BSWNNhclU
N1JOCXMuJ+OnbOhqJWm5Lut/7M5gkJVZsjeodqOmc6Uo4JjbNH7YXjsJb+fxLW0TN+mJW+IqZ1zg
d09IDEYAqtEbfjBENBdnt0OawDqeV4xk5g89zpYkODf2s+6AYifwOtXQUzLvMmDQzF4jr4Rv3rI/
WwZjz9KNTtnjNQjYPWETyFdRfGxld4tc7vyjBmL1/j6mk+7vWcpV6Gv+iVdY8erDI4fCgz+qVUzY
y2GnZNhXHJ/xrG6r17kEkcB6ARSHFkucIarQY+88S+vQM6TeV5vF6omv+PQSIDcLRnNHJp4TsKY8
bkNx+SlxuxH9dAa0uBIniux7SoiizNGigt32VkiDBh6D2edMMDY57Eg7sW4a1tJlXxkm5lfIWIco
MhYREzNOrYbuLPzs9ngw2jDo+veFYht3ft2k9VVbpXAD3nRGo/4xmCKSemywrEBCBQ3wJ2MLvVKV
O8g89JsB4FkbuZXbE/BLs7WTFRWxAxwheK7LToA3THo3K75csQlxMcImns6VFIfyUNspSYYf/8Bo
Lrzq1JbQBeaYLmcaegwBXa4uDWZ/eIh/g1p6FTNHLCEMZZRs9g/95pAkrEKIqpP9GCb9gbMAiXE/
NFcFFUvCpxO61bt5xFGnNBc+SYfohaVkeInccQR0Ylp7AR9++JqPOCFyGr4jMXvcirCECvdoouvg
dbLaN1EBFBfDunbMhn+JXrGja6SiGWAZm15Q6fisLFn/CVPMXE56qCZ8gEuEHtTtOZEq2ImWuN0O
awgKjFZyolbmmOti18qLsb3h1BayYkFBjYeXYJX5j2QAsdZ97D6xSoZIw6kRlV+rJR4+Wbix72Zu
+upi7K2ANTlEGTIVzDxJ7WOkp9ZWMH/cie2T3l+cawDbnDii8PSqYdqXdXBZyy0up3G1JHaMswsT
FRHNfPTmQ18w1C37OEEmX2YRiN66MoEe8Q6M0YeWOJoJp/03bTZDU9YiNK29QiJENgSmTinjhgaa
LKsxwzerQ5EuvGKg4cmSUGE6k8T8tHEJVMtwST89xkaHVuR/k5YJnIGTDGXF9F0SjYvKc6U4jmvu
KVL3CJTsJkvUGRRaCQNeOeZwyFeKMa02dBePcYNhJVhYt+g2btK/eop+WvxFB9Yq/5dGcmh1zdO3
AzBWqD6dOO4L3Y7qyFdtiElaxFG1gU9I4q0wMf4OU2IbuZF8zjRyJYvSfpCVmEV3svFmAFV9rUw2
TotF3f6Bxr5C8W4I8LZCPWsCRRaT5+c6U+b+Wc1jOnQCXjOLhXqZUYiSsprmIa4JPKxCDwlGBeGq
Nwucs57QppYwQTCvlzNVLhFVgUQQVbdmaW8aOTpBQWCqGl/J0wtCcq9Vn4kIRT6Xa5igpr16bXx+
ANia8dgTU5ljAW1eArYHePGOYgT34CAqfvk8egKLPJQwBnK9d+oe8STsd/SuTEFicbnRGs3srLXP
uwLukxjsWuusv9ATNEpzmj0MvobouGVFJ+jg18VutmvQIRV6AjtHRYC1VqMVVvfy8dX0mldLpcG1
yzx7638T+E+cMK3/ToSGXI9ydUF2njHRUAIfMNlHx4gx2Z5SGOWFeze+hXf4azeVdncBx2byEr/u
8Ltawq8jx2DUtRX7JPIUahLgqSZvIepvKeOc2uCHIdo1tFbvhUJ3AT77+t4K5pSjjN+llrnwCFsl
JhIF4TEqt7dLCNHNyEswOT7r3tiLA1hLLika4JGP1Vr/ApmN45gAQ6pg5OPiZ0xy1XGkKfUwZnAD
tadcwbHPABL8BMlCMFPRY1j/HBILIgrqfx+BT4xnh2YxLLMjm210UrHxDiYpE397mCxZCcM+7xQj
fNGHZEndNjpBxWVNzfuJkOOfwNKjEmOqIJ6zQERA425hpQfvduYy9b8CT0vUGoqw4LYgB3ZlazH9
pHd/soSFr78x3uGB8/AEHTUCEIKt7WNre7jRiMNnj60fMlthvudMCuaz5h+X1G7+/gFhSOj0GsW4
hV45xkH000DJxz4ghrKYWwYxhgtPKxK13XckdFC5rkpLhITr7mc7bMDhLutXSv/KFsieccd5JrzX
sOsOoCmk8JnSBirjXr1PSnMQ3ohNHhbLtDP9OQF5dcd3TBKfnzPEnG2ONTnMxGFfR9tMidhda7mc
12HRLd8TmXUswUo61aQAT4os1RLaAbySYPZlF+irUb+MCg3ifjykMUHnhK+WcggjdOA0lk5PA09K
ladpRKGUnNOZABRCIUni4qBRD3Vw4Psuym5yf+4IKT8OvSaO43fHegZQ54rwCwTyn7skIZ/QZPWP
Q3gvSZPZKHrLgayHfSlpzHwEFiGSHpRpWG/npq+dPOkbAe4Q8vN7WQxngAw24cvg04N9gAp8OMHy
KEqXDQ930UNcF/m1O1TNln4gOly9gaEdQq0h2+kifAspmGGGalaMzODk2TMZa4Y9D3S0NoVsfEWV
HqYJSxutGCUtiDjcyrmitQGpAWwZ/cFXqoIw7lfAHbMswWNCdkIBVEf9czXAsgqQRGM7smOxZmi0
LeMqkV7VsTyrjSRy3amUpgV3QJzJ65u3E3arN3OtgwL86+8ChTgEdM8EKiE5qX6/67ypNZxdlm7I
tujess43HpsyWmQ/P6MMYu3oVfsdCm8y7gTZakIY+eJGFnSCaeMiQ2VUDrI+OE4xKv5fx9gNq0BV
36hktpJ/NSoAMNFdPr0NVqO9GfrUcOx0tMBAX/BHa1NSLbzqEJK2yor4+IvmlapyNVc6mJDB7MSP
F1UBEBG6l9o83vMUisZUmss6l/N7h2fx4fYvGC438+GHNq4/EYEW4sQxx6+4FM4+q956WsXZyzq9
NKBD5JhusQQZLvcF52RuMjqgLPtS8MK3V0dvrG3l8k6RhhgGfjlxRQpI4Zdm8gKYn+LXCpBzu/HT
KIYM7QFn0Okk9jLcEzQTe+n9rNs2+BV2E6n1SOj6vU5HHuGgwDLeVptKGRBRdIb9NP+jA8yWEhIB
oXXvJixYedu80+a4Wu9wKmL8M+B53Rh7N0/koBf6zODGCxk1wuUBDUOhNmg/alxAbxFdNIeWsR2C
UtNlg1ABbfH5WhEvkcQO8NvYZMXE7X11ka0FeNjSALxrJffCX9xQVyAilm8hpN7ozw5cBbfdvP/s
yeM9tvMhCWjj0lXj+FVfEvi3QB2JcirGG3URkSE5+y4D6PL6UmLpZW2623sGpp5cxeBrPdtCw8W3
kw0vgXs9bYNqFmlQ1mkTA9X44zb2rdeYEGzBiblkb9kpmwVXROrC+Y/T3V5gE6a7l/m0k9ylDZoM
+ngVZVIKWymPLFqrAKNRKQb25TIEh4R2Ym4LdUueYgoNMPE5bQiS1f80TniNmgh1DOH8R8TnMmIe
RAZ6oPtN5RhjsUwpLZezAvweFxuLnBFtFumS1mMkmx9CQEV28ildi4Y3L1aKoxEdsYg+ck8TWRh5
X9vIS3qqC8fByai9Q0F2TYH7untmNjipatRqeFCypQJoPz/nYvgwjjC2rrAO9/kYfnqfBiGt+iIx
qImYk4oW0Xoz8Tl2tKO5B8GlQTGRaU1H7rjilgf1SlHxqpayeYnSWZQeUvbORvdw8rFfucDAR0Mi
KTWUGoeHM//k7+2u8KDr7t3YAWOk+SsbBSTCpdDfMnHoB2RxraAkv6Eu021+WNEp1SeedCDGuqGd
2o5DsZIsyrPjWR00dpgRvaaZCDjnQfpOXuc63kheEtwvVP+jA6rvBj0ICTlpD3Cp7pkEd5oCoROP
w7zesDAR0ERZhYUL0guepgntXQp2b9Ix76FrJv9IxAM7cC2rptp4o7ZSJVG9GDotxD2fP45PT3Cs
g9sreDtJNANyejDJaDXKDYrZRhgtP20I4jeG5lmDVGIKODGOuCzbO6lhG6NtU7qlH9wXKRyZvfZq
cF2jjZtoCO28OkHCbkeZer3KpjHg1+3qpB06aP43rAwbFZydBLtVW+thca1zKTfwQ1pyc9VbULZr
6ovvxUX98+iwst4t8sZ9zRi6+ig2/OyQBJXHUwOhuJgt97R11AYqx2sqgq9mizB/00g99lVXBWlA
zMm/1T122UU9L3ha8IsDCDIWXzHK1ajYVijIhOnDkTFFe8OF5hLN/KF20T4PZIo2TDn8ATMVYVUC
whTpveBgyAE58JPZIr64BUNDCxtnb9EZk4RUZyYUFH//dER7Xn3CEIZzTVwhYwkmFMHUIFgwu7ie
q0tk+8kq//PXizrWUvEIr6+yawmadYiIHomGXTfTN1Nkswol7hBK61fbA95kTJt8DJne5f20OqUe
2V1FdIEeOPDGQl5EIYFn4OdcfCna67Xd7uf3rcau1T7GjyMuydOSbeIguNVYustd2/GGxo7TlOdi
4IblX5L+IeZTTSYottHYL1igXftxcV3T1VF7BNakxrJxG1EqxiWXrH5xvyFfbcLnHsGo64mUR/9R
6bu9QxyH54/leMmDsRZLjTqF3F1VD3tRYmdpBG6aQIur8sv1KhHUMNZCK45oxtZmmNaBDEtThAjB
njew58UycUkHk1qlqtC8WiMNkFeqcjcA/QDpuCc30RrghQ+tU4eWyGKeYrABbQrBgU9CXVs03ByA
3XVXk/7pt3Us2XpCsw6IIhuZgyseYKJFRs5Ktxi/oBSNDb8JiHYppAZzn6zLMoByvsDF+bewcqc9
/zgenynntNK6t5wPgmIuS0pFFNNs7GTHOQpHOnoAu1tYB+8Rpx2PJfibSPdQu+K6bFhHGq7Bz4/q
edUOkmxYvNT3CTYLKieDXSn6zMH8+LOg80mIWaNlmzqqyed8RJtDCCPEIfZ4jIOBb5E+6B6x/Lfw
HxDXB02x2ANBKO2s/URzsQuX0YtB8w7WGjaeHefCuqQ8ag6IfsuA0iRsXjDTN1EkAlvKqkmxcmuj
9xUZOeOTxNSo6godaAT+RxezdCYsbq8TezEtLlCJPncFb5UA8L4ePSsKCtvt579uvrST3TyW1J/2
YfGk6qtGz4nQ4o+1YqQFhMH5xrPv7ubtbY05iXqM/mKW8ixBYb1PqlnHDoZoYe5pIrLcWLwxF+Vr
KeGgAtPeUIuyusD9nsGPC/GGwVPI+kE4ANm1YxcwPqwrMPrYIlVG4AElEF4BdxKLZ4LOgHDzxuIm
URrNDwb6WgsV7rXzCLim5XcuARcMGMg2dEM6ef2ex2shyPK6YfzzlWzsH/ZTo+BlvJ53/baz+g0G
Ty0rmWLikM1OkoSII4lAC7jsQqFdXU7iBNQjmduz2LaNm5BVZ8OgPeq3XPxij3rYPXn53VlYFeUf
GYiqMsCg4Vas9tyOOCUhwt9ujNU5dm8/xgEVUXCDymPVtM6etm65lGPeeM/VHw13YkaTXl6DPfdZ
t2bVqF52HvJdyMgkJZU2R4LdnQFIL+xg+u4X4AlgcabXaP35vCBHOBUKDnCdKIEhcTqUh/gMkQWM
wuLb30n+qoiRw1YDKyz5NfnGT6gvCa4zJxoIKOCHb+trjEWpYfW23ZVpUMXo1J48mVxhGOi+SESl
3ZfSkzxd/VhVwAlkyf9QcEstGknQSiusQ8hc9eiPIBoDq3L3DcqQxi0nWvjK+lYVdwiIs1QKBJT0
zL9KH2J/bprbkCHWakUO2wXMyX8RQch6KHlo5WL/eh535Edx45mtatlRluqB7rrWJHBYAQx1Na+h
LFOGTE/002PMKAgjuLG8gSYW5wdSwjMvxk8Mtik8mzFpkALj96ayaixNsmy4rp/3PTLp9+PQZUEK
59KxalvJR9RoW58Q7rrW3yrTqGoaGLFx2LYNyOYcsZoUtv7GIQOyqBugzJ6iTDVS5ScZA/s9gDpS
nXpCnTMRKTtVeIw2W7ghGDVaJGCYyGdwZjD6FZAobWLC6UEqk1Avqz8BOte/sA7yzU9cc7IeTmpA
87aGeMQiJkSaV0F/VWE01K83MGVvxzacSBDBSvt/NYbN0pe3t6ByywGNZlJjZVXpuokkp1nZsIyu
Fi0//X22jPcutIhR3T1rK2s60FFyjmMdr4F5tknAHs9kSVtw+pNX3jfjq2xWkDz/5vZa8TqBwsud
e2DmbqhB2VJ6lzd7OBwJP2+UTtOgbTM/oynQjhjNZYDp/JkoWsZW8TT8vJba6lOaK9RjzNyrYeAu
TveOTuCbwvJfsxkDJm8SkJj9/YHrvp97l4oKUX+3yDxEyrhkdZVoJSRaxw+KMOJJ9J5O3HF/Tfe6
spzjxU1SEIc+75jaCy3LPA21RCyVuc0tVFN7beur1oY1qLTHAfmYP/zrMuf5wTQy5cNGwJg7dSTA
FyzcDngR3WcoT2k/okIxLN5VulnMWEogyl3SQFYjgYrszPVMjAS2XmITdJccyRORNZ/nBOpxjPFB
vtv4XQemkLGoF9BkbFwYQnGP+hPaNI0/yPaQoFIaagJ3CsSbisLqWW4uK280Qb7SZ1GT7FoFZE+f
5mBe3TvgrdPc410LC+cmCxB7M2ZlFlx//w/xIfPDWWfnl6OBbW8l/tKnL2n0qqkLRpVrNASzrnMV
ycMQ3OtTfP5VqivhJGIs6+o0GWFUsDO5z40QuCtvGdrdhBY/vIYbNEiRz1Zf+Q08MB0DbZ6/ZoaZ
9DrrzMi0lf0ijUHjNLIEtlgHyytyPD/Y2NUG/8juXtevIT0DV+PnFo3UvI4pQdJmI7x9kwKudz4a
ylBUt/a7qZhNChDCmk134UoroAsQvpSJS/Xzh76mFFM53vSLTcGxNfNswLFL/4qH5gOSdFMnhnba
oDWK0SrUBfXD8zm7N14I9MpxPgmWQgTAW40KTnAdFVGvTwxcueGDk6ivrTkPnrGg8/7NIX6BT+ej
1moWqpcxn8EWAyfJw+Q/mmEigkV4r0G+zksaDipOKy7uK6wD1RgF34l7i8fFDmDHGuHM8k0MW1MA
ThSIK8/BcxiE7cZDouySmrhf0cmKP7rp1RGrVRKaXQzlGMM8gYzfqinN05E34tLzvQf5Lw4jPWh8
Cc3MWWh+JCoZQDH414TP8HyB9rKfeIdAKRCo0+QF9Ql8LyQe8cb0eeiBKzpdeRD2d9l74VaduLsQ
LblTRpCv+DJA9zQxqivjEPzBKvilqFMCgYGOqhopPf0vqYzPV35TyStkMoazUjfP7gw/zoLeZb1N
85gFrahXo2A7r6v97gEH6ra28g2WalIMCO//hslOeGzOBr0h3sPfBmE4+38dQ1y5M5vNJZBjbhn3
Pd0bLALzn3nOjlwQAyocCI/zXPRS/1s+kOw4eyBHP/RYVZus5C+ndepzZEw4Qs2R6kGfpdRmVHYa
3afXWurWxRI62b1s/FgcejWO7JXF705ultfTFpjORdi6PjMLBq+5ymPwqKGPH9gYBqturDBA9KP0
EtxJEcnoXi66F7ferpwtKMRXJPTxoHJd5LXv7zBGp8zJMWsxqnT162dgNGY1G9QVQC46JmSv6fRy
35a508eoCMoxTOjbO8s8lQhAeAIsli+PUiNXZt1PJFci3EMC0vk3PoC4+Njk+KY9HnmMXYEMcMq1
s2luhp8lNRM0S238V8uwuKIBtj+dknL1EkS5NxmlMLF6ELw/26DN2qBI9o6T/wzVeAk7Z65kMfD/
4U9W4tbUtBYgoJDpbY4PC7LK7g4yeq0+oVvvxfiucXN5bXhKfgCjfUEhQOr76V73XEg0tZn9qzqO
lUM/dNvFP7726AzboyqOVFA1rjG/zU+bVAoHFg0i4rqafU8lw59Rb8pkbLaWP9IYi3/4aB9Y7C/3
DgriLQoSByPXf70BudOazeJeRu5uNDk4TgpaT9HGWnXyxRCRfx+xyRD5N+ueN++Tdwe7MJkqtZVr
goimGBw/rcdipQMT1ieaoymL5bZBes8tUVgvDtuFll6NWuMUWcKDqdOiD8vqMcWYb0W42jLXRa5i
LOhKfxbihjzRb/C6hHqMqOFsLFZnvJS/Xh6j0qaOgCDpJ7J6vKZuLjqObw9wcCOY3dmVoA+Hu3Xf
Dk7gPhX3QC1z6JxDwGCmwgNTFDQrht5LVl9f9e5Vk1L0k7xb2xPegHLyK1nsBuGmORJ7NetzbfrR
62V3FZK3t6U3Iob9/QUqa3jwJBtDuy9Ua530Mwvr80zOhbJAOlqpVUbMAB7rVpy4b+X+Mqmf815M
MbzVXzDQ1u1eM9vMljQVARw7AUlZAMnoKwewbXEThZpogce7FVh35Hli9id1kbKnRh+lNoTrbo6a
bfzO9qnTz0Hcre4bgM4padynEzcaT0+/7kNfftxhqjDNCKInIdnAodRGVbTDDW/Yaep/VQfagLEG
rwXtQuFrESA8BgfbFKHrGhyiR8Ne6OJIGLQcH3v/XaCL4l+98f7VmvT+0v0frKrOyQpW/BcxPbMu
d5q2elmZppKtikAPDhVTf52zMXGH5H80DHCm8SIQJRcHR8Vc6CdIJf1FY0/OHW384+jB75IZbnRt
AAhmvbugCkOBvDi/1M7vDWPnZ0VJWSJqRB/VbdzscbqShbN/k0CAaY7f2WB4RsGgYY2lKdbGfSto
JDwAgMUzZhJapd3U0YX6hF576zHBrzQLN6KIt/XjniSvPnMY68KM2wXdP/SMHPMFXRVNVqxts+B8
MAtm3tBd7QRZyB1vE8P5z1V1VVbf/sDf0sEwEBBBb4hr9cEI31vLMKGn46vTGLa5EjmnGqlRdzkH
pYU9kh07Njj4meT1FFkFNh+CxNqdt4Q9xwaaetJR/iCXYEaxNwHwH7zVv2o+/6zN49L5TES5BzBr
b0P9PdhwMqI8RcoJaReK5IJxk6OTJyhXauvpi7WxDMZaGntMEpLfUnSbdF0Mja+w1EQJ/Zv+nFQa
nvLJz7bfAE5Sd+17H9Yu6NtMyjb0yQtCnefgGZfuRQZYcq3eOThjEn5OsO8lLcIZU4HcMycDNxLx
hmThqPmT5L7JHRXEBz8LqcPLHsyXcoc9d8u9Icj0OQ2bLlc0WerXaNe6gJS/1MeL7kxi7g1ESvov
K+saloGg4wz/aPKrEGgE2CABJwNHUY6HON/aufYWSRQRXak3q3CGwSTBn1MdSqo2NBlv4Iaplb+e
XsllZ4jQNeftnb6CxLrxEoEwwnlhBaY/1dP2V9GsL/wW5ek1i0mQLE+uhF1tp1Fb0DGP/t3pz4zT
MfgV+NR0GT5ndAcpuTSRyeQwteqcqf5BbvA0SlxZkrhFZ7ub+9n6suAYVM+L6m5GOPni+1L3LNjw
0nfZF1kfwzxSPxpORBIvmS/G+gdFCDX9fiXC14LnEuNeWAwsX1CF8yXMDPvrW95jboAbErqqUGnJ
RSEGBGBFanSNCtfGk6wdpT1nUP51hsBD7ZgdmueosoKxegf4W4xCSS/O75Srpiw5vEOoCpfXrD3s
LNqfrDjIneGxWbyhj6W3Vsjs6dkxRSft7IpUDm3EGTlPR4qylLij4cOkV+kHVsQsOgeaLOPazjLq
e7RUby0seWKUMmGBTICqlyJ3KnLSW9gV5zSM7pkojXHBliiPWSkL1CGKUvYRUolVg0l0W5K5mWcu
J5zFzi3Q/jWR9f6h75U/3dm2oc0H6UKLLqNEIbGyr025MApZXyJBfzRpozj22c2dt6gIlw4VR8Ss
BEK27Afn+GvuDDsi8bFwlqYW79OJmcT5SSTaHVs2RhRSPwwjLLug7pgKUuAFuVaWKypF6XPQ3qhc
fkbiE1NoKltlQjRCVyhvgqYZOWbe+q6WYbZ7Vn+yL8g/2Eig7r9RhktSbLcGAM/bGtHWOZSlgJrf
MANk8T6/TXZe6r1H2DbpbSOWNe4LKq9QNT6jB2gzC7mQXEwuJFS2FL/vapeRyAFmGteQyQSQtRKu
NIbG79NP+gN2MNswT44/SQkRD5xBAa/YPRBxZwQaK7E8NVwCtG1LEfAAAQTksPGqcvsmd61XRcgX
U/oclrMH5VMJJJ0sJaIXXDihwqhyCPDBWQO3pravXsmcbBdCBhXyAQT/T+kEA0x+irQfbc7nQBEC
WLkmREj6t1YutObuGH9x87ahq2PhKmozpqLqdCA2LloNhPeZLtUkpW/e4MmjY6AH0ZIr4tA37ODa
9CxP6XYQ84YdHEJzGUB7bdilxu9lj60qQ5OB9oKOg1iDeOgwoL3l7YaG7ncuGyYJoS7cMGVLFdYE
HGr1QDxftwU2XOaFXXxqCs1UQFsx4Jp31a1onf25svn6K+4IKdtLcnd8Ash/L32AjpDnwwN9yC01
c5qUVcPPqHM5Dqf1gfS53lK6FedDEfM8fe+xcOIcY16krRzvBDh7+7i02iwztzvAhDaPm+M0h/Y9
YGQbf9upsFTB4fQaZ8wixVWYN/ZyBO43ktYo0FQ+fw0cbQEdhdz13NW+42w+gZk5YaNg7yprpCtn
GjDbCY77r1oBBSOAFXM4jCBwsO2G5DQB5RxupyTssGBBdh/4o+HrySFu82yzNf+3WVGt0gEpGJkd
/aag841Y1Onrz/qLjlX7YsNUKuoGQxe579Jujgjz+UEnweTg8Swdt7IrH/hRt6GLsXEll5teBEaL
L9vVt4DnKHZ5qqJRiwk0ZctER+J+0N1fx2OfcKQQ9HG4p3tmz7PAqNw2XfxTLdAztYsDQeQe/GL+
nHJgnl99iEE38VE1gqheF0t05vvVF8WK8jYlmkKdx5UKaY6+5WcHoxXhwRs2sMFJ7C5Ijx4R1u6s
mnWW1+wHkbYwnm4rnE6DFMvy4LTfNwOdAyHnUmEpJ4zx5+W2lfpgiFOjATI3jhjkMconmWd5Y5sx
sv/C2TdoVHPt+S9m0n9++Tu5sxsNtDbutjOjdzlY0yuEuQNYsVRMmh5tLD+aJup3I9cEJJAbulaD
Mpqd84TJ9ciW+z1zuLollv1SR6oVA3/F1sVoVt+iq9EbNRwqZTCXTpPM/EqziV+FPavA/KztNEm0
c6OHAEv+x3a6N1yGNz9qJcoZfbLaERjEyRntxxw+cLf5W1M1+VdRT3XBNa09xJVlRsqrL/5bv3K/
jcJ/rYLs/uZAFFB/vYlw5nSXQ3IeKxkkXFIyHda8AFxeyFxxPlxwexLc44+DJoWoZcHB/V7d/MQC
6lerYKvW1SFrfk+DmVXvujVaD/SpAcgbORh8jgjOiwjuqVzZlx6BN1jHNQAc2Z3dsAtBECXDFn55
O+yJ8ZmCIogelMN6d0V3jCe5cm5HxRz3OOyht53LfWnxJIxUlcM8BNtHzldOFr8R9pg1kqrtt4PJ
2+A0RZOuZpeE1/CfPMoy0I4ejgNYsID0H5hCYGgsj4qMC36LY7vy592vDP6fnAMJ0IFkn2gx/Uad
VkONUJOIEJLEyPZNxjZZOY9sjXAm7P+tQ+KHiSXTDyiyz+KS/8oULltDg1HT82S7XcybIUU+0wJX
vp3AyuzJ2UJlyWxUwSwldD98djkyxDdVR+s33GZkVlpjRuuQen83Zn00mQBaY8sJRrMKxfE3Sa1z
JbWarhyrXEcsMUpDm2FLurIs5gGBXXerRDpAkZeg7CmvHL7rw9tCHbo7Q1GjIkEO+gHlQXawSilX
uSNmo5qAJCtfPXfmdRPpJmPLyZ55D+KZ1d7eA4piV1im+E1mgrECGv89hIF0y8epUUWuKU3qODnE
8QQnJQK1nT7A/vspypujVU2rB6DLfQj9vJeVy/cTv2GTBF5Ads4m1lzUwpvpV/dJcYiqsMDH8puc
iMKDld4UTunVPQ1F9wLfr2x7zVRzJArKeX2guKN+S+kaTCTeIX8ZuwMeFN7zZHm46X6mwr8b/HYa
MyZRzfsYYPZumUyMLNbyq0FzUzgJmsX7pVb7Mr7t28LIix6z9H+OoJasI9WgcgruXbnynUkPSDpH
RMKSCwXVjY7ga86gJdkIJRPwvHNT9yFbyJaDSUleDdkBOU6GicCoi5HhHXNOSPmzFg9IZsPj0Nxt
QM8lS1zpbW3wDvbT8xvFZGcMVzo7oAHI273subZyKakFnFWj/VeQUIOjiUdMyZ07Koxn5NBXTexu
nP8YCMr/JQRBotHLJktH/mRBPHmMH4iXLWaZ0AGkGzvCecEDvUWB7uyrFI8Ol9XZ8wnU35Jjeymw
k+zlr0/oFrNr4GO+y1Hn3CdtEbuEOSZ9lAKDKADeeFqksPTFb85SvnwsL6BzqS8XIaCmaVNiNkpl
AlBdzmpTcK0mfNB+uEsNyqrZtrjvTVP46ggYEj8+4UByAJLoWQL94rdcfglLo393tznT+L8jTnrE
i54ZtobClCIGWm7dO2i6HL8eQXBHvwdW+NtwAMDCpf2Bu1/KFmCvXYIRNQWhh7fhFm5lq4sOXpgs
u+usUs7hmJyT2Uucx9bU5846ToTgQqlps0YHi1TRe4D740nFvFnOhM0NlqYuDsDQo12njNi2ygbq
4M2aT3Xm4EmV6PP894lBbcrRp1ksL4vi8xYaFWzvbi31o/ARz0cOd6m0NxWwtKlEtiagZMxKru/0
4K6RPrlDrdTn9FBh2M+dH4Iq5eXL907PcouJHBaNdxmVcXXcXGobP4jU7vSDXv+LNmjO6fVMr6Vn
Kgdms/9CLXYStz7yiga2rcrZl6sqGHEWt7R+tsnGQIfFmT1UbXe55ulm6d0GkWhD/ZiGXZ4ZTT7C
qFMahTzqcYYxN7xMb7Zl7zmAW6kqsygq+Ap5FP40vGaJ9EgvURJgx4IsWNMiPXN+0iEmZqBQk1VW
i5yC6ZagERfaNo/DeIEUAeagD6bUCdShXOrxOTUJhzHhexOfoRLJscqzNcQ0ckcNAXysJm6k0lmb
4l1Ekt9sqKSljuMG4rBbIg/3ozEboES/b/f+x0yovXlt/UeEzyRC9lNW441mo2quJ2SOBc0arvR3
y+RgqmQgmx0l+en9DnJ7im7hpfpMFL+tzT08lPD/k8Pn42wjsMUQWNiP0ugeS206umaVF9SdAjPA
AoyjcxJrL7nJ4iAcPHM3itPbcZd85j7y2L5vX6uGrENoXfrb4JxwYT7MI/pgSYM7LFW7l+8dyVTv
aBdVFgRkVCFLTiJgtFpZoLbnOI5DfetC8DSDQZb0bjkJTFkN3xWOIzNzB0FJjIyds36ZtKV3NrZW
wuZWX3XKNRsdP58eJelzPOZFe932oIYsyYs0I0LvyIHXa5dyxqCabLzAXQNyOgLHR9ymqv3xdizO
HpGgHDSb0JDyqJOLdlbRB20y2AL/bz+G6yfo+eB4ypmnCHtTfrv70SJM5A4q2Vf5MiHEhMBprara
g3QEmVs+aEA1Oii2iskzu+iWwvn8vFqzoks5z3vlsssuWwbsLe9M7/QxnsUQvuOmarR0lNL9dykl
2Z+wOW3nMvYNdXT68o/YN7peRktwAHJEoGbTiNzAcaF392LmxuATqLT6BbHMhYSXATdVPG1XLSuw
rKHyApqSi4lZbUFOyzjAe+RwyN4UjcmO27+qXXKof+PIELPTahymJF/JW+qOPijmP6bNAWuTnX4w
mjWXcSXfxqZS0RcfWPvo7Ze2VZiRfjj3MSdYwgLqpoLkc2BaS2iGtRi8ZbLS+R4vxLAP4Dx1KXtw
5dNXxLfmqtpHdFI0c8vqUIxcbb+ebfeOx5h+qRyEA5AUOHBpUrKAEf5F3WJiLY7DcUTX8lKQhjtu
ragitZ5Wjkhaw5naEfniH/puEBLlLGL+XhSDl+qCqxa8tgckALhPuuvSGd5o04QENILcVysiCOSP
EBPTXuaEeMOXvmpf9365jpgM/9/GalXls07M8Aev1SkyjOkJwOWaCO7thfgIseTtCQ2Ecx+hcntx
eaXLd6Fr1oFsKPOmRAq5mItOPogAYTajiYiVPuXK5ehJN3Ko5Js6ZnYu5m9qzvvpVxxxtYF3Zqj8
xBbhfLGfYs8PpcwvlTpO2KbK8YFE1TZksDt6rIEtwdoBGJWFjYzDsiQj/MWdSJMGk7FBjGjhpzaV
N5MBmIKmM8oP1ILohcnWIeKOFU+1bIoK3I3Z3CVCIzVvfAfe7zCSw88MjTxsHJj9SPj0wjTO23Sv
JO9PflZMuy63DLR6SqRgJ8AHT+303ultA2m5/cvIQjKP2gUz0VIhgqo3kqpvggpJE0BA1sN8LEzi
2x/W7+rQQUkgX0ka8+y+XC0OFTLUoQhGyKpCcp3vRRXeLIBhS0ex0pskjsiALRyth6EWywRGS3a8
nO081+sbw6tOkGU8L3IheTqgf5rspXaRyr1lDYvluesGXUHbv6odfZ9VUwuQ+jKGJcjvO9YI4tCa
vfWsIzo+ISUuzRA4FNgSGutAEne/Qd8iyL90Zd+/Df7yY+dRlt788Muwit+OaLdxHdcOnwzFelJK
Z8ZkWX9I6gCpS/LZMeZhWWW0fa3eDH6OTDUhjFkxum2bwcuKbg/2cYRIsDJjtoudzp83JFnQ8PQ6
RdDL5inxDeMe9Op3NAVkI2YUttfD/W73OOqZ1+kjj7yVU4Y5ASOQuZnuUMgKnE02e4JEs3MpoqcF
dh1O0rRHc7mYIKwytg+iOwf6PHk5m4Spuvdck2fyxjrcynG2FGkY7I3xX8bXh7QVfAkn91ESnU7m
FwcDdys3INXG5RrUv86u9rVNZyFebFm3btXnv3i+/ZzOi4vFaLrEdg3z+GecNXRlHPEZEHoTSJeu
gP29OQTQbHHFWGdIOsoH1Mfa68tAHngXytJ/4rHw7l5mHXadqKpOYvm6kz7ljtK05HuBFn9yVCZO
EFp+l6JmoFYLogzVHtmo4dkzuI4QFWW6VImXDYTF/WyMhM+umNYbx69ugzPlQSj4PxkKGyguXZF9
qW9S5Zytaf7Em4xLnY83BkZ8NefFgT4r3vv4usRbrLkZ7hZpgYtQ2rKOV5+e8f4fs9jCgzlL87Om
yoExQ4Is5hwF3y/TtxnPWp5Jawb5HdP22wW70b/cQJacdsYqqBaNKEWQFJBjeVtbt0nqqW0f7Tbc
+RRiw4IE5LCq1ToyTlanvx1BPMDOs77ezMwKB1CHjF3mnhe7XAstJBJad8PUeES1OKFfyOruXdC4
PRd2cHQMTzJEK/Rk6k5wcLBtQ/fhQqGXlzddZoHbvlFMwgnNFgicChXMpxnT6PnExWRum08708hk
m4PYSTQ8yRKS1pDcB1cKWvYsJtwa4SNqKBYvGVNsDKTzEkBGV3ccj0UhYs+usIkJFamfocEjj2Y/
wfdNKvG125K+cw5DooFm/aIqYjeQEHZZaOCstPhTGBlnIMpeDbtTa3rFldOuw4fy7pnmot558GjE
+X3zVaTYmtvmLPW5Pi8B8ofLMRsEvf/OX6YAKp9QDXpJcV+396b6KbmFNJ1GFRXVRc8VXqarFswg
1OjaUN7J4EL60E/8tpDsFE8oCxxTbYKjbV85YS+o0gTZqca6EC6M+A6NfWoMc/TkFl/BtufDLwGN
4RBnql/S23qZEKlhSBtGbTnuuui84fH0EJpUztBAxqCxumbe/9EvVMrTAZqFjjw3ZoyLFqZKSR1u
bi8CLHCYLHDbaNCGoF0GsmnCP06kSLwLK/qg33sOsDVez4KN+LB+578PiqxSuDlPljFHO9Fkuf4C
BJyD70yHdyli7L0xrquNQgEzZ6XyxddR8s5mGk5lWFGnkvDUyHHMue9VG4JDExQy24DM1VqlSRyA
6R4p3qfF/4/HWqzGHdoqM9XhBdRUdXSXdDd/GWWsUeo/YWBzTcpCALbSQQ9gDaeKzjn5vktD5hGL
iUYCkXOrVF94quGHb8CjU6r4Zn68lDfocnIEy2Zjin++xJvnPNJKwbclel+ru/PPvfq+A7MNVgVh
IuDCkCluF92jyBT/iVZIdmRiuAhQMuttC85WKmg7W8MF8Y9xmXqxadXCfG8A9I+Y7iSrphV96RDQ
oS9NfgfbPYDJUVkSJqZdjxiULXdDyT3HIIwMTCUTy2YrlTEq+qsh10GxMzkk+/BWWlK6lm6mt9WD
EXYsBeWnH7JOdKTzxzZ6baBvx8ZisNYOQIZe/uqSSE8M0YaC51M/hQtYManvJWMLKp6D7ORObFIb
l0TwhdMJZcLnj2yoIM/RJAPQVw+6WwVeBjcw0Ja8dbRfErXk+zfODn0Js9yLeLs20Tvn3XrlYpRG
rBtcKazrSmPq4oZOpw3H/IlrIWnLIzofIBKr0Rml8BOIvnPI1S/VK+eQrXVyQFxiOyKQVVKBju0e
dWWt9IITcARz43+nRgyPfgN0tT70+23w5bYugsG2bflWC70ivMPLfiBA0Sx2yEZpdkyCHO++0p74
0ilDZEYSEa0hzXQ1Aw5hxXf6048Mm20dgR+BDaI3xFI0jyYOaAPGQCQBEMVwVxsFk0aPCOUAGtYl
YDe/yPpkrmPamJLs9mh1KsJ6UV7m8sO7QKKj4g0Y6x1oJSLK/mIaR9iom89YFxE92wjQKQMifhw8
dRjedq58oST4ajDQgcWKKqRIcZ7ZE87uS4L2X8kBDm8dXIQ5uGE59OS1q832R3zH9WjZlmYHUDqG
Fo4MnmpR9uJGzZBuYdNFLce8+C9WBq/pgL43BYpA5S+JxgoddaRy3CZ4i5pZm+S6v4OQgZmQBDr8
vB8RXwKe0mGogJAlXJNPiUcuZRazdXgz+43cYIYwG6hPGQVakG2B8rnSIf8Yjg4ekWYYFch2h0Y2
duXV/NPQfK5oH2G+VsumulQvG4dUqnkUGPJMkEYf2m6Trd3rR6uNl4zxYFbVn7hNFO7ZlEV5vng3
ZlOm9ZUXLaD+DTOVJUzYJO6ZjOz9dfUz0NOhoQGzfE3bedYSqQkaV4Ek3tB+NudjXZK8QSdZzXdc
0rbMSriv/RdUrWd6ddQDczLKUDAKAB3RerTRhPjrE4pzP1gBPhbrYbAxjMlG6m6zblArzvAJg17N
9rTv4MhTjhxLRlkfEDgvX3LE0A2XqiNNfUo6SP+Ao98+dZ6NpNIEMutbdSpFFvk/3/F8B7cqgoai
SG5uJWuCcj/skCFKWosW8EQkXMqvt2TWeg659tjRSW3JuFUQyT+5mcVnSWapSqDPVq2dewcfXmca
+KWOT6EuKryC3w3yymSEuVT2tVaQBXpCaibXZ+hiYyaD8GzaPBmAQOv++1yEuX+ZeQU0x+mRhadR
x4YcoFUFyIs3smt5tqyc9Bd5D2lKldvZYqi1AeTvm9Yusx3JOQcOAZNOhjwfZe4zFDszCfuzYuuW
KR+fJ7HA3JNZn2SUtKSgB7eIE4c3MMIELcXguxp2BPUp+OlgIhKLR7gSwhHnnY9vJQlY5yYgbmuP
Yxn2LzkRQ3tCdXrpC5kyuRZgLEp3TF1PF2OY2GhW9AgOtY/BwnrRzmhmqjJbhPRr3Zwtv4R8pFPe
Hp1aXpC666JRqrneVn9QXQ3LADPjzm5JBjsA9LJKQHfNfcm5Z7wyIls6R0Q3drTi3EnGdYvFvB9L
bLSwPL3PppBqjT9RLHBm4dhUxFAdOsGKH/+ml4FaBpT+l0GFs6ToQ+Ek1DMW+nnE/pD6+uS1nfAt
YmE+K7RGpcxnsutCvdbMTFdu8tSS8x8gp/xUDcS2rkBAfPG0E4TzvQ93NSJW1gawYW8jxHVkeOBd
uSsjExaY/cghWQ1uYTO02ioKXW/Qp/lZr2T1GqFyRj+QbiCx+urJkGFfsUsomDh1L2doO0jj+nKU
VYwi3tZ+oVH5fuj9Tg6N9aoB9xRagB0puDggwRypcYE604KHEOS6viec0nDeTdJ0RHbjRSnaI1OU
G6sqIoviqUdNp3KkI+2YcsO9y3lB0y5bgP4sPwfWp555wQXwWDafaezBKkUv89aRcBSjRRTgjabW
UCXLAt5FS2lFjbSA0+4CQSiryCRoPlKY7BiXyGUaQDRfUk0LrMCfyIfok8Lu4YsUpwa3Kk7bAZZ3
sHR4uvzH8MoPmPcXGNna1iP5frfI0dCbe8ec1d47VTH2UD3mxH+G6LUeYNk4a1DgE76S0V9syh4o
c8pfMN9iaY6yjCe9bVpjRtK26Q2e1349GorUJ7VbSLToKik8JYUDf5de16+f2eAeCxP2C0Jp3QYG
OMy0UE9jSayrvjoKFreL0FBlROyN9iMRLG8FscpVzujHxNfvTGbWD4JvcTB//PkUkmCED9d0+LUD
KLmh2eRX2mAzjO2iUMle39Gdp+rIvrAP3hc6y04haXmhrga1P/xDb/RNif8ettPONMmByLlMbkWw
4k0DzYpoWDEeiXwanqZ4DgFSLLlGZ+8EKT5b73azkN/IQHKofIcXpWqMb8WIE8YBpajDOAEdK1we
F8u7wHAj/ZdwfQVmUJ2dDS/+doqTMG418Nzk5DFzyqLsA51vQPhbTnHS5S0z2UsRmk6oQcAzXdAL
nEhyYhixrUulwv2EotIw4OKKpQBRF3mR9JXUXC4bcORrshuBS6DR6qyB2LUrUeUJ1PZLNWqjkUAv
K6R51hx0/pWAO948hStIwPouRZLkuBIIOdNcaF2s07xK76gW8rUWMCgkad9IhCYzsTuoeEO6jJuz
Rj/G8eTxsWAw6T5f5INQaSqxewFy/eKgn07GKZFfH0isSq65/5gJgW3d3Gz20JDnT+sUMYoKJKBY
SkkBtX5XNgd8c/xD+Y2QDCxxlcvTsCUKjvxzh0xVLBo75A+WCUp84uP2cLN3SrvfpcobpUOZj3pj
s+cXV98jyBgCDJ3305u/wu63u6ShmEg8TKBDSq6AM3NR1XHlgDTUd4+n+ZKfk0pdYkYf+VUmcZZk
FGlwwup+JXn1NiYG43QlQ3/sJAID7cCJzG73coavYzorSZ3Di/LUG3qQcVlth1lX3wQZTWxi2/2v
Qov7J3YwtMUK3HJ+R+tR/07piR1AGObfW0gn9etOjVSvrQxec/4G3VSrsBBfoOAP70w2JLmf43IY
DqjUgctxl+jU4YLTpDXXWurX+Gf+OomGScLCcNNsiga3B/LY5Ipxp6J9RrW87EaBR5/am25GIWFF
Luu0P8SfPNKwlG/q3VRIwpzH0C3M9rvd5YrvOZ7+81VsR4792rKXC4b/bCFE8nSJVApF3yxTTW0u
UQr7PDm7i9EUw7Xmei0g2lZudUujvkHJLFvUNpOmKKoEExv/cJ8Pz/Z+ueqKuoOeIGaS4vB9qqTU
4/BHX4othfVWPQVESkvmhXSyA3Kr/TbFZB8J0cckfyrAbblz/V+ionP74qVtvgYB7q660bUyRi6i
qTtRDgurhYoZj1ZdfyD5AM1NQg+dDPtvlTyEvh78+5zNVqUrca6pr8aMEhS0y5DgHUPVFjw8hKnj
uImklf5bXl2ec4NsIpwNo8wG6sgmJeQyohI1xuAAotYDhu4vmWZIW7NGWP/SEXX/+wk9v0NibDmo
i1jUEfCqLh9oT8gDSHItWQtMxpZZYIU/J8GKw/qw2C0aqnpsvmieqyY9SOOh0mSy+dG506kHVJmI
Sb+rcoHT3BHQkpq0vQ1o+XEzh79/6LIIIKt06/h9ufiP8NoC+9RWC3IJAj302Ck9MvYrCoHk+dcz
V8v8nTZw971uo5+u4fzuaiVfyqelw/2YCI8dypUZXMAjAMutK6I4h0ehEad9xPN9LexHTiIc0U09
ThXRBWx6W1QLCeDMh+NTVh0poZU3EwtjJ0epINcjTdf9qgK3Bj9QcgJz0in35bi02TLgIoY7xCU9
aHA23dRDVDC8Px2Pu7CUXafzsyA8jcy2/OBktq9GZOENn12+r/9wxZK55lxvdtYdDw+PIQp8RPwR
zDxqvqdL5dSI+KI9OYVKxc6gzNuZ3LPZiRvM5Hl5IeXLDQx0T/gJNyfl2cBNYoUxDSUoT2kK/9A1
VaPZkEvP94CksAtWTl1Wsqu7M3MrPn/TbQiWC3USvnQk6R6N4P1ZtJ3JdzlPVKyqBSodom0dLQd2
pqmpwhkWsJCmC0UL5+TyMaXl3CdsoksD0W9TlJeLRdlLeC5NaQazY1HNoRptiARNNMQiwyZNL2ss
fIIhPxEqBeNDzibdWuw3GmFaQ7TGGYvmXLZ+PgvI4F8nkxQJ7GAHWnL5i9ZprWskzZcRXme/QuBx
Z6qtLr1eGFzYMO882K8xNrouRYWfuL8+5v01VTVEXPyfs6OwDDhTWbES1NeFoqa72KW8zvbwKelU
e2Ra+unw7oUtflL6HsIoPdCNNHq/OSnasTPGdh7oiiutHI0jalf16PT8Nwd4nUQ7n1gGVA0LeQOk
S365MMQGa2UIi+sis9M2WxivXj+Tf5HWPlMp/wdf/LgmSbl0ANiiXE7bBv1Sd7rAC741NUQ8D1No
86arniFxvQEeLB1dUvisJbvrPJf4BVap3YUU9oI/i0fTsyduEZ/WjFy+o/QYcP5OEjomKn0fljrd
ulnhPhoNYf50+frHrMD47jPJnB1oSA1N/ZJgwnjLEF8pLSeKHHKbLMKft2kdZwmEWcHv7LZ5ZkBJ
SbszogAsXH4IrTwK50sBqI5aSHwaEhFcdFLnV3n+MM8lChpHvL7JybVDUBdeWaNmVbMy1KEldFCp
lL/IWsh1qxDqLR5fRhvaZRctDrun29TOKpO2dkAcPSvyJBaQPeyZy6YjyD3H5u9MiwkabEYh97Vo
TsW6Zfx1rj8CvQAYckQXMcZdxrsJBw8k+aOZBp87v08K/aWsmnevhgF2YvgDgpxCQ81gVo9ULDX6
3E0fiAa8HpO3s/mSLfSV+BqbOX9PsOEcYqkfaUCzEyho+Mw63HfVyla6K9SiefWlDyYl/zZD/Vv6
i4+/HZ3v4OwrgVjvlyn1fae7LUIWA1iqxJvuL1n9s+HzB5oxVKPWdY9CzPGbT2hAsGeKu854qZkT
Hyy4dUkwIPo/ezFjOGHfR+NryrhEXumHyDNWgA3X2GIrEBAplNjo0izYyPVJVg3wC4QPOMXwBwbA
moXhXFJGNV8oybsJZtCXgZ35YM4/x0d1lfVqaxT0i2SeLqxA5WVPP1DoJoreNJv0QixAbjxLyQaU
9AI/Xnuk+O5skXiDwOaqVRhbDD3wSBhpi4pv0rHYEUpTiy3QEJu0TuU92HXItSjY0qzQGoUFMKYm
kO1TsMkVJufLEjcaMi79Bj+QzGEpGH4zEPSFTGlCJTooVPfeyJIt0P+4pk35G309FvMlnSUiKMcP
9w/hZ76HetuM7wGTZawCqiwnXqGWXj1hwxDOltr1Py2tB+argutBYcJh2+xjrljcUQLo3+2eXsnt
QNySHRpjV2iAu4yeZIQO8wWdVck5jE4GL2JiQ49kZcArjN2tXccgajGMeCC5JzW+roJ+/yVVEpOD
R+gHJzeDb11RZN9DuGHrLl8/NznZMeqL2DpCDXiT0lB/1q7yNWzX2+2oJoTqXAep+0RS3MWWRl18
2Vm+vauLH2zgjH/99rJJASjUsz1Iq6UEGCSIAVfMqlZDWe/Q1Tiza3fPqDWU2YS9Bjqm0f28sbIB
82F0jLlxLxolZt3P/x2MK4TXtl4gsqWEP+SN9woNkkWtM7QOBikE1HZa1Wi5PmVfci3JsHB1NtVc
SRkDrkjcmSj3E3PLuyvbeTa2+rkkpXk6eZ+HlMOA66E9np3B/5SBxehwHUTatv1p7wSQHARiKcc/
npKLU9X8Y8b/tgnEmU6yY2OgKQP5LjoyoYms992K8lrMBEq66LPQ248njOjuDI4ru5mYeMPPRhAS
uy8DsMTpQr8fbgOqrZFWC+TZcbVVqf6EanWQgjeMnMEt61h7SyuHQjMtfkbHocll1uJz0o/5e/Lw
4aUAgWcbOZK4DfpX5/g9vaUhIOjHgLLmOqPwRzZoQce9xYzRcnZ+eogRwxVkNW01EAyv1SjInuOI
EeQSZ4HXR3jtfuB0o8E159CdkvHNgbHeYKCgWwa7jq7N+gTkHKuhKNS1G6Oa/m9H5uMcQbbndXLf
LZMjPFLzoITgCsk9jnLiq6ago/V9dP8P1s0kBroORNNIw7opwGv5TsEGLqM52jlmRsLgbBiD8zEY
MbNLGwYGYYEzH9NCTTmcK9CaTF3Nzq/ZKjVdUS3FOYMlYdyH2ZySeY5GE/U3+9TZ48Qd3gDkHSBg
zh4Q6VYgA83n4Sx2aBpPnArrin/XeA257L5LDgWaMSa+g/hf++Y07CLou+QuAC4MnJJ3LBVTHJgj
HX4PK8zoxP/+ZPedWkNCj1Edh7FbM5FhyxUzSibkqwY3L16JwWKJ0oR8Oh3L+40fDOwlNl8rU6GD
evPb7WhzALDuf2U2YhwudUdb1noC2ksSK51UUh5lrx4X3r+RMlZdJG92/hwdy8PV5DYN2E4TzcLu
xZ5egNjzTR8P0K0Zthe8GRNrbER64AO2bEpJIu6bWfXm53Vzxcy+f1bKT617fWV6PHcHbRVrFBX0
SVXwbrmjUfu1au8vDYs2JjE8szG205+m9/69eMFm36Iet+PYpHkesNAO5blPINeszklIic694MhI
lpnOy75H3o5gkuVOUZhfpCAc3WwM2JhE9d8ii0BWecFNiOfHpILE/onOzalxyeKdRL3KMc4OcrYx
xnn62Pw7hrqTWzVI4KthUZeAcu14GOBG16OnDs4KkaSldTd+Pu1HUiVXa32uiKL2Tgi0UUOXkPtc
stRXRCJCz3w4rTo5BxoLSKNSudlJ1tjxvdMY8BizLIYs3c5hSDLyhWtcDtRRq6zdCyXUZjqRM1p6
/soSScpeyRtSKAT2ZYKOB8kjyElz2GitsikaKfeJ0McYNUQY1O77cUYOr1ixqgQQwqG5PGfInW+K
Lkbg4p+s1jwyzvuF1aVYcuEYDoXFl4tUd7LXQb7xQShBNGoh150w4OSZc5UIGqxF/pQ9sTrTQr20
uuxSdZhq+1BJQ6HBnonEwzVU5Ir4VejVlKgsB9qYQboTfDc97zGpo/rF5i7NthZn7MZ3q3D0fBAy
gAryuM3JjOqtBMhut8BwUS2yMZkRRxKijUfkoAdce9E3J9b6KxfrGiKxPrXJ4x4i+6weGQ+dmY66
QES1ly52ymZn7TRbxS4IC3CfEvvv629bRCP+/SpTG1wJ2muPj//zyLiL8llw5/h8LY7Yb4LGwg3t
kZMm+aa5TJlhcpVE7TnCwW+39erhlNsJsKShxyzYBaMQYdJhRmWON+QVt7emrkN3D9wwd+betZMp
1Ock0aI9ghOB/13D2mAPNdfNknhRgm2hBUw/VKMUNYc4FA8CHCMHGaJKEBKV2QXWXQnqWDg0SeET
x5Yd+KFOYp7krXAybSLGwqOtSDVqgD9KUq5BjtPJOerCbUpQhjSb26HA5BFFzVsefm8NGiQgdiuN
GxVs+UMHE4MB7M2/Fdv1X1aLB2h12I1aCktUgamuTEIVcruLiIQUzl+MTRgUmULOyOR4vHpVHU/q
74g2d+ERfpWrQWscOy9B6DffGRc5IWko8ZNtEaErPb0G2cgSw+9GXLAPMFOgRnbqbgkI5F6Xcu+a
9x2xPoEFbbqmSbuO+1jerzyl2V+qoGTeH6p94vC6SmBI6pZu8UTTglvelkfF1HKPrdRCQRFkqZrL
uSZpMdSv0XSVGms9L1nA7MnqyAEhKXAZC1FulYYFYnmxvyzrKUnYhHypn6S5XsVg/hpCZ0m8npGm
Viz+W3igsL5GdWWwqbrUJ6LN/7KNqsD+zTHjYy5cXtuPrAmTZakw9AkMYzUY3fadcotq/uW4UJ3E
VuT74LjIuoE7EM/qhQfj4SxQPSzVe8UqwM07gXSMRmWh/ZHC9Pa2+cvoOgyN9UiC80Cczn1TchcE
TqT3bmwTmArN3u+1mIl7kwK0PECMw6K1e1NUgEsGp86M7ddKZnHzB4uUhyIESFGLPcNH7EABOWUV
AZ3EhyemKpY9EuaK+Kr0hbJdfywwWb/q5LAOHkuBzNsOVev8B4Fbgfc6r/yJEUp5ZkeypoR2poPm
YaXmnelBv7pklluWOGecfeKz7PiDq++EKirjgkYDeQiv9oxYoYR6cbIMobFT4v9lOCTJcJ+0F1+B
kyrExa2fDhTt2y9W5H6i5Nzmx88rdbIsPalM6IKDKYni5TDGjzJ87fNwxgqSQP8I7/hJQLOTe8nU
aryImUgP2rBgXiG0hjua+ZueSlWM/qmrcHgS1Y8hG9KlA3Surucl7YfVLXIABdtByr8iw+OJYWfI
Ah2qczDs9zEaLu8mEaM3j7AqU2DF5/aFmUhupcKK8Y4hnJy3IcImYgLv4n2WI93WY5YzSVAthfle
8EFlSlX82AvoERDSavi3C77MpR7liVKXBJ+KVTatEsHXMJlWxOfgUAfEBCvv0CVyez7lktwJSGmW
7Oti3WHeu89Ay3T+OwKNhh4s0NnfFaoW3iI9CKSqLLhnO4L2XJxqSvmLUuONKZenUu8z1B5JMkr9
hrssecXhXkyOwOWxc7nPf2Fsx5pDaWKGQ2nJpdK0QkRT9VGnacBNGUFNpapaOvLEdot8/dS4/2yS
9vO8NK5iOduvU36mQEVTsBX3f3i9n21LNTbszFXe6wLVDzeWX4yvg98+hsrG2zSMLh2jKFIv2tZF
+T5RHQjtjWYFfQUAEI64/nySzXIUxmULNSIbWJp0Eh1RQf0skNdeVl6u/PNQnc75zEmDtCzG/SbM
OSggy8meWTw9x1qNXKASfoqzu/4/UDTBumqv7/FQEUJ+C+kWO2gr6Qy1czFG1yewGfDV1nsqM2z7
bsn3k6Rsb1J3Q2/QksF7FoIWRv15RxWRCh9OUx/g6DjsD7M7reyrsHVN6Uk/i37Ry0ARtChap0Eg
yjId+6Cd+YVsWMtXgk2OBuJKX/wqAW+t9fUnl2cMyNRopD6Jbiam2v6Ec5dK4zzlbzqOMFz7IXXg
k5gq4oakyJN/teysszE3VxsIm1j1Qy9svU1/VXuO0LMwoGqaS4mqNHBeMV+ElLWtMjxYK68JjL5Z
GIKnlqZzo6KIGDsxjnrocSG4M+V6alpwNWmxftfUUH4yLTvwrs38AWIBdwJY1S9XrYoYQL+HCDy5
InnYJ8xABdIplVToHGFSsdn0lt8Tu4NRw1W5SJtEp0Yu5nKqYaZGfEnHtTBocj33cRun4mUeHxhu
0JY7PHnrClYVbINS+YWTBRV9LyNcYixu3vGN4b4u8Dbcfpg2AyES3uB8MvPxKfRkvwmBJ5dcogr+
c7EtJESaifK1fMFDaXusMwKBySJMNuzTSiPfbX9CYVsKZdLYsGHL7WNLDCXj9tXVCyV34nwM+/Gq
4oX42hfhkSAvGz0vgLSVyvLQVm7NMtiTqAl7nEaUmGsGdMZKzCNd73V5pkFL0H2pqOZO7z1jTkbJ
pAIPF/PdXjOdvrY9dHpIJCclbd2xD4dxAOsGxPHJmsWtxaMWvUXOMnZglsDHeCtgIQV4x7NthMO3
ZGOnJz/EODkRBN4EHBSToEhO5S1JxE5Ep3PrQxSlgHfkAQURyJpa+HAvIHJ85dSDqXQeNIZsKF2S
8nroPKZW/nBBIlqpKyvR7HAh6pxoSj9zlTpCxu/onm5nJDf6bzCb/BH8HJmhRxa7ruhQPh+m4nne
0jG7fFP2j2snUIMDOGAmpUYNG+2ySmzrm6q8lml/DOBW0Aqc5gzTdGl0cq0jt/dURM06JIIYgBOb
+xzUhnEA68net2929Xn3QZluNBT514n3yAxOpMV5IKS68vtCimNWKWop8u2kpxSMK9roZP72/L2T
+QvOXhjLLePip+vAPsBDu0kkyNvxI7P4sVUUAzyQpKk0H7rQpImJyvQH6YXJ2UG5/6OHwu+sRitb
+qrMYY7JhCb2gsHHCqy+n4WAESm8knxS5c6mcrCMzmnWSBTJHm3MNntcQEr1D/SrzZJCoBpFZ0i6
x0XrqE0UpDZdY0bmfFLnSXbolMqxZ2nyJOQPtibmXs1TaR0G3PnJbHr6zko6jnTwPo6yG2XhSm9g
zBKJ0HvfaWUs+RuRFa9hh2bkJCOGytxJ+fyX5+ueDFs6B5QPeykeVcQtPOv6tdbIYwLNlMeQtrrc
dIzcAjLsFGR2rN8zGmnLYZN+CmFqqnqglIzdNXWDki7zjMY0ZYaEodM0yJcjpsaEH90s/GhgWYwH
Rlo4ITJS8epfHFIDhfYTr/yoQdoO/S/w2kcPoBhcRiAyG09wfI6nzYVU/ccx04SPYyKDYmow9Vig
fuVxevCx3uYqsZtLdM322B2e8MU6wK4QC2HSeSMSuk3vAElu4ZyHGjUh+74FOgMgd8cEMF5Ofccz
boksS1CczuRFhPEQaOZrqAi4yBB8alvr07U62AaPued1dblCy3qlWCng7WqonxSxm2dPan7IQvfx
HwY23Vt1x9h8s07s2MYE8O5Fqk72N0ZCN8rfAaYfcviY8H10l/HkM+P4DTncMRuNzAf7w+fgKvuB
c3l3A5IWn0VW700xt6K0nDUvKIR7mD5d/hQ9jGxxtrIZ7GjuDwYSn3bwTI6GLN7N7V7tOJOxFoi1
Wcpfy8w5YGTIcWpzS77gAUHIPW3UdIS+FeubGk53bYpEeWAHFdn45EhMN9NfboI1Q6Iz2YMTkZov
nN3iVrCHngO6m2kRDkaT4/HQY3D8OqjpkyhIYNFg0VFgZ+jvAC6/M5Bw52vxHfhpW6pCe9sILUGm
7EImHkxe0oRcaFMYj4L287v1CiX2YsZgff3rzXmXyNwL/7t7kwqr+9uchBkZM6PTRPqCBIbW8ECC
3DBrauA5CGZNEGpcFsUiyEX3UJnMys7z+dHjYgndPx/SNEvddD3nDnmNZoiO3ZN8bTVgFoZgwVwR
+Vkyrs63PlUUEwl7rWVRNrEoTxAhJvPPwjyA05svO96ppx1Qx6Ygy7fYaCUDIauIbEMWVm1s8Lsj
Isa2WLp+AbzLTbJ4UDMz3MdMQeYjlnsl3Eui5k7V+Y2ryBdfVWXysU+lKz53OpGjPC9ralhUhCAK
yZf458+a0R/sHdnWQoTcIMuy6ZugCdby+3lNgw5yFNNe7Ql5dlAWArEzFBLj09FIKZPeLojPUTCL
mkqeoG9HxBy8Shfv3ZhN083Ms153x/SCEGG6ce77HU4XnmChYpwxusmfWnNKvfnTWuspButo0E9H
4RhPNUIdtss2UT2X1WGcupSRKXGM2gIUlS8khDo7bSmouz1/7xmozmKIMDfm2HZz9vMbrjPtd25X
fwYwuHrXzaXEVFkbiKcx4s+/AEQApSwbIEwcFj50POD1vSrBYKnYjQwqnN3cPcSTxA22cyqydkX/
EfUtiqV6D8zzgNwr3DHbH/BAExr+7vqBYvVuTkVn0Hy5YW2OSlyIz4NkORFmEcXYHH8L4qeT17Z6
4Hn6Ug9lJHwN73NTMkLDhKTMuuKemJ41GOWoN8zg7sUHjfetDZlmnWWRjq+lZoThoJezkHPGJiDi
ANePYh+EgGdGfogkzOh03h+BGAg2f4BY9Sfmsd1s00LBlK4m57y/JTwfotvSTRNNeTpI8lBmQ1JL
AiYq6qEDLPq7mhGj3zS+1zEFt+5U6/0otIoBONxBQjzownXXuGHjyfAvkYiqPJPrJfIBat1lqhI+
0eNBlz1+HXYef7VTe4cPKToVnOClTHhlgZbMQ9FkLRIalhldLShg1JlYjqWfSKjgC6bC+2AhApwh
Mhs79+FN/DhAxuTT5knn3dC8Jd6p15lnos/KLUtPyD+4xyMCJE0+SlYv9WYbcMqlni12hOfAcjOW
rLnMPjPNChlEs2Hh31FogGt7wAjhOSVM/gTB25c8nCWFddjOtPapfJzLAPR8m03ZS4bYAMLPUNnE
hTdTnvmH0YoGZIsqM4bI2PciN7s+3yGH5PQvtmuDSZEQfa9ajMN93Pc1vkWo3seG4/vnWRcgH6+j
Gapx1Rylrqt3pkJsXTkV2RBuLws11M7JIN7L3KvkFsgkXDkfrSHCN0xk+yUSImV26aogG2R7KeHi
lApfBTZKpJrCgOL5RBmn9KJ0Ajnf54jc2UoQFBFPuygpXwzh83XUhcH8vy/wHs7CaRcj2tpDo5DH
UKLaes4XdwK5C0Rcz40Rd9stDPBxEYkqG05nFrj/rlR2TMCPaG0LsCkaB3HCd2p1bNs8vz9LDZab
W3MvR2axbv8IGnB/3SSfeK8Ouula5LYE0hKSslUMplSK9nTU+B619k02JMy+6MKi+Vwc7D2gcV/a
djNu9vMAP3zEZ+Qfi1LMCWrKHN4+7JljKS/XTtjTeQsvUDRJilQYL4e8S6ywEnknpzwlm3V+JwXy
8tYjPcvw05FA+iX6ZrC9M24gXgz6fgxfdAjpA4tKYkTxTTjXzj8mxAN/IbIgQ1gjHb7WFHm1oHL2
nwThPOw2nSClCOpg4t9T/3c/CuxOAmXfNhCM8JvJdFX8mOujetIPuKQEXvr3/GyVTt0iQ2BDE4VB
bWopYXRjhkUgptqLbzJbQ1wgn9EwjfXmfjgJp3l2ms03wrvWqnXlFvNhuhECbzSxN0uR4GaP1MKw
ow1s/OQwFzCCfpnrWMI0dPMObVFvhVEynC1rIycC2KxmPuirnRTzwAP4A+9kKG0wD6ltydR/MAYS
BBqtXFzySjkDp8iCJ/zDFzcgpFoHRyzvY2vMF2S9kuJNWYCUvtxScN02uwsFhwpEvoNRbQW4Nx3i
39fxrDhC3cvCCtjOLhEqVuwJrAj7XQQlc9c9mKwmmKSJYuwVZlPItWQc3hmdU+fZztpDsRc/CGFA
i/EGJLlnvDoTCCUqTWdgSrA1ctUTEFf481AqFZ4RDDu0n7A4+vJEcLyUD/j1aw0WLkRBm0fI/lAx
PLolZr8QiyaNN5LJdttaBWt9ihzQOs9U5cm0hKfo6gIyiakg8C8yYSIzvSWYsIaZMuXhvSH907Of
RLSM38uzRkxEWCMt7SCaILyR+7IcoFwh7qpGfQVHFMM5FuKCjaXirUpHw8T44X1H/IDaR6YQJ33S
UXUSpNG0+f7mUK/luearZHfjg+kfqbpT/q24WA4jjRe0N7LidMlGscdZ0uIG4wK8kN27+5rFJ/DN
wI2MBUn45CyfNCsikokl24NWSQ4Qe6Y7RZjNNScYWZp9xTBkOLKhiRXCWIW/RhXDDYJa5r3ms1XG
/847Orxz9WpKFQWd35ZyX+4S2pm4bb+UvnQYwcq9SyEGaBTBC35gMLwhP/pKMi9hf+v4kl696js9
xwprTVTkEUTndSZl83wstfzu6hb4Zt7g6R7mBgIeuD1xxk+//auJVIB4MsFzzUPklUFG9z3nMv93
em7PuMSbhRWgwY0CHI+HlnRdEYWnjxYpANElpCT6H2rR7Gua1O6tgoNwYiARn3s+/R+GuUvB2dPa
fMK0Fb2a5ZV3yfC/7GhseUWzisIJ5jOpU/5xjV2IqgDAW/11PTl/N8fGbiQ/5qn4bi89YGeoGqHH
sUSJS6eGlD05ctrlx9IyD2Mjk2SkZXAkZAZYZkymF6ux0GNEVOTTsM79GZwbwkLmWyjpdvP1Lq+w
uMTRRUIOLJtgceDWqrXBcxexrTGn1oOwuHmMQjxNi/FcUacf3r+Wdyy5O1dt/QdGSJCpcsEUW0Ry
8by9OhAfeqGtHrWs4W0uOSnMKU9/vJNjVWASJulJiwFlp8UCH+2ftS69HXZXRjieZ3pARWhXcm7c
x2dF4QJblk7Zhror/P5djjDGuSvvRnkp5CFXRW0hmONy7N/AeRionkIE/+YOdMmStgLBoSkGVoBy
gvLbnno/sWaE7dIBCfiJL2n94oPkTjbACVzRC+KCNuD7r5x9h7guYd6+XiNBxVU3w32mSkdqP+Km
LCnBvboZDaW0hFw/6R9fE6x/lqS8F4ltUraMgVvi6+qsVkQIbMPaKHQdwtjvNTJXRBTEemdu6VL/
DHyZJfVbaMboBzeLNsjkBVfe/lkryHcCXxrWZmS8gCccLvS5E8Knt/mub7oCgdUrsq2Zg82Gbt9v
fGy/raXSWO48uEVILIzMJUzOll60OUx8yXl66iI2JAVUgP7aIdsIpPQNmhoBP3e1mHmYe5yH2lnM
GDGG93kbtotM/I4jOgZf/8jAFgvJLnedG+lpCrPNQ5K5+BfXWD418pf75RurPqZF0X4kXZcfqLsu
rVwOqei0YkibpIX0LGgF68xOpAnA40VnR7vYMO4LbbY/jDMCXFfeWWOCSYr8lpV1+FnGRamjr7MC
MYJ221xornS1XlJVc5aI8T6Fzay9JM1wO0yGB+Gk08CQiIkKW4n88Q0sm4j2E07ih3tkaibPG5rk
gNYPip+6Q+wqIoIn486UHHw3t9Kd4yFDSAGbX+kcrZc6sytl6hhomFb0QojekwM/XPP8iBhS+zcg
NCtf4RNj7a4B+akG8Jjdi3f5RxMlOXxQZFU/ezUj4/LVL6rm5fcQ8LD5vlGWUQgKu7lms1sPYTr/
nmcm2mElERXkCumthB2a6x+hnLs6afV0vqEWiWS7GOc414FeK2GIqV/3Rn4v71uK/m0zp1mFJlyB
vPoLvddJhaH/eN+mCtzajJXJOAisc7lWS02/l1UAxGYfj1KROqLL/sDeL4YiD/wH+9UpBn8FiM8h
f3e0SZg3jzdMW1O6jJ7tYQjBMBR2dcTrOzf8lZP39WoOTwJBA4UpxXvNp+DmamR7e1BMK2o+1qwk
KwRBNYvMXtahltPCk4GvUpk0rghUCBBsd90Hl65EDLZLwyWwIY2fj/XfrYlw10AFZsShMFI/C69I
0j1tohN7IFBcOsSpvwwyrdyciRBYG1PvSJvjJ21TfP5i86MH3UbTxGYRg7zSD8gtEKoA9S6v8zpR
J2QMe1MRNjEWFLeQRqfkAKOUnjGl5pRuTXla1PtpUcFWPFMrZcoP8M4BQnNRcyw5xXUnCXbL6TRD
WFMSpOykB2I4SZe2WUOahgEDznlUOyB+Q7pcGg9cPlIxNy/fwM2Fv3ERQS1+a5CYeIhr/bEM5nvU
B6OPKRyXz7POjlKQh1wBoVYxEZ+ioD5mx0It2rfdNwBHDzVp7iT92b/cZXE9E0FGeQfuoqn3s8G3
nOt0q/F/1YWgQswIUDQbQJKr+QUR10xoD5dBnSR9DX65zswJyAMlfg+q1jfs5TtPz8wA6grkEv5N
6BziAW4cdaS5O8LKQM+18xkrdx4IKGqHGSc/6npN9xasqLvhM2UDEAkXHYyFAWFzty0t/A8nIqDa
+WWl/mHGV1DJ5OaSZZ1rGyFWuAPGPozk9Wt31RJgoqZ+aUOAJxCPA4N7t4CfwCHS2RB5Qp8s/wg+
kcW2phP7J3Iwv5YOOpfdwv8yp5mQWxVTLao/9Hv3RkBkMdFfOPd1tFUJIEFvkJPFU1rfkG8PQtSc
6RLEOX9TQnXwVDvBw4fG06oqhXyNpdVq1AMKwn0hfEYUxpjcVQ9ViN9qWN4vdiD2SgGmVjLqYIOy
a7rl3u1S/w24eIUIBjZgYHWPMk/LOcZpeBfB/4DHEKGG0Sk2Sy1jIfiMb5TP3fXSLwXF3ZWOVDCD
rla94hDPht45bCkweeImG+6HCa4mGhF9ysXaBvjn/GdhVxWPlin/N21tzaXSKnOsaVdaB7+3tOAB
yfzwNbe2ZoSyqO85ViKFbxOp/QSMyJ0lItZ9I1u9cautVn5NI1xJxO2Z+coew94GlSq5TDVr/6Co
jhP9aRP74QwnhNMsQ6+98Jq5HpJPU7SGwLbiSvKaHw0G7I3zWLoWyQEb16VKUebZCD02tgdDJvun
sxaCapjv2Oh7oaUBcyZIlEqUn+02OGL6pxwG9AVvXe1LiFnqxc+rNcyROhzcLSiHPSzw/2LX6jdc
P6GBUxXISi1+W6UAbk+6DEX5EuUVnt35SQD8OLx6Zw+Cwg/AUlfeOGE0gL66BvmRLR8rBFVsoTDz
FEU/C9E1ngxBch6HW1S3gkbNUpB5dRcpwgSgBSJqb5hUdjW084E5EU0YRvn3nks3qA5hSVxSbhex
iWtZOV3hpr+Ubs6c/pK0YPieHkDqYXYo4Dgey/l0baJr2npTLQR9uC+rbF/tp5VXh/Sc4/PjRqAx
6AUqx84/9lgtUMzey0q68RTdUAqRMDOOvzeGlIgLFUf33csvU8UcviHWm7Rz8BJDYhLwGpWKJFll
Drb2/NfhpukOy3s1WgJjvhIi+5sFN3/LCQ1q2kvuyPY8DzJ/hgkhUc+1PkB2WVCeZdxHkN27eoKh
36s/8blOEc4d8p0797wMh5HsT3Ncw9zC+6S/LLVOWgI1DLujxXpCQWlDUbn49xVaxo6mTPJDiLVc
JL9yltMFDE7vM6tNYAz4IWcHqWX3HL7vV/1OgznI152BI8lZjNquDpWJK+/WONrJdSnAakpDycNd
s8Y79kseZiLy9Ak2LHqVGdTia8w/k70ZMdMPLYWhQzR8Knwq++W2yERRWdwIemHEznoKs3AdUrJc
NWtkPqtr8G3g6GB6nXSGrQffLmFac6cDRgFrKgSshpDuXT+DRJIrWC2SBd0xYCby1FR1T2JqNs4U
7jjfE9QbRSVs1E4w1OxAtTW3Xn9K14PPTJcKGTPiIpwn0G5hiCkZB8e4jwLdSpVhUVHqnQhirfX0
RaYqqhKaKVPbiqwhwEfaLENOy7+QCH80orsrJfqcl+RjiNyhRNhfcFuleQ8R6OkEpjmUbb64iyBC
VhozjKMQcDESrfMDtiU2CIkhvcebtdW417pSpafZqEKSMon1oLzTJr7vpdAqWfihHccAoHNtTX1E
TBTqTIONqMPd0tu1WqUvUUYUkLSxsWelzM9twhpUTGLyPzFFydYShK2k+oaSI+Ir/m2XTBtK8/7n
84WihwX4zuGzk+dv8p0viwJG1uXJ/cmyjPa1XOtk4pecrowFrGLwOqIsZvKnhfrXn/chvCoo6zX5
gNbKgXVjc51GI3XqIyszIPPSWZ79yqfHXeBZ6t23+HOd8RTyUg2pgChEWfyyAVuip34rUma+Pbic
2phj48PeOgGHX2N8X2siBee8UjkiYdKLX3AIqeMLfsvogDgOMITFvEOIKia1wPN7okHaGztGFU2H
gavkwHIgIE4Y8DSTXmF4UZkRBQqmJA0ANU2FUW+Y8bl5y2SNlHX5G2RlV14864NNrweImZq3ZI9c
TKm2vj+q6gNVsmD7yLirOQ3pPn16SuQ+8X+6KrTebm0qsIdFkfaWbU5kGdrLpYaOmLvGDD2k9aYw
blQbeIEvzO2AdfDs99bOirB7glCMgREo9/YFtI1TiJXSo5gGvcuitYQBgPLANdeMplL2ImOpeaaZ
oBRE5Nnl+PLasov4JhZwfCsyuAxyV5kXJp8neXM+ShxpCERmoAiw+zrJiIMQ058OjTP7zh03XO9f
+RaoMBAg3X4twp6n3unBZZdTvpuyE8NeMb94pFdie1fofjlPWcMMK6Cc3UUqe89MhANbI2smL+iE
hnesjOA3u085KNpZ/SCfHUBEf7/7Uj4Yv3u4HhKxzAWycbgYpoYlb+/rNE6GIOpvxyhZqDDbr0cH
4xPD8AJ3BpkENsNyoqCZLrswAR0DJlC8ZpzUyzf01X+wej1hvyPuxP/QcZMiCxRzIOcR++uYSvZn
FgpU3PP7bHHbqEqUdKzRzDNklQLcCAdqkXOkCqZx23LtpIW/ISkuDMqIRj6NTUUPdY43nxoGVuvG
IbLfuvwB6tG78fGMQZo5ziVyunmI5QQ1SRVRHKj+uE1zSwNsz+NoCbUdAXuCw+RZY45NFoMKCHpM
zDxD26kNyCMg7Jn3H5a2JWmMVLuLxDYEIVkwG/RrRxu88oWwX53v4DrF/w0gLF0xhzMeWh4Xdvj2
7u9etSwuJ5lL8aNxbhNUAg7P5gjK0g3n94xtjar18jZJ5S9Jdsfx3DqQCcyTznLbYLgJMwHjfY4m
cwwITJuRpjp0W28wf1sFbkje6r0E8HQM279FHF3stohSqiBXtbkZP+eR9kL9kyStW4aYwYpjw9JH
/TkzZfymibWnN/OiECkJsjsmWya16ZiWZns7pqeG+GUJl5WSGC1awaG42TMA2u140AYeLKb22THy
qPWWWDfiKk3s6eZIqTPA7okrSx/8rzakflMt18a6dU6se5qjcqR5913sdrIhoWskbuK6xwApyrfE
0PKXFLO5DvuPuNT6fgbMwXWoPPuBolMHBnBwVRDxMuy+TKXByFLo+0o2+hc04MxoFN77jx1ppAwx
U+Djq/qlFkgey0yzJID7ZkG4Y2OR/lK86tG+Qx7NLXmth0/JbzTIx2LtlSUKpMU1yt6laH5HrbmB
MBpu08p9tYRDbN9Qe5JZ/NQig02pmcbRTJJ8w0hMpqugSMgfHJXA5GS9bWb0eEJAoQ4rKnBm03Mx
MiAm03neh26EWdNreFbd/pGsBuUmQmmeAVOuIqB9rn8qTrBxAe/3xp4omT0N2gckj6cqXN135sqS
ouCUyn+ThcGlvK/g4k6iqzoonxMc2bc7CzYvJ6291B3Zm/qfXuSefAswgZnhxx0FxsNWSRvyoWsr
65Or0+ARSowjWp4imSlBzLavi8cJauerqROuFE5priJwwbqsDdg1gQvDINNNvjOFmA4cNKRGnnUD
0GGzmrlQmsmcWXmWdh089Hb/Hl+xt+CfdN/2MnwRymjVMOuaXQpuY5FVU0jF6cEwRnkENg0fEuE6
fPeAauQk4s85k0Zi8RXAfS2JwMo1eOAWEI0+ovaCycUz0FBrHEKpeG3tV3KKFpPxkA347HV71Dko
1ZkqtO2CY4kRzPuVnWf5Zt0WUk3gVKv5WN3Q1zu3wDQDLXyuodQ5kM0Twy07gzerm2LoAkUSjipA
2M0A74+/i69LCjmNR8BYEdHEXEK0Cq2OBbmn9Xmfm8hmp3Zovh3rkEzWLaL8dH+ErauXqyu6TdB8
1pT+HuYG+kyl2oNhykbDnF90K1ynWVYB6myQ/EbNYlqYutv5O2ZJFdbDRydOpuCsjbLrGb3OfB9n
58DdYa16nNt4Y/HttlsRJ/w1tVqVz29LxaScWaUu+hj+qeo6QLw0cbjywc3A7LbssbK+6eJKYXGC
9RhTe0lip/nzy8DEpjdY0W5wcGtC3RQrQG66WNaRQRoMF05Ripuuqo+esdWEUUEAvCGq4nc03iO8
ew4AwEGtphmsYsW+Q4+o50pXxeFSnf7roq6h9VzfAiW4QzI6irGAZ19brNqSXlGmJ9ythl//+8sZ
a3hl+tp0msr2zmcT4NKaZxgomIvXxLThdY0VnMHg8iTyxW8sLe7HDyqpmk651IRx+y0v7S8hw4pd
ttPDqEpzw0PG1PHmBwflrxGwV8qAWYNAAAMvbrUst1e+WF3SwKKPPcKWmPVeiO8cSaF050iqs0ZI
k0Va3jf3fCBuAKd+kgfU+cA9WnwPYkIM/MYRYVdKkSwqf8dhuG32IBkVczdqIOkKlfO6LS9LUUkL
I1+cr6SkfO++KZLBUe3hGSMGQkS3WMNDxjFeV5HAMod9tBX2Af2ut6pSNqmSTSTRmoQ40NTe5ktH
sYCZ9ov9UEsQqkG6wjHuwfMofZOvdZXzDR8rAQq2uHdSIAalPHP549zzSMOve3XODqGg+7wYhj9q
IwYCR1WfCTN/iLyrJlgrOtpdNqz6TSmzA+uWw1b2tkQymMcye4gHKZQ4rUnir6LBfiGhcSkud4h0
kdW43gm5cN7kiuZ40oJ29jwIPSJBoPpvopHCNrXyMJcQM/GVlouxHMrHdJK8u4Qlw0TPQ+/9Ho4Z
Afw49WOhgyKhT8Tq/DIj67AzZewbybRmFoFpcDYh1NaS9jdAOnHedVTsSPPr2NEdMofu9M5y0kQs
x6o7VXjLnPVKhL6T6zHygB2LCN+Bhlx/O+o6TThp61exap2svYY+WQOVTqSiwkTRmTEWomkbgsDX
HmUx0oSGVDjAH7Ni0Rv/F6lEepeztBdn4y29k06qrpFsQ4B7xnP5ioaIpdbnuy4W5UJcizrYODIt
zhn5JL6psRAgJ2jttqRNTFVrRyg0aKJNZW7YlbKdgGBpHDEmXuD7136ewxawlq4Su2gOpYw5dd+o
gRsW3UJO64DLk2mza+cn7JG6fCUkHtnFOT9GD+HYZen7ErJ0FAJEH6HVURXHJxUw48uL1XGipOdL
fZx/Xapdc6eN7iIBf0iaUKsf5TPsoZsMpinnV77LYsokuY9V9eHjpv0Ho2eHFGLJWHh5O/LI4gtC
AbitfHjAPRLhIEz+M6lN7pLyjDnRIUBSQpe6l6H/WBW+K6rzGPINFQve293+0WrjAeen7jLbwyQ9
sxuQZTXH0ikbejqEHXjxils3LAZCsxvMOqhzLcI/W8mgoFdBtrw9vYlyL48ys1Z/TWYbxoFRGOdB
m/YChmwG/9MIu5CUPAa/Z0GciENiRxoMoi61DDKod6eVCbcJ4Rd5tOUANZVoIQUSiGxK3HulPpa3
v6hvglsIla+RiDVXRXzTE/d8OpIUvo/YmJjrNZfoNaWbh6FLVpBsyjAU3p5Rf+ntV154tF8EvGPW
uRVN6HwsRmzmysEc0++O9+ecTWDov9xRKUWY1PLyv22nEFM0csSxa+uAg1/8JpwsEUvWR9N5Ep+y
UoNCEryP2rWL6JbPQUnpk5h3hfVr8Fd7ZPiwvXH5qH1Fn6xyLb0IkkPZL5EtBQBmsrnVQmBgY1pR
YudVXDfoLTpUJkWqKx2NNwkdZUxeLu+Y+EpCt1uIh7vDbX5JFVC4L+YSLXWcdZJnJouA7ikoQrcT
P6amJyPMNvCck7UqL5h73BXhdRLEWl4V2z7UrGSuXyMD6GwdrdXq/KPGjJCIJawQsNWaH7FnPZo9
S8FaM2io0oFRJ3Ap789yj1lX1NbORLQGVmamvDzwRUVGSxz5+HyG1Ei+PRCi+MSw6t/8VBguU8Su
+u+VvON1KYfUN7c1YpUSt1O4F5yCZ9ecDRQojf9pNBMe3tUjubEUHHDtbaLT/F0kN9AMSdD443M2
VZZ+goF1ZC6KGL2NlDZe2JzI+RGRnLd+qvuCSUq8i5QkPTa6V9EJeBidfDMjAJ86piBo+MAS0WkA
Q+9hQcQb72QIp0iyNnxJom1/fDkohsG4CEPlrtMZH0O/RnofSzAELWsJt77jvSl/eMgN5AiW+pKJ
6st/LkQqDhuVXfhzwg4rzTsBhix0V7lelJnAA52ARiDdfG2Jr7VWhuGOoQpn/dzIq0UirSAgj2cD
/uZCxEBaueI0O7CgZQVxliE3MTwBoPB/5Vi7S4G/Tw74zplDviUu57RhO5w0c5cLv4PAPGvaCxUN
7pRerrRPlm4/1W01Md603B3UvNSsXtFQYXJ7XyiYYNvEzXFa1dzY6ClueIKOo5lqxiSlwUOX4sFs
+fFbPGwg8Z0z9pPcSaxzpinMMqMsI+W2npquV9rFcxOg03NKVtkXwY8LyOfvZBN4e6lLiMjrJjjR
9si6+w8EtlDM5F3EVjYYaNnTQD8ywakpytBfK6K4+XI/wMr2yi+Mn88CNJyUtxQACdIO2Y+bRVx7
6ogP+tyxVTYyVUZ6a6KvNirgDO+jpYR/CXMlNZqxgyxVyQoY9E0aw+WN6MJCcJojIFH2BkgqdkYz
ZoM9GRq5s0VQAigMZ3+wEKTqksMDqBy9t/+f82pFKitKYBjDT+cjzXcBunzPOL4w1TTNGiPxcKFC
GzmmjWfKLKr4pYhMY+KKxo9wWLQF15UsBb79pUUw3HvCsLB8GZHlxMzd8HxI1esB08GNuHcg7Psm
UuNAbSImT2NSIcyVlTPZ76a9+e91AT5pmxV8PdE/e/DYc8pDhYuRvfpOf0N8bPF9m2T3cwfzjqmO
3WkSmbeu3SCebNct9K06bNI/68rn9wClt0ZffOsXcO9jOOJRXuT/PPpzXrQmbS8e4BoWptkDruAf
NOfKY+oWedUj3LUUsRbYosdZI3AyYeiYuRam1CK5qt5HvX8i3Di4YLxiWUrqVMKDJBNEJ7muF202
vZNTf0739wQtR6DVP5Lj4Pfr3pe6M3/HFmFYgJqRGzs93QtlcLWy6VXWX6UT/x6JSdVJS0v/jVaK
PhjT+9XNWZNKO4Mn5fjZt8fCGVvvEz10TbyF8vL8cszdoNJ1gfePc3o3qLavpLVbFEY1OScgB6zw
wGwG1Q/HpXNDd96ViHGA05Vy4cwk1MP2Su+CJVPOgMUjcr2y+qjIcIIl1GU5qDbzDYWVz2ocuKaO
kqiQK4ZcQStbaQ9N6kDAzqkGWp9O0ond51NJvX1AD8N9YcemmYKsoRpQRpg2MogJ4GDG/ugYhnZu
pV7NLIIWDyqwOyRD5fznROD+6SHlFy90onVRL0wrX2sHuK/0cgYN8gFl3WVOlLPR2FBI3zqZA9oL
MLd8Fz349xsqKqvGlvp5RDfjkfcKwtIGKd/vO1o7Pfyn/C4OH39rYI1x3pYAgK8HIyM+1DYHkcZ4
Wsu8T2G7sz3aNzKyp2ptbWmWyruSYozDFghE5yPFXvVW6w8tP2P0Ah2Sw9f+8cBetGVd1CrSQQL9
iYBjrBM34/h7un1rrrSRSH6yK3ziNZbDn5h1PJbDnOivHwoiAPGN/vmBhCDtSygeet+FA9RdIJPD
spl5aQ/4ODvfMEYf3ot0buYNnzYrAAPauCP8f4OAXJ1TTw9jLcRJSrRNFR0wSdmSiWVbD3a9bO4N
4mi98LgDo5149suUDB9JjSFG59dKP82YvwaOSK8knOeaRyLtiR9UJz5I8jReKFjySvx/bcimerNL
bZ7A9uBWHErZOglfxTdI7La13Xilsm5L/Ir0eK7plBUTt4eoq3BEzcXqZYsJD9DswTvRTCijKF3o
w5ISHLIteWwa3AwxwhaYygeYgxwZrjrNNnzPdY/N5H9IeJpY1l6llNDO8vIB7ApvtHiC5D0Bj3qC
Ydi1jayAKr0qNYrT56Gq6gk0PmPtDhZn9m+2BEDMXbmQ4BeUBTtQEQC/25Bq3DUcmgP9iAZmKXzN
7CxDNXoUHgIWYQ9sER5jehn9FVL5ON+5d4rs7C/plKYa6lurMET9/xz9U60nHANIlW6OJoP/uaLn
nGsO0xrT+ji6pLoC4FN/r46XQKtXdApqqqTFai7/iwHxy5fYlqdRMbeAnNCMLJPI06fRYosszInh
2DvOwBHL7JTDyCURk7FL9gIoVybmiv9I1DNqvriF+J65/ICa13C2iMM+5p1QbERITgtYnQoSnj6I
8M1tfB3CT1vf7R6YSQGyD2JEEcSLSX2O3iJWmQQYXnaHRMrKB9YpkKNrUgP8eOEomnriV8o0zcNv
fhzd7eig+tHzz146l3t+cr/NOq16/cHEW+g24jLOM4341u+vMS4Sj6CxlARiDHbgRZ0CBBTV/hHI
c8quq84sQ7Lk7NpGYIwJoePuUR3bf+i3IoYiaA/EQtw4YHcCaLOxVsiX003pvTxO2buEwgqAwfqh
amqtQ1EP1K6h6O+1Y2FDx5CwLspCBT4cnNBCmQB8+DYBwjOnTTlwRkjQazRfHYIRjQVZavxyaJkO
aARVU0W5wCGpD87gaP4pRLi6s0kSN4GWoX3N764e3TF5Geu5cUO80FKsssYR9TU+geWGRjEFhm8x
t6uGRWq8msaxBBG9aqrNFKY4FaZGCF5glOEwQjBVeFfUztd0yszZT67h2yJ4j2mkGnRVkiI/9xcS
QFxfgVdlL4x3caaArT01Nv63wr67ObY6j8NcFx1A6BrjPPs9mOYhUV1qa3Vwe15MsazugIYTOI9O
FeuBTaGWOSFXrhg5kEzALDT8lGNWsJQM7g7ntb6EBnsktzbzTuNnhvD4LRznTqn1Yt/UINS7MZew
mGDyL8IHm2y4lj1K/RYUr4febmuNem2Aj8nww+HwPgzM/lJr4rXaZ+cBMPB5phLyUY7tFAolK/we
iiOCpRzxywIeDuP2pjBrDzvn7rcmHbe5hBlQ+oWRs9HL6555WNxQzIgK4NibKK7XSdKweBuwwdz0
F1AP3tejBkVI3YoxSUxUak3M4OLeqPddCtvFrFembhrZ0AsnOAtoyS1AgceNZDkbQpNt2zzLushR
M7FrJZijWcD0NwweiapnDJW9rcSkZPHtvX8cQ3xsNaPGB+D4EJIPxCWS1jzjZ1zm4KMhE2QfQ46O
lY7XdIB4Gl801my52pKw1ciIG8IKSFMQXKrcd+D4b/gNmAnAolT0SyqlWBanPP6Buhyi7lSX33Tp
FMYZUKtBPOS7VWYhOfDo1JzOzGRnbonaEIWQZGUp70tB7BiDX8kQQRNeuJT2sp4aNSQGjMkhSK6q
fxrQ5/4Vz90ULJUXJx91V5J0nyQ3lVGLoFxRsog+bkY7UioPeLR7DWWbr431hXMVbwyLEejGlWqn
OlklajdbLpBK5DTnsQQxPUt5hT/geWvHrcSgcmkCCyIFb3Sq+sqYyfAibseNSgoaBZeFNq5vGjvF
dQDwlruQBac2+9LowLc0nhlTYriXYgJoncoCBuvkVjLAT9hOzdUeq9sZHiOdi8VLjIgahVAb9Eji
PEuYFPAwytWumdFLu/ys+tYmtShbNRXJTXKqVoiyqv4OsYr7D7rVKpNR2PLvIr2fLo2vjVFnOKnk
Y62q4/6cajH7fSdIoOC4Ft1qfdhDxm94yj8CiRjnV/Xy+xEgtt3B5W+8+RdeH78esBBlI7n+BWUH
LEMZCaGXzkuEJ3yNhEdECryqN0Ezlhz2QTLJD7+EBtSD9gunuASqGQfB1NmeEK3y/0SJ+zutoJ6f
xbVdm57YpIsnMb7QHZfKDzPhEzvHsFzcvR82Cw8R5du1oRFdkgiR7B8h21LEiJ3VM26OMm3dw9p5
zXK+6yd5FovW6xsfp3PW4AlHbwqT52OOXwCd6BS3/27H52XHRLj6BFeW2+RhFWT2YjHwrSoIRhFb
+e470YRpdUsQedHNGyN/G9nf2Vqq/9ZAcZZ7PiCVcrv/kFITKJTb/f/1Li+CxUCXXPCV7V+Hp4Z4
b9RyC1phVCrHQssC5s/+khaDT26kcD+9tKrq0IHdjWeSZhTeeJUnmxtJp8dOi7v8C4RDpp6+E2yf
eJCZz64zLxv/e350LY+RuYYdjVbnLrcqGOG37nORGaeLoAFJC4snQbpZNhsQnqEFh4rBkLAm1rWX
OBiwKFWafvL+ijuePvo+UOv94WYMWOKs9F/GP+CbwhB4QsRGS4c2B3Uw/dCRd3pxPS3ZTPsNxCXq
pQmESNxIGth5KY/AMWbtmzFUHXHU4mmQ5jKMExRpIwxIchBdkJ1ctziNjMN694nN5J3YQSdsJrkQ
ul+ZNd5N8kFpkfa7UFvbsqfccGqgrpZXN9/aWp56aYfo2cNy5F4fJiOi3760i3NfgCHZFKV/Y4Q2
C0eSPLCBCykgehEnbo5Y2yFfREO3hTMgcWWd9xZdFdfiXWcCZjk27JJ0chy3K8VXQDRllqce7se+
aI3UwOZ6I/TDYomWekeObj6GDpjhF/EXP9ht2z7+NgZc15UZl7kCB8zFnHN2NrLH4CU9u5EUGCvm
qoy02u92AXMQWkxcDSjyAp0X+GEh0eYpa95AEUBT3Dy/zL7mPmLtXLJbAwnG10m3/Maq/64oLu77
/VfDfD32CsfZ3WmHmWQxF7B8G4Kxs7QJnYHgJJg6e/uPD/TBz5kJv5+o4z8TNnOxWUIyBNeDojkD
Owo1p3xXQ8I1IXH8TC0ymFaIxc/c5oFGq3d5eN+Zsb7eyMLPcXd6VJf6+YAl8IWpMnEvvKcDtHCV
MjRjBZFq7TcZJkN0UyAvXHvytzofZccEXEoOvJAXOzmKmfqoVFhCMBshDr5+pfKWKvCjLdkVTZzN
fYzoUuaLak9c2eu5+eu35Kw6zHstVTyNzAstClLKwpDQI6MCypgIxzzIJ7nBLPLZp19IJ8kRfWQN
NXDJAZsRQcdKveBjGLDxFFucBJ0VRNCUAVlO6djVbI0f1k525iAgSsBtmNylr4hTi5GVrKbx18/L
2q97VXxraDu8SVqYZIrWOHwr9b+Me4acN8+2NQxN1qDDvHRgiIRnwi9EUkQjwxBlA6XIBIPLkwJg
SkBsxazpTsQCML5LGxt9Luv5jtG0tO+hhRvCxmgHHn/TLXTSy9TWzbHq7BcVZz5CgO+EpB5eaD8x
VQ3ydOZWex9b4c84RDseeX8eBWrq0zo+pIDylEOA148aHpzlTlHVpfAllifeDLjfJ6MoRR7GXBPa
oq3TqwKgWxjkAoDO9rGWtWOa2TZvEGYy3dXJ9V2JTMgscSMtGWlG0u89Vo4T325YGMYhaf542Tea
r+GH7y1FJnffP3GpbWe0pecOvtruMvGcq1HtM9MPK0cTurzzqyLVhMnyybu9sYnW1/7bF1DOa5mA
QshlG8pqx+qN/LHApyAn4l+gXrI+0mXRxj+yJOX7cyzA4tpNDQbvwb27AnnNLjIKJA4MZnmtDPC7
cHAy0giPd6qdopdCNp321bx//RxDmc7YFbj37eLDtrpbD8W4HLXH8mZaCPQ3HsyVZ8VIU1K7/IEO
v5gG5GJ3dJcPWX9QvY4yIvu+GuRGrezOs9a2uoTDMPQDVhFLt9J9E9LwjgBSNbmf73GT5z9Bw0+s
E8NJWB5x6B0P3eeKvgHP2Nw7hYR210PtZpXiZuM7xXaiJd6E0nAIpy34NWtqVSszzN+AfbJzhMb9
2JI8DuHjs/DGXo24YyeingMXKU/QiP1BmEsram3Yzynk4p59cuyqlvEi4aGk8i5nckLl5YGWLQEg
knm+F8bUOvh8l7b6xJkHWda4J+T39WGbvBooJNUET65PALn92/EzgfmFhN/X0SUizf7feA670ZdE
A39Ao0DWzUjs04WZJPNlSLeCQNpJvt9f3eCmCWCqA4WBIM4CN8fEJcAxJVIq4i7SuvH68NE2vatc
kR+5U0KqMfQ8aiL+T+CbXuVxdfGm/aoofaplw6vAwoPAVCeg9rZMggkPSU4B91U3NYm8N37lOq4A
KzlM9VShyhTcdYYrxw1z9IEGAiJCL/C8ZbuQEfh9qa1V+ZkS9MCgTkPHZ+b4m+ZIhcQJLpEOIxen
TkguRsIuaPmJje8QjhEJuY2sg17kF46sUcuKf5vhCNwh3QthbhRKMD6IqRJWF2fXXwiRSPPCI1gZ
wcjW72cp1Xu4I9EwK1riRniNhzYmg4eIS07y+aNRvfc7Ggt2PM4pv9EAQUUYu0nLxlQAqV1Ytwao
Xe3wwl8vSX3mnKAijWwPnfo/mF3gS5dWPHiLigqFWgnm9N24xgseSxYv8xhs517/rq3lRze951eb
dt6IAxSo5Kj4Xj5ETkPQAa7gjL25CeMGAZPwHTqW26cw1icH05+hJ+I5n6Zbt5KLLebKw8jh56sc
uWtRCVwwrHYzsdtPgb9BrnSr2bOtxFT3Fig7/lHN7C/nO0IHSbhygjKp/cbniw/uG6gEAnUTHuk2
j0nVQkAC+B5tQnAA0HPHIHyE6Q07LTiI9h3NCOsWTqXxR32vW/qzVJS3MOQMNcmMvpMGksBAhxXS
ZU0D2Z1qR2ZoCPz7aRZc/a7gAxbuhKDICjps/VBMGzgeobbkTkKEv4Ka7WftQ8l6Zfk/OvHL3JEi
Txj6xfZOHks9cq0MY+ewfPvaQ7z2SY0AV0NBi0U17qx6N4XbjzM+2Sr1bMSfFYftwzibJ3tGoGwd
VTpYFtNIhTXRKi1e3cW68ObKXt84+EzuG0S7kp/U94hudAVbaFBO2bjL0ENDTB/tGv5fSIC/JJnZ
KiOUQiMdivxdbOgqYm1vLB98LSqGfbXcmBOTNCRD2xu5IYdsnmWhl8NzmiUZtmasZ8ZPG7sAPWbb
SPMXud33vlGoijI62YckCclDf9xxukLFutnKsUqfQxllaP6O4Rh2xAihis1P8iY1I50+Jte2WvEy
TDGXau48tz0dB8varz69GfV8nWUmzz78d+3KD8Ntj97CTFxHP9tXeL2kWz8ThgdIv+EUjVdNGNEt
jnxqNOceTAvEFG6RyKX6ixrEtBy5OLSTPhr3or9KgSkm+vsCABZOXeBzhlNVZ+ZCuOw/3hUwXXq1
0YvModrgrB1hd0ugafN0eaSqrd0VPaMwKl9HIcX5eE1IRmv5r5obaMGJ2j2iD65JO7ABG0wqJGuS
/0QcL/y3T2klJrEqpo/aoOAQmHU6jzXJRPVYQbs8QcqmS0E5Ov83YstIJi7RMZu1eNFItlewuuxg
5x6HK3gXCWc3x6J3aT4O3FRU+xzgxTSiU7HweiV10pgdAVFPV037vcacv3UL9J968zjAmaTeMssM
fdBdY1O6ppz0wjTxpaISldmoydUcfAdWGPq/cd07aSRYw3BWdxhI7B36i5dluZz8zkfbOloUMExc
u9vyxPH60SXoynSkgBhnnVXAnzW1jHCRULDvCe6ea/1BRi756G3f1nA1lgeEOWckrqKok2whPnrT
3XyjgVQDYa5eydMPfeHJsfnHzczQYIDOXQe1q4noLIHYW96LdVeeg+DVMm2B8mFfLeehjr8xoDAx
eaPRj52K4ptgJRGCujTNa16o3jK9RVTMOYyE0m7/h7O4w9wlZg+M5UJanb1y82V95u1gC58H3WSo
kHfaaXocUnVWLoq+MqZraSNng31f1LFt4HxKYPXbciumCG1/YaJTyc7nTfbn/bGaJKGKqY3URvV4
MJEUeqpJKHvIWyeke//juSluTzuGPmmXLrc51QygXwAglPR0VWoCY2ZGZLK3dlSbIh3mIhUlmgSu
xXyOqnaxp3K1TdfQ4e7QOh/xlJweL4IFv2dr6GXAHOyhAwpzT2Q0wQcpx+7x02disYXQk2QiNTj+
F9apDQ95XMRUdFShfB+5P4/mMIcBcy81qshp2Lv8Jf9azx0YrPMETwayhjL0RHuCxXYoLLKQJqzu
lDJ64goLgnSyvNCqs7/pppPOuUxbUm5wgLoTA2hd1/XTWHDGZ+8pB4GAPy3r4KkJ7MnIStO8VkDz
CG+oDkZd2v2hEZNlDkJciQiwm0AZ+8/6bXw2x2XFP3/rIKfeNDxreZqb/R4VaZLWtt7aYPmbg3Sm
W/IeRxGq002nCfYT2sGjsIUvkzuHJ/S9jHQOs/FYqver9gHfrOlH+RRJduBvV7jBpzM1D/748y7D
+QmJzoPWScve0fXcqFFxLYQFb+yNOAMEnOmKV9xfVwlIPnpf7weEIC+3bdHmoXkn6N81woK3yzdh
H2H13AN74IFRm8yaMxNO1b6InXRBNAfX1funeIfQFsXHf3N4ciantQH4/XEuNh+2yWf9N0qLOSvz
N+f4B8/mM+z+YGGHJyL2XHwz7y35uIC6LuM0p8oB8Beg4zvJXK8B9LUEzgNcQ2BkFDcrZtb1oy/4
HUVp1+y7opaRYRF81eFIJKh3FCgdHzRD01DIEStOeeNcJQVIS3xxab6H7C5zhV6tj2hp3o8mK0zX
BSfEtYj2YHDmr1ceY6fc+OTMZf+o8IX5T2FyegcWzxJ2ID7aaGPCebE4pA02DUWTqc3yRb8mKXIx
jty5a8xV9tmo6EqcGktK6NOHZ8dwjUi6f6ffNKarHZL7Acxmm6a+G/DG7Mj+tJ6dG5GOw74oie2U
rRzDlz3NIZoNcMWFqF4K1B6uUDy0Zn7GpnGkb0pdqOrYY61FGhO67xQbdVAJwtkDkOM1D9+aRBsh
aqctSG0BSWFiArLetRqfVvF2BHWlntNg61UslE1hqUuAoIG/ITrMnWtNcCQ8chkVAeOhbtKFTbMN
1qsGNKKqXq4+zyUTTgdEvuU385BQgdVfu9wo/oaNc8w6Zl11lg8eoGgL5+iQeH+kn578wNJp1Lpx
FnbEIC8+D8SywjW5S2QwQxhckjs0bDveRMMQhlg9Vn2wAtmjfrAHODUUoBDxDC0q7TGoxT1DEowf
MqmoidjbrM8OzNkknsEbT2uUSeRIuDxV8bga3LWtgN5DEQAxVToO1RN57mof8OGDUawsKfZZc19U
cWdEh/Ht7uQ5Xr4wC6d+5eUXvar8fEIiG1Kt/BYz03hJdpf3HUj5Wd8fikLm548IzaZxUnBkaTtS
m3jHahDnjAWfjKU96gy+IZq2eyEZ9WxMsN3OXjWg0PU0q1qRyZ7mX4XF0jUHgvqLfAyam7qSgQG6
ASOOmAN7iEv8NZAiZb6pbvmH3V1I0SgopeZ6wW38Lm2LcM0pVJrCrcUB/3Hjv3GDk5d2flvW8Okz
mtmMwHCqnl6ewnNRuDG7S6Up+3q5qBhYatD0oR7IVZmXMgOiOIkn6O4o40LXMyccYU3XLt6v/NTR
fFCrwoxcfUDW0CtAiawZT28qr068k6AdRpzesRy/wvZRaNzBPQ0B0y/HYj+OU6P0Jc/2Bvv/aTei
8sq+Xf4H4O2pv9jcHVfQkTAv4IXjiZ8Mct5s87BKxIcJpjIxbmd8bHibJXsqtZUBoifthxNI8nfx
nXLNUoLlZi0rE9Dgq62PqVVc3zzLC0Ch2Oyi6ik2w3L/+A3tE6y2yU2Jdk8Rz1vfqefFvtYsm7OB
ZcQuCyHuVZ9sw6h56EItB5mtWEstC50Ay/5uCx0fi6ucLZlIbnjlLnVeJDDHHe/0gGKmyIOKX0Xa
uP8q4fHUaMk3+GNxZ5rIs0obBI7e0yWMpyO8njjE0Nub+Et81FAj/VsSNnCd62fDSlo3AITa/VQ7
14E5nrz0C/d38CifYhkx84+0opeCK+PcO6UhOnTAapZRLXp66auF82HKkOYsNrDM30ZwMxkQE3so
1DyJ0Z6xAirReRm6vpmDkCLG1YkBvFs5dJHvwj/YMVbxveu7WbotmzQZb6l64bSfTeE6D7Qau7TA
Rxr2guDu30a2R11MRQimvx9fXRDvfpsNrHoyR5G/VJp1EqMpOV5rKNBt7R+hqagRdOv91KRISLjB
/EV7VhcLsQ4sRPZkbCB5jpRjOiLY/QT2eQrXIme11BoFcDJz7MNf8YSQtajaHhf+EmMr/mFsmPkZ
aBbWWJjzpWp/X26KYhm3eX7ClD9yLBfEusIDnPPi26ptlJM4PtncgtaFjR+Nl9FSohXFjYfWLf8L
7KMhygABecVQSvR0BINqrT++4bowBL6VcDDIF9DFRYA7pupT0HrtIgiF6YXtHxfsnSDe1bbRgyWJ
TNIWFcpG+CIFanl96h/Uh/c3GbHGIVyR+4BdlgXPLdFhb2P9qD1YBBCwnW0zb614F6H9LdmqtZWO
aCQ6a2zfcQoyoy4XmV+f0AfHbVENPvFxA0R/kc9/IFG4HlgCdZK3doq71BbwlCfSFBrj2zKjMZca
Rj8PZCA8dci/OgXTPbHcbD+HkTV73rKj4zALszczTOzsHOz6NqNhzBttouXJ28g0P8ScO9l7H1mo
0IRtwXCu+wBu2dE/J4zpWNrHPd+q73tpSkYhS6t7rBnZE4Ce+w+7LTWr0Z2haJjeu/JgBnnpt+Mi
jHtTMbCVnaLiVRXibdsTuL+tV2pu/y9OgTtzNukjRyWIY2u71ZtVlv78y7W/fCg/uze1mDcsM087
GHW7NhHXduz3K3z6erg/fkGM9g2dfuMy9+y/zM/RhkWzWJiULforw7QcefrEw3LqQhh7XE4T6jq4
pJkgyZmosTH4gbFk8n1fH3BNnwAMr6HW7mR9Nmzc2BWDG59r6ZHiopihidxAKrEqK19vl1rmwHj0
nR042fByVXl2pwm513RVnWkCxzIfN8GTRvr6hqk+eD1dOV3BvqANuGeq5HGrweRjjp9DyE1M2Ami
8c5n/ThxlPQMoMLiALPirL5uOFOxyw5VT0JUKk3SVeom01GhUzbLo+6b8WKX9iELXmurHhB6SG1R
VLeQGHoWSp8ywQTvnEnRkMBryyp+tUdqdnZnxxa0UDHLcHimN7+m/1dtHf2aKCIVsjZ/ZaDo/HbM
DDK9W5EJv4dyNAtUYQIf3hrGDIzKxbB7+oge2zqK5jGcynHT9VP99VEgO22n5h1rBI4373/sovRw
jDfrjV07sK8GbNE3X4/+KeAmHx2V/ETL/Yswkxs/+QIwjIaVCEbLHSTFil5yA3c7OzhCnZvGZGnz
TADqyCNueEEYMn+4RNBurdUU0ayWxilkeqNeljK8B7djV+/81FZysqLbI0jl83+KyYpf+yLgK0K9
vaFdOIy03H/U8emSpoQgEKdjCZQ9oEz7TiMetS3U4dDP7yVyTxGjwWu5gOlM5jHG9uAxs5r9TkeN
Cc9YjNBNWCNzlodsFUNN0HeoFxss8xWXEQvPvwnpzI6K3ZDhn6WjHcjk/X+CqAv+OTupGoGxq4xm
5hFPR8fyGqkiPIDE1VSYs1KoO1e6C/FqnLLA/wJbiy7/Z6wl+M1gNsYRVwEsKkxjHtj0pFuH4ojF
g1G4Rl1Zu6V0e01bAgpm11E1OuMAzUr63Y5pzvRv1GhAcvS/WJ47Pfr7NH26NroBmsAuqYxitm7P
qOCjRT2zR5XV+KjxDK1AZTaeJqU1Sh7WBZYTPNW7mrFnKloUQl9rlyqeREf718Rpz/nxEeuG5zn9
wBxCstsTP+vs2/lhlNG+6m1macjVx7I768X1rLj6TqGyX3jf3CxmpTc3TOYeFMVD9jRJcnji/hxc
LzbCv8xUXUzskkGN03B7YXOMJfBHafYmEpLtutLjHOn93LGpPWFQnsiY/4p6VBTsl72dF2e/xtGa
Odask7SSUMdtVWv0lHM7iyu/wmjtrclXIuB4vlCzoVep6GYfJLpzz56XUFKJc3WVufG441i4iDPa
IcKC4M9YUNPR4NmeXK9NQOjR3+vkJ+GzXI1rNZ/IYa7C+JUO6FZIiwmo0trYi48fmLuvZLSSnhi2
3KqLH6mki5PnDP20oA16uhY4QBm3y4WOhngauZzrl62spk+6qkGyuAYQ2nsIcj0uxTyYTt1GvTGM
dElldnI+8pxPo5LnbKOGLtljJMJuG0lsT/hQm3h4/1VfP5V8FwGvWLGHKiTuY1GYyY7hVaQHyp6y
/fDnDYfb15MbGRr0dJrCpMwhUHWiMzEJm3vi8upUF7zT5X/ps1DfX6rXi/J5IQ+Wc9Ma60VxdDld
afFnGSAbtTyu7cxedLuEWDOTw59rs3FodQZDxQSx01uZlPi6lucgVaiQsCCCiHti1W3neRI5vi1j
sPr1oL7Z55r08OgM6gFFXZjSAKcbADFuD9IfT9OsX1KHUm3RMjWE2MNlbti1NxJaLNfPlk7lHfsC
+P8lKOj7WpAOpFNPiZa6oU6QUgphMvNjaNB5ayrYK6JLS9n/PDfPLz/o3G+ILuzLpCxOOHDyJSXB
qAgdW3480G/BWluXOfsSvRliDOaB2iBt0ll5kYLWK09dNkKx7lOcdamAY8tmesjX362e+BxvXXVU
Pjfxe74hrgJFXxIVrClSsg2k41B8To/LwJYt29Xw2cjAN0/LMQIpGBLaFhTCxzwcMivBLYNyMHrM
tNqrl9Fw5zt5vDYw+9P+z4bHiq9tP08sZsYT9mUjEn2tzDCSU4g3+UdaWoAnMl3oHPUOHCYApDTl
iQ1L2pnZ5reANxhl8KYCk5edXbrP5QgFTzNCSlReaLmu5y/MGUuhsZsvE/VDfWWWuGmYe6Cpi5U8
NZnegGNzF4dXh/IExnescE09cH4XI/sEc9o9nUYYzQ+WcP5WlnDjR4sbQTeku+9kNZGjchGJ/VYA
WpCLKqxuKeIrtVzTnB8Qfwmve62paKgKcspSoYcVUFmZ/hU5q32mmhYUGbxRTZMy/qqI65vI93st
ViKk9NmcPB3al5LLaGF3KCvIy7i7iV+tKWw2OkSFJbZYLXCEYRLep/8qDhnRaOv5yAfvyZLaBJt8
F8Zltj3BHTAcv5u6hpismCJwgEVWqIFddyA9VKQJLhCX702/ODdHTfD82KMaALLRvUdrMCjXIWXE
sgboX+13Onwmz5xS3531DKh66vdM2AzyejXWBl66EyHjNTRRc+JFbDUGpSRIf+7GfLymzZ40Wacb
mzC/mad6SBFudF1GpZjEmJZG+TwnhK0TpNSh6FWA5tcDi5vtRFJ6ChMQ295C7f69EA46p3h8RRxZ
CIeeQp2P5mBBmLmM9yoE73wphHwSGlxk/S81dfgSTOjawAksMVara6p7JFlv3GD8H29/Rf58lhCR
xiCR94XuOCgAnFcNEOcPf/rQQoW4EIAYd31sZqH/jgnetyeeeSfbRJg7JejLyQTxK0GRVZPZnRK5
QhBvkh01ffUIWFbG3eGinHcN7qgz6l5zpnzsLF03/ljpIKzOwqt1cFasIDwVD+9mU+yp05WTZynD
ZcWBKk3J6ttj5cyCtG5J362uLEphOfJDXDNg/8jBCdE8LMqQdhSCUx3qKVhuO/nzbkPM0levUi0d
vjqa7YrQldZVAZUYK2mgrJkg7Wc/aqCVg82TygE/vuDvlCukzGLlRQFEOlYVcJDaGifexz7RhVb0
+zZ+hincFgYpxGaRQMKjkDl7Ju9zZrjY9hvClDG4FcjC+Ldm/UOgXv3X7V8eiu17hrf+wNSDHrwB
LIc3HvB/g9HiLZQFvoVa4Pa1HllBDHlxfNGWLCoJLGP/kEqsJFL1s6Eo09nZ//X+R5W9BE4zlURL
WxYuVKS41L3qCYJk3scxv8TGZObvuCsC8HpYbQ5i61dpFBYLSMe6LqKlmGX79Rd6JAXjmIFh/YC2
DATNQPu36+dmEPcffcKXClINs1u3OWw4O2nRzzlTp2Xq9QLiGEwhhqOdh5tdKRKS72o1ELuaLeAN
V8Lqb90qdLF380wUCYOwI14B5SHF/MXOrZVxWIK9ney2o5GaABtOb3k3kGSZpKmV5eyyNS6VqFfQ
oSWcn8WlTGXCMq/QXzVq1uEYZ3BW0C1cCy1Tk+fAYxxbbopJrW8jy1tXiW7xS5mHpoIdyoFCzqad
qlUmWH+x0UyfpbbxXEnxNhPBHPDPtyRpRfWq3RYkckpx2n40P/FMZS/+ep1LITL29WOvlIOSz1+U
JKN1YAYJwj4liTZ32uMGgiMif0nB2M00V5FMMqLoA7p58XLGqsJFvAewFHND3ebjsR+uqk2X61dW
M0zXyL5BCNILYl7IRqO3HlJLC8Nx37iAWiQDeLXPg5nQvRk6qULkyRvlt1PAwDUYTI+7+aik67H6
5lOYl5YqV3UHfHJgYnpKqjhj0c/lJrATyY25Oil5fJM1e6bal07pUDk2Nq/tKMGWIjB7KgZb2r3m
WUOz+9BpoqATmjnZnd4Z2KWhhWbEvbIk6dS70ewRf43aOJF3HczzAG7+ryk7IKL4X6TP0dRILbNW
vdrymzxfBSBhcwZdRwXHyt/eYjmbaSvLPE+PGmDkjIaGFErIvbqYhLkGOY81Aq5q55iJhymhmP7W
tXlsjUdDnWJ7wVIC8FgBaxSUt7wHGTczTeUO/cyZragK86IIB0lvK9sie1+yWOaiMZwbuL4hDjqy
Vop++AaWlOvcQURwoSCJin7Uq+LMCs8MXt7GXHfdR408Gl4OUnujvbiSPb+5tLMNVizgXjZgKApG
U/3wC9hr0UKgdki9zLP7VGe3DoIljC9BI+k1Gj90p6AAOnpPoPbPOYDi1016GDuVgV7wSmnT62WT
9H0AWBbO2bpi4HFLuFUe8CekTNx774SjKgTCsqe8meFevnuct1+ukbhsBdj7RPUL6h6S5TDUFwxk
sD+j17KeyfgFrXtQr27IOajKhzBDJI9gPxNe8HQXN8q9KQXNc/9I69aW8kXxmxITqgdKFkwd6f6f
iMcF37OUztHxmP3zzUgprsUxd1owqgOVCKD3Jq1vbUuo8VJzdofFWcpUZ1laR0JpQPAENq3vE8+D
GV30eatinQBNl1DkbIn94N8YKm5N5K5SGu+vTDtRuATfq4toFq6jB09oGXrKRJyWQCuc8rCK7+QA
PSMwCx+jmZY4911ItUAsO5gjCYpRUAPvYnEWwGMEzCugqZVzcdSTSaI/p1h/iaQnWwtOi7QhdMOm
xay7WMAvPLslm/oljWd9q7z/1Zy4zXKmjsZSWJzS8mK8E8NOc9knfheKO511YFjIqX7uLpb+p1Dt
nBV7OdqMqwvUzjS8RvUDr2M5n50fHs/dJWGZBBfTgn+W/qkCwiD+FTQc4JLoMsPuMecD6Ihs35//
p3C4e3onos+MONs+ZGr3gMZAM4Fui04WBy4ikiyUZsYtw1Ow91if4DN7fj3WriOIoAilZU5ZvRL6
4IHfi/v4vy98AXsAjjJEa6p4AQmiH41+zy6GdcEOZEMwFS0uijfXZ4O+x9QRi5/B9O9egUmge4zz
RF9uBdwx2dJN9z14Uav78ixCtlkM6le29Kz/meY7qTa3JLBe9fP766jwkuuxH38CRXmGSoUtaO04
gGziGa5eSerp1fjWRJcNsZQi1qgVa9seF1CjnoNoB9MrKSb6Dd149MZXM9kcsy6j03zcKALWv4Kv
p9pj1/lwMLJG+HXdwBCjEjTBhTfgzLh0S5nAOhep8xw7nqOAtpaz6mepu2lD0+Da8OZAe44GTMPK
5bfDK1fhNCW9CYZIQ4wYr9siLL15nuU1Fqk8WhfDS7rnM/Y3ZMfb991QcwaqcLo2p29JMpY5un74
S2vbhVRB6S3pVLrwrIBpXmvZXpvLHXnWVOuuggeDrmFnaYdfcMx6oh5BFoOm2MTgzjtQxDDY28r3
v4nNYW03nrpeUjmjCXY6hXdhWdmb/BeS+3FGIbOgn7DlEny2JHoDFQ5pi/EbWwsollDRUXt0EIwA
AEc3cWFdTuu/q3yzf0LlKGjSv2DTnB58D6i718wrFpz+pP4P7TU/byoHvkjAqB+XwJB3cQZp3esH
ucK6N1usPR5xo8Nx/vH4Zq2dK8n1qarTjpadpJBYIzIWHw6AGev1luLjNk/irPbg+UiGwmoeUd3J
e3kz11Z3MN4WdHj0wc3+FNfeXAJsQrK6O0dub8xZZD1E7iwNXfGY3KQvCgvP9TcWqgnr+dqJZjXQ
Jk55m7rQiVWiwtrD0oJZY5g1qsFyovMfwwLu/qAkQn2Lo+myN+NzolP+YjmqyrpeW/1iaEpJMbm8
c4YKLx44ve1kqrXfPCP69gIvtWSUq6eP+Xl+ul1PPe7e7VwNY0BQDQ7Qq7UzLklJZ7MTi09woZv0
84SYyIFidoC2IUEBiY95tC1QC4b6nJeHeBwwtWwsRduolcQAO8jsGdeZ9qQrRLq+sVQLkoKToUYM
au+nvZuQpe4exZVWgtl2lqXwgsQ0OVEWZD7SiOmenegaidRh54jLRLsc1W+2F3Oa2Ls39gjnQivA
wtKqeB38FoDtBHELs4zWfTm28p1Dduf9kmaVwyVHa0fKZvuQ2MwlStR8mkdM09EJqowcSBWKKJmF
6NxoLMQOQurrtEZB1a6JWhx2ZZCCDE8qqksnPd0DLLSjDFpYKdjXXQCcZ5wr1v8VeIRbOOHA/CHy
BlDdp5lPf64VEHXMgfjSCz3NzyyyzFt9TRwUmd2mfGzXxsYS04TtDP/lnfZGQoycl/MG0pIaixJZ
VfjUbiOQtEEJ1fdlQafASlBxhjwLt9QieV9NQglnE8MJpJozNDX3vYmVD5p4eWxP6Vv5vnaoaG/D
zuOHs/1kBMVG9e3YK8H8/EkN1n2L2g2iioz6Jy5tiJtjUHsxd5GvS1G+othX1ha3usu4RjVu46bB
uhd11jlmq1Z1ujEE6X7GEK6LyFMbKAPGdO/cw5xuq/3q8EZ8GEBAMoA0wEfXZSzJ8HkQ+vp9SCol
MZi66xDltfhDhPtepPMbm0+ewJyT1JlHIKBm6c/lmlj6b84k+M68BvJEFKHhnEz4pTKD69ds+Dtv
uI22wLeJD6fc3x1tBWw2DMrXwsZpjEgDsnr/qWH3c515zSoykoAlHyROiU7uFDI+e0AV6gZW55zt
hMQfyEKVBoKfDgR+68GhspSfL/RYIkcJqqW5XKVG8LSdsgGH6cvjEwA2JwwnWqzW1yf1ukheLpj/
bJbrxSNhd2Fv3NO1LvIuARvK4Z7iRzDcnBrAtYU4iTkcEAmownWWobCWWqxjCXOdEV+O6NhNHyd9
SC5RdaOh9rBY9SJJTArNXU6cIlUwh2gPy0oyNIsIUbC/bFUoP3srL35BMIud9lei3N2gM2/s9mJg
ymNGWAnQR6Vy8AFvxqgNRS6iA+cseuyQIT80cDWmchtjohbn8S3GhVA/0LGH1Y88VdBjqLDGQRBL
IkUHZGzGuO6uyCSopOm9u8jJpUUhvS533mVTig7Il3M0ZDLmz3Sj2D5cAI1tgnq4FuteIr33Z1iv
CZs0x8vPjCsLlhBNwwWNUdxQx4eWuYRFFFASaZs3Wsdm9Cj0Kt91huEkygZsm5CrVmfN+V5NviUU
qDYXSit7pkqwtHehWnVVjZUA/9BAqI1kPTCufhK1JrDwLrcVrZj4EMCapbI2dde0EmW+3aa06cOe
kszvwrGr1zufIH1k4w123YDijqTByvXrtY3DHSsw5T9wTmlRTpz1QfTuuBZUzDK+REpVhAy9UvDX
Oj8aRFF+uEJK/Vp2o47PT9UfNSKTF188WUMUdIdTB5UJk0EetsFDabc9fyimlMrro0zH966txfTp
SGeg7DYHNPZf3UI8Tu4vzfNU1SeQ7qi0KMXXfUVcfYZ8Bar9Vr5fSxEYZOwULprwoMG/uxmGJHa9
jO9c4lQYVEHGtQy5oauepe3PU3fTRXjWcjXFQ7QXKDAYlk/GIXPouUpmSusMqmfnSvWrBq1XmxAF
/GM+B7mizwvjIXZmyWT7udsySs32TpmzAtE62MUsnHb8XmjSBF6XJTAWm6bBiBc7a7OdUBSHXdH5
gip1PWFJeqT0tLlkd/yVxtgXH2K5vyBzAmdsFouL3XArmZX6QGq9DQLMLfiodumCe34ZetZ38+nf
rk3l1L+TE00PL7bIw2U1EczLzI5FOxY1i08FSrIZdn2zT2lxuUt5WZG5+yUDskcHD2PeqU0h/BJf
feQ3ZV+yqOCkDThdqIurG5OUArt30SuARks2Z8TNvxrWEzIJrmh9ScaFJ0G9pV8h0CMlyh4vphOf
O9LdtqDl1qVQTEbmAqSudoL+mQ02O2hZzHkK8WFY5mbjylVSXdqNA7Yvqee9C/UfZFRVSpK8YDmX
7gtfL5SQAc8FmGsKWDAapzFpMLEeRRrjX1FkSkK3AQ55k0gx/1UklNQERx4q3xBN1NWoZ5ZEo1ND
EbBJMx9Z+/OPbXWzWnsmqKCeHdYarKOQjLiE2dSgMMkQoZtEsUcCWaJHA7VUbOZx2Bx7BgDc2ais
OnTnCxiZJsrvGyJ7w6I3djnt2NOsZ7OSypVRdgJZYhusXUMdOtJhVIbjxZKaoVK2+n8KzXG0mOJk
dgKagQLoPs1fzceltfP/EWqXV11CiNzCTZuXdazaYofvFjewBMdpuQSvRzZ6uHYPvOQfK4v9dsjL
icU+cAlpNXcrDpHZ73SDf0M4HY5Y0tILYaaR1Q0XUw+65GLPE8712nrpC1kU6BRlZjHkU0ZbxXsy
SRd16Z0FF8k5OlL/a5fprwLjzfo76eXc4IIy62JdRdofdISmHtwZSOxJMzJMmqSLo9JSMwFow3x1
HirVeX/Dcu/rEUPtLQ+3b2VRR6xjRcBM/BfXTUeSIs77tsEHx331sCxQdxA1dS6vjx9HhfS0+sAF
qzuLxytbhzQkmL1DfUNJgj4uPD5soSTjK3HPzvAJMfk0Tv8mHEislt2uIdXQVhBXioh01XiQNQok
HMBY5qTZ3K2p8tHYpZpPrG9PwqLhV1Dno4iLzreBC4nj/GjJdf9vN0nlInk332iwvFb+F+x91far
S6l9r3JK43anfdKBTF1ap8K2JYtVT30Hbt1N9XTFLetO+j+xwWT0wuiz6ZEbWdJJuZzi1/xRbZKB
HMu9+M0UBkZ8h7jFjVPXVw8tY9kvr+tsYQYfiNgNGviaW8aeKYalmGtm+cCNd23a6lC5L+uT1Tgo
dH+1ivZdEPg1CRZvk+RnTb2PkSB6LxFkiCr7Vir5bbovF3knCZ/YMe4XVNqoREtjctrjyOeLaLAA
rPMRoaL+NURd+QFZGz371MvmFJWMZtDtFQjw5w/RR0DNSgsTPKCMDIb9T79zwfqrz+ahado0moQw
69gZkwxgD9mFub8n5ufWLUq+gwoWRSUSiAluHK9spZ43fmxn+Kl8U8aw4PHSCSQOtNvm/kWUUpYN
Jfm16agTGAa1Uuuu7kwIjTXsXWenwL4Kjf9uOq86ROnh2JPe3kJHRWzhNCIh4Cd39PEI+PXrVp5q
IfSVTTx8ndWWWp4/MIsBl2kXBqyg20fAxS/FmVGAMC968ZfznsnxHVzz8ZT0+6S1A7F4UehjVog3
+0RoynAFPiCtpbiHDDPcqy6S46cyD8cyoV4ogPVwZAlOuLTry3z8HdheGnM024zzpllG5IYMTEs5
Ly6rlXquTYNNShBj8S/Ra7DbzlG61LNK/uEH0nenHrF85fV0n7/fFm+UmqvPEvk47brfGZv7Nr1/
TSm4Z4pf7bL1GRBhWzBQg7N0nrIKw5WY6eGBN5YBlj+bN48j5cLMTajttbMibbtWQl2ai+edmMmb
pAZDR9EFmRGPRJM9UG09djwfnfAea0KM50txHNPkOG2si37Kr28F86Kw1IvWRsVLJ/41MhpX1ZN8
r/4Q5KYJdPV7E2hnbboAfiYtMqTV/VYBnHtfpQhQgh9ADFsq+6guo5cvnZWkM2tawLzC8kAvUH8+
snrKFlnYAKmwkAgqOBG5m5LBimjNbhifkhb+PzxwbXXi0Yc/WcarIdd3hceBrcKH/7BEEaSf5n8u
ykODVY51+i2sZyJYojlSeok8P/dwgnHY52JhVnp2XZQY+NBOI7GBWAlNU3F4+6SrilhLfbFWE9u1
ydYJKCXVmxETAQU/hGTtTn+rYPejAS15Bq2aeyqy974iIsIH+X1CAJrUjKtAM1djtWtlvLkloJIU
elhtvtqU97Ouj/4d0AQ8wM/nTEqWXnslG83qyfYy2XzM5dte1PEpIoNgiRrIDI/6nB7Q9xMafNam
PqUpCAg1ev6JtquExUgsGZdYjtXGiQAKvHQcsfynLHJpFd/a+sbOuYh8MCZrdhDrzBeE1LekZJRp
PcZS0XyIBgH7WSPrihVkLO7fgi/I2b3BqAzjRI77+pTXDJ0diFZlWmcZ5ZN+RMrYVpfxHeMUQ38F
EBZCtLMLjMiyyUU0vD9G8Qw1CSpAnkj1UhxfFZAd6Pr+lVSACTvRy9SzaoZ4btFwp7WdT6dSYGIt
CmR+FHc/neII1FwRFgVMe0chdsMVnceYDVd1MI9TOrCPKAZT/tn5g/E6FuqFH9QYKegQhYGGblJ1
/uy4GJ765d4sBOzZRSP4xXmYCSeyAo+VAu2gAj1OydPVVIgiSJBvIwJlm+pMUytNxsbzo63Yiju7
0xO5iXEgIAWjc4HIdlUhqB6/yuAO6lHTuWqz/I0WEGd1QfbSSg1tWmgs/DiveejPBh7/K8Er4Yqb
ZS6RzYNCinU3e69HUM5EZJiy1lEeAtzTAYJfCDIIXgSTXH8j13KCPFgGb1WeSDZOLvaepLlvCt6V
DcOKf8T8zYmTdyMjKUA5hDa4ql6HK5R6Fw43bSAGhhO+ieKkgJHLVWIeosEdG6SY670ET196pTfk
kT6tmzkJq9lxKPN6qwh223TgWEm4vxuIbAuolUJlpbk84DyZ+PedowDUdJqto1hGaIC+djxzCH0O
le7ECnY3Vud4Z/GwcDWHWzTEyQLmLR+63kD2lOSniCkSMzzFkA/Lmn+pL6eRmRbKfT1Y/meLGmgV
t7xO6cjazf1lPeweUQfC0mS41sPyqxzbxo0sEcy2b8G4Cc/TVSX2AeSsIRfMSgvlIwXn+dTnFriD
Q2zviiXPZqbBZb/pCfbWNaElq3XBx8NBiEM9UCXnqg7qFciX2DFVX2vJpWQ+RmeS7fGy6lSiB3y9
leNL0rDBoeHmp+0WdxVMdxepn//BA6rJxUO5iff+H7yiUlVh0hpozO8agNql+GB83rjRuZmdpahG
gpTYQuh0FEAPeqJNAK2k8vtVr/Z0wqo+zWsVPKcYy3uxF1vqN1p0uiUKl46nrfx2YWSIfgy2ikSW
+k6no2rvwfIsVBXKCp8/cIzFG1IiUJYDqQJrqqudZsc0UQ93WDvv+AYARJExj2sydlmnWIydlHwz
XpCWqNSJcwSul+737/436Zi7LYMsZWW8V/+1PM5rkFKO9w9a622mrJak2CbiAjnPIExSn4bppxB5
4JQOTOkgKCMjUEfyx2LbjjGgg+n9MxyRFhJ2DNwzAjDpPrP9OYezkAX5fDzah8xNzwOhNmpBl6oP
hfer4t6Xq8UP7pydl8Oby6dguhw8Lpw33mv+qmg6mjjFAFCEobe68KY1OP3yW+PvsO1XMPUeczQR
QjL06ieioMLyRHj5wGwlSt2QNpBP9uqUJDshhlb7v9b2JgT6L7LcHcLxucFo0382rS4podHxUwBW
YuFxJFtN2ewRjwyvzZIGfLmoip7DtxfaHl8Rifbvvu8smqjXfFPhVoiceqjzDfgBdPbx/HbE9f2z
FoXeV67vE+/NEwEkRuLBE/G8xlEDQJxb2QYHKCBpD3LbSQFB/oKgJQ17SXYBX3caDYT59Ivlho9W
GxhSmeoBkXCJKb09Ck8dcls4yzTDHERIvBFZ7q6BZ5GgTf9Pq+izIPHTwOx0tpBSoZgP6qf4JkhO
U7tcKd5ZV56joRsS1bY2Ltu0Fab5pQyFT34/5094XY6eNviFzhdBplCymVz2nBO8NvL9/Rkh7dDa
JEl9mRXudwXDQnLWpfYqti31+F33NlYDug8vKxRIgW1PXvLhFunOtmH4Sq1RFhA5/WNw+y05J+je
3SNh7tVLLxDqAJg4cg4CtVTNvx71prR+jQaNGumm1Cql8XyZ2LvJE9JVxsryaw8ChNbY9lDWprzm
/BIV1GJ3B1fEMz6E89mmvTlKM/VZ2geE0ZDMnQpY3YGCGC2lUEZtd6CoO1X9mxtkTni9PcaQhR3X
lDhRMQcFdtXm1PAeeI2lHPttKcJ4zw8b8Ahk5r7JBXos7OJi6P8zwgZwNkaJ3pkWI81NFYU7tjP4
zkC0BJibMP5kmiXvHogKtbJocud9UggTZwA8p4/SgDzIPqsMCezRNfmEeueH0eKa8MjqQKSCJ1SO
D49VeIi75ORo5ywvYAPewSZM+oZUJHs19TOHwy4TFfB9q+K/6e3m+bWDUUQvSqmWaUWk6hduDj/l
DCAI6lI+qDQUPe9/LUQrenPt48rgYy2Id++AaozFbqvsxFnf0Aw2JIpLbJGxZg0bHMs3IN/v/ECp
v14Sab/vPBonUW2M4cdj9IIWZ70qQjpJfSwfZPc32m2AYY7BsWTJ3h8CU/yCCoQYOIUbrPfyF65U
WMRJ7+W/Zjo/G22bOjGoPCa3nldOYObG6CVdUMaoHIm7dSQrQZLVf1yqkklCQYjQezlfjT0myXeJ
RxMBPNegBkszUubZmppw6JpS1Ko9EDWTgcLYsf+LPRL6/+YtZPkesUhf/oltakY7RqBSasmhua/Y
AotfDEqPaJgcgFAEDPkIiMXEf3h3UgdXqOsVWOVPn8jC7lXPfw0foKN0EXWBEY7CRmgTVJgv99gz
hq6zq5BVKkjCvVJDtk1K2qwvxRTru0X2FPScpRJxgJ+zHgjCRmX/6/5xbC5Ya4wx7QuTSX17cc4x
IkAH7TCEFVMv/7YjlQeoDi5C2JoH0RTtSn4hjp5kQijy4+/gB8svWFxtEL2BqaQmB6/vO4dgEFmc
q6DQwGdc6HUiIhgUo6b5tMCVlSe7JQRERZKUXUKhAKVxmI+70hBX3/5F0n0Eme6fP1i999umEZ2m
UIk/BPrQtTXlo8rQ5PkqEub/4zGj+QSF/Ufk2E/WCY/+PyBNPkijcwRUWYarC7c7l5JpWaj4pcz3
Zfwo56JLYYpuoGWHYxaXMg2NURvJkyYyjVYfW5mSFqFzN6vxK33+DXbHH5WIUArJupUtkWO30AAY
hDVg7fUfmtZml7I6s4M+nRO7DTaUS3EyykqNdOythHLuEkKZIEqy03h+k6pZkFrpfYYyUszwBp5s
5ap8L5XQzakD8xVf7PNPGpMG3NlH/ceuJglOFTGNYci6T6YNbLidZ/dHmbwvFpfqxe63euOjkiCy
tD3rpAjJPqD0rVcrxWqg2fSfl5zlWgSRMeYEoI54ijhnsUAzvPGBD9ZfyObq3nZWmwEHROpk8s43
yLfGvcZzoyrZHW+sh1Ztiy0Y1NuC56l5olMSJ3h2i9OPqdToTdTt9R9PJmy59mgs4yIdH0MFrOrQ
2W1FsW+y/X0TWcIZlxa7JGhaR+EDqqzOoRcF1wBlD+PHt/Oz0nUH5kR/5m7JdgDUApmUBJ177eqG
anZENDVbObJHioRvP8HUzR2pF2LHPGD7X5UAJqN0jDesP38rdYXWVO1qIVFclHX47Xxak4GhMeLH
SoDEb/ruDQf0BA733LeNo57JpEypmX5YC8pqbdAVWXinbcYNFQ9XLCg+H4Dg0y+RkOJsvtCJ/+Hq
T3kbNJuechMv7pzrbe6JUotU6ZLgfwaBWGjKRxP8JXU4CrZUisRaEbR5UTbW6ymYRsJNTVtMzodZ
nYyFMl8S42S5EYvtANxGbdzs7Tm9dUzPoslLZoNfNQOx9rtRw/qKwJY5DrpiAFiUYBQeQm6PO5Yy
F0ruv4lj+ncYWz5k5PnYBs1OqAaHB8p0kuWKD/4LiQxB7WBPXr3Yri5AlImy7JXwF0hBkazBFSen
Wg3swBMzMX4mMtJh9I97rLiTcq1qYMT3BK5+OxgBGh1yX4kdjyO50IFqXBEhMdA7mTiu5kPwzuR3
KHkAZUfjOfqhBNY6A5g5Ew+SmO1Fi2Zsf9DVCeUaM/Cok/KEUq+PYxUCtTeYA/Dge+dc69ASKrny
snj4uuVZ6AvE+GdxSWi5OOPFVyhkBCVWTmWKVrDsUSGvs9HtBCWc6ZjyV+FK8dLuYGwPr0bsFMFm
Hhla65Sos9OM1ka47JYElPM1hWbwwQPahAwVkquSJYzgUZXcVK/RgqgWNsS3iLXWP0PXXWCEHP4R
4FhdEj/MhYEXstX09iMs5DO4Cje3HntNRH7DR66KyFHRjtpqO+XwIXxQQqvZNSx0ZXcJKFkW8B8J
he7Drm/1B/n7y1ku0+7PfQS/BmdDrkx8UE6WlRt8QZWFDBcG+BvLQPpCUsKsjh5uA9V0F88G7b0X
optLOAhJkLm4nWx/oZUGmzG9r/+Q9sKChaCrIBt+jHxJ3K1p5kFWZkuYX1RQv6JLnfsrUxkFCBep
laer11P0znbaaCmqZxrH9yFh+sv9kGddGeNIcfvuIZK17X9Cv2fB/tBPR5gBRfRXeNDralY/jgNC
UN21KoNpQMYJjd4lXkSvXh+oklmi1evfWbY1v+GcuSsumOvOc2dthWhdUx2XzDD1n4x+fTGDj/FE
ARpK/IZxSlIYzQ/uvf2BbgwPeEdXO5OFdDMH8XWm0vYgTmVgi1L5vd6k8B04MOrwzQLh0mN3S4eE
JRLvUYLZ7DKpwY+5B0PvldMMUE6glDlbJfScRZSjz1Qq0TEJ3W2jPrKRwwSzcn3KyZoeHxPN99fw
fcpN0h8Qq4HxcwzUf8OcCK+uYJnDmMOm3x4h89hdbj3xzkufTfb6QjNf8jeHNXI26m43mL0HZhBS
4ajFEjO4L97xHN4J3Q+vhuOvKppt/YdT6iVR18nn8RV6J+Zxr+RTXlhcEtMFb+i4+RGOOnb+iLnY
8TDj6B7tlG9yDlmkDNRvLlJxMVHJRTN02GH3hmQ5EbhszoNeGY5i00pbAJYXQlMMnYsGRj1hSSGF
Zp22b0sKI3KOeAWAVDg1QmrgaYmJ7WtJB3pAm/yO7g+exRIYrjqpuDFV7s+1mjcaCzph7PS/90qB
zgkmGznXxiNsBqyxLllxKgUfYGi+p0lmcey++ZLP3v4V5twk7tQCy1DUnAonqu+icZQP9ya/4Emf
dHvDiqyfKaANyQdvOJB6G30aRLDuAN3Kk0PBDk+J8zsig6nyEUH586BVuU/yIBaANTzzsLqAQGbm
Fisqtqa2LBtNWWNtuqnnffbjg8EwaLHLckPHCLn8R1WlQTdbfJ/XLLll1PxXlt+su0U0Po+LyIr7
Gl7rujDw1LWZtn/AESDB2jsNMdxUxGpCFX9ViV3A0M9DI8S+EZSoeEKfxwm8pl7HPp87sGBDgl5e
bCSJ4ba8icLj/CHBKOVlDSR+fbZxK5tOUfcpp0OwzdlmLOJP9PRgNi2W2uxDgciLtveb/Ty5gPGq
LH0JVIMo08DK5Ra2IhIXbyBSnmXJCfjXk3fmeifDxoRROyrbzBXIdOlXz9sh3C1EDItb6zTNX4hp
arHLXmTsumkLRtUGrqoQ3iFjtFFqFBK+RsZxx4CcqtMKEb8FlKRomDhchtAdqyI3FzQBf+JODQSq
TqT4z+9lur/FNjYEmESFsNis+wjxJ2t6lQTkb4FBNAmx8jN665r8ccRUNmOfULx7EcbyOOy6lk7k
IYcNgbkSc9x86lPIuQ6hxb4FPgzcOTFpOX0t9gUqLL+U/w+9Ab3uBen2yw2/YyrA2tS9cS3y53TR
n062dBz6qsgyyHZLMicHVBJcGwk9RmpMcTTwEWkxLOr1RXc5Brx1Bbl82DN5IxCTAk6MQv/osDpa
6+Z409aDAhvQaCmZSU/SuTRV56lQ6mTHScCmpz1S4pc4tZOdHr2uCBNmfajhIRtBTHvppADBJAUY
SO3oYqipbRcEHIE/gyVgtQv+cNTK94uQswI+5PnPwciUYfaSLMlIuo6trThSoW5lkV4FXVEkaflL
0LltqZb2EPGmhDbCFiqDtNE7OrGruEutDgI6CUmcs26ACdE6yA4N4FM0i/j4kWPiMB3LdBIPA1ut
6c94EXIvJK2G/F8LTQLnbE0whW5bjTZOZLuu/vzKycJW0WB8wWp3lPOv0ru4MCiCKligi71PBV3L
4I3IpOcoqjk5UX1NqFhf1V/qaNV/4lSwrT4eG/mojcU5fSoHy+Lrv1mgxpLR9DPwakmiNsw/o5hb
kNpCKXE1+ysS48ICvilil0rjagyKlS60TCOLwJcQAW9pPhgxp/0Qic6ka48oFWHDiFhgHg3rFI3F
GenTskk0S6DRMedNNJzeBZgA3iVMEtuTDJ/A7NHPXAWbzSKgC4WUy3K2qq/2ZQzdLbx8a3pDz1ps
dKvjIfcw+utXb7eYhxLWxwbhGuV6eUtQXHUEFTlajDt6310pP+5IpaLjrRXRpZn278Jz/AMTZ0hR
6LcIZx9Q/gzfUKEXtwmvW1pFDIsxQYpEtxyt8glNICphKciLDgDJ6B8iK1ujn4CB2FvkNOYeU667
K4iYsl2CD+aMrQCC9oG8q8tpZHNI7GMqzHoOyzlhgtHg+KNRmXFLwiqHxygBXsU6xe46OfX3UNI5
fsFOtQOFlmGjaEs2AGC7EJJTKVZaF+pYubSboKjqLt41kE2Sl5fvEQxuF3x5bZ8l9LXESi+etRxv
0WkMioaUU0M9Wltk6EWrJIHaiaQdGu3e54vm0+cPSsjujJOoIFS9s0bgNqzcOgM6I2YHPQWTV7t7
LBZP7NgImPQ37+n5EBKsV5I84OjD4ezW18542WHoZoCkqQd0se/4NHqgQWFyI6K+OF38w3FcYzRr
i1LAV9tLbZQVgK6MqwcE93MssexUA6bboUB8B5RjL6zksSTodf67vl45XlqWXt6yYPGRWEDD6a7w
741Y3EIlRDxmHFP1VkmOoHr3yJ1TJc8N00bwZkpHxX+Y7j/aofcIxb3niFF2+KtwMb3ZJxUH/7j3
73/RiBwf19woAtiYeVnflTXkTBYc4+A1Hx9PDO4vWcpHlPwkGXjuMaKy+rx5jJQxJtGLFq8sGLC2
OqJFx+zlgCiHoT9yAYP+gEvlJ4M8oI92l2SPU+ISAXf0ewloxx/4SOAfere/hE5GgOF3vEUx3P2E
IzCs01jEB1Op1oiXZnNSA7vsv1N3JPhnQmxdVu7X2dJcLiss1sblGwBqXUIxnYdXmAji0E5f5zSO
RhOxmCKDzubZxykyfqsMAsatMM2LN6240YzrID3+9Y5rf3K1k9n/VySJ/IcoRxqHS2bzReNKGEcm
SnPkZDqG1Xf0tPvS132h0o0Y+ah/LcxrYUUVEMIJ0nSfIxwI1Rtt7ShhuGRtUqJsEinPXmb1j7hQ
MqHSAXX+wc46dafWQn++ck7CcySea8v9nZVyqFhCjb+5JB3qeMAPmbjbVUfbsHfya3hOr99IpIaL
Q4nnNhOkoHaCgjCdW4nX9XBEGeQseGvQbE8INqldGcIheI96LjVxZitDLO/OLzr+y9gJegApNmeR
WXQMVOjgPMbzwq6RVskNxHMJbcKCRJX6tQZmLDk+GI82V2hwP9/EKez9HAcoRwElv/CeH6byR7rJ
DMq2qf7gJx7UCi2idGYMubL9Vo3SmSm9HmgmoFNZfPsLpPi478LYfLp/Tgowzrj5K0O7Iyf4QlKw
T5/lv75HyRXcfQvCQ/jX05NGR38DvJtloZCCdIDTtxmJC6YoPhd9wfZZYdh5Bz0ezBM0qyzc5wc3
Bwphz8B/cRMqsAuzSrGJHfF4Wa+6J7hD89/+IVwG4kgamUsQYUf9cDOJbHCuMGxMqiM1sFeA3iM7
7qlGTrfE3ohfbbnAiqYlCH004BKRWET0cyFY5mhD4EC7n3pMHWZNN3s1xwl6v1wqEK9J6zFOBOry
h7E5juTKbvWMnv++bxArhQ/rI9htkSCGmQG1QBb0O22l+ABrfE9Wk1cRPA9swXroj1cPpPEceq7j
HngOr+8qnQIu9b9Kv4hRZw9c4lx55gc71KLiOGVeCYMxdT+4ooZcNuyVMG/jBoTspzSzrh8PbLEN
wjnEvzpSPwFzHc0QRTJ4XzLI89Mr+bDKBKeHcDojXh+ORdoZ1jv5AuqWtbIMoptaJM88cZe65HeB
6C/1btRy3oDwmGsaZk2thl/HoohZ/7uV5ToK1XfmWrhJUClpM7qNtB4aUdd6ZX/Bbdsm74NuMFOL
Xo/ViUarLKa7Baxnwpk/LcTyBeHta4o2WVEyZhtZSAFZYcAnVd+4MnN9sDXVgs7c7cDnXIfke8py
+yTGv8YNL7ASiKyskYBzsfI5czXrIUv3sKmdX9c8mz+psXUOfEEp/H5oSfa4BTPL6V4aSCoLVRep
Q8L69Bxi0ZRXqCw6GeZmtM0FvxSrGoq/KLyKPAoXx84YoIyK80QCi69JIG0lfyGA+2NkK0IKrU5D
s9XQCxuS3Feh78hf/zFl/4LjcrqndpPCrsqVzSkfCljAFp7/Xxgn+fqZIsVYjOk+8O3nnMzEu6pV
dBFCkedKcx/aILcdiXknQ1II1hAvfmaL6APZFElHijsMVB9JXKmeeAnOf5D9RgEQiB5Uejt4BHyn
g7tq/Gbrwd5hb0/l0843Fs9K0jGotnIUH6sZDA0yjIsOzI2vAi77EF3F+LdpvyEZF6rMXFPxtDU7
LurYdrXg54tycVoTSjQrynUNhfP8GlmZEWyV6O8i2sWHxKIpVJOiuFQcWQKDrVyq5C+JzxkCY9mD
GZw2tTfYkc4I8As3RVlrHi3FEHbBhMiATOoB0G17oc9TEEqCYLr9B11en6Gu5JT4Pfic1MjI/pjV
QG6fD4TsS6SCxFzcUwwP/IWespLmbMVeAhdfu+031iONw0kv5VBY+ff4jvfPKUS36508qzNf4wDe
hFEnUOBK9jNXXaaQCM6GqrFQZgVb4hVSRjCAkKSTkYuHmOL5norsh5WWv6EU95sitA5KRPQIV7IJ
BQBoEPf+14LpqelUo6HcfGwJFYaJxVtq6UUvccVIGIYKaFMpzfAq8JD6V8mZY1nvQSuv2JpkOy5R
JfKB5cZRfOd1Li48itT9D+5rZe8wTcJdWmYZKInqQx+kNfJpQvEX/w+kV2U4hcCjThuvaSUq0RyX
yZqa5JlYkHpy7hNTzDLbd0MfQiMscj1X5oDh/RIaTtzl9EfUS+y3gQmmIOKykJBEGRlzuR6CTfPj
zY3u56DpO0sqDfkD0TK1h1Rmsz77f4Z3DlVZQYXaSJKvRCb0E0/zJmcGOYmd9dQYbvako8F0h++z
ybEmoMDbRCjMpqGj5LOwMmvNpklE/PL4bkGJqR74Xjq+gSlvca33mxTKFcz2tR9LM29OiIWEahkj
PLJ3l2mheNDs9mpw8ee3eOheMTrNMNBlqBl3WJPPejTVL668HWBzp3A0RpwZ+P6gJCZW5ME2jKCT
+TOIr3N6zUwWVF9N8C6UXHHEa47E1MY5f8QqE59P/cq3GFn1pDidSLdP3iRhsxqylLuJPhYCF5Vp
G2PNmEzUkO5HumIMv1vxqSLuLtBAemInKMD89r4wcnPa1qzTefV3l+s/ZoB8KKlWEJenQKQJlrwx
j3qB2+EVSr2xXwDzUsxZNiBVFp/8X12nkWhNzu3vZ2+rGR1fRvdzV8FdN3ZMXTIsILOMtSKQ/iQx
XQJOKP0A7uldrP4sRcepRSQ4JlYL56n76WtKupz//0e/7Os/3JJvLkgVIckuStqUO1PbRD/DO4g4
q4DxpR0hJReCGoFdjHD+ZCJMaKc337F2esIUpyousN6RIdXTpNf7Lf8+51yreFxK2i/2+IibiyQj
Tx1vEOSveK4Q2zoP17yaldHtUwOlNvKyi0OqcACnqWPK6jTSyRMGSgoGV7Lm4MRw+D/5F1UGTq8f
c08fBOAJO7pKdBy6IMijAFc0LrzcJoclD0z6GloS3TFUshUyb2sOobjAmQSIQy2Wllx3br0hnJQ2
mpVBvN01+AX2vrL9EiYQjQ5UGz1R0n/36J/x3eBAZqLR9rtMqspiimQv5utgWABv2YplJlxckkKb
U44U6NUh7zZzgVuoxdwm4KnCc2RE30xYqD7saAIPEcFxJ+zYV0kZbnP0HUARk+4lY8qFyntv0f/a
ENXQwUOc8eeI4B+BJwEima/PkAzFS3eVBn0wwTHRhODEh8dXvLDEEc35ar4I/1NZywvgUgbadJwZ
DrbE1X3kq2U5txxMssEDp/PP5qqMEptk+ByUifpFq5KIZGS553dnQBViTto0v1MEJUdsU6kZdpuP
sPPJNCir9cQxCr+clr3d1J8W/DJre/bFzG/rNx0lSjeagTjKTuuUu3ThGQTh8BmDsyLBgWiikldD
2jLYWYcxAp/dbn/lFpeKva3/bj4FPbYsao6FTpCtScmKigGa1HYBj2wLr8f+GQE0SAgb6nD95ki5
Dlltkl+m92oj3LexEpT6lYDnYr9Oi2HYER+8joec/+pr1rSXoP4tCJaKJDk+SqdnmVh2t0aGKcab
y3JRPpwKxSdVUEyjvTPvONwOrdkFI4Dp2DYgzjjHNxYlvkwg6z+si0x1/jfLRTa51+F8Ug6PYmoX
lpgwh7lFdSPQZ5BacE/2AefV8cl+qVRZfMUcNtjf14w/Q61S3trZLAGVpym0rIspBf4ZDwSqFO+I
0QRRVDXfabMD9zgiA84qtkk1X2nmKUSodeShwJeIQ1jpmbOMEi5Nw/ZYgm0FYfJf58f0HjpGoLvY
y7XnSlLqdz+pvI6V189x9OgRTK0LBac6tO7pvlG49ZSMHLnAkBog1j9MLC+NG4+gv8tnJTh/Ggu0
oLbq2YqFjBs4qe9hyGnDDjy9Hu3hIkA/WWlJyV1osOEcTVtvzPh6WZijfxHsPHh9MDdluSWSDq6/
DhLbYJ0jinHyJrT+FVFc6nYpp7pzp6JYidvVuhwPQjDiyE2Wk/v0u3411LM4GwGPbPzehodXtib2
3tuaAp4JTPOOc/y8vmNSr9F6jZas2y45IeptVwj5vgljH8pLdb4OKDCSoCEKYqPnjZ1Vtr4qb0aC
6mA5sek7zVa7+YmJROwm+WhS405hCVYVQn4r8PDkgLrEKjI/Dt8TVyGQpsiWZeJIlZOIqcOxU8pP
1RhngyCnfVnaSPM3B+WjACZyb6guzBoVjfK+J1KV7Mo6FVz7p1226vn76vVZfL54cF31DGoztvIK
FrpqPg+4vdUnvCvX9f5vMGk7v+AaPzisUpmmQPkovOBr8Fc3u8NIpBfwAb2PbcEkgCRcFNVindwb
JD4WhYuVQrRLAYU9AHhqswn6LgINx/jt1OLELB3XWOun2GKDqn7QoVZkqua/RmzIfkO9cK+1gEHV
l9HZLTRxQk0OwzFEzlOPlGZVQTIA2HPwjrDRJG5wkuGsYyh5Ody0t4uTliXkObhcNDtaoP9PYZjq
gMNHgl47R8o27ylXZTMVmOK1wwGoNWUbQT0lwfg7TqyxpEWjRZ4HySblgMZnnwkuH2gYmWjqOuVH
NUZKfEHgBAaUssjNEX1E3nQCXqrk408nE/zrM83Zelcvr3wXTewQmOLTA/rlzE76OyXpPdkmLHZR
kLWVQKe59ONEQNC4rIN3daar96XfIDAd79QcAqQva4LkkCeSGnthRx0d8n4rJJla21k8fMKWqXNo
+WgSfKYxi3ztP759PvMMQFIyimO1o7AgudvyqTaZM6SlxD3ejJVZ8BLscJLdhUU5YdAXYNx7TXv4
Si7E6OA8WlcRnzonwSj8ofKNsILPnGJEMF3HE3j7o/iz5w0ZdhbGaHZE8WF4dFxXggaKoRAmkQdm
IAbGGkVt5IXLMrZ5+/rwr8SrY60YbsOGpcq/hPQcy2RI7eJ1HHDmdN4mSOWCCNQPEhS3R8n0ia7J
9WWDabWwQDvb/16EfvRcAsvKIw9QHtUQnUNBIZ4YhZVlJIabZUbqD6dsJfkMTQkDifcXdCTVj8HW
iIiveEa1lKcHJP7asf9NiV6ob7pNlUuQUJ0BulUp/7RyKXMhrWY/aN/HTJylEqEPm1LDKeklR3NH
7pwsEu3NXrA48O5vVcScYzXklKNd32wwvCVhHOuAFXsPtFHEd1JL7WHV5Ye5k2Aitecx9f41NZj1
d7/XQOTeI1AvoDDZhJM270sef8utFsrsx57856F92DeUd+GBYEc1wUTX1CyzrYmvnj3uebST7sr1
mlDsrxyHkNyg4+UcHm2zBXKNyxSzWExcgGJXNX0J0fzdsAcTyZPYu0BdEhXWn7zuL7X5W6x+tcYy
jTOeZJNx5iLr8e46BqbI3yVWQiMGUGKuqr5Hxgsx1/E7UJxVGomLomm9QmE9e43gXqUrsGqAd57R
egCjmBEdi8rqk2R5ktwWF8xMLjUeBDVkDgorZTmLELuCAtbqvJdXzjsyld5MIQl8NdNkBD/6gUJ3
hAXid0vVdnX5Q+qLyzWRJOa3tJYwPoKwgE/ldqr8T2DA3/2URqnF1lTGBdd0Jj8n9HilhilXc1Rj
mMvV9N+wuLVOYRK+rYkta4BNBh8LkZNQTl6aMSHn3XhI4kgKkpoU4u3bKKUDmBcuRafI942fK49O
SPf+xXh4l2XiyAKERGlg5A/2riX9O2jqIMY+ycoUAaegwWWhh0dEEGw1oBXHErVV11LlM8im6RF4
c5YHN6Ka5g++HcnPpgYYXv3pwKxpk7+AM5ZOm4r8Yfa4jIZopwQ6f9G7ZFNPe+wv8afQ49Ax0IkC
YV0IdN5YA0MSTI6zdq8/cwJXDb3XkkxVk8FOaTrMQqnLnPQGKw2FL9PZjZkd85c997JAx6rxMx/s
Fp1WdMXHW5N35m7Cm+TFqYkcuf7mMZmSKNQyHV86yjCwlLGsDTVM37c4Y3IwlbNmIROmh2D3yuBo
st9XsfKEtIpHLS/BvAbcaUgWnkAwwmYOcEBvDgkBBLhivygNlPmLV4rlyRkiNZr1s18DGi/i9ESr
YF8TdKANbet41Rdh4lmaUItSZSZNKvfMEzM3uduFsGHsS6j+w980BFz5S/bdaYENhjkfpDmXq/1B
rv+Tlx1fTlVD0SJCUY6K1F1XGaqxY5gZNY9FXkmZZ5RCQbZCW7V/ftLzDF7kXSuZ/hO2j6EkJlIg
FUrTViII1KniJiWVhZDLKjlTw/kGbVdAkhTyG443LZQPSqvOPar4hkAvgK/xPsFiB//TjZgYy/Gd
xipIUmTsBijF1jDF4WH7lnTXuE/p0V9YTf3J5hgGPuvBxMTCqXtQmBcKUYErUnbHBEQvJI2EkQxA
gD4lgA17OfaMUQRgwBnDawlydOHozARbWDv23DcdrOyYth0NyI6A5K0FX8eSK0MG74vMZ6IrU87P
I8dUCD0Y1XOVZTP4v3pCnfmbpE3Z89P/PfDLLCdUqbF226GhLeKrR+pyk08VaWiawyFRAwIfqyma
DIR6bRdSuh7FyH7aF2CVJxyt5oYSQqngQUn1RWM9pcenBxVC7xKROhiRtKwRYqJPT7h+fR5U2Qor
I8AqWs7jMmKB10dyqtuC44vek/N7VcElyGA0AdudgDFu322sPGtiIx7LIzR7NhAWsZbV19BZ2Cx7
QENTazaqZoxxbkjiQ03LkIlor2iQhUHGXgvGXRf+1n/ltbEb/zTGVXFe2RKdcH3LyVP7JNiSDVek
Abihapnm734VADVtxLIDEemfFHEX3PDP37LmPvgb1fxVAgBnLfPcH2sij196r3HyzsosHQGhsWz/
JtT9HkG8J0UadtFZUfERRkmFmBMv+TRWimDzkChaVyij6NSphlLLBa+oUdrYpGGPPr7TRzDKSTgS
59fcyjkG/e3N8WeyzJGkkfJ8A3jw1H4cq+RJViM1dBdVpxsGUrCT8dRoNzg14hb58ngaQ77Z+f8f
axMrTpf/GE6VkjrsXpsaHxPJaC28Sh27wxMtb0gcN7KF1FnfacyPzxWHCVCCOb2+tyV8dRUtB/wX
X4D1d5W1VrA8F+36mTKcR7WVQNBWoms4YzZRyvJVedeaFDr2il8qnWWWlpdvUzlXHMpfiYuWarAt
J/t5CVZDrT9+uCuSxq1e4gDCQyLFM6UBve8eriBdYalQ8ZZb2xN1vaa7Yk36PiUddySCOtnuVJ1w
VHK/CURE/PjwEF+0GecjTgMJUA8QWUFV/2TMMpXtKSzlV+jd5zSDif1Z4wi6fwmUXWYuR+JCuJZV
POt80LeLfHlfy6wOwPL/0Jn67sDUe+8xsqba0glgxCu6vVUBzzp4D+b5wun6SyLlJ3WtN/8zUpzG
ZQcCJSogUm2DK5MOOGmfzMqvg7Q9NhaRh2d2TclANXNPu6Dsm4a968cokEJfrXOD10NAvUSmDfnh
TEWWU8HZE6ZHA7XexUAeo57ePtI5WOfhk445GfJWY+qE0FKF3L1QzlOifbp5XSFAbeQXWx/XwVEq
n3SnVzDkhh8lswexds++cUknytxCoy9U8iUjwqQ8kizaY0xoK/crS8WHZUafalQCj3fhqGPtbmPY
cTcyO4xz0z/oPJo6m1fhtW3X+CMabD6/BFUNOnrKjCNmhFf/fUdiLvtY0snKmz8vCBYW+ylHSUsl
iVaabW1DGLjhHAc4beo9HsQFMEijR5868halJCbeyEHRrYuwhA7BKEBhuRAKv/1vLeLt6DBR9847
5Z7YznUrWj4BASrE2bilV5vZqY9xa1ciBsrA+QV0D6D8mphtdKDfHWNYUS8ZfZmGadnsLLoqTDdw
lLHll+ldKdh42BAQeP02lQMud9buTNTeSm5SECk7tXwswaM4NxdLxX47YZBZn/EN1X4zSQO+q0aQ
oq0kyU03CfFgBxrAGBM5Gye9Hm5DTaGgVAHrAcLGhSeV14xbPGUYjaufTB2GvXFDh3CZqpE2NgFv
e0dt7uCXPl33MZGM5LIfXX3qseG2riLhDAe6VmSVYJRY6+gMRFuRpqBbsiouHPQobCsTONungET6
PkzCVmToejZbP1ato4VSfgl58zrA65op8w2DYAurKfSj376NUWXWmJWlfMjIq85Yl3EZDB2PjAWA
anew1AfG7OFlWud9NomPU81fd2Iw8A8Mk8MbcLr5Wt7DPYsjvM6vamos5t1OJlBMwneG9qUGLvfG
C82wcxwJy9HZPo1mlyyqBAAwMgCyK6Wui4ktTYISsJ//hXzXkMcXbbOtmF0x7sw7q1RWmvCbzb3s
m3ZkIpzxwH/z6wJIUIpPHy15IzAhpJIQu6DijWvB+3J1G3M8cmrOJhaCiNst8f1bXBJ7BFVqBcMM
I8SdDw7Nx22Nb2ya1NRzee60Wt4+DYhSXMTbHjJKmyD3rTTzyt/Z+Sih4+JVn7RXvtsEunWlZq9M
lV5OZAqvr7thXnioUAz0iQxFN9+4Yezb5G1GWIVg+6VP9603dTUMM+0ratnTq5Bsbb0+2WXsFsxa
grFW9+sgeqn/sE6gTMtqdPjSjr8FkXxcpIyzBDdVAkD4y9Inoaa4uuwbrOEue2Gyw87tRwvSxwjx
NLkvArksX+6ah9hm+lIHm6aDvyscAHPldDkjLgBRuAT+GN6NPiYCTWoaEZHKH6tHLQ5ieYC+g5Pc
82p9YQNur1Ls4Ttrh5kzeiORCrRn8IHXUebo0/KiwAMM6A/16naazYaNKG/h46rAbVy4JELoUrMu
0h7Ewzez5d6D3V/wwSxMSaLZyuKuY+tL5TfeD2eWiKVVKGOUro2Gyp4paxXqglXR8KnEmoJ8MWin
Boi92u97Zjprrt1l9ZeI/HVdrXF8Dq9BwkfrwFDS9ng25q+VvkNe73u0PNGkFYTbi4JdOVDd6TdU
mLNRV7LDV2flTMIv2xPGJexDMvziy1PxsnJaCxeY+hkY8HeFJwiyLwsWpGQV6Q5qcVuq+WjxnrZM
XyHGYwalSHP/crBP266vsQN5u8xJ0T7yOFRUDb4SLcAqCSpU4zEdpAibQYh1TuJMLfJNzunIqRRi
G/WEX+lmgDJj6CzEw2DFnVLEelLt9yEPfS/aCTyGHpKUjYvOJUTXvNaXv4ejiSi36m2W2PxJAMWr
wpJi5dMe2FlX0x4yRxQyedLsZ6LRyTU5n2kDCahIgLEKFIxPKSKcC2Gkf2LJBIdjFDg2wDx0sEuO
rvhHNu5s6WbcEAq4RC2ocGrTZdWfsGsusdvs0KvzDvFsTqL6WvU9E0GgE5Ed9iII0unIMBbmq/vk
YCyDg34g+PZbOpRrmWL27+hAhpQ04Mm7H1vImbpzXI997sY55bjqCqK4MtXWb5w2inXLYdx5ostY
VWcj3ULlAD73UzBXB07A/6GhSrdI6d0D7zbnTL/Dp5aNZUelHgdQCLP5R8hbdcdr8C11pEbTbJLs
3DcoFFCA+Q2MOkADhjTduHJjjTwvSxs6l9r0ZF4t3Syasx4BIlpV+JQ3WvdA1FBlFUzIhIHZFn22
H+Jk4MRqSmGOdZseMxekdjRwqfMmhwhhtogVD/szlWzT7jb6TH0nq9+GZSfO9y2+3eI0tU8kWJZd
gWb7lqIFIyV8RgTxCl45LJiu7nVXSCWFnXZsoFqwTJvvktPID9EwE6Tai/dT827sd1Z3thOqkJZ5
xmxJibXV5IXULrn/fRwJkwUI3sPRgUFN+LUgltOKFv3C6h/YQ98uW57h+xmgROjqaxBmNoHBtLmy
MxG/+Uxa740m08j6qSioVsLa5sbWtnZPVUv0f6AuqYXzyD+VqavkA+VJ3ndwXelejMWsCQUuaYQH
nfJedy+K4qUrfNRzmTd3vHTTg9JxAxHxcQJl/B02k8xLxNSOeu0S/JWvRgI0orlX/xy4pvne71RH
cOCqMccvfZ6ASnjLX1xiplrFRH1Gk1ka3SYtOy3quSTnHe/QQTMVRKv0QLfzqeN0TQyY+6lCJ5r1
iwB0aMOooDi0F40wnsZSkv8TZvn1ktKlzKQRTiNmNvD6q/gVCyFJH7khdpcPLtWw2xn/LsvqEi8L
YxHQx3Nm3OYNGNrgAAoGs5mBtlHlOzB1RoM+9hlbb4HRKl4uy8fqE4mG8heFsEnGlxkjqkOrVm53
n0hhBwg75MjTbSYN4CRTocJyDX3tgoLeuHCUwxjdk1IPo3rK9u0xjO1zftFDaRvqXdl9KBv4LHGf
i2sui+cof3zX1efN+qQiily5nqfxL/m3XrztXKN91nqTDRkYN/TV1ZLGfsTNtdiitTQs4y6QN0Cf
v7hx2adVVKh2a8vfqMTl1kT+M7jO7vLc/h/Z4rDtSeqlztZmi+m5OQIgegONLBCYQCzvQKSOOhdL
S53+6H6cN7BlT9VUstWwD0atWp4+ZAqXD7SymR2IWEYYa2y1yovNQFn1/nyEX/y9gNEc1YjlJjlz
S73WbSTuFtpRJ7CzJXlDNL2qQ2OpR2lrE3YUOPrKl8qIeUmE9Un7skIwi7Zvq7pp/sfS5qtYclLh
r8Po6s+6hHcFBdzABDOXUe8uerl4zITqO0Zv7wG9H2OTvOEZKX57uV72zVB63Fofap9fBltJ9Umw
cokU2Pp/sb/EunahChChP1QrTCWAzejPk/L/uvZ2n98AOI7OweQGwb9HmmLdqp2eEWc6RdrlYy0p
UTqg1sGA2aMLrfiznUopOy8t+AlSYCwbbVWDm1injo8gkd5enW4LhU1u1eImoeWj+sj57AQHmGFL
5KsNxnGU/NdcQEuO7LKoAs3U5OEd1IfBhMsGQqNm2RROOFQJJeCNlxmcucwfIOKgEDO2GN5V0j7S
sDob8vQAPS4BWFNz6zH2x+3QiwZmrWyUlsJT98oK6jxCrKKA29fQx8u2mp6WeC0EGTFWgGDgaDGj
uCAXpx9GUrrMe04M1ouH/XFl72EJgSJJdBnNZa3gBxiogiLKffXFKjCxfxpexcJUmfsRNmm8cJau
a+0JHIPuAkCTKNqHUA9tA4DF6LQ3dvwjkh5YgLKUIGWPON5bjYydTaDYuu16nexS1v/UcS76z+kJ
VS/xyjYSMzxQ013SfafEpnq42IzSGYqW29Agpn/R6RPQ2/8nBKnd2VjJJG2JR5G4zpF7ScndW3dG
Ka6rZL1qw0O9PCeD7NI+CFFxOkox5YSnL513PVAG/NaSyk9orErochs6jlBJ4kVbtTIV1Ofam6sQ
AGFpJyhbOTFR92uByEkyIeIgXrDP9NtPUl2tb9WuJA10y3BqO8eGH+/7zwdJAlWT8Y6oi070Cufg
oFWE1cDwr0d+vw7O2IBJfnXZAS4ZcQ7qAWv3SJeeTm6hYWZaDOJP3G2Qfdm9W3VfHxsC0AezSM/y
I9zxyHcJ/ht1kn7fE0D4BY3uX7tHTsDQpsTzUUgGuej8lc0PLuUVr91A0eGTA4uRHPm9skzL7vZ3
4+qPtFa39u5KVt2vg1jwbH8en0fSdZEz1n68k1tscHSVRSAy0emKoG7QhNH3lGTnmIfgSPKgJS5L
3F259G9hgazFGoE0ECWj2Ru8t0FwOzqr3MmoO5cTwfWyqJCKFTu6shu74YDHXPhuZ1V7YWzJyfs+
sQtWL+gRcdqNixLi/YjWZt/TSWvsJpwCAyw4FNEpvlhKlj/wxKPcJ6bcolN6+VSm0auhgvCy8ugi
G9AUe3UfvBPNYAIlKfQ3beYXW3ECv0BOAjxYzUK89T2sNKEbisMbgmlJ+vdw8c1FfCNjoSYROcHz
Nm3C38XM2EJVlNbN9FpYZt10FBbZzp5cB2fldmnAjhdNAjQKh+hw+BDv9znvOMdONRlvCg0VnOF4
IpuOWfuyeoKwF1d1QtescJVA3ETWo39N4vFKToOu4gw9p2NIy0r5OwBxAcZb2FE3LWFyItGwCVfG
KgE3lADD/KjAUkQVI38KYmOoqvf3Ufz26yU4B0PZWLimt5k/UGFZo8Eg1o9HCWmo5WA6g27tVlzi
CzK3U/GkFzCabSOXVnQ2l93FnKJ9cfIQ2HNRK18W6S9+GV7B4qwyval/2BRhAKakvRJMTwmrvjw6
i4eaUrTyDG7WR/Q7QILSQCh/poZVSL7a+Dr6JW6fcKRf51tAX1v8HAlz2m0oxuTCfmCt7Bwb6BJB
g5T6lGqSU3ROlHIa1d7Bx1jZ50u12Cj1o5w4PJ7DdYjj58xKwL0KP00V6tu7cvRjp3gudY+5mz2b
wgtgkCBNu7iInM/RP5mfQ/qvB5P9v/cfwcLSJmwxSjpDdyJobssskIAL8BoAx67oB2jnE+WE+ukW
Y++cZUY25L1pjP5UdBtvqjwZt3VS8JMSTwOjXF+5bf0Tdi/HEQeqlGX1ystMH+dyDvVWK2BpM0+n
2VIQTi4/xf/Uozten3WR5exvRJ8FDv6kM7CSakuhHhV7BcmakbqSCjIQolXZnI2dKwhFl5iyQDFn
mLLbOXkI60yi5KoVbMKxGm0GN+5cBbQAN5nrRZHrbBepvhFOnIp5uu3sMNWQa6C+KF8wdpkocVnx
TP+UelaDNQGHBwsQFjKNNu+IWUnm5wz+mA7hf/AbxabGkvQIA6YC0WseNBc4lEdO0DQK2dr/z/Cr
RZ/XNbtndl63/Qg5IhM65BL9bGn2iqY4X82RLIcPrbXqlXAzIB8dQy1VBLFYioZ/bPyxEwFKIr9Q
KaA6A0m8C8n2YpWHT+bvpbnXmrRiKgc3D6oRGaoDXFttWat/vtLvzKvgDf5AnYttDLwJpv7n1gX6
NMA6rQ+g3WZD2u521mc8x6QaD2IT6I37cIMMmlLybo9WjKaTpvNhsVB55VzulH2/GtWzUxUy9e/r
LBTxUurDjqNit8VmkwLe7neZ9WqzcgWlt7DHnvRIpWawjNrGqPUzywUWmLbU8EmW5huAsv8tC1k6
bsXK4SNWjGo2Gl0/J2jy/dDWugfeYUALLcFUKPPCCv011bMEI9/9cgrfPxA0qJWXe7xEAd9f3zpU
x+1Js+7rFTaY6rm0dcdl1plfmEOEiqaV5Z8wQvQyfJs7focoxtF2Yidb7ieZWftTJNWRQuuoGz6s
dKgFReH5nb+Cg7t7CVUjgeQmhJ0T+HkxWhayNoe8VDxbyF7NtdoSy5xPiAy9LnZ3UDuyhwGQd4IH
aZnB54/QSExENRlx3AxPnIQe2ozWjKgeB0TbYWf2cwVIGVQqKrlB55ON2M1QWjsLCYVKyAtkfLer
pj3aEduectIqV2k27UqVL32fhexj9Cr/doSuJIp3cVRw7ggKwqhxE4zXMm173CEJzxMF+ih/wmn4
iqzWH+e19EApJN0EaR/YReN8OrevkjPhyvr9HkHvLpanrj2iPLnFfvV7ZHZfdbhQk5qdkQY4x7Lh
mU5V0MCvs5sbucwlNCYwY3It/oSlIArxqo6s7FNxGGnDoq3cmx/1YKoTppdvDvgmqkSitkir3iXK
5tHzp/bLXr3p5mHGvZb7GxeHgn77O7mj6s9bVSlm4JVuE3Zx1WdEfB9oBvYLtrxS/eDiZ+qQnQsb
NsTWjEigTEi/Pk86XJztm9kMDXugm1/8eFdEeAUFjD9sQ7FlYFLjNPnjxJEKL7cnCJHuJde23cN2
uD64w/8aVbOkvdiJ3tF+cxBSOL79wv5/+1yv1fsScciUINxH2PVIzG1IxIzCmhQKsPWegKO2UnnN
LZFNFScLVuSOdoFUgxLuKLGnaPG58cm8nNkAE9OTst6qT/F1isqxkIBy6m+C56NEUfzAXu1trgmG
+pghbrpkH6fmYIKAuotiyjWLXBX6L6DKZ4hhBWWa9SIzyWKC7ZKZo2oiKDpQ0hIfcnn5p21xDyuh
2gFfEK7j6kl4zbEox3N71k9Se8W+YxyiKbYyGlV/Rwsntweb+3MKaoE1PsV/LFyJPjOXQ6itmwxC
RDg9T2080SX0iJ1Jksopb6cZNoYViON6JnAI47epU4f9g5f8tU+7nnQHPyVleJxaamQd3LS/0vFN
3gpXOGs94cC0bn+UFViMHyeJw2oPuhvKqlRIaiM6mvYKacpeWG8givF2BqqJ6YK+reDBrUcbcaG7
C3lgO2jWFicbHDOUDP1IKTqhKzglaMD5xd/q9CWocpm2K3gEEKt6vL9R8EftTUVys+EelFPDoQjQ
2ECvF3nGnl6Szgn8nuefsaKXNyBQqnMeAlAswjq6N28K2oWA8ktHd0YkIFDVHQ7V3odWoiuhMR+b
GnHiD4endoCgrwMSAJRsokyJ0HFVQc0fyw1nWvVNZzehh+aj9SoHOYAeBuYiqPU4TIsOVIN63uBl
xC1pF12smwWhpYWxFgQFERS/VjVNqcpK8H1oZxNIoKLMFCFZ+sduIjTnAKW740x1fIHmzpUirnzp
ZnRmG7hbne9T6KxQncB5GLs0xOLdnaVhV/9rIljXAq6D5aE8ZCbX+lfKNa9wl5Gw/WjzIcHgB+hG
wCML+0puG6rAqgPLWleVOfo+f0PJ4xfaRk7v9ljJ+dxeUt3CsJ0ty/DNKbH6yJBxktb2qUD/1AZN
3x7pJqpElz5NC69KU7Py4ybJuduAUeAMGgC7DLOF/TSQM93Dw0SRD17uYYH9a5ofAGdshoJTGMU5
vMcGXvwDRI7/br598211ouyk7F/i6aQqv4DcRpeTjXvLPehOFqY5HGBkN17MGK5wVBGJ1pA42GLK
uX5+bygJnq9wm0FVLdHX1rzF9uKihCN8UeO1F2L6GGqItWdw06iDWg3f7k3V6rSmkVDq9Bu8n8wc
qpCCwmtKfDRCbdpy+WJZKgzFcm5yloylB1LXH/uGMWG0SKZT+Iefiz0Pcvv+NkFaonPyZ42UZRmG
Fs2rsZL4bj0UipMsQaMv1RQasGQ9f27m1DkP53MActtLsW1SsztuZXLSOrfO/WQAXkFVxwE+mXLx
FmwN4rhsMFfiBMNq+3VOnsN4CRedoizpYyuBqmBuaMGR7mrvmU02iINapavte6qNSGc0SYuwp+fR
hz+0KKOGWSYn5tErta7CZoiRS00yAsHWbh6UztllGYlAkA2EEoHQndwKm30eHmqKwCgx7m0qZdIW
22Sl4wcOBYQNP9xsHwjLIh5KF8I952lSl56swD+EbrsqkqXtGXWrLoDc0ccIiLZjBESfH3zNmRZJ
cXzP9g9VuBHaoCwBYOEhh1zifpEdxMR1Ativ9PV/uhCe12VDlFsKkDbsFqQM5aVfKnE9DUW5uquy
ITuW8TN38qbujg41DtU41qeoEHH1s9NmJppdT7QUZ3+QdGE5d0oFmq8Hiq4hLXNWOVnlzgyPMkkj
iIAe0yAPVqj4Ip+LhmTxMLkRxciSntSc6p6/ko7Dv/ImjT4+XohA0t6K+5I2ncn1mcu1tuZBK3xl
Kr9TwONQA27GndQEN6vlftMZ5OTPWhTQuvWSuMjWhiTdfrLkR2P/mgzFbdxoj9GLQQtFX6wie1Eg
OovwyWjz7F6TO2W8Ha6slD72/60lDoU6Ks2RN65qE9E7zVOAVg0bIvJSZC/BkvV3VjiwGZJS/PqB
Qd0YX57nWT9VmW9shl05mJv0KoE79sj2MGa+8+m8E6OZbwfot83P2bUzE7Xl+yeHb1ud7YHSMs33
b5qNsI2Af5tAdlJB5gHRs3IYETAS1S4PMWdrjev0rvRTcgeQWwe+CkD4d7dzo3PV5FpZD5shcfDE
5p7gf6MyyN/44DcSl+5JtvFfVtUQhrpgRjp9l6I2Cjy8K3KMaP2Gr0o5hIGeZW6ahKik0amP6XrP
H+da4T8fu9o4XZAcGBcekXRbZVxxGR+HMu3Z3+Q38eOHNPlQU9M2GP87Ou4z9Xgy5YgbkkZNUqKB
1/bibiiXqFEoxAseqwCfqOXMH9ujLrGTa3wRc/KcfQQCd5hfWUodZ6e8qfow3QROEPgC39R+sth4
H5i1pDgMqxu0soRfqq7D9ZS3MyctmwWl4Biv3/fbiM/0KNNIFrbAUOrLAyO8HttS1EPNk6y/DUsd
Yj10Nq6fSz0JzPY077wA7W+KO3eE7zX0kZE31TCwxg+p0/A315U8U3mYOgY9TlSNcRaAWbuVxrOv
zogGijOXgFrl05S8rVQOHwvH2ExlYv+CpN6uC77WrQnP6coLCGMLWjf08apdErlJqdh0UGd06KM1
z7MdGevUUZFc52mI2nZv0/hzehEQuSnk530G9K3NbpRUF+rczZDzLw2oNX3mURME+pNjapWD5wsc
TsYfhJ7WPoHSB3tFvKECbMq5lG9rHQfsKEfeuNAyY8brXi28xcz1RRNN9Cl7RH/1p3vDGS7pD5uu
43L8K3YX/1DzLB71DzZcpNHC9a7PDmUJ+P9ojr4VrtH8IH0z+rX03Ywz53Wb8DcqmRupbQGshOh7
zXnLE0sueZ7BieMgTPU9taU8LHdKZy+48JUcqkh3M5voH8ebt6rd7IyFVcmli/tHtGXctPLCXMNC
VOtfDe2DkfT7uHxSP4rN3GtbTALbdpIlCWGwsFlleZbGa3J1JDsmmXBK1+CJAbFt2sNXZVKqRd3y
UNtpxMpMR0J+b50xFXcEKhQmEcCBZNLazTUyf0XDZvqG4n2YGuqSv5ssmIf3hXh86JxrE1pkqIcp
1sh0tBMUtibDgDGud2voBF3n5tO0LTg6R7SdCyH47PdhcIt2r1WJtUrc6t45VhoneTKWpcJHFWrH
tibfYHVJPW2WzecPyMPeylTum9RUydoawwgLsk1fuXoNTuQzg3XXSyzd9pwfmY8eaphpplVzMuya
bsmIrM0xZVaGJ/Hcrk+b27NPmZLh0CNZxMws8bpn1JsATJed8bHvAISq+prLxbxShUBjNdvjwq/v
2MWHE1T5LLg+tRwr7/qDn9ryljdhKxyLeDOT0Gfi0/d4YxNyrdUw/XYHwKisApgoqnmTEyY8/+lX
7Vs2OfmyHfpsZOY41AIpZtKygDyQKfixZfJG6OrwDaDR6/NvruLNIchv3Q9YzukmPpxllQpP3o5n
ixlOxrfoaL+xI3bp874eRKrQ+7jK/b2KEasTomAIVyPHP9XT894MhAPpFxtIbYcRAKjsEVaB8Uwz
bhujYjEYWiCbevmXY4jzWay4lMahqk/ExhojYTtQSNv+Y6oxDWZqJTy9ot842fLHe7wCesWFfJpT
RKhXt/FQJzBBnOZF+egt49/CfNiZ+SKmJnBYe+M6F538VG9NBDbI+34ZuqFHlLSmQTDyqz+SMqoj
ACbAnuFtsw5wzb+GkzkjPmCaY7VN68iJQCobSoQDqSzmYDY1YCnRgyihUlxsXmWTNTGa4Nr8Fod1
eUI70m/a6QdpshVGOUdwg3hvr3TT/sCGZ12YBqwECUWB1syJJru/NdoibVHCeCGFINx28K8KIjtH
KBUHN9Hhfg4tcNb7/Q/qIUSt7S1AugU9WgYkr9jB8yaL5QYzfITjKhkvLRU8MuSroGkt/dxFLyhu
1y59Rri6m6/PVyciKiqGRsx7OVKpS9DesBgyfmLkfD17anPIwA04Kkx1iVpam4BZDXa71daichGu
nE6BZOEmLnQSjg6XKfUvsFyN+IEzCyF4BLoFs0KalmRgIcLBTgkU2V4P9kCRFrgdcfPUxwZ7IPY3
QT5vzeTti3hVSe04luuuJPo47q97RGmdtmRT86bHfgA6o+xqNuy3O++T3QML75fflOnmQ04Bejdy
YIrVEBuHSmYmLhdtdiHxhibi8qlvFmfwo3wRoqQYkKtsEZXu92JOpGxW0WRCDNcnst8tXbR2OcDP
1aGy+46cKdTMuTcC0TOMTKUtdcbOd2Pjoia1AFEIDObE5b/05be19qBFd7rXfzfWRVdGTXLQ2Pr1
TVXr72YE4X3tiLt8Hz/TirZQn76PskNYRsAJti7PvjQSz5JhATH11Mg6NUmQozXYOJYZiVGB4xpX
b0AD+RhxLXsvK73/KzBldPQEhgqXwpmz9HSvQqFJBqAfYDVmF0Fqfpifn9V+1B/eosk+hY3vtmWY
nmmBIGdiZg2t3lQcwY3eUUPKTADh57tqMbioQTx23OtuNG22sjlWZFJaJ58otGR8tAuPQ/uFXrKc
9K9XDfMq/y8ObXJ8/hPWCFIpPYoLoNbvxJ9+lTyVF7rRWKLxLPssJ6oxlLGGmLgJNVoqYxj/5WIk
skXIYPRnq3h0xSKodAijOTQHJyQa6EhCQTkhqstfx613F/iURFGQbpz5Z9EDHiU60x4+w7ZWiCld
tEubG7RjWnPgk3+0HuVJxSK8QLTeVg9xzRVlX04U0FFt/+30wo854USXw0VXWuCcJ2Z4k/BIINK1
prBNT/celuPqfNckv1W0VWwUJPYfujZVbNC6GXpO7fXZeIM/7QjZvM+DQ6LtvDsAx6HFrF5qKv5M
qrCyfCoAH52IPFhfEnYO2MvYLiHn2LPfngudwAfabyc/c9rMzeIqLSYDncD6SR0ioDPVZRGU2qHL
sS9OJqtbMaYNxCRpqKVJ60lMiRRDAzToIcZ/0GUgHcYl7zGmu6zODvg2dR2X+T1pqIFV1HyWorwy
zS2d29XRSOmKelECfxIrjzeNfZ0QmXeK/SfV9pV81OtN+xZ/iI307YrHy6Z0RbIwF8wKzwmI8hDK
Jp2MxLovYpspA08wT3q0gwif0mOspMFuNIZj/MInCtO9bCv2cGCB2ZMTAtCY2RoNC8Buu4NIlVmW
XgdshlAGaoiGSxBv48f54vA04MeFjGEDXbtZe8vwdNYjm6zBV5Lfa5b3J3/ipwnuvgLAuwy4sywJ
Dfp9uYmKAz/50aB1/1r15yd0VK2E1uy+2/ILfV7i2xnmOv+Shl9fkZoKwhw1LKbfjCSVi14VGkDL
xxq/mT0fW1GUC2EzEZC5FiRpLMU8xD1U2gk6fBkpvV05bWRSUvLdGLj8poFg2frW1A/o3xgaNsPI
nlCzVMUaoBpwEPuk22C/SKNwNQ/vK5m9KIrZOvR0GXcpKexnlYwxUmpGBFq2tdzp46n7XtM9DIt5
o4solezfYJ4vcXSN47j/denJVPng1+pedcfKBTB3kkd3LqUSzF63Q8iq6/oKR/7JZYvpVcXB7yrr
gTq8PFCpoM63u9XC3/n/AMncEsmG8TFHuC7IY1Bd6AnyLGAQfBZ9793gBmGO0sxQwZwFNNPt4p4e
sqji/dZkv4Lo1R8ozsQMdLdRglmeJ05besgqWYqUfIdR/Dw3qUMp+uDXJ8T4ojkXXGb/xJUcQ8fA
fRNHl+2ZRtNxdYBCDbTOZ8ESsq8/hvOQtAzUp+6LazEVJCIjGmdrabZsppVx3jCp2kgGXqJYVpM7
kbW0Wmb5gmvsxAgL2tgDOs+j6P07JQ2hz0qZpMA/28di/iOi/jUyI17Q/hPJzORdmGku9C2Dpyfq
y4c09YJr3Un27RdewLugKoVkrM8I2gCJHP8iNGXJ8NAj+2y695ZNCDOQoxW6fVDxlCO2j0RjDGUf
0Qd9y9PwqeXJuxlV+00UjnONf3fFQSvNCHOTSK/iH0/X7ung0dpKahRohhrhLExcOsdIZxdxy1Ku
xCqWw5i2yyL8zPP2WkOGzantUSQK6DFZebYiif9rIYB8WQts9jN15/Uuym7fg4VKFOlDvH+6HJoU
0cAypbx1yOC0Pgzf8z5J2iN4zysq2+FQEY4x/RKKIaqVY0RTBwMrh5Pt7DqQFRHDm2/+BlcZZoSF
QpH52tHrpMAvKyLlmRuxIbF8H8UluK1GTLLRdEnAQBsBkSeTnO8FIjPkXZvzfHghSnC8XTAREz3c
MvV5Leqcql9zUaRp/ikGi9kCeV4rOh/gxX1buvm/pyulxtOe9KzRL5zWPIbgv/P8QjlkOZzC1pGP
CxCz36Oqe1x+qQw+sU1ia1WPbrFfLtwZ2eWBvAJPaOfTDYOx30Rx/e57rsQuIMiuJP5iyzHhzSkz
YsQZFTeQfa5HRAqHEie7VJQXmwWrs+5HgrK1m+Pca/gyzRBaZJQTSVc7Te9qk/tr/vX5iHKaVo14
Gy30JHiECHllwY22wsACyLOPEtpdHC1gxEEv26kwSDUTP5OpXYE90XIPsNBsLY4+1/vFuY3TWJx6
uFYCa1moaED7Ob6wZuipThj0N4xrUNI5OOq1TbJthtzdnJbUdqbDse36NM3M9W3hcbIh2l3sifxH
3s+AiT0N5gL5fvU3ToMXNr+ryeuv5yN3S2G8m19MajjG38s/U5BWG61JSUMQe9WRNwuDd/4bLHzH
xTq36rUUt+4CyEWiRvtFvItONTCSPwjH+ibiITe7D7IDNun5ssOuoSKhL+8yB9tKR4AGveyn8+Vq
wkDw0cYh7/vMgJUiTaCVkv1zw3klTKnkIw9VBDRlmGGkWrmAP1mHvtInROcaeed1IIPgCx9iscom
PgUTBP2JjaS1dWEeMoT8JhduVFkHbeIhZCw3Y0Ip8OxJ8UOu1QfpsCXG2IJ4bgj2bVST4JUWJf1U
5wTkfm/FBLz+WLoodjDHeEErgaw7iaOcc/P1WziKPGg3E3al/zJkeOYF46BNwuBqX2IFGjneEbjD
bnoxliemi51dDjXgz5b2hP63H1lxFbE1SPHF82T56bp6xigGCGlP339s7/8zxo8KBsDw4LUrp+si
AiH8g3tA8oEWvP1l5wBWHS+EQl6Z1ZLRMECYbq/QgmFWzak8uQy4nplFWsv92O7k+JLPRUIwAfyo
xurCkH+mo2mrXKnpNiZmcAGp7QFq8/em52AK/9E+Oxq9HSFYfifTMBQ+/o546rotngQiMQnWsbCS
mwqgDAGmxjdDuXChKxs2X8lLPC+3xwaYar7u53cKqSZq6kbMfpBHsY6t8wDl2IpaFzRZUwmfuHgB
eFabL79aLpTNN7vnuQX8ohXBmPNzz2qvVY9/USNMwoXdcN04NxcFTMTU+ilO6T5FlKQlu0AgoxJQ
g7gOno6BZqo1Nir3XVkCONGmFc8DISZxlKCQhvbzMDtm+CJPb/FC67FzXhhfPdK/xjc4LIqs3lFO
z9FX1tMfYu+kA5jw2gHYqT5JtzrmlLHw3HizLr8xQQX7VwnBH8sljC/xj+ySO2L+edr7R4q3JEYO
YebGZWw0nOJhDQdFmD2/xvFi8Biip13yo4ivTL/P2fawkUsTA7gaqFg9U2aGF3sW0Q2YLL5PlBF6
VCJZhJIvGmKA1V51Xhb2xdYLiURz8k1ovhGioffIBQM66/VwQQGtg4X9A4gnRtRrFaDOgwLKJcil
KfnRXMUIdYcqKsdpS/mr1wEBEMqfAudhCM428czJSXlT33E8OgzKw4zylXfpu//dYKzKY4uJaEaI
25pyygI4nF41FT2DDZY0BdJN4GG38PYepsQQe5Ybgw9aIV2V8jwMgKjQ9Sdqj6oPzH6oZ/GHRphC
aVG1BrPUJDIG2f08G9CV7zBGgNV0XSewEoaiXwrIhDZsslQ5jtjiFMrxNKXUxHR3WZHP6wePwK7H
UFL8fiASENZSnMaBKQ2VJvbFKKnkS9ZfgRvvX1M+VVe9b+gu57fBmIkUFyePnBMZL+D/BKvWOC8N
zvMMmKo33MLlT8IcTFSsat0wjzWfEF28JQIC8h6agOzGFtf/nP+SLceJ9RyQ9MUl7pzxRU2zq33i
8dQF1CABJLMNiV6cuhdGc5S4I6ZbZQkWYFan+ZXEqCBamiqTkkaX+XmKrYCSzxsbyAWU22YbKjuH
gXmUQpVWDS0ouwth26l0VgUcd9agn+UknrKQM6gijdMP1fYDnbYsjaj9JXPTjS6p45F2/GcBXvfE
kvlmlEw7zTUzePN6evuqPwcs+CtCIURlwqo+AB2+SsouM6iun6IsEH7O8CMhKqwpih0Rk50lkcv2
7mYPsuKncFSVWV1fD5ymfOTcMFFfgcTzB0zOZVrlPd6ST7bLg9PLil/v8jZ3OIaJUPbiTzYNpY6N
V4gsrFurLpbxVQ5E2ICSxa1PBRKv9FiKSf2+F2xYR8mGMs7ubFS4LNluSoS28w2EnihdUOjtSaEt
ps2Pf+P9zORbi/WklSIcJfIEz1PiILaBil4OTzPg6wkF2iBtCoNNMGt1EWUlxPS0Z63YtuCocffY
wlQwKXf2JsGyKW43vphZs9k9iMGN+HgMDdaeruZm9kDIakqzrCtXzqx/7Pd+2CQ5WiFuL+OH4VDo
wtkdKao9Y7euidsupgaUz4jWH1aR+EUxzztn1uCO3qHO79pIBukBW2RNzTsaOK9d5et9/L66eo7U
dGVGyePfKLiGLE5gJiCH51Wustc5BdSSbcDukT6E8N+wlEGVD1z0xVzvWVgHelj4Qr/KpHk2fNFL
UpBd8gcACbapAvXj4bIiNn6RkDTu5Wjt3jXiikogyu3K8fGjz1VbLSzyKGTk6j+VgxefFDZcne6Q
w6H+QXAtFnF1qYAL+3eihPRJyZAHcQEHCTI5vz96WD/TvkXnWhZ+9qjaQtOTE2wdMur5PJxDybY1
wH+eROnpCozrT9WU2LaLA5flvIGGbHhTaq41fFG6LNY8BHlZAxvXjjx8F+aww1cZ/rM3uZQ6aZ3s
7fcgNSrdoIAqdoz3RW3MWIN/OMGgCJxl++55hwKkMGxGqXDbG8svRNjq+c/6xTReZhNVvS7r7AXJ
Rhjba5hRK5xa6KGmUkB/0uuC2TG42HV0Fbh/6X1ibCr7ArsJ8kuO148bUI3H6kQUr7K+Qvf5bMeP
9bvPCihojriwhdOZhGardmfNE3v99sfbeP/0IZR7raIkIGldqAQZsrP0JoAAzILtcSRoq9F9+2o7
Prqr54YdxlVFBEwJVyPwb3p7Q7jv5FgZwgnQcpS+PWTFznGNH9kHDZhYyX19nKfeIbmK3gAbXrmy
8+Sjw7/CoQv/9KZwevkPxZiGWeqdNSuD8lzke6SvoynIqz/NLJJP2TJjj/jZU6PCKtmNCzK/OTRF
EkH06j7MEP9JhLdK2/+J7pWwPqYfEN0p6hZTRPX3yYUUfXazbBBzAzdB1iUBA8K2qVo+T36I7F1Y
9nb5yp3DEVjJ9xaSWSoKgUZml37ZD7saAcprB7yy46q2XA6jyF2YsxZ2qPtwBa68qNPH1JVURvyu
/udvTRyWpVv23Y/sGuqRdfJkBqrZVHFXLGr43r7CWMUHI59p9W59MWHtWVErsLQRzFfjpFcQh5Un
Wip10IgpYjpFbQExIJqg5Q/BijjePoZbEWxY2J0TbFG46zWk4Fi6TiuceZccunSdCtIypv2kqZ9x
i7gezYp0+QbMjisVwrc3GUpmmsZCXGHbsTiK9EbQTT5TtHPsG98XqhDrVkb7rDNvTsZksLlv0l4/
tUMjwbeflTCrlyUi79O/JjQDzzmmV/V0N2n+2jJlIw+aLDie0iVPZ3UgcAUZIG4VeCqMeqA+aXqL
87Ro+ZicswBaqY7Rk+7xA04QOZPcFmpzHm1UWwArt1yEMFvMWGPjqqkLyeW7y4TQvSOnUVtewcYL
CurD6uEb2IxX2DY5bDCH0U2WcS4ubp7RME2LHQqymTwAEb+aykAzyLoxZUeG9GnT6vDiLsk0rTXg
3ERqPNrM+h8v5COfzaEf6OGUdd0f00ZHf2SezTULl7LjgF2H8xmXmSDUwvc0DlMtfybh2h68deV8
HosP+izaz01TPZPAbjuhxIVXa0J5XuYYw2TzNUy7fIvdwQNHaE9f9zscZn9JrNAOMueUF9crlwph
cGN4ZpKXKcQlJCnOS4lkHfM4dzshhtJxF16Znmu68cAqLzcNOWeO3TyZGnCurDO6lW0BMTOOIsxB
UtcXl+CNoo0gUpZ6nya0BeOiWnogufLqG96vtDcrc8CB/zY6GlrCB745XunqCi20vTEsBec4pJaE
AVClZEK1EHJ9t833tBLeS529MrM3TRf47gHvdeAK6EbS6yVO6lDrEe6vVdQx0C8yGhilm9QTXdS8
a0dYQTbMc1mCrmkIkps+eeAB/o83Ni3U4Cwg2NyLyEnWuTjSM0nDNToOcfNbmJFlB/yRlk4VVH/K
bXkeaUQqSMQrshD78DIudrwCjF5cIWwjDiNY5fxAZ8Txbj9pQsvVz5+Lctv66OeqhGM4GhMtXFZ0
xYS7YdD8rGWRAQb7Z8z+BvUvU86geOuE93RFPf06496+3mTKsO6jn+DfcMsVqXuy6D7rbqwjM1dA
dhuwUOwZy8csxBVsVAWSj71+JqeyyOluZE9m3i7pvLkfE5ROrZt2LtRjXJJFYIK4HqPx3DZVTp4Q
22dM+E78Jx3B1tfumWg4qpes+SfxUhVGo0Doa4q1yef9jB0gIMZwpKU2aOzqWBgqpGOrNnSoAXfR
Ma4oMvLWuy4FqQegMtT8deJquoNiK7yBbXbuw6ZDKrIONvRMbAPPc9Vq5EcJhXEugSXk7ETJtV69
nGNkGBPvYavovLPOcg2+tEDPpNJySvCNRB9yDzvfPkscGvomDur/sYdPwhG6DKbTUmJWVvnksSkl
uJUdK/uSRCCMJco+wUrerzbCYat8MyqLgi9Qljn/ig9zeXaz2sFOYw2HmcN+g1vaE2bVEImfbhPF
NqtBLvh+sGSlXCNzSJ2wyDGqHYBY+Izoiq6olLw/QsN9dwaXS5otv5qm5AMTx21B6yQgQvPSa+Tb
zH+TeIRNb6/dhMmOM4XbDJQY6OSGKYxok6fIHIH5RVqjl84xLqHWfA+8ie72GP+aOOcdbrbStp3c
1D2q2xaFj0x7XihnaDaNa2tFyuUdXR1JAJDb6F0KAIwY9jw1+7qdKbHIYVDWMVahTZnmVjEQmmP2
/7CeQk2+UmbgJ+qFQqt+9u9rhmoUZOugA2BW8UJ3HAmUnOWQ93JGbUZr2Ud4cEVhu9tkRx2UlpkZ
aw9xq6LXSj/pwkUTdCBSeeC7biBW8DTttI55mkVAtS04iruT00IK5Pl/ZBsYBdsP/JWRS0VHe9qD
zxtjF14lYMIVwwWI0HcN1riz2gyowGE32dmoSaqlZfv9L1oBHgyrMIyk5bnAS5ffbV5D2zzG59hC
x9XtfE/xt1mr95EbmxC/qLoFuTVIsWHjeEGhlDRZkHLYdK6vY4NS0d5Wwm2GgkSnSo8vNdWlTQuM
ex3Vh8Da9KyqKk5nF18xFrNs/S4+jvT0BLVvKTA9hn7SI54CVUvv7lu/EWgaKTUwgUPaDX1R+aaG
uFKuvKEFFRccC6dMadmZBU4NR1daCEKFY4n1Q29dUl80oorwskxs/erMCfd4/W7fCP8ElIhNJumC
wl5LGC5Y7ogPP9Qq++1AgeWPE1VXdLRlAknEqxEpHS09Fiyf7XJU8LGJZserBeDmuklJeQIjXjyu
WKMczNdjbDQZqD/Y+KfdUKuX8S6CDlfUeG3bxCo5rtxU4oButnVKffdsAzvtpTDX1b67kCYk4+Eh
mzPwYzci6FzUMj0bTJl6Ij1oa7Bd1i3NTXbIRdSGXULVwgEgqd4Ai59/xnDiNL2OMT1O0oZ0ZWCu
mV5Je6o3IzifqvyN7G4zHyFQ+YNnLlbv5ETC9SiKP2f0W5K9X0V6iYlmNVODMGURbSmzGiBCHLOj
thFCchHfnd9GQXhgiOyWsGATSdDsfhvgCt43x7QcZBzw8Jt4jggJRmW+lCR+RfpKCM1HXQa/09tZ
lrkAUDElz5zimtquBm59ehWnatzqG3r4ROzNziQxww8jf3FPoRTbFBTRA4vk/LfzISNo57/cDZ7Z
ol+pWwBJ3Az5HqvWskcOFytFDeTTIvV04hSdvnQ+vxiCa15tE+jB0k8NmkdrS9JKFLXXiqv8iYFY
lN1hlq3GnYcEtkZJGcMJvse0BhkhGqxzU6yfJ3E2bpEG0J6vDCeK2yybOGGxZLUXD3Cp91cxPiS6
ZxhsVIrg706vJeS5eZtAu0g6cxcVPyA+50mtuHA7MJUTZQOUzqCkwpcpCAWriXhs/J2IBcBH8/92
6L/XvtIGf+CgypyUg5Ez8je95jUCOu3nRdWqG6/rF+sgsphJv8e+OaxudcTZ+CDEnHw+rUqYy1+C
/WACH5u2aJzTjstKsNyu2vISygf0VWk3NB5XMjPLSub1TbhejMOGtewJQtzGltOnAb1c9sCdzKtf
ZwnQpgANBg3ZnmoD2K0SkC+AKc8xInopjOe3BbZMpipYCu0ItziO5dbGAr/LTPujrcalDR4Fstcy
XvCzIxeG7PNA9drfSrUC1Lc8IbZE8Uo+HP36qThralFPce28quoz4nA6+aELF6oPikdWKNBkPY3Q
yNweGWJ73maEpR6XF/RN5Pm9A0iGtF1yznjMi9QA32v0C8ZUL0CFEb+axeykAzbxiKrF1rQ5Q7nR
9luJVj+9JjAshIoQWrxitubFaterLOkdCXbbgCFFg6Y3jIO2jxDk6IwNoXi/IdCln5rPQpp6yv3F
fuedg7TiDCcz9gLX1mLrDoflsNGZS++Lt4RE8rwK2mjXIRGVD13HjeUv8zRLaQRxs3mQZ8lRp888
kjfy4HjpPkm+tknDfc7KbaFslfNgCv8EwHOtlxY7ahjk11j31jLspKD6XrJag0FueBqtiamJGNCV
qhjbVlBIZS5qwvcNZ8SVK3FX+KN23X6DH8bcAfev3Nh7YNIud5AyM3Al+BZzCbVks3dD5F6fOYR3
jSipFEgmUd9TC3BJpb86f2++C+f8Cc6pPOHmUf34ptTXKzc47K9o6RZS00znOvQjc3oXqSbvz6cs
KeMQ8ofmmEFaHLUjOPUCKt70RDme/yi7GUDBbyV6oO4Zrz9x7hF2FgVDxwulDct8ZIt7pTQHenQo
/OT573LC2tcYNhekeMic+jPqy8vswrQq+NvXp1fY9hvvdxpMpRxbGYw8dR2pZieQVPEXwYGtDSwn
RtAqUxuKrKZFnnt2XAfxyFP7NYkFy68KquRogIB0M4WT4NhxSPqB5tjOZ4f37CD+UFcSKrKn4ySh
Tg3e6Eps34fgGwPq0u7tbTAU55kRMB6TAFDistiivg3NE0w/fPx8DD0Hwoqjn72V9evhZ9pEyvwn
5Yv57uwS/JcX9pX26YPEbBviWuYdlqmae7KTeAXATvKgZu65c0mffV7Xq3k2jJTPVVKUpprrGzMz
5a/3tTwf2oj0w9SugBi9yNRNjJ31QME0u25Ooi8Qy79o/Y4NiozNqcBAF7iGFx/vHkAksSzFCwoY
Q2KDd4seaLj+zUu2/jkqNM3SlDqGYkL83GtIdUEIPN1Meb3zRUv1Fm+RNkHatrUk59tFYQz/9dpK
mv68IrAIp/10n8BzecOwKmZGqP55iZJ55NUc/s4f/z4oMz1qPfgjBx4Pjv9Qe4/cQLUPZaT47YJs
Ehgo8EmOxjbTTEgnFlnuGMZgUiOURonS8kRWpmjEyq2tOmVbEzdSOup3tE8TG7l+KV5Ss3gcz8ji
kgv7pURLcFRLDRUKcmmC4g53D4dNA/9JMKJqhIz8dut8u3ZNuwMmqXFru/niBpyzieOI8pZMa2Fc
Q8nFn1QsmozTXfk/CuJDsyvGaqwaRKg6hVy2Jg3bOe8Yk2gpyLv7eMJFcLN/X5IiFzaqiyq55B7n
mdFQx8U4e3vGUPcyGvQbOBuVLMqF5tlVD4tjun3t5B2+KS5WtAgzBI7zyt4Q79/qT0QzhdNISpn9
d8CzknLHhKwBJ9sqMyGlmZEvVhuc88w/Ff+t23yNQROT6G1laTkSyO9tfD9KeK2V6em23/rd4eUu
+Q5qNPj+7n02nj930mq6vwgSUQrDyuiVzToHWq7TtogN4xNMl40jB0w2CKL4VDSqOzOKnfUl3g4g
TmSqtVIAb5nvfOEqsbigT55ki1kWUzCifWJhAWVbt8/itg6fcaGca0SwoQXTugWDrNYqTvayUBnc
yhKuGJ9nY05/LRuRJW55zaaIVn0WXbrH8ta4Dtya0j4mDIwIbNfgW9cuVYPGlSsPeNN59hyeaHIK
2paIAb7gOWYaDZ/judD6MGytTlE86WfDRR2pv75thndcfPPuHyQsV26BkzR7qTb2bcAOkcB1eTfZ
nfOWbXp8jP0XnGzA7dBpu+1zvMkxzRtk0cKgDnNKsa6R2bCZ/ibJO7zNnkDAUiJkD1l+++n7ZuAe
ggFU6TFa5Gyc40xKlOBvfQpBA3mgJ2yKAg1k96FZ+uJUEB+zKeGqT0Wa9nzWBh0duyOUkbbbf66E
RUmaSKtyFj0rJXNJHgtkhnn/KGBDC3Srv/GxIbl6X71vv6gU+grJXcnwN8LaaKr83lUrjp0RiSAP
5iSXETqJIcyo1jqBUs+bUIV4sMZv3H18chb+9sPq/6SmANfPtdGjIJkyzp1sUhgL8wSLm2TuFXhf
Cg0/qOEfIvu7HUdfUplYPOogdETd9z7ePwjS74hGuCm1bS3Nl1OQAGcj10TOIGN9OQeNTR2Xr2xC
GCL7hULRlG9ICwo2bPJJxGHp4C+DcKxuz2wFRCa1adt26zwJDdGfQ8TvL1MhS5zxvBOsgysSbHIc
GTVv6vGJMVmExffoJP/u43FH85ERRYGfrD0VrymJZFSSlmtFvIpeneXgzkcobxCWy25oPDWVUW5X
vpY5mcOvV46dr5k0s9sgjBQR+GCQ+O7dQMbRrcCBi9qA1LEViwMC0YbFK0+f1OEFLtSzg2kqkeEZ
ST3D1sRu00x3/ydF0tNOg/5qHZ0FBt57jxmgqLzRXXaJbS5mXxe+FOpHEZNZeWC1g+NNfmc+OYqB
kor7wiyvzxpWAvzJl64UJnq78ZPWu1Wm9YkvtX9znKjUxJrSGKg1caC5rBHDNwi4l2qKM6EZdy/J
t+bhVgy1YIg1TkhN9VagyEptcmKCdcI/oNPdgQjoAMuJJ82/FYu4GBe6m2uRXx5xvo8s6FuD6XFY
V/7dfmOYUBi2du0Xk/w71aplSoisomC2KV3UhDXioc34Spb8RrwDqKEEzA/IaxmVLvyFd2Q6uGGl
82dnusj9Aq6Xg86W01j15FxpysEZvwlAnpjRXnjr2uekRADtQ1UdKpXN4PUfJj9zGZsZST/Q5aGl
gNdpPXkCn20UYTS9BKHQMspK3KtGg2Tcyfsy46iTuJamcrs/QlALNuB1CbYbOypvdDBmz2vbkZqz
SJTanGqjqheKzIYC0eVIrNo7vBdDeYGUrZygod6DOrCrDvPYU5LPJWwk2E07+AHvCsFNa+zNDuaD
5+ib4nQcfdboinKfm0lQzobgoaPyi/084AtpRQ1WFTM0eFb61cYCvAlfDIbnE+t6vQA99yP/kRDQ
16v8bgcjpG+8NVKt8SNVCCqY5L+XLzXwhIuWqErxQs70h+LjERbst1KiItXmWIUSF5+Z23LiUWjd
fB53cdHbgwnwLyfcg5xzBz02Q+ZQBekGUmPZdFTqOyqUwf8G68UzEMs8HVEIYJBUZFpijn8shD6J
GGcvgi5YJxvd0bGUSRVgeOS+q+HOQ71Fntz0XE+g3LLqV1x0ePLSfJpwLK7HIR+n+Es5xYY/WrTp
CY2GwAMEMpNLoqJEj3dcsVfeI1dlIih/4G+rNL+nwUDFS5sQYM/zxh5BnpddipTSGRzBqLQ2/GlZ
DgjKcRW4jmkHPhiybQXy4hWVsVLaPOHamm+iMUuH3EnUXnNT2YWJ/SSIj55Pe8a88eao+kRvZ/wa
VkdsNcWMzPJ3yA8GkA8He7SYmTw+5HmOZ6BIvtGXgKVSaEnK5qGUjK5ugZ4n2gePEC/hu0GwcwSN
tVJWEOhXxUBOqdWG4c/wRtejil8f17KSb1DtE/8EsJajIXDNG4iPHckvbZHh5wm+pQpWsYx/0fPC
hKkMo0ZatXSsGrRE6woGDsU4OaxmZzoAPDOJ2sUsl4KMT764h2wmz2cMRUMBJfGdkYCJjicKg9IY
82X0jB++xd+fbrnbkiGFkqqnNyIG3nO+hTJple0fBLigTxw0OYxhiaTZOkTWlq2NADGacKOXIYoR
35kzpKsmzM6WnzfWUAe+IFQHtYxKQQEh8+XhYRinYHguHSzZTN799BHHyzyb7yQ6wgqdmcKw+eBI
jBBZmdBweekdclTEDcljSpAdMJzUzeYXS4lcGyqQYsWE1MDHKp11chPc8Vbg33pS2D4eKZ37T6t/
hiov6GBjtw539hZjIB/GO2/u3L5E5eW7orb4EzA1a125aW6tuUz9sz/VY4F/pQsnVFIiFslxz6/V
hfda0+sYBoxfskLIFzhnfMU0PPdPNoytCJobQZTm3PQHqNCagSYks3R4OQ/xqTE6/9RYN+REHiSo
SWrvsvAnlSWrd+DlthyXGV3vKXHQh/Otr//dM9TNOr3Q+zgnu42uSbkmd2ymY068618C6KnfrR6/
u3phyhVzDqDcCeTJ4nD/KFbhyqA0TXVH0abkhtn+NjlqUjHs1MKj6S9J9Fc+wp2EskG0hwliKQcu
AbaoYj3DqjA+UX1Nlxhe2fELW27KzDPNKwJz8jUwgvB2VS8tOI1YHZnpOqZ1lGBFePlee71/FIWI
RNleTDmk7enIzQX55UaB3dQdEZGlwYz/ZhYT/QPYHXATJaxsypsH5Tezy0RBaIwuHtP23xNnzS1q
8r06ncn6URb/TZT7RbPsSzYI+jQhh2cm5b2DrglrQ4uUqaP/HnOOFSwip2x/XnFdAo55VsJoCFrK
he2a4fti7F/8CTCiihNDBC3EPzYYmXIQMS7kCgKlm1vPLmtSN1T5kDgJpm58jXROd7mACaxJRtrX
ViWFqM0QZg4l3U4w7voXHI+AmGQFhL6/733Wi/quxaJnNzp/YxekPMhZcEh1zToU5bsonIARJePt
6pC7Q0jmIzn0/GVjofJ2snwgboDgWr56QqalA/p3KUu7p1Zy5vlTyEND7C0VayvCkYLyqvLrciL9
buO2LrKC38WVnFcZ86qk/lY8WuqyUcwuISf0McSYjfgIQpqu/NHIC/Kdyg05GsHzVDRebv20WPBC
a5QmYG0WCxnZDNp2k18Zyp+65CE6sVxzdR6o1hDGblWb/rBlPqZJRZ+tDdzSeDEL6qNQDfmr80QO
IN2RG4SVI/5rNyCGI3lHXN8iK2NwMxCN7WVo3snZEKlieGj4gGx2th0I+vq5oBMpOgnJG9z468UT
c3YxPEJzblAI5hMkV5hfm+9JAR3GlmHSyeefGBCZkGUC5SK25HI3gms8y7IXmX4m1uTSz49ePtDj
fRlKjKK3enIf9Y2BDW4E3E9S5KaVjHUfc/203pDca5o+NEa4wU45KDulTUH4pIBe9fgXJ0rk41sn
n4sVRqYtVvS3TyY0Te7mqxFvzB1vGxfRHnSVY6Pf5+NTaGUCjmeeJOFCm9lw6p9ABjSEWlqIUMba
OQrwRUDXQjFpblMO96XkbWRLs2Vmji9CZGbb9hiUj86uMKd2qxmH49T6M3mXjkvsLGJ6i/HJO0LD
qk1KRL7yXiLH0qnmOObIpAydDbVc6XozwoY0W3mC4MsGy+mV99oNaF5h4JL7NNR2W26DGEamqGjP
NKBSOkAww4hng4RHs4u4LVmJJNGwyI5OCmYpHcNI+9xh3efhzH3VzqIMvqvvLGr3Dp/5ZCy2W4LG
4xXrp9ZDkw0ZsZTFWbhr3XNAIz9bBTv9fHeB1KrbZqU79Po4DxoNiVtr0Ga2ZjVstJ2Y6QZKvcZO
P0PFGwg9Fp4GNcnysO0bZ3OReeA3vFsoF0yUr7Lk/n3dcWSGGFyynOQd0namQdH+FvjQ7U1VXJdP
L3e0NKBbLEDjfzlXqEKki6SlUI3jrRXyb92/+ORYjUD2fTuts2eKoZc5po/zG2/0P30KM23duZnX
0GwI5d4YYX9XUmM9afsrcRP0b2cqP4OL6PUK880V2rgv/MYOA8r71K4gko64qj+cNcyUCEXM86tL
WWJBCI9TmnIB9or1Gdmt5bGWzsRC/RYy8smgTxOkeDxZ5TVXi2BiBJcfumhp6wgD3yVNcY4ZU9+M
Y4eH4q06oAAYBxgPSjtxkvKeutRm71LE6jkwHiOG4EjOJCd04vc5VNnHzVKkY7v3Lbtz4zaC0GsC
NQ8pHM0SkBq8TS6+rVJQjygRzwahxLsT90X8is0ygHkzcUesx0K2hVytyTFpHweLdZUFLLCBfPOj
Iqq3iyBtNfTIeHHvI9VHNgPuaMXswtqbZwR3yT4MoZ2KuFnbdi53YpNLxQmHUhAmrF/iwugQ4C++
OEqaAcknDdsCmNZ4XbWkfY58seuKBRxXpK7dRCa8FZDEbMZqQ19VR2azmJ9w7EpHpr7OHLMKomkG
2HYNsp9ihdMAx+jkdBmCkUPamt59oMvaDY5A+GrXdGKd1SFYvufs2fBAWtAbmDt3rkE65b2nqGBi
2tS9FprkaMDyAXWzUUy/eV4WDQtbGz5dMfZTs246/sxjstTPayWbECLczRpjyjcwHM4qg/QBzbB2
TSG53DK2UzRVH6HQA+AlnbB3GG2QpzredpC46ACt+p4uPxr6pc5I7lW/MXokWfy2VfEmRwdq5YhO
3fA+UB0+zUhJ6zmNbm2JX/hV/f/1yH3I4sjuTH3fEAPq0fXA+CE5+JXn5kYiuMC+zzlOES135yAq
NFxJI1L4GQWj80laQLKiPak5cGfU/tCDxfHYcWTPnzRVpwbXCJsGgN+e3mZqoBQU2rGX9ixeIilG
n6kjtdmHRi1EdSK3wsnCkTLohFAd9F8iVLJv5LpnHMkwhy36ck+KAjuE2hI5Roa1KwM38xmWkwyU
8Lar94xqlIQ38Oo3wIwyirWLy2sCkgdZntI9aHRtAySc4OLa0wonhDNvLJ8GD1hWt+Cci1IGvFlY
tGzvhHbMrd7oc28TJWKJUqMI7yIMhJiKHRQIb7nPfGI8MvFLYJAdjkSn9ers6EBqnH1Aqd/TSQCf
i/IdlB75c4VmmmreOqjG5c+KuaDs6y9gBiZ5ZvESbMUm+//I0APhV0wHdjUd+oYQAxZoX6IuDj5M
MK10Yf2jHmo2zkWPVUK8vdyCtL5cQbZdNNK0/MBGOzq2CMjKE9g2QuN+PvXqLqfzqEazfZwA8hQr
odnZAGRWcs5an8QawYOiXkKCy3e4Fqheu+ISDtTni1Xp6yCiiE5MUsT8Nkc9NLoVpXkNDe7aOIC2
5cbJ49KXZo72cF1aGnxuJHmnc8UL/rgfvG1+SPPhjFCQVClaik40g5KXtPAo9ir594byGM+VYDzx
OS/vt9x8bUBRPBYWhj0otorgiMH3dBBgBWs6np3kSGXwRIa6qJbYor9xq1lVboyZboHtrlzCw+cq
JhGKMTvd6/bkjpbiqzIllBDqJ5PLDMd3LAWipbvCzHboIowD9hMpaOdVnfuCLFiUW/Q9Jxxgwu1i
imLdKHIoO6Ie8Hx5Pdf9sosoI41nV6y1mnzyeS1xcRZmNc3flDCWLQZVTArtKNk/+IXg1tupsqT6
xIjqog3JPRhBuQbJvIMpYOQPhLlaLmcKOsSdoYqFlrVSeMWJzDOIZEDSaSELLLGyKdaNv+1G8HWS
2dqKe5K7xrQYR37PKA3otWVyuqfLLCmZiz3C2kSa2iaR4zM/e8Go8mxw/1TOjqBTr1NY3VWTpb/+
93dycOwtP/EkzWMWx8uqLXAZgH6Hcx45qCnz3cCclBPZJ8bTBWcN6YXrnNGtc+axOTmAsswz57ow
HiZt2JlqMWHydC6LQhyfz4MLsQGxym9N8juNyP8AziMrGPe0OpWZAMzlfBni39d+c5pNCpXCqITo
7YRoEPRTTboCncxi4v7kTF+StdtU/JxDm19eT5pRwSgTBe02bUqBtXEMPyvyfat4jRon3v3oSmUq
i9G6cbjhR4km9AuhQ3J3vsRf0Y9eSPxifYHOpMVUaO1aay4cw1/s5k4gLqSrvuB59SB6YDyr/fC0
xSIuBsAh76Mt/7hgQx+M+RWw8y5CA+tyqjvkJFm4T4crDHxLuBzj08wN2lluVdWhI+1eiaz/KQDA
ST+lhLQHnr4grHjM2WBnYYPmi3r6w7XxVgUmmonpvQahsZGgxmh9EpZAOIiqiKcDyXZHMch8S1TF
B5Mcxs3laxnEBz/Cz0Y+gFcB2xeasnBk7EIdpMhNjO1Pa8TYme4TDjryZtPEpkhAHrU3ZrEP/eR4
ubYCjn6qtsTdjvPNdwNWC/QYzEDSOtryQMKK4DKaZHSVDqEvmXbEzDx1cI0B2Lk0JXAXGD9lZFHD
BeDKNGAOrVP/0fb5DSsl8ZWsTxko8aZiw9zxNIKpzIbrjBwpUkIsuRiV7woY4Hnsg39zW0Bjj5cm
pF3l7TaggicyIefnzhYM9s5XD2Bbc0rq4NXtjzyVv1z1ox4RFwSkZsgtcUU+qSgXo0b4dKrugDS/
EPLH7HWUfDOJyGxeDzETmGNmFA4fIQZBDSdaRXF4gtz2KTYhIOLfDMCiXLl5S/rFHMwyCEBvt80e
IJsOJ1TfToXE/MNw6tsLsz7djGSGrj2x17hy+KkOqy49lQvbWFPkJgDgVlOt5h8MlY+SHUO1mBcM
oax7XSf1VUjrPtPujIwSmkfaybpgg1wba/1UJuGt4ESViRFyF5r3t0l9zl229pLLct46BrC/N3aK
WPg5cHTSnozcRuxdBYywXl+wg6gfvcCSvrxDmP0J/fH1kp23j65ECLN6ekmjB1v4qHieHzSzoC7I
6mptf6dzPccSU+8SoqeHCCEiaRILYccVymFRdyV5doNEhNCTT9j579PzEWcwTjQdA7aQwDMH0RZo
wVSoWmTkQJDIeOwKHYSphylszugd++Jpzq6KpIwHiV0YzG9S24f7u9GWAPt+7dO8nGAfJgVWs8hT
kFJYgp+qWBbj29537wJCmZ7enNDw3Dx/qD3NtLXdq0xQT2jKaFS/wS3tQGFzhbh7un4hsXfB5YJ5
ArjPkrX+HMzkp3FJwa5+ky7YUmb1SocNdNaU2ViSx7uEyram8wWWBrqVFEyFttyI4gjVKmYO/edf
FBMpDLsw05K9vnpgn+tbFYLMbUbr4MNt+tW8DHeWJKgWV6ifhy8nU6zUehhA7C3DG5+7C3AvG78s
sLOzrmxXeRHpdbaeQ4DJrd907t+wlwNLUDer5s5JExy5ubJbpJR82oNnlf28q00IpyQqpWqDSOJC
X+G1ZaCnDOXFzoYbuO4v45Vi0cKzIJ4qovi/mBgqxFVWNYa4RrLoVJcN++O7K1HgLf+XLfu2iVlx
g/cdl3pVflRI6xqWtdcz22LshCX6/BTI0F/p3Lca4fAh6Mc/WGdlpyK2m+nCVV4zLb9jppHw8/BT
sx7nKuS/mZ+8NabAsE1HQRHvOpN3Z47nvn+DQ9MkMn5inwZ5FldxBxWA5ODj7ryOoTggC0vw1nZj
l0ML2+DewKRpBMQFvixho3ayruwWYIQwUw/k8upojaC3U0cRJKjtpP07oHQKkOoQ/QyNujv0IJpF
q7Ogedm7r//vSxUMAawMbXXm/U/bzZmULpMet8f6z9Nh1ZtYHlrEt3ovfVyYgcC7U/yVhVK+PUSY
PG9hUW6UTJkg6OIPcEH7If5byu8LGli5oCCTOk+Z6Zk2elQef+5uSWQCRJIq4Iphqq/l8GYfE4yV
jStIYYnn1Oxht64CbLVUKwL4zWEV4YDexUdROYqX2ii07yRhrII51O7YD+6PpCwK7TYSMJNAg8bL
zy77M2XvKgSiezFf/B4XDbL0I2Fkl85rKEytM0zvlXYmCgR726ligyKUiZZ3nWQ1DoaioQKbVjoa
c2pWi40x5NU9kPEW+5bEP8ATbfhL0X85Vsa259iCSVhOWPb0VG6+w17CRpEZMr+55Za+O+4cdkE6
lbfcmjyxdM8SKnwPcQgQGP1UQyE5XTAHmKvIdRic3oW1Bx5dcVoW+oJ0L09uvOZYp+MSMNp1ZJ6I
sRAhP6V3uzhEhN7RzklwX/84RH38ajlhix808jU5zLR2hYsQnR0mra7DAMQL7UyFVgtgmOvh3TJ4
lq8D2NCgy29yNZWzbzE/1AFkylEc10hUT0+GFou7+sMmmgyvWqtprRwLj84G9ropgttb+X+hHnYW
q748LBfl4QTEBar2vflboDqJ1eh2mp1TcOe4e/zl99b0LjSUdnwLisSdhWkK/m+MeWsZGbhmJI1Y
IE5gDKejjYOAGAmHMyflFRrw5zugjz0p+9HxCKv505xQHvKQwcgsYX8aHUFl03g5j4Nke85GigDA
aQI1bZECjGviRd4EtU34qcclhr6tefBDi99+Oke0GxYF2u+R9YtuQXNSUg+pN1akYhRLHtBN4JnD
BKrdiMIsSqLB4YitVJoRywH3fwJ0T/v7oz6mKavaJlfP65l4Jyp0FO0KdFJPcklhbl2dHnznbxG6
g0XEUFjrEnpDxKwoUVHjQ/EFASkkLNR04FdaHXPeoMhAhjURfekJmJl2MZHCpNsdceXNWhVos2XL
8/6AiBVzNnhoQLfufGLGq/okaxsjs6MGFk2SwCcSgNPCxIFijyXRAswUiXQjeKXQ5u59F8q7kb/O
6raX7ex48ckXJRfqvaeX1if8dTWlMprOv1flqYGq/1gcWHfHfObb6jppGRmF2at9VSmFYIMU6Dgr
Wp49FPU2XiNYpeVwcBUIt2kqdIuLvmxKeA86W9ESWZVa6d5IpUS+esMYkK90AfTcmYflLfM/U7l1
NY6AxhYEM45MGxIS458ysrmYKfy51xkXkFgsexqsRLK/kHC81j8QArnjiJ48J18e+2KZUg9b7qk0
7LiHLf7wMmj6NZsIJdLGSD7MfkLwZRA1TgrMBUAZpmMBjsQREreWrSi6PBIv1rFZQUskDha75+SA
kDZy+FPA1u2EwWiza0QLec+SaWSrz6G3ZrA7B/9q7QN3yy7lhIXAxBwcpcE1fek2DQ6Rtdm1hmPJ
YBDrcwmK4hdZcGpqllH3MQJsisSlFzSEUCWDvB4tiU4VcD98YSv/k5Cr9G6MPj+/uBTXO/ug5XzQ
JnlPKioOj7viemAedcskL1pPgyv98Z04e1p5B0+jhqZdyYtduvQnIeKXNDVB07T1jn85rs9vs2Dl
VfHUcEgRZJpJYCr2NkRRkGw3DnTxs2NHksO27L2+3Mx+O8fSr+ZVlcLS6OkiZBYBnErfn5CX0tXA
P75i0uPSA63q8ek82ZUDSgdgJVuhSQ82y2fhaJc7aJx6+/q+55DqBSRBDtMkfMzHsvl3lnjHHSZT
K/M7o+AJuXOqbIk/PiWW8hJrUGaIJ7c5EewyC7VHSDj0p93SbdAiQYTDbBXiBdHQu5p7fdflVKKB
Oe3qtviuoRZD26zMzQwCBcsvYuxqF90a/A9GqdBho4LxkrnwuRp1ujBNEHDUjOG05iroOekjcUlC
Rq6UZhepwKDWxczRKjMzZ22TdE7a4ap9dSuRnAM/vq4IYpg/y7tCHY0K/oj6I1ZtmU1cHPP8l4ti
tIOY7F9M1UlqS6Q+AA4hk3dVfTs1dIyYF+oeQ7Jdh4X6m0Y358eZiRQOQjq3FCaTequgFAX/qIX3
3aiqzlmB7XxRVlIteVODfLOvPZvZXN5EZzJKEHN8jyOxhBPAlChdW+s1379EEsA4ZNSXBsVpYuQu
Rb/jm5DMG9kx1MpHsnB5EO2jYYLW/SfcLM6ndvOSslZ+svTgyk/VYClVYi4R+CMadxCQIocFuODn
Pm4fSSsbluSJZeMiEIm4Kvfbp9inchJwXDmUgN2G4X4x6k0gEDSpXSNfuRGcEQULoP1kMJN8/7pU
PgG2kp4706/itRExcFqfdv4o1Zn7QQkmLee4cGsVsAOFQVUjUKee5rKTPVf8wN+ZoJtm/BqCmqU6
g7eAb4l9pLRBWYGg8rgZBZ/4mCWKN6ACMYvrnCR+IGwLMk2jdWmOAyOvRagNHXP4aory1w7scref
B/RTJZc6QyKDpx9sVxF/fqp51RfF+/CHLYXym9c9H3nRfDh9izkILLIykUbP10PvWZVb6v9w0w7n
+nrsK4Glei04PZVI0TEdLHEXXIvDz6lLTymls+GmBcN0HE8m/L54twwfy0OhPs5EY94KFRKmXL2V
VfzYbIX9s0VTRJLIo1g2QeaCIIapQd7YGTfJ8DhlwiqN1u1pDr3UAH9VIT1mNtxkUbGfAdAymM4z
OYa/REAGWvx6C14DWTVAufhMgiLwTsHIn2oF8Pjkce360hN//tp5MOPRskIpTFDfp35lMVCjEh18
/lAE0Xh0RmfX44/M26OWiYf24tjzq9eD+poMf7SZ6zVzVUn5lxCMEIXCMLCxsHIxNml6T44RQypF
FOHe8n5bfttE0G5JRqqe614gNMwFjjtuDJOnWnmwv13eUrCUs896ZumSIJm7Vw3Li6nFkb3uH3fU
pSrSvFYigQDlV/fZ3JFrjaKqLU8FSlDq0v8XsoXRCWMVqIy1XGHo1acbrHCCwRXn7gdatf/+yQd+
BKSRDaRul0v0WBpCqS5I79HT3kxX/4HYY8P2YbfaFNfFZikafrJKz2cff5Q/J+8TMjsnV9OJWYQJ
quRNohXMQ+Q8dHKTgMMngKE5fL3f2AUoRpUneb56hbuVjw6GLCYmhwEzlTPnlgsFdQ2mwzFfdTBs
TR2O44+O/Y8POqRCUWHcRHm2anTrlI7mg//g+tSgVACUKjvYtghpXid8bBZB0uMx1wPTcvWcnVF3
XIRXDy1lhK/vWEKhokt6Wr67qTqWH7iV6g3GpqwQBS5TrDCReHAkXBDBPI8K/9mFKN9PHEtCFr05
wd5nsXxjk/umQfUf8FTZgdRez42PWNxQyf1PqGn8dV9ZwDg83g8A2MJlPP1GoatvrjKq+he9VXhX
3enuIuGRf+iuNf2UmYcdfhexOOy2/LFNK9NBxVdFoWGzVwFN1bweB+gEMZDVrv629uA0cwXYlH08
h3THF9fUNW4hxBFRINrdpPf6ZFKqC+ZIxL6fSbZJjHrDwNkNif9gAQWq01GBC4kUPwc3KPGvzxHr
C8JBTM3hCxqs0lm5C+LVN3cbNfR8FAe46iEJirMe9JfbL2QiAtxoS0C75MClEOPs6j1PLK79aRxg
WiefBJDRlC6HqwA49rDcOzOywwiT0FPWy4EXqvObGcVtkUgRiJq2WXUdy/GzDb6oz5ckDL4nRrA2
KFXfpWiZhgMgaygExhS4Pv+9DiSRTCjdHFHNu3evmyqrssUDtY58PYlIP6a9Cb5xBPbEF84nhvmM
uOCwtQDLHfeYDaytHHyXauA5iu8qjphasPJ9kqHnE7E+c7J9V9Ulhh4GmcLQ1OLCb/tIayU4bUg2
bWzKYR41zDunhBi98Qdhz/ndnYVFv+beHtNN+qrFSoEKGX4TDh4chDj7xMBGkMygYYxjKUge+11Q
ZZVRdte/5r1Iw9ryEADcOy2qM/FeJUf3ANrbN6kBAaa0HRbNraqWNOwAyVir3njiHOQW7CmvLv8m
M1XPkGorfdloxkX7wUj0d/k/yi/32W7wSGTkWoueQN3mu3wM8LWheITqICUn3ocEBps8cOTJAsFT
7VPFofb3aq3GeHZWEpXh2sIv2KKEYF0Ye19XohH6VLq7JzoVf8DrAhO8m2OX2Sb1qeWn9rOaBe43
RVmERuWi70ogF4L7yWwbI06/x9Y2idA98Wls2tgIPSwez1ar5NUqLZa53BnHU1P8Hh7de0J2wbnl
T1l27WxS4Se+EUBXWfyXPCc5IIDXi04hwG68DFvhXjFvLHta3LtbESf02CN7rvGRSxN7ET9An1N2
iCCWjibbyYvTMUZ4Mkn86+eq2/b9UIhOoFvWPd83Aq5w8cjgexxetaqyGnMyGTJYBTwOd4FNvzDa
FkiItaWMbmZQnxDeRryfnE0thCRPwfvHHtAPip0TMIEFoBXKWSnojzrsNhx1ckYTemOBI4Bzp0rr
s/IgEGn5pL2iw11ILAZCdc8hiAazXRlsXT+UcWDET0L7ouDNa+pnkfnygG9pvwad8dTrziKT6CYV
zU1zaPO8eAWOmq/b+LioIORogtk3u/MUvOp8eJ4ac5LHdMfI9zl0O7IUkifs2BG3L3TxDGyHDCJR
WCdBNnt23kzphzQHnBZMJO/m958H7fKkzs5hiDqpX4MV1zaSadwoRwPRuC/ih9h9TjN3wyoUAigy
qhYBCjv0w1Dpey1EfCXeIp2AeV8ytI7AVztTeuNQoVJuvmMC9/3QS2k/CRda+mZeKNwf0ZmZn9G6
7eNoqsw1J836SugaISLf6RCq2/BWZSSWOPx7GiN68K+ckZIija9MHAF9c9wX/3yZlfaS5jgNNbz1
oVsX2SLL9l7vYlF//4ZUnq2Ioi1slmp3w5OqT7NCn5syuKzGOnvuYmO1ozGB0oZzNPsMAzXrgM1B
rApGTZZ2N0iTs6DKOa+NMpiI9mRMG2VbLtme4iRd+GPJuD5RHYiHsGzM58JLRnKP1z1HD1Byq9Z4
d41DVnpXYwAWMtjqoK/0vbLO46HSZoMFNC32C4Px44LrI9C5APk6Bg++teWnLHGkqfUQR+9eDPFD
E0t2JnB7oJe1uokylsoJxQgRdEP+0NVjV2oCsjHhnlzBxoDUHDKJ7kgXISI3SVPkRLzITNef2ig9
e1/Ke6/JSzGD/URLJR4xytt6iVOLGyq7z5L2XEJEzZ53vrmwomSexZ1647jLlkibqtgtnXRfT7SG
d+qcIiBkMjlseHyPoCNyI2YjlNrE4QqaQVf9j38Yw8Ynlby8i9WqfJ+VCE++jib0VPtBMthKOHwn
GGfAFdecutbVDZW/k7b0w2NyG9Dg3Xxdzxqo+ezutmkbHzb/bc3yOK+iyBp8u1OClVYFg8baCcxd
b7g9SfvgxFy9CE5lLpnaoCkaz2by77dkall3VjBIfdNsaCZBiY35Lhpn+Q4hJ+bQoRfJUPxzJIUd
AHjMlRQbjdnM6Z3O+G+idPvxM0jD9D5q+pODGmE71VL6ZV+HrOMd/DIOS3eucowM6xdnkxqUkkKn
Rfoy+6O/tCNNhJJ2CQp6bS78TgbBBIXJUeEM25fmE6jk1wXGFhHp8xZiv/oxXUeP7mbvVVurxcbQ
0LX56wcargtCUnaKszf90xb0SIlNcLOEBNjrtEVPguHZR4K3xq7gg33l5948rxkelEF6VcKTMZ81
pQPCVP5XLrIMj2mduBbzBMQC2jzQoY+ZLPe1ZmCMI+386jRCH0vwVjjkeOQdCsbG0L+ZMrmCik/p
z9aJlAoGsjhIVCYd77QHZHRb8CkCD1WXjmY+YQNUImUFDS9ONFU8d8FzOTIKRgUStoFuZX8VymGu
WcpgzTXcLoxK+C8LC/DfzsnL1jk6eCJBcgjz4ye2Kwk0N0XVeDe/RN6gI1zULhI+bGQdTNRCA4xz
yzLCcS2CihegLeLNQH/IFYATuKDiI2MkqJHhE8GmaOGZIMK3LNh6P0QBmiMWJpuN2YseEVRQ1OZ9
HoLdPPnP7enL7lay+ul6G3x/grQzGkG8w7Nt9jdkxtAO2QAHwPxOhseLvC5j1FAMiIQ8ChgtwJho
Ob3fvbr1orBNngp1Mc6t2Xa81c4KoOjm7buaeEeqGGrr5VQG6RPuF0qU5iBAvG5dIIfIz7LvM2vA
zy2uxJ/bO4pB9pTDcs2SBMpGbT1aNCvYPACkKQZI+u0BWbVDtPXIMQJ/s8CXgLC0iKN2VP+Takkw
atqPuh6szN8iYcosASUo+pUY6ZxczDhgvOEEAvshWQd/0Wk22a1Ex2wAsnBwyRqjxDAhFCgHz47A
3Tfu+h9enVWiAo+9xBYHdEw1/wd8Eql7i+vGD8dLSMT0ySW1n6vb0Gp95T004JvG/cuVRqGuw3hs
gALnnmjNw1DhZ/D0BkpAaVrS8qdRwc0FNCUpSZh5LbT33/tUWcXfa1gmdycqHzRYdDrk5hCC6rNV
gpVSfwQxBpbqUivxP1+VAupA+W5bQqOL4e8exuQs1t9XP3yZAumFfwngCzmYsYeSiKBiTa95Hwsj
/Bz0ZzUe6HogFGaTRHbj9zka/66OXPMXwivLsI2HgiIMDrTwV8G4NGingXMFsPElMAxKBC/9DB2Y
Yx5TBX7dWZLNTuskkuLqboSXAcxIfB9hWP9Zt+NGD9d/N+ofyO94+yuItW2DNpU5GTUYgvTkzi4a
k1GCd2AsQ5BJJ/rfEtvMcBKE9KI15Y2lUhiwHJGR+ME1CE6Ys510/DiUYyHx2gUqy8FovHFQq4TC
o4fjVOyUZO6ZCeSA3mTpHklTGLqvfqBlj7/z0n3yJeMYzsY/61m7YWlESpQ5lP0XBch29JM1FjZP
IlK8MCK4aPHsOj+LGPV8LLKK8thXRu1rVsZlnaaBIciipjMay0z9O4TaDAQXHn1zaUiU8zABbi8U
2e/E1haKeg5C9Ei+WdAE3OlNRs9T3UvxEYkfzCfLMkBPJyl4flsigKPHD1kkyCywI4H5ZRojGunI
eh5YM+GJJrOHASEMJ70xNWCcrGMOeR+EWsIGB7ERwpHEXd1lMnT9EbW2X4eF5lPveVOxKSpI7xtv
KNs1WnmG+9gTJ1INXH6OKTgLsrsQVnljmEcTTFdDsNonQcosKl/gKuJ7TB4o3IZGKPscYqZ8HsIA
KMqhMzEfeWgd7VOJYNS22l+Nk8ILXCV4374O0b8yoQd9+atXRf+4jNOZigeeM3GLj0djS6aTZkFF
wucAtnc4Wpf0OUQljnSxWX/4uS/O6bJUOjD0ZmSJ3ELjsyNAXO0UGpUU9Kt/8wh31kDWH/sy127Z
aF2CD2feml9qKE+7IY34/W57ks2DecfkGfsXre4hIGaH2w4FMUT5ohFKzVt1yuuKVrYHpblP4UGb
bEzHiv7/e5Br9VioAAhZiH54/G0G+7mr8aE8NPyyGHPfbab15WswaN4Vl407L+ErxTY5hFsSnHbD
G72gqar/HbrrOwfKR+EWZfeWvq8ydivtlZTRerb38/4lKQ9IOooYkf9sI8zmclvPwx5KabJXvfOc
Kv6lhntpBAJPn0AwYzlwO79Zej7X6SU+ayRRJJo5ZRGDsfwxVal+GBpirBwvCNnZY8gFw7FGRfCm
IwN/09ODiXx+uT8T7T5w1Vfa/JlGNXo3wKL0PVIxDSHe5o0W0gSCE/CGtU2tv52n/QRFRfAS3UES
oIij1wYFCtjDyZ4dZZyiqvvgsBGxXBRHt5vH4nWa+puFV2UtjhGN1/CCPYZWzNrmurQr56DLnNyK
KxC+xhGUGflI6M/UGA9CSWkHFZUJmVYMY8uSUmG6FIN0aXMe4Xh2xPWCCRohosbLaS020QmPFbnn
std5Xii6ZRPiuLN+WNKY0LRJKfyx4QVJAesi6I+NIozhqeBop+EGphqjAC2UceLXo62xbvoKVaMw
tl2dfp89jfz6iddJ0R/VO8lxX6Kj/CYTuiF3DEkB6JhmO8uv0yr0r3SDhX4nHXe5apobFJrM0JO8
Caboa33p9MYXR7yS8b2z26x0pJjwxIuEP67RmqzF5QP0fLV3Kb0RyRgh00Wp2DPYcCIBN/s5tVLB
eCmkY2l9K68TRMx972uTFgxDzsE3V5AFNnMMejIus5mnTxkLVL3/daLVLdWi964KmNZlWC3Rr71r
jT5Ol/GVLe+MdBNF7Jh7aaxoC7xGDR7fzBOPkZcY6V1xL/KZ3KpYz1kBu7bsP9mkHczOsPITnqBr
+asm2bi2aYjGhpouagc/Os3RJMl2n5to6Z/glidOYy6Gynr32ip41lycxBAZ6HnzUo/vp63NepM4
4sN04JI5Vvirm5NSCBE6dtGtQFBza862cP//4Q31Pw1wJyhCk6MPnG7N/ntVmVQFMZIKPPi1dF0x
NCgTkNTXfisrW+OVRF/SNzRT6gFEypCOlwVVvoWY5rAiomtqDc/miVDWKg4axNjL51X68L68ALqs
YhWeeoR0bEEV5wgv7ky/cTUU/LbJAP10qJLbp6DWuLKK6dXMlOfmYpDohX87ERfrFfJwsElO9Dz+
enAwDpm8FQ6rRJ0ND0AwAK+BP2VngrUfyt/ONbf9SaS37o2/juIPyw9Dzjrlja8nReJQDO2AQyPP
0twgJZUffonmA2NzExWsvTpzv+UKFvhK+Tyl0wey3t1kfRIvUBu90zYnMwMTlvldy5ED4v9r1wy2
2cpw3bsKRuKtn/jK1ZRz/YUMGbfs4ah7TiLqe8H63huUWxUVPREF/ZN3/qua3R9CejDTD1AjuqmA
XQrOuKkgyLOPjDCidTL/vfgey+f+UREEOpKE9dnfO19vpHwRaC0PCySFseQ5wWb3KnlTuwxQOGY1
nbYvFF3bxj4fEgBmm8xTlftIiblMesuoHihGSpT1/1P5TOkdolybdQYpO4NYTcsGkCkLzb3R/p7g
zYFaaoSi9nHK6R2lV25T4D9x2fiAYHPA13iNc9bPrqIPXAsOjRt0XrnpcaWp2m8Yu1rRNykmhybN
f70r6f1gxeeeDqZpHU5H3lVtA4wSriZl34GipglJy+KvfoFBg0bYTU0Sd744qUYushqk9R1i68N2
p4hlXr5vM6K4DPa1vCaQfFsRWR/6xGNBoVdb+OxI5tWAtUbMfoP1r7GLyh5MJ9fLonL10Hxvfbe8
IxH13RJ2C1Foh4NQVo27Va4n86pUErO7vARQjbfR374xG9KDoKZ+hXYiBFf/TiadLWOMHoY1eol8
pPdGu79ZJnPt+oODs67K/R9WPzeNFq/R7h2g3kCAghQsRCLM/Vl1TE/UqQ4+6TeyAYFSx9HYYk0V
nHMdgmy0cJILnhkQ+SkueF/kheFyKqMqDspI/4aJSekuCz/GPaPdssA9uAUhVo6TcU8svHxlS55S
v5V5S/YrYUl0zjCT/bkCxxoC6Ym5pR2r4t0TCaT1cqC/P41LtyiAK932OJonZcaHZMONEY0mTBnA
wbIUShMIwfN65AXV0S1NSFjkfJOiAPogL486WK8KfopNJmiCRx5K6k2ek9et5WCzOt9f7czpI9rI
Sol3tsohqRYHrWqFM2vzuq5vbKDXkMlL5Yr2/4gA416dKQ+fw4KqSd5iCYF2VDKBovIrZTFqT+vW
VJ1PC5QxW3+Psz+9CZEfKJYdooKnpnnBQnGCgxgC7cdUW1xOF3QnN7EkU7SKXnT+syjNYSJS3r+b
xoBqx+UzzqI6jLiahYM7idjAZ0+93dljWqbD+j8G50cDoWpPB+RN3Xx/T40j0c7EIsjXT7q9E2NC
AvJkte6dnP5lKOLyYlPNI2HIwJeagbDGeBieCMDkK4QgKZHPJtI/ZBFuKKL7xWORuO7CP31WOBKs
kBEfTM7KAVDVoxk9t2Gxc4/D1mcDHoLSjXI4tJZXb3U4reQcXQmcLONjriYsu++zrr3rACYoyXUa
GUfVCIL5vUq9kFjGP7IG55qMM9VDLkayXN9OZfsrTrUMvtKZAQtzIp4mdVYhk7if+nBacRZ8+h69
gvYFWl5mgtjeBdTiti0KebZBgKTF7MHud0BEWT32FZYvVRTMFnU2PUTrEev5uki6BvwXzOrxzT0y
PLj8YjMtL0oi9+u2yvFPfzI+BpDqNqpdWqKKPv0UCLeNpnRNFsLjP16Ohdc0ltotvk8l/Yh/BOfj
kLpjEqrt0gQ8fWbl+ChQWyWoh0G8KEvJw/zaQ1QSWR+ZRXDZsHh4YbBfHBLHc+JE2cvuuzrtpe3h
aUr7TsoyjAqPXR8bLSCoE4MGpJwOrk+VNppptSN4ndWTzOpE549gV2syqvkxgpC89gE5QGjbJLjY
o20m6B2njy+PwCG9zWUANnOMd2H8iAnYOwKVRqX1nafL2zCUiNy88WCX7h0KfLQ9uIkHdCBZX3nk
YylS5WWK+AzHRMvxAD/k7nEjIydFkaMpYhPSpw+dd1TPIzgwdr+/vhctugNB8cRbIT2oZZz7HdAS
HXykdK45OptNYJHo0cTn6M+1LeziA+t5sJi2sDEoKE80FsHySAFdq7HcJmKonyD2AgYU/O9reyQ7
we13vj3H+QsbSaL8lQ9hQkKILWee94Wfs9R8tCJcLhtVyZkXsJ9voS7BscwcQA2LdU66ZsKw3jdG
Bcx7fXa1kGlcU/q2OkZJ3Kd0gsCyQRmCmXxI2/CAHzepegnCe8SHnoSvuOwqqbPc2M2wUeASHlY5
UPlhSU94TmSUWqSjbF116aTjqN4Zcy51Uxp0J4cIlOF7WbRV/zaG/TVgtUD0p2O0i+y7S5H+dFnZ
m89RLPa2BJIrxoU5aCPDI2cZaLhZDF8/xojjK6YEP3Cyj99kSkBXxCFlQGl95+8ivAQ10183DjpQ
Si8GlHtM/ZAKt1qhSopfBgbepHzBq4pCkWtSALuIeBYI/tlSWoGoTiQeYh8QykocHQQmW0rHvYDs
o8E+giH8qqB7K0Z81LJHDfzTa6W3FxrOXs1bGBX3MNrIgNc/yzHUtbVD1myhCiOlHA33/+5uLk7k
4OWoq1MxViK24voySUrYM0i9YI/qXBxj326tO0LBSutS3ubpJCKb73QqcDr5CfQH2FxvOxyU5Fqx
t+CS9rtAB2jn+dSO7Ae3j5/KovNAfUFWDf9saJImuwRDA44WJKJIwLtm7Jc7Ce0uICYPeZUpBWQh
4bAZxBlrwrz1CEENXmfwchRgUQ55Fj/O1q6iK9//V0sMlW3Kzf5H6xInsAxg42sks3Y0BPQI1ofC
RRfwbgiVlqF/mFoxbxX2leGG6BepXIwEvUJVERcFVHz0XvFj/yG0cfcSlQL/uC/q+QgPnTGt/gez
jtjc8aXzy/Dewa34oTCtFPoKOlfQ8mwE8udTnvB+5JJCd3RoKZs0o5LGniQa8eesleiCyZKxyzvU
QGgReaw1I9hFXpUiqgL34IHoxjxcNQhbOaVSwNCNMiGyDtdM6mweKuGB177w3Kzpl9jqRv7g2H0s
wCqckLn4Dnbh08Xo2lgRAyyKQG0tw2K+/JhCv6wjX9OR/jr85Le+Hurri+i6IXcpsMUIHZVwKrCy
c0luqQS0+XxKMxPbfiKcjRZsSS9M8Vg0fzQSfTykVeiANcubnZGeqNfiDsCk4CYvxmeYVj0yl+V+
yyh90/flbKi6i5IsQDZMp2EY2MpbNklEY6gBzKXUzHt3R1trY6jIkswfggrPhNyPL1nNs0c8/cSx
AxT1etlFdUfdu8mZgjCVFZtX3lK86lsJMmWmAzJY4p98h1+cLDYtrOySToJZ2clMWJc2e35C6jQQ
nvPcO5S1+t1JaR+pkbPX1LLT9jrqpUBkcmDGz3OqfcyCmGNQwXwPxHz+n52GAqtnWMcYDiFC/oUk
RNsdvycJKVVcFVDB1jUoufCMH92JjvbXdUfwHfXALgk15MLK+7wVB+XzSC9fF1xx9T2nHSJ+20Rm
V8v1PY2xLNvJ6WPDE6H37vJvtP/rjiehyQkuWN5cZRsb1brIwBvAuQ5dZ9rw/ax9jxtSWqXWuNfr
PFL20VYTF/AHYmxTrUpBeXknRiKBiHZDL8cUO4QQ43KrzYxIo1HJ+lly5VDisdD68K9wwP7NL0ZM
UInFkWVQLWX1TIDyDDtN60eB1hUhFXg7X0ZLMf1rxH8vde36hdVqpKV+nPe/coLWvcElH4Q64XZa
i31QKJvFNDLUJSJ4+JZBziTM7PXK8M0yZGJT/xkEw6Wcrtu8W53mmo0plDFgrKzju5E6FQQoyPXz
3DxSPaJLyKyU1JsCgZ10oqFvHiCMKfXSlr9JUB9PFP5QvhSy4e2N44JfaTbfSQuqexI83bPTOe/B
boMprz70gQsY5sLOvfGWsvIYoeLxBqzuqHbUTjQ5UcZ7/UtUvzwQ4s22Wng5D7UO66tciEH7O7Zx
4o9MKHVKZWvnFKmoorpD/Vh9ABU9tqNggv68OeCUGoYUMEdBaSbQ5ZZ+pRh/sHO11SsDS8B5lJBY
Ejz0/yy2bi1AhKIM+SgJs/86FfJtQH/+YiuDSFrTe7mI9QoClJqLhxCz3Up+0fYJK5ZGyt9vpGbT
1ijzl8g3XBahc5x4brdDW50ZsZCusyq19qLZmtBxLVgwYof4H1XWud5c7ww28n4UaQYGo6bUiPok
0WGxnPMRxOCJs+W4dkVVVguurrEd5BoqMo58etBQsLA5nndlSdMgLE3rEobY2xmyHQU0HASpwx9G
2+bYgxChPCaKjDVkzf/8P+furEh3gybvsppuUyqC4/mxZcUmlleps6r4aFuOLVqm95pv1ORO1VhK
LNG792iAYC1GewJK/Kip25UF4KttswXY/F+N+almGxcuP6D7eg3pTpAKBG4tzxTvL0fWl+QRrO7V
ttSzL6bda3vGhygHwLR7JLpibDZ4yVM9I0pNyy1TrktVJ3ryJNsUSfxH2oc3B+AtoztwEMtueurt
1RpNJafMgq3WmtU48AhQqnZ/8opPfdDfrCMrELAzu90SzqzaSnBu5IGAtr6N6xN0ocC322Kjr4cT
wLIXDWBfWe3UypZ2pSnzZrkxTawQrJrU8cLBERb9KVyHMwkMAM2TcGxV+ouf6LdOulcyzyEJb0jE
N574VgdWLZ9QqH1N3p0vlAzZu3kHkckm51dO/2nkMHlzTpFSy1lvfauQEWY9NcRO2Rml7pxnWD+L
0frMFrQ/c9UpTJFuaniyFO0Shc1oOJOcPQ+wOtOlW4iOVcC7ia/NytNXhyKTeDqmwDZlYQiJV9+q
FOeO0dQlRZSvUO+0DewCUrT9bRrkq8BNZbmElf0aYzti1aOuCj2s85iQCS6a0rutuz3TJoa9tdhb
TOYmK0p1fmWKPoNxqcNoLjjibyOgo/cbqYTKb48xha1tr3JLJJx2UArkOsJPPXJ+JFb53B6W52di
MC17iYdYJOzPlQYycNpZ3QiBUwVK96gVw7Q7Pw/6ySb45oZAySS7+n0iwCfo7Zqs+AmM99m+P9t/
4K6h+Ud0QfE3QkLytLHz/P8c3bgUSSQZOTKZZ5rAdcwgbXfwjIQyYjFsFWBb5keq5wZyPmRnHzzZ
POCaKIr4d2z6YQ0sEAvRyBh3MrK9BrnlV0CpkAY2ZY2ICSjmIf2QFSsncg0N2HKC7sK/UirftQxo
HRGfalxh0mNi/WYNyw/EurTkLspnmwqW9bVEPrURWpO0SMDmysXZWS6W8indDmEumcAgi9w5R5uk
7WyEQWi38Q344aGf3cZ7vHmkhXI6gxihMc1Wmqc6G8cOdUdC1rY7TkRY2BsDVrMQniqHt56maa4e
mGTim6i+T0F9qPhLq3gFEGszATYmWkA22Y5ccQ6gfX6h1ef+XCuKXuPrmRM6ymSUkla8nBuxwLhc
eg3FNJFMKZ5mMsbqKI4+B9tXn7YED7hjL7P7Z/c3NiCFzZH4y6gjOn7LkqULub4kj3GAITkJtCgc
aVBZqSAdBZoJNsQocoTG7l+8SgQmkQTwsSRz6kd5RK65wdggnUQKoNspbyIsZb3pGqnsogyWjvjW
ZwQfLcIkBC/+QKdRkMuC4TQIsl99RMgpLFNVFz/x1RHLsEKpwuJ+HuHqDpGfGaCgBP24BzoCWwTi
3cY4Y0mY58WGY7LXZ7Zng1vM8yFqLov2F8Ki95SaanJ0klK+sYhJapnS9MNpJb/PjUmVg/p+qZM4
qTmIZbxZe/t7Lg7rtBbhxHXIWaHEXr8theM2NDD1Bn4mEz9wubyxfxSnUJ0B8u/0F+q3ZnXSNSvu
rtR5LJ2WU8X1fSqfKqHwyt/wLNHESQ0s7/eLNnoXQa5tM0nylATgkZTRxtlNDTSKiRXwCCLw+3g1
6fpblQOBHgyaGgNST45xBcujNhBE/6QLjXOwZmSLdDs4LaA9twDUInZG+TNk8tBRLjVrAFOoEVG1
ZOcuuOsx4k61qPnrY9G23SDKPmrydP0++X4W6Bws3ITWaW7hXhyATYalhPVi3v7VFQl+ihEsiCtP
5zyVMVFmDS3199xOGWm9p5hYEMuRBmHcguBc0X5kT4xKy7OSR6TLlhY8fhXHpQ9nV0q8La1ruX6z
3cIGP/vAGKWwZ1VuWtcNJkEF1vo7pUa9rlRZL095wJYhZnsTfWaJ+gr3JJNxv+53raI9x7oOhhW4
e9v7RU5wZ59J5IeA/8JB8vGOCjOZLl7F30mGIhghLQPxDqC4JbXmYtkQ84YmqezjAerSwHdAQzNI
QeNbCYCu7XBkJEIKmpCn1hjnkZClTB81QHHV71dqOdSGCo9WitAj0pp0dS9yg2qa9paOdCpoz13L
miGpJQYDZd1SFyo8/wHWpdfI4WjTzx2sy5c1wQkG3O3ER+1k56nhr/OzOQxnF/EnmXuyKfc8mVLU
bnxfaqNuLdvfA1wB/lHgHgVyQvAd+k/5aS1V4pY0czoIHZ4PxF5m1WcW1eK1lS7YBO8apKNHFMJe
ImcF6qjgpBzTmAkTx4mpfgwGkLrNbBg69tQC+jQNwsWmBvHHP/Xbg+1NotKgbFBXeAPAewAK4yIC
VWdNROe0JOugBQ3oUjWCcq6K04brOIMhIYPnDBA3AdIVNW671xQBrigY4hQRXKlDiMsMljNsHzEE
vi68LHg4/mxeeFxueTOSkdaP5Oe59dPrr9UEEJiSzkv62Azjcsrx9n7c5sdzKrpsLqxPNfKKCPfR
BQcricB2EkKnYuD9N8/UJYTISe/Muwat/+3GBr2XEd5ALVj8eieSgol1BBd1piwLApfyBOcttr6S
VtCQ6iCCczpxfyKADyfKRMLiuVzo1loA9tSbSHOMjvMQNL4tAZQUE3DWfkRIbIYJKBxsgVCGW2Ig
ijBo4Lig+n9L3YgeHyF46lHzor+YbyE9f1vRyqnoEKXVf/D2EoUzdAy0/mSIPHq4zo6K9sjDFwm/
gDxq74J2Y3VDNZID5sNp1oKF86y2KkQ3Eg00PGHVLKkJvxLOZTkb96ExyaHu74fPrdlnro+PcF0z
Sfi3GEozjNsEfOiu2+KhyzROE9JqLKFrM/G/lnEWztXk6Pkd2LkJyrnkgeGL+dRDeQridBEIss/D
1OWKKzZfpM6L7s2OCEoPOStjoywjWawf+cSbSc42czwsUBBRZDgPJoLVyQfs/YjHtfBtoLESpBKy
9pGm6BoxSnxF7bfY/qzZemhSIywrL5q/JAk97KxVNQ2aiT84OVqG3Gg25rflR9OaBKvhk8UWqPLM
vmxOJCIFvfD5BwvXTghPAcVcuwsfAB301ZldxfxJOQnMEyJdfbu/uy/9eGmUbVVhzIvghD9+8YUa
dTLnkFtDmq2P9FDIVdRiaG1eRcdsiU/XP8r1rEf1YTG3Y1pkhhXlVMkiPs/oB78cy2FtbV4YSNaM
gAmgauCeFXISuHz7C9o8DFsyyAaY71rUmXtVIfFT3ylHKSgQS8ID4v+rm8OJzD6TUw8wKSo1QX1M
ssktxkMCTWMaiy810sAU/cBH51QJwCxPUU1HBn/eOT2YWCznT31ne4uLZgy1aV+AyE+ETPycZVTa
QCR+TnkgNMA9qE2AaOSS46NiKqOaFOMuYQFy2/joUxHc8SP6aVTSoEt4Y388jn1sSnJF1lFaLkfe
ws6933dEz34G3h5QHsf4GFhC4ikM1wtVdJCCpbHv0h9T5IxiGhy0X4hHuUVD1TaIDYPQO25eeAVP
W9bPylchmGxEF26NUal7uel5+NR+/6Rh2r08vo9XmXq06RtzVvBKh8if2huhae3gU9L1DaMHr5lV
uQxM0VrEa9bSovf0DeyMLPriIwIxCpqQmmpouAzjl5hxtYNetf/DuBnaIvHc69YCeJ8JROEwPAmf
OR/COYi2Qu1oBb4V5tYUvdDiIO6cLzku87JRKDpjaAaPbceSIr3oMi49cw0mTE/I0Tnz0uZDwVkm
5RqLH3gAwknvHquw65/iJh80+Dg5554nddZGEuhlPKKxu7atc5kEo1ao+qW2TbKzgFGlvtNnVQ6e
ieK/4QNW5aK8TYqYiKW4YbRhv8HorHoDwkNgwtOo4bTH0TBSgDM2GvisLVK5Gm3oTzMBwo5nABzb
p6bLPx6us9isGqcVF8tJas4bWUL+M6eTNr1PERL9y9ye5FqAbDpMJC6u1GonUBVtRnkfOJGBD+x8
9kO4X2p+naJ55/I0i67Dqh6c4aE9Su7Csx8RlNwFqQcdPpx5jmDrWd5rGpKBJJ/PVSIQtg0faImr
jvN1ghxcztuPprlDr+bMAoA0TxeyyVpnzYeWan74cNRwm0uUfqbztBu9Gny2tcPOJLZPlxjE2a13
cgYs5svbjunVucxGN6ZjdcT+FlxBTVvqkM9An/IH0a4kk9IraoSl7YD6CmA43ii0BN856ugV1WWM
rGCbPmMCF86VrH2wIKukWQil5adLSaHagjyDRJjxxbbMbTpH3bojzGjfILM8+JlCx0CkpXa0LyhP
2kSCUxkz0znenrxF/iKfHPCdHbC7m5yLpoT6SV8M6e2/8faz2cnXAU2rshkX5VQpakn9A3FS9/5y
J3qsuBa/8x1ug3PoCG1kV7y8CaGio29Qk39UR6nPDZLvcOgDuSskACF894DVholDQPUhqxUJQ4wV
Fd9N2On7K4nWJvOlqJDYNFy75wHxiI456SOM90o2QYmZud3jYRElraicf1vQ+k2DMyCGvxwosW3g
2Sj6Eg0j81VM8EBrLaS7EDgKWpAMQsBv8V06aGqYlG3iNPXzEM3kab9qw18Xn6Ar1YlxKDscjO5i
kaNNEy9DF5v5uSxV0fN82QlvnGKvDGQw9Lq2hRuZq9gqWtr38K7hDW65yoBAnLxswZE781DrAYVP
fTx7v0bsNTeipDUnLFlerkWsOp7RejP0YO0U9vzsECqEAcdZf9Edpw8MJxHm0SSCQIiw6I75sU7u
fr1IWK1k9SRkgLf8YbIC7OH+x0fC4yT59YvRR0QrUSIzVbiSscHvbq30iW6emc741LaaNhFT9Gdp
Ag3vESZd/lO/Tg39BymUjwezt4dYkbPkzWl1q2x+HSozwWerj7KHrp/ZMPfTRm8JyuYuTKZiHCHy
LVH+secY2r/xkvK/gX7+hczYxy/1MQnEcH+8RAYy8ftiQaHi5v3RHKOYRP1H/zZwmwGMJD88ckGH
BroeiLEQuBs+nCoVISHLcSXy+YvkalDECLGTOiDPO9CeL0xiJBZez37T9tsQRke55k61tZ5wTIp/
PAT+mZAHGQaEk5A8QjIgYbeYJnarivnqP3zLkJ/ci82P61eFubzD9OPSPUf9JyB+tjPbF6xPEhTa
vHeGYFhpatWCjkSrseRRkJLIFT4hCRaboyFMOjvOdVbnsIDc1K1B9/rOKBY/oqyWDE5ol8l7/ymj
nfSDUDuT7DZyGsjPZNLQPbvVgbwQezSuQCFrBzKYHbw/TtjWUTOR7NZD41c6/VF4vMzEBqfYzA10
7MbseZ0J/4RK1sgI8aMxo6ByxbAnqc/Fo0i0QVNAniAmzoEEyE9MTQy6ztvwZsww9ndeSubQCAHV
856MKVUmDTbT6aPxHQ0ejiKkRacTyByhWBx3o73u0fpfK8xTN0ibxyB3HpWmi3VE2C/mlOCHoIWM
GHy7ljSjay2qKZ6JF1lekg02N/nbddc3FV2geOFsWDH85Wzr5kbNikTENfo5oRL4vbTxzmfd96ZP
IVEIqlshk+KcDRe60u5YTqKccqhbEE8YLSEMTBFZ6KH2Kl0tNL+//xQzlhXQlUlrNcELoWoLrAik
Qr/g6hR+iZEthCTzXoxRIDbJEyLiWLH0KSWGfeUh0JG7kdPhBML6CZU2utxqZ/QDckqj+pJvqMxO
Kv+sIptaYlG8GZKpiYbyEE3bdJTUwObNkrcYHKQW5GVRZuP/NkFiQYzlqKnXpxSZUVf/lchWPga4
eX2shB0xrbc8l9ED0e+oLusm6wjAubcKbCaapmH9GprzO3LH4UaVzVLxWm87+Bczi2ArE1ZhQj1T
anWgAb2SZll5LEQZuq3RnbqOBZG/FNhlBmg1EG11FEXYagPRTWsPCA76DWsLPMMnp4Wk7oaOue9d
lC64BL2Kiq1soKBfGpso0tlZgDNC3cpEE0kbum+gQs1JckbLfHhiI0f8TzpORMpd8c+fHkgEWDRF
935e3XfOSiu4i64aGHswib2jbd+5Aez99gGhnVNfUw0DFVwvca34nLMpkQv9+HB0ybZzbEbkEobe
MgQcQgngWQK+cAe5o97okKs8Qiq7ww8U1ehtULSKlIgtwdqWXghkpBL9bINmTu6S3H4iTfBpr8Qy
8Y9OUen1wPZJTaaA9KwJIlChRnLOY0Nv3XMBJfZQF0hSYi63tANaGZvv7b5JC6H82AdEA7P5CvyS
XxyvmmPJGgvOBC6w84/dvFtwvXNBKl/YmYCL5efyMejgnc3dtX/JNKi4Oq+PUyBdu/lhJkR23vTl
FqwSVcg2gMNomp5DuidaKUXems1AIiqHs+NajOoODbTprdaGxA7w/UTp3H+nIHABAClRjC3GQSbk
9K2MXysBijFcZOcGbgclunMOPLcvY9DERDpX9lmXfczku0hjcYNDMb1aZPx67baTpOyJSGyp59wP
GxE9bAYwFs6LCygrAJAJZq8OvXcTI7viM3HOCU9yZP2+e0AiElhXBCxdG5XaZ0YkcGBqhJ5Lsubo
MQPs31R979iENe/6lf1Johs0BI6kB6I9mwuFDTQeoggzCAr98NyIlk4LVNVpUQ6EtTBBSTWcdtJk
+HPwZoD7X6bTCOD8qTsG4fjnXMN0ntwaAxbB1YX455bAh3XCPjzIfRA4CtVayzyXu+X6MDB3AZtz
Mz0LLAsIs3HQ8ktqtE8pE3OGcytCdbheBo18FM8cOdAfI2svvkBIDbOnws7tR35iopjkwVXe+CpN
jo13aHz8G2QreJ5jeffSdXCUYNUHIp0nv3pRm0sO7mDHDOjrdm/USMnsXIEnu4/a2rsnNo+zP8M/
/iM7INS6Xeo8GsVj8CneOzqNpYJNqOT51Z+jL2d9b8UlHiOJxBLqYl+w4+EtE2iCCBOOmmr/Jjcd
L45zlm34fLNAQhsoh5k+brcx3oIq0gHGLHC6ePu/vrGxY8OtUwDiemBwptEKfWCpLGHry6SuUXC8
YtS86O3kggcThdA4DyVMN8Odqv/6ccmjFutmo99q9uUt2CUZ29RBG6ZL0K0o9V7BcO/8o12ymTth
Yz6nrV0Ipdz+YpIEXEAhjja8wlnjBr02X7vpRaXbnrsrZFZK9EvWYEfMU8z7+TlLMQqy5txQcbKX
oj9fyLetSn5uakqVTRm+xVojgLCEskO7Yo74i6rQi73MZel3m51+9GNv3AEcekGtT134kq402sWp
RvplyWmcH+x2BzynJJDQlldTkaqzErTg0sDeafTwf/ASBRI0wyyp41vu5nCA/8+VHHhbGwclWf9K
ejHNXrl6dx8b1tJ42w1eA57D9j1hP6FQj6ouSeAViTVd+UNv0Rzlp1fq0W+pgSO7AhiQl/n5gGLn
OjbvuDlf0yY4T3khNhOQSXtqBL0jHMxUlAz+P7XtE580Wqo8o2t3rye8VMj3cpMhj5spSiZ+6fJk
Tgra/vTkTmx/q4ZSbd66S2iur+zVvqrEkcjF5FichFffC8a3CCIz7QYlaR0qA3/XIJasZYGgGtr7
tHniE0BkX4+exMnqOiGq4W1cWzrlrUWxWsssG7Qhdu7mOxoBXJTwgwXV6Ro0HSl80AAUYzFebhXa
1YOXvuARybLggMjG4VTGWu0rH6QsHtqmSGJOE+xbPbLJEZdCX8+F9rMCKXGP0lCvnyx6TcGp9vVv
3PJ1FrcpTD6+Ny0YuNsktDFHhR/IM6uIVKnfjZbDpkKFHjTdf1RPLaXqV4ZzWm6Vga0Zmm7d9KQa
CQgTZEDgC4e57letcOrAQAm9EgsYter0ZwNgaMBblmX3r6WcpLNo/9LlDTAdq9NmRTPZeKWGRSHv
I9Kk22wHGek/as4oO2BcN/wmquh5LEZ89e5yBL1EjGvHfCFT3in7yz+LCKboYRekkiwUe9uco/Fg
TWbcY1ZrQJ3vbeZuQNzaRxZRxwR3oTWj7ym4Bk4MNpoxy9WcYU1QZXj5mZhYwBIhSZx+WWPtI29d
n8Ky5/zAaMtjFh10P3JrryCdAX8ipPLkwPNgPeJmZGBNtWbx4scX+yjvxZLzmOrwvRUShs4M468q
Y6GH39+USTLgxo2Q5cJSRfPfAVXTyD6n8JWZWTeVYIw4xxNMvu4GOssHKwRmW9ttQ/uxqlgkJhQr
EZpnkJGHsKA1YSoOqAqJIJiIrWtBIAySjWkYJV6NWKvs6+ijC37CYHCXHcfNkMBagSJIq7UQogNl
DUa9OJjUyR30lEaHRWQVDb9FiZflIVhFS8lPSKVjnnyYpDFNA77s2Q0uJu1BiG28NDPQenY+Von5
st44nYDdZ3cccSWk0YHOJRPFUNQ7k7HX9fucnVvjNIOxqCyQo3hQUhl904REp01KznwzJP9vZxIj
gjImjOPxjdY9SZUQJh82YB/vsPHHrI8Kf4FIR6KqHa8Uu0rH5jdjPXXgDACWGCmd83GAq9IV/zBz
c1cQHjbAZU3PBzkCicdEo6J66DD5OLhzGjIxJWP4OQlPjPgmgcRJL6WEt+QbJNn2Y3yAVM+vgr0z
xKIdMY2mopVXlB63rV/D0ZB87RRd46bm2MzyhTsptcu7jV9ym+gfLvKh8n3IfXvUW8jNlsMUL4qc
fldgJcZYjmaECio2U9o4CTsyoZzBZRejGBadm7sV/CaTsOYD55Go/TjnsImNQd9ysCUSa4mHyPHj
zWt/5GOz66o+belhaLUwE/a4WspHWtshZxELKCKZyYU1ogypvd8yKqyxFnxu1ZpW9peamYKPzKAm
C7HBY3Rb5asoQbvXnRijRN7Cs/zkYqN35qAUv6PxrF/Bq4LlBfiHjlDWklbYyTdt51cdwCBRrt8B
3fwE0q/DHrozH5KIvJeEUq1ZYorzy7xpGJCU70D8SwWu7Zj3RBCHwMsVgcXg3Mfs8oU8/p5p8/PH
ztedihFx85Zp0P9R46CXBXZdnxwEhJjzN5h98Fy6d2ki5Xavg4+jbr7avhJyfEc5qNJbe5+UJX7Q
tH7WtMgEjin1yNAMN5pYI7k+D2sp3lAkYNhwnIz1zDVS9juL+ENs6oRqWRO9b2ZTQkJhPWOy5xEn
wjc7YOrMV0onEkJmu6JoDMcvGpuYFZyTW/6gAlwS0W5pkE7jk4fm/lfZtn6AFvehaA626fu88K2T
uYQ7XDNsKZqbedJFGweoHI4642plk0C2YtyzwojqY6iidPpEoDtqjrXaHLsFiQGmGwlGaxQhQqDQ
gd0wOWYBD7u7XeSUv7Hds0eY3IM2Z6nUrLowfsNKs8KsA4iqh6gqWwQXGG5qlCdHiaaC+UeBi9ki
Xprz97gQCXvbTWLp2FQOQIMZfdy+Efvn2NMlw0Arpni2rQbVGtEusvUNfznwZg/zzRZ9116b3ntI
o5A54meQ7e6nYFFPJQ6wpfnomlqiyuVE5YNoRVt6kZWEvUXWWb3/wyvymcuW4GarmfDMXuZLRZ30
JL5NfFvxMBot8FMoFg5HUlEpDC7bQC80WpwHVj1iY7F2W1KRjSwJJ7TorbB8tp9BGYKIfRnddm1z
IRPRMRpTGGeO1rXh5xzTceWBFzPOGG1/iPUYFC2T69kYYMMFI1FsDOm0M2h/aIj5/Z948XvikEiX
bFKXJHV8fDqaC/ymrmg/AgHg4b7QmEQMExJFRkTKfIWupyiK+QJzjvjFTEBUV6cI6ZaCOA7uMnUt
UL/k5SAXNOv8/dHz3mqMolV4YxedFGGAwg/HzCsZpxUjVmA84mR6V0l9/h48wtZOVbVXjZWZBYoL
tZew/2DLONrS+DRfJxkrCi5xhzvocHSfZndOCoY/dLZJRGpi9i2MJ2uLxcRl5OsLZi9XGOMKyLbQ
YfE+ETWyd3kK9sc0DBSvsbPyKhd/c38dZMT9LtxbsovEa7nOiIjwbBsj8LOiFzY0Lqv2Ou5iDG2i
8PRzIju13LHeAYLehO7V3H7r2GC/wQC5aUWnDFMV4++/HWn/BAKmkl5gT2+v9Xpwrqj65xWrYoQr
+sWBggIb2jCx4NjK0lkOY5BifX9tPt34mDXp7GQG6rTVyqKLCCEPInGzwHBYZpxrtElf8ou+tpwM
/B9W38nnbOjN9QOmQ6dgTfAgXvsNyQVj6oF7Ufva15amJ1CXRC5ChNbhLCIOsCSz1PQ8G04Vmnwt
X4ujJdZMxYXLFFudLXEF5WI0H43zC0HJotmtzUt9N8VsDox650DwXghsYbhH1KQkI7pc1KwQ4kRN
Q/QIZWyYqEUBLDuHIMhtV06hzWMIplcX8TZflKxyP2TSTj54R2/A165n1TfMhkV+TkQJDwquI371
vTewflSqZlvChXb8IVGIU7DeVawayhev7N7LFOQvfdV+cVlVNLeFHE/3x+hJAsnLQt3dvRBd/rN3
y0iigWXTCOnHUHf4oHM5u6T0zedIn5IscVtcUE6yTa5xSRpvt3mlF2eBQPrHdCZwg2LohjVh5vyM
8FoXmxIIovbUgngQowy6A1MMWJacjQQnKfrmuc092QrIwI8dXHXijI8EnwgBCsEJEIYVC/F1wmG7
aZFwHCNOpmaZfnufFQ4Vsp2LGA74MSE0zYxzHjcdW0jHfZRGGTapRHetQ6Hp+/WQHUog+cD0SikM
7u53uYh3V2I4tw7zbjyiFQEZxkTeOW4brA99BO/SGT/hFOqqr0dbBxJNdaEAuIQSYPl6FlzrX/+W
KpI6chMBsPCKCrAZ+avxZsOrJrisQm98rqV8Q1Bt3yZbojRx7QrxUIjYZDjmeA0zJ0FxD8CQILvf
5KC38KopbVPZJvvld1k72wp2REBetcNUcFmbdUUjMdVD0jB/80M2+33G4zjsruwh7J9/lRkVb6qE
Tt57hsttp9OKKDGBHPm9vEwsX1jbp50RxqdI9DtabsmzREmvWJq4Jwv+K2WFx6xzmOAXxVUmFVU7
oorBluKJRgpdI5kS86PLfP8Rl3KBTf7RdSoT8+DQIzp0qg3dezBgtknlVHbRJfvVKpgK+HxCDzca
bt84XUr93MVAoQs0UFkgw8m9yxgKitStt71R/8rIQ8IwULGdtGDzVdjzqvpelsxhYdj3fy2aM+ca
tOgXKOssA7L0PlcrHSk4vNctG6G7ws6RvM1E8JMjlAE+9WEPZrc3C90pH2INY03DA59AQy3mp8iq
k+bUoWsncbhgpRB8rOXQtn1Z0Twy6XR43hdFBuS2dgapeq7ZxwDmcLZMNk0WlDS+xL/05c9BdyLH
dFaw4gmOVfZQZB7Rc8i8eRRKHwp2TESZKVU9zvo2zqLhTKMz7ehSNvbtqEmCdY0hn78/FzyGDQ6A
hCo9+pPC7eRPPqv8TfZQpSNBdRQgKWD8CQtpEdK1gBBDdhj65yT58XqxXSYInR3tEBE4kqbY5rqy
c2bRue9UyKtL7ZKmz5rkcKj3rHGEcqITxW1G1U02X4vuS4phwDB9pdRfKpvLjOghpLJDwOdnzpna
5mFnVL7G0TaH3F9/AX+8+/iDhdHrJF9F1UND6Zb+4ALhSqJOoHPY9H/CWEwoud967KsP9SIzemy/
j6QGHGu/pQtrbqVkgqNFwyb/qfKRq+8ApD5zVSZNNT/KnNI7IkjrPnVxvyk4SWje3WjvZ2S24+Mc
o94WuV3J+Ecb5PA4z4cO2BusrBmBT/0mMpUvwkdCtc8lBBVvPh5mhgrXW6P9GCyWNMDmJZeJkyi7
iihFmmjZSsL5/8L0hZGRhcIYQ1MWgG2YePem7uWVRkObQhWlZ/52l7Ak6uXiRatrnMDnqnkUw+0u
hM2jKsa5dN+kMsIn3cOqMwtJHZ1oAYyofqcmnb2ypsKaM1FUx2wHAJytAn1nHgF7TmKWyFlMr41i
Jf9HcwJqx17A2RznDZ3z3pI25OyovQ0Y7N9fGM7DtCNAmrTZgmKgkK96a/szLNCTJwTrTZ201Rel
6Taaxa5Kjg0ihCmr3YvZFS+PQIPhFi5VdQ6G8ZpaaZYVCnfUaGg+qAoeAf+br8UIlefUL0iX/8Ya
7qFiAQy40pFakmxfN+m8GMf/HmJu31ZzGLBLHJ3FitQhVokersm15V2ubZ+Q5HggbulMC6gh9Cv6
e+1l/vcs7w8PYW3Aaa1G5oJd+x+GtiFIlvs/6tD7/NvxCS+KB9GfvF/ZcZ1pRhgkd3yTJr+yQ7Tj
47RPy+3+r44gaTqemvW+tPxXrPL2sGZ8Iqk7m1lS47Q3CPQJ/FIxiTmwb5MgjbHR9Qk8sUDcR5bb
+Ww6huLZQbEhAk/XIeakPXG85CwR+c3ldw3Hq4wcIy18H7MrrK9FR5CrkoxBdMOG3Ne1kAQu9zEN
WYzL6PrtHl4Hx+dfhGDJjZURL1gn/wwAIigZHuoNxP/xTpzXq8gIDNiU6jMd31kYrND4LT/AMlzG
nLFls7NEdTu3J4CTq1irGJcE114jVGrMQcEQDLkVIfkozhZFJt7qMtBCLyg1qoxOg+Hj9mL790Cq
oqZummcsVEYoYr3R8YFFIFc9dZeDJ/Kuoke+4qdr00Dg9RI5dO9QBuGQ7VM/PObY+gLwKTrB6VCT
h3sF8SC3IYCE7ARLM9wrv2WrZRp+VPEQK95rLA6OJ3+RXwGCOYXILxIMQyxDIpZ91mcDB0L3yjXq
CIZg1DbzwyCnbKcS7DMduPtYjiwD72ykozOcPHrLkFpS5Hh8Sp1pnDjo4w/gOXsMR0Rir1dVU6Al
JYOCPA3Cym3ggggpeov0fzVHN7RTveVFjshncda4yYZGgst3dfn5pSijO85xECKxwH2Eb2ciY4dx
nFyySKHEWh8kP+OZK83KJB6PsYQ4cRaH6d5O7FIUrz94VgpArJ5EQdozCH8wzZnFLCEidICWhWyF
i9zNoqSLo60Je2VFJoSIpERYvWPUYhBmwUGng4U1A05Q0og3CbnCP/BnQEdpSuyQ7IGHG6SAWfu/
fgLJi9G4oIvEkG4jH3IDIjMyWU66+LJN/MLXxV2IsUNE8dz4A+leukEWsum/eptk8Xyohs5I7tDO
oykEKFmKQfpFU7igpovGrhD40OXDtK5zCcsEOMR6l7QnidqRsQHmrWm0QRCjlcINrrctqGDc2d9C
ore1iW/vMYarpbHHNxTGaN57SIUA5n9Z4ht1cmRsLkB5U+TWib2HgIlTmrADZpCEU/RAOCvyErnK
fAcmb/IjtgtK5fGQ9DFOsPPFkErojyp4dO8LElWtT/TzHBUmzkMPMMV0hhXlBbhup/NEvO/hMa9k
kXe4DJiPaifH4FgRWu9wIJ1lantrgfdlJau3Qx7iHb5x3dQkfy1jcz+gXh12vii9pj+X0oBAH2XJ
qQZi/pzoG6eUFBhSVAJBeaHTT4g1LLjYcgrwFzmPRBov9ancjKXHp9uoEgQm4yDWN549v8pAfbnj
LstmfPponmim1WOrEL+6sGc4biuJYMEMJNgLr4i7/D1mKAwJuCXVZu2XZDq7quM25Wk1ifiCs3nR
xLyw7bApUoid8o41vT1+Xy21khSHHteL0Y81Np4VC2yL0Mv2nCkAmOhYFA/i/DhP6MVm0H813DX6
fhTuE2TjXpDQDicbNI3Gw9Hs2t/num/x5zStgVValiNv5lMm9boW1T09x9ZpvyoDPJxrS+gxQNeO
5T2rT0YsdCn6Ij5Styv9zVb3MZ80kKt7zvUJHQZBqjxepdMtf5T4+RjY8iWmcCU3Afa1bMtA6VI+
hmIFSFbhzmSvKaTgcxy/lhl21Xv6ANq2DIv0ufbQOmkuS0tt36NEPZOU+OB2tGK8KoiQA2sMw1Pl
eX7V5M4cY68pGdcl3HM+jNcCCu+z4KBpOGhBwWe4wmh8x/TMivAkEqKFbyks5t6dG0Rm/JRpQ3O0
ATpy7bho4a8sDvzmqwjRYd30QFiQ6jdeY1D/1aDVdTURbBb+cNkcazXQVL5EaWoNbzqqINtSF/Wc
HYIjYh0OyGJxcevO8rQHw6xqrVf1ft9BgSJo7rQ4zY3ggLV+DWyVWGhbb0keRoo+t9lmFetWY6HT
KU99TXpvMhwSha0Ap0iJVBtvy7FmT4gxUy3EUIrLfPkF4w67/DmGc3lFrH06riCQpgjDDbnL46Gd
2fLZFRv4uZ7Mx4Uq15SrAfpkjIvq3OZcXJiT/eeAz99RH42HKZObUBxB4KiN9agG2UFwcQb2+p4l
V5Pb8/RpmFCSWgBP383MQ8ECNqkvLmSfAdwUiyt7Yp8xJCLb8Kz1JKWRw7dTBax50hCbXWiJNrrz
170iQzWY/Orl4+eIt+KbEqilW6nqA8SF05eUWBu6/qablUEgLkV0yX9H1tPwXNRKuGJ9e3CdleEe
1PA8U9Nqj8VHeqN/JyHuss6Zab7KyWHq1pY++1E75+YJZzXiQ6yFNu4Ha1yIk4OHGzi5do+df6WF
NOkMdroTdbkLuJGAdiNMicbtvW3vBz5e2XBxufUzr4Fv+Gn/WO5Guw0gY1vY7YepKQWloUtp/x5V
UIhqPQQ45bCCCSAx2knhcCZFlEGUfkYA+rIy90RkqFqcpwFiU1Cxhrn0Kt9B0Nt9Oe7NKw8XlNYs
hWdWicUjgdaai3FOcj81sFiryFLCj+zf0eMJeJj6eTEXuuStgRSp1wh0Pwo3BtmVjulW/UmXOrl3
HVHoy72RJN481hWWMRA9Smxm+FGAcIQHB/vPZILbzWlHRfwsr5X9sGQV0VBZLSc9qCoPfaxtC8oH
12S2DR8N3YZR4OUW4T7njrGLgvL6HDfztpSVODmkae49xkdOPz7Pjyo+6Skv090+RA3O4rK98EWP
w46H9/hylBQlRDICdbTw9I92wpGFsDzL9ad6I105Lw3+uuc4RQ682/QDzqyP3IAtrACwdVUBYJE7
BbZv9XqU6+R2NJzRbXOQrPej8jvtz2JnZ3AxlISHqC2vDZ9uzgm2wEbBeX4PP0yQURClE48vE2++
62eEdSXEj4WB8IlaAHjI+DhSGab6n/3uIQOg311E35bNCbHuffD84Ys2Gx65jw94W7ERHOOgHGYZ
zoJ0o4hJ0RCaW7nRS196SzRVYhL2U18uZbFIDwRXPXfyNisoNvOCfLeaTUe2uskiss7YG4KT10GT
YR9ga/2CszFY41PfMdHc9qc/uiwIqjmSDllQoHeQAq3qncWiW+2fdIKgBek0PIqQEhvPA+nGoh2u
XDaVXHrgzssqVDLArshprkpZNeTzpIdYiTYpMVjr8Ice1VnZq6NBc0GOJPqBzkaldp/LX9AVY3XX
WNxj60Jepjd7c2WHGFtSTl4ArX354dS8ITlfP7N8/XrN0Me/H6GHdiOKHyqfZUU5XylaFLy+4d10
hFtuiKPuI7H9tBKGUWpJ6kNM/04QsRqDRyNUWj6libtr+lKd7jIR1nmII/txHjC/+vFrtvRy7pS2
QL1LjPV8gPQb4iZLj0YMZXvEZfsuwETNpeHQ3Sl0Yy3l2xmmVBABuT7ILOlZPO6A7hNQ8KE3idJ4
P6LQC8TlHpEZmcXROP8IU0rTh0YNb5vHXU0Oae0q0dorAIF2eeBM9RN+dickxqTRL8wa9rI5sPL4
nvbPCMRH8H4FUcxBWtW1yHOzfetewLll323JBU9wcJUkU0MTQYdmyRYGcRAvN7rVf5xukUN3ib7R
jXMiGAaJBxguaATnCzkD6Ukk8lN/vxdSnz8cFb9fpm1LNmYKFwAWu2IDH1IkdVNT1cwi/Zt4qrK2
F8C5XPTnMwaOUKHSy1ta1Xhk2Eiq2cfvaEh+s8Hc+y17hfccDCITy/Ix1hoQE3wKbSugCjcfhk4O
2E2emuPo6dSs+SIvmavqPaR4dvAX2bMdlI9HxMbYjKWBfeDvAKsi5ZbFp+rTG+epAJLQMYJC4VW+
1+mScp5npHiY1JNIeVkMvTNzR12jjLwOLxfRgQ93gfGgpcNtmP5iCMhBVBfZwQgVpLZpOMJswsLR
zwm/tVck0uPibNb31oXIf3MipMZubTeRwTNzcbEx/gkXAbh6mSW+G8i9AqA9rwKjS0ZZE87wI8bj
Z0zgOJM9Q/TLb3NWw+4n77+SF+TssH+fCE73VwQdnSzdLCNuM0DnSUnUulYOrGlcFvQNLjpSUowd
l3J3upiU+PgJWOuhxY88Y5bQuiC0HsgvtgKBco8pPn+sUBG+h6dhM71YpkdNXkGyEija1sM5L//C
bgxoHzZds+zsVqLBatBJAURbgDHUVtCFnmQ23dVipFo2eSmjjQA+jlVNGdMeu8WuaXRyeSYgCT9L
6K/AHk3Fh6BzcoqTwpWlfMZX4Slr/2d2PgwNTg0Q/PCGTnRK8UbNBvX/KApsO4otcQdUiphn/2j/
tIM4qd/MK3ARH+/sVg7YZgi2qjwFrDzbj00mO17Fum84MILQJILOmdwXTIGEZRsV0ZrOmAeKltlx
kVaarJ3WUiZF1Ioioa+MgEH5R58EDkRi47HyUxe18acc6FmSKSswjLDCvqIqD7SaxJLwteA9heQI
gCQcVlH/Gnzj7OsrvbD76gumdJFKznmHvcfhpT6ZYygH67PKDPfL2+AZv6/bhDgtxQ3J43EzHtgP
S5YnaoWWpDjjCmXCjVHPQrY8fpwDEQsKhYa5Y0M2cY+V8hTHjhlOw2NtCQifLJ3hjQbmBcPL3+w0
OcUzRL56A0Sa5ror9V5Bw3A01piVyPi7GhTKkhtUeQPiJKQuxOrcRlzQcov3Ko6LpVciXsuB2Zgq
Y5bf0ACSxzzmV54s120Pcyr9p1viSqqljGmGdINq7iXwyP5Z+5ZL1mvybDw5TKBXoeYZ7BvYX8YG
c3ZGiRCvwdzIwLbe1RLGpIu4vrtNhqli3ED5gdA9rtkcVY3hRyDauyyl5Qmpm39aUbxbDHTTvlJb
SHFxU4th5/X0ALSgmtZmc5TnVhLvqv02/W+eFMDl44QVqh/vD81m3SKmV1ycoVHYNab9e2wdMP0N
pLJEIkP77C9ciAkDSVGfvbyRufSBAuDcbIy0s0aNasbTKroDt5ZVObDbyl9Xyg0aDxW3ozmQX8db
0L3uKqOWdHrHGo/H6LmhKaP1n+r+Ef0LP2e79H/UBBUh5RQaUamNt/ppVHHHSRTBsh0SnumkOXEm
mvruyI1NT9NmQ2iRoJpr1VcGgh8JcvsCVRwLPzU5lD9Jc95HPqxsTlXtUpbJ9l9Z7wUOH2Y/j2ZN
UUWOq8ME0UE8T4zI7v3+10x9O0eN5X6kiAJYv8Mqd3zTXTYTJkEvza5VWCcWF7iRpttayoxpIZQO
ss1/LEFezy432uHUTnpoWRbEbPv0k3EqghF075EkptCtllBQiaL0mhdBQ2BBD8ODp9ba2SMzrWeP
qqDr402jINIB7sE8zIvUdk9aoy8RQuUwgojVF+WR6u3k2CuLkRffxyh9/T91B+Z3u5xMSctbCW8y
6+lQVNqadEXfJzHVDdokzZena12NLXZzQw5YTuqlkfFStIZMAgQb4N3w/OAfQJPQjjhles5mOkrP
/PoVlaJZND5UCzV7h6wg5C3bl8mw93KTXkIPNuDV9tkzSW0JOYvilpeixErag8LUbqr1IPa6RuPY
SWtSZVdPPmRQ75kTfIa2D60Z9/QvxvU8cdZQoM4wb9ZFot4+REIIjrpJfjvBahDBAQFtQ4u+rdvB
8treIVWNtZFvjl8ACYIgF3KwwmOwNUKYrMRi0cUlaD4/zkH5QV4xjeoMxmzI6HRi2I+vvVmUMWPD
gxwmdGCQgFPbmUEB/xa5bwb4sSqnYHFJ+uyjxS9sETQl7p62XKJa/v9gEhIpe3h/yQ3ahax9eveS
BZrb08d+I7EfyUa/ZXKqeEW70o8U2XBHw2poKoFYBjD0PuYG8Y9EkrFN7+rBeLwdwLnhTQsZEVXt
a2eUObMeIR9bOYH7DqkBs9C2ELKOQaI9iDdOatIM6sSHXCQEyOq07SfmxZwa0PphHUdiVAwnueZZ
XAD2rEXvcGcAWLucl0ORb8NgmEx4Bf2aunUnFX3hDk2faKEpfoI/V8M5/BqJEmqi3E1NuMcmDwEj
/p0BWZOXVJ3eyv39ZvLcyWyQoECEVIUt3JizaDE9mATbpNjUZ5tpwquGwPiwIZL5J+chzy7mbtWT
UhAfDWuF5DKMlv1xxOd0r3eKPqw4AfYfXdO/aS3AwGgdFT+yOC3MkS42rUg+Jeb0ZXTTbeTclgTp
fF4z5LCuaWXboYM4WwrOshVwU79EKh25GCAFp748bPVyw4kTNW3F72pcl4ziTaJPeXFOkG0RUfc0
zz3OJAMh41/cQMy0O5bTD8Ov784UfvIrnFLUorjAOkDVYc4B8gZhHPDz3sd7xJ06NSTpogj9ON65
f/GMY8yuu29c659w5dhLOdBBXgWwZ8exfWmlmHsZ3hQunGbCR4kBbL2CQAyX3M+6ZDNwUVrE5Bg7
mhSBFC0o3+YAqM6BGjKydZ2/ZydUiL6J5BJu+CPGo53SiJ7ZLzn1vpY3ueNGg5EmuHagHTGcJtlg
7cN9B8IyZSl9CBBd2Js/PIfLMHV8V7n5GRazWkkQ1ujebiomtzyWiWs5ruPEWdN0fATv829Rf3yG
zJhnZv4iIUxXgJP5zDAWEL9t2IgiZVK53wl02ZwJmYo1XcViSbEK+8uqhrcAakIkzh0tOUaWfiVM
31kdfbi+fFMZTKAJQzYsV0ZFKlPHajqc3sCiSol7/wbMgYm3qBkgWsp5pHeOoXpnr6WgDf+kBmNi
0xXSoBTFlzUmm4/mbKVJ9lY43tFanVjJf9SE/FPMHjwVf0W4bD18j0f8iRJTspqAhl06mt3cCgXm
35ps3Ac1SRi0zXFBdefigEt4pvVCriB4o5YVhatIt8qacsM8vfkEGEgY09WjQPk8PWX71lIRRCEF
31iNTcPZpDY8BC9dLa4QXHbXDi0EODP393YYrkpKPgVSS5fMKA2a9iVhjbJCKR1n535IOSRwDwrk
MZy2Rcrd5TisEHafeRRB816H5SgTs2b3C46y+gpzAg+jPxEnH0EVsjT2clkm0PThTGY49OOLQsXW
y5kC1aov8mSvnKosxAvXUSRWYeL613YDN5r1gtx8BtxrKhy39rmT4LsE6PJphhghEBtm50oQbHS2
iLYGXLBxKTq0CdY4R8TILs05T1HhPrtRm2I64XEcA+TtRx/vJDQrJXzb1RQS139ylMHEzZLu1W1d
9V+bpvf32+ck+CpHLowwvs+J65Wfcnoz2rhmq5WpWjM0zAcJ8Hif6C1GgYSsPHKAkymY+PuAX9bq
bN2YJdhwoJvN0unLMfVdBb7n+v2UfTfqrGFsOQvs37hw0rY4LZQoD9PdAQ3wm2w0xSYUBWT11Dps
GUf7FnUnSJkrogPs/gSJnAwNdS9aFu6Swua3AJAC2Zz1IASoM9sJ8X2bIzzdvOA/bSoHvBWNdG8K
fkVN7SeHU6a3YvpQxzghfYDcR/NVEOnciqweySNBn6IIZxMlnCNaRncP/hrL8Gneac1/XXdcgtdg
zGC7cfE/nVZ6f/aTdo/6sNDea0mvXeB1qQ1pkRjzt+CF5rjSU7+ffZ75res2gBBt3p+eV5yPs6sv
BL9U48kJ05jAbYsgZn1/+fFsTmTgAFPu3BDWQiL5XQ+Lvi6JByPtsFsOq3qxnn7dTyYPKMuVPt5m
aI8hh5MiFYtce6xbRwr7INEAcjKmDQvKoh2gBgUzhDxIgKCvSViiq+/Mqlja7e7znXrSmqoelqdW
agFGinXr5APpVmsgtDAVc9dkgtfTm8v0kznfHMm3p7Gsod3lZf8RQxFx6uhSFbMx97xFgXCg9e83
0eDOEjha0kY7iwdjtxoE/1XcZyqN486jZPDmOY1YfwVAj2Ev82GjsnYfLRKg3nARI0copNcryzbF
hbE0jNp4ZGaek1icXnsp2dhnVeGLde7PSr/POLensU9O+DzSaYQqsPxsQvmKLaXeNgiW0kOKmK2T
6ddrz+4hjDL86UG2cdDrdfJ7yfCuTR6/cOuLiFi/FGFHCa2Cy/NIIUrwaBfABeLi21jsi5Piuf+D
l7r2dHhEltK7id9i9LQH0ozUzUzBYDv8xF2wgsBmYuItj/VUhli5Zx/p1sQ0JT9vL6F4krNFi4se
hrb8czqY7GUcE85/oNDVXS7JsqBNJxjytbAguG7S3HJU/v3YTtNOW00kUZ9XLvof2MqPamnT8P/s
DOkAyvI1FC0pjRXYlUofZCVGDa0Orz3nUY1xLtk6w8AHPIS59Ml59cR0EPozXi9ANGO7TWeFg7NV
DhmB8gla2Jkk+zDiWHSneX8x7zQ+K/lcoFDB3u80rXGHqvvJeCQxTBkGEX48H6/49eTAb+VZG/2p
64XGfeG5lt6whfrSQKm5pM5kC914Huafe7br8v5e4AvdsF48ZjFmOPgQuRoRbP65S8EDjIOTsJM9
I/C9oOdLX1ySHGa6K/96SV8YghYQJ7+21u1hBShfLdP9li1EWNvxgl2b5Wb+xwuHBso0+OFfsudL
o6Ci4TCc9zUTheURQqRnJ+ZVNEl7Hc7c7mlPO/KTC5JxRnRVIJL5c4tTzH7XM3F32cA4xacBSTbF
oO927kOhOnYdl9HB9Wdmwe1eu9OY8wUTAeCgX20CTO9N96+xBpeeKaNyLegYu/NSZ+tfK10d7Fnk
J5rXVYEA+q2gtgJpSx6aaGjDAeHeuC4shhwvieyXgNZPISe5iF+GbiBQM9gnc7v5TWQKSMjUs/dZ
1YAiKsFBNtJ1+hqWKw93xxi+WSoI97k1LfedOKwthtu3uYfL9ehpeO+5kbfuoGnRW2WYm1xL5/RF
loSJszJ17EEevxoqHs18SA21l63TW9/P+E5pRcWvUJQdH80wXrtzrG88dTyWf69iqKu4H+dxOvDc
TeMgh8lxDvkjfEXLMKMRpeEV3kokFLUvtxBDvFPGVUOPSA+44uPia4dUYhg+73gFJEOLoM6SJwz+
nJ+Icpyh9z3c0Ct9hw0hfdLilLKBzUdw/bmi4v+kBnp8i7f3gqzaUtmTPkEJBzM5dSyyEtZowVdO
W2VMXOXcxMd3/pyr7lcEAPIUeDCJUpvHJj449j/Pd5BWJuBxbMos+bkonWgUtmhUkfVuXzCpHMUl
aVndxda7hJBU4P768qhwZN6h8PkI4VOPX8FWUoatitbO0GEOMYYWu0zWrexI2lSPMFhPOIivQ1vj
JobI4xRUxlJ6ImpucdjADTsqq7bPyFO4ioRzsGMPHKqTtCBcegyWRg6xJ+ZXJfSksqQtMb7Mj8Vz
/Hyu5PsSL1s6sX1GV+yCjV5WdTAT1TxGzDiW5AdlmTR2rO5hlYP2B8ERQmzwwVdt1wU57EtScMpO
fcHIr3jFvKxzR1xLtmPigKyxfnFikfprTuNZBJciHE3kKNSFY92BR7aINAF6YhH3opRayd6Ff++i
u4HyG4qE27/yLdsIhLvMhYirSLU/KFdPnrvUFlbXk8jdmBSlbNxoQSGW8vWGt3+Quda53FS/MsGV
lrH/wlXA/PpgLn6aHDnDpcyzH00Ix0w8HNIBSME4NmLy9DiFfgfYgjUwH9m9lsLkRvG14vifWpwS
/dG6aPgho4jVmfjIALY8GhBA4LyZawxN9wq3u+hQuLO65R6uYG89s8PL/iTWUj7KrYOF7RoKQiPv
jsKrkOAo5GG2p80IZADdoNrItH1N8U+Yzt+eO9p2ME75JfvD7KmfajaeIw1W9cwCMF51paoIkrKd
C7NnPD7WlJt2xqqB8zrXlAB2PuvFhMoWZs63xmMs4xjisBq8mS9v9R6ZsA0I2roUacXpp0gIzldZ
fyVQr+O2xEkwQBBzjMhXUROECb1lTYukZzFOiBUUDnE1mym41h9hWKGYjh25GnTSbbS840xTi1s9
4JY1qJSoUr2veIU7z+ENnFL/Z7J3lw2oNXtT7RAxOWFVWglbfSCRBbD2G+QTSZ6vKY6y2u+6E4JD
dr4+hNvAWUBh2xXzdPDiiJnXh3lRG0h0udn6tUZZWmuIF0CjZMRsGYnnf/YwMlD3azJbMuRer1ZP
epgTrUMbMaKq8L6nnwchBIYD0id3fxk5ZUqycpXblUopmqUs459Aa7oRTvGO4VK9HmFYHrC3JbpX
5nHXAt3xC0nNC1ipv2GRu0Pe5l8KMcTr5+c9697mhLqjcPFgaJo+eIexYLT7YE8uCSSGQIYhFUFM
6Agfkk8QZzhZ44OL973bpSUw/4UVJLvCPji0f7sm/kipjyWb3QmnETd584hf45o0niRkwxuN1VkE
yJAs+e/N1pUautm6D9syWyfsjF1CzIMfJE4I92+5aMgVnjzpWuTRVxThrARPv5F6CvEXFN9JhFWM
4Qlm7+JwS7JYDqe3W/HiZyRV+436vOwU2k6znDaXplcGNO/NFmAmWmE8bB37RdLTKkLVF5vGUAmN
d69a+/ml/dWxtkpUnLT2osPRDrekZ1kEzRaZw5ptdpZ8IYt7Ce/gkqYxHpEIC+Piop+QwTAokOPw
QgcGp2T7Xg8DFOEHCk/3AHgNQ4MJSewPhBU62dWgN5o6ggW787hf6r/N/Xm2y9guP0q7iHqMZUuh
g0HRKMF7H9We8w9YLB50qL7QMq1q8xOhmC6qQZW2r9Gbj33PFxpWD4/YDrUIm7pt1t+vYf6X+5gi
fok/RUEyBNLdV5772p+5i7g6/WuAW9eDMTKwx/UGbfNKRgAwzLJr/PbQXHb0kFkETO8oxc4n/PGf
FVtygzvM9TLS4ki3l2fgwL+DcMzlqOHwjl3lVt48i3QRGQrAmr998eHTWpkIQeTMfV+wcD6bw7px
SzDAtDfsokdmOi+sGDLkBlbUL54uh4E+q2u+7lPGTaiNdU3xvtiAgFf7egOgMGZMHh6wAJD/I2sc
jAO8tjqC1nU0oJU0TXX3DyPN/bzs8JRkchDs/O0W+UiCvOyZ9L46AOFZ/EwE/c/C6r6kxaeBpaac
1ox2Zfb6L5ZYdhpoq5BnEgdaouyoaML+jQhCd4JzZ8XM58gm559IJCzyqv460flLuc8qwbgZfPJo
0MtHgYYusGHn4+41Zye5l9+kif0lMlE0JQ41OC3Qwxiagd/NazA4KlchSKSxZQdcrrM/sGLNmIby
K/Jile9/n1c9btAE8lRrQghB8vrktEFc6nM0HxqCT/vKodaN5qAky6QPfFaAIfZ1AoQ8Kb/1VVBM
qEAwTJK/vcLy3WmRGPSSyENe9qe/IY/tI1JfMbsx2rOdd8J2RnqAYGLVmAZvLkWVkGlKRmooMk7O
kk33AJ7OhAD3h08A1kUIKNPRicFraW/ZDOful8Q32uhEf0ejS/K+F8jiUoF8f5vwmbBd9PybGdK3
r4kCqSWO4U/YUzNONz8WkzLdE3YoGp50nc1/u/OIZ0FGgDln9haYqSgMRjcMQ2WT6i/lmFpBt7hX
qnDwSpIdxdyXYw+VI5RfLSXAqeUu9lLTZ9cnCi07jPtU5scGJon26I95BX432BV3RSLoFzxfPQgw
X0PaPDgGalyNTvgzRjI6MKL3Aq8JGbOfmEE7ah1tcax01uJKeqi7V4JfcIlIMAMnL5mjEvAwFm5y
zwQYJDwjwFAUvmL4kAwiQX+N1RDO7LXR/8vCX66azXQTbVQ5LxxopLLrtfhV/aJkbShlOmYavRAV
5drGaqQBQPokyakeQizBoRLwEhdyaYw4BqweXa5CtV0OMNJ2c+d4YH2VOrEinga0DuXIYCI/vIM1
37tW/HSdReAf67bGCSxCcWotA2MTWyl/iSchF1sZmA4hFoC9ubID4feBWoCvxM9a8zpedSAC2yUg
CPy1zvjMkswskdUG0lzPdiqArzfhjLRLmOtflZDlkm2coSH9Upu3Gc/VQd31e2RN4MyKe5Ey1J/w
1v6C6/37BLT8VD4ofnJzF2rzt9yMGCofjVNJlen/1cUo9A/5ugGsMZ8fzQG9aBu56W8Bym55NWaI
mRSfWu1TT24oX308XSHaADgokPRe27YLYVTwVk+IpzbmtyCe9ndZ5qD3jQC6pgbxkUnmMQI1b+gh
6IxaWJb0g0ZVHyGH4PJACXvsLzrJlol6Qv2zW/1vnqsPdrYuaOO5mMSZnafAoDuh6N7muIP5AvfP
4bobI+gP0fKa5wzqwQQVVa/jXsGLyqv/rrgbC90kk2m7TfDL6dzf41RMkFhNj33IfQzJBlJPCsug
HvZGy9XTeTx84/GAhFwBkSkOcv9uew/xlyNOBxLjw1FsVjiJU87q3xTd2YsOilw6XwPRyaumHfKr
rCUjHRoGeqJSlD/RwVPaowrGvkCcmj2+5ad03lO0yQO3K+VX+gW7Syti3+F3vDge52ghXrVRDmSU
NbA0UKA9HU0Ale5C8prkoudaJKrUkesWpgDKegkjLRoawyHyDGZzk2j499Ru0DUnfmBYQH7hmJqF
Q7TusLc3HIqqCB3aVdDG3CF4Teq6tunO0j/UF+q/y9amPIxNhc4N7PcnDK4IEYAikiCy3YOFWYHK
zPNagLUXqYFfL2ZeW1zX6MBbJW2YkNIXnzoxCZg7b5hckKmNwEYG2EYfsdHOSbjpYw26RVEnCLYz
D4sSULbkVrhgfie/jppt4XxY0j74HYmUt449D4KUPaXTVKqwHgpkPCqYpGuo85Ah3j6pqSpmnNGj
Xb7zCzBTAPmuIL1ulpVvKCYSKfen5ZrmC1wyriMFaQ1KACD1qH5WKCCTf9ufJ4rtGng1eb5zbDnI
XwYhUhzYSRRSUE9X2Ekpwv1uwY553vuK5R7XL+RhzWWMiHH+C2x2ZYfPWFlucO6oShd3W7VcK5MB
Ba65FCUpSMJIY0YeOmVuWG0I0h2K/sLtXP4UFuaNs0o326XydYCB6T8iHXm0X+tAANfbLzT3ga8d
I0Pafbx1eQZWsSjjD2DijL7zNYfo0R3ocw4n9tynCHngw3yq5KMEybwPwc61y0rjlx/zLTo6HcHW
SN0MxRAeRJlFwZGei2sGgTrj9VAXB22i+SKuKWihc3Ja236x2IIQs+Ja6GgEQTi4jEIC3+nBj5eU
lX9HQGM9KBZKqlUDj3U9MLOpUXH15CLEqUqmG17Rptqq+PgPnGNmOZKy2dxjdHeNQq+P+2Xog/D1
RV/cfl0EebwLn3vKwQmqXF7qoV8Ec0xS66NGUuvPxqPQoRYE9VKlfLTTMUzOXGIv/bED0y8TRAaq
2rlwVX/9Zuu+KskGNXzVeHtIMMdbB8Eb2e+LFx+NcIi5RKwNXXM2cPel9V9IFTswF5y9W3XhebFn
PMm3IokH/AcVsJqpDN3lhZmokg16qMshLRH8BT2lu4+3zQ3u8phCYjIdh/TxiZig0xmSOWlxPMZC
kVkFWmjeIN2wZXkxEGtpUoK26uT1bumatmnEFlAuV2T3Qx9WDCmcUMikGbMHI4rA0Czyih7ZMlvC
AWgUcO5ih2PfL4sEpcMu6xbSbMY4gyc2S4eYsGA6sOgEgrCROxU9d4G2SHG37DUtxZBrCzr3037h
1gDbB1MJnyYDBYEPL47uP83xng/dLmU3ZBGOXwgr8GwrGy6p234MGiTeANar/WpaqLOa8h8Pj7zp
A7eNEPNdFOQkPaqdq0v6LDW93q5nd3zo9AOXLkSlxgO/D2E9kicJZVc4TPqUoF9FtBVvd9384da2
GZR29tDACEzaaDpDbRvAoUzBZzE0Uzb+S4soK2VyQDmkd0H1pe/EcX+7umHoHJ7BcVi4/O6veqi2
R5+Ew5G+SrXzHvZcX/UM4p7wzSpoJkAdT/2Bb9z+fARNZgbWOTmsFU+bBUMkbSiYgRZaEMp9dO5n
laXgsQ8LZwV6RbX8ypWOi8pVr82fTGY68K3UFG5wrQFTGlmxj8iEGFRblr19vijd1IgUol4Mf71X
fyukewpal0cFwKAB+Zzz8PDl+TaWUnY7wIa1Rjg7Wk9Fnp15X3eWB416KuTqP8EXRKmxUyXdBfFH
wWucHB8gV6Kacg9p3ZMPLTp9gYuasyHPyU3hwIzCVbFNQbF2XkeWC1uz4H+WTK38FiNM3gqmCJK3
wwTr6paajH0b/72x4cHdUDZntzLV3WliClfxAZARJDMhhvr8/OZP6Zo+tytaZfAuv9TEXUu2erqP
HEM1pYE0JpoaWZgdsqB/jeB6ljA8JzO0fY3xeM6Q2WlxSnvOIPFD7xXucjOzg9Atv87OYPv5NEwD
I7px9IxT6bOtA54XzBkmObedfCQSqQ6CjhqT/dwfIhLBJAELVrOGQGYhT1wZQTbfbm+bQopFvOgb
rTI9Aey6n9ajl/TqO+M3P9OyfgCaO4lpLDKPXtpMS/9ax2ftq9E2Dg+pJD2NtoaoMv5Isowe2aK4
4jtkkkie27V6E+FrbCaWClaB/WvJ/bEfMolun9yfjxgkDHyhbZiBk++SWgWLW7oe2NgnmEesMGEy
+ZObY/H/dfSSmLfoTxJsxn0fKbhgitzODES46RmZlnW2jgTBRG21kyX+fbicxRk5MqHCqRc4UjQp
0yn9qyEPOQ6jCNoORgAwMT6WTEZD7sHDBVf/cdFOYvDknf7DpAbXGX/9PGTG0H+1tzFAofogrOU+
8OObrbP97537PQUI/kA+Z1l0Myqyce+4R4KRQpmjN/YId8x4vseuPZx7p8kZywtz4qv8CdKc8xd2
vV7AbdwNTeVBUvaG2oOQ+TlZPVRFgXq2vNZupEliVJueT2jxS7+sqido0oCxnfI6HlFpXwjYFyCU
iGDwFWo0PqV42dTDzm5mn+EyXSumEvLvclCyjn8wE+ODybh9QZRneBxtW5XOPT00gVQkcjvTEz4+
EVEMt7ZXEMLLBpZd8Bac4zLwGbX8qcCv233gDR0V0O6ENP2s5rTpNR1HwVPkhZAKoAPFRap1ndvd
C0nwO1R3qVlpvSpPOpSwua9oq95EyYi5m5aKmeE9H3YQ2FXm9yRn2q1BfZTgKyxCigXrWj+4wL9i
iwbhqrS2WndbZ8nr73n7vpkZ1MV2TVTLUzXrOFax9LmEOt0PcBIqGYWNZgw56tzqFpqNXwgiK9oo
7Eenq7o0jUqyHVPnqxgIJhL3Ny35ktbxk9qWMsKAAxjOrQojqKy+2BT3kPPtQsR/RPc3ky5De06j
JjMVsr0M+gMI4WfNgwWUvG9z3IRb53KE3kKt8kRZNYcUHsw8uTZ2AgApuxfA4YWopxUsMqk9RcQ1
u/oYpAVgEv/jCWV6+kxgaBvxb3TUa3/weFcogrcLIS0ez1SS1O/E6bLEMMI4BPaIc9z23zvsCZzk
1TWjbX6NQaSPoYELvyX60/pBgzVcTE7LOdrvImSBXSLOkz4QlYf9l2A4e9E3VlJEMi/TndVAFvKV
RjWwDf+z3OBy9nGQfkEzLSKM3SUZokFOCwOb5GvO6ynrhIrer4GS03Me56uPwoy/Z4wiHMilw2ND
i7DNRDw19yczAiyN/IBi2BAGFEHz+312CXo/2GGIWuS6YdZpF70rmEoM51OK3Idft/jTYRbDeDwT
GWbOgijVFqOCw+TnscRVI+H2k80tsDZrhhXYS3+Ur2TKnP3+RTv/4miwInK+oxltDrC5EBQT9uQQ
rfC74zBc2/claYr+IeebpNnPmOYJ9ZMAaBzYeDOfur/dwoW5vVEng7ING7rgzEVEQ5jvbwN/7oV8
pZNlF7Ir20ZyNjqlmC6HPQTrr8yaHW5gXeBTJZlgMkiJl1+LibvG0NlvfnFNpvHqn6ZqAt1/kN+i
1grQ6f7EUVVGtB8/bLS0Rzqs3RoqyfhTx+CJ2yQoImaLpkCo6er5qqbPrVlUEupHN/9WCmFjx5cY
vRmoyArSFNhMGJle6wozhjGGAojkFL0aVYMZAtb79C/6w1cY5NggN6rD2zZ+IKGrjrod89vRVZp/
eEhzYMe1Je8hmc+Ou1RgBPvb4eOqj4HoPANaGqnqBnYteQcY0vlwG/nXMGJkQ3xmdFAOzPIEDl9T
p0OA3kUWyrnfCsvnW3Y63AY+FTnZ141B3LsWj9RhvpstG66UPgeT3hwFNkNOFXUAPR7cMkuTVCuW
33oUSuGnGNaLyHi6Im4ZBIuUFJhnMvgYbNvfFtzsbawyihohedvjmn69s7Ludal/vAYDHxPGLLZD
Hp2RZmgOLIkmBvFANzbmYijV4KvCf7yRYmsBLNsK3+D8bIIaRoLJmGasdXBKnWxLV2QUxzrh3nyl
D/zpvEaFEEK8usXrnzK7ije5xH1XqkFpIrr2SotRYfLJiMsXkG92tHUUxuYTp0O4YIwBYtv5e+8M
RlwVwqCxQsXPmWgbtWhJlATZl4FysOH5t8R95pCd3ZW9O06dYIjwbYPvrOPyaxSMrbOsrLju+Dxn
6byH1/eC+O0l+c0RGw5Isml3XdPvnEdixlzRRsjxm3ow4Q0vCIC0VGpLwBiW3Apap7axJtmjXG23
5NKgNSC8C6adicWEgYGTDySJDbyKY8CzADcGwbwrfkFJkU11J1QnYPftAUKxuwBCyHwEG71q+Rqv
mSTqZVMHY3FrGKhTlAcBVcem/r/Dpb1K/aKe0YievWO7054Alat5uJuU5IFxO9OSSe1jMu1097kh
KzGLEykkzHK6ewdCSSeZmKBp0nr5hhg/uf+8zePX0HghnPd0E9TpRVNS2sNFrK3dUEAESVI4MlLJ
yx9d94HS569j2vlcePycJ8/tlCq7L7s7hRrRYT0QCKUW2kGfuRfjn2ujMKsoIqlaVLMUd+XOvDmA
hHEQETBp55ifR72H3tE5oOClopTWMsd+4J/seV+oSZms6NQZ/q2QzBERXAYm/+GqrIFCkXUgGwte
/KwDhZmecp2XrP5406USU7v+PLxOQBvzm3nRe3/5XOIdZRee1/Zj4MaA1ZaIpUZy4csLJ/UWmhs9
LMy/AgpuHFcYRusSF38Jl0VNLKlCn4T42WHvT8dlkMA8LEPFj2Zp72tmA1WQRQvgf2xku/y7y0jl
K1bS96/v4EsrhBueSuKPGBQ+XImzyB6QPX1W+ZbQvm8fAik9MAd99WgHoH76DfTUWyTHZ1tqYC9h
VuKPEhoYFNz5/zq0BW8HeUMVjGHVe/93m1OeE2j8Gwc+nlpJ62rCnbi95Qk9Aut85urnJNNDYdRH
GhT/4is72QY0HschO08/gz19bzwnGtctMDgHTcAcwPKJCC40bmebaN7ULDVqsC8/MogPiW2PMQJL
Wt41wR7/gy3MriRDdW66ZqnVxNu7pM0UygpRnF3wjBuYJV+m62zW51nF1Sg0YHKUd4hyPK4WZ0Aq
6MK0nrxqlzJINkiuuWa42lleWe/O97KdTYCZQN3zKElCkvmkwNpgmE5p5EMXTQfQYv6MwoBNodfT
e5OQSW6eEKe8bFh/MzoctBZiRy78ynTdsLLdPgLLnCQAqQ8JTOYIszo7Zt/ZMx32fDmVIB2F7q8B
4zjRj1eNYyuAdc28U48IHFFdrvrO13i0B2gxkC4aMWC3IEu/vw8PAz/MmVMn6dYinDL+7j+joO02
cC8wXgIDi+5QFGFyemEt6ibwhOjSvoq5Ouu/cP1se1RqMPvZibht9iWlt03mJ+b6rROpIr72Hc7t
LS/5mbvnuidl7o4bNgPRGBmTvHFmUdRRQNKmuI7PXPTc4QRRmPOzIihymRj9HR49e7Mf8eUfugVf
ckOjKsg+maX5zRrURgy7Ct5HI6G74LLktCUZ+UJx9Q8ABS0oV2E8zxuQRJP6YblEP9boMb2W155n
hWZAfUnXoqC4X6xJu3I/KeiCS5fJdQVIK4gXTpUuhTCNkjEk/BPnJyKWZPMTVA++IsfS1jH8dNxv
8oBxLBYAz/uq0E0x0voevGPoiAtWqmt/LjkIJFt+iLaMYr9T4PTFCE727ZroQHaewEkwJh3HeTMK
3Bj+l+s5PdJHXJOZCE82JGgDyYfMwe4ne8+FtG6e7QaRxWeKxEIybdHXSY70yHIIwslk9dGowcok
geCpekqJpZ6ZNTZyl7GMOzf29RK/ACbIzATSejMmZFFTZAbwqPzMGfzYvWjjp1V9w4L3H+Qae5YJ
kiEBdXQwxNCceHmnadD6gITUCFZkwDcFMbiw0wycdpNRkQ1wvR4BhdDY8QJ7Sxlh5tWKYVwvne0I
ors6IQPNc6qsVUKz7QV9wyfv5hnA+yCeof21u4KtJnCaa9JUsfeNrJr82h2CHAqk3Wntf0OmKNOM
VQEf8nRB/aR3ky0faiM9xczE+HJ4hYhAPXH3FvmTgUKyl6qSc9VQSlUDqMkqnC7HkPNJUiu9uvi6
OtJdANup1CwEVMfrN6PpHaYCtHqmBHi+2eUa6Ih0zkgEHflrGZ/rmH9J/JbXOLYo28knQSbmjm7t
REj4A9MOgnKH+5FxMhPyXqfvLzYqr4EryqaBiKQpeCtlOi+ThniExF4TbAwUzX9I3OJsIUoMjQ/S
UUiQkdCr4qVYumAeRl3qU3tZqRb9UHfL+3ZB+fZEm60UiFGZY0lCfk9M8I0Jxg0WFeGzqtJ12f+3
NIIbdJahHBVVp2Yd4PUoRdjcFGDeSLmZziyYpMj56QC+kirajAD3ucMc6YfgwXaglZ++ka/W/wUW
7omKiWTH3OLsuD35N+i5KczzyFZ5shehhD5cv7d4cqbg76WFUsDjRLAumo4QbWUW9RLSTxVXvrYF
CfavLbpzOqOTcvttx8Kr5uJroflH1XmowzNjlMawgTwk4i87WAA/XWG+Kh6GKc9FBiwVBiqHVoFe
lZoR6DgtS+xqvpJCNlCixpV7VqK50CKBMHKZH7ylRFfFx8utxKPtfD8hXaneWmXhzQ4w68XNz4mY
5PCElr5Ay0oDGCVE+39ZHOL7Oo2fuxf4PPJ0mM6vJYE/MiyRY7LEJ25k83uQGMm65thSnZaJf/AD
Ddj5trU9Ashvk+9plT11UGY+owzIpvf075q3zB/SMyL8iS62GeJYDGWW7Kl4E0431oo+a6dSHMTu
AVqTosVq+fzT74/I+Ibl9njyxfaQVqOWfcPgxe863b9qNIZU8BJIk8EHIFMFXDW+V9R3iQ4yZziF
iGLuWEl54H9KyMtLndPRzX2fY55yRcHSR0i3A+2ByG9e1L542SjpZkSN1gqgzjrv4Iccy1HBXCkb
UkCu79bZvylQbQbgZGxDDIo8OZByqPTCBzulOI7xJc/snaNfeGvPOKNWIQTA+tMM4oUJn39ijQ8k
vwQni9QqiianLZPT/zNYS90AmlbJJ8x1eC9is5Y5JH5U0+YUv+hWMqAaQXBACAEvU+UarpEKn3nT
8DTU2SDkUfouUzUuqjuyKyAvULqwkaOi0ME0HbeK1SziazfMMtHOCMw2tK0gaB+RyWtAWNKxd/7a
kUrTkhYj2Lj5+X1LPsk1tw7c2dJZJcASXBTXGCBg1DhJdia1gcF1sH3g2FwIAgAmsCcoDZUrWEBb
Da+RDzZ+TraPgMCHromCkBLJI/TLb56F7c/0bjJWA3ks36IqV3Cg6/FczPT7eiIlTJRFDTX5uLIl
wwzlhdQ3FCpP/1RPQx+io9I9vFQI7Fgg0bDbUcX5Meo7U7QSn4Dt+I+3PxHFFfSSUOix93R93S+C
bCLaEW++8mMQ3iUKnN/D6DtptcBCIlfqu5jcRhCshWODX6xDsDb1F/3ePjOpndg5lkMQTl5vRJyQ
Rwe2I2pEcVu+VR/xQE/biNOzY/BUixLPv+Oop8geSBgxnWcHUGnKjw+zqgvLah6/KqJwn2pVkZ1E
giFyO4H4VJW+nYEXkeNLqU6TKt8rkpVCor5zdeSJZmc7NonZParnhJgAWJ7HFMm3nGxs9LSPBKFs
RDzGmifpc9LjS334SnmnmZry96N8qGiqnu6plm8OHWX36j+XQZVE87Lo5MPxLWNRvJ5S29okO+pO
qwikdEkt9U6QSGNoquN4Ob22GSAys53pyJTgNDqaAcsWgvwwha2hSt68inFvmiuMLz3WseoiNRca
aysSnjKgZgLBsqg3F6ngYxwQd2MrbhxbEOm6nM/aB6PBjflu5s/ucCfy0vyQGV73U7HcIDjpVCNf
V757B0j3gO5c6B+PY0+nthxI1zpt2BoPjdRJUOw1kSfJaO5zallXXhidZ9wKsWDFyY6FiyyLW9f7
Q79MFNqZ279dILZ85+RC0ewAk5oczfr1E8Soy2e7FAxdUJR1nkMmnUSrR1x5JfPKIJF5fi1Z46VP
JUI8AHsPwnUNB8US8Ztv3M3qB2KFYHBMYJA6lS7mv91JJEG9jQ5UFKgpdQfTI1iXIQHXuSrMNoT6
ERlt9LF3LMGAhGvavMe6x+ircwyBdj27qzSIC5RVWWwPQYKwc1zH5UrX20VwVQfp6HJ0U7A0Ce4W
FLYX5flSfR2S0clRtjWZ+sms1nBNLbQGACLgZl8tHuKR3lLSye8KXd+glFl/icNoX0uY1PAFSknJ
pV3JjXVECT2QWeYrdjufAYXpfE9P6cKs4uilQytVsU5OyzbXg0L8r5PELzkDeiWB+WJMKGnRAhq4
c9RMerLiUV2n2bxUldHAAuOldPuzBHhaGC4J1MDBlxjMoyLt7xQgXlaJcArFv8JKVY+tIA1xjoGC
BvBTOY7vvo3xyrpI/BmOQX/Ma4+XznxSh2k9O/PD7lfDLo7E2RvwDAZD/v4UzNxP1u3dC3I/JbG/
qCdz1VM4qggqVPr7wEeYLQSbMQBqEMfzpfBb1pm2AT86tcV8gq79Oay+jk48PPb6VoxhVpJDw0FM
tKakHhzN+HsByukFOk/zmI9VlHtVrEXDuc0nSMBlRHLikjJz4OgTjilnEEHGNGH/GE1EGeTZkAY4
fOJmHHGYzj7LySKNrsyqxQEa/R2vnyycMKkv3VkgMA2vNRZ7Y0nZpoHMpOidOVPbNi1t9JO9XtWB
xMzJT6ntB/FZRidMWbCD8mDYUo2ZoPyB7qlNuYaSPQYE0OXkahoxXhaYkc9nMgiceWvwaUEQ2UIA
nUvM0KuqB3Khsjh9Hd3H2v9D2pq9DluiE+xpK8zk6AhQJv39DpELno1C5ZbKY8rhO400PIiiDz9C
KEOX2zOA2G7u6vOERqC3HAxuI1y3u4xVuPeh2xxmd6I/e+TY0F2vRpGgLuNr84snys4g5fPzpn/+
s6z9njJ3gBAkTnBZzOY0SYZa3TVpAlYtNsWVrYUufc8VNv1ujiLCd5he/HRPcx6/+PG0p2NLJX7g
TdbmcUtmQpAzYMyMytWAvRzxuA6jXCLEXYEQzLLe1ujaZi7adURMTK7X3FUc/aytmjh2gLHP3lsI
aQay+oVrEi4PTl+4YIgEOA3DZhh05n7ULSvO2VOh5Qj0fbMh9e1SCZh/gRJgdYTO3rbzhM4BAlfe
ThfxQlNfdXhWZTW9qTv1/CIfgYWxmovDJi8NkeybrtaJuqmywOGk/Z2q9o0SabjkqSGAAYygCPhM
AF+HEGAplEasqVGh+rwajxHMfTuR3rhC6SOdas6TyZQtDXSQA8vsEo2cWQR5KmxcI2mITtK8eSNZ
z/hBbIvwfLeG8n9jqdxPmuFWD2w6km4Mqlk4LX7AgGyVfzNLybPP+b5/sAGKxCEbUxd6uVbnilEp
QvFQ0/k5cyNA9wT7WYXyp1+jdlsjrhJhRnttZLeSo5qT/W3EGeTGJgbfDXtqo2S4aGOqZ1IuNx4/
dX23iCJoozgP/SYba805Wj7aWb/f3vOlnCIDS+pz+BxK4iJFH8rfZa04jTpPct9DKuiAiAUX1lWO
O+GfKTdmIGRc6gO9fMFEi9VaxmuXO3Mb4F1EUEMMiupNKoZIn1wpCGNh60tD3WkmyQwOBHMh8lYv
sJKcG/RL0wHOBENX4XSkHJthodtva855Agg2JNUHNXJHa0ZD04Vnqgbm6bEJoVK+RW96OPqvETf6
l/oMHqgWQcQp9NPxiVXlYhxYAbv/UizllrRvFvHR5j1bH6b5jybmFXE2Q7Rmk4y2w2G9e7scS0N4
LsZfMjopZKhJCpcxtKlA9TQetus66TqZkXqJ0Hhc/RWJrtHcixDOA9HwED8i+CA/QOG6FYr8Byqb
Nh2xMtHtxVhyWFaLEH1jD8+I0EBBVEKF8KuWe1Vqj3q3iRHGE6lC99MuSV6SkIg9xnvHlgGM3/8x
GMgx+pEuHS7j75j8OyV+hoVHY47wWc5E1K8y8bfsYOaTCMauTdFC2ILJHkX8i47K5y+M4hBizKAU
BHJ3qpXXi+fzhSi56ejn1WTNgPI1ot/hOHsNglOFiqCCmEvmJEcKxxVAU5i0Xj8xJ2LdWDKqco/P
o+SmM0lvj1RqpRNs+lpepfaJ2PObwvopsCeGALBdrPAckD/D/mvs4jYmBb9b/0DCSj/pphfYlNc3
pUydZuKcjzmwAKdLmg8elYuo48oZQYt2AFUFyFoAYDBiZMAlYU+YrniwQXORBb8AA8R5+8LI//QY
YGMvAaFJmVDybJ+CUKn1DUmaJl+FX8VdZ7PiCLKt5MncQcbzG1ufdQRt3xeIzvUU1SVA5uN7Cm4N
GhZ/1tYRvwsnEBRWmrx7EAd2ysB3NEa1B14DfBZxx+gZGera2YfVm3Kh7aadvW3Pi+Fs10RV4G3D
W0SZ7n0bcMaUlnP40TtwfxKUQedaBx5xoFgkdZ5FrTfjtNia21UJiOJrof/3BmTC7H9eXuJ+NOet
1R+hlCE1qlsOI4Yhz3AV/x2hHq/1Yp/O9GqSZi4C2nEn6lYxmC+0F7gj5sEX6ANv3RgRFOo33KJR
3yru2fVgl8R+IwXNxXxbNqFbHFULMY/Xw/P2K4A/njGlNyqN/zqWkrKDHpCjQfj8dQVB40QN4Fo6
xwNSaTvPJI4pgGPwJ9oedYt5v6F/WABn53bQ2TSCLE5JMOnuYlGnZxVx5XNkAUSGn3txPgTxLhm7
syF1QdyAYdk3LpqJh33pQ9/qJza4FHW0LoabdmOHR87h6Q9RIcz+24Yy+cz9iCwEBjYYOb3zHZZp
CKRijlfzkS0KCFKOAgGqgzqUy2X4WaRYWl60uSAU4ugb2EI7CmO904xycOUWS+2xD54irZ883HjM
st8FVICGXydt/wc33Hyn5dxha/6pa8GQI8PlqHU8fKMIMKZO/jydlKvb2NMDp0oJh2gCRTLcjpZ0
6UmqT7c0tiaV3XiL16cMppsVGK/rvg+UmO5diiaf6cYNKvhjdJYbng30crvkkOA4yvYKDmwLDGoz
q8Qh2ubmTlAKTt+X0TPeSMA1wHg//HYYeLS2q7zUJcLf06wfAb/F+tz0gebrBFdlRPnNT4iC5sfk
6oNRZYG6AvAVP0E30a/xqFGpP+xrNi8JKhideBFXUrGE++ClulT0GMbAz0297npf6l/gebOOcaOC
JSlUjyoMctS+QjXSEPIxm0y7/XW+FqMGdhi/AHcgDX2kr9SmChntAbmSpM/osfuM6LkB/w8nIcHg
w8rvtkzJSqgORhbfd6ACN4dbXXv4uIksKzt/NNAw6JtXw7ge8gc2q6Awtk/w16otso5duXRY0wIc
9ednw0Vh7F9FXYcACuHwK5NF0t9XHyLWFH4rIQY3HdKJHvcYOH2XqXP0Gqc9o6LxiGKcvqYXygce
PfCpDuF9hQ7gs9a7ma/XWAWq5f3na3mGtioxYlm6wUsyqBxu9AAmTHTWk8vy6oxRrzu+Xz2UzhDz
K8IIV66qTPGEm1aWtpUKuJtlqjh4m/INDzMDT+AiMWT9zEt1jevKjtcqvzSicfvhb/YnLbp5YhcL
y5XWR3YeU0rOrL13HVqAYP8VNO3CjQcU1HM3QcercqOeX8PvRi+xP+KAEkgsGSNIrJR9sNw4hgaH
4bMGkdEzqv8XB2ZZsoJ2REMbkaa6zxc4u1Q1qt6DAGbxN9eKUaR6QiRK4IMpSDBhxH58rKp7V4jc
pXsAN+XnXWNU4jWzPraVInpnCgRlc4CurAL6aHJslydHlRAHWGGKgG+BiOD86umbqyTdkEu/ZeZb
+x0FxXFBxYmB1cCspnbM2OhLWbs7TwTRSr694W0J34xn2mcittiIlNHWX+Wz43kmZEy5+0UsHhu0
GRFoxJui+mK1pE8lEcPZsEQw/J+yxLybUmpYJxQjxx00aq0eWuxNenCBLcLuP85fApGhYWSXB/Vf
4uaxusmvQ4XWAJfuRHIfVUnepMzuZ6WDGu7SNDKAe5X7UHwUuhN62jpM/QS2IuRCbFPyUZtqDrNv
6IlwjqnDP0V98BmHh7Hy/1zel9J5NGz410tqNW7xsuMrtUmIuf4fPvAiHyKuNRELl9MFZRpuM6Hi
XuGLDZQ/z99wqR1SJkGWBf1/6EzbIYOUN9ib/YpR6UgdSdhX9MPk5xxt7LpAq6XzBeyDMGUbFaNY
1f0Nv0jzt00/i9i5dH/aAioEYinQseUFuua8A3fRl5z9BNMaVSYfyLEn1YBH026QNgCLuG6FJgPv
/Uq8NrYq1LkVt7jBYximNZe+mo0T3wtrUA/7kgue1tWZp6i6h/dltvm/A3e+GuE4htkwsYmOSBt8
Em8oo9ahDkgt2v/h29lIT84FhJgCKbwFP9N8/b6Yd/5xjR6DHZJcjbvU1FJ4+oWDsBTwbZHCU5I2
yhCWhRNfgIrYbp17DbfgOUYRoHavQnjwMy82L5hBNIAliYwfrpmDMVO3AKHO7cRZmCrbwri0r+Ip
yc2F+dPw/G9DKTxyIXnHwtGWU/vOHYX8J52hxKrsQBfTc/fQ3aVYArn91SSgFtDSOUpNuhG0UGXH
pVrnyLgKZMQcyU5ncxBuZic9+Szt0dtMIX4CN1dWACxcALHDKzRZhkQF5/di5+INKJjHbnBzFxx7
uZGXJQ0c0e6TqMryQKe7AHKjof+1eybswbyDKOHfgu8w3/odUf8Uh85e2vBSnrUVbcNwAJAqz0Ld
1Q0pq+IDjMTXZlw6n9O4ba0c2qhpxofTYrHrh5XREiru1zhp6ZGb+TJuHmXD16GhcD174oVcSNkP
/WNzgTDUg8GZDqfNe6EccHLBkHTwRRMCXK2eDpRYhVlZUykwDX3Q2eIGIzaCXflkdCzZ1Fug37Uw
IN6Q7KZCotE5w/xsxi8NjQ8pCf5azNl9HtU6CNaQy75PXY20Sf5lj9cNdmDlnFz7jDsZgWyhuq1v
RxrL8sz0DK5eMrIPGDFbXdSlfS36OXTbZyJC+np8nlAoVBZbN4DIXyYvKM+CYxj/iWqypkY8Ywme
I6zhQQcD2/XQ/UwgQ4pobew+H58zR9673c9IsI+XT6JM7BfB++naABhCE7PiP/BZxElPvIXuyQgI
KVb8fBiRwazDrzSE+m/u4iuDL8RHtDCeeYJXpcByd3BsZ1MwdaqTIBhy9JOGAL167mE32bO+jDvA
BDzWyuAic36ykVeu8xWvzkZaLYD7ZM/536ddwIbwL+6mJ+3YUkZ8rvnPW5RlH9mDWWoA5UcXeqwh
mU1ojh7sY6KNMJmeMDPE0vlVvfFi0+YU3b6KBe5zTQwq7Ibw1daaO11M4nCFkwjjY8JA7TTDjcV4
0jjZ111apWA42g8Jjnn65+PN7Cuz6JIULqOPFRvoL9ZakdW6Z3xMOAd7LbvQGfYc2aIeJNou1oCu
gi7l7TSn4oGeLRDDNIedexaHoxb2xSHESmKc4/TwpO5HBmrXYeefCdlNT9R94K+pyLYv0jRtHU1Z
V+hw3iO0MsyII6fciU5SUAmxKu/hNszVCGK6USreYjM63Jc2d2O097g1OCi4O/zlePSK0tyclmX1
rUbDsI7BZhp+zXOHsF1cqYSJZqvVk+KPc1bty6BnJIRvQd85E1ln4jU3nXPcgz7JG2ud5JOaen0B
FsnWWKj5j0nVHVTec8EDCEGj0U/4nM5BJPgGb4Mo2WgvuPhMLWRfQLAoEgB8Lh+7ZjiwnKVipsao
7Smh3CFd3fv5VflPEst/bJka0oR6pePDQ7EiMUoMpNya8l4XRfvlWL7xEBqmLkADam4069W1Ouf1
oE8aXN91Cnwca84jNNwbGCwvs6Wb0zAkekktyb5Vorcqs9QEP6mKjzqvPRBUTWBodxU0yp343gjg
gtLq2BVBoHy/RQscIX0w8awlZAVdh9xd5VeXpClVk0qpfvP/UZSfPTMggPqrx+a/tl5b5NMYkolx
mmatwtXDgOuh8p7J15T5hpPE79IAoNDWGHv5/rmLc9KdHji3415HEPd/kug7L/GAsvvH6zBIPRKT
UvHeUCVpn34lWBzbtuTOArxiJy7++Mh7hZuk0rAWSHbq6nOeBNBHMwDuERGS63MGwg75WIGCjPSt
lwm5YiINgWRqMht91BnjasguMch3AL6WaDtVZ1k0y/kzoc94PWg+p+lxca4QSdzbTxO0hdG1oc7K
5tGTHlEYzVxDSeWqFxnMeKPducIpNYzBOvkVcKwF+Qqwrk/XYMX6dKDyvQd8F6qlUSD/7O8hHQqs
vsNwcZLLz2Uz2jAAzBgiqvZ3MZ6QT6296xQ+/9j3RlSO+4ZZ/2BBnEvpPsMmHy0Az51NwVq1oECD
UeM3ZeBqUYK6VunkAAGbMzES32fsigZAnialX86WfADSsUiS20YSr/j+hh+WvN8lwpDBHx61hOMe
ifoC2cKxGS5wX8GDKXcr6ESR6fwDbqK+ff7H3MD/j11KLPGdcVqezxYaUlAG0LIgtJIkfpLX6PgM
dF2Vw+aZP1dDkGjSZ6Z0myvE24MhiqBe8zO6mmZeG974l2S5akwlHjg4vubLuRF+TuH+7utiUNxi
Kiamz0cTssehLeqR46aBtEJgX3wJMW0VTMV6diSBitoa7gM1tIfxFgKUJ8Zh3kpP7vnip9MXIKb/
oZxii8UmsfhIFoAdnDQ+eqWvYdZ3y0W/xu2DmDm6eQDLtx/SuHdq8QOW+cnyqo4gluTWT7INCtdO
ta2KcBKduwQeIkT0/JSkcI97tckUiLhULaGBZg9sOcvyATXBsCZ4dFvuj3mwEz5OEfyuxrDJOxib
EJykmnE55t4mvskyjW6GC+e/GV/gWGVkx8XaYf6ivCY/EK3MJi443WktNN4e1f99eS9pvT9WKk1M
gaNUxj82Vqy8V8lv4tlcekugWQzXxj00THuyqW+8pKg7QKrkEFw+HvkfCDuhiggWY8Pe899tvXlI
U/bBfPfu+E04qCmGoBxC5nYX+/3nFUe8ikGyvJQL3xPOVc9DsjtSXCChsTqgV64ypwumgB5eiuis
jwvdT3W5oUiR7CQ+8DEQqJBmIKEZDSDnto1uvbxOxZQfQgnAHw/0QVx9N2/OkR6WOHBB3QN85YOY
bE4TCtAcm3F/9hey+vc54Jc8nDU+IjXUk3eebU405sK2uzLq9w==
`protect end_protected

