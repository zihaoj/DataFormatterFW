

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gFPxhRrTYv6VaHVPGAiPVy2YZ6S6v5BzuhWPBzwrubAT6kReucnryQjohV6YcQAEW8yJvtBp1Ysr
C+Bb5OtwkQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZrUOXlzrvv6qQpYJjywdImSGK6eXCI+MVQlcEaIaqP1/0j88qHcz2caBn7ko88g8r0vYZDYOxV5n
bwj9ewbJDQQ9ap8inJ+mdTFTKMPo94XSVrTA1cg28DUpjvYCwKrTbA1ADYh7RUYFbkkhMydUo7LD
lH1Uea4TZeH7p9fvCAc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KbcSBrdjT+GWw7UD28rW1gOX3CWu2vBfC5H9w+FelX3uG1bnT8AS52Y+stg85peQ62PdcFUi3fwK
NXs462r/hLo1nXD5F7+p11ru4OTbASkxrndcH0xh437UXtMIGNy4kESqx3cwYEQPIPbRIRHzo9lQ
H9EeuRfgapMIwrwKfCXh5gP57kN6zZB6sonyIx1xDfWBlHzocSUfgxGgT8hjIANluSQYpSfuUlo+
dEI3dEYoep/bAM20bt7RM5pEkOJajAoAtlMCTYREM5sI9ThqVmwHm0PxWocsdrpPEQovhMXL8bOt
27757RGtc969a11Cl9CQkDFdiqII0115hijMGw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PdZa1nRU9Vl9CFvj4B3l+BUQbX3f5MtNMaAyCvHevFovH8IDhuKgsO//TZN/V6VMR5YKx88nRmJO
9ayU3n6NN6JGyQ3D58SFXa1a3OL55wVnztwe1sdhcybNUAinICFBWGz/HG3ewmeUDTJCH6F9JROD
zSKXdw3fVdzQHjJ8CBI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RFmPg+ESJU/XzKxI7CxC31/2b9ui3jWsU5VwZ0xzon7uYu+V6+oXRkduShPEbf95d7/36KCCl42c
DIZ4bKmOA7sL2G1GDfX2uAXELrSU6RP0dLua5f4h4uJ51pxMoZ71Og0jK8qBTgKG5/XNcTiuzcSx
J7dExt5Zvipm6MezAEpMNhoncMZMfeEsTHfNvBWH6oe73a+ylanQijwvhLoY7BQzeOBhwqx8DnjM
9rOxboLIf08CAVrJMdT5yb+t4+XQyBrBTrAmlnTZ5Wd7nODE0b5llIj/BG+v00hD030OPT1HhKY8
8XcBy0JYRhwIxcQi6EWvXDTos47nlnr5S4eXhw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25312)
`protect data_block
m36LAfS+x7yF9fpyZsEiNJah0kSyOesfkrY0CCCRDOhPilnWXsVcuTxGWQ17LahCLJORG/UoXbzd
H2tbPiW2ORJCYrSKX2Cn5HYPm6bCxoK92qW2EN/bKje1MwAgLYwe8MnlAb7IdKHwPn6c6GBBklpe
Pjp5KghVIyeTIktQvCB/jJjp4xp4FU6wtor5uzUnRLilryQRqLWfSs4owBOKn0Yo1C7E28CR3Udu
UWDNzDFoXhvxGpMVsFx5n4SWK05bqxZxkdJRLnYy748IFwR0r3O187pQ/+VEWcIlzMSpP7pe6wMl
GEQxEwEP57y2377ulwXbaJCZKLfUKhVIyQL1SZgqIVpczWgY7QQaxwh27Saya09BhuLnh0w2AbF7
Z72O+Y7pQcOMjXUuDaQOXRZ0iLe0Be8H+8xA5UWR0ZHRAixeuVgLLbya4rchKHn9UX8K2MwJ4pa2
J9VcgLmH1UYj0oSF6oml9jfWsDsSJTOo3HKbiIiEXWXh+HA72cqzwTETEp0+yTP3ZwH9dtaww9Pc
34snJq74F4VDSf5aeRr9HIKv47FP2ZSRX00oTq/1jtiKDvFdlblhuPCYkljiJ3jHzSRdwBHusb3Q
tcu+gEYEbH2PmRcfBevXo03Dv44XVe+vOim5JVpSSgt4NDFCHlc7m7FF8mJF97d0Q7FIgLd2ogx1
CTOQHrRBjK5oe6af2Yj90ulZFsM0Z6Xe2i8K31vsbEpzJr4S6xa+XFCnBIZO8cTNHsD/BgqCwbY/
IfaCajYOtgm36ROKxqzWie19Ytic3JOEPB4UftxUzW/NWMFlT+LutZf8pT00BNkrZtpiC0K50v0C
3jUNEHH3MStMyCwNa3Z4gm+6NM7rTM/AHkqow0X+KF8rtxG3cJAOwQ0DxDNI/If8I/B2YZcKEdiF
pM/DQTIXTq4ECWAvVt+qAl+hWMgIN9YNw9jySj1H6/PEBkqlcR1YFLsKbH49CAkaTS01EoXYl5eF
oZmcTSV/RSG7hqUtKAJsKAm5uYXI6qF/mj3WBj2ZG8Wx0w8wKQ2QrbgzstqyVXMB+nXqUaHWGZeN
UAgiyzw+iocVJKLfh9SZ8dNyWA3fn4JPdpB9V6h+r5YGk5Wz4dQxUArNtEVhYfFBQUPcqJPqj58i
p3WRkWOI90DYcvP2OoBqWki7vMyFV3eyu2D3dAX0k7l6ywEk4DJxwcxM1m3Nrk4kbk7G0Zv7g9C7
cB//uFxSGQTpZxGWGgpKiPG/MG545FTlly3EjQWmNdS0qZsjhx3edTD4Fl08Q8Km9y9q3j4WoQCV
GrE4PhKQRaH2wtpTubwObpis4LbYgTBx6pQnYJwbqU8iMOjEHX2wl+tMVMT48lU36QIy7zZloylO
rzzk9/uQ4+3kMnLUMOUawiCNg7yVZ4TKj/e9wNBxsptQmV6zT9hdkvUDgtvUYIAlRpWJtamUEezW
CXR6lf5WRH3p1kB4OcTrtl68aCwtTjwAnneNkXEu/di9Hpw60KJGpj8Lnoe9g3bkVExDBq+m79tk
yuZrIGbK9+WdcKkXeeuKcgxYpoxscrLaDhgPfC9yxnVxJ2Zq/hQK+5rNoOIngGtdb+Whvz9Jbhfb
q4EinlaBWMJQp/sQmKHyRMc59MNbgtJV8NQ8xA4MptTSKfJI3xNoCMxUNQ3hM+hSpSJscXV5muaB
MGDvHx3lkKWJPp260J6PmCgEhai9eE4JEGAYJpaZkyL7ftSrky3XJa5M5zHGd5f60aeDs9QC/ANT
dIdOTmPN3n0b+i/eohB2I12kCKApXYAZj9LR4iER/yXc9Z7SDgyNeP+KZAK/eRgOCXopzahkxctJ
VJHEYUgL6IizznVrrzmH/gYfEoNM53rSY0LJp5e0OE3sfNyzT36DpF8KFvztSdtvrrNW1UI4whUd
8bvvXPNaYcranYgpNTGl5CmUJQKIhdnz3uT4A/fYPPbVGS4RCtOFsFf6sEX+i0vpru5tnPWfeVns
UvpyFfBtO5NnI8jUGGf3Ai+MgS+XqrXcnlBycVT4WZ4o5KFbLOo1n86yZT25Dge79QSDVW7U3ZJw
oPL4IXMTbjoiXk+ELEhj6tERJEuFxkwSVKC5e7Wf7sa5OVXllyAJeShMTFxYGy3MzXbMvwXwdwPp
hJ6o1L4A42lx4o+di0Fcy7cFEkrYV+yGem1ZN5WFubHpWXzO49ezao+MKw4DvGodxefc3WK/4utN
Ymp6780TC12X93aNi3hKJurqw89jANKqsyK+GOzPF9F2PMMIIycRc/CnuPhcm3sf9FTvrk7rQjI6
YOsZbU6bmijcqxcpraf65z1zS+LdyiToT8SSMtbb5/lRC6N3s40pdFCllMhIDBz9vPDR1WUGMCGK
PZHSLJ92VpH3HJC1xDllPl4xz/PKQ4glyuRvrxocnoUCnLVW+P5kjtaCqtbiOlWyDNjPJ7MwS5bX
rac5qJVjej0nw/ij4F5uVBvHt3ccg5Rgb9jA1/gC2gwoUXOvghOJtO0gmy858BedNZN7ZGgeLDxt
AqEtHTNme4e0gyXTC7UnjCeFmrbNLpqg8WNNUGVQbbxe0shgVZkArBHRqSY2EwUJH4UrbwarU01U
Xfe30oItpyBcdM1ZqDCGGDL+7ZMSd1Xj7zEKU/3G4PhiFniRORs7XKKLUJ5OX+K+A+SQ0BowPJeV
9Wl89w6jHaEgGKcllYdDIv1pPBWOfLDpGg7nptPvQqp18tWxMY1m7plvWmBjTjGQD3tEJ/v6xAie
QCk3WFe6cGCkzLCplne0efHVycF3GUph/d+JBhvDnO9DxHynx6zB68j1CaRcKhPlfe71Ttn3VzjL
WZU6CvGvVEn/muVLlhn0wYug6J2W3Ut1LxWdSWLcuxfeKZTp4s8+FEEygEz39XY2OrqNkQVmsuAx
87wyg8cFtT05xXrh3etQp92SFVa7VBRzOIEGk7MiEiFO0PP6FteYOFQepCYOzII+8hR1MFHkQyVn
gyRLMMzg+pk9+074jxlCxwbL3cLlAxrsGFFr0nQp3t1NTIUjP3E1iAkKM+v98yUP7360vuYvpxfN
8eqqA83Fb/hOps2z6/kF5k+XIcY+aGOX4BkZxrhm/UATP0DVnb0KZI2JC3CvNT2YtFY7ZwPd54px
P1uPBLCZdcD8XWPkVxZLQwx1JVjPAsRLB2BC9pLjlynbcnl4IOH4/uZj7hD6gJEO9hdUa4Kc4so2
YBJgiqMRtZn+EYtt5AVCIG+gT/hrco5HkKZ4bQU7c0AND9ljDoH3qc4GhcOdgszyqGr8dAYU9EP0
ZqL70m79Nk1JzCn4B9dM39lkaJLZ1OQM/8puk9RqWXTn2pG8dTQxGZJCDbS3LEGKrHr6DvnqbJiA
yo6SaHUbAIy7yyhVXQvLU5A4Jl+VfC75TrGCtsk9aiB1qI1rkmDEj4VjFbdp7JZ6gZBRs8f7F6h4
FWCrXwI5/CAqFcDvdHb9+auiv3s1wW2LZGvXKiLRhGLftKPhK/tg8NeC6mzRaWkKWVHG4ohk9Scm
+d6MK3qFFRVJiiKzQ7VxhEmu4P8+CLi1eeayAm8mE9l8WkBzuZZRzpuukuiT/z1IklkEKcQlTRed
OBe8yFuLxnTX//H/bgq1Etih79WH6olUNOcZTy39D425nVYgzLFGqjqYJQ5nHlydF8VeXwiTaml9
5eSopF6X4yns5yi57aHoQ4SWftcvvt+DaDGVIT0ySGTH8vjPOELTrp4MnGMaYfbKv4Y1neTEA+94
iiokteTdmAC5RwTif1nR3hbk6CgirqwQpBQiJgYau+Iqm/oiZPh/tF9CenafWOBnGwTYkyyQtOm7
xO0CrPCR8UX6tOmGkEalN5RwY9gJd5eFIyT6rxwIuE5YK4DbKq8j3yf81ESMmvp2J3wMszcNmHgj
bqoG1x/f+9AMIwTTZO8OaJ5kVmSCNDeRT+f6c2FsjD5etBtCd6KtCn4Mx4PvZ1+p5QBYttb2bwGT
tMPsB225R8PmjG24UB89eBF6OESjQmUd4LdQM3AuYsTOTsq2PBXUc/hX2Yjoephr1QG8p/BFsFyr
+iNozuNdUCKLgumL8uEl6f8bcFaLlP+FTT/4eG0PeuDWnTN8LNRvr2UDKEYKTGPSGDH6V7jkcoH5
erlVvJ2Rvw4aX6k2PkbomaWzKevrZxPmv6768fggQh/b4VitWSu3zLEOdDJs6Gn5JvUJvEOMNcf/
psbliKaShFi3HcqyOpssnQIXjZBSWtExoVfoW95fWhmF7o3DzU54rAOdeYhTmtX+An0mBnTcfqCY
bTuPuJfflArYYhNZ0uFkbr/iH8JfkKEeLXbdv1rnAlN15Qb2+Lz4IIPI4fJ+oO9peJba111BTQII
Ewqeha8Eaj/zNR1TbrXuHFAFD54lDq4/U0ITDSJ2UxYOrxA/crMtuRwaRnoJQStwQhympNF5sPYD
P+s1j0Lb3P8QwpKDY5+ZHpkOU8H6ntZrnm+fQIu4tEuJygiBXQSoxMe3iL6oBUoR/9y0RiDeqG0D
FDkBGTyMgYdz6hesC0iGpcgI51bY31noW8B9uYD5L6pB3tYEw6DwvUlFLveWShYgVy6FsTtd06Wo
6OkJXNzIpGE9BmWPhDpK2wAZZUmA5iaTBec2jGET+qu8OYwp198v5mqS0Z36dE6bYJpknSUNtr4u
t7VtIgsqFUuJXM3YVB2tUnd1ZCa2iyShkWZyKpfNx9SQVk0Rvu294r93zHuRsk14wEVzbt+5ean4
8zFKGUNWHF1WJZLUZBGGiYKNCMgwpLYF2B5glR/FYjdzemePeV6OfiM4mi3Emmb5J+I7iSsBlfds
N5q0/eA+8IgTMWzbkOHMQdXodYARLZz6y3lOH9MUdnYFnZPsP4YLkdFZvp5TBDX5OFwpHRTLAmxj
u7dx2So+8zigvHiO3CLsxx7uOVgHSjYU2VGcgh7JDyvsyON+ZCJJq0m8balxUmW0i4jPHch/9EPa
7jWskbgRDmEiem1gdiJf5/AKFDUX6UzjrCub3Qpopy4jZYcSWqa4MKkcZZuBPNzxVUpVNJJjXcBW
cWE/OlzXdADn9DQYCMAqs2KaEAuMB92gMI/8NG/lchT4cpZrzRzf84lgedFHLUNC8/Z9rPmgSgAA
BnBLr1pMx4jN9kDbSahs3AB+HHfpLOZrLLz87AP9h0v+dBng4np+aDX4FPAA89GYYJCMD7+VTowD
LWemdAFpxrGye8d9zO+vj5m6ODwFHkgGupG+txkYgy/26c2UDLkKqWeuQLUexaiXqIAwWOR2qVoi
Emxk5zz4fqNmMVc8DamAcEEg/Iuce+jGF3GhtJpgVvwWUCBMYM9KMqmC5sJeq+yVBnZNH+SyzcuJ
VB/3GFUS4BM2LJTV/9x07B1dyUgmb1jbLLvprHSdEUk6OjJ17YgThaIdHpXl7mF4i1OC4SOBqPC3
aXDlcUbLxYWxqUIlQVdMwToED+lPTD3Ui7r7EhFLeS0j2jjCjeVIy00USM178pdlmNw2NcArbpfz
XKjSJ9Lz1QUW7Ninv+HyFGGkpi44S6oZgI5vu2Ke9YitIhz/ftvU413+HB2R+ZwJaZ5QdtKI3+gU
poruUPEDhXaJuNCjqUsStO7J+iUm7SYNKCarStfU4VltWc1k/fdUW401/nPNk1CVqKTIRIsQXMf7
bHvzmFNaKxduyAL5HtVU+hzwpXzMVwMCCfq39kLOiZJrvN2LnROsBKqdlXxhwtbeLjJuvrnvcXKM
UEfldC5pCEdGn02Ig7Wp4jw03xMJk9PD7a4p6ny36GJmqMna9gDzfPGOJYXvdUY/zBUDIzN/vR32
fovFSWHhizI1mhJGX4w0j0s0uqJq4A7JC7rqNCMkCVcl2Z75UNlRFC6g7KYoz2tKDG21DJfuoQjc
UCCHJR5PyCgDQT8PxmdgqA6S14xTYrI8AQ3Rl8F3kGuTtdsJunamAbwv0/j5qquxcJFZO6L2czzp
GRcneN2eqYNz4LJQDfTeczaH+BR/CqBEYWkAW/GYbQ91eGpFLhvEY4pSmFyeIHBC0o8L2/8w4SUJ
wVMtvJd47ojkkliyPcjTgTaQNrOPZ/8+iidZR8mCqE1AIT7ZjaXPUGjVMu52Qoo5z2wFPG16xT6h
/iCLRL8FFTWy8XNuiAe6mIZvwgPDvP6QHnxkQ6Ehx4lTzr2b459uzf6uqDsNKudzlbVArDMeyOmW
p8kwWdG+2OlWbYR1dPrYjBQ4gv/psJ0YBFykkvSLlS2chhs9gwpAeOwdcUo27OH1pa9BQPMP6oBX
QdATf7eulyRJvUbb5k+65zJ8ejXQUAimMaf3OwcpCrx39m9i3zupJx46CRv8r/fYAkRVDvQvWbpx
kLwxbgFHCLB//xbD1odDchW5/dYFqnMIuLPvhIMjvl359/8X6c5IA/4hK4PTIbp62C4iAMYPJcS5
CKQeFiA3cv0bhp0BK/Cfsjr2Q7aeVBs3jfP1r30Kyk2h9KZHk55yN5GEFaF+CbstyNnmqUajTotA
BUYfcfqJ0F4Eytl0JBlf9ZEgtPyEro0+b51uiCDHybDjQPDoKARR30HQvjBnDrMGpi//q2Dz+vs7
vWChbZzDoiFxLeaRfudQcy+kOzS4IHxfZ573VJwD2Vlr7BgCzispsC905Yv4KB0I2WuGG64j/LhU
RdgtiQIEAuMR4J4P9vEZBkd8v4KnoEtNxlG9vVFWzBJyvGaW6fy7/xgsQUfQZLsrDfpH6RyTLpQD
2VAEKNzjqvth/V73/fIBRAjxpik7Qa0yanVU1L1soShyR1yAzC2L/WZAye+kzJCjTtsFJDy5W/B6
3LuKPMm44TCKvZG9+rKOMoCtj8w7bSwuIqOh8tKPF8EL+21uVlunZHaVdPjyD/PpzushQD7yQ1V2
SuOaVVI1rTljrpiGW254UGe6GQX2zOS/Y/BfdIpE1q3ku/Oi4VTa1lGgFzQi4Tlyo2bnag06r3d7
fmTD1divyxUFROJdwvBRhgUJ6TFStyDow5ZwtP1ijGLucnWW9XnWm1kRUqs0BEeJ3bhgkODgLx2X
pvIlS1YPyaCyDeGfeCSjA5XhIsOPVQoqqZaxZUpVcHyVz56NG8OXjnLhMxLQZoBzoX81cRSoFxqF
Abu6cI5H82p98gDv5+YLTNkqCIurAbTd4PMo5P5wNAbWhplql9SG+U+WEa8FzR8i3de5JBqM2g6N
k2KmdvhDCh+ezjGro3fvkuFXRMFbGT1MQNb/PrIkXSmJSA95f8xk+eMYMNQrDAeKD5Y9r1x5mWGW
uBppt4qROoMfuFiRsg4fsjeUficJVWeaRcuJSBTUvNA7UPVw51NrB6GAgXaLDyK/gA+V9Q0y3OGF
zs0NDmiWTb9P1Yc/qdqAXWjoHivy4P0doMBtcyJNbryDHZuDPw9mrlH5wMu0NwNyu6DbrKOhnyS2
l/qjt2UOm1SQHkqajYSLHJcEmOkwkFOmg0HiORk2ELO0qhyW4fUaAwj0AsITNWfGb92TrJQHk4de
5ur4NQjrI6NW21oKibmuASBzm/rPmQ1qohWQ7SJM6j7DSr5k+92v4rUojPWno4rMdRWI3IJXJPPT
ZOQqxu/3uj9E3K73Zl3EI2N78H5nC0Pp5ELOKcJFxk6/9mcmm18wdDE9OaUZFGjUSyrxcZG+bMAh
46M+u803dWl3as7p+scZWF/d74eCM177A6tEOhs0xunXhdnCUwlB4cW/0+NoilSCM0ZejfjIlceu
pvo3Mcnpxv7AMfZ0aHtq7sXvzgz+m2arnfMG+5YHjPlnKHMV7DBX0bJT6Ydvd6vKp7NR+YyNTS6x
0y3L7NYb0HG+QrzmjVwH/0sdnwvUvic9dRNlr2le6Vw6JFDsF1w3IbdyudObxRZut6vfr09Zi+gm
totHEMGLLUmqS4B+MLgRyMRXMzTd+4Ztn1LVZ+4Ym4kKcaxbhaZpAqYcAakso0U9V0O032DhMUwg
3hhJO2Wa2vq4GsP+mJ+wbwg74tSp0HYRyyaBCn0CAeA2sqCFhKDlYWciT1uaOrQqwqFfEU0x5y3b
L8OzVkqciPN/XFIV1iNTHE8tSHJ41iRHj9/MWVTVImODhiYHZoCRH/7+e38u3pWKuNEN6CKJJiw2
zjNxfOFBnQopufoVAZ5IbIhsnA6QaxPZ/Hj4aa3v88VTCh/qZ6+5cND8+zmI4s/ScLuDk6TMmDmw
x0p8kggtn17dT7KHCK6nodLeA/jcaTcHA+6f5vqz02AR4g0YOL8kOXz6rkRaGRaZA0w7m84QY1OE
6dsC6arxtM52SiuSEdsaR4xPwNB+smh2C7cli1MHl0IjwE6pY+ZrdDrdvcTuTHrUehqwpc6LQnRS
Lmrootixmfns1FIliQ8iObEl8ziBc4GSBOAnALpXEU4AuVunlxFDlhSs3nYbqrW/c3zqi2zXmUQU
0ZHPQwLvx5awiQYlYmPl9nEOYBcRL3qxtN4YlwqIP7T0yau3ZsPzrnSLHWI0Og+nRTWpWxRL1VYd
xV8LBwjyTOE2v9OXMKOIZbuR9ejsRV/FDg975btMSuTFymeAcBHDZTM0mAzfP+cZD/Y3Z12qpXbv
V7vsCjKuM8m12uGAi9HtS5pAjxQ+ra1QIKkEtrwvDU627TPAbsWHknr989ZAaAxABGpTH2N63xy1
v0fTmyki7xiS9ku+OylRebnDDxLOiC23niNUjhw8KIq58lFwPREfDYUH5F/w1c0O/HKcbcrtukZa
flfKqMnHyGCY86wo+x07jlygwXtNxMtvPE9haCRXY3UIy8X042Yh9CzwalpXnJX98q/VWBrzcreA
/5+3Co3p6XT2texuAcylXkm+z6JdbwHMvEbMjm5S3KliKxkYWCUdnkWvsY2k1N0KjmuuhTL0EaM+
LGHnEW+05Ka4iLwQqn0D5FqQmIxcbIks+LX2AQtCLIT5veDgBrG3WUpMICZ9crn5ZAl7Ftn6vaib
SZqlaz5/vLMIdhgwyDxbIIdXpDDOYA4Wqjkxf2ILyysgDk2NQyjiILpMmrcRJZVoWB410GaWpS8D
72xK1F/8JbFwAicG9/oawWpsTfCzeF46xsTKJqsGgn9lZ6FjMDjgBmstjyJ9N460FBs/9ElgVElI
BA4DX/bVHmMIUX1F75GFvmMhdE5HOIoRAXI2jRkq3k08RUFAj7l6oOL9UZxUxJks7DA9cHHEPHTa
u/rtCOZrh3EU611bIOLj+xYUVw6/5n1COMd+xcIgCwV8cd1xDPBVf1fY0lmKiPWmKB/WMpZNSkGl
rQUNQ99ld2dqtseaW8AMJc8R6jsK/kLlq0vryBYlvL2NycCIVtcsST07f3LyzT9UFbcb/ySpgcY3
wBrV1OIYYV7YJzjB7OjEQXN0PmeL7jTRKcvHoU6MKHkgcEjwJj0naI9774YilMxPcTFk+ALENAqO
K4OY6+H0FKUH/+krjqMZeccm7UG6ky0q9jP5VOpVcq8OdCnIwuajE0aPlRrqpn50NeXW2B5YNHo2
quCj8lerjg61OuxY+F/QoYoN5jX2BmIufzFrDTtBdtX/q7vu35wPwIURaqmNCc46P5uR6NRbxc6w
MEjmhD+Mxg4eR5XEbAmkz3H2n1Yj5XfPxS27VZZHvXK0Jax4b6x8kHEWAk39VjlhcUCykkdgXgCC
gSGTtaH6tfeOWuJh/vkcpRvx4p3mC4CBVVfvhpLbd0l9NTQHu3v0h02bFPY4JPQeylIFyz33PPJn
zpIIqiCXxnpkUWKCp0V1f0uteDx0BW3krzt/oVB5wdit3reuQDNZb5VC4SzQapX7wamXH6f/97Ry
9PuiK9GUwq5B/E5n6OcgrfYIb4pJCoXGl2K4f/zShbknsdhwA6J1sPuBKtTtwcDz0aArvaTvtfk3
+B9JPvYIUilvo94gZ8zZutJYKP9T8RoM90NrA9mbgRcc6GqodS7zDqTmY5ct794RLHdu0Q042lZO
FTwWq1NBp6l9Y63v1iFoZDd8Le9eObgv1onINT07ccO2yhXZhMiyI6IHJCXjMmYlaUKbfWTI80fz
0e+LEdVSx5Oxw1IWl1o8XqiDgE0fcbu4c/1yJMjCVBJuGBwomcZ3fZiQKdM7kVyxHeF0SkCS8obC
bqzGn4EoxX30JwpxTg4q1Rb1XedNrQA3d2K96kBsxPdsp/AXnymBfUKjuOWrLVAgPoFmjrdbze0W
AU31pFbFlmd2xXnFLml8DHbgajR30o0PpLoQ2evZWiRI4CF/74pInZC+SNxQYS0yg9WMo2g1K9NA
P/W+JfmDuGU2tX886CXTPLiw1AvIB9+RpZWkJUM0YXmEFM+D50k43sDnfKDLJUiYSlQdi/5Z8vPe
6JPd1yP5RMDzvZZNeXpX6s24JKiCHyYFPxKY6DvY12qBn21F+nE2UlTy43RhfokkYLcsgeR2+XS3
XnmLXwR34/4d6tBfwymZHn8KE9SVyKm4aDJUVLoWkKMys+NOPHDkqUf4pE0V32U2NEV+cpZrkks+
mqjLJx5mkWyz0DSCoY8lFiiHuJoNWa/WvKs0vgGAcmN280cNfijBWYpXF0AyJe01b+yfGTE/Zxvk
7LO99HpWSrVZiXPyoGKw4HPW99murdDDso0zVhoQ28l6g9/CnJ5b6qF8HPR+N0HHNsdP5PsfGDAs
GWqI/p6sNcD+Wm5/VL1wtu+DX/RGP5RiVgm15lOt4gpWdKUQrJ7TuWAAI05fxv8raZE4AshhqPzC
dNQkKVCf/Qh6UtaFCOZ+UsaaHeDqnbQ3GmKfAa4H6lZSsX3AHGYzqn5wdMUMnH4LC/TaCs++lxCD
3/rRx8OoZIfmHhinCkaEsvQuCWntVy3GfcrfnJa7xCdIZTxukDvxNbrzHBF8Pyt6Df/vzKH89/Kv
wznmqp3ndOYA5dzY6XQiq4c2McZ1RIeXtxSpqgKMjds8ozqkkG+pktuG9pc+7UpZkSJGAIo08Vmj
ix0g4VWYlTcgI5f+be1p/BBKEIIJssZLAFLsMAN11ukzqWHSIxmhB5uScOPhFO3TuJhs5rAuU6Up
T4YTvw54wmi10Bq9SQPcu56MhRAbOfez+aEMB/ETr6Uc6eASYULcDRBhpzl0QapNUU8z2i11B+xF
odCZjY7OfUKP5FupcxaIXaanYX7/OYdL7YVWyRlPlgEAqc2K8vgQne3QdGiabvznDU7cQOIgWLZO
I/rFwzoO29RaSuv/rKifjr7N14eo/JQYD+6FVVkMwfX+gyP9p2ATfC/sJeHfOFexpnkbyIU9GXZ3
tigRgFHn/9fue7dXPnH5Yaj5qfsiq1RWnVh36FmBG4qnc6LoWbCNw64P0QPj351MGjy2TJPWfwsf
tBqHFed5slRlCU1YO4k41uaUuBs83L3W95nyhD93PtzyPiWIWKjS/wtwfDj8ij3RDvno7EyKQM8D
+WA1Ozqe6+Vf5ftKgKgVQ6SlIPoMptXbqq2lYl0n8e2inlBpnJLAHSeG3ySpaxYEenrJFSnwU0nV
ZI3p83FwNP4xiygwwK+DmCjjPJMvOqJxtDGRYoaX4PwOV0j3l/Krymfj3sgcV3hZ6Uji5WLyv8dB
uh3WDlVkHE+CV1IttO9tnlbKMT9G/n6R04DSrmKWp5BFx+/l7hDdxvYgX7kB/eqoiAKnI+plvAQF
NTuNilvZXXPAF6iRUu6B8hz4Fmds7hvpBZgb8qCCvpkY3lorcTbeUvPhYSsLH8hgfnT+MkzvVXmg
4jmSQnkXDG/zZt5eVTNCDE+ODXTBdioQrAHPgkVRJEuAzWP2+qKjI0nwCzQdneUgh6WA235wXX8j
7JS3HE//zQ8B3Rij0l8mUJnl7zQT4hx9UafDbJ8L7aGS41gxGMEwn6wEOjAHt+DtS3ugF7jKBny/
uHk79n8dQIIq/T6s5TQ3ZxnBNtQJQv2ae7h/YiNLDOtCuLY9q5ZCXmKWMbdSnR/6JISSP3uXDTNZ
Usvde4GJnHtq1FOksXVUyS2EPEIpwdqyEBUbJO3IdzEE+NQgUgJYMc66Qyos6lO8lCEq/+uXZtL5
6QPpQEO6kiQFku5Q89b5NwJGd28NHEwFL5CObkMMaixXH7RZT1Ne/NNk+Z2her/wsOq8jQwbeAHA
vir5Q527afwbVCmupj9yEfF4qP4pcAyk/AhfVyeOOfnntKzCFsAZYShiHCCnyMVJ6RmYpB3hWdi1
LNK5aQfcF1C4te2OqL5ZmSRZRloKohltBOZQhsa88kUMgFbG49nCIv5UOdxRfBka7I8UDcp9UNgo
6k/makbVSXDvbFxbAQdtFiv+gpGyhCPwj3+H4jjISK/F7tU6Pn6sxG8y1myL2IsV+H/ZyLH/MzEF
sHt04Fkp+NCwpFndSLUQZ2fsxLlt624r9h+PHmCTR9NsznBIe+qZ6WuzSjZGLRkLigtyBOnR0J1p
nMsmX65QKl7VVGKA6l9vAkjLRRI15rOT4ZZzFw1peFaS4BOf6ftjlxpzFOTlB3h3SOpm3BPxkBDW
+gMHWqKXCbsZPr6IxNEL0xldqDFGMwKw8WfT4a5Ry36jiy/w7vARRAA5FOjHOP6ErmzhbGucBpio
wygQaVUNIZN98y2iuxwdusA+JcPNw8SjkYFP5eyup76O4hmffwzU85PeJ7safHQbXHkoE39mcQcx
+CtUa+kuh+9ApWfpF0BbjyH9D0LUnpQxZdjr0oKoopPVsqNUaR1HYjc9iEyO2KPGQoWyZXpDAqM6
ntYE5wQCdcP80hyuLEGfZFp1+DNNre8VhjZ5JA/gSpxWEfUUEL0StNIH7w3CY8xeB4cXu2XtCv1K
BJcNR09U43IPN125xc4s5ZH1PIBz12QZaMrYxeHJ3xrY0bjsWuDkfg/c6USZBDBXYcVkpLLNE8oT
VTsQxtJFLBxs2I8QX/Ey+vUkSZrPSkX6VmDpzB7J109hePeaEsqL3NaspGBLFs5TKIgHMP1eMwfr
Gy/P+hr4r+g37RkU3DB5WawFd28cnW93RGu9jL5Saa6yb2t81b8YoanZpyZE4WDJOpUcw3AFr7lf
9L7SFFbEZRDRnh+jBKmsXClOdHnAujcyfqyQuVolvOoiulNbfpODHkTTkBZoNjU7B7olBMj5V70J
kiDHJe5PT+MrwNMKCdrAQE4x/utxEbclwqGp1kvJnZ0lGhrAfo9gUT7SVzS1mxA5er9feTRToXWf
U1UmHz7t7SWnbY5LIbQ4FhP1egw4SrEvZ/qmO0qC4q4DRhlMUwsfQEmf4welNqrKKMdFBcdbZJpa
A3Jucto22yTZ/tBHi0hh8T511c0yYtmgFtTIrr1rxrTA7XaJrdOhfdQ7uzyDOUTBIB109KdKMnV4
QWLOA/Yxl5igXTH1s04pAmeQrtr/fbZ+WQdt38GmGVZK//U4a+2Bs9iN1ortkAfhOgFrBb15obkz
A20tEkuaUT0UafOZBmM/L0myIr2+UijOYlCBxS0Y9eSQB4yMxrSOmMlW4yygIZyU9ZMQ/iUVc4gu
XcQ5tF6DBIi99Zc57KvfxsfzPqK30I6mzcCnDiU3Xf35P1L4uWciqmLZgwRheyVa6D489pZM5E2W
fq7lZ1SxhXBvFqvzGri1AHAtNBUrr0IGeGy6yyXOlIhQx8nzAEriRuqFm+O4Ezv8eJ7t3jy/NF1L
d0sg4FwDY4L8knxISBrrs4oW8Bq69YzGoDhgZJQOhvslvQpq7R74zx2ydcFDcSIC95ECSlH3IHuv
yJW1DQuf5BvBf4VWUh9OPte+QlWRFyTjBjEn9Dtx7ArzSSoEn4XEUwmJMb3VpJrc1IgUXDnxFXIA
ZGVQtFpP5ogf01s9u/gVtmCjI92cZF53inux9iQUd8cQ9+m7T+lbmOwddmVOJoIja34vm0D/Jc3A
7QqVtAPT+D0K9hvD8gp2P3+kEYvpPRv3mwhtekc7A4f7l6U+WRV6+w30wU9DDT82UpHhkwUQXbhy
PAPcGDzpIIsFsN69BShh0r3+qdxCJ+/ei8yr3AOxN0Dliekd8M0uiPKzEiUlOhBZ/czP5QQ0rvMx
bmrv83y970+gabnyNEi7ZYMNyXsQzcrH6FSB1e+6PUy/UvzPbaYWJLuPfxwFtc3LLhDbOn6O2OIu
03hANtHEc71QSRS+XIZZesr5rkdvn9tFB3ewcZy7FQw6GA3KjxNGGfOb0P6ROCT75ibpWsG+piFC
T+pfdbnTHTYRw7MW/HF8tvMQcm9LbkPpuGY125Y+8xKYSEuiMpTUA7i8pgdzkF5HcM8iCFqXcS3u
w3bGKgtL5fCQ/mdGzGUqVT+dbWirkV6wIdBUGuVKxz2QGm65WVCR1Ikld6lggrQpPsEdsDQSj3K3
U7ZzwaPitaNKQ514KjRY+kWaF7zSVKBLj6n/btCyF12KlFisEV3wU1U1rs9Nbp74lnDcjun7yM0f
6+JBF6kEI+ZbevH5x5uLDg4nrCZqkWkdz0oUd9M+S04GoU7z5CQSn4eck0BRyVOiyZf598Yhj//e
10cCLO58xAy0ZaVWG/3fjFb9xLPQbXFgEmPVHKdzqE1dsw4Qm9j+Ty51mY//nWYyU+osb7NGvzgF
7iFP567quaMRCHzohYqNV0Vc5APwbNGcWovFKGilMI0lhG/WHUY8nqfBQpIiEnm01LB+kKY/ejT8
ONa/SDRxE7j+LCCmjsuYRC8o+tN2JwsKH3YsrVK1Ei7MmDgm3A53STJ976rNLQ4j2LApG/IDju2Z
IMw/L2mDXyuTWeY0QDYJmCVHw9AC8IeattV9aoGy5QuDU7asGUr1UarlJY08kiMq0SODpCMQvd2B
o/xuiBpvII1rSLBbEMAj9RHnSQD4qrGgj2z9Q7MQPwkxanAEXzm4WEbobqC+EHtsPFdE5ryagZdi
Lyjsyj7QbuEuzjVavh2InvG9OVzvuaJP+65LqSqNNSxlwQuZyCivkRypA9nCV8q3knzgYStnZ55V
AB7HoBJNjDcDTUOvNu4iycmOFE6rYZY8xIP0oGDJw8emRoL0/ZMT0LRwEen7UeVC8PyNtyI4O2zX
GGTNaxJTNXKRe3p/Bt7K8cNWreKFEAEEL28HUuCbxnOrcJQV/zeDLx6bb1wBzllK/+CtCHCoHkYa
L/tn6ZAfnV95gaYjKZ0YBnaAZtz6uAhjIe7vdY4HtlYN8Sfpl0YAaEe5BCkBuJE0dcN5e4tTdbrR
raPHc8t40l5YcoLNt8FVfGN9aAsa4IusHVpetoF+w2hewHUrIzVH2PTthfg0PdnAEGZqDp+K6FNO
Jw8TDrTeJeAyAC5sW4f5yfBE9vFX7w+yYQ01RlzVKpADU2vWEjIBLRj2N7Zj5pJgcMpVUXnzfP9Z
Iw8g1jYSKJrIEHla8opGRdaOUYxWc3sASIsODuve7z6zWlOuIURtAs1pV7WS373PM4WzN1mvTHXh
6VkeZBwUiOjrUpwGy+sU+CwpnhEQ1xKHZAcxxlYUBgqHjXUoPkIFmQRzBV3MKxiIOR7Tkg58H7kQ
fCfVOsSl5UeY2aXpxXzFilSVOMeagV2EQze6/13Lj8BxdlOFnindB0ToLwt0BjRYu5avhGfXK4OW
bw8yReJTXgwogIUyv5baWlNXedwx7Tuklk8eo+YItNDgVSO6IK0mH5TSNiFHHe+5YBP06lQQxSbK
e2ZC/puhuihP1rkCgdGgLj2Lq3cAG23v9KOIsoXFfGgNAwpP9a/i59ka9tYyZpGrdUxlDszwY4pu
sKKqAaIEb8gYIxv298Gus/Pw4vgShs5qOyGW4iLq2Vt735B2t4avAFoSyuFlZh8UVKWJpygSEE8+
txfjttb9J6r6TMsXw1wJcpFw4bvUePqmH8Mxy1bTmeu+Odm3q8pHEy1UExjunSRReNxLOq9HAibt
1WWI73i3UVtRdDBjlwgwrEmlzqxnrNimaTVp6ba5eOzvZiIxBDQ1nziUEzz0qhExGJzLnaKuIeKn
MtacdVHidOXvQkXHuWjA/0VNw6int5UrXQTqca+V4E5gEfaxysGzCqaGi1slXBi9QOpotEq9IjQt
/Y+uwZs9BIvOIck4H5eBDo+ykQ+Hh1/w/JMLwaVj2Q+cX5PWkLz9l1tG2w1ACso73IgkvSxddaNq
yxbnni2/59NxVucHUe71i/VxNujUssFDoVdkElKj7LsumR3GFcajNWBTq3+hF8JRV7zPFVdlfggl
4JHXigMhkEkjlwB7fd8egqpJEhlvDB8Kak806psgcidJCjzCHLb/Ld5t/NcU3aDAzqULWL0zv4LZ
fm2RWEBWc3UMYxODNXTCjhb0np3yYpMTHOkBF69DHfsCdFlr7Wg69jWjHAMxFsmNeuj+lzEMGsJB
3Haa6qomZU0DC44WrrZMmy9Jafs0oCE4tThiGHPpw4lwJ0sBprJ370Gr/06SiXQf83P1dOTk288r
g5x7Ffg+unBCWizY9AkKm481/Gv3nRJO46Lrj16Fnvh1V+Q5X0a0z+VzZ2jCzOUHZAIP9DqZH4uV
U/iPnavqinNx9zAEqtDCJ1qCPjEhtZU1HoolfnqH5wWDI8yUb/51dBksSyeG5MnreEDNiW+0uxE7
6/WPXOrIRuefjRuS/xEwiJ0rThGkQLMloEXSWpmM1SBADCPR4gx5b4S2ravZh502SCLFaprCS++N
Z3AkyUfbcM9Oi+mXDD7GoRml9w/LTNnWctnjouiZH6FMYirYTQEAFEb7/axUx1t+9yTSGlSOgM30
YkM7g8Xz4a+hi6CYOFuskFYk860+qr5++fGZh4A0MeESAisuFzb3sqqQ9QWZchHY1FZGMwKwPamS
YuLwpQyDILBAqHrLDFQF5YCNGkQQP1S/GyPbfoSZ658EjVbCRx8a7x0yAocjxEFMKHGBsTAkTj6Z
dDOpYeMqKG9suhfHfLiEfd3Oz4HeCzIW/lL5TjO3sXABIBQJLEMYKv/D5lvfEPwpgiElO9E3ZuA8
ecUEvzGsSluDtn/UyyqpIJB5tY9o0UjHqb9zmdg2PzWHCyI7dNKbcXnmZrvLX2Ez/va2BVJKFx7e
AxF9nS/WiO5zaFPhWho4zgejpRm1+JsiU8QtbSBOvNkKRWJEBcXXd2+GDyx6Zz3b3fFeO+NWD+Pd
rZKMPJZd0tQMRf3PPdVIUQoHI1kAXgN8+kXtVF3Vu0cY7KCaf9YvXadHPmJoabOMvDcIbgkDmDui
k+Sqe1+KMXhVpW5mNrLPygxQbfqtOMsvrcV0wgaH38nyMmQBOVVVwFFrEcnPShxxqukIPkvPMI6T
5/+Td/sV5S/rSEIUChOse+8xwTvi6qaw2KcupUxNqeEO/k7lSEia5e1hlgEIrsvE2K/X0fUplP/r
nrhIRcSc52qx5NyKTkjDAPKNRQn3pu9Y6sB69cG9aYohTI32E1mjYz1Cinb/DdWmwr941aytYlUZ
4Ilf/sjOA96YnbJcVt+y5V2eZOSlu6nFEpxTRDMw7eEqC6Ma9TQb7Z3ZvWGIOKX07+LWlGUquDxn
SSZ/cl9naLdQMrHXy9sOVcYAzblhyFqwLi9TN+622t8IR2gxD/Nl7Ip0cfFK6/nF1LwF7DZJbQj9
r002rIdDHa4mOBWIRxA2htC/uuAwzKExizSKTeG+5Jq3zk/mm3lIyfiNzfwmWw9jRPWvF0urQojw
cSKodb8jztkPGNfW+GIQUsMURjUfvdhszekyNRIQZci3PfACd6LpksRhm4x7UJ2FGtIOy5LTlvJi
S3xW02ignU62d47U1i1AOtS5746Fdu+1bRErj5VhKyhabmIr+VHBNlu96b8rwVOTf+LD4HAZBYLm
Ieh1YG3XF42nx8etZFX+U9kpRthAQFUnYXWlgezGEtUjiI8gBX1diC8ogHDz02xOm8PoUfhdwx7e
wTvN3DLSofV17MwBgTzIZVttBML7YxG9zsDBXVckGEjWcSUuM1Fo5VVK4yHHvlXX4OQJME/yNyYN
jAV5tX4XX90YF3cZvDptAXBPkTxEfqcFL/gesepH9wPfqIFE9AOPUTjoeF2osz1iErplBDtcn2BZ
QLSSbtdOeam7ppPENdQhbX8vol5lp6W3eb7RT1DB6bl3LWZigmZAzhDSd9q9UxwN9Iiz7EtA21f+
WIGxbftDj6rbExE1kdWoBGpxoZydFyetkwLW68JX5i4tyN9W/7tDdKJrnqeQ1vLh1k5hKFqQnePt
zof+WCYFOynzNX4zkX1MRnI8p5pWaN5iD8j4aMlIdJVpjzOjzLPIMuJ93UazSPiDiLVM1UzaBFCA
8Hn1dmCJHCbPUuOzxME/mId9YY1hbAbSN0S06TSI6V8mnJg3N5X/MBsdTk4ZjD0J2pHqLJY2iro3
pR0a5oxM80/SuJA63hSgYUd4b4yzL6XogAsc4YpzwldOsVtq+RkOfIDz6+4p0syOJse5rdWhoDaT
3+h9Hjdyo2n/PJGhlzPw02rgHqKKH/5k3pXiMgMFvUZyKKeN0XsXBlcmF8OE9ZbkuwCWBFvCIhlw
CBoIx7+KoiqmxvYjiGkGCG01VTL4AsdOWmjBj1m1rjGsRzOTBvwEAK2WQwrzPwUgWPgk+Zxj1HVz
lr1uCRRIVunXAkQl99FPLxRqBOftLfEAqbCzYQAL1gOg/v5OZmtRebPKqw3LnDr2+S47XIbRX/5A
GTCzJ92XSG7oYFSms/pOtEpiuryZ5zWZIBVaVE5EWNoUsOm/GZmzODN4hTl9xggj3JMZsXzSbipL
iiXMxyue1+CekJNu9I8KGVAXHDjTCqYmNDioSydYW0HQ3HfDu1sgOXY/wYXz6rwIcRZQjrD1vRYh
4BEMznYRGW/HbjHE4j5lupCtK7l18ycGZ76t4HghQAN7JzUsY9Rqz5BREarfYSbLY2k9CsGIfEme
D1CM29tyW3FXo9HlJx1J14BgdqnopMtSxC7p4lC3gBFNv2ODNQRQ61wcYlacPgsflxUIUPkDEL/x
e/srW5VYqWTGZf0M3Pn9s1/c+JSSqBk4gzJoMGcKbwjbdE1sH5JqNZRpq2mu5lTBIE9Oqsgd9NWe
INlRjtLBzukeDL4BqaXb4kCpBCLWNeLEnQjgQNia8aXVJD6akV2NHqLg36gd8dView/vwETNXXKv
JSXrMiuqrU5P26Xny8rWmk0FaSd/DMvKD0JCAKPv9T5I07yvnIj/KDGAv7dSiu60M90jevqT4WxZ
ii1h32DggT9oPdQ4Qj4W4g+oUFUUFoZK9b6KKzCCh2oEQjmjmd7v1sZ13UqirXlOMxqME5vNqMs5
8C9cVYOAuYnRDV7Sc5jipsLCRCJQ5rsRG/ho/TXzESPJgTzUB7lPDLl8CXdh3BP2AW14MxcPoJ7i
zMeIW480UaJi7dTP2jK38JQn81/0TTepOm3KCjCar2Rut11THlbBKd3g6ynhuYo9lxY6N/xVrALf
NDjyHtLbQpipx+9pLhEoCGaKmlDlS7LZDwSgoduGbfGkI6Wur7wwZd1ss47rZxa9CeGrC4ZlWhce
ptey+okufovv0jc6tbPqzUCf5gTUcrRd3TLpBiZsqDagX5epqU8Ej+MAKC7q9YxOzAphYf1eohQ3
74VixMMGhFMT2u0DxxGcgbwe6okoDIdN4v2TdRY12tQu3k2PA1SUM98di61/BYDADoIsQ9UnxkZz
ZkT++Oqa7bRPBjFiO8AzZfaJ8xPPUOHm8A0ClJRXl/P5epP6zplEJUKORJDWWE6hIfWLTNpmB0IL
Pn+/o7VK9ed/L2MBbu9MCtWGg4CWjSiF6YSQnIW3dqZ+8tEMcse4QKGrscqfMkJVlgyPRYSdWA+C
T5I8CtxEDQ3XqkHBHzJcp3X5WkV1TR0OwaMHPsgNYSwDh34g/tV9iTWSJZZ8vT/MFf0bRrR2WPET
9UwUeVZCOHim3j3boD8WLFRyAQCMHPOoU61uHC8tHecVnOO+knryHJXXFp5A9jZw1dbVycBnZHGY
o0JDjvIjd7G3isCP0eF5WaUzBx8bBEMR2Az+6whtIisOu2aeYZzN0KwjgejvIFt4lOe2bU2f0Z7H
BhXjz4jasabITL/f7zz2h0vJBfu07VnGHNfxFbRL0/dGh1XiSu6ImMoVviqjQMTHoadswqS8+kjB
RdX6+m2aTkALS729rfL071c7guWlblVsBWnAWo8vJmG+M+DKv8+TWynLwGZBS9dj2BDUhrlGPPTw
nXrPN8Zro/qB7FopIzUOHth6+xgtFwStUxMLsBqoWO7oabpVSKJs88yDfUswFHRZKUdHuiyrLMJg
CY57C3wLXUWUUxWZONy1j8cdnAq7DqZO9+GCkWOFFykAmcRoVYkWiaLhV1EBzBXzWe9hTKe+mwDu
fQoSfHj18VWLQDtiCxdC6cGoE/2uLvJVtGURUMuYITrrQGZQSx60fE9ejU7uQMRY33AUsjQyigCI
nraWheROjq6wdKaoKtk2orGoTjfLa7c0WqqAhOpfSnyunndB3u9XYHDJ7dVuWiqQBBuvSDiP2eQS
OEkWiYbr6clfnpvPL42IiWIDjGiMFV3ytQT+Sv2zLACtlI5dFo/DYRiULMg4QVzVyasotqz5212A
mcWWvl6A1A/g/3eUo1r2YVjcvEEgdjJxOwv/dY+vkEOP53p/9COYhPq0QLFSmi0K5D87lh0uGzgH
3cq13iR++CnjFDd624D4rlyx7ndNA1GwdrO0rw9/LtmaxUQF3R1Ojm4RCG/GcLPzkzbnFd4yJWX7
E8xboubtny+zyV92/yxLFKdfKc16pZnMpQ40Y241EGFrflh6vTwv+tlJaIdcE+W7f8LJ9kw8ap3Z
wn3H0o0SYNgRHvhSmuLW1B3EVA4nlhG2gue3YyNO1mu1p6H5n2cVDHR/j8zbNtojg+RCvATDQJ3L
A5UOxNsa7sEyZ+5mq4rmPMt+yA29I0Mc+fK3xXbIWsN8YzodOVQspEPN6pIjL9T6awXlXEsrMWvU
+qEgtImEi2nH7Q3d2O3/YR8GiB4bFATrc96CCEN+hrYiEMTqKFkQWpzH3HCvLYb96MkVdr24LY42
PLlKlUv3rrXvlu3U+V6wLeDIo/ZNES6cM2GlbNKco757j0mxaNdtUnra/Te7PSZx43k61mv/zGfY
Po+yGyHsNf6LhAyoUmnTjq2o/ohFATKwGXk6vBYaIPDwyyAFZRiShG9jVUAgoD63Ofct9gsfMZLH
wDZxuZ9ytzIFHJo/OuPmPb3rFOUCeh8S/iZplOnTq+6o8eG/HPL4tEv4avrMLHfzK6INYLvpAuAg
jMhNZjQnodFuY9yvySVMdVQTphl0N9M3qFuVDz9PiNDmQSbA8q0lo1iweKdgGtITSi8zPjsnvBNb
G29NgwwNmP4QhgnMrGwDq8w5TFQApSzL024bY+Mp2n6YFNaSOeLgZVopqXdG1Yxab9HXYY4/a5IG
d5b14Rr7lWn+thfsOtlcFu6cNgISGqQivAChuGE9MYLjh07dq4/VkpOk1OP//imwPNjPU23yOz/a
yVGGsyAmprL0dsMeHidHQG6M9hPZvaTiLOGgroTZo3SxfC4nGt+cKL2QdZbDrPhawTdJsGMx8Y4K
kwMfiBHcchz0CgnE04eWpdqaFfDbWcJ7EB1UVEc0oKIn7n1/erL1EEkFq/xzYtMbZbD6KJqNWmba
1UT1wO/vwZf0lazqBxc5mYTOMVDJ5eRsHE0PfogeytoeFM6n2tbjUxEumlutgDmU/t7F2ujGGwRw
L6+CAypyskOzRA8X852IfbtCqQexae3pA87qr7Yux21EcaEXkcni/ipWkUcuwb9tYdUhbrNn/Jh3
Y4igujGAKBeU1sUUzLVdvli76bWwHXhJC3XpQB77vbpxxg/7J7ORvoEYNn6hsQLY7kBNows/kPAS
E3BLWGo3N52tnfcpwNLUyMsrL74U+HDP+ECKFAHuLcIndNlUy8bAKcTHRbZ2ODYArv/WPxI0eBwz
8LZLncTnFJbXgEgaBbx1ZuO5otrgrNU25ETwnsKGXD666FZDAdUSljY9QxT9qkPmEye+DuijDXJu
Etz+Z+eEC1QPAMMRMRW+aETX+n1dISvdnEpt8j4kYUINhQw/FqFAnwZaGbpEeZ4ZCzXA2I8H/67h
sxNcso6Ef0ePHcJNU/YKqT9itQd8o8bwi0d2VmNQzFqdZIUyFNC+9PGVua4Jn+wTatOmEFI1/ImO
1gLSA453HfyWLHN/X2Kvho6XuWTmz6oqgBxezP3sokYG17HgbyLt4+tsug1pJuKyyNRH0MUWs6rR
epoOVvrUvew+Z5OY8T4BKhMiuiMskuPMIh28nS/cmqHCYO+yJe0wQceYeiHbyjkUmX+lW4PJku+6
0BZ6zstGdJ6qzWkLMCwfycs77IBkrqPPvMal+kinQOzWkXOh9dD6MlLm16VuOHoKWKlaNKmjCsN8
ob3L2YBuMfeKNqS460w7/8KxH0IEntMOBlxvIH66bF9ue3eA5VEMT7ILAcqFQakvaZYuKnBDgtTi
7SDH+IX8bax8cgYEHyrRijg6o5GD9BckQVUvcPtTM3L3ir0LprX++8aQgGARtBeIM3BMqsyjZ1+N
wydEkt10JPT28rcPJtKckGvvfrD+YiroFKT03RAfFlSUZ+kPEMpuCMcQGlrn7L9GFwcGO1g6XyaO
5w5x1dvpL2gcBsk8oNJn/lrm7EWLdV2xr5bKCowK64KcUKpcGHebGgXA3H8lK+uVtkk8Bn1EIb4K
PwOenT8fGVeBZGoEa/s0lqMMY7GGEmA2Kt9HJWlHHMJWZPqdukMBmkvDGYdhE6zR9ZgnlnU866Co
uxwrrPDvzik0R+XtWvJI6f4xxoeEaNcBG174N/XPbgOU6+WLMND8V9CnrA8bCuUbyHQLDy75Jrg5
nUfZnA6pgzRrule6BF6avWhcAU58h2LOlEhInvxkqj/HCg2+y+hxPOMndvLg8Phh3Vrlxbs+lkIv
HNfNfwxTf0XO287azS8ENnClTEchdugeMRxB7D/l8Hm5DsDoa+CeQyqJAnNOY1eW9XonWKQGfYYV
gtiycQHfgv4EGjohMPpUgwZNvnZWGYx6rn8oASVfv1Y5AiQVGILz1vquxyogcJRB/NNMwFxDcd/R
AcxUF8kz9pWAL4cM1HhYCQu4PRHr0NH6LQ3XlnWmoXfrR3O6wcXrAFjlO8L/iiXI02MFofLms59h
a+or0YvAHcJNZzBUfg0CYqtl/WHBa2kJLIZywapucWYhjaSfFm2F8ofMiDarPAss9YPkIJNiHpBw
9EB4xKY6kXndWQXN0JRJ53fZyGpP4pfj1rwvXeLysFqHbQ9rBI0GrjRj50QJ2To88sXP69adCd+h
NfPl0UuUUQ8snXwH+rdbrXjFPaofZBsGHixPmA0Fh2yN7fWXqUsusMQqcihxaZsidSRq91nXpIJ2
qFLbUAkK3hDn23oKO7NrS66tfC2cEBc9jswdKInT2uaaXgQHHtM6dFuGkQewzo77XwqedpgNC8Xu
ynX9U3+HlnZOQnyrci97XeHpConwi5GHLVAQffaln/Yuandl+IC47E5fM8x7Ka4By2aPXxqX/n/V
WaXahvFzAQw8VscUj8l2t9+JltUnQw5Xpm0imnBjP5TIsnUumMnQltA3j9W7yCBpolZ6rbU7qhcw
aDq95MPIH4MkGyu3iT/lMEqm3feqnWfoDGx2hFEwt01Giv7DZFce3A94qMlLUoZ4RltnXEo/PIxF
LS7SZjUfRRlnK6mLzQP1Wyo1s2nnJ8AZNVix5sv5MiWFCkOsWof6SdHWrodwvFxry9AKp4T7lYtp
ccstreQ4YokU36pa8+OLPVG5oHV1SIyS4LOvC5c5K5oVsvVQfgpWsCiqDdPxDYZKs96IfOeuN4wD
/vvzFhrjN3h/A3TKjqwHepTvPwj1k9276okGjVdtXPtwsLE10gbmo8lym194OpxcyCwGS2mkPza+
FqgX6u4rIvn/ag3k32k3JCcq0/un9db38C2c2umQaNCpIOllndbKlFi4MFt2fa3j0V8D4fL81zhf
iEAqdFvHeL/ljApHrflo7yLc3OnbGAT+/r2l8DT5KNI7J/pZ+A5XHbpOu+XQfX9Ie5A1LgvPEdaa
18hGjDSiDCSNu8YlBS4VCelmVnqcbgGdhnI0GQ0tUS7uUb+Tj88pgJ/+frrnTCHXUzsGbWHgUc1E
UzSFhYYlxgellgdjhboeGNwtm/QBS9ZpRklbJ8fhr94t63S3/OKLuSl+RDRRWtjCMnnt1k+lcDpf
z4g+3j5XecMtBe4f+SoW/Jvq0YRLU4FPJEpCvMwr655Hww1AoBGYECVKgmjuH22Mu7EowCQvwJDh
qJu/+QKfUfT1X0SRGzCu2leC1d7IuiRDEMIVCZ1mb2fUMbcBRXNEaEEOoJlPS5ac8olLwaNLNvXc
/O5GlwnqN/FBG0u5efMgy5kfT5w+fjzPz9cQEVcp1bMQwJHtwb6rQ4P0WQy69VWRDXEiP3BUMlHO
f2t1JgzH8oCg1G8MDwiBQMrTdKVStusHr9VyWeCwKjXMxCK2MeAvWG46ppOyL+vO2KSqHy44T+0g
sy8Ks3NuCCjp+aU1mTRte88Xa8Mk7VJSiGQA1Y40Qgn3jopdObqkmdjEKUQ01K0MumQ/eZLCTZAF
RxLV0BAsxC2qlASUlYR5JYeoTV0EQTOxCulzt7utS78SHnfeE7xH1XRrvsutBKXOlYTxmCN6R3wT
nmPsejIGiQWJWIoRyajCtJEij7XujhB1SCgaDQvro5GOpwpnIsQQaDzfneT/oUsMMDLzMxv7XkmU
7A3CEPQrhzH2sjTlCTqpBKa1jBD39tUj9afAOlGi258B48QFGjoQJH1BFkQhy089jT84kwy2zHWJ
ketelBG47UeBlVAzlfzhtrs906URkUxVghxGW3oeoZn4TVIK7iY56zhCdmhnnkU33Bx6CzReZi59
dEHJ+G4c/ma0BUD3ZkZtpQWMtzi0XVA+CaQjocCBYJc7an68QAS4K6FRdCeBFWvaBgv+2t5fl8bj
BjVyNIsSkmCpdQiUfzE56nEmbhI7g+I0ZmWMOc1DWMYTgzw1Jl23OFAHDlxeu4EWi2fPJ6WD93Eo
XT0a/ci+hXT3X0bbKCxWNWYYSWbsV63fUk2+iKr8AClpMPi29pDPXyVmAtc469HaygDwlf1F+KJ/
CcW16Hd62L52w72HihMbtLx5D0AwIWFbH8LkUN/6sMtiE8LXj3e9EoJjC7zCp3fy6qHXqiNNs2Ld
TK5BJIp1VZG/TwC02KI0DPK6y3dmq0n2yxmZC2ZdyC5WrjoTxYP7bHRIE1zdrh4Cyy7z3Kfcl7I7
eb4SIHuGjYw/0gRVpJFpJhnOm9s+1m7tte1hLFIwxXxfAdoGTgP8viulK+ZrzihpZJYxnwO1h6qX
4XW2ciUZxMZvUhZgQbgz/3EdbUePoamb1Vh9QqfwnXC0zoUTwkI9UhlEOyUbg4GVU894/vhJyVkL
4soQTiyLqp5Agt9RAKEQMS6sDWKg+Ii1TCaO1kWw4+rowXv1/B0eIk8gXM2RqNSUhCluYyYqtavK
sXD5zb41qEsA3qOx5mqDxSepoYGDlwLHYD/rwus/9j1b04Lh+8dtQZxNkjssOFP9NjlzU02d1O+a
iWPjWr+XPrrpkeTFUsEQnCbWDEiy1fayMv7vD+Yt8wgxES+eMf1V7rSNjBi3TDCYwBuuPz/LqkUI
tJUyOpisd410ECZT2yoahrxImtay36BUCDaf4Kdg27YGfsBlnuK8mPpDMekZ2fGV7F45qks9ctHn
6zBB19Bas+/vz9vp5ula0eUnyiLisG76SHJH4FDy83f69Tale+TZRE1DjVNhtBWAdz5+crQ0kzSd
8828NsMpz/AtkQTU2G/9TMgRP+WsLTPUhRIgoU0Y4OAdWMpFYG8Aogj3JeawYEPuWP/D7tl6eM6+
oR18znZxYH39J4+erU41iAh6pDBn/GdVfoygIOJPrsk0fffP7gAnKha187FT2Vo8uf8GW+3d/TKb
gOktUmX7QGUD1k+pV0Cw1zz76jBiZbvhQPj1DDrPa9Cow5IM4OhfIoHQ/77ZmM/VsF997Lg+2rvP
UFzO6C/JYZBkty8BCspbD90frK5iAH2uSj5XsX5kpVmQmV7rT4HQBg95ClbcBzDXTNf7l7CRC0+j
ceASwX9Qk330RLENN5NAKYEfxCqvcA85UYFeRjLmIKbrImucE2oaZnfQqqh6ZhSxDquSQhZ3lCno
OkPZFxITYPkYcTmFRExQwXU+rELHXWsSK8Vm0ZualC7e14y1c/wkCWMhi8jzS7RDFFb4cmXQ7Lfh
obCduva4tRbCBaBGFvvSUDt7n/Vs1ovz++OMFvgNy/JTyv3rpsm+bvzAOJfqxbHzDlFa9H8rvsr0
toqpLLvqZcY+mXjHn5XSwPEJxkjALyTfqYiyyEJIkqWU5dlSkR4JjQwAvhroLmfQPPBdiEemWm90
6WSlHkTowWT+L2E+2M/rWCandX+zlZUaTQ6PNCRTtnS3LZVBKTaFAWLhHhRBFScULqyQXda+uznE
GmmcJYu6EYbRiwm4hGJjWTRlt39Z0F0BhpMU+9qR5e8C9B6K33y6HRje/qSTJml+3gurVQThc4iD
+ZMGzzSy5qHNyEISZk6vI6KO9i57hmeufR36qjh58IJa3A/1zqD3smh/UiGI9nIgLsGyhJtvEl+f
I3fDby746ee9usAHCIOMHD2lGZk7M6bU6XBUYLEG8SjKzWPMZ4Jh/XL9gTLLI1KXTq/5hNPKcK1/
/nrBCbRed1sKpD/AWC2E+9mNJIw0YnwSVZ8ebhM3diWl7k92vM8Hm8b5m0ibhVBIpZRgLZHX6ZU7
pzOt5DEiuvI6pHci3rPNdrQ1jBTVr+flOj1H+6pprW19Lnpr1pIuyfI+xDcxpZX/OlARlJ6C2heB
M/IEMOgo6VB/7fbL05V0HVGzUGPTntrD0FcFfeNFRQKvXXoM3BvaJdEYl+TUDSNVrGh+uZuyuC6p
ficb90YOUyCHJRFTJa4xPJj9SyGFEYSixV9XU61aiBNbPM5iLLokQZCgGcyCuS5hfEuv6ydcOwLo
RHxrySzFVPTF2yZzVOQ080g+asEE+e/NaDaAhTDepoab0UgEiArPxuUVawUabcr7l2x8QD0on0ju
t/LY2j7r4novk+IDuZvCS27D7QYuvdkK4MkCM5ox2b98ndo38RboJXYMfwUi+Xxq15xvn1SzSTMb
mi4wcCWcFZGr9rjPiqNO6QuKr2RfRoPlysq6pc36On7uruAgoe10kkUJPD6jzHNNcLmfb02RLeL2
PImDMnyPSh3BbUZrpR/ieIyXE2FTtQSo7Lf/u4zy+TtyVbAiVpgIdLZt6+AQ5i2Q66U+ofx44Svj
4kYPStw3QZ2CHHtumthQnejFKP7yWkHzYH0S7b9dKGjzb5+GmrH11v3qjIQrLTz452563MJBhXNc
i5Y+ZwTiKv+i2s89I6rO1IipXTptxvGahxVvy9ogiVw3l4OIOGUYu1naMmsWpwuOjbGhdW8PluXC
9fOpZJrhxPODWYM476nORLfB0vKmfH7OY81hB2AbqSLuYZBt5Lhhscp2PBOc0EDTWMZsBGKuW4fj
LjxvYWle0mDn6v8LNPKMtEgboZ0mvpBPMDLtP+P0SOU/tzt3O/+u5wtitpMhiIh2uYlXTeJ9EPpe
8tF93aKNs+41Bmro+H+7ZhPFEIP28CCCVZHvWuZ9SjRZdAYMdY3Bqd3eGxz2uqZXZ8XHXJEIcJc0
bB34upE8lqnaiGX1poZQA90TrOuDlGk4vGuN1fYZ5iEaRNKmhbN8g+lYN5IPbnnXHt8PM9+R6X5g
ef35a96pdmgMDeM1Gv96UoZcJUi22eZjX7iSiafMfO5jSolZj0X+lR+MUciXhJOJpTocUklf6c/d
RnbNuq0GVz8PcV/1lv4Td4TezmDIJMpncN3ilW1Ottw7oALV+mTIF5xrJmNXpL6qXHtgl4H+67pI
qPbzP8lgeXTqFL3vEEWFl+C4OfljYbUlVVy0L8x61HJdOex1eDh4psjGOyjg9qCB0Yo+wJCUvtB8
FVkm3Frcfi+FyIJXoygWeydTQvH++wKoaRlm/YUR5tp9qCJ/dELqMZYpQG+Ll0liq3ECKPtdqRrB
W9bGOZb7KOtQPYpu9OZ/pPCDksS3wwUKnUhsDB/McsyNH/X3T8n3g9opSzXA/77yYC0kmDna7tNg
mXvQ3Napx6Jl4FiS8gw8gEKU7EKasp4szPW4uH8rf0t+fAfL1oAzgFl7TO5PUQkH+IPP0ZXncxw+
Hek/TnYbgcegGkeAInfksZMHGHoSqsFplCsy9A1aluG2kYiwIisyfAdbpR98TK4elbcf8Gh887y9
EYBMZwKmGRajZ9YxSaHyihIebvSmIHxseXc3JXknXMo3uxLqg2abpxLcSI0WYAPD1zPHPHJ+gJmD
Z2rg4b5DqhMfI2eg3en/mESpU5NXaOp/FZfrPQiXR9Uur20W0GPl22zLyt7CYvSKr2ONe1vqVpTj
XtlN7gOGK4EvWWvRh7ZFn5wmweRXnYWgKYzPbiB6duaVlufyaBDcKroRYO9GqryiRbQb6VEiJR26
2tMR7sie0xS4oR7t8k7zCX6CG7n6vJzU94eRUKg9fURAEozNMS7MSvdboUfJMs80qTmfBqVgu0NV
hUyFFDOC270gKCYb8RyJFX1oAmDsV3qT45DMW1uKnZilVWtauXgdwwWgu9KEBu/f+m+R6VKee6NS
3Yrj5d9n8DuYyxp6gDSx5QcAcrfjD/t4mcHCgt3TsdzU9OW+aPsiJDiN872j9QNto989kPJAXj8V
9LpX/Ebf4bQ+FpRdn4iajuql2PLusGlbmxdwnMdCrNd2k04IUSOLJuwauCGLyTQLdJkeJSZFfQ3b
MUy3AARwcHtseVJOhxAqgeASuhiTCxnQDp4JUe+f6nc9AEodNFZO3Du7sj+5Laa25CakixcTaC/K
yjLHjTEyPNTn2Ifa7mJQpJ5FSjNicHHwOXedhO7ABv/0We/E+cX6cJjRG9EglVRkDLa1zi8pzJZP
m1S17pdbYLg2XP6JkAHfd8TYXVMCTPDSwPH26oPeRUEVOUSppQ+igO+Z/XjMgKlQ8KyMePrAu405
vdrY1HVKRQTyT99dxglSZgxX/o6RShbVrjgKSe1j7uQgK6znFlSx11WxFq3ksaRIdPibbi1pybAk
v2GYiCxkiIuB/CIcp6po5/wBK2ZGEduqQxmF5UnnoV3O2z0aeglTrCc2BtSnlys65T7ZqiFBTpwQ
iUospcKbT6xN4gvGIaXCmM4KufwR8KTJgnJgrM7qTN3hwO61O/Y5+PRyL3LPX0DBhXcV5KC1cS/o
NjGn1GCkQa05JVvRjie1pr+7LZW3JCQaGkU8uAofc0mosbbAqruK1LO2fyZ6EA4864G7vL9Y5Gcb
PJZ3L8hSfmXHyVE7XycDb9wCk+XLLKfTNLd5D/FL3rPN6O6T5+oVXhin5RIuTLif3itEq1SXnUj2
ThYTmlXlOCXdjx6o7a3k7zQTYUr5PiYF4oTv9JwNuqXR4B9Rkiwk0BhmEuo511DVM/E9pLqrYJ0e
RS30ViALQ8viIAlxrAWgA1A/kDPC/OIY7czV5GcZv7yl0f2OeY1a5rk4RKloeUzKCS97pdTVlRfT
2IlkN29dyCbhRX15pjMJjCv7piLsWzcBLvcyzOSo3bOmM2XYQuAR9MSd/P0c6h+oXjpklynSfeq1
yI+OnX7Jp2Kzzqpp78ECOCjVJIu5+HcVZd1TxBxTJ635Z6/i9thRCn9HeZnkuXu9WuUDyzyoEWk2
qZxO+wuKw9jcSsbIOTx1xQQDawgAb7t6Z6S2e6gJ+I2fStDirbWom0g4J0J/KDygpM0k0Z6gysoV
g1poOQD2Kh5gPJWW0rsbZDoIULpXfRNJxYiBltuZjr70w7S4hUiJE4X5I9DFvg64mhwpD16fU4Mq
tRyBz33DCHk7B+qf/c5p24IJFj4JBqI7sGL3k3a9Ho3QxbA/Of2CzsoOyQEagIMpt7IDw7Zpa+6Z
H6qS+EDLtwYHiYYKQjeowquNX5EWAODeYH4L+rFarc2vUJNqWPHMqoP0jrzCE2hdyMTSJY5kHcRk
auPCex5JMvavYpmkZJ/PJT/LtlcwsxhgIUK02p5lN7SY9+s5bktol4FD57VRu6Yx2RE3L1LZ42j0
CBxlEouAazoWSAL/l0ZAocVRbqThuhUUk6G10A3TEU/QfcYncVb/MfDgKk6puc8qPnF/uWH5hqUD
ixOim52oYUyH2V2x6OIGONPpJjirGet9rLnPHQvGsDoRZuFzes4PavDpJ2DmSIjLVEBxQRK69BXh
WzCTOnHSQcOnQqKspkuRVzT6k83gH9Lc0nyOjgA+/QUfE5FciylfTeK0P0BwphDU2kf3NZnCwII1
17Ad0kF+EnAD2bWWERvSWLDUkxdlhVb29WLFqDpqpCF+URRPhU5mUzLTPQx3lIkwlSXo+aZR9U7Y
wkFYiBxagS2l3w/o4oFrROe/5DXCoOzngBggvnNq2wRa/iBE13tC7CVMDy4dCryQ044e4+u1WZi+
XywHHzFlUJHfr1Fa6j3kI20FBznw0c11AVFIJ8/UnZjHecXah7NpZ/XEFLAwYU+8L6Pvto8yhmIB
Si1LWNN6sy4FlP4NNo19CJeJ32LdKJKR3d6lrpwtwLiIGbgqA2WJ9Icw+gBA2cZrfsIvS6+9Fxc5
bacaIoRj2xMQTJsz/tI+Rfp1vtWFQojsdqcxkmXAv/n2/dYrTX3//SbFoPpPiheMs+BfA3b5RfbC
Xe6bsCqNDINxmHw28Ttz8dko/+rMC9AHYdvE0tfBtvrax59RTrDn47NWc+lfjd+DJANjq4Dp4yUp
7EOV/VYZaR4/XPRKpsTDSlOynZdmE3w7MDVKm86FcNXFU9al48eX8ne0RvML4MmRii0RS7bkyvGl
ltpuR8PEpNPSKPUh38NNDd4bTPyFUVboAU1my0MAR+XKD5EFWSJyBiIBKSqCa+ufTPp7CTsBC82B
mQqqCzfjKJ2YSNE9BQ6oRJcU8dp226v3e3sGtlxNRE0huTKH62VVvsEBhVwD+pX4a1tdhHSH1r26
V7gCXhLGGSLh9V2N6z9UTlD7YtxWFawjyEthP+DNYLF+Lttpip4PN+ccJyNPUS9L/F0+0NtXAmPb
nCYve24Vg00ZZyC5e0suE8binumf6uaQ9NXoRwje1VowC/R9m/QwEpo34/fEYTY7m8LeSJWeMiDn
k4Iye9WSwrc7pkSdeUe4/kaTE4sRcb8FUjSvGh51KlFH/DeMs2hNm7ri2KCjwTjZBIrhIALurZ4H
hutIOn6El4QF99qCDvJ+1T8hkZbyxI3wQcqh57fjaqk0Rt5SC7nS+gWFoT/y2CPjHidDjSupJ4xf
Euajp2rJZRbwnUmYZYQjn0/CoyKhg0fj75QDLQFvjr7xL9QgPDNcMgOeOWXr3rT1Sk4sPHqY/ZWj
74s7xqzvWeC2A4tLlcoChATqL7fNeWjFVgQpZP4ZI8SiOMCo5Qv4a1RNnkM5I/pmH0ZIbxF5vxHx
psriT8nyHteBE2isF9sg8Aml8Sl/RVMTr/azWGMJzFSDClvih04+bx2DRQ0QAKZAiGHu01/89WTq
qkwS7erYK1Jfv/Sy8jo9qjO5LgtNc5I6bBgzrfSbyS4LBurpNqyIUW5TicZwP0Tp7SsHANXTg3Dc
InDD9JXg+fGCsx5IOpuM2NIJHH0Are8EwFAdRIYnZDORVAbFWgWuYgXJIJmPlzw5T3t9PYglsKXN
Uw7GaXpfHS1s3jdM7a7IqDphqmTsSITRbFN2fDioaNo1Z60KExIs7QDZPuS5Jx7WaKmluXjape2r
9tTiXga/4hGPyWYZtLFH9/QvWGsLlnlpzlg+AKFuTSO93UDnMhAiyyKL3tYPqDebpI+ZxoCYKdwH
tNIst4UfR6DxMFZRoK7wgxdORKLDRgJdnHzTzhaFnWLkyi7x5N7HtGNtUokRiTrpiD+cO+gvFL6m
qNMq3DSpnLvwFkylmJnyEVVe7ywIeNMo4/SVAucLuA159FyFK1Ydn/lTwD18VAW0ccTZCy4rqR9F
f4YBHsXirHk3M21BHmLzn/+GQszLrdz9YePgSSLK2ZWISEZB+yIAUp9WfINegJsQYez7wT3oDgjx
fgGTgMD7pmEWFVqoJ6uHEEwv8rHBtRL4HDk1v9MHAhCJ4eWXe1VjH90qx5VIba9YsSVLnjzdbrGQ
8Z/b7HF6tM6aBHXKndarznwm5xS4VmbNiCCvEYSF/yFwLO4fBV5Toa5jDxWr23hZ5ttCF0Hg0sTc
Ch6PSeFpUKCq2P0unx0trngoCte4pbi/CPScnbsJySFlF5uNXBMawi5nbelPOzVQg27SWOXySj8f
n5lSzTT0/iJmitaD83vHjAUv55RLjf20Jz9TYJpibjEg/Tv2ShIjL4/81XS+c4aSk7myEMJPtaQw
1mHlrLbnITJSSaKxjma9VZFr7VSXVN9iyvR4nhXxiuw2lBvhcFUMLXzHNVvpNPoF1d88CfFt1fh1
Tir7mGqtm6oaRUS1RKFJE95FmGTTecjuFxq6ElHO6Zh2f8TYNBYW9GcDP5nobSE5pW+dt9q6YcIH
+3wEtndU4EU/1ysX8WHqIt0rDk5NkCBrnYwETg6uPxS/SjOnvtUTQXLruk8pmm7cj5Q5tF6Eehhw
CW2WRtmREfLTWQAMAXQkxLmpaEJjSXqd4/pNxWk4lug3QIOiLGQuH7/2V+JmiuObhLAEInuXxKTJ
i7gvC3zNLT0xW1xnhsiplGU7TGvEkfV8sZqdAQgOwifWiH3gtmpDZhwlowCEU/P1X4DEW657E6IQ
5Tq4uAyKQK1bu0zRPpOQCOPNNHFPeAEDiniAgi4VXQXJT/vmJ68QhLHYLfkCLsei10x+eFgh+KG4
NGtGyx2SNQNvedfCr6Z6r7gHxj4jRG8gVWKGOhe+iMpVSviIPLBf5OQmKy9LAP0bP3yPMXBe7psC
sbqJZotO2t6PySaOENXcU90zkfxvX4mtftBq3dhrDNJkIi2e3ubCCw22FBw3JPYa6VnGmAxfzhwF
GaPqGDiR6pSRJ9GdH0PT2Q9+42lBJaLY0ZqIQTyXXwGx+XIunk+PVbsDdzno9CBuC6VzeokofawE
VtzaoHf9H3RxN82cGSTuwiQvDbiC6DzO0BLTCCsY7A0QdTb8O4Q4NcnLovTRLbpsAyF8xYzmO8up
PMhpGK1vnB6GNdxiUaZXZkRfF06iscnj5op7yzd2dfJTDBSr6rwKgvvqAAfd29fjCO2uF2vIWCUk
EMCh279RlGh1outmWniDZieMSfZvxvYGXyjqqb0FfnF1Q4CX8R9MAPhwIM8csUn/xOz3IWJfDWJ/
saFydmisCnhEQ5WHPYWyHSGpvzaa3ucxm0bU/AyJC8ZBP+JkF1sh+slnsiyS7rGhXh5cXpah7t6Q
c5bwIFRfuP41lt8fAzzfFj0lC4sdA1V5mM2fzqMpQugPmuMWHOXANv7dJ/MTv1wJsf4ujIZK/KnU
npAqfWVI8IGnKunE+WmkIqkKsAI2fmBGUyN5M4z2WD9KaoLYh/7bDT0J+R77e+9IWSBNdBGh2O2P
gz+x7S2k0GmM+YRhjasJP6OZ8rf5+rxDoKial1PO3b7j3K31Nj8JL4rgjKRomd8ZTUC/rL2IENzw
lmnTdUVkDfiftOkYoQFHXtosC5l6+/Y1AUlvbtj9NYGwrKTrmQDC9tLeVXidS2ICAToKSel+S7Ao
Y7x4Dvr9bC08KB1smsBSCTLdO63uYfCSBd+sw1HOQUOXcDHCOGmpW+cRMsmadZmf1w3mSrvXr57b
fB4iaAUyewTue/+OJS/GgECLBKY2iRbgmQRgS1/dSMQPw/q5YC+OBvNlIF4CyJ3y/7Ff7lA6hfVa
5Gh6My6O7zU8xEvuWbW4qkhmHhhkIs4Ri/T3BNy6rZIOAQiczwofpd2meg2vkg/PK4wG+VHZiJLJ
zXqrlA==
`protect end_protected

