

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NLuPKxa5mbHmSJxckEHjUBUOWDk7twAsALGLJTfoesEfyf1h+MyHFt0EylBuknot037Zem3a4g/8
zqiJpRTvDQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PZD2wWu+M5aw+j7eNGC0wVwZ4AHpsd0CPVCpF47C7xJo3X55KdgUsR5H/ybZtMk92enNjFrgbF3L
KLt0dXzbb93KwOc159Je5hTevnSDKsuPBBX0lFHiAF4XzieRUgqKA393lNR1oHHjtPcXU7UK0+IO
OzAzlRdUGjlDQbtNdcQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HouE4V5hA7QCiWy/ZOPsRu3XTzmc0wFcS7HgRKGHCsE7XwCF34feUK6Bn8N3dH2x37iQw0vfk66K
M6tHX6VRefC0MyimGFx5BhRdZq2+9JmDppfV1gOtGrREe6vR2IC/KcusvwTIiR6cQOza49aJQKA+
epyhS70PBrDp2VBILQDMeZvSj3XpQbsXPr8Q1JIB7enfz3ztp6rC/LDFPOPZe8YTRh24WGrzpXce
DAXUY9s6WN8OKURansZYbw0UNKD0cHLvro5mUb/lNTGoehE+Rw5R9VbAnGpd9pq6Xo7PPFVMpe9T
FezLXjjYSVXyY4UaLu9/mkvg/I686Ex7JR5c7Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mQhq1J/qEcykVkr3796fO9gQDJzaYdrlMC9hjsMGY2UKOKUbTtyv4tG77bM+PRHomfZqg8iU7uWB
GRXGd1YHbwBY/Wo99Etxtx46zOPIBoU5nFYOpTJ0bJnLbwgg1pXJxkzA4oOsNRCM00E9Tz9jDYcD
u7yXVYNO1n7TbdSWAho=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EIlt8tLrN8oiN0Z16C/INtbKo7UGBZMOz76+FUKU0dZcfTr4khTZ5FEXDc4gJZOM+wM5qSdRbQub
CzCPni3zASJ+ELeVlFnyaBW04E07carlE5UDdrotA4p2LXk7vZzLcnqW33R6DTbUogfnDteQ90G2
rsl4ouAA15HIZj5RFfE16KQtkxJiDGIwOrcUzhjmqqnH0+oOfSHDJeWV0IASEIzodocR806zCuhg
XzX3Z8z59bnwpkYETnyBEOLgELtERsBiu7XiRZGnW3iYQosufAJSskrAoulfqggYHW6NCOFZhGQM
6C95at11rwRxl3HbZnf/S1pzmZYljP0ZGBuLpQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11744)
`protect data_block
jewvKosrNdJZhYNFLFUIYe8BKZC6CVGaz62ivN5nRoVZc9iTivdLlr/FLoq494425OAthIt38IlA
zltl6eipI2FoskmmX9pP4etOOUN3R6tTcPb474w1OQ4HLYYA8406yx/FXDPCK69gC8H3qka5Kxmb
sNXsv+adygNVDSnkiTzwr9uo8xL/doZUlO63+v5iaHe2kEV2o1Aj1mOL5ANqAFdaUE9kuIOaMJc3
ZmyEZmnCc3EkzP79v41MhCNERnrNlBPCLecOaU4IPQkkFuC++s3aeLxD984FSE1Uy016fu6ISJxH
73sE8u4/buPf1EHKPzfc+9/D7mimXuuqwMreNV+ejpfQ4p3z8Kgdx7jb+VwJKmNWnZtW1SQE9iDx
F76YA2QMD4iKDqCZf4sVWxz1VESiruCzKQN0VvDC9VDaWBkz1IAKD/1aMX3IhD1tLaTdGPhBS1DI
EhnCEM0t90vRbzL3wj1nl5ZpbL4eOA1seBZY9DHjfk2Q2zZWUDwfQ4sJ1i8GmC7oDOZ9WVUwTAhS
CyHiElSftSS6kffr37TPbD9tuImZ8v+182nD2nCcP7Fev1Wkc5Uo8Zx9+XLiY6G0Bu4zV7IZgFIy
lLpi8B97t9KBL/oAFnivjhEIrCEk2UFlU62jcg0hmFLx6/eyqYM0ibfa/24hkLqiJ4EYAocMvIXL
mrO7rVcQsz0mGE7FS7ZbBz2K7QLC1zy0/Kwz1MMKYP8JaU2ET34RiOghrapQH63iwWxxTxJ4E79p
AldoWPpsESJq1piiHK72ryvPIFqtqapH67Fw11SdgsNqr2UxHt0aAxgoh36UC5lJt4I9V8pUgU64
Z4ahIp3Yk4uS0nuJygh1bkXGi78h7ke6Q0hSdoOs5jwQXJOb+kZon1gLZhMntzo3c+CwaESG4XMP
x1NVKKNmGTIMxz9koO5WjgG8ncq9ez0XELNCDqglOxAUtiIa/HDsnDu1aE9Y00vN3sbVBOnlY6v4
qmUQ4++CINklr/KIQulDWDf35ZqNe9A61My2uO2OCeYdTqVeMcWwi69eI4uCkRoH727Vrq/cc/k+
aYZi9ZR0vpOaoF8DTazezXX8X6BSNY8WXG1mvS+HgZD6IPXmTB2C0SyTFf72xWwkW5iRcz3qqOoc
GKzhNjVzec+2yrih/UGoZP4yqHRDRhfXsLFwEfJkMHB7rNPVyDc3nz0M9WlHvlw4z8nI2IVPyS9D
h0TWNcftSnDwm3jgdK6WzTrLXgg/1MkXHFPK4NMfatfW3v4y+sENwoFbs4VeyqMvUW4LHJU1CW3c
/aa5sM2ZNsBqmQ+R066JauxQ4nVDfvUJ3O8zYfOjtB0CN/gULklmt7l8ONdoVOpVAkLe0KHnZFE+
3a36LSBJOoAtWonUqYGE6IpLC+XdGSUtPE5FjZwHZNhGaFga9Mi1II3MvlK8Jt+L+2xUzR4UXVgx
hGdgHhJdWpASTKN4Bwwi7a0AG6iDBbT0XxmZ8bBDvO9WdWLbzajlXfY/PxhngKTmeemcubNUxM7Z
PYhWFMHXp/qSr/zHInJGQEFgzRS3nosa5eFYxXR6Xl4oBShz2pDQO955mDE3d8Z8cc8iAMXf2dA7
Xhm2PMvzuqwL6rxQgINwAq02ZqApE2VX52brcnxmTnWnpG9Sc7dQOMEruLfy+Az4KJICNOQSDiKp
USuIv9NCsNbInVs70cL14Khn7YxP/ufzG7iTcXeGbEs7RV4zyYZcJp66ZyPMlEPEtbno/hKP5AZB
XIr3VZI4rEkR6n+ygMxVEiWyz0KERvxc5PmSplQ2zqmVhP7nZI5MXPqu7p+bDWGqsNk/xdG6QKkB
K3R3AWZ4c5WMmHla31usIY8bJtvD4BB4499LNxFPGN8oRPL9r4g6RJ0NQKtyDeaHXYgPrMNL0V0j
g2AUziqfbanmkruYQ2RASZDToUXuCTTD3ZLyKBjjNBjmVcdmtpvqVu/7RTLo/RL/IwYT6j1USjX4
VmtsCwv//rCDowgX2ns9oeUcY8TzXQZvL+jsVRvR5q4FZL6TW5m9o4F6DYKcupvsFKNCgAEzwveY
y2DrxKtVeHxRNEBjv19S/SXRPw+QFzWXxfPhXO3y3S83ZkMVzfVs0BcwaEAtf+XwEZ7p8YbW83qI
DmQSAVhrSNfvrg/ughyZwts/fDEpjs7r3s6lQ+sNXwJBDu5X5hbLCQS4In6V9xlfqoRPv14lG4h9
uv4L0F1B8toI6uy9OukIW+mTszV0MtnrMbAiva17cxrGhWOrtx7dnjW1BSxkyax8IVtuaufaWRZN
N09e9eptMDZ813o4HQg5mWWlWXN6wSwRluVJCRT1gGW0bQSiFZ6SWBZKJKqHYKzYK4+alsfiwOkG
iW1ABwPe8BE/7DDC4P93AlFyOAEVp/2xjoF1rS4CUo9Lk5V3Wc5av1wZvrSkh+/c3exzaQCM+kUR
HIThg18A3k2Ptvx0rnu8htip5JnCqqytwahEpgV1aA6q6jP7s33Cp1vM4u1iF80hZVrfj/e3X8yY
C1F3bMi6RTjiAlbFJwrpuN+9dAhuob6cxvpvJBrXFJNaLM0L/VXTC7zbg5pQQGj/FWrfQyr/K6SQ
POBaywU3S3ts1Cfk+9cYjHOPW7HwCbBOkDAVkSZAn9gjfr78w2Itou8rX6maBF0kOMGAWHObENLE
uPZV5GFV0IRW4iOuYCqg9h9uifItxGfHF33sUit36TOuwHfNcVRLOALgzcYeqjiifBYrO4yM8715
GlU5Q+9DQ9OX7vgLy2wVtYb019v6N7tandIWXPFMHFA6q4dQZZ5z0YxQT6eykLNhVcQrT5AZ49Hs
xxb0D8lotb6fQfaeteUOElqDbN93o68FiTmr6WjW2WEvy/Kc1AUGJ8RBTRbPdIP534+KEU8SlE0j
JdS0F8EhlbvV6MbiLZQpgcKXqK17AMjDqAewA1h6PUA36M6+jdCPyeCubknOlcXqtUUPfpQ89K07
KxUx8qSgs8hXEMFTdCV6BDEdEtgAkB5FGxME5+ILMcZlAl/qQRT4PzzLg+TTc14yqepa7cBFBAW5
caYUgmWCkqBEDBY7CN5ZSozNmmVZ9AulVQcFzRZz7SCuKT3hm1uzS4GGE6X3Ym6pZ833mi4OczTC
c1cS8d+5gyY3IRkZAhmyOIcdHzWCwxQl7k1TKLuiY8gMOLEk8lVr+ioH1ssqG9pPI9albuhpRHew
xNuFRIb5jhbU3BpEPDpOnCEN7ULi/blxJl8TPqSjV51ik1KYi3sAPBIQE01qyLlZant3Ol/DRXUP
o7HqqZ3NGL/ipnMz/ZNILPxKZNjut+uSGHUBoYKEsb6qEXbcMt5ok7T8Iu0kPw+rZOLkzVYThJnT
Hi993ZtACVZYgPLpcbb5ao4z6Z3l9mBd1+O6BkWLXPk7jR3jV6jIklIb1f5Vda8Z8sKqM7gFcoqN
Ui8Fbn5k3gBmjGoKbMYyXpLDcbp9H/n72lbbkiw2rrFoFrrJA3qv09JGwUEpsdWF+YrokViRBhzH
sG7adXOb7vOlXqS6X9JacEEFO4BBxJE/Wj6MwC0f+TeiJg5FAAoVExYj8A+uVYZVpB8hAec4MbyD
/r+qR93/CNhTnbLpD6MTxKxFj98xeMu2jpijmZEzfIH5XYIdocuAQwRwrp4EcK3cWCU7zUMDxte/
O6u4AecMp6YzdTSOwKOgO0sLmdTfqMHyWQeoCeV4M5hZL7w+OuEFyVxeOnEywD3ZqP4xXeXs1c4w
vOsEOc6necdZLSAh1PUjfiZxTSMDaT5IFJTLlDVj0zszRQ0GoVbhX+5bi060wzteKttUIMLvG3GP
BrDbU4qLsBRrT4JfX0VG5q7zVyrUTg04jCMGnNr4FsZi4QboBblr9p7vajimGtT9nfuWuLDT1BAd
w3/KGvtquCIOBxw3nyQ2yel9zii2Kijm3t1V3o3fZLwL+WcBKlWF69tJzItpSUnt4t4dLJmIxSTn
sGmECoz5yZaQWHfVAF0m5GXkbBbBvVXd+zHkS2QXmuyC0zSIMa/+3vhZV8w1h5VawlgwzMqxKe/j
n2cYXI3cSjd+zSZu40nRD/BSUbCcNrGNZR7ymvlNV/3h8ERNvIo+vmnK8T/XLeTYiSV/I7r58Oig
aatM4OXMjVIQtnmR4aSW8aTV5lcnBvwEWAbCTwTMPnxGvOzcNx83gvyVlahkQRB6uQpdv5g8fCej
fS3FAYde4Y3oeTLZcgFaa9LwfotTv5K4kB9UFGs72xmp6ZeBKis2tmaVRbIY83BCblR+KiYif1UW
dj1AOV0k2xEyEu+3Ehkf5DjbBz4uGeoK2lVdbFhZUhSIlFRuiKaw0NqqANxiHJ5kP50wHZxKzSj1
NH2NPLmwy9IFbukaTaEi57unUKjbgTP1MpBxX5ZU2dKCvc5zQ9bxC/SFd+dE1oDugQ9Z/0Ub62L3
oVFuDhnJYZxrQDTWFCKUmFlAFVclNkWv8tK8SC1KNUvNXt6VR8QORmogtxi5bZYUhrj7yb/t0ZTa
9np4HRjrxfLP6Nx1OIytGc5p9eXv1rE082EQVtHV92go+O+bw6v+gvp6+mMK9/6RIdqr/1S3XOza
6cbIbH+xy4q2FfkDP21RejE24bikgJ9Pzd+W0+J5Fsh74GGqhBF4gY0AC/rC/6XArGaL7oIDKGaf
6gge6nMMErh/PPSnESpmGBTe/21WcELNGCIy949XIDIVu4Nfk3xn9hfqW0shqBpiXwyUpx1IOpmJ
Me/3E5KQWO3OVdyMCucr0mrN0WiLI56or0KAOPVs+UoNGqkElhcLlXnvLspIFmxafjx8sN7+BC/d
pvGNephDkFkmawUo4Z42L0anH9IaM4cJl+O7j+zTWK8+S8ZLymHvBi1A9xd9IcIMtoTSoHvyQ0Uz
W6VAoDP4S6rd7IxVNdin7xIG7ByS9IH9mGco4U2n7BU/YycikRoKpJhB22XAJ4hIkTA6CzBYxR9H
TSnbLCQ8KOu7kTQQZ87ItGgTxyOR2f+9A4MF8adOxiVRrF2Dsw5lJGuDnwuxl/BXSA4az9N9Oq7I
2duwqZUAAv1NhR8ayiJU6s6t1gJ+43OJ9uBodFGLgiTF82TxSYoIij9Kkktb9iFLK6u8ew7emUXL
GmhB5snF30WxGGjsU+th1epH1qKFIWAJOnImswv8F7DFEMBWRhxtON5mk7dhT2xu8coWIfwX3/3d
c3RwYCHEcVRBSLbvqOl8pcoXCzLWv2iqcEiiw7zWqU7ieWn+9psK2tAsaVPeq3kWpiPT+qHyhzEs
kWc5IbNsKtq0Vo0cdU2e2RLyMkQrT25dj00EZ+X03gA3vFSQAf3Fs7PmU6ftJ3i2fIX+PACgnLiw
1/nbgz1YhJ5I0LbU0yzCMX6Yfg6cfVdoS4zR64w7rO1NYD9TGyQAm9FgxtgyseTi8HZf4YEGM/s2
rWpdL2AYVci+TfQBsDMERNow9lVqmof//8BYJUKsD0AySpMBj9nhtSZhMOsjECaxwuFetreYc7HB
xwIcvQPD30F5hPXdhwIjXBaaM1puJiKovo1+4Vkzoj0DVQYMgBdGIm/kAgQVvU0Yg7ucTR/qmUR5
gthR7SGAt8jEnIxSKvvNDADIp7qwo6T7PO20wt4/vbGJFMVKKC3ga7zyNr7a8pgbQkMFFm2a4nly
3bJ+ILfz6f08NuQwaZbid70klLOjUkLsICBEw7xRHdn9owwqnD3eWDzWZtqTrhiTDxAiJtu1cVgu
qMuQlnb8ZaDSp+j3fsQo5QjEw7h3p1TYDTKT2wqHmDLR1+S66WCdxxAAdcEknczHRCk5cv+Rc8uz
5grnKXVXZsPyJPKjyT3flWGRah3WCuD3q2h1tHaX1l05fClqfiShDr3ESqtPnVhpN9XScrXdPZcJ
w8lxWaYrPbVVVmwXcoUxyD8gHtJsxOPFwIjn2nxBlL2E6Bdm0+btYvBOn7dpT7Kp/GDgOUrlcWsK
5DDWfsvH/xDQGqCMcQ198AoGmxPPGHArnDqfw7vK9nfOAytkDBDt9cyfxQYV4OAbFF1+wxmVhYJ3
yTX/BBG3Bqu55bNvkZetIQdA8eEn5XMJcwnOxUOBsIhRJ0RnGtS5I8B1C61mHEsgshHsuRdm1H3i
GnBkAfCaKXhUjjm4CUMhoElO8Wryi94JQZ8wnIkIP1I0AsqA6RD5rrjOeGfFlPnBG31oEv9uCox9
ukAnZyVb9sOf83y5PPmH+ZBZzUBS1r07kp39Ts+YM3U80t1rDq+uUjbEK00dmrmCPPWx6NgLPI9J
Q5MfK7sRh3kZzbc4PbtimLJUY37ZvbOymfLHxJbxqSu2tvQ0TL7N/7GnHc1zAkkzhkH8qpzsSyXE
UAVXHsi4C221zWMA4ELhdBm86g5zhaktZDHxL37YsXVezOe64qnfrwEjBG3rwwjwXGumyF3ZNFZJ
b4FH4OOKe11R/b9qbcWKUjs1TmbyjW5TJvi+A3CFGivYwPNMGIIN4Fd7sxwS472MNFDUqanUMnBU
QhvuUY3Ya2/Av6RW0plw1MXXQs7SjEENtJgpSFVUGgiB3xPzr549gfmreoT21NwADO91Le/+Vz02
f3GMgMjmMwLglRYhesYYUWQTxrNdlEktOaokry+kaWIyVQq0fH2CdPSkUlZVb63gYjFS/GwlW3Jx
MtMP8ESHkOj8U1tKynzxhlnlzKpb7haLDaGf94IDe2PVApJrD7kSaSpiov+f1Y410Keo3BRl8Px7
SsfEOzQEAiJuwasFhA40Qo4cjn4TKxpaFEAWwFyR+UzogbEn6lNLndQdnxRUgYoCVIqYYNc8m+lX
io6aL70gmvRjCv0r/hSfmIyz1B/K8oes6u4Fl3a3Uizogo2mMDIb7J4tjvxYZdyNzi5/SUktOXF+
v2k6Ed2zEbUYBDTd12SJO8Goync2C95LpG56yJSDh754U4k4uCD285FulvdXrCkOEm2rAACzT8Is
Nms3B2JEDzrIDTFoapQvw+iYHIznxKbPtNpryBOvkbul3Pk13b4q060EIUHe8l5oH5vRbmovsIcr
nYGkceZB9PERvrxSfhncFccUhIfLNaiJX4BaRMLX+B9Wo76wg0PK+ME+JFMtCpLBymfnVgJIil/U
3gawg8X7tguvKf55sq7fvHp4TgGCsscE3cob26SmkLByQu26h8LTEPxuMfwXCoZi86zbCZAFk4N8
xSqj3csC06a88TnzVQ+cV0iNinTobXAzNf2YDXICeYBCiB5hRfzkqoZH6uwT/dgYvBTBabpCJJq5
7JS9lsQUPs0zEILpQmjAkPkCeYXBJS7P8JpuYvlC1RwHmUs/RKOnpsN5XDHYH8pjnb+KH5mj6wol
qCukP97bZvSFriy2C80Skk58oB84/M5ycUYyoaNUt+2P5Bl8PR4uKbqdgCuXoAI9ggA9FipDXbqD
8L0aREUVA6Zp9e7Ml84H1gbVSZh/iRzH0FhVYWJCk5TWtMSj5pdVOn3OBjnx7r/Ih2edkab+js1D
lVwzF1l4NoaYAJUd6qcPmEmcsZW79K3lWWTbb+SKh+qcbCLVldKPVIGqYIFsZ3orXdkdO1VzZlGS
3ajcNQGHHd76C96iGQGyx+bh48L9VfJcZ9RbsbgaB1M4bwVKfGa/YkrTlwttPCkaJHEMfwYjv/2q
2Q84UZklPJjlsJDVnGUiIue/n6RPxT7dETe8CG/bdO7TNIj0NSdDHFzh8T8PDUmsgAFoYEK5oPOm
VV8ETU5Mqwh6mSf/DnKSgwQla2CmHDrS845Xo1QL6fa0dzdJsaAUN22vhcjkqVm9e6cVNHDsb5fK
Ddq+yDf+NfrDiCc7ySF1oaDuKsEGJ7UkKUv5WdwIJ2H43LhFgBaUGEUiitFeuWmRcSTEDptXPIK7
20oYC1poLNEpKzNZRQLnwRX0H71HiXrrvwx8E04gd8oO87sfH/3QkhNi1WP6I0DndGufE7JddRLm
SxEKb9yfLuZNvRhIflmeGRHPYUWFPKQloZl9dGWrzNISD5hE8vIv/E+QsETfp2jB8FJASzB1WtSI
HSQhmoHR/RoMUI73KWZTmsoyui47sD+KK2zRY9nW6nb0MwC9psehbYVR73vjgIoyQHBAj6t5yQzd
M4rx3kp3Nm4TTHB0gaEyyBRpRsUJA9OFwl7f94YNeL2fGw+JJGhaKBHk96fDcjiAXbiAy4PFkpJ6
tLcJWaNnoT13DWCe2mdg//4QmZviXqzKDFzRAiG7I7Mb2fvvmNg3qHhv9/UI9Zbrgm7tjAwzN1M4
7LzJBt23j6KF7/nhpCbKj55LYePdyHCon3JS9THygBaEVDOoq6eaQjAE2jXpYmPiFB6EXrWivBai
qdlrMPdPQb2PBUOSJPrVI8w6Fhbvuey7GAibrQHS465UnyblvhD7BUaMOVTF644DOmlpfO8IEFgC
xaqbJRT0lV1OxotwCAXCaJVe1li7HaUHPqt4JsFovk1r0IQNcm/xVGe2ernh0HdV//+kVah3HNFi
T1fK8LL/97gwPSCVPnl2fUDlnfs3hQ7jZf13suXeOZGeMXAxaDUxIAiFRCfeX6PzypT6W+s2JQBj
i3huAIUMeftAqbLqt/b+qg6qPClrSma77Er1cZoBMKywDftLtZFLs8N7LCIcnVRAYQ8RmOyuxdaN
iOXDAG2aSwuOB/uIBJYOxgWq+JskuSBevSLABihqjt7oH5CCBOOt48DCbaG1c+vlrybrULNkmjiZ
E6UpiH8vKwxoxVmBGp0YQ3v51IFjV15/AAhhDpHcWrvDGUDiT/OmNsOF2z/8V1xolllV2LCAzNiC
kvbluO5gKzzaaDthlYe9Z/5LzVA2ByMTj/OkV3P7DQDeZNKGF0NV3c7hbWgGvJCO15s6/OG3jCqE
qD8pOHczLHG1XTtIyk4nX0tsKhV7NpqM1hV3Zqs4zqciMOmBhITLZZImlcmLs5gTvGrhit/eRVsg
RM7iB7B16DFHd13zXQtSdVUDEfNVPvgxLUWodajq3Odn51w6LHOnEBlFGkE+wxl+q0zQ46vKXGLo
7wop+VlreyGhKdV9PEIU7fvt1Ca0y5mDqC44R0TevKjRl81yPLnnQxjXOFXQaysz+e5Y0JI4oYV8
EAGOK7HoDs+CkdrXuaeZcZZQz6lJ5Tj6ReIVCuql/BJtojkR74HMLbvvi1jgwY0BkGX2vB9DD6am
ZV4QyNta4T2dUhm54qgOTifYqY4ivENt4WWyybWwjBexOHWxuUd0FM++ml+1XUxULrK/+nPcuKeO
OOTuIe899BnlFlcUdMY5556Y/pt8cqSyW66V4stBAuVBm3IfElN/mXe2d9dK/eoNAwicvMrvC7yF
J5ZKKD2RWiMWalsqPUyrFWm5C7R3d578H0P9eHTBkvy6xKR13GbzMT0zCA+Q1pIVyVS4uEtMUzEV
mR7X0Edou3gbNQzaqgo+9elDRizmmF843MHCnKiDvgADIihtlWvt5zVMuePeVN3YjGRknSV5Uzi+
9wJ00boOgtqU0AbFzXSRrKonLNLgbq7lrwslgeJXuEriu7bugSxXmO23LqUBROGHsBEZDr2Zq1Pj
ntudf7X2JPnsiQuXyk2IKcnOMz64X75ohgQrtnBE4dwsTIEsKaby6eKey3Qv8MBK+BNBmU0aVg2M
jJWNiAyzFeefHAHIG828kLZ6j3j4BikAI8+Hx91Bq+EzGFtgtS5RBBrB7odpbcvcANzoMzboHv9w
I88qHBfmfrETo+wO0aRbmLkg67m31XqN5b9De6lisiCrLJHlycFAO1Oln/Sg2tgvlg8/pDTEsAWw
ht0bRA3nvZTGg4TdDAl52jx75LHl1KOaxbD+qW6iH40HUUXO0m3V4QgeKTmCh/fNmOPOl+pj6+hC
zctTZjAEgVPwkz0A/+yYhHzeorZ/ARXzPJdtHKchbwmwhdRu5KsUPJr5nhmpZs/MJ1vV449shSHt
xjR0PTCybRhjtX+DYTX+plIpRYcJLybA4lwbNbn00Id2gZKahxX6/veSHhStCGJgGjq1UH8CHx+5
DbTC/TdF9CJVoL8VbSCKTLoNY6ocoD/ARxkULMk9yC1ue6hejXxdB6js3YihEtSNk4DM5nvICQED
yuouLcHOjp4yr6/r87GIhkF+wYjNIQJAEAOSlHXQ9FX7pKKnrNagrZqv6me/Ax3N8rvbhdSoCVfu
j0Qjioc6MMGRDgj1NSS36GzXPnCg0tpDtSbuwjae708+CcQQSb7uVPVVBsPVwaYkEt6hzMTrCU/F
d60pNYhysMsUtpTJBNTWAyhqwEldO1YNiMSOXNV3FeZhTwxYlphcciSiOG0l+jwuqms5uchGzJBR
WfLS0bLN/dgxIR0MiwzvEqnOSKwin8bylDdgLcjpmAJ3nlGBWifcUlyxmX1Xqp0hj3CvvKr6VF7l
qfZOh3VSJxxe51Z3scmoyeai+dOgnE1xGYjJYXYdVBqw/2CRGqgRVWcfNq0/qS9ypiDZ7ZyQYHr0
k3oPXirwrMvvoVGanbJOKk2PWAyVaICDK1yfHAGlyEHO1w0F7LVJ9/cuyo2KqQBrs3hkMDVx4w35
egGFh/Pj88am3muv4iAcgJyL+HRD3dXSYysHfVTiu1P1NuxnHGqPgj/0Br0bJvEtNt1M/9dykAsR
5k5jeFEEE10wdgkpNt/P5kAiUPJHFmBPse85OGpydaXAzFRTso7lMElG8Rd7QqTERVfjMZbDRLkJ
xveldcIHZPhbVuEiXMQYAVIEeRSA2ZfyMKXTtlCoRYvBvXm1cbdsrwnmbMfiZfNjbiBxBVfL9K+p
wLXWIc4l+nBRuUwZx+x4O5YdpvhnY9w1bt8KV5lUWc6/UAk8te4rxPeFBdfkCh5pJkT+3QasNqdo
hDnepKOoHzsI/64fgddrSGJzUuL2v2tGbAigsDa1a/fEggDnBJhhWQtbe5cE664uSG84RqRNlNQ3
yv4LETd1PFQc9BMSeqZvZVrJZFRpmAIPI8Cr5cdEPHQCKEFwb4xRWPjcll/65z/N4cZo9etkl+GA
gQUfB45dHb2da+PUPnuh6xaMhccKyRMdU+j93o8t4Vje/dXa6NVXmfgrx5BOaPBxj1TVC1zB+fzg
mNqUStHepluhLQS8XjAVlyDEV9+4a+NmNG/oSqwAslD9prBz4JuLwea91AdHW+cGLGp44bAdes/4
NKu7ET8q1ME91WUD4GyOjt5YZJT0tW2UL/Uda2+iSk1rqDoX2kknDZ6+Rvq9pK+H0psnrmuIgvt2
maqAwxuKvMKzM3m4+uu2q2aEV4fszkJLsSxPi8MweMH+ugkIIKpIX1q56Ydaui60H7+0I4liC1QN
qg7bHG+yWZnLqyEF12o9Osis9dD3iZVI4pQb4+T30SAwKDQGmonP1eRMbaIKHy4bAHKSZtK9wVQm
1nLOZZD1mIO0rvxyQX1cfzuxKiL6CrJnQcXorduWy4mQS/lVQhCS+VpPm5aKjAHU23V2KWLufblg
tDvbZM+O+j+l0eZVgTJGfGq1E2FEi4JdKZ7yyQa/IT2gEhKCI6yhoSoRv7sEWOvbU5OGBhHRCsAK
wUrfK/qo1at0YfHxwT+yFDqz+QgSDW9MlCTPFKQ4+Y+psgAjznPzqazM0fpGS1dnuNDQT7TY0UvX
Z1oGTzHlP3t2w4cdIjlLzpy0hvQ9LC5I7ICCnDSa78CsJaWx7CQEQNj0x1WrYeVBSyuVeArfBPRj
Z5++bBAMvZYuzbFeQCJGSxtabSp+R1yZo2z01k1HKQkF00HRLpo5LNpEoXQVQzza/FvaHVQuZv0+
Y4B7WObp+xbdCiutjJmLHZQEWzygqRIxnAJE3W7dpM+qonFHJkgIcK2Hh67I3s8KNLv4pVv258Ir
N0teMlW0yXxCWDJnMV4+/bpRpouGJv9YTFESwLLO/xwHGNijnR5sOX/XJF8EXn+WueOpJK61ETsR
MIJVuThOaoptRK7KfxbfD1W/OneSwDcEtnx7ABgoSM12IOKEGUGm6gax6gjHX9UOdWoMef4Je+1q
l9nDlAVZa3r9Hm+oPoS8VwkSvD6+sbmTfJS57H0Ct6+ymnSvvxdN+j32XSWCAMOuocSeK4Gd8ZDr
tJ79BudBWH1SWukvcSeYeC5zZlC6A08jrwrS81h6IAKDjAxtbYHqc4/HDYQF+RdX7mVtlChRl023
qhAvcRZYP3ylUqOVja35//dQlnxMvBzCIkXuE0PLK3GNqXZP5j6jrfSj4EJ+4PHqZX41wLBWpDam
7zIqWFiPyf87SSPo4Eeszwdbrmu2zcRmszaSM2JZLcxICIu//42YrB/JpHAJO5pR5lHRWgzgDG2h
oN9bHFGK9cwHPpfJjwIRDp01vK+qSQK71Yo90B0Y7Z200bQT3A4uF3M9JnheuG2ZxreaMoPY3iAO
6RpIRXky+rTnuvCFWDTYT3IKfi92TwExYB/x8Xw4HL9ETjJvf9CFdiwa00XGhbfhqFN+8BEPxxZJ
vRTGDIDEwuJ4ekR8KgNZTNt6Q+r7YVhdUwsTob7T+wT5dlU70wQhPJqGrUlZZjGbnb/Zl0UaGDml
LFwWIHCzn6zeuDzeVzdh8xum58XMjJKz0PNun5hLt3GqiKXv0gCCmwQL4Rvw2szx7CYrLzTIvKZy
4oXEgTM3cBEsw2wL5HPu5Ipz0VRhgyZh9G+FZlWoGnrgAAGPUOlis/xV4khfEqV4vNPYZiT/NZUI
4TCVxVFx8CFPWnFhAGVWBILcU8J3NHccXfDjh9jAnezW6PDCg81i884yO5jOdevIZRf9q3GqsuxU
m1vF6mmvYQg/ATU8+/4NLGsMtCNTyi6fOrgc9Y8SJikZsmJtfo/KYYl/h/k3qAIXivlxNNXToY1O
/4sHicpsJJIEaRVmCk7+RvLIvAATobOTNKyGB3T6lXZEiezr4piy8TJP89ugNU3CEXvqKAmHEMsD
3h+PQr0mwTWxWQERILPdzr91IdVWntzkem5bdGoks2xWK2lEO3fMxEQ2nvCFdM3Lu1OTx7ZpYLCJ
FyMmEnbe6dqIyew2B/XFcpGFnAlWBuLR+z8kWXncK9i3ilqSX+9HLzUNkRmDf7QII/wbZjO1YSnK
S5oXF+1hwWwq/QTvK7ASJsgp1/8EOebL2TXaMtg7hwhvO51NzhZUNGNGgooqPLlee3gPJ+QMQnga
a3bkeZXIMyMl2rN7oF1WvkGgkr01BbQbQqo1X/5+KJ1EAQMMPeuKhCs0eml0YQGNfT952rUWS+Sq
E6qRrROy1/CuIrUW4/yF/lopWTvGJOWaik9DdrigHbuOqBgekLfNBuaAz6+hiKJCGZfYhHYw4qq6
+CDaalvKWcH/s7T71fsvdVqHvRpGV1LF23hqGC5B0TGtSIxy1VtEQ7Xh7KOV2XdWxny7ZtDeiX0f
Bs+LVbhoWiwCkDJShs3Y2Xmc0G8tjFn//5huurM1F85FnXY6hRPrL9eaxVL6IdxaJfjxGamXCahS
qQLjBQ2iS7KwTIrSgcyDI0h0Kq7Ve+0d8/FBn7FrnzfBJdWEg9wpnlTZ0C219L9UNJTAnOdmh/gJ
YRy5MZrVM+c9Gef+L1JJ+UcuUh5wBJ+i4s3F0MRSHScWcdiTUhhcmeUtjGRRXyhCHHlePGLcSXqp
GlkB14/DPv6EE5vGg3P37GJdmWn9D0ziB+VwZGhuA7UAhZToZf9HCYrpjmIBCkLZfpd7JpxKqwnv
7r0O42zNiqcQ6O33PrZyVG/M0T894Mh27C4HOIUaRLfp7g1bJm8Rg1t0VR0DmcTwUd1+NugQZYKf
Aqv90gLSwSL1ALeu0R1KW8TeolKSM/5qdoK+2PSvmwVHPUoIRvJWOk6xhtI1gcvwvsMFL90aHPkX
G/4YmyHtlMB/u8TZXxuWmjoiISrOI8bEV5PAEku434NOOXhdgxQ0VOe+Fph/qGiwa7sSI7wPStCO
H3jksvp2JZzvuieoL06vCEONH4YOU7f3B3Cz0hWtE/z5TyptAx5B4ZexIZM3qswkzqg9zY+FW9D2
eN/Fn1GzQbGiM8/mKk029TWVozuZ03osv3sMVG/g6jJpy6ghaqgf5K+rMQJ9lmfrRl1LciOQ9SGj
cHrrVS4gEVhXCGr3x1Q0VyAkcsMq4ySLmZ5VLnVWR6Rt6B69eUpoceHM8xQyLVn8U46In1c2hG+4
brqeHbl+HHcA1f9vyKhS6cNTb+vF8+sLhNlgH9t8MtAbesV10PhPh/1zU+8JDSvsyU8CQLORHFOX
vCsIMenr3U/HM8ZrJA4KLcn5AmXy595TYbL/pUMvzK7nuWlOqHNBAmL0h/B/1AkbiNEeVy9u1JxX
lpBUlnR6Qk9vvTJIw4okH35k+tjATnT5YYrd+u2o8PFNe45T2dafcOB7nNDp2EMUGpXy1Gt+4Q1p
JN/T3FE6n7NHa7KKchjGOkFwI6FRDUpk98SVKXl3ezeVmdJs5EsiubRv1+AZJUDg3s2cdEiQ5cId
82jYwoY7Ua3BXWf7N2VWchIlrWSAehmEuxBONh5BJHbp+0VZaZsTIwyY+JZbQOE6hIAi2bww/0Wd
Y4tuiojDeRtNT81exPegvFM7DR8raRYK4pn3PdpV8xWhP2UHA9WzdJUxvuAV5OsANiNhDXUukP35
uwZzFX0dbj5n4wZgV1OWXSIo0IhoC+cTzji2BEZVUOaIDath8ePleZgY1EKgQelV8y/I2kA7f/mg
wEvQgXYSYYaEFfprqWmiShz0r5rwiCkGzJYC3PmtOC+oPNJNtsNAmepwVlfQfByOnIvHNkeF82Ni
UtfNtZsK70Jy5u4wxpOC8lnhLkOgxGtRex/L086NcgrsonLS/OPNsSSCM7RAizq4vppE5sJi+igI
UdDLqigNa9vDWa0lvjrMu1ld97kf/KCokzScWtASaqXrdRQWaWfjk5bKcI6ZR5k4ee/80GT/rL3Q
FSbH1NGArNqMjz+a089Kw4vnOzTY4wAImisfo4CnAvJPiWZ9WVpXpwaRlKyoJree3QXc67no67QI
ch/e6T/Q4PwC7qJAKDkjQOIp1w1NZV3cl22TZ1TlavmbQauVGrRPD5Vdja+b6c3w/qGxi6ykBeBN
lzTiPY5/p+4QSrlrE11D2zrCq1SRvkhm/U6L5LKRj9e9OTIzX2dPc5M4acck+p2LKrL8JRDSQAVQ
NyXt7t/e1d8Ygp0Hn1e7LJsfk9N+MHEdVsWCJtcCX4MM2nqxPdQzLybl5W6y4GNd1L2qk+qSKYGz
Zlhqv/htF/AoPlGCA0lzdyNlDfd91DJveO9hnUVjTq9wM/q3ADcOUK384XCvOUzAP5JVUDfqrnXx
k8DVX5pqDyQ/hXTXUJdtjvNlD028teKgO1D4xP9xn2FPs9w/Tvzoyql24sYik1t5Zb5+zfqPkO8Y
RW4TqwkqBLmO9YMhHzyk7316NC0xDZxcYUkf1QAYss4Rt3eux6xBnRmYdps+FQs6GRIrDJn4vWHj
E85UIRXiVA7/WY92s+YZM61PqHP5Zzu2RR4X4YcLBdNFRqoROT90ixaIVaZPxcyIFEFE6vTXAHzq
5kC9JRzFxtF9fR+Ro0HOFtyosDqbQPnXlME/WHtE7fa01JlSVjZJ2suyQrotHxJMaq6kAnZg23BA
JYjETGggZX04cYNXhK0eyH9nlX7AQvf4VbsedrhT0X28/imtBWQiI3KQVgqjAgA9RzwoB/+P2VO2
4pzoO7rQAnLRRkBBaLgd52YzwPRzcI5AnBn1Voy8jP6Ai5IQq6mbsPe+qXXyExA0BbZV8ThyyBs1
jFU=
`protect end_protected

