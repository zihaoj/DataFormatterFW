

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AxFQN/XzhapwiOYl8zfwy3RzY1FbpV3RUPtypt9Gb6JkMkjIFIEcJns/v7uhf01m7QjiIwCR9IPR
MqvLFJR6yA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cv0WfVYQYq9xeYkhg5SzPGd8MXWOq/NS8R2LJmTiT76lT6FCRSKU7qahGenfPKhSt/W2pPDxOnwy
QKDLsyXq/6RzO8X6wo5Fw1vb5xHXW6hZYtTdZ2dOdfgdUM7rwhSvape8RtQyi/g2wgTJnO5P622m
6KqxQOIhyi35BIQat4I=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
X44v/UcBnQMWhqI9HgQoPEjsAibE8yDRkTxDok+dtek8+BA8WbfA8n2Ea0ob8R8z3/dyix1MIYZv
LUBtPOX7DvH005rnu5HZln3SPNiiqaXJNg112ELEhGSVwSBNaH2ToyrLODgP65KS8rHB02QeUy8N
A92N3s1KWGWyaKMa57pYcKbFkRub4vpUtgCMdexD9okFsG0CsKo83OoOlUtj0hwvpEW+Nlc39Gdu
Z4h1hX1/bYdX6HJzuJBY+x1ceGcs+uCK/YxszJL8C4i3EvMeUwbnXlxsqcFFw11FZa+zbwEp+y/6
96KWDdCB/sJRXLRVs2KrOXp2HdKMY/LoFiMIMQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EuumDHg9FSJKKyWOGeuz7PERXANvej5/+QwBuFfJBojZGr5PUCf0Vym46P8lGXMr315q/N1jyCVe
52ZuI4uKZYzdo1jGKNjaDeJedl32XB3+dtKkpH6d7byLG1a449FvIoNPbYmoGtDQun72ABBd7Zi3
MED4hAS1kJbgwpjXowE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ej1TiNdXyh47z32+4VcSmxMcOknMBRJClM2CA+BB6CSKnFVpOPCmUQGcvJ1gEmAed691xCYcirPN
ZIywpNAGfzwIwwrLwXaI6gQ3PWNLJwLRhddG1Qz6WwOi+TgMRk5QT4Cke1emGXrJROhVJeUdIMPb
j28cFJFHrvjCHikDK6BQowxG9jnkLPp6v7R7j2rGWQAruTQwRjAVIgJ+yOqKxMCNqUJAo/h53qy6
5fwjMPZmP+ItP3hzRa/g8NiVLaE1N68h2W3TPRwagyS6s5nq6gUzAV+F3A+o7MJ6fy0PxyarNQg/
YPsgtikt8X8TZwowoNF/0mDybXHZv9u02Uwl8g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45264)
`protect data_block
l19b9NNFlpeRYFBPeQemw9C2SgCJ/NxHMsDgO+Whi2jZyMds9uyENPmo68q8EQhWCEMefXB/UeJ/
odA4GAM509a3Pj3O1yeF4EsIRpb0qQnDqJU/SFFugw2CxVpJbc4ICBSKOGbVMH2rpF1gkn7MDusR
HobYJDRoMqhRvQYCuV0E8iaFH349kNIYzTHp4arMQBoYudkz75sdLmw5Msl2nv/y/b74PqOwPlgL
RIgv3uR/udut3SB9Up9QRCGRmCN1+gC5aQ6w/YSQddX/YuBWIxj1dT2szPe2YCwomNB0+QBcMk8X
K7ubpya968hJG2FL061QdQJIhRcuQ9sJ9tL7MnOS8n35uIFETYkhcqiBNNI9n5RHERcQ+qmazHPF
POZHXnRezCaxopauW3URBFNwW2CjExWyzYWnWODVRLpi4br8cEY8SKXvwyYarmdwk+2hrMImH1db
Nppn6LcXXbJEPTK/dzin1popC2JXH6c1LKnIQyTJzI6NyF4UiZW6VHP5fMphDtpb2RAZGDwchf/l
/uzspmxPqjrrJEPd0E8UmsGNTHWNs1GD/EChsP7V1HdkbVfnT38kWQuYzUoCCDqbUsH+8KT9xieU
MfSdXYFLlli1hZVyBXUvghX+t1L7IWzHhDTVTAIX6JlS+KWxTXcyAmwORHoru3IEcrjbzSXWtfY/
eD6KWX/Oh8wbIcQcgrG0g4ENCPdLlQ1m/nL7ZNfPGE7gyeEH8lX4/O8emv6kTWvRvvIXeowiKq1o
SnKrf3VLSf0o/lPqsoqh4FcF8YFJt56tz+QZjjklpy5JPawt+e7XNz2B//ma3oDc2tJS0m6r//OC
LPvqx1/83kJmzb8MpZHIg3J0bMlayG29f5zhmcRO8/BQOlL0CB5Sma5n4x0oHKNeW6CgAnVN/Nnw
nNEf5vSCOCQwwbOAkM+vKwPy4KY/eB3BFuAMqhRHYjPFILOH6THeEuq2ViOttKUCXgcN8VqdA2Io
FgEMVZ39vlqrO1Mqi0zVeZ48nHADK6Y3tyl30/XR90MHL93ihgCC0+wNFBTyN5IwEfhB0SQL4Kq+
LIP+giZW+llqAr55z/BBIi1kpkA9nTgapABMELaoTutZQwxzfDzFcjsxCX7pKlCmKIPheXAbzg0e
WHyDgKIXdQArMUUAVnIjXSLhjhCztdh8jPHQgWLZAsDn/v1rkVqH2Ni5sVj8ArVHWnmAEQKVJAyD
RIaZjQYYut0UNiBk6G4RA9WNqJhPn7MQo/hTY0FKbYGU2umGZfLLdWDOk2H1LMCmTJ01cS5kufEC
VgEzhu1aPRCIpCb8N9FPh/N1vgmCO4dqp8qHbC2GK1JvXK7/J4AAyf3CzQnyRAwADKncEhFnKpWN
vwF+jRTkUlALb35NAiLkSSzft+oIpAHyxwX7J1IQSgT26hNdMfTf/KrjZZ0bhSAvyJ1xggzfQvja
O4eYOwT1Nelpx7q8etbbjOqHudURJ2JK/LZoE3LjIdPkw0q2uZuhYWJGw8iiKzOg7RPrhtBLVT2I
zWR0RrQtE1xW5RXT6ry8z+HH2Ukk79Xw5qZF260ognitEK/SkgaUToJR9c3Fb+XNuMZ/lZCrMVT+
LbiTAAJwbsW9sQNdUJA0VLUR9XOqHH4WQtd2OYiT2qA3VQui+bTrWJML2fRrbcJSydvJylm7UC+X
SainRjqkL+rfLIj7bXHV0om8CpEm/FVvOTPKw4WcYkkGMSPurA8vZVW67zIKtji7bwg9VnfDfS94
vy6sWcD3jr6KEHcUhsUwKoX2Fu92CwcBU32WypkTNNGGvnzwgr3SSffgLpwVcmuuJnlgthu45nRG
Xa9BKM3W5kx700YMoroLWboDuETanS0SoZdUsPBrBPCp8Nf4qEtJMMtsV6XePWc3i7shleap6xJk
i/FMKKYBZVx//lz+98dV4mPd1hxW6qvB4MQyO4zBonypNj7y6Xwq9gd0AbNRH2mX5ELj4qEkNpn4
ljygjbOmcOY0oKFFor6FOJbr9K8O97sMYO3ug3X0HQlE6XK/S0Q4u7DawFm6rQwTlUExIxdMURy/
n5zV6XtW7xAbCIGkjoD/hZvYlf7SODN30cueayRkxgEc7E6DjkxTlFQ2Ytil+bzRCE6hedKG4b0Y
Miyzh0HJJoGdAA9eZHr8Y7XAsy+zqOAwufTUC+XRD/ova4s4dz8UYA90v0Q627+nRiV7DWT4FkuO
K4UXNj81u3m89pgQvfAMvzHFRQYn62anhT5lNGncSfLrY1PUT7X2KB01LgPejrtXmfN+mxMFldlW
Av/GIWPPQw7PnO6gfETwsk5InQ3iBPUmHdnSCXVLuaosKoieHSp3BD7UHyfHwGcEHD/vbqYl9WEp
/XZ09QGMkbyc5SwXIEh+vnb0d/4dkWDBGO1IusjM52Fo3fFjD/J0Tz7gX9CgDh9B3RiAJ1H8xiUz
Xl9w9C8EDRLwcBIYyn3bmCc5WszzMM3uFBvoj+VF3IYZPmOBEzZXBQEPuWrmy9MRR6vTXmLO5W7P
55XP+tMvz+LzhlmeH9fJUtk5WF0tuZYmZuxKkNrhi2hJLQewtTWaTtIZKNCGmjMRziH8Ijq0ImBw
vYcKuLqOTUoQLdUmB7U98XXcmzlUb6hlfn77vgRX+jVOAKZVdxXk7BFkvtbOA6VlZFMl/JycMycJ
zVkxik7LqEft7y4D+9U9yvcNfeckJ3oMrJlBHuyFwEx8W5NMexZfsmwSyPLf+3IRr52Bah9k/ivY
ZsooaWIiRn1IVpNJskXJsEQPTYw+Oic99UAohRM17vgYrlUIjuWPDBtbUJTelqNDacY2K2HmIcP5
wCQdMFEicVnW8CgYihnbqnMxSOY4pH/5D5hgpH1cQAzRBX2jiCBAfQt1xALN6gmhT5efNauM1Ipq
wVxm/EFMy3tXDijfiygcC1MwMD0ctL4cG6G5bU938RTeYYJUsjxkTAe5kdrVw8CcO80buP5nHm5Q
Q0aFIMZuGPM/2BBPMU5w9P38feOOKEJfonM9HOpxEtLtTp0jE/FXPdwQKEX5N5kNacFulepdP04l
mxPsV2LyDPeRA8CGbWwOJzoCaldA9yAhgHQesf4da7NU2sgOZjZ1eQGrnpdTCYSHHly5TMtd8Apt
iyqSVYRoUypOqGBwa+JwHc2l4KiCJudEkpJJpetM6A8fKgy0+GHPibVAlMd3w0KphVU7T6NO9SF1
leP4G8Wej3DcsYbIvG1HhWyN/zooSk6MRhf9qWZnE8gTnX+sGvg4Lt8DudU9TbHLfgwGvQ418JqM
/zzf+BIFiCm2BFeQMUKsJuoGTBBQv5Jpl4GqTIMl8IyA0GZ313LhZnGLDqBFvyftQ0XBHlJSLa/S
qldODybl7fmZkKSW3IqkXDjXDvWfo/bTBaYsEi0izEB90VU9M+YZ3clcdlDVNT479JOPEcQnrxSH
SJp1bCGXV5+6tkb4N1J8cEKqdmcj+xc6LAfhWfdppmYqiZR9ihZ4tcuMdaBsN6z05dE1ITvXC1KQ
hPklgHJAzbtyjYMKD1qLHlFW2JGqD8FIIh0Fe+XqJSYQQio09Q5GcyPsKAeFZNEjdEQ6vSDP9s90
XSkPyxHQCbhzH0hA03/EAH7OIdpkfU1Pm3IE75c9eYmEtAWRZHp7WO5N4J0sACP6vSc5FsoKmlNd
cEpylyvaWD0pUbQdzxYFPV51kB8SIwj1cuyWxrIpNtjPVia+7de4XrcU2jzwD84MCevq9LcQ9LVO
wmMlf6ZFZpY1viRZIqav+odBczWZWLu5aRixkhpExcmqJT/6CTzgSfVOOwSEfxC81V5f/xPhUmuP
DuiZMx7FgNdkSZd+UIlOxMM6GrCqgEbjYhPCdJEhWYkQv/oe605l7dR2EtzHYtEl8VzpGky6mll0
Xc7oJyYvQ7QeFM0LwdjP/8RwQU3fkhDvX89a9VAr4AtZ8QeWz3ECLSGnBs5XsfSgoFHzCRDy7U7B
h/yPkqWYHS6J5+MjsJlQe87JXxVHaqdyhHw9lrh5PjtWXUV1Z4/EPON7bbFv6CqURgmYQdO2EAnb
BiAdIWeHsW4dkaaF5Q77l8+anEVF6jTnl3ps3GsjyZepxX4n5Qpc6MgQzsINyzXaiNIdoKH4xxgY
TJuy5Icu1ZgcO7uhok9zXCdd3Yd4bSEYzXmXRkzQG0OKsc5JZaC5B5DdViiMfgm1Q57sAFRS1pEC
oljDCQ3ky0UvUSicCPEwspd23KyZGBajDngLPk4jPZsW3HbiREOf5cNfzZqrv/aQv4WyEEvnlDD5
f8YHxyapRfswmYdgdj1dx9i9mKM1+CHT0CXh0r0npXgmfBtKx9RHFO+KelDl+n0fjx9IBpDLp0Ya
fKcydMZ//XmdA1h9xSB6k42fFUkVqFq+AnbBqKm8ntEPbx6gwnNEw1YqDeGsqSDyoJNVDrnZ93Qn
WXQY8/tM9t3CbUgFeCj+Jm1f0yrYfmgdoidgq6QlcEZjpJOuqHpi2zGZXLOQgM7h3FkluvI0ocu9
TnkoLDaL2ebyJGW7oLCdUgw0e67dKo3r/vLa1L2VCHswKuQq+BS5gpaQ2gaAQyIVbw2+KWNBo2VZ
tOJR3pBsV7szaYeqcNhhNXfR4Fek4X/dsJ0PAwfpBTfsf/tk9yDEi9rAUG0h5CV9FV3IpL6HAm5m
2WP0XkEjc6gwRmWqs9XQl4CLm3h3uLWgO4KVNo8zH2DO+o6OtGnpEridRhUXVSzQBcJ5b+A49Sy5
TcDbKBly610Lolusjf9GMvjCgQYfYDK+tAbQEndrrWfFuxK2uaUvvra7VK5WLrsrDYBs+jmuVat4
nQCmy8htxbZgvno4klY4oqGAWy0tnLTazWEd3UW22KFv5p5W0JQ+fFMBtzcVcg87y3uNHwHQ/nPu
xIEBi/ofDPRRgHW7UG9XfzoVfmF0D8xNmCw0Iz3CrX3u6OS95dld1gl8Ag+2h0SHI7CwXTHm5htv
V+p4nxzYru6LlivkajYjX9jNr+1Qm7MGslW9GnSm4D8pWtEZwWB5DqZ8XT8g8EMBRHCqCCcMr5Q5
p48FPeb6w4T2uon/EdoBpCLbDBOTqS5uumg+RJyFQ2jrzHS+WBFeuXQfS9z6txz3M92c8Xp46TZZ
Pr/FBIwm48ZkPSn+vOsE971OWxl/kKAX03ly1cR1Y5rl7iA0W3NMpaFedzvCpV31DgD2+w62VzTt
B4D0WFLkSKOuvSUD70GiorVaBC9TY5yyn0YhasOxv4RDRFmDHL7eINGkonI3WseprnIZuCFx2ZGG
rISB+q5rbrnnk6a8omqo5xTGgfALzNU/M5pYrpoCUhsZp8Zv+/fC2nZNcedEFTo/+QSsiLXm6I/A
qwwdTvBd7Q0Pfn0ZwW63u1VmB55bS2286aQUVzrOb7nWahLSDJFSlPcXNNEOW/DsG3wuMJUJoL78
z+7y22+BhcHCSMbCCzPg7AKRZUTp3zu3VweQYUydUGI9aFKfU/0yxW92YdwdLdT9DA/gjLJCCipC
uC6+30M8yE+pzqMUtp3PbH/7UgrBfM8botn7Q6j9ZsnAYYxszLCqOocvfs1UQ68bJGYZuOuwhV0l
W2sJqjZQyH7tSnUMjNYbLBbrrpmYF0tZZyxZrwnUZfBWttdrBrUvtejOVNj3YjTn1ZooqieBnJ3n
rL/FMqQ3ydx0S6eP73L0aOv1SdIa8h/cifKAncu1sKV/17O77QmIQ/FZs06JJcO65xII0X68/nhI
FRkggGTU1RnFOlI/J7D1kcm9TGuixWz9AdqyYtKJSGbrSmbP1bb40/01Zn6PBZLF6HOLeNK4Z5kx
zYO6UYpJEbUprLcuP9av//scvgqD29dwavTaIxKW4Pb3hH5bfTnZkxwN5phbqS0qGAd+peXsZCgq
i9JSgIuIrL+11YiPC/wzBv8V+9raVM3cXpQkO9aAmfy76HBj+X/66QtTViTuB3QZvOGu1cukBMXi
qd/o1LGaH5v6z+Bbb8MwKhsvzhrNRESUR7JvXAsWfL6zcxxgq+mKxvKMko3UZee3K8QiQ74IGQrh
PEwBnfr1FJl9Y3/fFWQR+t/lIpYnt+qGX1N+Ct6Np9Qhw7DF1mlbEncsLcSRDqON2fmx8N3MN4uZ
6E5vqE+aLsd38EYt6RfULzG5vzM8qudndsd5iZO6nrnH+d1Ec263SJcCYwwcjw7dDtAVSSH3gxst
M401DG8usGUOm2vzQKlvwL8krMNeRhTo7DUMOpv6R7r2iT44xNT0UeWulwabhgfURsEcbg7G//Cl
7vvVOs0iY1ZIJEVDaE7ZVCxJS5SkhwqX+TLTZl72FFOxxgKSKRHMopTAbxVWG1xntIhje941/uu5
RKYcQEtrBi1+Dr2gP4h51NFyfnKYdiVoXI3UhnKmP9EO7P/uqpUrB8EvL1Rd+tY/q/2L40WYMf80
eHJJcmNl9RcWAtozy3u3EhwxqkO/36VkCya1LtuhYMf5tgHvWvdwMJLbZ+FUUrFXS9AU8dB6ddwh
ldzOn1BKBaf0BYjuKlRHh1lj37qUpnOLm43hNnhwthgSpa220uerZz800UvDiKgebfhkArXQ7FAV
zHkgmiD8SaWCa9anEWMS0/woZlIzxp3SR0nL9n4ymOhptka37WC6m87E2K3o6fevBFzUDMiHv1iK
dAUbWJ/CkxHnLjo+gjVdAl+1Qmtshqt/6LbUEXhIa+WNO3yGo4gdR/BxmR/N1ZOyvSGDtUPrJcWG
hqmsahg6L03mWNA/uQ3BVeVpK2KyTxXZURlHFxiy1kbOB4hjJpqYXblEN3BsRzU/BO07t1zGwO4+
xdBGR/iVBLglc374q1AaOMTqzhaZ5p8XjC1oTm2gxkGrHd7yB24uLD24HdQv9EucsLJP38obsJUk
tngWdDdNvo3rdB9hH6hge/ObDOTIK2zfxMBSU2tGCCxVEy0TuowNwF9GbG3GH6Hum45zrCGRCoSI
Jsfl04EUE9g0u/nuUfVqFzcQMwhKttkPT72cHj7+DqIj9rtocopCDpaidyy9oBBLlqjioqAPGvqm
XvjIzOpKLqrMSe+BEh9R9rMMAxkYFccl0og5aJhwIGnCZ6GPj09A0Gt1E51JV/mQWpUHLAYCkJuX
OZp1ccd4/p9OL4486JIT4ScOWUwL3Do8rqP1Dwix2ZqWAwyNyPY0tf+sJQ+1wWid2xxc3YEeoXLp
M562xSsrUI+B4OkyUqHLZDcqYYNZc8F6R5vaM4TsnurLm9aMn4hPA3gL9Qyl/5UF+4ufKYfjjs5Y
haeJqPEh4L7XOCZv62oVrI4ohZk65jKEFk4JaOEi0g+iDlRxvJz+mdpAHdgplsuVew/iA5Slu7Kg
48cRyke+jF11yC1bSzNZOCvyyqkUMEIO/Uti4MTfRbyjjaqH/v7hFRIy1Ul6Y/pi0BCyQ3G8tpJV
AHXybToyIsRR6wF5WIxovEjPLzHYdXB9aFRgodlTAbWwjowd/3jB9GJrTHRPZldp3pV8qGpmokQ+
z7vHWJx7vY25jjsxFRqNu505DvkPS2LiH/lQaTf1XU3jSJJV8ZrYcrWQfVTnuxxX1kfGNSBZBkUt
Ii85sRwO3Kqv0Zenfqt9E2jQ12NI/QurX/gJPS03MA/kcdr5Du+w5ydw3ua18rrp3MJkWfZKrodm
7nYn4AfazM0QU+WwBNOv9BRDqkdvhOsVut2xRwtrJxM+owsk80tLnAg7I8Qx0h/m2Jm6+/fweFpJ
M9Ziohcr8+0yC57xS6oDK1kg8wsBl+pMn7CoUHQAV+SAg2t+gbiRVN1z28/idR1GkEOtSGf2zIeS
8yr87NxOaxjMMZ5DC6o1s3W0I6WhTtrUrjuqZ3wfHWOaTAavSbhm/u0m/6oX6YZ9hXBjcPkFVmpT
Pm3OgfP5B42aPcCG6mmkTcEbXT5jJhAjH67+7JyZ4n2YSbkofNxatJSIrG4jK4wP6k4tDUtZckWX
sbC2AjNw7UBP2ext0v9Fnd2PvvwLjX1hbUSwNNcQyMa1/TDAdFnVvMsbiGSLnJYuUw4MTl+dMvG0
DqgewvVYvDb7B5xdrRA2YEc0uFrQOeR/ctMsGT9QDrljguNbHyRE3YOTwQpt837XmlCTz4FiJbRh
7EL+DTlbOIrByDHCZ1pqTQP/UX5nfjgJsPiPZzk0QXWqwRaiTenRRDvqNkaU4Qrpw5xjd3aqz4UK
NCLbUge0c89Bwzx92RuRF8d2taA30x5S8m4860VKXUxySHdq4eThc+qtJmjiWWiqO9rxU7xul5sn
ihLjmBjuaIT/yRic5SZGc4JlikbnGoCs/wCmP/adRFf0RfRF5ieExFhJ8/oN2riH5a3Z4TUsGdGT
YbZ/REAuX97tXRQK0Nu7e7dHiuDWNo0pVM/LjsHtpV6HwF/igrBb2leO8S2hOgu7CNK6ERSNIYYb
+itkQXFIucZjm3ox6Se4Uw4fZk67VdYt+/Fvo5KVIzPQxGvyjJcHqCrvVjWmFFagTl0Ape5e0QBb
YUU5FlS0ItX6IsPZFV0HVWI+jbo6+UtTfTx72iBaAPnXiUS6lW5PyHMbdrCiNzlq6WBRqkdPnzQ0
/PAtpGBhbP2KSRK+f733Lc6WSTSfJebAcrXOGulUymi0liWFWDy/X47gNWCKVA6nm2JYpiUaL/B3
o0Tk6NQtam5F1wMMX4jVUQtbf5Dyaa/KfJhMDwXTrFPPDq6BT6Dxtnc26+D5m17vCm03plgOie84
2cNFdAVYMykJ81RwuzNlSN7FBTMeqEMROsF8xY/XkAAQp+L1O6MRF0kNbeK/1kFFjeQ3uE7cNDtd
/oN4SYceya550c8donL37BklpIIQTwEwNXtcoNYI1xkzHW9RO2SaEmuu3QhGhmJgOQKtD0nwxBdm
aJxkMGjn63k6S3voicIE4dohJb87YeknfHexRpHh9I5r1pzzjiar0KrfsapTqq7tgn6vgVZqMLyO
VhR7tE2KoEdlfQ2IELG5bIA1eCDQEwkrqsjgpdl20YpiGYnJy1GSjXSCqeh3aiBtxm8TvYeI/Sit
H5E980MuXJ1/sLP5d/ZAvPUlJZJrxGqDU3WbvR+CjuRVrRjyGD9feM9xYbsQ310Ejkt+UrJvlJHo
MUV/vjJFhpWphbov3/SR5QAuiZ+Yc8DQFdM5KKOWXbozHc+AGr/F5nCwnINRTA78P84wPwLMAac1
5AEq5yqf2l+xipC3EYrXjpFfywnlCBHFctNl9jreYa1lbPDNtUOy4KugD/OyvXSX8dap36PW/Pyr
L6l3rwHk3g2SebZ0my3lA7Cq1lGrsWsSXkBc9TvGHXO5bc66Zbp27U3Zrcebsmy7DV1+Z2YCP7kY
sm/UyNtVBBiGP8DTF259FEl3WdB/h9fKqjvNG1pJ8/wnG5epWAKBhusX8FBpSsQmXwthhF3vQe9n
z7fqCOr9FgXjb4YR1eeEdFDLVcECR+SJBQtNrEM5+wlTJLUljSVBVWlunY7jJESYY7AFaXAsxP8H
M9ChfbHwWXFEPJwYr2qbLrSNYmY1QEMvjyw9Sl7JjOnoj0/AWhqluvtbAlgUF5m3M9AkiRId3U7Y
c9AIvDO1BSrARAdoL8D/Iw5Ddofk89djwu7GqiZHfiOrLLpznmnyeUihwAZcijoq/ZrXU9ctH6C9
saZGKW+YkS1rTWlF1+V3rjdLxlutqZK0Om/E7P0THZGrpGuvQpUeTATz8pnWcGlsV5m9HimTv3Bh
E3aJUtovpqAzVoPFuYY6seCbr0+EXPO+V3fvhQXJdct4HxkWiR0fC89yhyPk1F0UMGkxJZk7ujjT
W951fjkUSHz39vL/hKb3l47UE+B9Ia1yN2pRlsU0pq0T07l8E5dVr6zSV6QQTFSieh2QOL7pHO8m
kqFiSTMkcmIlj/2Rl7hYw4iAh4Ukt8Gsq0k0QYyuEvmPfRq9jpIOf/gpGvZ5LcJ/QL6/A2w/QrwL
LF3ZiDhcX+5F8EtfGJ4ONe02FnVe9pebfPMKkZeJwOXQq9DpyzW1PKeNOYeb+XIiFIq9bvUPACi4
CjhTudlGzC8SHh9HKl8iItOYO1y1X4LswyxKpYmNU1XS28dhHq0/w5eoxqW2vE/FxMbSh9WaMvZx
R3elSCzzAudxnCdZ7ZnqXJiDI/uNX4vthThyWHnvUCkFkGPTfIT7sIC0cIDkMPgss7wHkVx3uOxj
aOO5FrOD4EevNX82Rz1JI2MkxKfdQfn0RMwOunuX8Ni9YWWE88CgAvi9OPmjMNuETwQNWOp5AIfQ
ojlufnYwPTtcNuPJgcNwipERgqVisIwSo+5e93asv8nqhAGQmeHHUZElRGL1nFKWY8VZBEEzGA7h
k+15X1aFtR1sS1XymGIR66bat54MwBB5mgmFqLQJhivbOewOVi/jBvtgr66r0pDlPaYjKhQkHsD8
pl7r7PCyuC8vL04GK3vaU0eg+YLDHMxTbMYFjqquJTArvK+6qTnrDosHcfhD3CBiQC9PcNpqE2fh
aKWo8bEprtDMqJI/+B2qkg1WO1jQjLDaMJMkOKDjgKdAV8HKqZ8m8DovmRbERCXmArRJRHGcnB8f
Byl+TmSyWLQtLXawgwwS2xvFK/t6f2+BuWJnz9xTOlu2+7YdDI/1nyAQ3Rw9uNLqabA4L4CKZWwR
C4c8wE3uwgIp7K5N9b01t8sNYi1FBP3cQUMMSHORMiIUvWZe18SU4UOp4srbQ1dV9WJoC7JWUZXR
zq2fjNTgUbM52kA2fzk56gFgeeygxLC+YthHNyZdbslmkXpnvwc8caudBFs6BqK9OBfoYTogyNv0
3rxkOuD1m+f3BB6LqGmSGMMCdPP9mmgtXsSV/xoLrkRzFqsqsbA2/MvO+VM0ygEUeeSykTGJtVui
VVRy1mGEXUBDpDIDbyDm5cw8X0cg68YwWJbGnuJyaraU8gXT2IdAU0BuaAhqkii2IlwqUKt13TAv
lim/qdnj1a1H9pb6ynF54WJUJ3AY2TgDIIriP3b9Fx6wapEvoSTfTq8iQzUB2f7ACziF88IUAQVp
kuRefg5U5/eKZyMoVHg5UGTpb7sz+o6IH9ZCo511xMtx26KbByoxzUbQeWuVv47cRByZiJOGYUKI
qj9k1HRKMvUIi7T4jewqO4REAjWsvw8l92Nspx3wkx5aRj41U1j1hp+C3iMvDbnGUu6rvHlLNRHX
JcP71GzcYQvricAfZAGsf8LaC3BnEdCTEzSUOjXBbT+7CeQcwjptE+qzCFRL8HWekOeNvCgyNa88
jb8/QFPc4mo0MyTJQbMw/+/tLRVkfNT6YfxrfUr1b1qFkSB7Y3o9x68+tI1wHYlQgyyE0rBeOLum
LKUwmMRoUw7OD0/OU9VHVJUpwX6rrtLqavcQ3LThje4zmC2gfygXtwULHI2LrMO+pytmClTxZK11
seVpCN4JUwHQZTdp4cC5athPwc1k9SwnWyEIFsFr01QeCj/H+jUYosf3LlhaBWQe2VSiqwnj2oUn
fix4gyENU11FRZ1rId8n1pIhhe6aeI74MqcZfNvf+MFExrS3V91+oT8Kh5Aqx7EnP711Z08Xdn9p
+w786shzgvrJE0EXHraqSxxZuwJzeSbpWd0aRUEjJzHs79k2QsGQtfjr/CxmK/Jr54rfpGjfS6AD
KFoJrl1zZ/4/Jsaytiro0SOHyWidR4ETPTfOjHBDoEdI2an2yWsB3LiPMU6csPBtGbCS+JqKDy9X
zii+XoeYo/q2wEqbwdX450qtYjXVfeAv6SlUSi2LWEphCoZf4eFB2hYRoJNREWMb8QCU2JqmMalJ
6sWrL7xErxQ2XfPKl3ACebj390yB6IbCtbBqqnBo79JPr/5FNN0NGzNT0DWBRsa+gnp06yz8ppMS
xE5QuNHvzQXIbbbLYtrSKHkuC8O4g3HMMDGEjjtTzThn2VvErR/Nl3Xjwwqlqptfbq4AlY+Kvy5Y
UL1/VYF66QNHr5mkbTdZT0DbTUC35NY3sm8mWvOQb+iY3g8Ml4PENGoGJRLtiBFJBHYedUsA06eU
BW8B0HpzYxo2VFTe3kAt/earALKelPkX0Y8PIHaAV2h5da5tXiwHtRlwCBBpI/i8nxkCRpPARNJP
1U0tz/rVvKs9iAY/AluiBghT+pVd9xFFMv9SYU90dUGWhu8nQ9xj3xIKWVshKbdq41I2jySxOHLD
3fTr31QnhJs5Pl7FrtjRuR0lxvpaJFginIoct2gVXnAjVaE2484EYx37csDXMIE3sc5oBE1mL2tL
kUV19kpUKrratpn/Asy1411TXLh8B15TraJfZnLvCeYOHabEgKvG7P9WLYIGFePFjBYgMHVWkWry
YNdWUv5Fe688QzOAAQXrtHP0PfWq3m6KzCUEfzNnEfppSFH2vXFe1QNBI1ytbK0CwBGneQBviDfq
WG4hE2bI5YrgCZmZGr2BEPdLm7GevZTXBDn5A8ReJOXt8G3dY8En9663BT1WUumPU8k7fGEk8+PM
VEZRxQgqOk+UEnLCSVpF6P3OO+55luzWtnL+kf7J6XfocKOVuiEHJ+S7qCN9eewWTQ2thMBavb9j
XgzGSIYsN26/QKSLqTxfw0/wKcDcH9YQThIwmwDGSAfe05RU+zEvnmjm/Yt+k5rLHrQnkTZSDQBs
SpooVWlblPdZVpoYo21DMsIpfvXm7OVEaBVStuKPd/Jjnsev/3x2z6wKMQAN7RYnwQ5F9ZA1MsXX
JKwMzhLDu+meP7Qtqr25+SyV9hGGmWvBSZugm90QZSROlhpMB29/PahVSWOJ9STbgf5gMFybIGSn
YJbafUMc2mYt09zkRFLp4W70y41LUJ2MwCH0fPkHYAjr/6mkufx9+fHBaAYTka1SKwjLpGARY2Eo
Q+YOM5H0GjIoR7TvGXcerqOulEojalnEd4TEjXSjalmxtnTnZUT8Rr4sh9+76ztm1RyQMgfT5UzD
+0Jm3K61dwFfnG9q61NbbirouC3NU20LbEHNGLcp1eOmPRzVew/0l9b2Mobi1OYQ+e4cytPp0pBN
eR183drF6PPFcj8qo3qtbFck7a602BVZv/+NnGyjm02ZP3nmd8liblBmo+a7MVb4jIwW+e83BpSy
md1ZzfazgVmHSvtWxSR5SOa2C8pSbRk3UkeQ5oacpOwbKyrTXJijBULyjp8/zP5inkhp6gSatb63
O3FxB1Op3FMG0VhvEYb+7ytlUHu7EbtmQ6ZyJHPeeKg8zacypQDBFYCpBtvhXhJ1dO5rP9AczOod
w9ZCzmrsPLGOmSMdUXdUr7kTkkrgMxPACjj5msNwGdXm6n18ps4nxcFNxCKV8kbma6RJ/fOzp+x/
HamZKXwKJtVMkPffprrps4o+OVnRrn9NtSH1oIBihUS51Gx2cS4xNXoxZWmP4MvtOm1403tLTIgW
TcNUFMX6kClRQ3OLrBu6a3IsBdkC8hHilyxI+iC3HsNjMBO0sFZJD1fTLZCWfVJZraNIswxZ45qy
LZ+/BM8O1s3vFM4J9x8xaTmPIlnvTpKi7vLs9AruV3Ay57jpeyrbE7XD6U5JsGMhTxQVuGrKpFwm
McWNfWITrAg6RYe4T7UCCj/Wg3jf+lAqgH9lzDLPTbh/rTidbhdUitsH+hotngifZ9gfpfV+1MHi
y1y6nd0ujYDgdiha4+iR1E1R+7qEUo7A7vRbONRYmI4C/2gSS7N6vPJhHLw5F8OW4Do8gCTNuBb8
DwN58ld/CmKTiVRvCsJdJfXnF62gl536wW4F08pNkOuUvt3uFzpLl1GD+uTT+IPXqWiji1FuK9Wn
bfFX8B7jQ8zYeyCEovTov+wOAB9XY+8upTqF/3j1RLeTIpT+q5nfzfc5YvwkDDMbAL3mH9wY77yM
I6UaWSOVLvgpHwD7zaQAkoQhLREHUmC44w/QWH97+Z8ZvrQmVfLx7rA3jHOSal5unrjTgfN9tAxR
DNjS2rxqucTAJWKcrFzFIXjs6+ItOCAzkZNZT8HQjLvOFBUQ/oY9jlr5HcIdcHZc05MF0bz4lwC6
iSrq1N2WKGUUFPRtRaWHo7cUEin9laBs6mZP6l4Axvoz1czPTctEavdfxrDipJ3oLYdo8OxI17Kw
8INoUJSF0gDBx6GQ71sniW21i5SfENJ4dQZoBN62J6yx1wTzKeO8mnA61VPLQny4j8O2Xp2yFd3V
fcOyxrwxxs/hJHRwWuKR4VYe5Znc44SY7YAVYbHcC4dbMILAG+9FMHPJsOhMfRhMWb8G+jUCuKrn
qH0W/DLbzW7p7lwHOWbgoR0+bcEx6Q98YNh+xVJ0xJdH5dIlqN6sMY+qWHOkXJ3Q99XGfe4HGPnA
/L65SiLaKHFTF7hLePp14SyuwIW8ugm/UTmXdZtw7uuMRQqtU/s8YyUwqLt35AOrrVw2Tr5lgYxL
tFlwfMkUOq7MgmcdVKJxs/K1zCo5Mz9i3YjRI+sqjH2VR40xhUwa35U7ZyQXIKXB94bB/KHb5TeA
+E0YmCkNh+vUhgSBmgdXVk4KdXMJfLZXJA72H/yUNOD4TG1yiAdTqJRqMbzD5aWBt63GCxfPtUEp
Cf2tUD9Yu+Ar8M/0uce/2M+x6GiUjUkQAgEyhllrEc66gsZ0G83F1i+dC3z/e36iqpCUsC6n9alV
MdtthVlNXyzknacYJUHVbFy2L4cR6p/I2m31XysAVYbCiw1QJfkER3vyVwPCWvIWrjO6z45DeC7P
GSjYep5cRR34bjFh+UDtEyJ/rprsMzdomJL8ftV4xPAMeSEojlyuJYIGfF0BT4IU9rRaJQZpVjzh
RbvtypxGRzTg7h/H7Bhn6QyYJfr7GBrHwTV/Pruxl1Mt2sspPxid755FcVCYKdx5JnI8GQkyax7X
8hzhwokkodxX5YeUT5//QEcwOwnvm/40rgI6ngPOTcGZmegPzEgBDsMYkG7pjrO1YWDDXk9XCs7H
T1V46m4DpRf9cHrpFkRw1jf3TC0MdDlOIAJSMY8tWc7Ch/Ha6w1lSZZVigVpn13MQC4DJ33GO0gt
cA2ghLi72g4K3cMZYdFdp5RTIwqVsxJ8Yz8i7k+WGZ3TsW8I+s10sPhnLpRUDEA2ab8FyzRX9UI1
oGhtMjlOQv9/kDYCN8GN9PWQTFJNq1PV6UZquDvT1EpS0WGlqXtLfwZpwQxWoCjSXMenfvbjz6NQ
eMHQTTUy+nxckDPJg33QPVBLBVicCSWUq183C9sURl/O76C8xgZM3zp0hMQBIeVnfTy0J6i+hX25
Jn+D8SAXlaxo4lvJjJVTn5HXfOhZW3HXLtL4a+rOTZ+YLwndf2KvClTqquzv57VpQWTMmlMTMiHt
ufnrwPQorgkG7hn+e/sGpVDM3bHZOznpeImFUoAGYIORy3mEr0noc82aVS+ThFFWttjuDvbfM95V
68kJfq0xGg5aDLoGLdjOlPWcK+QOBL2nu7JZ1ywHqbETDlLrcP2T8FdVQvmbUtIpX6X+MVchwS8U
fhrpYpS3JlyvHfuU/YjBA+7xhCPElTEg9JjQ6wbHPBMUnaiGAb68MAfDIJIW/Ucy1ZOLhOdruRyh
FC9mNlCAIWZlwoZFnEVp2igSj9UW3F5IeTkAanUwpL02m6/UU7lLW3vr7pFcnjsPpOGOxe76Tez8
eKMudr2/HpHjvzXSlLlzs//+h0Ko4FAw7oGw2jZ0YU8JfI5ojzsjKXYOXC1kC47lxblrf1E3QcJX
vkAsAXvEIAq75FgVTkjbn6NPLHv9YxUOvg5imu/1cZXDpWn08tFa5+iwgsPZ18leGxxjxfsHg8/z
qoxeys2mUW9baDz8CDn/VMCq73DKXC9Hjwj+Jf18Aib7sk9EPCDprbpW6iYsnf3sjeyWpwzasP2t
G92ZVxz7GY5jxbFI7weW21LKsfyyqRmmUlIY1NDOLKIxNKl0cIGI+2OjZhRS4Npugxv6FIEYZYcM
hQeKpByVeckacoFJk/5xz+FWmWi043ktjjltohn6CtPlG/R+dJAKafih2SPF3N8dZS3eeq/TmFsa
pP5wRx5F80SboCp1IO1jEjYO1uo00fXSjisS5xQK8kzSbWo+5IJbTWrWlW+i0JtVD4PH4bMj63wc
/uDn6Bv6/bXpih1L5ITRYz8etTyjjtM2CZy3aVOjyLF3d7Vb+wtEr3J0TZHm1DJfwz34m7fwWjKn
44O3fHXF3axzwOGF2+BCXZtxhleDNEYdm55B27nono501X0qzXHt0PK5xSc7RU49e6vcEZwWqsda
TitraNcupGTioH6ZxVRFldGNNuC2OIeDx5ETNNv9TBwwrTdkiCIzfeqecGRxgWmwjEgOzIT1y7CV
N5WJncW3JgcDyKM4DsgTr9FYXCs5fbwSQRIzzX7WT7x3XTAuf9HPPzeZ3AJEOF7K9vREAMZXRYFq
dZhVqUTHNDNmpwjQ0nmQ7fo8D3EYcAosX26RGLnc0+8xfmdnRipLHqxKaX0hWm+7K/kOkufrQsoi
pJQtkB45WfB19wjwQN4w25lMu5XGWcJBqRtD/WFisqeBCKftZTSGCT/swcFxMb00gNUTUhaRgLtZ
vjLvlWGzyw8iqGwKJf8U2bi1viIzChxXxiYy3uzdccS1JxDbMwJUq5SGjbg4i3+ieUfs6MO7fZ44
4Gkk+clgQeF7e9oqQQ1J6iFTY6LAulldidRONsBHe6gsoQX+JUtn3imRm6nelYCYVHP0m/Gan5fa
g+pKjrPhKfywj8h9jNo9OKHtyONngKsAVp7umOQBNTwAvwgjnWpnaoJTqERXHLwSniNOemnuv2tO
ASAO07XDGOM2gbuGOPbkgyMnUBk8oG77Eny/ZFrM+cN97PhhvTBa57vE1Yze7eqa0fedjoDgLn1i
qDHq82U+EInYLq5+3pdhGC5AogbY0jc+w4yRx6JTkHdo9a2uQUBQ9D/LFkxJWrlvASyi+TzNeygd
g71yV5IObipPiCG4o6MCfWBGZKHex0R+l5LSy4AzzkmJ57+w6D2TPJrDnK1QYmh9zBoo3gMxp/qr
SH6+CXGF0U1VHWI5T2OehQzgevy1Lxi4xPQu40lsiwanGHoMSPpbubNeYBSY478ezPcWxYUOcXZm
8wuXbSzz5JfNyhAkoVZ39re18tGfmAawTLuuItimpN1/vEagAJRrzbpll30092Evj6mKAx18oVBP
k+AbCUs0zjFAcjI8eTLyuGvESM2BxS4Y1VYaYZZNEVaAhm92vZv7Npbmv8hTzPQT9f7youBZ9zWC
nLNUIy5sLVBh+JS7fjQ84hLCFlo0xTaagE/2uQsCxFmBbik0RrgoK8xC24pc5Mbo6zipMmFd0VL2
r1C25D/NbflsHNK9ybmDmKjkpQWxES1pW+yWjab1Od8b+FV+NwO5lYiRMFv173sIxtAAg1aw4vGI
ZTDPTf1rP9E3d9fhL0fjwVO3BanpbL+sCQ9IEGKxj+VlDV7aZ1z4YfkULoqsR2mAACWdYD5s0E+V
vQbQg+Pkfgx3G1+PrN10VPrO5009K3wyEPs4/mWpPUSdUvnIJ0DiEd+0tf6FjVdFUwvFjQFYl5YC
Mn2HqHGZRzKemwFdzD0xCzPIMHTW7mVD0+YhBVTj7Od4yE6vb+xilUACIi99HWd559pVTsAMmHro
/xFzpbc+0reO62YY4OuX9MKPPlM0uFseoSOxHiJ6pIncgf8S9ZSvhanIgFmJUk9t3DxUV+2uyuhe
XBeI5mJwNSPDa8ZOtid2xYP6qdPlek110jZcyc994ZT78lAFW2ccNcVRbIXjuFz7uS9RsuAiEphP
zfGnisGCxAY90qIp51Ng8bjazJpGTuDu1KPxzAoUtsQNIRood7rGrQonnVrBBuh3JtdDc/StPE6z
kACfzlBYQg+DDqBLL/99a1zBhSLR0MxNSic49H2Jckmjqp8rkSqE7oodd4H/6dsNtl74nTzwKVBL
9SFxhaKjJTUqEThfaMwN9yW67e31lhbWjYA5ASCK2XyqO8aaBdF8ZQYqsEYQhrJqH2+vr95VOhnS
8m92YtBfwt3QayIaBAEMpK4ziEwEpl7Ki61uGJmbDeUtNqjyNlo5Zde4eQhZBvdIEsgKfuqSQf0V
U0jz3ZpKOC4Vk7Gd+jCr8PrsOH3dnZ0ao53EUoCk8CiajOCpP39p6s5z/tGux0VdYuGt5Swn8XqF
x3JYofTH+caSKKkW374o77kHHVx2cIAdqOtdBKxv0erw5kO61mXyBPJStBva/dzJhNifmbt+KBTL
ETugbs9muEEGN3ECwr1UMz2KW4c8Lb6WIOHidp0EEXUKF5Fm/P51smCT3CmZX0x2J+wTfyNzqa1I
RKlvE1V0bymDJF1qvbEISzlSLluxkC9u8vFRdrvxmglOMK+quYnacgVF/Ks2kI9IZTYLtu8oNu3W
XjsnPc2tyhJr7N9kpzcHdew/Bkkj78TN71kIvAHSsLvq4XVZYcel/utots4Zv2bVxmU8CnWEEs3T
ZbCDKtihKYBfILTrZ7TvrPBLmjKZTSrXf6CZhk6VVsw2myE0JN+gLZHGyCOHSklSFsqOtorBwcny
3N3e23MRI+JrSHw1MjUOQiTw3IgL+Z7gOCL1LkIYvGlW2++g9y7Kiml6QIWQfX0j8zXwScvBioOL
K4iAMkYxZ2DDJkPFUsrw8nm60xTALwpSd3Eqgqe4Aq3+0zBhEx8AJGb7Z50pUZO/5utaYU6JR1iL
f36SIqj+yANWzYCIzSsvuQNHqyJzXLAJkIrvlQCi0GiT4R1Gw3LUCvJdFCMXDWLRJFntSWuYMBWp
dXDeFTuWPdyJ9vJHbX06UshpekxlIA/JqWG12nRhpoScxHT7OEnEdeZqNCJBjdZ0kD7mmhxiVJtl
XwVNF0Ks8A6mII6LIfJ2K5sji+0va3vghFSa+W55/+WYoUg2WaV/oXWUkK5uFxgWXn9vyELzGIns
/TyLgDUu78erssawr+1TTxvWFRK605/Cw4jeywcU3ido/J90M45KucJQXXYCrk7JvNNtdBqSSGg2
H9cpesU04D5NZmtdGKf83ovgge9G9L1nLF6yNx4HdrPdeoOnICgITwzalJTcBc0Dm2hD/3K5TX4O
JYZlW9eVx7YDhzKfwFBrmPL6PV3tWm2SmPhzQ7DiZbtAk93zC4Vszi8m4SZwGQlBRqe1QjK0dQhL
Fbp6DOuCoRrjJxlwwEz/Pl++dAt6wXCdE04JmHkXhu5zsSFC1qVATJANi90D2b8kbwey7bhRLvN1
ETdPG/O01M76gsToNsScIlrENLcbXq9U7ek1CjUveUShcwaH3m+5RPbi6zoPOmhT8kHePGmD1kY0
TplzHFpJopsSVy/Sai7PoifXN+EGPH+sd9vg0EQtu8C2oXS5jrwU8JEmQ1IWsQl6e6FF+HiQZEbh
fDabmTkM1IQaKll8zzawyCysOjNOQGfmIw1KrMLQxFhs1X4TQq1VpY8rp6DMIcjqiQ1uiVq5Gi/d
6Tl0JxPIcKChBvnH452OA8WTKC7A56siQM3CokGcIJ3HXG8ViLZBEBuDhIV3oeM5+iDB/9P0714I
SMwGpkHSdq8UoPfOKEc5rynnROOmQgRLU0Nx5t+lqDbQi4yjqMvVR8fsVHBinvk7QMyNh8jPEsp8
flttZFNq3Z3DOQQ6cpZhHKg5mfohnkgwzhfezS8Uu58RrCbVScDU0L0AI03wKfjLoc/AC0LCqv69
hp8Ogjgtv2elvecYbe/c2rQy6b/NxwnEVgTgFQKWV3rO5PR7wRlpR5TqQvknSjER6GBRVV174bd3
4of/akPM6ZKDemwSgxcjYPlAPDkwqFXzQTyQhIcO+O7rMQPD2dPHbOPQpfPJZUe7hm7edNtbY+If
O1p9pKI1kklNKovQjrhDZx6X71MtyrcvX92Q4u7YMYHrE9UFvrzoyFwBGcNocuK3vfKmtVBjOkCA
jisaMbJfG3tnF76suUsj0HpihE2qLZnZOjW1RDNwNc41F/bsVzVm+eXVlpoLaAaHr0Hhw9qg36wg
xx9lGP6MLNpmeaWDWRhx3HR66bKVeigYDLlo2t5qngE3/GNQwNpts+gv0082+FidscC5RIe1T1wd
24EdWaOUMukH/cqJO0qt89yFTe4E5dqb0OSOH1UO8xAO02FSNeCCy/1lUXy+PG65yDvX/KMnG6E4
QI5RFneqp/zSVL6gvl1y71xLTAjWI6HR1QElUKrf9vWLzsQTZSq/ejgpx/TWeM46jsK0xIWnELVp
HWeYrhRxkuK+Wxr0xoEF2OjOSDJzg/k0AvWkpPQRo3wqLFSb0ZisAY5MU17YgfnpRGyl7JrAEYYw
xQQ7V1+5wLDVO3HFMVIwqf330+byBEex5ZgHkY3mhfOxriGStcFFYK7CkVS+8xd5EGbY/7KHWMdz
56MFCQ0syVqbj241h7GjR196uJEG2mDFrtTDpapZmaROoS5lamPH4mkvjaj/ogDbpH/oR9D4V/mm
ZVfhIcBZIutrFiPnX6oas5hWeTmOv/8IqDdEtA2qEehRN3nNaja0XDkyiVbNx7zJazlaMgixrRrn
oQ4qCJ0rZejXkOqm+tQA+WudBWkQM4ofCZJg+g519rItju0EmlAlTS4IiDUSV2gIZglwpPmFx8j4
DGv0Eq+njumuZ1iTcv7OinqLU8OPDM004n2BzAKf/Ccp1zOZLD4CVcyVlyJIkVlXS1H+yl04rE7x
yy6zzs+c5ppcscE+RId/CDzTIa/+EcKYZWn/mQAlQLmSfL1yLqZmp8GZ9MosEXVn3LoNkifAP+Da
K4yfXV0RoxFtBkpXP+GWowWcxzi2QVgptXIGKyAyjmCuD7Fd6vFaqdpc6Mjshrgf1/QiYmDkKM8i
239z4ge2YD18I66LIl4v/Jt3+P8ob/VAZgrF41it7DnS8u2c44hGbEawcFRBX+npsZf0FObf/3p9
9+m23HCcS4ZPVdhNLe3puHSRtaaqu8A251TjE2KwPf/1gDFNoTn6x2KXzz/aY3x+RjRBfOpiBIiH
IAFUgUXH1vlp0OI0kk4siUF6xj3wFcp0dzTUekLkmDPsXBoLZStsGk8vrlpk5GhB7Fs60ihz+VA4
FeocwfvNEjx8Mxf6GAfo4jmx0G8Hsf9UCtUKNQW1dmAXtfDZD3REaEJbKXTVs0hEEy69z7UEO5oe
DTJKICf5uWvOdzHO0cH6AWNvmAvGAREX7Ej4hIKL0evhZ2ROsez2d7jJ7pNBESTWO5wwqQcqoKl4
MghcMdCupMA0lWSrVfAo81kq3oplcL0byEknRGGXn/KAjtgdHJAxmL8aqhR1eDalCdy3IU5tuoQw
oWxTjc3yyYERMp4HaZVnUiWISQ+7P2w10zP4ToTJhfkgW6wVjZz+N448TXynAUPF+ka7GuCzxTjD
+e0BPvp13qsUxIrvGY42JsdznU+E0eR64Go2dZUxQ2+x8kBguq1j0AAByMUzQfbdukWQUz9mZtMo
HxXqpd3eV9/5mrcK148eSWZA+43zAp9g7jIEqGCL4gRxAIJrhbdwxjywP8S8ENLEx72KX0BAEId2
xd0J3DPZ+zmbs2wjfCFmqHHg90LhuF9TgM8XeSo8gy5s0MpLwPHL+8gWWgRiWfn7XBj2ymyENkID
tZ1pJzS01gVrR0Jiw47oCmrVjTpbRkRz6AWuUEADGIrtbIpXVKBg+gYqRU1N3+MBOS1D/b1z/yB3
LDnTYRu0YI31CD29Hi+4AC2tMP+JedeeoPXxPjNRupafTKqYoCIYUqM09+Gk2JOxhq4ujthSHJ/4
NsrdDGirET0/lGMzWOXv1To20TZGXy14lSI4ob+sUNDxj3FOuOrMqS7r+kfYCtL4Hrewh687SDZn
Py+AKodComu1Vkt+ByONY+CgTCt8DXqUqaFUanF/QKJF3rQhkGVyhM0l+3s1ffiYSOMyaJNr8N9j
DWA6KYc1Oob06Aa6lAc1INPU4wVpopE43BY/8eOUqszN95TMhjW8tnhHIqLNM+FQxyW72TuexGjx
oqQGiVoDMUNzQrwm+oV83Pp3y3xstzaKRnVx2wVHf/ccPV+WtgnDzVTOJ19BSWC2s8ADpuk7VbkV
CmHe7euzQcRb3AnIhQZtSkcuT/Ixej2U155llX2lZYxxmNwLu9BYeTvpJJQMGIyk5U342sFmpyim
x6FIqPjKK0DqshJiU/1EWKk2ixgFb9nncJr+Aure6MQIjN7np8UzmG0ooJS/B75HHJFtOohHtcdX
E2p9yPQacuTQTe8R+TI/K8rf3+1rgim/cDXyoxsmeDNhveEIn6LXdtsGvGt+NVxMcrWp3jzIfPL4
jdcp/fEnoV9jBGRNbQO+qL9aSEuWPM6JTykQon0Omq5u1lfbhuLxt8R8X+c/otXVUWHrQg/cqtld
gOlqcUT7k/6KyrnSGSE3Ip6ZQtmtQL2jLrNsdbvjnjq4l2XWL6h9b/yjRcmLSopWYZ1Jz358Is8Z
1ncNt16qsCo4IfNgs/eSL2iOvSi+GLl34Rup9ew7nF625PtGrbbMi6Bc2jZRwF4V85RZBLe+I3N1
hpqtXKykyBpOwfk2rP6wI06SpVXRuaKuGhQ9nJI9onR1p6rThqgCJH+KxRDk5IFKZJzPKn0c58H8
8T/dlJBbaifrEhc6NUjJFLJonE6dCNutlC65ZGxRvq4BUZ1bYIobaJr9iEyWM9raufZnDTePuB6a
X5GFW0bfU12GB8tPEozOj0sGyfEta0AAUWD29fcHKeMXk2c1uR3XuHwqa0LMvYmPzvc3GHElmqyn
MdIpob+P/1LvufiYil0yENMvFt7m6LESgcqVOb74R2PHVJPHt1kt9ovJzWmAEeS6WlxaXIlWNI2j
L7lwCKuGMd8LrR2xogXXxbM2gFkwe5q5fezgy95YtION13P+Wfvj5EH/UA9oJXrhGtBbx/2wzOA+
yBQCDfU5K6AYK/IpzzWovPyDRAq3+wgCqOAOxF8poL60rFO2yzHQhnIvBwLfg2YSdAYhh2Voq4ZM
66jr7Kn167XyZyVv905g9EpHL1nLJ/VnashE4tjzWtxT73WDcv1TWCaTzuqZzXxG+6ovXjP0uUyT
Y63cesYJlTE/HPGi/J7JrX6MeV3TjXQ1xzzB5IHC0eueXrn9yB6ebJ+faveDl4K/b+aSaNiZCElh
yoqPY/Lkzmef0ez7Rc9Gp8+QstXV/xxI79OB0GbwOhLttZYe27/p2cWIQNKkSofiYbES0LX+WaTE
sWnPSRoUzkbA6iL8BItk+wnjmCHCrkkwfwamiaf6ho6CS3gfG6PEmuMDhQ2GgH6zQBbxY89CQsN7
fLX30SZOvNbN5LUOs6SWl/q0ZP8nY8UgmEsv7ebs84b9f1U/sHGaL8Tek6PJ4y/41R+5D6Xeevo2
yGfccejYYf2QsK7j7ojJcoeqd4OFyfqjlmKgc/9h3JmHLg6jJvFXVyUI+nqMSvykraWYeqU/Smlp
NKuNYvCVUwqdUpeKJDKWA8GBDLKTw7WyEHdBpjZT3kK3HOl2VRn6kkmEsU1Vc/so9XLAbLG0aLww
C45Zml9rfFHsodmsfTROVj5q6tDkKRWY/3Nezjxa1fKldgaIECmy5uIjd/M4d1PjgUW/Tq14Ajbj
Xh/imL7oPFUmrytbPHVHjZo14MpxsdT93hRS0EfBDTH4YejbddMdBFY9RIVJ2CNaTQRo83itczKj
zNKn4bXY2bCPItxi7Oc6JhYepTUL4rEk73TOQ1lB/nWazyTjoqI3Rwyxh0KJAJiL8V3yhks4Se03
5uO3jITr+WQV5ZEgToLObPBXCdIAAUk5ISfa0sF29ibsnfdnHAK/mlGuI5OxidtTuNpSNwAUQrub
PJPVOydUwNwcGTwiWaNtpNc7LKnADDEZfxiOyxb6j+A3APP/judo2Part+bH0F3ayjA9UNNgWvx6
Zp77apa/uBhLpZXOEbAMx1CzKEB4F4o+nUjKPxY823bu9dfWop9CzQSi1sxjmhee2npP56axOi5e
MzeKyZMoz+uA0xNMtGN71FAt34zCHIlwpkXuOtP+AxzljKQJmyPblKTdYa+SR9tPOZ3Lb+7XHtqa
2aHbuIWDZwL4RS6SFKbrV5fr37C75xQL1uA5fUdjuK0mPdZefTu5PccBrzSooSl6hbW0bCMwSgZ9
hbF15aJFaQJ1GUeAYhlTmW9Xz76JTKytrQMtls0oEhk5mWXf57Y7TDzWRi7wOqk7ncIeLb5HKu6s
gOlF4FTLDB/+4bgpgjgLXCn8OL+dIHa1/z2guWOKZCJflutyz0wIGNmRwdFGhtj3ZkAwZyA9OcX/
w31pLFIssuTZ3/v2grcve6dt8Mp9+1U2VBCmORF/55/yCHxlS/5whK+m5dBoYmAfSC5u5iX5E3MJ
BDSGllNYWNb3kScYCKfcfqvHfwgydVqhB9poRilMoUBePP6tP2cgpEKkLY/CElzRSj+halPtqJ61
fVyQviIc4wN8GuIn2keepM9wUKuUaS6TA/7ok+uDO51H1HzCRDZGx8tArgyFBXKIBsS3xamAMBHf
TOBZFBVrE6PiRHHskqyfPEASJr1T23FVgFUF/n1DTx6MX8GdgwU6+6RVGB4fASP9Ds14yyY2ci+V
vm95FDl9IXMymFVWNSWtwJURBQ92nQzadAbACyUMph7ty4DuS9gB8Wh7ZM05BPlM47rEQ556QKXl
sobmIWEgKUm9+RDlF66sxRAdkG2b48catnrvtkx5+Pm0OAdZQEiJj1zmdgHu450wOBNT62M2cZve
WjAKxiezw04g7Chmo0PfnMn/lFY/Y6eH16WnDcscOqvNy/p3MkDCUoDq7ZeZ85GZD7wboUa1aNzA
73LEdtDmmfc0dXGrHKJemqQt4vquZzkUp0eg28d2EhWbYKdsBK+uAmYR3S6S9k/zu38O1a7Gpzkt
ANZ731Yw2uDCrclMfDjR8Di7JuL2EXd7CXooontj+5odB1GAzweRla3cI9ledSqqIWBL73CiXSpk
0QEYiqZxl47/WFLAjUa5GUULk5+4TemnCjRRhoGnVQRpvDZyD1sOON8KqSaYYh5JU8GQ3uHy7Azm
R/zQ4zqA/IaytA3C1wOiE8ODGwtg+0a37Phms7sPISBOunMsAYNUs1rd70zxULMipVKkX5/7hZqM
kQC97Kk2E0tiWuqtcBr8XV2vIqaRrP/QQsuZ1Gkt/tqg4yghoAJJ5aNLF59QR36pReRCncCU8Y2t
/5IgDS2ifuqwr9daGOgyjKaZNALSOFEOBYoASBOYGCbmkHSzGXMyjbqXJGrefzKtqsTkYXhbWVQb
lEo1Jz+trDmMh5REm6VzdtsosIYB0Q657EjPOInlod3qqbfKQnifa94TWtEDocipucNnaBXmeiLI
Xm40VjnFChOkGJcNm4jG6XlBRExDUdK7A+NvFbORpDdh6p95QzmA2dBgo4gfpeWZFyckxiUhL8SN
TLekH1jGjXcpWG7gR2Msl+k440/RfYHW0UVKuSWmlLa8XBDOsmjFCFmsobRHgDp6kgeFzHixShJs
Ph2IZIt2kXMaEt8/tGvXO642gpOj8fAvzdb8LRffx6eDwhe6a3kZgCOhsdwD659fXQwp6FoFOFzt
X+ahGwPVSboXW/H/jBoeemKaehTfByuQab2M77h7pFOP+7YzWs4CZXtXkGVj1zcSXCIOS156nIbW
krsRUHf6NGha+OZb8GU/a8sKNnlNYKaOft2AM9z8qm1mppTXl7pbLjfgVji2u1SdG+nCBQ7CAtMa
F5K18/w/pOD1zCsqTGliKn4EzosUT0AUNz4U0einebns/pr7bzKIhc9PUeyqlFEFu5Qv5IhQ7o5i
m570kFbnb7095eVUxReOHXp5i7Ux/JTYLolKeP3B7YpfAzZwKldah0iwWFZQRpXEjdzX3ZKLqe1f
21QID3PyijWzJ7dEGEW3hGU/J0aTYyKLL/KsrlHJ0BPcry0swmKX0baZYRnpMuwEnBymBS9Mah9a
3QFQKIG0QHiXZUsmAi/fFaPN6TcTHJK8RGZd0l+SXTq1VxWkCGdlaNNpV4hOmoUfP0Te6VeFMHS1
Zi/FgHjAXVM/xtFbJi57g8tiZNCYinQIR9Hbs6mY96Td4IH7nZ2wg09QBBkDcADTzGaLxJyj3yLF
0gXUVAiuJWsRxh/YUiOrb3e7kmUKsLE6JMIU5kvWydK8DW7z/jfkLoN9oXonw7yTBthfvwNM0QC0
8q5z9cu4ZKTcc5b2jEz7kYlcJR4sk6IkXb+icdLerr964IFs4a70oYWzeD28y8YMhd7J2r/1ztGx
yxHxHM8o/RmIDWiBaakkQ9VMcmyGdBKjkWnFlxfshHPYdk5SOeQi77597NXyGf9OMBYg3y/RAbja
dCX866PRzStYRKRbkNXESmmU8SftWUQTNzR0dZ+j9tQrRnvefccblk/MdJJHQs28ALE+wy0V1axY
1ev0v65bcIcDC7qA+oNw2u4kogvGsihRKxgRQpP9EbUky97URPsNuzpqYnkUs3YJh3c1K0MIGx6d
yQ9bDgtOplMLd4EkSTdDrcQRofbZ6pLSEO2GWtAcAGZ+8qYiYo6iINzo6wqj6fhHW7K7Fp8W4oi1
hatzVtSVg2vOKUdD0OcVyfyiA5QZcXFGT+zQBfe1acdZPhkCwxwN7gwX197LwdVr3RDUh4HsTG/N
c90W/pb67yESuA5k0SVWymbhXO/OTxE1cz3rmASnMZnOUZsM4vtzVHZxcP7CFVXd9IoamP2vV+MM
mZtIy55tl3DyoWFL0b0Pzr7Jc9sueHPBaK78crmFnYbbR5Htre+LMdQumag3YGk2udaFbxxcIKnP
JBlu1f4b/ML3M3EoOfV3S9oO4YyyDYCjRE6szSCgzjtybNtLFTycn8OdFbakuqFQeITWoC4KP2iD
ODbzldwk/xoM3EV19qqpe/wQoOs9+yjdEoMMyErBkV3INxD97LY6B+3r3vzwhCtfBBRit1byCNPw
yI0JCi2QQvRxjZUmvoP7nONE8Gm/VFyaR3+OVBMKTRrQq3ZHV5X0RvZKqIv0ckStOZnYX4zXnXW7
lmjlrQjhXrFZ74fb28xNniNGMeo+A37IaARxIudFhHSDg3RD1YeJaTbGzKRTKGVTHCIti4lXK0f6
QCpIViXHpoKy3C29x2jXE3HyjXQrcz0ESw/lXpjqfUySfa09w91GPj9L57pluAseITJd1MUA8WsR
jWWoitsVokREkQ+iUjqHJRW1ytti+fw2Yb/utRQV0g1HTt2+uPDfcvvGk3pR7LUNCv5b63Vd6rsh
ghFM3EYsIoPGRp08cEe3WWl6/fnBJkmud6n7a987jNdIXfuNzlmIYTYSwiUruJnNR4IDVfcnY9jj
I2LfIoVFD8T60y8lGeYLJ9rdrDszfZUnMHNPwSRg4x6Cub0Qm+B1nAqmYT31rj7Tb/WMsOr/2N91
jw4+uAGRLHAtVMPj2e9YIP3ztFWxWForZXntVoRiNFsU84tbkhQ3PhjnGKFmiUO3eGe1bbFIneqd
OGP17hp9vK+PSZzgR8KoiwSSBe6Kyr4LNMzbcmpgl4Oh7NY0ZNe2MAih+Ymgez4rjFt5THNhyT9d
2C0Qm/7towH1L45Veej3pVRd4aprJSB8W2ik5F8x9F9UAmgw9MQGD+MHNe5okudqho5InN/Yx409
DjEQxRYsuDoiSsyiG2ZcFPn/RXut/bNRGwygxEAJPr5aj/Sa+3k58wkhPpo0877Y0yajqxlYyKg9
Ac+WrFfaYK9Bur9s02M/QtLopkNF6Z8Mxto9R8yREstaVmUzNTxnmg0KoYE/V7yzZ1rfkxizka3A
7acQciEeU1QJ3sBNPA91OpukruT9Jwdo7HYTa+7QLk0iEEmjp0RkLoX9edKWptPZe78Jckx9M/Lw
LToruEkXwt+c6Ajcaibnwt6AHO4+I6ZWAb09g/VsYUWr1Bw9qzCAc5VsRcn47Un8+sWEOleAiWlS
SDE4p0wdOPK0jdiVsEj4b//0hXcuI0fu7w0X6ZyS59EjcucNQqjOmXy7SuKQNM2D7hRQ2kBh00BM
UIoUC61OKDW599XzNMbnKm8e9cANvv06gGsjtIXsN5qDMaTtyXFCj04XLUWNm1Uk8tu0msCvBPsG
9Q113YHUcs0NzI9KdRdbuXoh9WKjU9L1SIdXkNhjrZe3GLoe35my23eaRTZIHKPTYhqaopaXFbTa
yxI1D4+v/OAZYbB76lfvzgwc9Q985gJU1ABWCkuFjwwik7qmlakGUMnayy5/ueTaJ1BWDeaoIpO1
A/crAF5ZCAvKVM9il9PvxsfJSeaNbwYHYcfTO/idqKgr3YMzlGiGo/qqgojEej9xRhAnwqyEwp7e
oNUKLO5ZVa7a5W8guDuhKCPRFf/fEw1i2F5oEo7T64uV0dkJKvlXoH2a226G5vYuEDp3S3AWXHXu
2SYOWpP2UmDa2FPzhklqtoP8gapyYPsa1eq4hy2seea8JjGxq6h2PBwLmvUfYY4sIR9zTqCEY5LR
lOTajy4YOW6eVvMRb5LAgo7BP5x4pfpyKgBdM1U3W67KcWbuJuK6SztlCMP2PFec8S4J74jm4h3j
hvrjlMgFNuOmMSnRzsfw9WqxgrRp63GtwT5pGORmg9BojCCMM9ChNQqboYAvVEExCGWC4jABWVhn
ureaEtRH7Kx/04zYwxUiz4jhqqkDsWeMSlXbbQG7KjMJSMhQiUr9kQNBZdNFsGgRFWk23vKqLn7Z
B2KMJv9Hvdw9LvQY9zJkk8FfMKlMCpXbH32rQ3lGXNYCuZkwAIW/Sw8UA5UWg1B7crrSj5aIp1wB
+iKQrcQB3uRDxDMmlVZALXXDUh1sKUSQ/uC1CC1OQxDPinCGTUM/ya4U4uoyFFS5/aW2zedhFR2W
yY7Oi1zDaW90W1AYCI2GHSqa5UXtbOLOOwtBlYbwDk/0XnU1fj3o7cQQcW91sgKehOSJG94ZH91r
m1phNyRdDaMndYB8+6Qfs7gLFzG7pF8S24UZ1Gtq0036u0V77hYZZH/tpZTSX5N44kJccQ+y6D8Y
4Gc6hfzqOe+gEyckQg0CA+t19AD410QE+e4DGffQ9DF6KuOPoJetnMGjo011N9vRiNUR7RWyXgaR
IFtOiJP0ODOOnzqN6ik1npxa3FTlpjZxDHXQ8/IHRj5/mbeEuItjyAl0n4MJBTHnOBhg8G19CGfV
a/TFcUxoLbEtyJxKhNVnH9lJjfrTCpA4TMWOi5YCvQdN29G5PYIhIeLhujpemomywzFPz7AyOUDi
Tr0o8pjcQRrTXyeC1QboN6InB/ea49hce8c2yTIprnNxmdnqO+HHQ+DPHyaocj8Pd2h4EAji3qWK
uC902acQxLBGapTsCV/dHPxY3q1vOdj25VHbRRLE2ELA4wKgE63mkzVhe5XP67VEtOwgf8Oe4J0h
2NrAHzf1RexHjF/rFrouiP9M92WbWKnOZGOggHpQEYooJlIwEXQifFdBcrXiF/bDraxUT9PUHnxp
J7JYj7y0JJJNQPpTZd3f975ys93J1OaHM8znEZiIp/WazHjairePbabtkOrim7nD8kU3FXjn4KYq
ZZImnilF2pMnbrY2lOLLZfuBNzTdZlw0QCg3eL5aHQTJbVbNMXeluObd7uqhrKjTrSgtML/NweUG
O7T7v/zMVqDQ7EXsrORtoAo9yr2JuHrVSakwzNCPKg04Ett3azyomTQXEgirQFjZ4G3Fw88KDKO6
IYekcQkYkYMe3KUhdvRskBzcZm95uL/LZKuzlgHMQjRsvxCrigGf5QLZpk9+vmcfUlefAABw5b6f
9RZheCHz3GjWL0Bf0xITjfVdqCWPwRatqJOBOxKsAzob1EwWydy7Atk82gKdrIb5q8kDXWoScadu
EpoCJIwAGk59qMT8rsdQFODX7DjNbvTk8XbicXtA35qn3VZmw8TNW98a0xw7ZjqHUmpLMCn7YxbD
fbfl0CdLVFkoysk4MDxfQAf0TcfpoR9KAH1md++5a2/JR9ILaj4gJGWc9Vlbj8BUPA0oF9htnIPv
1b7xuxK6ffttWrwf0IoVddRbCasAfHf7vXaGL80BF+/lwfFw0EcZ+CLCffMwOknewNtxs3v1r7Av
9nL1uSazFVHcsqaXLGa4EWo7yDPbl+rn9GdsI1eno8os3PI+HkToM/jVnNlIYjZbAVcWdreagAib
lc/dhkcnb7cZkpq+KTKOSN3c9OcEix2wkYNl6yJTl8IQe7JW9s9G7NVoLQC3TmkznQIE5TD+mkVG
XJs61uAZOn+k4JOMPjzGEAo2uhlUd+AP6duEAg5wwW29R25g+j8r/wH4esAtkP4kPX4dJrNVqa5+
KcNJWhJpBal51XZ0BsmL21MXO7w0xY0/CCmUyk/Tfq2H7BAfFWJcP4D6/MdhlxgGN8VmQKSkuPMk
5WJBxxovbLc27edlBhuzV2ytMrXMA6FbtDQpxqh9Ncyp0jLuDFV3DtYFYaUoh+MtsOBGsOwI876I
eXqd1+BARYcOGXALxNmIgv0OIdOTrMv55snR1m3ytCI/wO/O0M9MyfmRAiN7XnUrbPLK7ScR7Rsk
CCTtLTsyz0xrYrB/iAv9wYo4DnxQsrkf5aqGeoyRXf5Dz2+v9Oc/BrEN3eOM2/qsm0Fy5Tmb6emj
/5bmWAELL7l/ytlnWsGBVMqxENeR2kxVnWg6205o1JD/Zr6ecbY+qcSvsA5FSN+OjLfNWChku/UE
Y1f5BYAuW5cgIQ/CYQizSAQuYWb7GCEjBjG1rE9ofTg4jT6UKLMl3Tp7CPzEWk+J5a8sJiAx3Kge
/Fjcu5Sd7MhKeYQV0lgiER4C/WjZTKnpU38t9EOXBV5cZx64bitUuSrr6T2EgDwODVyJYrGgGZIA
ejV6JePBbVB6KBV42RqV+UYpGjjskO+9xjpm5uFhIw5jvrAOpOjndjPUfRCX5ALd6Kq4uLo44bnT
CEtpiSvi5slbSeRlzJYXwa95Ba0DTN2+RDmiWLRf8o3vfBuLDUWrXvUl2uPlILoSTEe96Q1kEClj
eAWfF7LWNVGfSZ02pO2MHlpAqwIHpT+/y3invOgkUyweAEW1xAPC3iOiIggdU27bRdxIQU+/3tdw
OnqN7GoK6TTdk2mwYIc/5ZQ4czq7n3nQfdwbasmwcJfd42TD27Csg/6XXtTjRaydgFNtq+vzSFO/
xIDF1NdrlGQXO4S7u4wQtFSGVgCQnUCguCLkZkTk9KP9UQ/CB3WxbbqotqRMU7ZAkExlIdYWQbZ8
GyzxgohT772Cho1unUqR5Qy6X33C7r1HNDrio2jffu2dUqHdVKj0bqBcS+HF1tK3ANbpagaAJt3h
7x7E7ft6HIhWvnbZ2p6a26yHTM1VSxLY6xrw2m+rlWowv2wuHtYCFedteZHFsYF16bUpebD5t16B
CVkyWI349O00pxEF0/3X5KWXaSboU1rpA0pyvpJm9XofqeKg6gwcw2CdNN7HMGNYotPxy28ddm07
VO0D8FmlWUnBLWMP5xQxgXAcrTKoIRGddwm+5lgmHGpFK8ANxq9yv0xZNhgXcymKYMqj+Hbc3aCN
V5B2nZ8Hs7rjxIWGb8Tq5wJKrX6HmBNT5f58fBHses118hdKuxbeJ83Fb1hSET3mMpN251hUArP+
ZFGuVSYl0JC82fRW9B8iSuDtnDhmylDsLQr+U78vQkocjnErBn0RipcrIUPicgObImvTLp5VTHlN
pkJizakhW1k/fdYEj4bE9WtIoEHo3zhBiMpRBUvxB2Vu4Mm0rpT6BufmQds7PgMDdy67nXR1QXta
Bbnd8AZy2TpOI58+OjLOVtF/pKXbUoJmTBSgCfh7wJH4nQ5Zvr5xznWOdPEeHmYSSNTSQqmPz33K
IpRnWQ5j4qENIFKjGhbIjyugsY60s0davh1kttRsi18PbazEQVwdvjveKzIYMW5XaUOV7Rr03mVq
eS8xV9G1U9f9mKho3pFWBv0XY6ora8W8pgku18nmmWj73h06ymh0rEgCA+tBrCd/po1cmGZp0Ihi
6ItmVKvlG5A+A1n5vKBah3UyqBMoOR41Q/B2D9QwRQonY4YrKsLONs74O/g6kBkJbdOdgMFH87No
yrnHB3N3zt0P0FSsl1QVdcea9E6u7CImbXd7NF2dl7uUp7EedgVU5HsSVzSEL9ERhGKhXR46cZqM
vhByGj26o00icoiXPtWhl/LffwIUbiAj0qq5tZpd5+84cBNmBs5YKrC4wsEIfGcAe7Mvt+kzNwt/
2liqFUO8ykg/y0sNWW2LplUq+hOb3AC1qkL7X8vSPC6jFKw8CaKN4EbbBurOSv5ceYzWVeK5Wkan
iz3Nu0Z4s6Uraw00esD3+pDqiLJ1FavkxMBiPJnCJSVdPla+bKxxIP01aBqnYpPtRcmg7fXYHW7s
TvJLW19yC8GWchCV3hV1N7S/ZXYTG5/aGQ4UMjf1hOodP7tosD75X9aEKocCAhCAYoDGCCvdTELH
LFTgahKqLqt9pTbIrviYgZq53zgLfTVd2bE5CR7idCMlMtM7BUlxomfbBPm/mJp9yLQldl+icj0K
QCAwVv7CEBtb+MKpMzEnQ70dneDPqKKg4ZfGQcf3j7l4KEfEPUz3444THvLFFIDP9Qof36/W6Oz4
1pSzNmXm9urC+PTFBf7gXjwZzEBhCq8arBsnaiNZFm5SfwKHbTDq2ZlQVQwiTgnz4E4vCkD6jwxf
C+Bkd8KrjKuJk0PvjK8RpKs+znjweypK2DM4kfNis8f5o+WSKlL4bu1PlUEAkECA1Mcl0H4kOUrl
fSXJb9XywRGQllM1o1Pp1NvTq2BRLqdYk5f11eD/z8FDqGxWWKbpNLsPb/TUDo9r5YPQu71Mwzpw
ovVEPnuEosLAp7gu/OHGrrzNLs/2uWE+/GQAmnTQH9lhEGI3o8nd1LomWl2eHqSbfhoHctHDx2mU
tOqhAxbBftofOxXm5qhKVajBVUYhOHLu29tJiLqMEHSoOnhWV/IJQqQNX+VQ4P6dZhxcdhgpLtj4
ge0O90av1slDNB3lpCsK0h24VdfjeZfnZxVypMbdnXRK3o/prHYkpVDQR+dUYskdhhnwNth2slon
KhIdTZ98Q7rk1dnXG5UY2L6C2FiUt09YgQTgBHRy+5E6Lu7t2FvVtMqizkxt1Zxtpvl5xQEl1rM3
M/1JvWwjt5xLcQPR6MEvWIc1K8OtFFTWqbP+Bq2MNZvYRww40g1izZX8A4rVEJ4uVQORfqefZkod
B1GVKvra9IqjgWbSnvzm3/7k9ijwbeOfsWqfv99POdpc82q/ecfQvWf0UxGpCzu81GMySAmK74Th
ypdB9oSwqN+nbyook4FalTKUhg3MocRVw3/BMejBNVKeRgJ29phUz/9YwnsT/N7+ttfvjBSdmT8Q
SRWF/QOSGQEri9zVJgjdDkVz67WvrExr4G0AUZBr3/6fOy8H49hk3jZlAWKjMSFc0LOwc/lYY02v
Ur3dzrbi8roWZ2H2Ev7qwEgZSHd7oaENeOpxe/717WIfr7KOwWUPD2RlWJ21p+pasrJz+b/j9sne
NfsxKq+RQ+pN+RqsvMJt84qBFp+bw5T6nBh767QR58Rrp2Tx/myrpU84vUo61OGsnJrikf5AjJM1
U6XCSkERoaoxGtFrkmVX3A9uv52goljUy8wjppV04Id2kLmFRmbPn7NcFyO1NwafIyTuxlWKkOP0
8n4uDZeaRq8t78qaUJVbrUu17SZWy+bl9Hphg0Lw4Y+zStgdHWwjT+3ByjH89HXL14GZ1WvUrip0
r2hUkFR+JwogwyPAThMXoCst8I49z7yGjccsuE5SjGH/zvbG05kq41u73yrmpNVCtY+htZ+Ky19g
g9G+M1IR6IqmyguQO4KL9URR6GIRKOSEPqyAyTaroawH5E9S9uwAQVxpv3uz9yvb0AtnGgv4ePAO
78IZMCM5vNJCgXLXysnXfsSfDbiENGCeIvsQae1wvpgtfcnkqjGaGh9jf4tbguWmgFH/FaQZGbTw
IcaOe1A9yrzSa8Dl7cdIhRA5xJJeqCwhnv4ECvhiQB1urVc1wqGWQ3XxHAyHGoAn5UcuKbwAKAzo
G58Xl0LTchjyuE8cWswRwDa+w7XthwoARPZYp0ZrQVUwZC5NVnvoZs4qq60zgJRUBjBenDxPD9cL
k2RjKpMOzGkjn/xnWdZGxuOE+7tEhUcgy2e72jLT81CJOsHmBrh50M7gp5fI/2wH7+7qD0LLFYTv
AKClnSyUpTnyqfMe2LY0zSD+9X/1vv0PpYWv30U4lFhJ+I728uP/zhSvqk7mvdyf8iexpDm+WWl7
+k4o6kJ/0g8taSuRKzryGkNkMpK0wPLqUcC+rRoM3nYIgSCYe2MQPv60bSrai9A++9i+dfN0FVsU
HZ1KG2g27aG37tFCzI9smxDZF3je2L6/uu/YNpiuVZPMrknhL6E92aNMG4SXCo0/a1Lv3RIdFQK+
jgadOa0e0AtP50Z8auOq/NU3YezpyDfUoKA+OJoaGzAx5mOf4uqvi5Il8YeuAnGO8qLGTSnbbXnl
qgcCFn6iQ87pvlb/VdTDaXfGrrrRRKZJHYW++ofyOMn2D3RH9/nC/zyJcRAO4/f1yz1EagHCIqSl
j9Xnd9Fh+SbIEYmTQzOS2yzTlwSh0KjYe6iDq5W0GtRDtF95ldL7+ui9YcdScrqLlrqIXXOCDcr0
rKADyk6gwVpzZyPtEMjbuN9C4utq9hE4EUN8W/sNt2eRgwkhK5WqKLBgs7Xfa7wRPGOcYGxlBIvz
i8UPuC0/SeeTsLMdX6dZ8TFxn7p2HaxL0kc/DF2cWeC8VoKcjVGBptYALULPX/2jovgZFLdYPqA4
als8etASsnUEISoccmf521sFwmvRewHsKH3jkgcjnpEzLASQLmlHWidE86rPTUdah/c3VWXLRBJl
SZW8k0cHWWdMlySt0VDdmO0liGKe2gJeUy1tTii2lzlfaj4WT19UHfBWotfvOG6YGEkvCYwoavv9
T1mrmnDNpa3FcTzl13K1ObThOlkNqsOHGdhAng6tNUVP/wkVdFFFqnqgdwajogeIO9NKN/uvLMdd
CqJEImBySEDVwv6cqNuiSUAe2CDT6lhO3slijXeZE6N2SJMk0Xeu0pMbPCJOnShkWNgcQAYITXAB
6D8R4Ju8Y8upSDMVOAJlFVPKTNf5deMVlv+g7gNvIanXDuh0idMCDFbZXfM7iF6JCvfd03KxF0+y
sXV5Wfyf/IEafaKgByKcEoof69B9JMuORzZllVK+KzRQpXS0efL2+BN4V+nrV5flmk7p/UW2Z22i
yXmtsgYbDYW+DQmLXEb4M6vzgIddPkeU8kbf9915tZcEcdD1N8WP03H2IjwvgtTi6BqtN+2fAfuL
mKg0Ias5n+fIZpAJOe65xW0+1qiEFHSB6VBEdWIgfHHO1r3VB3f8Rp9oRpJd0NyWXn/S2hPRNMIU
zian2Y41ZrExBcMMdNsw+XIKSw8Tfa8p75LrAU17aorBYBQkHaTScBdyKtj33dUhBxw5I+dF9ZXG
O7bcTESyMTd0cAPasqp7Zz63QZgaC+lSOFWibWvNQE54mcvEen/4AgnwAZMOpXl7jblkRi+0K9xT
8CoBT3LiM7JrTSbqw7a1vGbe+RKy8Oc+Vgs4NXKvvSqi/oF8V3mCB1Blr/G5+qGxgbxE5CTRE/E3
Z3FVk+VwtI6KhRXdpvZW6JyLlqrR93eLPdAFGH5FM/8V6npg2RW5pdduBKeB/1K00ZNFbEMMrlXe
F1mPIE4FlfbA72OovXf8ZHWaleMCwg+xR1VI15lNpIp69bBPuCJCRx/3LnC5kMwjiRh0Ef+BbiSl
3E++ASRDdAP+CeLwJIBdcWcphQsOMBSGmJM58mU5g2P1KTJaAiR7SGEvaoSKDbCwMR68d/V86GqP
D62uUDF0pKkvh/6U3Yh2EufwC/Bo6OB33bi9QCIWgcRCzfG2rYQI8+Dm6RGpa3RyZzs0QDd5KxG7
tSdFvL6YI3+GCURxjzgeixNtJP4TOf6R9WFKrrX4Dl0aDIh4qVQsO9P7h4l6jwpFa/4UTVVeIW00
zhXzAql64x/ncvODKj6XSxDX28EcGbD+QrOIO5TSg1Lpd6lZ+HBO/ndYAJgat0a8k8DS9/UTSAnC
717wrZtLqAy6yGbuNu2mWvss4z7yFZOj8rNXwgw8p7WnYZGCij/u5/CVxF921eEUQ1VTArEzZTby
pJDYeX3B76aQIXgFfVjaxKy8A0OAp/9ftoLq/E77ItVfJblFzMVA1hLID9zvHrHmkBg0c4GOiBT7
xWdcCD9NriM3hP+M9HPcYD9JQzxQUtuEPkv2YaC7qTnzNVUTEsXbpdRuFMsg+ci5v9Zq1NDqhtlv
EzgozzDwKIe8ANcUGHv3Kn1w5hg/5izsh6B8Ex8vGwilFP6IFcTRZhqCilagi7vwAvEznDAMClEd
zY10BPiUH4Qz5GLeVLx1IjdeVhs5CNQlb1Kv1I4aBCvHMStmYY136igBD7QBRn0NK3MqGKR4gi12
C7SWV6Un8l8reLplL9Wx6yOsO6W0y2npOMkTFsuYc66H+Um/LpX3XZRlEK7uqzg6245jogoVcM9v
7TARJDHTkHFXupuCSzsVNBMc7l/r7En6EJENaf5EFirtr3Q+tn0i/MuVJNruGNYpxMaqKc99xUVi
rdeow8ZEOjKsh/8+dSOEPh6Lf27wyQXWLClk1PRmM2Nsv1yladNH/W7IZELQhoVyUlnfhPhA3XIg
Bp/w9LmEBEtkGy76Uzlplz7w516WcqGYykHUEQWuLxWeTnci97yB39gg9lJM5B9impSta+yLIK16
IgFFGQfTpXUsQ2RO97dv1lJY4y6vaXwjpAwWN2mHy2GZQJgaqmy8Y+6tygy4AMQRV8Ka2Cd2dMLM
B6iOEC2liqb2P4FPmHTN/JshsOzzk9z7oi4+LRTGw6pAXfo3Z4gcL2EnReWv20ky5XM8jxHa46JK
FLJoO92ESBDoOpt2Ek1b8ihXiSbzT9PC3hbS0pT7QUNECQn+zxvRpA0AdIB8jd87K16z3Sqtq7nT
py7kupyj023bvuo4lLe0Ce2Edac6QuBJeJIGSZdFuzApK84Su5gFGOvdv5bJRUCHXP3XabWcMzt4
Qa7Kqjg60lWV9BdQzKTgIIziZ/jYJlrQiPEAPibgRpK+GJ8LLJK1t/qVt+gyDuBrLFWxe6lGa4jP
HzUTSzW2StzHIqd8OUuCCnFgnHbUI+ePs92brNFhnQfyZ4VibFOTd9O06pG0z6gGflcOS5epGb+F
FRE7hV9arW122KrRPQUbJIFBfmrpv5RLp04KKA7Xsjbix9SZrQRbKVizJfgNZ8F4cc3o9pwLdn5h
QLOzm+qRURONOeKWi2oLCQ8sryuS9rN/nguYY8lxQN65nZPrjDpIZUb2xytQEZNch+rvOmsfz7LN
Z7RvzrQGxEdcUguDIkPgzMZI7oOhnHc0n71sPj2++bT3FzkcrLYtpwocG54LkwMncMdnB70PYgzC
PdvSSODTpj6+HtIQNH2LQX61kO6OvHbmrRGAbGPctzpBV9IM+Nw8ypjqqUieby/B3XQgEn4hua3Z
IMC3ZqFwOlfUTMOYQ3SoPKTKqQmbg5eVcVokipRU/W67z/tJ45pLCoebdYPejxKUrp4qhLBbWcNR
+ojASEmhTQg6JkH4apwqxyVq6kr2K9mSFpD3WqTP3j8+KQSK8VEOJ2WoA7kFVi2+tkkxOLw1GWKW
zdPcIj0cdBsZ9LKOrczFq5DSOTeZYjuuCzN6Psov85O9OnvTgUs8nR13yQrICBrTt65zYTNUEFjo
cUUm1QUwx8o9vyVvg2ur7tV98UYwSk7IDvx+oGV+MXAg6eFb7Hd8jSb3D9moidnjq65NcY9C/Mhw
e07NOn7go0+Y9xK0QZREQs5qmJRiXZDPrbJ54doBcAd4RgCT34+dPFFzjaHPBLvKWG2C5r+Gu3es
p3sTlO9FtorF/hCNeZQ0Manbx9V4A+oCRvJ5OGJUUXOw3DTJU3P3sYkNY5ygMDowf0t3e5bCwsGK
sBLwxz2E6RrM4/09dZ2S3kINSVLWnIbTehb4XPe4c5li/zI5JkrGldYFDBiY9v8xpjLfyJ1fHSWH
Mfh2v3R4ipaKZTLfI2kwDN/EZyiMJgVcqqY4/vk2w8X0Xi6aOr8wDvCvss3V1VM4XmxKgp0z/gPy
8mWZIsuBNp6EIv9zqwz7PamIrpuRVS+jNqoNvsCmR2HvbBRVwyBO1lX+zwPjDxjcdJN3DvdoxW81
SsgrhqEolPAALvANvmkYd2fWUaFyyxLKoom77Gx7DDB1XJN8M3Vslbl5j+2Lmq+eamBwDzSk2T+w
DF2gGmeuqEDffjuQQiSWLbtxQT67U97GTuFa58H3/CQa+yg8gzyJHJzissgGsqSep+5hSbsxNoUP
ihfMwVX0ibXwA7INn4eEKvXbAYyZcrf62XKgXHfWNxcq1k2rCm+ra0ckxeN5OhpGGHHp6QRliTA+
wx2tWZLxfpRKtc/+3+65QzbeFmLw/F26phZskJ5N+RFj9MJtUOsxuQG9Ny9ZL/Em9v8SFT0MimeM
28I+vNf6p6dnGMLV08UNW36zfKoqNOsf/qPvM6+uEkb5kCoafdkAPA5hQnmuDzc4lIMcny3rBfOZ
Kp8O52114LihioMjXh453TQ9NBjQ3D9CW0NSvWveNd9x5Ga8EX4aGUj4uRK/LNl6FbSgE2cXiwB6
6hCwe93eURifYI2MpH5UpbnAutTft+Wpu+OgEV4KmD7oAFHqW54NULzbaWO47rJx7NStJ3mOzRYn
MJcC4Crd8BLioWTcdUnT66PiQfoUDC5HGvWj6DVNz80r0rik/C9hpd7kNpiZmu5mP53pgQTah1I0
rjW6we9PflfzQNS+aCB+nY1h1+YfMcuwG1MGV6Pt4lKVxVHdRbTno79v5oSi8FZo9q4emVVwSh+c
oICxpHEkxAfhVd4wknA9baLeHpKP8wuajFDtpaLMEkcUHCMb5n5pdSRtdrX9OQMPCw0P1Aj7F7Mv
/TwMWOrMDapY4IvS9dmKHZyF4s+U+Pb3GIYBueo1SxN9Gyv0fWbtg60YwoNc8BSNe9lBZwzjriFr
m6hke0iP9jp4FxRKKthLIEfFEW4X+yCLlvHNl3ZKKGMqUZehDHMzZ7P1j4VXIHHSuGoEAHxh4eGI
dsZNMioXAeRxvCG1AooW1QCpzN1BpUlII0GgNXAtPwh3gM5aSy0XF8dL/g0zNJ0/i02PE7MR8Khg
8DRDnCYdqwI2p6edHKH0bSRJ8Dlsa0LpkJwi7M+xwmOpgb7wOPo6CnPUQhzI8eJncis3KHeThDL8
/Fqc8apYrNZDqGYQ3acoYKfQW7AjC0c01nFD9uj26cXFYlhQC2EQrrE9IGNcaKba5QzMYW+myaXV
iwo4G2MoCjjlCHeU4fb+nGCLWMmeAlVcmaKYeRRWyTtioc7iw1zR/YqNEpReYPmbJ7jRkV3740av
1gx+jNs8apiQlQZGM2lv4EHAXD958Wcn1epbMDBUKwXXAdYRR8+jmBa2Ees2kD6OLlN5U4CieWDg
MpgCBWkg/1y8DtITHuV0bOktBJhf/eT/Vo8H2yY7OjJMAXKbctzKG+S/+xfL/8RQSX/u2dAI+LZb
wgvsSoDIiiO3JItoc7lZvanOxorEehY7pfBqmrs4OEf4sG8C4/epWFidV4XgOxFfTy2FJP7J3jSU
baveCC+NheiNJkEIdJVP74yl0cWxWxP1ZVHbk4SPtFc44dRDgjdc+DF2+7cun9yR9uhmFWyKja7h
x5mpb+19COXl9qlw57ITC97c7auMsuduQemG+Xp902C7rdRMI1dDHQX2XPP1Kvymn2BJhT65V+2J
qnAtVKDq1hELBNB+lrPIu73p5PYFP/ZRBmt/8P18fBSyTC6FdN9f6fYEsiHz8MHnJO0xh5WDUFh2
ZcbkPNppVUpSdAdPCwPF2Q4K60pjIXSA9Ndrwf0sUItAKFkwsRXIVIIivJ9wWeNNEg8K2wed4GFK
juBl1eA+muLw6voFP26GR4Fr74c0al7VfYP7CCbk6A34/VTZpt9yBe45V8mNIZ7tCOOrb+hfg1WN
VLJWHGeBy0v5gr6d6mYcjXYa7Vnyb9vgOfLBU1Q1FzHj/vrdg82uF2Fn6seJO0+rKm4q5bosGXtx
yrWA/2J8MIfkXj4jHtwd0IKiwqweqDHQh3yblISr2ZljAG2xrv3/oUElNoiG28WxmgWphaLG+ADf
cU0QbfyN9BOLASwKUysbYebo6NM6G+3kIo7/DaqWqnO/rgoUHhR0YG3UYs91ncHuxrNS1vp4ScPg
NrkoX/XZb79HqrGNsErG87mVYboiJNWbTpUcXXrU4ue1xoqNT0AAA3Ve9c3b2B49zhe1AihJUqWI
zjMVGKJKODzCoW8s+483hjGT9kb0c+R+U5fPxnSyKVdsMgERszRcvozC6JJUv6dbb72Yw0dA4gjj
HzTxUfLgY2U6uzHkMY9EkA/7u62ZaNEgKgoIcY9A2QHsVyk0HJGrDgFllFboxHTHDX3ox4dyQU5r
0gkwLiR+SQiJPa9UctfzVQPDrXLrZjK0svJIqHKYzhEZydOGkP7UpS2dnry8n6+wc33uqQRFO4zz
mERmCbR02cRRBN4i8VlkbEnFd014nJQsN5B1iqTFskD+BHRaO4nNPGuSvEKdZCv8Q5BfRflzV2Q0
6ap9yXxp1TUjp5iaz5c6s2/qcPa1/VIYuofjMv6FYoK+n2ggIE1lAuKYa7lFWqGKt6UNEtpFG162
nWwvFM9YtfZ/pdqQtSHZl3WijLQ2sDg5niYvTXhH8c9KUtwVjTQL+TPWB/aStusUwpzC0GMYgTnh
N5Nl4SHnoRUtYWbPdjAncne5oX5cQ65b6MsLSBnUP9WvmGT87wtvYx5d/u0MiY3B5UNdGaWc6dFc
Xrz/P1Nl/ljBSqRhQaXlvUSepqtiKBtUFmairfzrCw/avZ93wYWmHD2ihWoLwfRUOaHpznGPqgC/
vGmrdY6foL1DBXQrBCHEQ7xNW51+0w+ucPR7QWKLX6+BwmiZ/QaUm/Vr4eLlyEzoQ+I2FOJO9+Xm
CPAgpDpz+TOKDg0q2DpNPg88Sj9xuk21MB99C7pr69zYeRH+UB86IlxgHl0KmNKMORb2DfU5NUkq
vEO7T3WMGMjbC1jNVGQ7qqVuLQ9cxbTYWO26wkTE2cSpB5gvpNSrd5BBvhXFpWqbEEoIN162lNEx
eBv7K8NhLxqrCTKRgBoR0DqNhQcbAcsCLZqH5ZsZCADIgPvjMhx7rvPFdfuJMogjLLgnU+f+91vz
OeJO+KPt/nRzQQ+BXjZwvDXKlKuIKtYJ6j3JMIb+UCqkg3an1k4Ru+GhHbExtfIuThIuWDVrRP/5
ftqFbgGfF0Q0L79MUoIjtvkrYmZAL5Jj5w6koSeONn/EJD3onRMnaNPjssSHR2fh7BgcwVKLaiDJ
X/KzSPRm3DAAcssRbQB08tGaWmenOY+8j3sFAaqEvO10v+IO4mwrlW/t20eXa/exLklBkjaZ2Rvr
YcyVmdb2pdnUfMBv1l9JmTL74cQmyImMn1Yy0TQ9HLBKzC10n3ivfDHm+8GR0pfB98HwZAtTa2rg
fVdDmpJetOVkSvLwgrxa/pc/5GSvTUSlc8yTKZ0VZSBZdWAD8Wk2Gfkg1m84I/olVGPDaUkBy/UD
0a/M9DM3BCTEzziPWR5r/em58nDv5MjF1mr6/s9SIweejrqSm1k/TWYuj0454tzQgkW9v5Bi9Tdb
UkhkJMMaTyHizKwfogK6Dz0Q3oueiESGjBVsgBwA9EO67/bdhhhr39ZOfVfJXry9lOE3tq1hZfXL
6RuMyYqHDbqhixnR2G3GRHPgexMsEDjKi0py5xjPktSFb4mVGNHa08zoliqvqEKEuVDX73C4JC0Z
yCpld2/JQMd1bLFe5h9EqTBJA/LgiyD/8rQvkGXO/2/SvH3ARCXA540WBRVt76iLu2NMgK02bP9X
Xn4+gFLrKDtd9E8qjCD/P0O5SsbZK24OHq/7QnyQImAQR/P9da7quGASpnDhh6l7o2wEAuN3QfA0
iHkIt69iO7DcoFeMnHKI/tyn72M0Dple1NkdRAPP8+zpnOHOuliotttRAve725e7IPjqvJXHGjjI
MlzhZynkHbKHAShqbvwrLqBnBBekSlhtWK8Dr5EcxLpBGAEp0q/meqpNezlJOWKZo9hPKgBDmn0q
NJ3KXBw+XY3HiDjgOEmktPVpAt1FMbKQo51MdpYVhe+RGIHipKbRCsixc1V1i7QNSD8a0s4kBR8h
cEcIZsKCAOM6bSrsNawJaa9Ff8yHi6iV3kXAfY681bktWLNYvAJ/JMafk8Eq8QSX+Iag2YtMbVGD
j5Q7kP1yeqL6FiC+NZQ9Lsy8NyetJjEkGyE5FnFdYypkas1C6PD+XAq0M5sV9d/Pv/WkLdIkQItn
YmFp+r88w8Yqy8FRhrPli2qjFqcMEey3YU7lyOJeWKqdOPMO90Z5mCU6kCVUQWePqfZjTu881NUJ
hIDRlp7vu7JvONI+GB4icxZSOG2uL9EJSFNrSum5VQc8XCZHSArj9hNGhAs4y4PTtbdT48nj0lar
DbuZgyOH3dPXSgkmbYQco53Ncpy5rm1Nv9K8xfnWrfMfbxkJYmrM874w7xJmQu8TGKvhvCjIeCnZ
Sa5kHp58NHIJ7gwVWjsxX+sR864zjlpUawWGgh/yYu4ozaoSxXE+IzyrCNgCyCfQw6nEhtSw0CwP
IW+yNSXugkJriPvas22xRCsrSheFLeUhHdyT5QyuxKPPKrZBS0rye7z+TdzARMXHv+9rnx6JUQeR
Wu5veWRGMQ3f7WPqyQcuh8FSfjW8/7A28/eKk/TjEKQF2lW93P/4Io4FDTsSZPofvKisYdxAmwqx
MIVA85APZPef+8u/+LpHhFhGyQlvpzJ285xCLjUP2BEp+bHZEby+h5Qzp4z90WcylAkbdutmoTVe
EODJSP9y5uEBPoFDoJWwfOf3LMRhOySCtO0FRruGrvLHGNiLczv8szehoNYb+kDakMR9V6VaL8OO
8zDy/49zr0RJmuYZ4pvz5wTfA75PflDsgyE6eIw26phpR7qoJs2gYJX/6FgeGwWR+7/cBSUMYvur
ciFeqCNVyoFQAyZXlqIKN2bdfKmeVtahSN9UgfqhljCHJJSsw5sOErzd0u7nlNoK8BNuyDH073qW
24eo74UW6s5X0TXfpQY7/mSJF2xOSIw5wjpJ0jHjtxA9ZuZ15PDMW3Wcv3MCP+ZFYY1NtVXn2/YG
QUQwe52L8bK0bAQFpoBb1Ilcp3nUIZ9b9Ynr1sW3Xq+VERPuoWaCOVRBAyrzDCd59CeXfqu17I5s
obfEZbf0S6iet0AQ8Tbofo0oJ4fRfYUMAXv8h2jGzKEA8k1aUw1svg5Hl/EqdCvh8CMYxKxZBNe0
kmsKn/0Qbn9J3Mj+6QrExqjq1XBkeMd1Dr9NBphn6WtM1PnWpL8mkU1atzZqqAQJD5H64SyzgKLY
ypkOEakcnkrbsl8LfHrJtyefZjKDYfivo/K5qxJOY3n/xI8qNfcu5+0Tij9++ia3dBOK6u+vI+9o
xxHiiNCVQTBZrW7vXjQm55VQS7jekZg3uh8HPjUt5+AO43FdbEFrpNeSs/n7X7G1/slvJ+xxsSLU
V8xyr4i7cQbzFyoilpQRzoihEdeklGkw9NUFxQ4KkXQ3wNkmpNAasoOW0PCOUO83SIv8eDyuLjRe
AfsSjMRSb9oTlA8Om8bplrlv70FQ6RCwcM1HXb3en4SxN+e/p4pdNgP/TGQmuDpDErTAqkjj7kHE
lU1JP6s38LPMfuzUKbBbSxmRF2uSiZLy+pLrxmUgFUTIl/oEhL0saEDRvUSQf4jGRpHhOxWYYgPP
IVqphccJUjLAJgqzPHcH2A8gvjvXe5bPMR+Icsjmf9v0nHZqd/qcFKWNjQVf52oPm8VA+WSCLvxa
hhl2aYPIfhYf4xsYdAiOTjD8hsFVIeKlmH25NHXeqqawIzRn7xzgHrUIcvH4FR4GUJ5wBt5bId3F
G8EolDs8j7oKZeMSwALYugeye6DUtD+Zpn7DirmcCBYw42LKx1iG3ZaPSzwTDN01jacQ9DWt4PRj
7/U3g9BTvKahIXzMrt/5ocYgZeyhH0Y0/oxkIWsDf2+TCbe6fm6BbVU7Zy+TwypdZF/U8JuLWrGd
Q4mU+kMfDvzJG36+AYWSgjEu+KvpCL2cl3DyatXq9gAxAOSWRWZPBXZGskDriGd1cVTi3Q/gUYSV
fZF0IWC7IBEsA/LPCVhqLovDoPZPmcMG2QkKeXQOBbMTUhNUG43fcLxrZ1hNSs+b4qmY+7mqwJnh
0ttl/YDiEmDdFzwe1zu7XJg8s+807k85NiCPi0WlSPVigYicpdQ01pHymz8s1gJe0JqhO85QLdsX
Ac2vGEjqR3eGmUtPVs2pzYRXD5wNylHug8AYBwk0r5Wv250m863iB3lRpCEB6v8TZ75DqSBpeeQh
gWJ0An0iLXSjzCehQ7UmlioBuN8u9Bqn52kTGXaOGiCMuCeXuWP2lhLAi9vdX5/3JLZsD0IkH9AF
csteprntuUBM7mJruzOe9fgpkZDSOu25qBqPw4XlGG7ZMuYoGZ3C0lC88TlZVWuJtRFEUcZNYwoM
VMnOr2I86zcE494BMtuAYHhiKcljLuIsibWCdHrIWPJ+G/t+0VsRezvOuv8NTNMQs5IloAMjieTw
RQ841n/FrRO9Wfj4OQj31SXXr2NtpQwvRV0IvTctMLBrXDK7YvHZ/CDE96UiWBRZzl6tIBj4JAfB
FG1dRcrBrlmh4PmXx8ZGa+kBiLykXvr6gP312Pe9R6pq/SMr08uR5E+effmZlWG7b9jZk2dLJsnW
QELD1JGyZWuvoGdryaScbe85qXAj5ycqE5YDEjDpxcoI9ZcC2Ez/9mG1ieVEBRU+ISHtatvzCMeJ
AaYKZKO3YCeykApGRRlZjDnMGZfpq9q/cO4yAY+BcOhnlN2vBinu+SImpwu/hP6O2MfwmpsS2hFU
CAXMZALSVwFgx9JY/8iEseb5WjF3HV8kZlPBnowngDZoeg8vKlIyuXQ2FqtVm9VJEElAcpLMni1j
KylTVw6WZ0mJY+Aet60sX8hmKTNJeoPZ3OGUUY75EPVG2aP7ZanMwjJTDyyq/GMmE6jNa92cgkpj
X7JUiUVx4+4yPS96q4r+1glHz5xarVYgY1eIOFnRdS4myUF8ze3tX75O+uPgVot8ZEVRSaQfv/uS
u+7bh4zqZ2nE5PeqSB+zU7GooUTJ7UzdsKv+PS1cieULqrqBSiv0RnMIUGZ1eepZIqpIaHCYjipd
PaxDUQlA5V8eLVtCHnKfniITORQ9z5Kk3rNBbWMzWUy9Bq+Byz8++E/XFIkHtENOSQgcxefQZZu5
NCeXw1g09WA99MBhlH9F2Suan/buDcBibiWexPSgOtpMKc/XtYTuvPPa5poPTnuQJmmgigpmaLyw
7Y3yeiNhZLq2iwbT5+1etBduAR8Pa4D0UUAMXngW+1M0hmmZJrkAiOnsAfExsCvFtx12N8wSV80V
rOcOvz8Q5KfKmyoOv8GaIbOIGAxsJisTnuVEb4uQFz3YNsHR6Tkpntn1MiiLtDglDL4p7c/weawi
5BywgeiStR0N5fecE8qjrAUnKAIO+dMPDHV5F6TcjUKk/rZ5eZR1JeAtNrsEBaiffKaRkG9hvSSV
m2C6sWdX7iKq5PNTjmhvWc3Ti0jC6WrnGeUmZjDOGETprBQpADv1R0WywthpJ9KipOvkeAXe/1kB
zftLRrUWY3Hqd3sGBEISDBGpdfX4ff8xI9ezRsTpkkzHmOi77UHR90x/5B+lMSl1ApMHOKoATP6H
73YkmzXhRd/lv2ODV+IEq07yJS008VgrB7Xq1KZefjWZ211IxpXELjH7LjeJUILhLAr7ygEYuOq8
aZykmXqQTqLeSH4soLWmrYcWcr9kzq0JRpRPmD+EudK0fKj4guGfA0BsU2p8SgKivMixeR8FOlYk
/qNaa7Mb1sPm44OgkqgoyCsnkPsnQ80cUS4yr/9H0ra2CyM698BqD/RQs/6Um5JVp2VraRLgW+E8
zYMAltGzysTw5g6LXBLm04s5gb7woPkMLcTCzAcG92YP9Drsnb+HTOsamVEWeywrr77CypjJGt9G
D1HlRDqAnCmyHAzGfAzjCSxmzRxiBf5PQIDApPNgRsJRUj8x3JGEO5GL4kSKAwgF7wF/JQZLEyv2
xZRpLWmynrlCu3rFI1urBPow91fWx0eynh5y7+i4vqNn+LCbn503YfRTHSdOPSsbmAondqSpjukG
m4i4Y8fU7W8MR27mXTXkJkV4cFNqmkShO6dL5H2IPq2ab7mtjvXh80qk/LycogPilh0s+LM7XW9o
bl99l+l9qTIIPT32KnqjsVFuQdlyzBN3OlLlhd4po6KUVThvp/6+DAiz3ljQekRG7vTsMfJU7AZh
weUL4tFoH3pOFfhyRtkrs3qolq8Aua8o6inm0ejC4HkGJXM4GtvoszsPwN44NTkgJguNE/qW1VY4
2Kqkt08zjb3VlZDlh9erIysUNZ0KpHKgR82t7DSQzsoyWYjFwTRO2OfvQnvY5IFBEnKTWSEZ1WrT
iwyCoM75WqGdc+jrmENox2mKEuKiKVi6Yfd7AO2gIHXh9liC5/pwPimgIgr+V6htYPLpQPmeaOMw
zxRq2GZUXhXYqu/1b9QMz2fzcO7thu1c1lx7Zfcca93d4gphAGVL+GDq05oidWCG9EHHrGSCe1+I
6+XbSAv3IS70X3CMUvAUY92Y4sLaMLFGtSjaExeNRutB7bO+ynw3G8+K+xj8cHqPJx3EPNAWH9EM
8Gn8t5FA4xQ//WCqazrgOHSBaFqsEyoZOB9YzPuP52JoY2zWzgvITdo1EMfyCuLn5TF5Ty1wscs0
TMDR5cLooCm0kBf6CCVHyGuQarTdj8ribUnz8rUDhPNB1sFNSQb5pryhNjmPT/ykXZmlRgU//LKA
UCZ7BoLThFS26eGdt72IwbweKk9D8tNmMvkH5YqY+LymKB/wppHBOVIbchP+FdA6wJD1DTGqZ2cA
ZH+GmYy+jepDTkJTN5Xh1ISFexsSBzrJfpcTVvkhoPFiJwyFAb97oMolMnkVCB7IxI3/n9KGqf5c
ehkfsXsNQIpv4N8RhO17cO0wtk70sCdGGPg8/AaZ2vAoISBFpRLyMzR3cQRgCa0gg63mIUrruDQs
NGJnQ5iLFvPmcZFlm2aI/upPYucbbVxgPLTTWgJHkmgxEllvHs4EVGSVXm6gD1S2Tt3FX+nEFed/
rEKFgQ/9G4A8sidEPxZJC+mKTlA8pAi25TOD3VgOdm5f7l2b8FeVPofJXl3dHrzlImLReTD1Z/o1
v+wfknuU3IZuMkHRx4Jpkh/j9vNot8Bd2H83WQE/LQXKg4deglVdmKeQx1Gv3oKugh3R1iejr8Fz
kLW6OdslEE9bxfiH60FYqEFMXLJdCoqWj4pbjLKqigEXeMUMGldtgncuN6jDxtXrxURc9Qq4x6pX
KjSJcmgmFQ11pFH/UV2S4gumPJNQ4JeBKtOFs7TBHkt60Q2aCsd0eNV6lVtTaLi3XNbqleFPlxXh
TJX5U+yRggW/5GFTsPvTEIXix2TaJrcycVBajoKZusq09dYi7wRlkS3YkcyEKWle5lNRr1VMA4mP
fHJXyRgD/WVllzC4PTLRWCWvIXFaZTQbNOjuKqCrvBTD8mq/KvjuRuqFzO0xfoxoMJR2D4eq49MY
KuncUuxLbFgfiITsgZxt7BViQsVtyEUDaWhQI+uOxmC7EW57gVLLyo8mp6g7QpY5ovBPI5JBbJ2h
35sy1WR0xy1T5uUtyEIVWvuaQvTYsByimJmbbFWSMIoA/oktK4B8CSpZrj7lxMV+zSU0fwtr2Mku
jJ7dWrVN6pWetSgNSMEIH3ZZuFpaWC3mYg3e5MdGgwI0PhC6ueCkNS2SE0fTRU/Y0dDkJUJ/Lhzy
E97aejECnoryINRdg+deNWyD79bAgBMAZYkS+dCVYfYnH+YUuXlVGKBdDBAv/pCnYsDzAjLIWC/b
I0ybjqFkTrzcy51K83MRiLbZQyzxBoNLSdopizrFAzkr6B+kZ7rhJTYorQOOhZzUJcW3vCHqISMM
l4StGHke1Vj3GtybNpQj5j9Wz2ML4KOISbv8NHa+Clb1L/mmbpNYzAhENVzmaJ+WMWUirLlHn7NU
/UiauiUt/9T/J7lowCXiDSy+t7LsewZSBq9GQu9FhylLL9pvcpU7k6UMiADMY4P4CgUxFLP9M8up
m5vFNGGLG8eW1NTNt4SVf7n8MjbCdMD1OY+DiPC5RG0TMQhyLkSk6zv7ae+3a72LRU4o7ORLsXdb
fpZlByxd7M81e6wJFQTlqOL90r168LVDDiMrjQrMEP57+9NW9rDR9uWlT7nFqMeKw7G9zNUVwXqL
gN4wf804lg3RBfs40yFpd1c8/6Ew4VGVntl8ps7ZrqDzZQzDG6STh+X6ZooUzMMDKJ2UqQA4xSsA
ksciklsOMxD5N81tfL/SJFJyNwVCoKh8znDo1VaOi/vXyJdy04lh/43Dm5ZPk/TUx+tHRzis+wrl
rEzlH3bqugI30Tiol4XO9+MRsaPKrjDnoo9XRIBATNh6VBy0tpWZ+b75Icjgpg4IOrcso/kXpri6
5ZqDsJImtVvd1bM3X6vqqmRd97/xM/Qn80zP4V+EEtOIaj/2r0imTP43M0H3zbwyY4dkcVCX5WUu
rC/LBH27aM39ctd6kCLJDo5fRLpaKPtEn+/rylD6ovs9v5d260xxcOoyzoCgggtp4Coa4aCyiZCi
nm5WeUYq4Dja555mg0OuCW13VD8UyLlDIWibV8ek9mcv3wuO4FwUxF9jxWqFtH36JcRFaTzZW+Pq
DuqAr/BtWb3KLvP/y9cDHUmfH7+5PhRzup+t6lRYMB92TMAD5/0bj4SmHSWBa95b9/iezFAhFL8m
viD1fYuqUlp7ebS1d+ori3Wxoydoi2B6HQwKan+K/+NYlopY1XmLv6Xq8kgylCAGjY8NtkHpnc5Y
zySLMeItpAq1cg2UAw54W7S937IfaKKwNV7u1Y6wUmbMpKqXZJCUodIdy8NlmoPaKHJ5nAuzn7gp
gFalvB97SG53ftNA3NoCtsRTDqarQG2tTQe5J/I9WXHU1VNPYyKsLncYGBkoXwuxCGO13/uQ6N0j
V0iQQm+LoP1LT3tSJaDLvAk6U44t4IZ6s7P3Kw1b8nsEu/tFKW5CjT8TUDz2vv+2q76cNLOIBX35
01x34A7zrSksSh2Tbe34UpoMfK3m9dTPTnu16l0F2sIncGIKbmIEx8U5AEYXYt/X8aUDF6nKdg8I
dXnIjgGnhTQvjR1NVAShjaJeL7IpCqfGzRKIMTOoHv4tvE15TRKRttdYr9d23XIMwl6RVrhjLitB
qBnk1ThXT/5abH/1A59rXkYnRZzmK9LvmL29sSouclO1RO+KnX/n5/6VeytB2Pw3wYyQLpO0zDn6
xRGPxyunSUvvdBiiq1poqY3pdjqzpDknAiBGUDIQSjhwfV2j67haIUnYys1z3Q97WJenxgHWRzT7
u6Zm/Ez5NEmnyzFlN2fDaEDSVhl1SwHRofA7fpcihO2PJHmInIn80mnNMrxpbshPH4uuIHwVu7Vg
TRwlyCc3Vnif5kn3UZk1jnOVO5Dcqh5ENpBTaUqzrkQsfJCAeXLN+3oVJxm14WHlsSDuFmqzl+Be
IwA+3e1N/vl1HThAH8a2vysVHXJZHpdnlXTQ2sAOl876/STjiUzXNK5LwRTCMhGYZF5I/Z8HgVUU
EXOYfTk/pX9U+y8952QqxU78czyaP+upQuOZNi9uUm5e8xC84Z/y3cVLWrMGYNtMfQQVfOpAwhyX
y8PWqvsUk3yttqU2mMO+8EZQ65mDtzP4ZkD9Y6fIMCoDLrdE70/+Ki+C4Lmnk2MFCj4bFATUhtHa
FqUq5TLMVAtrhQ5288Cy0MBq9hJ9KKaKfvyTprzwiovssC6UAj1HcenUIUSvaMW+05Tui12Jtx7q
AkQWKvYcwZ4kVTME+QduGpqikMa1mhFRHX4d5Hyf+/5qNgojSDWX7PS3xCk0x+LwxqSz6hbaSXTC
l4tkP2fhQDGBubyvK2sh/kSoBsI1bY+Ztj92XXzwCnpYBM8uvucavAcEZ/fn55kfPQW1D1B28BMj
4DUzVV1ldhOoqBLYl1DwLMg9GsHLnrLbMuskaesG1Rp0GlermmetirLN9UoYVCA9qs7rDfBcBRYW
IGi7AqrmJjbPsQFS5XZQwY+LzGhbkO8jMdz9OOuxXw+MI6toIqsDPJ60iy7aBQFiloijx2ORVcjI
ARVlS2MEsyQTX1Xh227hd24GC8iq+I4sV5hnSSumRTes/qKm9lEgugPrGauqeWhD++Pw95DYlA4f
tcoUZ8wXG5IcHFuMiCN389h9t0Z2pTBLyYffd/wj0i9RjCyIAWiGEM2Y/g0Fyas821c522nWtR2d
OJMNt17cx+dpx3w6Fd/aEBy2asE9y/AYzhe2+J99uEXgSKBs3g8pJesNvvQUUiCqKr9OpbHqu4ZX
ixDWGbPs10xpP0/PAG0uJDEHdLOnEcwJ2E3FBNxtyzD5lXAGMXHDf0xuZJ+sWJFWBC1x/7LJ5V2b
26WJBYeC2VyjJmty/pDOrla2c+h49JYj4+9LNlxKh8xD7SGEtk8/0uG+APhvykkgABZOYvFY9I6Y
aqZwueEjNQOrqiC5Z6+shZVG/zHohXr9+kkylpPb36v1rqQFbwXHTf4XckTlruB9FSa96qohi//a
zOCA+tdLD3P4aHnPcuGUodMDvchI34zwuvIO1Ppi/+gCrZYsv9vag+Flw3llQ3N2laZ/nT+jWC6E
8SHbrEP11/28OokT4u7/uMF9u+cQWkO+VQv47QOc4g8a7IWhMElzCqNistNUc1n3EVpfGRkB2W27
yyUOHvJPds7Gy/JsWXq1KDntzZUgXt3zxV6M2C0W1oV1PzzmyfOfRXWROh0Is1bRfK9qTi1VFTk1
ef836XJ3rYuC1N5owcd4jcLK29LN4QOMWEYQDaskwTBUq5hNd/3BTImIBHdPLWsOWnMbb3bYVE67
hgSUPC1zEEio99nK0XZvpS2IhFfVpzVwJ0n63ZY+7GADZSblxtrhKn5Lc73TflvHAimpaYhUNIAb
KIjtXiaR8Iv+Pov5yr86JeCm3vU74xTtcDTqDWBMWg5/UoIEKRm9jgBStBct31KtWOLZGRaIAmVH
oeWTpu7POnHgRbagh9NXWtfkWE8FIYZGz+/tbzNAGIuRNJGvJhnY8O2GyxutVcPz/xkRkNfvIO0L
B00lwDkHFOd1Q4gTXQy+qAVWPo4l48YLzH0ki7aZan3QAlbsbJKhqBEReiRJZCXOgzUf1w+Ulsv8
59HVRLLCAQa6F+r8+RTb3Alwfw3MZ6+Binesg/mNKqOIkYueVinzmZ9LCD/iHDQQNdBebScRLwXd
LXzVlQtAMGnWcR2Mf9XeAmzC0k7oGRRrQ6+iiW7JgYijZ7c9+bFEht989YE61Dv7zf0Xc0OBek7z
wBktMvMvGDpOvAYVJi3ZB8TA9u9At1sbNVBYIW+0NM+dOWb223AL2HyzcmIvBD2gcos22PmJ3Xe+
98bnc342V47JGOBSNuOBnbvU+Mla0fzTXE41EYFBnwsFsEmz8gj38UOGrNUEXYARWPSBiQTh36kA
k2DXZph4RHrunWrPbeVa9Dwfn6SFLnUZ3KkW1RVe6RKv2aDZY3te/Emup8KbSAcjh6r34lF6Ncwh
jtuK4YP5i8rwS3u0Ud3uAbH+jOSFZqgB9bXp+pgVA3wiApHBgOY9wBxF0epUTq+1dC9oxTyGIwgL
H9Cx7LMtEyQZ43hAI8I9nRPC/7GjmEy67rR2W/RnzOOhLYO9uuoydpF4uN9xhIwUmfL9r149czrN
sQOt9ES/h4zDPOyqVRUBrA+F5FwwJOVJJGx0gNngvDHkSNY0MCBzA42YH9VytYQmIEOCf5IaSZv9
IfkdExbBbqG6oU+ox/K0pLeGclzETsbWyQFiJhzo76ROaXhQQ4roczku3HqdzTM8uMz7TkexXM71
3nP1/Gr2wTYKBbQHtD6zXTysPFe9BHSThFnHeY+xjf3lxYxgzMB/OEFcffSZD1RMBitBqBQ8CIZ6
0eWH7Em5XGlj5YujdDnXsAIQwHJOdkNsDft1d9kN1WVqDykqteRv9FaTQrokY/5D0AxUjQcdTr+h
0Q8PxRx2aGIShM6pnB0tyxKOEo86i/cSTRvJ4UxLFUN5ghnYahKhO+8G/pqWghP+DndYxeoE5VHs
uyo0Hh+IryWbGRuD3s+0ugLu+4Ovd31lg+vmcUHNrAOCVRYgSM8k2HRvCFAmPHIjQVoN3wfGkKxW
OsrE0l4YIBTLMLAAqU+sDhwtjNFRWN5qQE7NPy4A/3caitxyeVdu0F1q9lqN6xDqfn9eGROjYtol
UCjgZnIruejC96bKZF0CvWFOGk6NpwNZkS90NdPTtQD5tcWN/qrlu7DmP2D7NmLt/4dUBAeQ5IaK
RcEUV8GvkntAoLJ+kO1PXfwJ1nMuLdNOLz0RrcpuBVMbNwlAlY6lO8w6rHrBL9Zc1R6zLgUoiQzT
/Ncxe0Q3vRgmodtmaRd4KxMUGzqC+biEa257x60HJKq+F51eT0CajHsziszTYyPOv+2geirY1g02
axg97jDJkNPKdf7KXiytU+gymAwT5nOY3G70NZl4DdSelIbf5ukC8AsLx9cr1WroI5hHY48i7lkd
7iDxVnsp33iKu8B4ih+JBEYbD4CjyylbbBHJoRGBv8DuoibmXfLOeebK9vo5wSrR4CaEE/VlNQvm
Au0vSh+yoPYI9C3xbBiU9SsqmRyyiBxYdDP8zNdQPItkRIKYOMeLnSoqTFVhQZlu4xn2gTH1371j
nUFQLSt5dGImfIm5GeYSSrzqLlJGF1EJrHdagvC2WqWr6QAaA3r5CDC/yfLHY3Nx0MGkneWfHunH
IpUqtewkBseiNG/xw4wuKw9HuNfwvz4gnGvwzd7cmMObFKQ7zBqIH1UA0XSIn1l1NOtd8Pkgqr63
V+s9KVJLpOH36jW0iG/ngaUazm6JIP0HuseTrFCQZNKytVqhJxygJlulAak4lb3sUqnebZIt4f0Z
3oCCQxdd7oqpW4c9RJpakusuxkgVdY7RhKStS5FRrDGKONNm8zz0+DPTrN+u3nrSxGoOEfy9etxO
WBIaPLQ88pDjJnMxDlR7KlHIwpZLEzj8qCitR6sYXRzdA0CYLtdiPDyMUSUjDkZ1cLlmg9y7aRbw
km79Eh/4151axkGZFRoqU+DktfX7sR/FQV5dlbHoJx/YSDt2K7SNA2avJnVfHlZfRqEdB9DAHzVh
9HG1XjgCcrwPUuTYFHpI3iipYNZJPdRbU2tsvSRGrsL1Wwl20NGVrEzVhEPcYCA5GhPE9yqXsXId
lMBDw07t+wSCPqcsNHTrPz62uf8gKkoYjI12aBfEJg1nwGpzKX/HK6aX94cx6i4h+KQ6SseX29bj
2DcN4Tn3xaPQpebUHWqsBmdvvU3l2CfgPK4k+bm7vWKq3G6lhL28SkNZb41T7NhLW8chvI1jcQy9
DQctHfdySZjumBxbRoU9L+lgdRB2YtKzPpWaPMIHPecQf5HUIyXTCL4IozvM84Lr2QKLSd63e5Po
IJXDtN1IaUTJbpiI9FJ771FKNK0C7V6iP/yMsZzTWPZ4Z7FNvAHH1k/pQ3MvIYNMowKWi33HZKW9
0fAIu8/DOdPhRtjlt/ZcY2yDNnONp0duoqV6pwhmdf23Tfj3tYWh4oor7PvS5nT6BkzJKBqcagd4
sUnrZu0Ieh7LbAPLdfSKsBM+yw+/RqaFdec4yVNpAFtZQ4nskUaDcgfF6fKYzVnAHGbGAKNHJWZa
txrJJIBqKn1/B7/fRgzP9+FByEOMyazbD5EcGHzTiUn9mHTsUUH6iq5re5E+YjaHrIw1lOwtmaI5
9CpDHmPSyagR7C3vdiyAS+5qt3qeNttpvysxOwSdwiOFF4bIk7Jo3D/jUGLNfJqz8Nhf9O742ODY
dK61v4I3g0PekMqpaRpqfzZIu1q91txTN3WN37Fpax+rRRcMkRMOkOkradNizehvrUurGKLAgl2q
e32uX75/o0P3AliVSce6zeBpdkiaTUOxJqjIabBUFXrXBk8zfgk3inY1UdIdemt0I2BYczb/ucgC
rCJI9MjuPWKsnOu21Yp0PpfktaLF2RVcQMu9GwvP7kfeORU9x1YOcO13xJE1sdmdwu6QcNKfYcGK
f3OrsaRtNTjKJ1eww/bJcIB7dCCRL7YvLcWR3144W8Yo/0sfEwpMA9PNn5mYuqODkDf9anWvntbH
IcSaUgKarUgd+EehsYI5+k+Ii3iQgxmx1djFwgXgjuZdIlVTEI1VW36pCVFg9RSqPOaMupOPgvJu
8+EVygxmlKHo7FmhTWwMGyIEi8P/rMZIYz9olQfDmQTfROuarKaE/S5w1wx6yq3ipZAuLnq876pY
xsEnrQCDI2ER2UvaSpJHfbqhLF6kcTN1wx5ZjDOSF6ydgY6+d1S1zDSNHkI6uJImOZNc+wY8sdrM
zBmk9PP/WIvBgYcjUyY/nC4BoZ7jInsChz3eaLt/R/LSlv1AwZaAN9d22tTU8/aOYD/X9w75RIF+
gdsQUAGyMmwU5qPMP0ddR7sFIsvgfWM6ag7abomECOhk/7OVduCAgAV1zwzy6dd+tZ8biweTphLD
Z+fcCWlwofJjBLY5r/zZE4O32biEWzDydBkUh6mKgVpQraaElgBijhOJh5xYe6NzwmjtVkrlpIqh
vRaAhd1rTTM7xGXsCaYM+e2y6Dyo7NmKliNzoNdm71qJFO5rbiCf+QW67NhznGxdydDpAycokOBR
Rascg4seGluIEMaP7J9jvBdP9yx7SxoQitj8wzFts58aQe6TRodtrEWgFBvwcyg1t4nSUf+A1g9m
0Uzs9F7sX72QQI47DLYYpR8Odjsr/top9T5sLf3vTZXHQ+3jIownL4W5Eyjzb9x8Wl5j65t9qKlU
CvLk2Qi3bTwGkBGFWsMCu5fQxzIdOQhfPfzvP6HoV9SrQNFmCM4ha/YyD85KlxvIcYzs4iXJBbg2
aHzz8qSbbaF94PGBlBL3IhsoBengqDd6ewZRkdgEb19OM3bq9rKT7OamISndXFCnVDM26WXiDEtD
wOxqxldj/24xNoARAZjpjsrX1qB1FMLWl6TaH55NN/3kcMq7LoJ73IEf7bGJaGL1SWPQpyK2g6A0
guPGtuDszxyWPBkKuxTsFzvcGbcEbqMcMgcSSx0mIpaYM3Ofwu+Y+wf3XQwrO+cS5rPOB7wXkO3B
OcI7mtN6HY6Y3T+0LEPOX934uGuG4WhGMFsTfGYi1X/toaRYXf/+ULLG3WqqFTIbEs97vyNgfTLw
KZOxNPJRyft7JZp9L7Vl9+i6Jy0TzvNkjbTQVIeF14ELqT2j/byThtvDqYH7vxvjMvgnF4Jsp3dx
NC0Vy5WHlTek3YA1UuJFJ6H7fEkSygdMmaZX0/0/y2EluN3kuZjLGLdXFCRV2TWBVdSKnyEEXGL/
N+IPx74XKBOlRJB7wJcoDXqMopvJM1WkUjkCnSh9t6/gAy6TC8c5ox1nsic2LW+BDfxhtTTFnF5p
dnvnuwp7dwvOYFVeS8WTJSa4fUmYwbIsooM6fPrOO7yzKqRTp1Ccd4+m62aRnALbNTCfuXhWllCE
aFCV8A2d1r6lOK3i9VJ57vAcjysqNi1GC4iUPqcxW3gheY3MMDmHw0bQOtlebz0gP5A9nMzd/FHl
sCad+Iuo5hpbXZEifqgNraVQZCM+2zNmUrQoGiw1PEbw+L94Od6RHPeXzrplQlyoKecl3Qkhwdy3
IUzixowBtzr4DRmJPkiDhd/ulauEZElCRqC5DhR5kOqY85enZZ1iJbTBSXmcg6DUimxcSlHOpZ2K
/4cRqw0do8QJSdvdE+CbQdYeodGOum0GOriJkTHE7BDvof4g3SSpOUvsROU0m8Wr8ZTylvF+SKYZ
LnZpCzNqBpOIV4U4fCocYYcLf2vTW7DksqPYsjylnI9DnuH+aNYMI07hhr3jCU+EUmAxllAd1d7+
VQcWektLvahuC2rJJvtk5Flp/M8apc1rbZH6ts0v/uA83PyjERmvzptwAAPKjZsVoEayoludMU+R
syYRjcH9kvbQd4G3i8eU7fly26yrH0kDmpi2+FpNl1GhWysslIw0z7CBiATTAmFrA7kwosOvWNih
betaw/JsKfSCNGlh5CJB7qV9I/kCU6p6/E/lkPxAk1SuXdFImrY8oigrGW/Ks+OWORrRTjZDx5dk
Su9jC5z7sh7C90hIs1012yskNdIuD82YgT6hOs/pFpnhWXs8f9YxO/eexQLSo8yWyTR1+VEimPox
/Nmq7yIGX8A+iz3fxs5GLWTdF69Qgzi+szu0nwvzTjqzCOu6pQlnvMMjnG7CJMqBXit38kMvVHGk
5S4crOsrLQyHZOveuFjbyoFTuJVL4Z3C7NLxcRnqF9tloumetEUzwUorYDVzkNi8MTjuSX8vbMOO
0aMIqXZhn8lXjFVuzLb4SMkyGHMSsw3RD5XgEOGQI8V2xfBIdk3GrihejXW+Qf0hbnE7AWXKlnnR
dRy/RSyI7KLIqu06liyYqkVcL7lPY70dMsutsL+GJkJ4qElZqf6vZpw5K/LiN2kVPSQO0EnJ6pIu
w3IZw0u2TpG4y9k/RvAVu0wspgvF5Y192DIzAZGF9y8k6pgOyucbtBTM8jXAK04nLnKsMRQLS8Qa
8tMDMTVOnWsz3JmIG+9oR8jDsoAfF1dS1Hx8eQFC7+lO5iSXCP0VNcPDSkyzLUubzaVV3hrWduoY
lVj67DgtIXeYwXZki05xu6uTc9eGzgMiuFJh+xqoilJ+YRzusA/UTmbKTggu4arTgCm3zDgz/AxN
M21M6p4yA/KGdqwNTqiwD1UgU+hIkZYbYGgZo2bqobm1Jf7wo+ZR9gQhu/qbDYp54NGeo4lxUL7+
mwEpQwwCTVOqgupx9oY1aw2X9++e2pYJ12VFyxO02ZkP3CAE1r/xFIxjuq/94sT+8UwCyXv0GlGm
z+RM4V1sAi4cU3paxI26Q34DsxzMS8DMTVFCZpmR9QGID/afr8Yevd48OWmTcaErhC6TCuCJGZx2
jkSn0X8qAeD3ZXm6eiBtXeFNzbyfPjS1LSaZ5ttnUB646NXh86R3fbysUm5PfYsVg83hVuCxwYPm
ImUyFivZHO+y2qJBPL92kZX/sjh942jqtWYzJ8KwLCl4CllT3Z04fVnlKK4prk5Plu+AzVIoFaW5
u/x1KHp8TFrvRWH8qTW6XGDrGMf2udF4CN84OAIlfj54tI9XfdPdE82DWCmwXzlqEnrrTj2Q9dhl
K11Uly0CngXbnxqsMe2kbQbg1mdueXGUrt9wK49+UrNHRoUb+O83kWoTCR9TQiqB6QAyTMzrwVDa
FflwqaTZqB3xLNWdMnKlDQelu5lZi99GGfppSHgBV2kAS2PwybaMq4ODhspikwfUWCuHwaDCPUfI
oDKiuuhgb8CrQ5yn1CpNsiYCW/CaOiBLBjtFuOEiOmSoXhP53Pjp6z5l2KGKfQxT1epr8vFhv8Du
q4e15jRTgJUGKMMlzOsrnnSPqrGkenZKO9jFqv8A25zHhVMMSDBijYlraWTCTM7ZwMvLbnzBp4GV
NNOhH01J74xXsMis2ejBHA8kTdfxbKrUTH0dmQvfygbnVn/rxo5/nvb+vxtz4yPEI6sRQ+ev8jzr
rq6vcAOvdvqqH0s4LzioDSMwT7z0Y+We2uBd1piTatXyU9bOxD/2ReVdyhbZDbWyc3u05BhgQ06c
v5O6sTJf/zFKo5DFwtd5yG/icKhz9SwDmih25m1uEz1w1EsRDu+mVSU02cdH3MU1jNkPbMQ9qzz9
jnDlSHfefnoZXX8LzxYV3Y8P/XtC1XnIQsoxCpcOEApAMZv+JmLr/AE+u4p4R8tdX6zSuQ3ZSTCs
BWe2Ci5fsDHEns6cZsWDM7feQZUfOwQc8CXmnS7fEM4xPwU9LNv3hVc2Y7Ou570kK5/lO2kaYYt1
2hrcBlpQVSL/ut2yEQ6AXOJVctBMPOpw8hptaMdLVU2EvGLnoNd8Y8ZRVmgT6hm9Sx9vd4i0CQgd
77T2pEVuIqzvw6r5XzpCqIyBLNibm7h6aeQvJdxWkhgOjWGD41jKB+Vy2zOv7u3gr+5IYH35ATkR
sWsuuHNw4U/wv7hgvBRF6xb3WIjwPRhdvYPuoElhujRqOOsl4EVK1w+jy2gFNxe50Gc1I4O0yZsG
AWalVJvtO5hjdwD0lkt6KeU9TJEtHKsL6RyJjYFQKnnTgpivZCluGW4cmRkqxAe4LFBOQR4ND8e5
7rmKnR3m3RwR2gcTUYfI6DzyqMW9k56epEBAVlfuxfBMhTSG3JBX9FmFG6kwPsoVFhOCGD8AdHW8
HIaigdRfa6mKLTCJV2GW3NPToHVyJ8Jye1gYbCJ9WnuKwd9auzz2Db+hIXB+VL7lXKoK1qcZPGGC
EnuN2zEoyt9ZmoMUb5bovPOwtqPjTUNjtwwXFU6rvvgKVdR9rm8FT6LNBRojg2QyyyJ/l3tLa+hU
Dutv27DeKNwPYVcM/ubWiJfLT9b0N9WWOTG7Z/z+l21SC3W3TMUTeB6T86UP5Ab1wHT1DYDIbQnP
HjWTU/7v9ITV+NFtBfSSclnxMdvR5LGaooVgVV0WysOEza8/9Mfh0BlxvaXyAjFyihI9IyggLxOs
CzXrV1BjKmS2ztt6SrzV4pGsBcXiJiJFR8da/26YwBRLxMj7jrwBdJbTF+2dkUZVxew5XgLp6+RP
FJ0yCskZowelUB30fY5NhqAYW90mRxNIyC1EKaqpfkGY/6QP2/K6bqZ4wZO0x/GwPxWpAvQapdFa
1tXu3oWriCacub/bOBdYREb6JKghGe9Hr0sDvgmjoZ83aa+DbEkWIOKcHd7vl/4Jc3rgTq5Zx1WH
M4T4j0lbYrKHKkzZ0sAUaRlf9E+dA1CGY6z4mebZ/LS/P+5ozhAtSsWqBmpFvqYU8wK+lM7b+i2/
OfwnjxY6O8TrgKiiHfJHSqmw7GfgEPNkOUhHB8auLeDXuaRexitNW8B6PezKQItmUbdl6vBa1lE8
hXeoFQpgCswdc/HHAgyjZpAGfl2j3LjCdSlP9bQkb5XZeRkAX4JEjO3zOFg/Qj5O6Trs3pbNAKC0
Rb3z+B3m4jiiDzMqVgMjMzdZMOVWq9VQRj4OWtqpfcV6fPQmJHgeZy2wKyzhnZ17xL11avc0/sUg
WwXVVWnIFBkKy0C6cMctE/Cmhau2mGYNQAEwQKMvHT1cAKUepJ+4KVXH/gDkd0IrPt0mtfMWeC5I
4fZOizvprTAmoKHYXUiW4wysHUhugAJWNgplKmz54mRmR5bli8r0mg7mc0ADZTz21aLwHw8G79pL
GSw6z9KJXU80rZvjprA7zYRt+NmBaZQlV25rags4tzA8zjzlfjfiFu98JXcK7J5y887YH6uxR6bD
s8WtcEUqXpjDZwwBSpyfoCDTgDw+JTzljsBYCy9gYQmVz1P/g0Z71BUa39QovW1vu8vQI4/qIQUm
ot6xEVIdk0xHXklSjRnKSU/PqjPqEJUr7LHinX2C5u+0lcCOS1xt8b3fG1Ew7Osuy0AfwP3Q5CDp
kOegTpfvbgEMLyMi0gU3cbyK7mTySWm2OEtJ+eZZqFgvAXlokUoaUIF/0pfb5PjGlst6T0ozU9qM
Ez7sE/UqYuhiMqm9y4JZ3A9W1Gafas9xu7k9n4SP8PaiLUvtpOdyu7qmqUWiJy0QdYUDlvHqkDLN
K/ggzSCbOLTzrOWMKaOQvLw55BYd8djM2FdTRCYXSdIhqF7so/Iddr5nyr0wBdoZaWKNil0mMBJc
/PoP9zblv5g+OHRKH/R6gmi865+8YE8GysfyEgHUy/jQo4pZQfCLPbpEBLBXjRZlBUM0ncxHqtGa
3wtLFVvQmPCoeDPVs32gA6mMMQwz1QySvjoOvY6UGuqeIw2P/3SEkGpg51TBDEAHBFG+8udzwc6X
yXHiaX+3JRHhJxiA0x2P0xaStZtk15lTIec3OOmWYhxHwh3cYYQrF7cSamCWf5na0UVQ6dwl12Of
H5SvkyMm4USYoa/7Vu1WDpv4k0vI8wPfRCe7hZKKuVMSR+KNQz2HxS0T9r5clUPVCBzWCEQJt0NB
XPCmrCJJbWNO0gC6S91wrhatRtnhT6fpRYZdCcdIC1fQTB0Wv/WggHgrh4M/ZtwqTQYqKJYr58Ox
9kXZssRGkRwCREeZjJF3usBzDZHBAHYXICOL3ZOPAcdLUs6HpdUj7OcIuv5fcvtYIVlc2FZBOEM6
BhsruZhMpm2g2gS0a4VW0TQMVAE17LytYpoScCxcT1sT8RNexXv8MlAVcInC/V+O4xi+xr9koj/B
WdSrfIgE5B8OXR3Eb0eiQc2lUHm5CKDvYuwWTTn+AU9D7EgOpKmsOfwh34iUComEcAJuuhT4hCCr
76sWXTgGaAnt1kwOR8vIWbKrbHv5+vFGbKCVMpZSHKeL9Yl7MxDiD1Gym8kh/vmtqoMVRS/pGlbd
DEj4hgl4
`protect end_protected

