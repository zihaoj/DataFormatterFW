

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KZGjAkLdR3kjLPFPH5iJsGRlx2kJ1RyIMt1tF54z08GdHl51la8ekAgXNqSwHm+pUkSxA4BlSLmJ
gvATujadYg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d7SQ8S104tvG77MP9xZ5+VVHUHX7CaOet7TW2Un6VEQKY30cW30EjDTT2OwPHtWSUDpAt7nyivp1
OifRs0kvgifi8izEVbFRuH/kLIEERalcg84H9yQjz+LVmXiuNUBXk9WZf6vFOBAlXAqmVrTG7VX8
IAua0vEHboqPPMEQJoI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sjkpOc5VZ+XmiYF7KtnnIPxnAhbs6+YIgOV3JBfy2/xXZFZiYr0fz8XXQp3MyjkLdXaiMdsN6UoJ
am3mV2qEoZ2ZDtHbU+SLmvSfrFInhb6PBtcHRPZ6CupghoMmTxbkSUsuaT+nCTASqLh5Pqpme+SA
pCk9+evw7/lHFdkSm+dvkeRbcUYvE74gGmjCSZHWU6Ec5bvrAPc/vvFVJtm6BdpKDgt0pX2r5B7C
00qY2RGtNvbLonEXOjfiHxAASF6STcROY7vI7TEQ2qZfcX4PDxk07r9p64R4EkVi81lqhKq04Ljy
aYTOutWxrHDC7vKTYQMYuxHa//0LTnlEgLkqnQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P0FGyCrlRNvkP/m5GQKXkrfT82yUReudoEnhYNDV6lUCpPGIfBe0kKt0N0evKaD0Vvk4+wE3IGFm
QvNXrBT+D/DaZkGuiz3vGeN2eskrvVl/NJSVDbCORE11zd5mTl2Cm9swVlTFxaboTqvwXJCpWbrI
5T2sOUizFjjMgUhW2U4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sbxBNj506Htq+9fXIwt8TwsCd7XbwXN6TWfkgpmPiyijyl8QEerDIG3Mjyb5MfQJccsqpgChc0Mj
2LezUGzRKAbgGZZfshGjCIb9KYhGhorzzT4W5OJexGdeM8npWA/aFeuIsvPnBlJqY11DgzzG+wMC
UWHHhyLa/yBrUMp6LW/Ko5nHSbyB3LcVCuB+/os8PZvJDZ9E/DIcBV6I/9RMwPmY7UlPUf5uHkNT
hg61kQH1igmywF2R/gKaA+NkWjQ2aq3+5Wwxu9sTfNKETbeSrKCQENhhTvip6mJ02jyiAbtEqIoY
pCOMfAUCHoZZnuORmhpRGjp29+ccnmJbzapEYA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8336)
`protect data_block
qaCg6nZOckYckfJh6/dzcovq1xaC3eHGocCB9v5F701ixxKiHx4C3cargoE1SVZRjHUwqF7ffD5j
1duUojxTWHmxI2KrbE9ICls6uWjAd8KfHn3MHP8owuomnhR3Alo2P9cS5NpF+3GoFAAtGcrMpV9P
CEDWhmysjCKYal5VtHOM/LQi/1fyOpN+7XvA9Yyz9WN3MxoBgaZWFUaRjlZN+6VBwT05GhqcG7XV
9e6jbhpgcaBsqu9cShmlTqswS3Ckm0GKCsyWasbji/ZTPBKBx+MAcrMzOOKmqztEMmcukZPLFzGy
LHL8L5wC2Vt1nr0yN9hnClfoeT19o3obRoomkw0vpNk2xTfOqSJrvPfarp2dHv+JkWYWejJis+5s
OE9dHhbOfx5J19E2jn8JZUqWd1n+A2aSvdXOE28yn8KSoqgA3BRtWvvIrrzLwKXZu+c7DahAsUnp
BgHbvip8CzT7nd0qGdQ8Sf6LysHJOHyeFympuOm5IPhrcBtuokzQDuYVpAxox1PxntpW2JGEB3Vd
H9Bq/TWvQgvfpMmtbHGrWj8BgoOngFU0AQWEgLum28+otY4Zqxfl5LGjMiMUlgmd6VAG1B7u39DP
M9JLt1nV7x59OoqkMO72L9voSxA2EBOJBwCgbjpavGD9D9i2lCBn8JjaphMKc7gCsVkFUh0ave+j
Vh4pPSAGaZVavamcF/IqkZNRihQ00jowjMg0sn4Ji7NnzW/IsmwJM1OQLfKrNd8E/EoAzLAWPtdd
JE/eHck+xwQLkQGQiVM3tbMqaZ5urHSM5qeZl2WIX2d+C+QpFLK3C5/Phi9GVvqNUtjZ7mR7pKAb
0UMhIxGN5GZQLJdb+iy+24OMqQEDRMXRXQ7qu/UhozG2059jdx226WuxusPw1DBGiqXTHHpFeEPv
CO7/e1pOpNl+Xy6Mt3pRbkBoEmk7jDhdNa3PII/+Zfmn5gXuN8xzqmSjD/c/gj4O0jNU8sEFMK2o
Y8fklLCEQIRnCZnrLsxY0t8KCmhgxOklO1zQm45r8eobhlgGfF91jIST9OYZbor76n56sA9uARnE
YzFlTKcQE0jLGEiwCmJJ01vxcgVKYG+iOZsbeaHyNK1GC3HbexuSQdGyL/dRhVki8301nXNg2wjp
VT9/WUpxR65NoIMBG/WvLROrxe9s7P+8Nh3DhOdCtkF2WmKbuuZcvyd6l8DwQHTHOtI/QTY0M3Fs
yIesXTHnmmzXyUE+bnPqT+xxIwRnMte0P758Q85bxeBaYXylL74B7EzLJQxGcpn7Lw8HQ6eZ53la
XN31vMjD4krgm/FgulFmVNOE36gyIhFgSJEzkrze19udW5lKgGBKs9IGdT3lpS0EHoHBaiH945NT
aaiA/EH0iceRGMfw5HqGLpCpBGl29rLrlks2GIaihykZVw1RJzHDFFPvjlzxyjdrNoACU5KzgLwe
lcENzIISKjUB12jUfOjWd0oy51jphjTNMaSX6B2Z3GJ7aX6VAzqjqWnUh+KAIFkBaOhvZlUvT7rj
B2uwSwFAll27iN06nyxJu2Al3u3fio5Op8sbqvBXD2Uhkb+69rJfhFH6nP+694qXwqHguqOJWYhk
FPAq8YzqFsxpVGv0rjDzhWW/lRV35GuHr/uAB5XaZjp0S8hjy053vNTt5y6g2vKaq9yKzqrcfgoX
3UCIbxpJ7unA/JRfZl5TKVj35RwVesj8g0AZTeHftH7gAr1nX30O0hkMqXUU8i/LsUpOhXdjtW6B
PNOtNoyiD5OuQHsev5MbmE4yv4atBtylXa67SF6SFJkaS7MsOqHgjjqiv02GbhKSOOK2ibBvFdbJ
2UjlBUEuEDESTNX3XGoFojZQi95q2wbxctfC/MVgA5C6P5X2Qkmhv7C1mG1t0SwBs38/XAiVBc+V
Yn/1YdJZIGpD2PH+X2Qpt+9zPUmI1eTS1NjhVkDqNC0A6YLZBoVDmENQaHVLTlglf9Fg64VGmLrT
sTiB2o60BUT0rsSDtNTC4Y1lLzK2mwnwzmWo+/CZQeWIHFdXy8HCP4vcgS5QulPxobllse7g99xs
jYL7gL+PSlUKjzNvblniwO172uRlbGrwhXUH/B2IEnULIlVUd3FJS4yA1UOBn3oHG7H0hj0mIj9C
eq4/owrLB+O6zK+tzL4DUnyJaiRTLlwgzatk3hAijc+esP5+xJoBcXdxucNeDHfDMBTJoxmYpNRe
VB548Y3BPbUCgR0b6qCFQEdLy2pQ9w+JkSfbUwGH03PwXRmOF3ZUNGyEpyvbTncLx0MQ2LxbvSKj
6E1iYn+FFbeFhFoqmPBZpPKUefokI2o6UhWdxQnVb1U7VMkiJATvvXOU/BorXWyLl9nPqZUk7FL4
OYIh00ZsYgUO2LxJ0Ec4/t7HUhHrSoGKqtYzYKiQp2J04wXM+JReu7q+gkwjU5Lw6/Sl8lWD7KEk
41t9qF9bw0V7ENMzJYZhNM47lujQlxsn88gdIC92mBRC76fRX+64NmOWmHvweMEsvDFUFqL8X8xD
VjquYhv67W/fNxwhNb9VctsDO0hRFeaOqyAmQ5Mg+p139iu8Lt3Pwtm7oLuiIV15khkq9VEDmLbG
MGR9ZiMIo53bTaDobB+OBSWjlEsG0ZgqDmesgPzPNqe5U/dEdwbmqGcMaen0lOjAuBS6nZanA+05
JKgiMKbuhQTuNYJPzstAo5qaAyXpFpKl0XpmL/ky0rLFtsiRi1KmvP3Qr02h6CuFtvFHGHch3Yn/
cH2iFNKndABIDJC7K27gcMLHs/ztY/hp8JmPCYVAYdQaHW6+09ytqLYJwPxk0u9YsJ96zcfBJ2Ml
e3TXe8YyMRohfc03pij+zg0WlIdC0UNJb5xKCMleEsT830lTJQK4JeT/AG9qcCDkq/rnPuJe1xzc
rdcOFkIMxafTOCEYEQh/po53nz1QHjOFxBzDwJ/oNYILSXPDQ+5XVVIeIXb7/1vROGckU50H4eZR
UiufKyk/mIADudhr+c9QdG+6mQWifTkeMiIMdcSVtBbzp5raE1/9qkODMrDKhvolC8uvU0FzNhXl
2iV0WJSIAuxRuub1bShzy7I2SlQYaMogmHRgMRhTMUcwIzg+U/Wmo3sCDaDi6/aKyXsvWIHM+0C8
syG9Mc/XXP3HR+Zrwy8tW2jjp5VjU3e6nma9FEj9juPpcqrHDd3cOc3QcOSi5iunS4kwXez3DMIT
enOvKgtByCILtuXFVzL8fPprhNc4cw+pmX4QUctQ4Mkn2jyBKlsgWs7unEt1+y5LKCXP+dL8Ms4W
X3qxGLNaxnHuowkCT75cIO/yZmBE2mE6x8Y8ZbDthPuR9HPjTPqtbXK5luXCRxwuSFIvy8VtagBu
+v7FcRbi2oQxSCXRr2qBNUsftUssgb3ChK1sNNYbj2F84eh3KG8eJmIgIcST4S1oMH4NecTXRN67
LYNCGyS8zNGzfpHAqIe5033s3LY/6FGAGtL4rV5D/8t/yRl2tuTYqXfmizXsjacju/rDWj8vToFR
zcCqsYsXBCh71zOvudvbQ5dRX2btR1LciLKaae1/87cufVfA6AGbRyAw3cR457hLfM6Kva5gKsAX
Cqt7Cr8hgpOwwEQeY7VNjoEJBRzO68r/nreoSyKwTrEtdj+kkKsM0137WGW7C4Hn2l1rVmxr8FyT
nvE2/MFIe7gMlo0+ej0caaYkiS+0bsRQB7l9XXzdJd3PPjf2u8PzpBICGExfnlKxMjk9/fe3Zs5f
9w5+at4YF/ESSelmOt5WccTJ9+2Hb6Fwu9KfGh2PCbo24ZySXkhh3EIrVZ+zS4CLL8x+pyfkMXh5
dk0BbGmsKY7nXEtYgZ8vcXPfYmCjOABhAchsH6kspE5NuVcER0Xr3SrNTnhrUZPK2TOJ/hTYtsfi
pwvn5teHg89dlCaaB7J6dH8P5Sx79AjhAPNpz027o+LjZ1b3hgc8togDaFyj+l7kOlwCPASP2MCs
7XRw0z0W0te22D8EWgoguHE+5c8wOe5dTcacLBzeusRYUfJJlCA5qRpRgxyCYbXosW5mWj5yqDWD
3ddBQgPtVIZl4wNJt466X4kHR4e1GGbyWNsTe1JPlnd2OtghRHRs9zZje2tjoVzLpFXrFO/anofs
e5DRj1sIBCyECmR93VqfQJIXU3cgTqwDeKjN+PHpA3sFDruGFapaIiUEvOy0cHsDWBaA4naOYB52
nlPGGN3Z48ZaGCzbsZw+msjhOcL7J4JrVvrmSrnygwXE2NhJSSeDxWj4aUHx8KXdO6uYVo5iD2as
khFI0BVrl3pOfIz4vi50RLMImPA/q+gW3mGhPAmpLuEjeJhCDr5+xBlDBMw6A8tr8xR8AABdNzqn
IFKuNVrAPWjfjcR2wO4UuifjvS3EKLleYbhA94KOab3mlbADOfO2F/TelbMF36gBw3/EpiZThpYV
GSsOYca2vyDqLgGeceQN3vtJegZ58LlozSSr1uB3bw92FBUdrSOFKwbHunv72qxHwLWhLV0jT2XT
pX2D1AOG2hmkpi4RChT3PZmu+NipDn7zypYSBMfjFu/KbvMzxJ7ZKwnvBnugfYkiod4ron5T64YQ
yGlvKmWXM5Sp3fg2QRk0S3uge9TsDyJenv7qX+zsA7tcEP+6GvVUApIropIamjduAeEoE/RUKuAV
WkJuRw267ZhRLUZhakgotafR2PvWLQuhBcC+Q3zWDq3i9sHztpPJ0MZr+RrqyeJjJGmMZcxXX0VR
odlYfInsl7eXwj3GiIu7m/GJgeBlAbNvEnw2xZ5UWMvOEYUvcsXpQKz/5/r82LmXIkXWa6576+WP
RMwXyhp7LYGxdXOcEmVXsq3Zo4ylPHgtC6WyELKtQsReogoQnzVdoPR//wlmsAGdmDj7zE7jE6gC
3InfOd1WBDbiG36vl7pUbOcB6wKGr9UKuG2IVvFICtyXErwLVtAimUSP530/srMqhCKR8ej8NCkj
sOaFYIjMpZFh38ERsehiZGRjZ5I7hgq3sVI1QvbFNjFUgY1u27cQrbh/Mv+aT5AollbC8vP7fEc6
0mNCdGkEgq92E/xXlXbJ1tZ/kCf4E42SZXrdCLOp42pUtx5vjFifUJFYCX1C/0stSKi+0pxsgyF3
TzgRmFiEXDqQ/CKVq7nKr6plQi3ukVpcWpz/XC63QnX15UYS8DkadVi0YnI2Pe552xNxhGU74xEc
oHUCHMO/zgYzM0vZdJsXWKm8aw567NXrHhYD8D0FpQg1Z+kXjxZkz7xFIDWlwl37wsBz3XYGNulh
rUjFFhl5zphkEcaKPhVzAbEPefOumFqMRLiTlbzFMeYlYZ+k9vyswKKUByEhjxik4rgcUGzpAMxM
kadMjdCAsrhAHs7qS0h6tKTyoiizSfnMNrGGyeBAZThkXZlL3nCElljTU/qYnd0kYwZ8/DGHLmBv
LlgtxB60m8eVY/g8m/qoySG784lmVOLU7GR3Fr2AogxKKrYMSSNyuC6WKM20+q0Xo6DZl92+uFZQ
YrfcWDABZzruxhDOKp8hzBYtsdjwXTYU1zVxvsqLGKi0qH9ELl1ev5O8F3aH+Ak9frXxlGMRq5O1
SBnS9F1ngBlWp8ecD4zc9oDpnOuqUKAQiXv4k5LcaIPzOOX3DaJM4+LO3wOI/tPJL6ln7gG7FWf2
3NX3SrvMRJJfmPTAscgRni+uX4FcqvXiN4JOoUAxEYipvrJefKMXhhgnPQvnhc7AvQIw3QFKD77s
4+snVIsoPvh57lON7XIE+nsi5DPb0PoXZBKwa2lIM/LU2i71tYfC/hz8W0zTnLlH+HO9idgvboY2
V+HP4NAVIqwb2U3jtBYTbssOySPbJMPUIG9wEyvxCN4JM0O2oSl/e7ipGTp0g7iSspZZMMpKyAnZ
hOyx8RmR8Ry5z5VXf4Y2lNZi3jDbKZWNOvPDI+a6tAhWyfh3joDjPlyWVzu+PrGJ/1dXX/DT86tk
KYwoxlFzxhSmbnF2V9U+X8zGx6fXd93tD6QfHW1Dv200z+Fz2D79X9fzOcOE+jGCUoFBvQc64ptj
QiBor0JIQS91oiEDIRexXQBmJhCTqKhAf9pOyXzg6sR4ycn0qtNVo3ApQAdCv8GI4TwDhtQrUSpV
HXji7Z5NXfXAk9366bMrqAjLDoiG1D0W/5DfuZb4mDAOyq+7OucLVn4AWN2BvERzyV1a4nd9cMP5
mQ6Qx5P7+BDAw51Ou1fT8uYgnwx6owFOZzsvTN+RxkQPx6KH0rTu3Fnos0eZu2mG4d8chojw7eeS
FEqWK3I78xPj/1WTKDKo8yLYdUQS+f57YLykKmjwJ7zjA1c2pViZSDVP54ij97BVHxiEiIzNOJ2J
qk0Or8c/SnRVySy7L6MjpsUEj8tnPW9CDgGTfQM5w8KPvpY2HGTkNQgC8B1gR9mi64xDdLGFCcsH
AoCNKndmqgG16XNsKNXcDzekbwVmczMMDGEo6//2sTmAEnGQ2V1WguwKfwPsqXmzLe/7h8opFAFw
QdBGHatyVHNmmpL37tayur63xWscYkqtMoTE92nkg/LlhBg/ZMG7x4IXQUzIhLbFt7UuIbJFkNG/
siT2/3UcbkknYo9g/VKldpVwBSSb1bu+uvSbls7yS/t95HqVO/NP4EjRK/FVS4wI4IhDuJZkm3Vj
V2UBbYuv4wQ+KlbBvTZ9fhLxJ5VT79NCjdq111+nAOMXYpt51t8kAV4JyoqzuuWNvtUkZirXsngp
I+KG2IMwEv9mLnZQddbJctJzo+5/C1XXIcIC05It9u3MFRs7WNeJdT6LvN5UVhggxz8AeXrBf1Ia
wCyqfyUxYsKcwQPS/b8ot7i0Uj+1LYhoSwi+xh4SuHwm/T1NCwlc6yuvuLbVlWu2CgCMDDUwZyI7
WFKW4u5r7N3zMK1gGgWO3CAvYdbLEpt2NRERDGeu5Rrhbe1JXqFYS/MSYqrRwDdJZO9QskpjmjxB
ANNUXNhwSgpKAgnt3TDDeth0yjhQQpUFZ0IAGYxJtYrCu8a7t/zqF2WLsMpUpbK/Mk/c1FL9SCNc
OkQOqWKMQc0OLmS1+a8mZLW7XPHEbyk4Kdga86XTpYhyo58vKGhWopXSzDVMuopg6Y18dGyIABUK
kj8mR9/0SqXVMNc6YV3xXF8tqFZE7xONvKmYVwiNnBoGcBramptIFlDCMfLTRtHrjNxGi2wiQZLS
/DrmryEzKUm4NRLi8EjLZ0oNvKnSbJmpLoGZkYF9uRjdOzXYa5eSrCO7jEGkkA5FmD9+lrssM4vw
3x4F13c9HxbbwnJhSDeDsITZvwEz/bW+ZdZGbNuTpM32bOJew6qcvBy28Zb5YAFNnbDvkVYOzgwx
LT/ucXkLbc/Ph4fGneKsBJHxTJLEOc+AaTvGZSofNj0noRBCS5Ni3/LSgXyQPeEHcu8I1Ic+AlgH
X/dbn0rZqKkE9PpUlgHpTaMG2KU+Yn/dl0KA1Sw7DepXc4c7kq93K2EhvJqY//XHJZIdVEMpTYL8
hZhd630tk+hopjxr57TmTCOFyuvKyx2UBFd+ag6gDvgEmvphCXgM/sIuiG7Bd4wczuXqsW95/6zC
kDNVgjhICM/FDrFqZswYrAXm378oc+c+nxTMG60qcHtIZ4j/4cnhNbNRRvkNOB1u2h6ywlAhtpcu
H8YMbcarXJuoAjKFohTjHN6BCgFr2wyOKtlcWEYiIJy7m5s1/p+yz6XY0GWqNOIiQFto5nVf3MBk
aqryfkxHvvlazNG6t9f0DtBjo3AhKCzHUACVzSfyCZYu4mouBTKB6AORpa29eADmoI8KOQIVbeYz
WQLUORPKBgA3VB4qV/zzAFwQSAmlfOm70JyPMr2tpNBvPiUEDwyD627T37D2pqLbILGADOwLbrEq
fT2FrluAuTcVWsjtdI7G2eYadgf8EbzwZmmd9KUGKmUUNOu9M75X/ojc7Agp4vg7/r9n7TxYl0Dc
rByJPnS1Pbx3ukXl/2Rg7SxnTwNZeejmCuy8tprMJDf1aGF4qV31foifSB1KcjTOH/8mEwOGNZum
uPRW9kQPNOjEjhay7R4ow0FmMbtJYwUw47z10crP+BsV/mZLk/Mc6IFACC1B9uD767abD3Aua1IZ
+ezv/uctRWyYnSle4Y7lcVrUFggGerK40+vFN8u4BUwwWu3nUDpE5qs/Cwlfhkpu4bG3bUSqS8de
csc3dOs8ZxRQG4JKFJvJOIYv9D7lrjazEyvyv1StXHMh7f6ya0+cwJBRkw3H3j1G3fyjhR7kyN7X
Qd8ZFK5B6jMw0q528eRsvf+Ix713th0h+gf092DJaXOsBOONLDzmCbDkL5lMz2qz5O7VCiY41/Xl
hcfMj454mIPPj3rVDAl3mSqnRM7sM4HjDlf+cIW605Ns7y4Uh9pdmnOMozCBK0rkQBQllvcaR1sY
FYlL3B+lVuhWxzh33ojfEMYYqLWsUVJMdtnvzvW99c6Q8PDnyFQLOkxYObTKV8/gyTuIUtDI3yvc
yhzc18UmlcaOZlEvKA8Lnx5GWAXBb98aOw/QjKuovXntNcWTljGsq2UyOIzBjvR2wS7kQzSxGonD
v+6R+WCvBBnUJ/89S6Ipt9ABS62xK8JfR7nR/D2xpSWlkUv/DAey/1vEJfdupicO/QlTcD6A+7r6
akQstLNoVqXOuYnR2RWsv2FTBgvKBlX2MMcih9yb829EA3TbC80Oo4ByxKEFkkmmwE8t/zJSbUoh
4b2P96gwST9zGOLImMNJVRQwAlVqjenYXyW7jKIUAxiCo2pjY+eIZyvI2lsC3yJlTELlWbjKJdZs
BN7e7wfAx4J2Ff8ChL1BzNalHT54gfbS186jkugl2hxyVTOXaabg2woLfwjMBqAX7FmWT7y8sk2P
rVkwGh1odacEHSHVnf2dzvPpX6ftdAZxKFZlAreO0af1e+SiZIQgP6xIgLYrwTmuSAMsNmOYSCxa
dlzvEZyBXoYYZuLSlA/dU57UfUNzaRa/cO1B5jH9pTsgXHhksGg0Nlasdj+ajpAjWJTtYrQvLILA
a1WNMGaJiYTGnqm+c3WALoShBO8n7o+SMzKDK74osToegpPfeS3QBUjVsq/uYHYiyH8aOupAMtbK
kGa+HB2Y/uxvWqXOnnTBvGSqBH7ek2cpUQ96RJ62bUY57jXv6vcbEt8KFLhDoR1gB2iWoUD9/tuw
CAzG2UOxqP52c1RFDNqoHbKBm3zvpvt9N4mfKQQCtQCuDDzEPL1OPyHgqSgTeI+gJ2FTlKuHXs1F
C5QMnVjB5R6kmBz0y5pStNEYT5Xwp2IhAsjf3OCdrSqWLuqtoudSYdfdug13Y+8G4deqc5CxGZBp
LYUcIcmK12DGtwTJcSCDYVPtt1S4Y0nYpsJTDp6269MWsPAwyGLaj27udc7vMr1aWXK4QD+bWk4C
J6TEA1PlfOdwbRdUSedq3JZ8aEPPqMIgBbimTLQHXHwPJU/hN3QOx8aQbfMD1ZrPqLNHGZSMxSER
x8Qa4OL913Nt3wUE9jPMGOcCP1A5YAPOPMm9I42seNTVHMuDaid0iOwXfsy9QZIYCfGMX3lDwU4F
yFTs8ycgSI4YlOc0o92mgzMxS/iMg79l5xAnAnn8a4VKD19E+1JsW3zobcXeliiztZjoCnU+BV7N
ww/nlNphhcThJqOnrZ/xVNJZp+SoeFT+qBhCj1FNr5JI8TPFiYysgsuqXUl9eEKAvy64OwuwOD0e
rqOV3DMDbaK++vs/4MvoOytDtNr04rhVmTYlTg3d8q0VVaOrjp1wlEKFSntm8ZH/fUv5f/Yj0PRO
nZz81B/C6oE9OYsAgSLSd+45WVJBmoQ0moES55uWx+G/ZMJTAEJyu7nNI1jF357D2yy5VLm21htt
N4lBWFcpS6f5vG8s8rP6qrJDZBfJu+lqpjd3nD+FqP8lWG2GNczaJARmy5FSWPV5+Z/mZSRGJcwp
xP+YqpbQW1eIYBtmQf4fUzmixnd85OdFcS5VAAlJX15OZtLG7cJbSSLDNvs9DCVC3tQYCdmrwlMl
s+/1rp9l1MIT+u2HINvG5AxranwuEk8WAr3BNEvyTGngduZzXAtkvx9XQ1f81tcwUGqgo8fUNr2V
h/2A1ZvzmAiCqip8z7F/osQuXK4uJQmLEXVYTgeZHNJ+6EchJ0Nls8IMUy/jpBX3F8nuS0dtij7B
LiOWuesQErSkfY+J+lbBUKUPamIpoZRSfeApTrDyh+7hC5Gz/wIjxyPpWG5+romyox1Ejhfu9I7x
M/oE6Y9LyadNIw6gCAZezfWVOjBiZyC5hmrpZ/houDWeLeTNrGAe65bDGazJb8GrEMO8hRUJ3cdi
hW9HPXggWq1FTJ7Ba5PKLXiLs6UoohNJ9LHD1d1QjnjYqkfrBsahUrFNxjVvi7DF2vugyo/0qrZB
kRKvKFOoDe5etzhkOH4UGOj6UPgdmU8Gmchn1pqJmnwdStRDnZJB9hyeMoALtbb0uGeTF0lKlPvU
j32tfa8IlMpdYnQRbGbyjNpeVoi1gSNd7kifOWD3Go33YPD1+bNimtGBkonII+FpP9uk5lh5YxOx
TiH17WxITr8BdioI/SPfFmMIz+M0X1CYqlH/f8heXarzwvJrv+OTelpnmOBhNFRPPIXKewfZxJ49
rclM4+1RUzBA9HPqmERVQ6cMPsG1t5zZHS1fD/z2it19wyjzEltDHDDCvcb0jRZBG0UHG00VFIuD
1V4QXXlRFjz63rjIxdcHrzDd85v9i8irRxphjaDTwBXI4c24d2+TLBZLTvB2J6UkBVSzkuXs3sFQ
JaGai54akQs4XFv2m6BMJ3m6pjsFELfR9aGz5LSyZaNBR2L70KzUzu2ky0NUxpc2Wy5fkEwNMIGn
0ar937KQy666di34vtQw72naRlc6fUuLQ47cNL4+dGornKeWc1U/4FGe4MaQo55dTZdbE4pwOWKH
xZYWqKP83X6GZIMJvV0QWTh9wsxwi/il1FFc5IUN5HhxRTmaH/w86dvHx3JaC7/q0k8nRMM14nBi
a/HiM7G/jYk7L+RTlx8i5w1YZWuvY4IhpXIEuzdg8p8FT7aWKlduOZXe2dL0oYtxcFOlclmcLr1I
BMSNmkQ5RZ4BuhgcGPU5Rm4AlCurhPx6QHi/wVdmUhdwauFdT8XCfeb2HP1IJwm4uyrJn0LS71aD
vwYVpRVvN4Wvqwm8h2w=
`protect end_protected

