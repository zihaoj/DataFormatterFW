

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YGdnhnEQiyXmCAlhMhs5C9Y7Cy+lJXMLhNBBLSL0lPedQLaoe5dY3XCmomiLTus8Yqm/GYyAKW/G
VVpuQ0g3pQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aN+uUud/I007VUdNLHNi67mI15MAqYjkbrMr31P+z7klbQxWm9CVsMmo2yARdmDsjdC+QWvmMBrl
BM/93uPjF8gm1iLWvV/lZ1tfnuNAqGZQzQcdW05X+NGrNanjc9YcRW23UdvAMv2cSpF6svSnjabd
hI9m6KXso5UHqU6y+Bc=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Sc5W1zZat0W63GLsIxrACXjAgjXjyl04OXcHwLJWk4iv/NLvz5CGFX2isK0NuFQ22VGPtQcHmGX0
sqQEMP2aZwNeTddY+nArw/jfebUXsinbuXKW0SH/EyI+VCxIqHP12yaT0OU9BzcZKA5wwd71fNGD
cKa0yemKRRS9X0xRRcBOYQ0sgCNHb3FQeVOyrh+EFdTfNiGsKQ8tB3BNCq35lTg/KRpFdLJGtRJX
3tMkRqkPSv4S/ird74Ts+yX+xCFDRQzTTdpjy7dUDx9oXZp77zTz9L4YCXDWBTsSkKKWb6J5vnii
D8ZdtAV+bgNhP5COAVMk8GIB6YQDmxV4ZONf+A==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yLoFT4288OmwXa2k3OOHBwJzpLpqXxW2UyzwW2qj5sCka2zlAK8U4P8WgxNwH0kFNJdI/QcndgQj
ETK17rtGEsyrfrwergnTwGO2YnYLtIel1Ew510zwE/y9dL0fPgWOPe4fNuV+U45Ic63jJW/okQC3
SnZso77vI6zqO2uO05M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PWolUVQUux4t4HUo6Q/Uab9b9cqpvW8X25n7UKXolDSNH8jiX8r0aWOg29QhpAQEOg/QOp32unYo
TZWzdNCUuSpJu+p4uiUd3wiUOvE6zdF2Htu+k6QP5JbXz6n1ylGW83GQ2AwgL7TG637oHpYo2MLp
obP5rsJg2IYPmYvOwXsHdSCW0knomAFBPAiTnASOKh2GOvxnzUwYklGB75dq2JubAhmycyQKKQRi
3uxae4bqJCgmqLkIwRFPpHA5EwR/AnC1WvDUh9yZ2hWmZ2U4HwhFJBgaYgNQ+UzgBCODhjEjmRrX
4/TE0+PwVC2OAf2fv6es2ZHAxxSo3LnUL6HTHQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23296)
`protect data_block
fkhNGlQ1DwMHavlj20RtZ6Vn1CGWuMOonA261sXY0+7bJSFGkGEOHZUeALdfEZKQXO6U9sP/IXpA
esCURr1GmooTdd9GDkwFqvE6UdsscHgktKdqIKqJGsrmB9fisAD8WoFfGcnHLrck2fOXbLykw2RV
EbvNz7vKvysQUG0WWU/yknLIfdqyRmqu/zylYup1nog+Y0x2Qr3h8YAK9SY08+0CXBba7LR24En5
Vp7oODQtqZ0I/RDJgLoF+vA1qPrGNSl56LzoFdcsxFn4UM94eC72RExehcN78MThwdC+GToC97Gi
SGCvvOD76pbosvzhrZFNf78WCdpltAkgP/wrQ+jmW75PgWelyQvNkpCo8Oh5mZvAzS8RFrgQp81D
sTWVXwGCPdHagdpJxumjvzA6cHRgrM/pM6iQ2F8Ihkp4JmwgHpxeO6ISfaaUrqj9l+XymWpubjl8
zJFbN1vlbLNo2jaGA3TIrVSRRQimFgbv4t2A81cNfeYwJ/E8GXKdKKed/K+ruxcx0c4svcUpv7ZZ
WM6KbIZUOBUCBSHUm6s5rebAK8CpOMTzn7jDeyEEmxTy6v7TsTzeBrbFWVvTIc5fa7gK0URi5OIc
0FBjclM+Kxaf22U26Vrvf2X9aXFCsghqg5pQmPavVOyi3pjbCqzpeu1FZmouB2T1ogi9juQ2X4E5
rdnLURzO7p833qae/H+E0crgK2duAjEI8imxyuHeE3Rs2i9zSL7i/yNlCAPY0/K+t6FZjl2KtNCs
xNlbVGcPAueS1JtjWZ4t1NI95Ry9y/l395CtD9FVEK2w3jZp3Nf5UuAgWM6D8huTUwth4FzxP0ll
R+nQwz0oLcs34Q6HJUkBvOGoS4pp0NNnmJwRwOBTk/8wZeeIhRR/L/WYRMpubXj/lgstSvrorZ77
l05O6HhXYhULDOSDSRwaedLuqX04RgxcY1t9GudoOIAEsQ1sB+yTRHnERmMuTTdf1FQJZLeGuuyn
ZvxS6aXFo2xd9F5AVsRW5ssNZxm25eIo/gFMss9joCDDS5Cx+l+fUNqyy7b1WOawKLRCEpM0PbyE
+ZqesMTTU2VyS8uzhnx49iPdMqhuzSchwOhi4ic/e+weJcgUBF1yR9K9RVH9XDQA7ejId5C6FqYR
qpDeHohmlt9Z22ipZoFD3etIBsERyprykW60mwGSpeMllhBC+aoF4zz0AS0JVb1RqxcmJv8h1Izy
e95JdhdysLxw/Tl8QNkYp7iDa0ZgiUevh2rHc6u4ZxxkJpX3O6sWaPPRq4zNyS9w9f1cZN75+GlH
6HF3meoy3iDdYrcIwAt1mnMoH5u65O97OEuprATjMmsAWCnJVkKjPXr3QkoLBEnpVW979RTAiXmL
qCEs83St9DEXkHqmCNgM1JsM38X6JPK1Ae4h+XZGYFRU0ikzHJ6AhJ+2zp/nAIYosZ/yg59sure/
tMkxJ5UColvVga9d287UhCd+uvP2FBS+qQKvUNM4iSBEiWRunJQL0rSifTBZ90isCZOfKYLRDbi/
MmOoondJPBAejlysLWrCOKAdjEU3mJzg4nu6b0GR+ScfUmrP7JZUHzF8dX7sLTJYmCh4KbHuGXZH
JMHxQiGoV8as7HULxk7ACtVPbpbmmmuwtTyLub3nKiBjprE89eFOUHs8Sh6CNPyjEdsjC6WGnuqv
9Tho0KGPkEOyN2la5q1NyfbysN4s8ChnuFyrOwuXfoTvBQ58dxJ7+FCn/JigWYWPyGVe4dZ2EDjU
6qI2LWXFwfss+s4+bNi1KRpFGPeHEOAOxaEMSZzx0d1wzTOxLUOemAnVzBdiQbg1MJQtrArf10oV
1Cm6o7ffOMWHNhG3EhUejujvBFA8W5NZN1QvX9wh4P4qYG5fsjy6PDMuF7eueOVir8Yx9WUdqiKp
OyFuSZj5GmHjGTj3RBALX25ZGM6oSuHl63eCWeWaGSabcdihZW9gW5DGSWfubuRNuCaAtUj34sXg
oPNZfbe9tVkpPN7BLhUZvY/QxySx2qR0OMW23Gj6jX9ZmV56D/KFZcH3Dbf8mxiNVotdTZq5bVve
Jx12kglazVYGtxN/nDefe7EfWPawv9mwrJ0EEUqhvOeB0LCWUmDNzzTLLSINzqVQRI2Scjb/JDnm
HbnDBngC7PjD0NQjeOaApVIeaJLn7SQNZmn1JOm56/c4erZDGUV+5okYjwOsmEtLDVo6u9wP7hj0
3AONh8ZRNsDYdcU3qGgUQE3v/oOISVbJSJYHx5CQ/dRKOsDzGo0CfU6AfjRs06MGRqbjiUJ8kutG
O4l8XFFVAMUn/xg6GjH3nN6GcpjnOPZ2xxntljeZwojjlDN9ALmveARxWJcc1TRd2TQVmNGd0fWZ
WVQncoiKOaJjCMn3GYlhlmOZSzgqCyBCbxmIbnCQb4P6quw+ZaN0iqqJ/BhQ0civklfltegN+xkc
0qhxDLLyYWNkbrJALlj0fjmaGpl3dFz5S6o2sxRk3mygxfRPtL+buUvFeSXaUSArewVhHX/WUFRg
1jD/tvCyvAKeZFuiu4joRSt40YlmmPbYNMMfK9r39V7zl4IYoqOYWOYIq33EOx5EdV1aBXvYiVIy
sgYyGhL+6tuacGUXf3a+Fngxd1kPuLdMz0IXUHs/cF54KOIFkd3zDgBgNXOn5UJAqNv7ITi3dBx0
eaNHPSPaQSGUkIs2nCAgte7H/eE532KnF3cWmucth6GPq7955MLLGjWxjxgGvwzR3ok8gpwXOLbx
A4/EvfCuf9tKcsNgQWnufI/viBXOaVuGuRnEHJz7kE8arWOXsZxZ4ayFaeuY2BNrMYxHHzxdKhXp
swYztGlT4znp97R8hlOsUKXQOeDFQ1/kPVpxMAGA17Xc8DmyE4Dd2cEb/2OA9nrMC2EWOwpm/JO6
wt1GASKi+/HHsXluyARno5ajxTmR7RiPzuiApVtGbJK8Qww6uhUpLo9Pvu5FhSSlEXQfNyeF3cRD
EklahQIPS8XBSF4Sxg3buWMM/texRLmXLjAvZQK2KSRsIuW41Iuo/k5jblkvwyo1k4t55iQO7Bp+
6sagwVail23iTw9lTouOKzxcQENEtR8OYU2dJBfuYEEMDUjKaxayFTVux9jIrTMjvh8o2MoRBeIW
FPXsBM2eg0QpH5HJY2djJEJIGEZZy2I8gMeb6GPDTj7/wjzGgby8Ai8bPgXGgnaAhzYg1azEgFd6
TCwZ2UW4WxqOXCd3eHmjIHo22hyHJEU3GAW3QvpbubJSvd2mqjh6UZ8Gz0/iBF/BvPuph1sbPeXO
0u368cqvYM1ZZpVU2o0cDKCKoE/h/nk+L8Tr3oW1cF66X7VsBchDWmB+kI9O2i3YErCVh2OSYVP+
ETE6rgDiTsS0U7rhsBrg73jL6iclT2s+xSgMnEDzKyU3N1hSUCqJ59RONbgVH+ez1EftrpGdJhIN
7ktGcZpbTkBZYKWXvrU9ELHeyJDjvhkRMUPoLmjmjmf3eA6st/ZurK6W9q5yggQH9k3+T75JHF3/
5AOaRh7pi+a0LtsPviM83/8fuKDzCCgdtrjR9ZozD2gMtUZqn4sYPg2WVZL9np34ou01RXHh+5hN
zxfL0TcslAxIF23JQPpSfVNINon09dHx2zIElgCes32ftgT8QvAIBe9jEPRoPTrldfqTsLS9fuUF
trNOgiWWUCh+AD5deqFyqW1VNjKT0pSeq2Z+SGyDPqf1a3w7snU+hfM86VpifMD8DR/S8CzDSLMG
BomFB6X+MPNgE2WlNefY7VnytmvxpnC81q3sfAJXiewzs3sqvVS4vMgurUDLSbghrxEc5KQZiG9t
WOTbahKmtelbCUWflOwCRshZCDSNRSZ7U9ezv+aseYFYk9hNTA4+bBZoHlNtQBVuyQlEpwcAK0Vk
R/95uMnkBXYx2Aaog9vFrrpf/Z+Agy5v4nK+bih10LJOIGZgLxHJaeO1H4C+zivlD/b4L/G34Vht
e2ggYaNrV6siT++NH2/lcnN3c4DAZPniZZEezO7p0P8677TkNZz7CB3azLoJOGdSzt7HH5pDLIxk
/2egda1udL4jWRTrQp85dyHcomIk4yI/BtIKLV/Z/cF2lMCX/+fpcFOpouIA9uZ5vj1Zuqpc2Vvn
E1xqXrBGb0S3SeCXn4QsUWWoTymJ2t26S3Tea5zPFL5FR/bAQgK93/h2mnGd2iI5iz/UQuSNvQjL
7E2EggUL4PouCTdpD3VyNhe9+eqKQVR/d1UErl2cOgSAguEeqd9IMizFiGz37MACGQ2fzUlp8can
3V/6pekBr1/MsZfapzKTtheG76Gn53ggYGIEG3lVq+c7MC+fIOJzgL+xYw8NAoMp/zbnVUoyvPBW
4hbVJm4bhyXk80PW89H2+UrmDJjEeqwbPqDWSWY0JRF9Q16sxBMUsvu/62JvUIQRWcSI9H0pZIF1
LVYEMQGqe+HfaikDV+Fa+FLcEbIiRnM3T2Dw3xtDyh9P+WmXesui+WMFbbhA05CrOzMpgAI2Q/U3
mJH3d4knOYtFUTP71mKEXeOBGYVVScrmGXHX2ZO3DWkkqHinoNl2K8zVPfAvw04lE99QVkRNLhP4
9fOUBGCMZUZQ5AaUX/FAuHPm1jWAKpN8Bsn82pjRhdvNVWkY0aVkTtZsPFEYErumAx2eiiG7M4uz
FKyfYnbNxZr824n3UJWgkpJ0ezs9ChgMGJABE4VAK+fuehm26xzZSxAIoonblTBlkAmJbjb5AN6J
sYBfcg+HGYdvQlrIVLt9p6GEaaXK9NTVIqxKlI/NARcoJvuAxCEj3P1pqeq8qd2U5XNh1ZkELEpB
U8s2fPargtjClQn3M02PuiK/O+Ecjj/GvrkMLP5m/LqeyXhAUzPJYc92c/vfIy6gdgBzOTNEBh+H
peDATHoNUgEmlM6JoyXxF1KCWRQ8W9X8sDOsj9jMHVUnBYYcNgkxIrUWxd1L2BOH/iYNaqoG5Y5R
bcsIPG5RjMtEHsZ4Cu4l8ZrXwFpyaCGJCRC8DPS0vNpqyQJ0tqHy6U8iXQL0mPg95X+O1RACiWt4
l24/I9DxOMADS7FACBRkrgTS14yZg7qmFWqakf4tWt3jqV/0B4X8oSLqCJWC9xUhaFaTnH2nr4ZP
hkAMVhtJjxpkcoQw7JRVoI8Z7et/8lCL3YvWL+EvWmzO9TyQi9cOvXooZX2m88vKxXTCsLO3TDAB
dERIWQGSTrT2XUkD8kwHf72HZfjWsgelqfOWq6d5FGPvM/Ek8G08ziSPQDpiK1hDDYfUUR63ilba
5PVz1MO7u7kgWAy23UNfcGR2zywDpgSh1Ir9wwZ/UYMmAXEpkzjTrs/Gn+mZz3blx2FufEoVXf4h
rG2NZzVOSOFSkcngHN4H3AWvU09nSgqJhBnPQz0FwwLfIIlyEldaoZoFNgd0GEsClGtxukqj948/
9EBKUiYGIv5vmqEwRgxNhkIDcKWsDKNB6+YtSuYtDEv1K55r+epPX98vwvCGB/gHtv9+/MRAKXlE
uEsni5i5+stjNWjNwfz0KdshVkRsdIduzt6EyU6lmgm6QbsEX+A9oG5Rtslz0ZG0mdhrbDMxuf4i
5kcoGwatImiSu1mh7kjKiJW8iRd0okK3GmOEhiU4UBY7v1mu1qjHoNGcHKm3PLLdKeRa+I3zMSay
l4ugVAhZhgRFCaSD9vHAIie0AuBtwUgzd+X8geNWTsaEn25WDt18vPu0R5hnIqiLiemcDxTiogJ+
++KYfivNUsK5i01MDTemiM+dA5YKY12yGG3Goivy6XGMdwnWKuvb3XpXHCP0rhgd59R6BzIx5vEB
qYF/831wdmyvkYhs2EIrf9FZhkZgdt4smtkms8xjjZKFaSAH5WgSX2Q1sdZNKNMNIrUn2yy4iJ7p
gzh0FwHcT6tsmNdSwD7J3kn2VjtuJ2zTJ0fKew1RD8vP9wsh4bSs31sF5dmamuRrypVpR8F1Zyfz
X3LmdMMXGx6CtfJ5/zfAXiIepEAMDe/B8MNzx9wOErtrtf9tdXVOyptXfgQAOXOjgSKg5wVLDoKi
6c05i3ET6FNdI1OwrMRKGyJU9DyebRh5OAP6gm/+EFhDzHDcOMPTJv/E/bN9+C15jKIQmE637D6U
VD8i7iOFUd1y2uvk15Z3T6Jms5fC6185D7I5fpqliP8Mb0P5tZKnA7t1dCWhUWsEKtLZwlwoK4Hf
Xd3dDkMDeqHS1akIN8zvUpEa6XjfjM9RRjrlnSth8GjC5hrcgg4IucrBrk5/9UTWI8YP7EZ1XMwX
KhWCAw/Dlz0AJeGCxNgR0HIDdxuyBZ2JttJMLMwipWJ3tcZ2DVEl/qqZgPp6OZv/zQwK4hRaMla2
DaQuUfrWuWKm8dQWeSSJMLn/ss89ANzutM5aCDnSUJqX+BpuGyq/tej7W1b2kP9Hy8RzMnbeNbhL
VfEv9xheQ0coYE+ufkCrodna22AQnT2LfcQ5d6373tb11aOyRuGEeGSlzN2uws4E7Ly84+cXmLrD
FMyN4ZXh6FQdouVfCsh+6K5oeTRlNIfIbmS9ahQ7BV5/UTIVH61/x5fbI8Hx7ntsM/IY+cfZhfoI
2OYdOmWvOEGnGRTY0xs6O4gNBSgIungsAp2bk60GgpC963sXdEWQT3at+K7pmZBiQYvRNsFJczls
JqvGyBYKjDsrvS/RB31ZFTh3uYPvPCzeplKGXUZrB4JTR3HM73KY77VHVhZSXgo+6oIZm8H9yhbB
FzbY8Stt4stHRtmb0P5/Tqi4x8FVKYFfqrtdh9WE4opgrjmEN46gO/heX8C9dL9VTFAFVCr0wtkj
cGVuSLIPuvtXooogaJza/y30lijNDy5Y10n7uUUxeDwqg9u31jIpToH7AeZYN7D5oDfkf7C2voY8
h8KN0n0/Nu5o9l+um5rG3/TmS5rxhpQg4NA2gCjYpwfu2np/4zybFuITARfJpcv87XJxjQm7vQsU
rxfpJrI3DWnRV4GHXZ16HSeFRP/zofomDzy7p8eK1ou6HS1yBSeKYUEqNMeOYcnHlq2PonbXNvjE
DmFfj2iyUmcIuXuDRdNMjYOrGL+TQ9qknxS5aImy6FYpkbCqjqQWhN1+UTkRak+sSXH5hcZQKkr1
M05GHki3/cc6+US7Mz0PPPb7TSWcTi7sD1CKX5OwTLsNMAGrN5h/KKE8lZqH79CSNrzfQUbaDrhJ
UsFT/44trzZGUaig0+vkEhM3yd0MQstTZncvmPeqVlhJ6xfFT6f4QWAt71Eu4T6MuJYVBcs66gZI
AwqOQiaP6VcmIv6ehrXCkjUrIWKmiG+pC/rft5j+BIIAhf6knFWPRm6Oa9pfFcJ+MEcpqXX7ujs3
bPFBxVckorE2OlIfQ3N4mkUZsSpGcNlSF0NXXo+yNhESh5RIVNyW77CHePPIXuFJzQ69rhsVyQTV
iBTgl0G3ShlBSsqYVtBU/kQe7qbxlk/b8xFPGXS5a3o+t1kawAY+1VOTkQFfLlrIT+0zR40qSvoT
0lU3Hpo55pV5CS+9AqoD4C5Y0bf5Rn6UDiT06YqyFWbqvDAl4k0rXX1Rtf1LW9O4G86i3K7BcvKV
tk8pPO0ocPI+PFeEprPGhC6VJfqWnk7zppkuDnPSpagXks3p8MGeZuI5g5Y8mms9TTT7+WN1cZvq
2n1FUZPH9imQFBTBh0pBurh8xzQUfTeibtjc8IGzFdYphTlgpJROy0Y8HG8kRUW0ob/XjGZe6UZZ
LjnDP/XxlDNFhnfYuphKEe44i1jYmkEPiXZ8Z4Cc3aTaCMiujMmvV/tf47XzUfehzkdTyfc5lzwz
leeZhGI/QDbeURtb6zx3SeequfT/BIpkpbtnDl2K4J3qbzEqHVGhiDW4zwfQc0b7rbYYvSvTIFBG
pTR3OkQZNGP29PK+68kdO+M5ySAvaQUIzcVC4pb3TwcDTyYLhWbs+G9cr86imRgyKKJ8UxuLodU3
cbWrlz4QR2pP+pg+zobKAp86YIbd9AD9ZEOEIAfaiPwyRF57NJCfWlu+/wwKH3hW9hXEflmgiVoB
yzC5dYRF6e8ehkSBLVQDxiuq4Rf/lRAoPjZ9W+KUhfzelkjgYr7W0V7PC4lNzAX4aWHR7HWiCC3d
ngOjzwSlG34UmI6oJmsJRTkvCaviwneE3CmwvIS16aOWJS7fos1Lu+PJNtnvF8DZxAJo9+Du6syi
te92dluD1NqsPOGvDIeG9EDvdiBT4b39HkgL34MTGk8OR1fC4tu1Hi9O9Umn5fqhgWMeDmQKGci6
0H3eX4/sXzADHnkCimXBEU9o/l+pN43kdSwUXLBLPDuR+xnXbZahfGO81FQLvsqwA0allrmgJCtA
PxnD7BfdU5Ozu+qPwtMZubR0Wg67/etvwVu2NkiGXeCcs6Ya/cIfvCajN9BtI4buzn+nnJ32gn3M
Gv1BPoJJUqSP0Nozqg9oEyNQyOu4cPgHhhE10zxYXLj14COZ9cwA5ZmhsF10E78lKxCkxKZi7jWg
dPWAi++XFnyQqSJubh8gofyWyumBWiMmONQtDCe873/54DfQgbpptVhhqp6kZ1LEPjOvZT7mYbTq
RauGYroStetScaHaZpDsmS4LnmlzvsCwzBtUDL6ZwyGsj7yWgLVQB1rfjNP5YyPb0RxXBFt0DR2K
yiq4LIiV98BTHlN8vER53BFFGeP9BZrkJo9eGvAD6S1mqlqZySk89s56uzbviHZyh3B5BLw68nhp
0ezuC7lx3gHwZJaBt/IbUEn0W/1UvgbW+I1jwg8eIOaICBTxY1WK71yKcjYUk942N+Y3tOXgHuHb
/HVYH/6aqbqvNAj0aBq8zOX/BXmvK7GZOrtmAyXGZb1qrp2SIHt+yWrxerraMj6YlpWmUnpfrTb7
20tJYQlcaguuvlTv6KA2QmWo769OvEj2E1ilqmddXX6aLoQJ51GsBtfLWi4TsKKfFQxxAY4yPmjt
ldxFJekT9JzJBoDx1chjOHzAGOfWi1+0Ko6mYS+dAZ5dJvMc3NPmTbKTlIv5yK95Z9cTgNxm4+6m
9JFy6lKfNlxz/6GEZNYlFuUkZxSX1pmb1x4TWPUdDe267nknJVijZl8AZnXtsB+lcqaCULWzJ7aN
IVQtG1tGTtXCRd4mx8uHHQK7nAkDIurR/5ltYgtAb5GooCO1O5UF7jyhgQaGOXcGK744rzO0cupd
8TUWa0rceMlSnFPjscajGcAXNelRioZmpP847pVhL3t2zV22v7gfN4RlzROx4HZvjIZI0jBZuJzc
E/KA6NRFs2gBhqtPpBC/nFP0d62IWNktyRrGla7hcxWgaeoSgK0vSu4zYGf9+n5LI+9NiaG1QORw
IYeceA9TEu2WOyfSpGxYCgNPjP9zY2A0YgCJQdm0kLZkkr//Q9SfmRjFfZ+BMCP5ENzzQxuBqLmg
dilsyz9n8pYLEb95K6qJjyWu7iEoB7S2magy+kRqu8jkDR5TwTv8yMq++jvze6UCTZrM10esnKwE
L74p3qs9dsr7HZk4TEgsMHYcIJn2bA7b2wS3zKvJi4+emoWubvPJh0sQAbJyCT4p+p30AU6jtmrL
v22nl+06thHo5EQba1fKI1mQASu8EFj12lG+NZcenL6an/ZSClI4xL9PFq839UTc0OS07pa07wmu
D4DVA29mBNeRIuHsly1W2OaSVpLI4ok9LCv70d00fHxqN5uh6havO5Ztk2KleOsn6504ReB+XA/E
SfSASgrf4UfB9SswGui8SIZYQyutXHyggKBq/xSu+2DytxL3kDyGqFxiqNmC7Dw5CMrTwmLerbPs
Ym+MUwUnFEh/CCDskAColNSP/wsCCUBQ/mqIkYRUa3dMa09crbBALUZourvYHBBq8HLENReEln9p
jcRDd0uq/Q0T4OHbkof8A4rE5eG9llmLLDOWyAkTOA3S5aXMFW6wD8VaWGOW3wbM4lcWdG5K7vLM
jrgjJ2LmxrrWUaPWChUK9nWk7tVsZffGRTFHJs3stc82wQRvpHRk3glX70iP7xcH1uZjkSwHG6JW
CP2TOPuoOG4XaH6SaZvipdDieE42o00KaPeHTfqKQnLWYos9IAbcdUIO4zIxwgkK6sIOAzgv99eG
pwLUFUarJDxrN563zwFveOud0rO5sJMM6cjZZKxV/01FFhBdu/LRg2HTfAJXFYTNfSWxtjzq9vP2
T2UxweA8ZAebk3nCJ2gYlh6MnaxkIde/+LoCX/Sc5sPklS+riTmN6IJJWgIY1BZmtlJqON4TE9zO
8OLWufJzapUKeyQYIg0F7mig60SuHcmx2diX7g2wRd+dpsAd+8LfybRMWmO408RdPAlO3mpTMWpz
i8OPOvjr7x6dIDRltIkA0SMAfjBZEOJ9AoSJolP0v5jOKr1fhKzdE/szQunrH9+8ZKHoKQFjzFVX
yfje6B3UCtNZHnOYW+O3NQGql5drD0Zq7PbPNeRtEIXU56t+73eo5j+D/ev8oV0b6Kp1zOCcWA2i
3nr7lfQAJ57o+PWdpeg0Pai20frXY+MXxvm8rrgMF3DkFk3TV09xb5L8G/28Ze7+EpPtTFhkojRB
SjIGzVc5xKFQ8hSZXQwB+EsOMqOMYJ9c5iMq387idDHNA9sNHLsF0WOt4FvfFzzCRamuz8+F89Yp
s1NxeYiTi4jAFYzjyJsA7Mahc83gR95lwPdExC4lf3a8SS4oixVN1BWO/0KkTPbJLkU3L52gfNxE
VMMPko4esJaa3LzlrQH793fplaiWqI8QXzxle3pYnjoE0OEi3EgtP7clc3gLftg/bwobKRWfBcox
qzGdwkMUWpl0ROQhIuk9W9Myw0R5L0nE0KtTzlxGpdGfbVijKGBCdnJBzseP3Wjv+AWAmO1Pz+Pn
N6CARXzLsre5/Zzi6R8D//kV4mrfutbcKIuxYF4jPbqCvW1vzvl4HMAAaajkL3HggrSNNQu3xO8U
OaQs3elktdizbLmECCt5cvAw1PghNTnYMWHXN5V9A1Uc0Xs5J8dPospWn/+ospZhvuR3fkIonNo9
OQ1t9JfcDTq0AuarxkbgF49ttK4V6dGCxmAQLBXDqY/koqFdLzzDU5FktRNZ0XN8g9EtYNdAw9e6
N7Ap3PabhtqYL4g0bxc/c7ROUFiFi88Mjuhr1TN6EaYKx2H85sDk/CL5ImdCAozj//v4J+E6dhGm
4IavOzt9Ln8Cu2MNOu6tYGEvAfwwP33cpek0UAN8XDVnPmF5eCmoc3vFYsDUdNeAwOt0f96lht2A
NDFEqkxR3+ozZIKZSlKb+rfIT2c33M4mnMehPwUsCpKGV69xInl3Sjh8O2IZo7zjGpdKPTG5xtjb
Hc0fTiFJMlX/esqxnQnaWTIEyPtvopEU6fNdujLboet0yyDPzSwYrJDhJdQK45ASb8WOC2asGpcp
memQuPxIPkJCzA5eekvK3gUzo4FTOpEINyc+6kcuf2tFrmMfy2IZCDjxxkzhYUHTYFcUz/20m1XI
PmFBoLz+pTEN83t7N8h2rrVR+62H7SOvEFPjiSO+wb/02kTRdyuAOQPnsjHhpimsQFfY0hLFwKBs
agXB43d2rSs6iLsffuN3hu20AGWG6tmKYO4P36cGaF6exLDb5OFCvCdADY+KHmyARp/HB6vrAN18
ITV9RZ9Fm+X82IArdrqMxMOdy21JjpDPj/udW9SfoisRgY7Ye1ra5wQZvvXgdvEyd97IC5vG27E2
0qgXk6kzuqlP8tSLannBNxrJ+IlEpvcvl+r6VQm+27On2N/SfGrB/lmr6hXqmrxAlL4H83k/SsqR
f7/B1CrVjhNF0NHP22x913OOFBpg7/WZrdcXBA3uYgDMVjxgq0Xfut4A4CQc7v1GCfS7UXJJELpU
OpkAc3nCU4BzKTRMcr4pS+k0j8JEx9Rz2Fwgh5JZ2JEnD0YKWXLi4Rzc2IE/Oo6lU12rw/apG1oM
OD9++OEPe+YqRbH56iUkACbxKXyH72Cs9Q61r05eCf7YFNUk+IyD8q+7mYngRsCy5B2VqB+cAasd
0iP8Gh0+qycE8ejv/Fy0vxrhhrBtNbOpus4ii6F/ZXgDTy7ix7S01poujX6Sqfqh+WG9kZPw+8Wf
+RGEOIhAH7uG58wwl6LIw3cX89uaL8duyCuuNSqoKF3zDtWVd5CbpV0bGYUifaVhzgnLb/qZ0DLt
iUx3Lbg/2LerW9oEkBRDZjmzKddQxYZXI15t5xl8bhZblOuVxcbuhYXEsgk0xZwtbMTF0iCOZkTM
3/6JahOroOiV5j0ejBXERyYWWoUjgQNhgC6cBydpKY9zFxMz+a1dOONmjy5HYjgvN1giIfZhM0Ax
AzMpLTcmgTZ0groiHNaFC9clDDYKZgTbX6E+JAyWGWh4I1N+v+nNh9Gj/krpgqvKw7QglFgD7fXO
DrjVVrQd7fhE/uCe9shHIIcW1ihvEExz20+YQuQh0P61WE2zKejPMSqv8RoqGnP27pA61Y80Eii4
+H3r5xkGjGRbDa1TRHLCkCag0l961l7PFkyR3z7FkubOl9UnL089xbcMO8QwLOfCId52n2a4lYUW
GSqCsLl+G+MkhboRvh9KDYEL5KHVvPIczkCLjAL4RZIIokwoYZcQMhG0u6e4DOUEpkAZUSk0LAqB
ngoF5xpO1x3Cz+uUMRhO3DysNo+h8MnUrh6HMx+DwmfiaGKR1VCzgNrD590Tc07h0QINrAnrOV3S
EabCxxcfhsEvBkCsKGNWt9Ub05OPJ72JAwI5OzyuuYhZWSDWw9Jyg5kjbyjdmAg1SKKnA8BOvzYP
XgBOwi0tw0xKg78N8OS3yg2ckM25Tqe6lWjITwp+XWakToiIhKlg5hD+pkzWo6Lq/MTfHHskQmQ/
NjQWzf8d3bMi/S/f/y7hzsi3jWqEqNsHJp7IRr/TS9iJUmdnFCsUfFzxjTHfokNhFcpptTg2QvP0
CE8zXqycJp9vbRUVGMJI5s7iT3Zk3udhRgTSCZzFjPkiINtINfljf8Vit8DeA3hMTm33wT8s0r6x
N7QqvyJYvyLHv73l2kVeHfGX/S2t/jV5WKBQUA/yaEvJ4ITtIqfTe3chHJsmdMAvb2ewW6ezHFG1
LP8IifOaoqL4WlGgO7KYGg6yZAT+dg+ZuK6mWdyXD7XLONcpHtNqFsMbyqDn7PxK92irWP+2MMYN
eKhbDmtnCnXgS02MY9p0g4vImUuWW2hF9MnoqcwUEs9lh0GzCUecL6+pNIE0vuqFWQm8x0h99BLL
vOrj9eL/nVZyc8Zx+OVsRDwd+bmD3VNcSAZuAA204BfJpaULRzbv9vWQhqZkiQo4XlgQb83yb2k/
sF2sbN5EeB+IaPojQu62IvimiuMV0JGflJnRWMiHKdnV3vwB4EM0UW0yL8OFG92wSvh0+QKAbRYR
rblABCZW0Cmt1HZ2u8yVsa9v8RiNagmt6siO8HPGQ8j7yGEMAYE4A7+Y2fOK5bPoRwtmeQOUgbbP
TjQ0rScT73wEDh7vXlhPxQyK4lmKRpsD+w4CKAofxv1brlI37tvOIOKXLL5qKQuOUbagGdKvsgAk
wNPeJ+Fwnl5rLUgRNXeY6Jq6/ya1NkjvBNUS+Ma5gEETuRzRRFw5rfCJSjwz7/kw+T1AqCY7CVPO
08ABkagWbWSb1z1xcgbUnhKclHhP95LDAabkYbNs04dOTHW5DK6DiSzoQSIl4pmHD5+UIu42902d
r7iE5cx16mkFOXRPi1yT21QIS3u2h8K972GTBxzUgJAKajlbfrB3oexwMgTXUpSFv3yFhurF9DXz
KHtQ+TtWW3V5LKe+16zi36ygQ4u4p+SXW/9cVZObT/+7xcsz5iwTch+H7kKIm67BAvR90ZNoAw8G
SdOSFizy9tq+KGXYQfrgx90x5WrAN88l+HjquHPZH8snCWj/v4j6uR5ybuiA/0r3l4THX+nMHv/M
kPi7ghOsDOhuQlXlgWW6qFe3Z5k0zRLr0et9eYHQ0OWVjYOjavywa08i6nXw6CGBintFXxBZdaav
psZTOfQ7YJpoNqEvw9/UYC14mKZH6O+VFn1fg5OlRDlEjh7yhv8I+4uMMVQkgJTH4Rkb8swckX2G
AMLC+gZ9Rega2tbW5JG1zjuLSXx4Q/RCyxMVwqOTIpkK9P+pR7ot0dwaFTX8ShSFXuRXCAJFLIIc
vUqmND2usmd/v3kXABG1VtObRSppcXaG05l9P2uMUKfuavc5NXXAUwWTPrsFZLfZj5BWg0wmQosU
RXbYvMiS+b3rnzQ+YwZlFxs5SNGaYt8uxsbfW1iD2yIRb6T3zL0wROHroWi1g3Doi4nPBF+vEy0Q
tWEaLD1UC6hI4o1OmvLc66pw7EowPG151shLuvXDbU8vkQJO8d5bgjEACyLPNItblWxTZbQGS/Wi
IyF9Et4OTJL8BofFH01uDzCdo2DXmKGNu1jbx8jpBrdbfBLRv5hj27XJpdEkDZVUeATbE5KOomu3
nkaZ8hdcTmCRXFtLspxlO8cP5MVpmFxgZXM3SI/VlWDXjtiL61/x2QM246u62bV9ZoNfUGgvypbo
TM2Vf2osuBk0yZIZZq89RNzMXuDG6kXqe2T7QgwrZ+rSQgoX78Lx9/20STgGgqBWFhBW6nG9fjTO
1BHd/gEc4/PMe05fq6TQEVYtsqTfwerXNAUWe1BqoePL8mt4b7Etw38Zgw+B8dIcUlk6smK6V+8I
TNRAewDJdYj5DoSez0Tlh4vlzu/fjMQlEhMea8CMCJ6iezVCjK0GOrkjXliFCYD/Uka+9l56SjR8
ohVTJVDm83C/+79CawRNmDQxcmLJzI9K48MxuvYTj7MN6yVQjya+HLQSU8OkBFAtGxZ5Vn5+QbXc
3UWcHY4agqy9VEUUmNdvuGzfNviddsz2IEJCcIWfePYyXcmmdpXVgpwgYUR+MLRjGVACifB89U/y
xNhF5zMpoyp57qbNEilhVgQRq6tGWeOlYcf2GsXpGo55XGWlR4GWv9x5jYnqDW4G02H5Gj11gLH3
FLva+YeFq20SRpSz2/wdcn/3yoIdXE0qXI1hTuBgDT87D5sN60A8uJSYk0BVE7VIUjnMT9uiIzKs
34Et9QRrFlINRmJGZvJQyArPeXO9TmQjaTAE3jDWdxtrKhh+RxSdmLpc1qSqcZvrHIki96UU5HWa
qDhk5nGQyvNdM1SlwA90pGdlaWbqv4ahsRByNzywGRGtbhn/h79yqm0/qPRtKePG6oJj1bMr3gLv
HJNMLJI0rK1L+6h2DUu6i1qgpcX/L+D29e3sZmjI8OqmeqZnBVYPvNlHM87zfT/XaHDMsYY1U3Ja
SbaTA/vbI/6H1Y890qGEce5VwN3QbElaaDnH3Kkq3rI3ImMFXeLRH/ToI+R1dI+FGEpHjN65qwJk
9q5/VIs2NO6fA3aphn+UmlRcv03ad6wmuhJyxGdhr3v1h3BBKM1IHRbjl71Jq400Je91WkopfKA2
ZIlb99B0j9eKHEqv7BDbgHz180T8gm8KEbX6iFN37fYfxc4OY8YYSVnCGsBKefwXnFaqeWXtXpEu
iTL9nPa1vAHa1eDb6j+5UAEsKeQTXZNSaZhxfKuCB4fmvJFF1IowEkxuQ6KDSdS6e+n6GMPvLQmm
L1w0ZIDzLUiJYNKB2+0cKCFTVzoK0pLSc4Yl/xF+oVM4pCE6o8c1fryBnuKGFqCCUQTRWkQrz3N2
2xvFdWOBoRNv9/3PnBuBGk0Al5bY8FhOHzqCKu7Wm9tKr2BesRmAyNNUO4o3vXgTmKSAfSwfIiN0
aMO2ZhohAWjHnzmXhNiO9R7OdR+c5phKdExJd3QQAFMRrXSz3S51Q41tFBX8dXEcw9isSQaO9qIY
wfOcHizBveyZ5eavUYYDAkHeYARVUYVf1sDjoX1s52eVd+mqFSj7fGAdKNCNDbiyWobT/hv2mfsv
0yXz104NKDrsfC/i1nBCk0NdYWeGPN/YWXHcdCXuSBceBwCAqMgV0sXIM+v5GcSRyUMQKMx8uFPE
BGJr4KDFgZx8no5YcT6GroihSIoQo8EoKWN0jdxrIDcNGuIJdU03hwlQ9NThhto5ucF97Rw2xVoj
VWVsAz4U1l4AdZ9T9GliRwuhvGgOeCfrAqOw2ytkOk4PsDRsgRo6G0S5Edt44Nh2wqfLhOhxRVwn
AhYBizerPBkegmYnhHQUIu0Z+N7+YEa4CpxSJdYqh+YjXDbprbNqh4UXax1NWYsQ+e/EAnAEGyoH
CUG8YNz8oafrU79twEqPfKEqG2C263XqOm0ChHVlee18pKum77w36KL9XM75wdYgvFCruQDKhGA5
y1CPKNr8y1oFBLxT5oJmvZF59/LBXvq0CiALvAqnes1Y50pGSLdXEA6RGO2mT9R5rdcoDyv6hDC5
m1wP6ZopGU32yuHklmMl7+HXZDxjXaOYQPG1WzAj4VprXYStLNyDdNaG0HHjMqUk+5zFH0pZxBNs
pbsyNbZe5XGsqvGJChu769mBVRootpXoVZ/xiSTEANh/QzEzJOs2E1Xgvt2D/5sllBSsCn0bEUOo
GxS9HuVdCSoRAFw9/RtFyPGX3sTKTuI9/i3i0UsOoHn8L21vx0g/cB30h3wxUox3QszVv4OPlzlE
Mj1OYqP8Xr/MX1rbuOFrahHQQp02WDbWoI+As2c/vGI4kUBs81Qzi3VgK1iKwbspEuQnFfkMz0PY
yaE3rc0LesxOF144YIFnKgqt62dJ+OuRGWxhCzMfRvyOFFX875BbPHDrNgq77/SMXnVPFqaDHq5S
dLgmBNiTqFGt//6JjdpLMbk3WSRQWo7KFSBx9oIKJVyF965ITHhp14TzwdKQGfMAdoxdDSsidmCR
TtCipDCY2G3KbJI4C+sI20rTQ1pDt3Guiq6nYsbCwaCbPsjoN89cMXRLocrbU/s3K4hGc9U8Q7Tv
/N6FoRHjgfokeBDbIMuoaXuZDd7cXSMMr0xIy+hFOphfPWctcZzsxwtfOGvVevYowaZNS2jd2xvw
l9qQiLFKLSi9KIKzjFRbaRQFTnRO+lwXqrASCiCT8jW+aw9Qx8p2FRBa2y0ansOExgptKkTim9Lg
2vYaqgDb8Y7MwhmNFHPZIVi3RVkwMM6QGtGjflf6srNYxtTkVDa+GTXS8oFcYY4+5vPL8vkcxlGs
/6/Woabk8cL6IV19TbKwpdRKAF9pKROekyeKGxr6dp225+a6hhBuhn7qi5blBskpy1LmJ94BzGq2
SKuPCtrXS0riJZ9/Sj/Tab5HSBsNcnoFjGx4mN0Z05Goy4x9rEFqO/47Le7LyqcYJB/FYCyiXQMF
+HnvF8ul6SotUZ/0MgOsFOk4Ug1Zr+4F9lbEe9/9T7jbcIiHMqXV0r0ZwJ27i/u9//tNWPI3hUXt
/N94Kk1zyF2MXTRDyEfL2jH9TssBYSf9Gx5DLtCN9OgBCfKB1Yhwq1epWI+5XT/6AHTn1GxWnnln
RQ3uQS5s2pfRAL6zu8YhTkoUdJddFGRPElLFBn9kdGLZ07beY7Z16hhYH7svvibvbns+YWiI4tml
ciDay79761MU8BpiiY2ZJvWYB+nK87ARk+HJaw4lvvahuYUkgmvM4rzDuJlpNY6+Q0cwJez5dn5R
vStoKgiOSDXhnN8/WpBJjqdG4mm+aqt6ShB1UB6u2NLGq9qONgOrMp0hqq51URmP7/yZR8nsls47
Ry53LDQjqFDuzqj42uqwIBHZroEtvH6NBoTztXnA24NZlMhHulS5c114JRO5gkj127uesIKYpd6H
k8XfNa7ZIvLvybhwp7AG2h2Rykv79ZZoC5lnvNvcdCzMkd79+xx24b81ukFW/rrulhSbJeI3laq/
19dm2rnHCD7iATDM809uN6FG8hieBigwtcp1CTcL4vmbMurbC3kmM0Zh1M+oq9QcXARmg0k0BeNH
LdCnYDLklYatQ7xA4QhT/y9msdBP0H4XQdBx+CDQgeCT87pkGEqJURGnWI38z1sOuWW3jZQRLzc8
DZIKjLfiy1G6dQgUhFhRrJGkAu1IA0A7v4LAoJfScpunAvjL3DJUVc/X2jOZOGCw40YsEY2Y3lyi
XlPRQSlidcaSZZPFjdQkncQjlBoQxvZCoU7SQvnKYt85xNig/nXLUm4LbMA29EWHSEfGjeqK0nR7
CcXKciuqFYUBD+GvFVojBa/YW/8jH0zR8iCd5eD8GOuUye3T76tNgwINUcfVI63QIpCNPqrPxSxc
T2MPICppw0Uda4fjZ6rZZwRrta45jgnsfTT6CU87BKvj6AX271x2c1o9jnU23p6E4eZPe1DBDI9Z
lNoc/UYb25hzwr49xWXG7LMHOuiC2pSUNga6T2xyEz/7UrA3ZGILFn7RUGkVMxlXCTVQWOl8PVQt
w3xCNNabN4rOyRhydDZ55dISqjF36YUsvxANY71Kv+hxLpn7wV74GZLwHqYLcxMxT+fO0Gx8QwdF
rwI1C2YekXI7rTW838a5sF8IzUA07pzznIUK4UXwoX7yjMRauCH9mqzySCLKpXbD6mRd1nOJojSf
aGHVBq9SxCPnR3U63izKjR1GpscAlF0RO5eA2pxgH7VgNVb4ynPVhF2zH5HjN7qCy+s3kH0PD/18
xRmosuhwqUguvrtJIUcCGX6Y77dSP/QRg6qgFfXpxEEpb76Xp3e5szLVDh+h+HGphiY8Xcwdgs6J
xBFlKBfdlRm6pWAnj2BDqy+2Qo2whlU/R+g7SSFawmO0cnt1kHG8UC6myc5RBBQNLoCEBHEMzpZs
l4ql2qohLDZJqzKILHBnQ/mrenhyNR23rj0VoKaN5WN9jgHf16QFbidvMBR6UZhVV9FtgoES9PJG
NVSH7Ypcpt21ThGSikqEm5+AaNAGijwyOY7lYka/QgZwKtwlFjHgH/oO2rf//Qb0pdAqQUSOpMyC
4NAZVgGcPnejKYm8e3itAqHL3XR3m0q9hI3ZUZRzhnar+FQ0eSG1oAIzoa9ZsOMop5KraUhyHBBI
LCQEGcj24klVAqvNJbP16Jpitr9OIIPXrcmAQf/e3wdYg5nccuT2LXd+s6Ei115COnxwvSGQqqh7
puDyxZk/1c1AJ4BGhArRCImoGtmkot/S9KZTWcG3iodLut2Lg/O0PVKPAPiQT+k6wsMI4aoUR6VN
EkkF5QSlur/JkpthHv+cUOncU+yT7+OUH2tCXYSXqhxMJ/AQpqjQAZSmGz+ebqX0B2O5EKtnl1s6
0wtPHLJ1+mzJuUNPpxVqp1MjFFQyFIFTP/vPKlarTg72sGJ+ZQBOVqUwCbdbNJL1b2cfM8LS+5To
/DW63qAom47s58Yq8uHXdyOT7TPsoCfhkvn9kh7nL96qdsEHOf1hfICpFWxVqQbFnlpvkiYFQU/8
Y+LrIcReAqNptsN/wDtkz/M9eamgU83UssdftBuAXYTgVSqVzZj+Za9oBMi+WfaRcDVIdEfUHhWs
I7lADMzSjtUhNjSQCzIIb8f4qzP2F8VgjamGR8NVQzhkfql1eUupOKgEd7UB8uT7dHLvZzOqqNQP
z/rCu2aZZwcXBsbtztjwVVfluz9EUfmNbrdbFJfYW6b/3jbYhGhVJp6C8lC2gUAYifuOJzaSbBUm
ScWjbBsdV2joBOZiAW9V/+rZ9Umu0AM+/vL9YuFrTdfYMLsm5QhGjaut1PnpFeTGKAPrv9+Mds2O
hK6G0zNrYr8T1SQQ57Bzj2FTkUNo59CJ4M1SiNsaQulnjwJDX5A/W1GSN4fU7IhbpO3hAY4BKB06
x7MA64sK7MXiTSC9spbohLAEpoikLpv9rQXNOruQ+cS3FpYwcUjMLno/xg5RzDc7r8JPDtgXHtkk
E7Zx6cQKGPYYjasYTLYRWdCRobsqggIjG8K7H3AY31ld341Hq11MNsqrpLSIBx2pLG3NHGnyQPpC
7EMcZ+LWvWTk2cdbYVVFYB5d8d9+FLeN5rjDPf57lrXUnLsLEc9g9t3mNG6xj3/Uood5QGgBbz/e
n/PrUBhD7Nt2nxan15YUk/N3wge5dZCYXtwnAWjubHmwNA2UogPUk39XH/EOMeqETrMSIVH82Niv
XACVUU0kiXHOtxMF7KWS2Js0cV2lgjEKHtBaenK83Li2vBycsd+WJBod3pmP+Um4Q+ftdxw1lFb1
BIvDCf3FsKSIbYfB6Kj3WV6zhJSrfiWKLyZXCiPAPBeaewvplYWo0RkMlPPRCE+T7A2ouQ1kVOPY
JAn7MLEfuq1us/fp+MyF1OVGGi/3SDNm5FmYKW36s6L41ewQ3z9LfikOHzv4/ISmTsh2z7NJfTR1
Oe7/3Mk8FcigI/A35NytAkNoYOjlL/66p3HKtuCmZRzUqKWSonmew5kTUV7bxE83mKRdJDf30jiD
c4EGfJROxxlQzskyntuvx4ezp0YROGNVaANuI5o9WJhJl0xi+hLlYSFVjATo+WjaUZ278eJzXhuP
3bifKC14jXHtiqpwJO0xqOCEyGmEGgqcjJB3wVXcWOGBJwPdseTn+4efg3XH/NwA1eweFpXpFqcK
CWZ2Sqq8ZCQ/0GcrWQQMpblcw3BS1ILZcYDaYXMhDyQX+jiX3YHobk2PLuzjs1ynMGUDZUjczLUq
Kg6KK5ylCOco571DWWDYPG8+aS8Qin+99deoF9L47diQNqIWUft7SCsKovwNBr71NVtvnbBj8v77
rKzpAYGVFa7h5zk/EIAoqAEvMK3BmquyXqt2a4mJFUbuy5iGjYLJnWrqGliGMdnK0d/tgE0jZlVp
KgDDAQAPJ/IoHRGxG2dzqc28Y63Jtaq5q1K8doWMd2P9gbPwoCo1xGphk1pDHPFrXxBSTNmDZ6jK
BeT94y5ArZKobh+Q+rVLCqGoCWeJh1q1EcoFc8mY/0B8hJJi+VxZsuCiW5w6s5XLIsj628qnvFSC
NjFkdFHAuy8+y/zsAlkK1P35+DKKSkM/5uSyHsZAH3Xcas1uCSAJ/SCXP0G9Rv61JGoSOeRCLrKt
+w9wGBOAUM1l42/qtTc7h3YI06lCFLxDne5gvax5FZVnZvt6p/8YZWXPVEXNlZwID1VQIPMCDdAA
PQAvbF6AUgJ2GdcY+MBhmk3Q9PGYdM0WH38fsbIjxzO7PzNUfP7iKZ09XHvLbFXsDCkS5/VcVr2U
1XtgdgNCrEg5lpn4Zi7GYBOp0m5xnDvawyi+zfwbJJCMuIhW0ZbNyNqa+LC0ss0b4rISm1cv2cDD
FrQu5IS61TV/RneTmIzIiq54qCY+3G/ikshhK0+5Wl1nY8y/BPz23ONpAQJpNcP+PmRSx3kFdXNe
swEGqiPzzQBCr6PoKtK67IRcsjYjDC/Rj8S8dxfTvfOyhS/xph6mi+mJUUPVIH9tH6wrfOeYLEt/
lT9QiTHrEBoaAgUMRY3T0bf7IY3kySjxKhvl0e3g0bHtYR8l+UFQclzi2vzcVIRtm3iSnD0snIUs
x2mxwKOkJKHJEdF0LdhdzVkAjeMTHvhWnLeF9Z8Zq9Pw12y+fEHEN+AafTxWFJRt4CzOVUngDStF
xajvqBJGRK3aKmQrkJfFl5cvzK35QKSMzzv/lDQ7qAncQPxDIB25hWi4Z/R9bnPnXCGP+jefwV0K
dgD5a9L0F1fAW9yHurcv/z5g9CDUoDo+cF8OUg7w/fod0hOGWahybddx+CA6qKgWtecwInA3r/pT
8Gj6bVERrpT046Sd45oDKU9voHr06ZWFShsrLeRWopKHoFl7kHGUTZvniNlfJyomqQxotdEM+Nec
PTCROfKMaFRJVTLUPrrqyva9VE+MJgWHDXN1yvWt/gHxXkK5eYS8bMt0/nrxNq1d+LIfkuPeG9P8
MhEYNhn5t6jvbPDhd3pRXyT3pFenrM7SzjfC3243Y3rdlKjYJ7ELu9+jVn+oGOCVuVDOyn1T9WVi
1Oq8afKw8gW45ZB7cVACkSE35dTL5Wp7mEWj1vUSBtK7Wi24ZgKWqnm9DzTbMSOvTXZar/N1g2SZ
NYf6ssIRUGC2PcEJ682NZzLxQmtcV1z5zP9FtuhmAkhVS6wIRSAI5llQ4ean8UlzcpRa9tCVHXgu
M+hvoE8zcMOejWRzGqVUCCu24z8QvPt3bdMjznyQJp/WOn3CUNfJ6FTcGyru15pBvxbS9Z96YIHc
orWhsc+T1v+oo97PTktKKe3sYAUtoke1waqQTPtfQoIwBM5GvwcBA07xuZYPvvmX3ZG2ZcUGmczz
5x/HCWPbhRCRSd8d/Qsrj+Alske0S0ZDbMt72crbf8v8jpuGhRjxFA/G7VUfQyMZugAuEMKglx7L
kzVamVmsfwzc/SUbZKTNVlodwo4YPX5M7J3lNeCn9Sx6KZs/3hFlfRMbtg6j7oMC2P3EWXyn5xjO
Z+FsCxOGEJbyVAvipRLKnd+LT0byrTbLI28/e7Yp5Nd/pkL1MF4eURMuJy03dWmn7mH71M6g1PhV
C9RjED4/MCGS0C7G1Duz5lkOoJhkrKIIoLhzibgxPHWFTRJVgmBUGENKq1yxE/DuvmfIl54lK7Wc
43+4MsAuaFskyknRFc1ZSayEzGFiSpGsMtxbReiiSO0F+pu3Pb+ph4Hed7bVFlWT95QZ2fKAwHJC
30j0gsaCHpAuvJ4nxFrzEuNhRMTAYr4s2rKhXPn4znLXrYuDmuS1AsjJSrzX9qjErJ4gZ86Av+Ew
WO+WBPEscwyRrB13eP8QPDYSHYhrvbrYWdmBoYD5fta5LCCm9TCurMyAOqduhJhZgjYEVapYNZcS
cUDoinWkTnk4MxaAteOm2dEPdmh+7bk7f3pPaviUj4eY6gCFTswBrcNqzFDDDVVLBVANiyEZELTE
2Oo4gwF65ciKV043je4S9ae4vG6ZfiQdvlffpY2WhW5/XX1EzwyRXfMb9sExkwddYbVbWuB8hevh
F5kqZ24792ZY2JTyVaGclaXEq0KXxCSJ7/NvY8R1XXQNB9aHHJR9ZlYGvHLXLbM31B+33l4rquT1
hB6PZP/jizoUzDhS5AmvVBn6OaWPNInLJmJS2xkVMoRcZvM7kdwhTX2pQXGc3BUBsMgPYq7RPC0R
klOSEJKInP0Y7opVw8noP/9Mux+BIiO8goL+36PoWrEqk0Qo3+EuerkBZMGwSzYgg2cypL4Q8sjM
+Dv1qrBotMbZfOgCZtElN02O1iJ8t/pW/Xma4bCpf2byZ/lgXfHr86zcN0eEF9LfJStZ37//RqOW
Nz6QuWzPLyPv7aXPAIRitv6T5wY297aRpKtJHPc8LXS3epDRW0Jniub3rkT7N4gq19nmG6Zbc0QU
CQ5cNXE6uWUgg1uL1+pPw164bZX/q6I0vuidUZ9ouA0Q6fy1l2DlT+gE89Ae7dm02wWVZlq27Rys
maRbBVJHRe1rrXPr1Tw0D0Fll6mjc6eHuELrXeURQbDIPE3NoBUSTp+avAK/rMp9hkCI+gi5ekCo
aqZvxokZBpKWiDKZwrztgEYq72bPxmMfy6lftWjKS6iOWmm7Y5w5opaFB92deAVvrcUy5WMzBAhv
ceBe5jxKzwrN16E7yQjMrbuhFbnh3/NzrW+MHqB93s7zvM/8wd6FQthsF3b185T86steTSl2T+3R
bwgUpoZbhNHxU1yiV1RjbylpLoxbJYyVUJQP+LbEpmuleQS1LbsbxJ5y9pp8eojflK6XImjeOdB7
/TdcL65ZEWUHuQq6L6YvzN1IK6jb8auMvFBvPsF/5kmYDGcxwZI+xCXAUVa0wBOkArz2YidyuVgY
k5VBbhSLzZDiA4ui30pClblNDto5WYfBXNnNPjOoWZ1MQbPliSMexKqPnRdo+IRIn/+GFfqFeEys
dlfkGBuS1i/WxEK3NISlSNFsbTsA11y93BI+SffsHjDRUNmP12n0IM2XG3uBso1JK6+LUeOqG4tz
atA+YOEUNODo+dlY+bm/r3DX3juWEMMF+TqAd//Pq8lPfnMo/KfhYcXvU4uPWjn8haHgUCUA09aL
9gA2t8deTQrXRJ7oMzVtj5IUA4a+D7S+z5YmUifYeZcMpP5dLiQWeG3uJZ/TOxfHV15H6OkQSJOT
yMMGwUOf3zNGzitHABXrFvGqtALAZdF6RTItUwKq2Q2REcAQLbJvPomSQDFT7m5QK939j1HIr9is
SPI0cuxjN9UVY7x6dOdul0vkDYpi3UrcJzRlL9AYKfLAm3Macdw80A+p9FxLsisytTUbLtanO3Cf
uDyc7uMi0et5ZiJcbnrAu6CuhBhBFgXb19OiCE2nQHhrTSNzyxV5Q/tP6G0UwltvpAJa0nhGNoOZ
SJ5AT2IvI+lKWJ0oPAPLYLrk/+UXUjrDqE3A1otZwMkSKsLrQNR4wMDwgCQA3J47HDBnGo4cke3z
DvKVUNkJmHsLR3LU2cCtQ63pzTLDvRRDtxdKzUgBrtGDQPEO3ACzcQl2AN8fhXhqtbD/5dp+8H11
TCQfAWUNVpve/cybcYDwcADB57GUVz/3sGIlZKWEQAmc3Sjge73ft9O1Cp7H1Bwq+Dm9RO2ac+uD
BN1wbW5FBS7Cf9YvNmHD+iVquYdYe9QxniH1Irut96DiSC16VX13nckUMYE9oaGd7uWuTQERGZst
gYc660GaxqFMA8YwSt5vKMeoQnAA47kfcpeyw1TSQ6+YLCSF0z3z7bRmFd3DsaSwzac2x2D3dL6S
8cbXu0zxpQ9cRey5qaY5s1Sos8vcpUsOGcqpy9Wnokx7QeSrCjTIAmKdmCz/ne+Czntlcw70MV4q
2rs1tJuvDrc9HNU+AMUleyykXIa1yI+VFjdkRpZS8k39tzXD5yGw1xbZILWYN/lyPYGC7tBY3XtK
Ey7wuTKQUxXoDsQbGcFhJlx16OcwnA/7uxzRF9MTtvTV9nXI4CvDw0I1nYB8w7sAVC6DX2rzYuJP
0q2LAaUOGW4W48J7RBu1Vwo+qTXox5+QMQxRnngJVxdnY7PLLG/tCShAwYawY5MmEdItcMBuCPJk
2a4e0Fgg6UsvTUfrtXiRpip4o9Z5XrDNaEGdxdTkj9SPDnnb/zn8FEUeT6GgTTpZyvtvHIMOaR4+
u7d+j9rijsyiFNILHG+tDJf6K3rtFhvacoetg1OEP6RXsdSppIr5QqzgPtrfRLfqP6Wj/1f6sbwI
ScG/RZYoSvQU43F3s0hIOaHfkiVLsSHtWR9p7kLa+vtCmCFhDmXtFC39zmZA9w1rc1krHT6Y5b96
rcpAuJaz7VIAyoUS7pguzAUhVntwpcTL/0xhcUWcXvBx9nnKOmxhd8eiofADDtew4cz7aG5FFOm9
0ug0V07PWY8DNb23eKmPZUU+TlKAgqTZ3i5V4s06JzR4FA4m8CtYA51r4JfF4Fy16W5S4c0rgGN+
OdtqPZQTdepBK5UPEJ9CVanwd1Z+ty7MPhdMFFWtFF5DJmdnPOjczMzaAB4v8WFfXCehn+bEotVq
YKtcioVhrT25o+9ZLkDSBadRrNt2a9ibQ9djO6IjCl4owwi7Q0mDTyXE95dfJ3mXLTHaJAe+MtuC
1QTGKFQC/kX/fN+iV46Z9yFYDiS9mQz4LDr/WUCS75z6ZHMVjXiobiEw0dg+jgSwmpBnvxERIvpd
zKuzR/MW9ZiA9b3HG8weTKcENO7ITfL7aLLRWCPeqCmbNKjjV742WhwflRQvEhBGv7INh7SMXrXm
tCgmLXsxUE6DsaaVJOxBpBzztibZ87I9HY7/mYnbymFeefsYgkk9yZPe0rOrKvogoKFz0ylHvZEe
jlhVmTd1ApldcLyXroXX2seCenQUb0x3NESu8RZO+dZMnxybY1uH4JwOrQVSnuPHCYGFrHXrEz6/
o3F0I37+nCUhX099SIK8TW1X6axEGYCpK7iJtjWULEquYR2nnFJ2JAtRECESZ+j4jW45ltUbqX13
KIV7pFBeQmDzI+V88P48RgnUvhXfEpC5xOSfP2WyZdgoQwIBGCzXdVS6Vg/BQ9Z5//XOkHJPdYiE
XTisVKGjQDHULh9UJg5ZcD3Na7jz+GfLDmjCH7wN/Ftmn+5XMop0flM5pNmp6zdulhCgdfIH+svY
3N7ugk/w8pWAgMyPRm/2j3j4He6BjVQaSO8Ij07+/ODltoQvikRbk5lEvaqxlMTHV9UxAK3l3oix
EYq/a8wrlFOqFh+NkRAfp95wZlM9WQaFfv6+WI6psEvf00dsFsbiS82JsgOL2y7A/LsOeGfUxsWf
c5OWVlOjng5EBQ6aJy/s1lm+DsCXxxEiVHC5csUT2TxI69igwvGjAU0JKxLybBZ0i8CYYT/7fBfz
A+3tpks61IGE2LHlReBSwnmkvV/Xb0yYxv3+s5P0DJ883vS+1O2HZLQNP53iDaZ+7ewES6ob3bQq
7WC8SRaEAvBAR0NBwIytwvhx+Xt+QfyBSbv1GUVMyQJxgxCnAW+lAQ1JTMRw2vKnrP+1ptOcKNfd
qzBC0rb8fchivLnVnw8JwgTE9qTpmWNfNndpcnuJbXKae2AwDwZz+0ytiYSdz3QqwOtJZwA7a7g/
VSC9FNEKUkHaKHLGv4qiXZwC1KDpoR8hspF3GZP2SjpdUM0TLPaaRsRyAihK1q+0CBMjzIDfP1KY
0SkHFtzBN34+eD2g9rquSscHCxjz2P7SY1kLKbmX+4krfvbiZQyGVKGDOn78TNYrOwpfmVBUZACr
jaE32dIPqz7EkIBzTTO9+tyDLZXQKdmfwTZNhDsy3zqmTL+xzeeVA+p6VUmBHSzSNYpl2cM3ije7
48KV0LsZOqftmFeF0jRZuqw/Y73oel49VH53Kd5G2u9qgnODl0Ei85gDMvopnNJK0q7bKWgwvam9
41701NfrQQ7YG9BDbWXpESdET9Q1N7MdkVNDzVdbM8vP0UllBBM+V2gzUbXwQdv2KmrmKejx9nW/
7Flmeu1utRpNgBypYH30c+J0ov360LNm1KjGSmlEfl72nCHy8HjXb0ylY5nuHckjLvkAvx8oLg3t
gJKh7K1/UK92E/qnViqpgDDjMRoICH+iXwOlqvpnWYGpcu89noTxq6m3A2Guc53kWbc8jJCyuXkd
KZOja7Ozrl136RAtgokI1/R08Wt/BB76M7Nz0KT8xSYEqhyJN4YxeH5mnlhmjwZ0htGxhyCrjJmF
d5L9bzCwIauTA2/kSnQE+No1c0pghoaykqPZ017Vto16nnkeqTYNtq9Cg0zFZUXLdTG4WFvDdO0P
6x6577pqMwMwcdFYdWQYJnDwfMNKHn49aDG5Nd/KQpG0p8TY3Ihhzp4gJnl5jTKGalmCLB9ELjgK
Oouf4O+yTQWwITNxZe/gm+Rm1waNZvTVzWdxd5Pm90tk88Srp59LHikU7q8X4N4rM9dci5S2guKi
I8XnquCtGO3isUL89LEw2D0wNeP0KYarnjKWiqbR2jEobMDlhoEq2GmH+Nh0uxtghLVzgGxHOn5l
8x7LHEr0W6+WncrVPD8zEt329DBB1VSLHw2VQ9x0wnZ31PVCVwmfZwIBbCmb2K2ZFd+OOYjDWvRA
Mma6c6l/wCnwiGR7TRk8+mdE41ZygQM5UNSmwD8s10xnvMUYbYTbX7YrHpsro5xDXmsZkfcRHGdG
4Z3I7oFiKBvLWXs1NxYbqw/+fxFZx90kaqDK9We7nCn8uBMWN7ouzu+GvsYpeHUgdlQdT/wu8/Dj
xp1C3BqYL/UzVwzpVjmR2r2eitOvFE3XXFJyrpGkQptbuwBXx1/PYnThvBWLdJ+oqQp3T4oQBCsz
sHUCfj8uow2xtl36iCoGozh/Rbp2tP/7c8n5uUuJaxiq2EhdH+aZyOpn3g6iSyosQCA66QDFEwpR
2orwnQqtV2wF6I6MtR4dz9s/bFysoTqDduYb5oK7wU2/EgnWcq7QDRZZFed7NOwAs63jp+0vlJR3
aIOXA+1OIfO6Z5awqsRuQf2O/nkebPUuQAznVtosof1u874GTevthNogKo0Q7teXo6B1XiBiMMIp
r5nsZhes+MaMCcF/yhKP6JL+5wvURb0EP0h5u7xJuk310BecO5QVxb/J2SNHl19dghaQOI+cybkY
T0rhTgcZy/BLCNuXPo7mlsLW6IMHT9feyXMQSUhM9IeeHNbblYZ7eXYS89Ya2Z3b8BdThguZ6Nsz
0ehywbiivPa9cSlL8Z2z0RFodSqyqcSebrcD/ikkHJHVlx04wym00YYCE7vUTrP0GR30hzK9lxCz
BCKEsKZlYuiQCQ+3WUWBu/yv2Kv4rAJ7qPXZ265tmN8pL84vCgmh8qKtZhCiC4DReP9GM+YIersT
xOnNtfXP+nU4d8V92vD8ODBihqJht33kGo3VOHSWw1mihR8cC8vUMk4ZMS7xjMeU28qvBA9gDW7R
WgRSW8jqtxb9sIANL9Rz54I+yujFGSMP+U2x+g9RGQ8h3mxAZxu4QeyutVPFBgd3ZjMXn9oWZ8NY
L8+8FWjXRVURDGSX5Taxz6dY9zCSTujk/J2b7KQgqpZSJ/JBIYTAp3HAqCAzU75fFUW2wQHy3bJc
o2dwHpSeXeLuPdYWFfH1qAxfTJienLJzZ1s6M+EgAoXj8U9T1sp5USFDFmhu/N2MdMIOK2jzuh6X
IkHk2wwTGoCr+r0OfiYXuRUfyLZbhOm3eTcnIfPvKN38baoFlIKmg4sEX4mlYq/KUkEctegSzGpH
sLixYXQ3wRjsksHT8CAp+E3sPe9vh1eFA4nBMpFRgRDnWt3dDiytrj62ozH7mFYqsH4AZgjauAjo
U9KmIUhUSQDFd+MhWig7Y+NB/mtzRhMlN/E94Q25eu5q/Rjvnk/GKeEN6dagxtgWw66ecS2154GG
CuAqxAzIs4gcqbUUma7mrk2j/qwBBS1HbQoTjgKfA0IFx26y6VoIzPInfdGQcudWIJmc7bjOL8/S
6GNCCxh0kvZ4AC26CihCJu+mznqE9gNW4BtfrvXJ8KYRjz11myZCG77kcZTYs7OdvNV4wr3pqKC0
R84vE6ImP/URpQQDZvrnQzjVb2eyJod/asfjPs8pes2bfxhVtDYqXXikfKvMO3ksmjBtATe+Kgpt
mevFPeQ4k7cLTvTvpk+Gb2RAeyMs9l/vLGj7jsKeUlmf1EyjqntZwuPcW/gxBD/hYlNryDVOFUly
4iXM6JXKi/4COy4QwmqT/2v5l7p9bEl8LdKptGPjfblyawBed1MO/FrxHbdXwpTtxlKk8fiPh9FS
BYm20dKwWaipqi4TKfskwVRjG9RPJtuu1BFdM2kHi61DKkeb+GWD9OeieYzxyu+ATUwbOgg+JDyM
c22m3Hs16Wpyt33VuiEaglCH4z71G8xQoIRQ7en8oh1OBOXr2hjBqBAiqoXnX8YW1hzRdLJMe6su
4qOBt4Kuk1EhsKs8TT/+PuipG2h7Lhz+Plbi1recjAbNcBi12baTAo6cT7JVWs0pUf+7XKhJuoCN
uD+QkUDHb62hMBw0VTO0SCh6A5d1uxB1UIfUu7PZ7QGN2iikqys4imj5GN90TOlGaaZQuWyK6UmW
aWf86Eiv2y8cHjvqJeXfucLqtKAZVJjmG6rHPj3O6lI1RrTTVKwrNQlTTplVyWC5RymMrvlAnGB6
RDAA9sYeSjPhFCj2tVrX+2dfxmNk9VkdjeX0l4CD/U7r1LhOXoHJhpQZenZa/it8VLHk76vDWh5p
Qap0NuwW9U7T3gVss6PlnV6+MpgfO6lm2JPdFkwX/Pbd6c3uIr6QyNyoYhxjmtERSdlADnDIEr7u
G9CAo00fsTjoDRzHBVYTyytuv9rP9eTwfxveMZaxGOvfMiVebt6DYkEYLn6+/LWBxpq3EeC9+TVb
n5JzMtNXR4joaQxms36iIXuGVlQN0fMDaY1icDkW1O7rc1x9JUJ4ECnC6IPfYvTNOCa6wXrHwXcK
DE+mvrp5Wb/VmNcV6lI6JG3KftKaECcl/+dmRyOLhyMV0gaE4JiwlB94Ma0+YZjpN4OunaTV1KYV
BewpWGBK55exE/Ag0LIACv/q2HxOk4NklmtnDLqc5id4wRBELVOjhipBA/Gn2swrZ3DWPYykbPOK
rMpV9doowlLtzz3G/gy7ukZaC7Itqs3jYgQH2pMcqiTE1Lhv/7urJTx5NPaF0w1fxBzVJVDFAvU1
fEMyGc4gl7+rYUoSw5oWFt5YP2JSpvPNxc1eTtxw8m9dKCzY/XbYGxfCXo2OjIyezOFSDl4T8KiP
fGAoVfWYvnKhjNzgZnkN9uQoQwWev1AXvE7D4qPiH4ABmJja/vo7WNRW/4o1BzrBRS0Mld3p3EHO
nltdy8Gf9VDVE3eWCiDuJt3+I6bgbYoUt2sT9aKsnax+so9L82+4pM7NziyyzcuENCUOUMfkUbCx
74BJaZEkNJASlVGGFydEaHO2HulLwRycx+svkieROaXeqPGVQBGWkwYK72Mnn1DshZjGYS4i6Wr2
ZS9KEwyTs8CwswE9ittw5NkGGv8pZvyWda2XosjQAuL78UiNjLIXKYQ/RpvImSq/CaXFuBXhPyya
5BzOm3c99vuxlkTyPQEQUMu7clMinjmuK6WIUMjPuR8iD+CPxevJcoozwEjtcZUqpc/vgeGtYsPv
/O3rol4cqSv4uXwSp/LNT4xp9Zz7HHGdlgoVNQuo/vfRjj3uWuZglW2UEfY836oijvefNQoOdJdw
mSHYtX1nSQ3GuXcGQntND5qlvxUSVYGLJSass3TjByHikwcRYQcT+i3MpV3dIUHWNZ7N+JD7TKbB
7HiOhjcUhXdWHZhK5oNLeqRKlKC6XOrla8ROop04B1K6ZdVHDMEMvANCy03sVV3FxoT3DISIW3i2
aFJASQQhPuOOLF088wUCTsI6KfhEqiMg8SyBxnGV56N2zJ+EtHEN7xKMhLygopF5XtgK7X8Ae9ru
H0IczjTtu+h8XmjvhRekdIHcg0PS/bMV0XCXNmjykILAgYCJwxcfUkrCIZhSgTX7kpTqh925S7/z
9JT8pMuWScRkVnKcgSyE2aAVBLpe01XgwIJh+b/pYNN8iPlJwuUeMZ0uYqd3+5sWQf/4t55/Bkw7
pUPa43DFaisWYa1BccUDq22zjUid1Ivr94gmQsJ9lB6Tkjx5IX9YuIDnulN+z9Rlinx5x/KFyUmD
6r54AIzKFddhhT+hYx/z1iprGY3MdGRctb8Jwo3DxMDtYSMFngJYkbYV7pwjPfyoROJA5iWFOj9k
oP4ftOiqnh9NPTAlEOEBIJHgX7CyWTJp1JWSykbKkrzKDQXe61M4DqPqxt1IuL4tv1Noh0HM2Wzf
CegrE9eDpMELenmSJy+Jo1SN6Rag1mSo0f9NnhQoGSuf5wpILzG97g==
`protect end_protected

