----------------------------------------
-- Function    : Code Gray counter.
-- Coder       : Alex Claros F.
-- Date        : 15/May/2005.
-- Translator  : Alexander H Pham (VHDL)
----------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_unsigned.all;
    use ieee.std_logic_arith.all;
    
entity GrayCounter is
    generic (
      COUNTER_WIDTH :integer := 4
    );
    port (                                  --'Gray' code count output.
      GrayCount_out   :out std_logic_vector (COUNTER_WIDTH-1 downto 0) := (others => '0');
      -- "NEXT" Binary Counter Out
      BinaryCount_out :out std_logic_vector (COUNTER_WIDTH-1 downto 0) := (others => '0');
      Enable_in       :in  std_logic;       -- Count enable.
      Clear_in        :in  std_logic;       -- Count reset.
      clk             :in  std_logic        -- Input clock
    );  
end entity;

architecture rtl of GrayCounter is
  signal BinaryCount :std_logic_vector (COUNTER_WIDTH-1 downto 0) := conv_std_logic_vector(0, COUNTER_WIDTH);
begin
  BinaryCount_out <= BinaryCount; 
  process (clk, Clear_in)
  begin
    if (Clear_in = '1') then
      --Gray count begins @ '1' with
      BinaryCount   <= conv_std_logic_vector(1, COUNTER_WIDTH);  
      GrayCount_out <= (others=>'0');
      
    elsif (clk'event and clk='1') then
      -- first 'Enable_in'.
      if (Enable_in = '1') then
        BinaryCount   <= BinaryCount + 1;
        GrayCount_out <= (BinaryCount(COUNTER_WIDTH-1) & 
                          (BinaryCount(COUNTER_WIDTH-2 downto 0) xor 
                           BinaryCount(COUNTER_WIDTH-1 downto 1)));
      end if;
    end if;
  end process;
  
end architecture;
