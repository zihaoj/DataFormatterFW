

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jYEZatDrXxapAXuMBTg/UWen3fw9jH45wq+s04qxsak0WEGzBxSyb6CIxWcWLXx0JgeRI50HAoCo
tkKKEVDASQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SIOOEYVCKgG11SLLhdXp668sIPddZmNOgZFYpDX1iRfAqjtSSdEYMs3iW36jQWf5T5v+mnILJApM
pP4HL79Q5Bh9LkNjwP2GSncUOsALh7pc8gWmOQHZSw/f9pmftP3mAm9twPOxP6A1egdfZEZHJs0n
mD8llCgwn11hCYBUnig=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LSxtq8m7OmwpRDVxs5DpH90NKe7PcjaeDXsx5fQqpXSvCD3GRJMhU8Eqc0Qi0crbUVks5Cg1PTWJ
0NWo62DU3UhWp7ZkZzsj/JaVQxQwnbukXO6thWrbM2I3dxpnDNHRzTTitw+pQqnyaIIRsiXDXboM
W0g6TOHskmIlxJXyf5TqrlhNafKtnFW2BK0cK7TBaQ85larBVGG63Rdnf61fJZoWOSLcXbcahFXe
JrROaYp3ssF6CtMpG+4ZHzZ8Ph5VkQTA6DUUD/7UOgXC7t9/4lp5So4Vaqh2z+SkN0/GBJK88BfF
qxS8L/brjv+61HOXByAPpYGYapkfFX3c2rD4ow==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PZ/qvWcxY9GbmjOQp0w4O8xSrXV5xKA9em5mXbDxw7OMeSQGVF9gpXYRVEeBoyZzxBKhrCyTOTEC
dIwV95XdkYGXJqzQ2MhOSaTFXDtSMNEfE8u0WZaNZQZZ62QHXXh48JvPuKmNBG0Q1EnjlV8DMcIn
3z9KAwodqvcqznN/E0Y=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tzN5RxGBWtX1dcXTSKGBOQHwqUOAsviw1vUeHmfTF5k5j8QHHWWjNV7A4WYfETJCpDW5Su5xT14M
mUf3cAClMcIKTGw5PShQPe4Nov9KELTWXkZkWaGIRzzmhYy7IaOe8p1ydIRHnMHHAW13mo8epZ7h
36ccAaKnj644h5sbPKSar5AKPnqHmTQDJ1oqobcB5UghNvkD/XdGqh2eKTZI8eNZ5vQRfMCLNGhC
cBRQNL0VlmEHz47k2EKkMUA1mxkd3z2MOtN3Fh73/OcpXGNo28W/h6wxzxAhB+bHSnMSd+XqLnKb
IDDWKvJpoQOfcfuV1DbeZfvhb9hqQzX2ubFu7g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8032)
`protect data_block
kZGZVVpMXaWUV1b5afWUeY92wxjrbOA/01f47CbxEpvwfTfc06qQFT9NhgMpptcuVewuUm1SY4I/
Y2GyerT5RT9L60MU+PmELMnP0jgjvW4hXH9bSA/ieLTxggvSzK6sZqFDw1mKA5ULecg1Ms98a2jE
NCp/GhYAPFdXyryDyuh1tX4T0pxi+6OpCUI1XiXdya/I6fZkpgPMGHu333Cx1V8kBKcq9Y4dYjfO
PzM/qcGY3IkLLKDXMdyVzMo5Iukl3uS6IGInOjfKGzKpSu1Ibcq6wS28VfrE2YDckmYf91asXOLP
Dym73lpD5bkVFi9R6+DQn99bk1N/JlDF6v1FVaZfGWnBRJ1biZztbSmbrTukMyxLCQNQcPRUbGWC
MUzgzJxZ/fEbFzhS96UTdRRnHgGIrJNho3K9Borwk8Qtmt6+KMaYcG5yz79pnyGSE/nUrG4ROhWz
LA6SckwNfv1Us/JRD1JLLZ8sjk2waMUT2nB4Gsf+j3ZQv+yw1Y70Z3P1pA7jq2kDfPClB7iIHDrj
gi7khWw4D6lNTrm/wwupIQETbmgps3bVXUpyUKWBW4EfLl3VabuZky7gY/wjUyyrS5rBcgjC1Fvu
I36gerBIF1gR0KeWlfTN+4FvrMBnOy5gVS5J+eDdO0ev9QR3MiFLbbSYVJ7aQkeStn0JHUQYILwo
Z97yjcrAnJE6DtXMXar4EnCw1cY3iksY25A/fYn9ZrwMFixRDCvvA88eXMz1zDifvZ8vtCOglQEI
HKKRhwmgS8FHj/OrP1YUMZCltPKWk0ZEbKxkGZmuUtmfxubVMx9MvoheBSwhnVdefOryRhK4IyGK
xKcqC33KBjEEZUUd54W8jV++sfIHGiZK/7qOO/RbwR7EVuWJkqtperaSgv+f0+PJhlo6QMpDrtMy
qfNzybM6BNdHQX61igXTHWXbmnUd7+E8ZJutfRIuWYSxqmjYUbt3xrU/fwcrf8scPNvsZ2SUcCMH
HjNbfVLsDyQM/XnMXtVfRr9I98aeof1JfFDcPbxjUwgJ8mTR88gl31vQJFhM2LYf8l2pCj4chaqI
IVM4VfdQhWr9BBrTagLdGy5WvNkcWWK1DBl3x2fBtp8AwBuDaUNb6Xhxi7+Q1DkdK/qlsZrADoll
ik8YAEJEY6d50oePNKRj/F4f7iWQEQbs+cG435wTJGoaSlvFQhIrjD6V7cAvMls0Rgd21C4ahxVX
w4soW1ymOclTQEg6wAYOn8fyIZaU/+yFecGn40QCye3mR4zS7RFimNUj9IWmwuRC93z8w6WSy4cg
7qxNcd3mizYgp0/Vc87wB9f1k5xGV3SCcQjEXuJnMg5zZ2uttd49FrhnDJmNZQa6UscJ9SOnl2k0
S9bQZVu+mIOzgtkBKhacUUTRUUQR301/0XSJWQM8pdImGz71ZfANTo8qD3omAinsT+DCHbp8xxGm
QUmfsLLcXjxpRZaHCWxxCou0OgVJdEsA48ptqL37f/B6eWYmKb8Uoi94j+NiTnHfzDDR/VzRRvfL
OlYaUMlOEDrq06WoSiOK75g7iJB66LUEIuL/IkY9GlOrhLXfAxwt6o01Ahr4fiFoKCyFMnmUr6Y3
4NDvPD5NX2RT1pMef3F03MWIXcOS+rohZoInR23Nd9hk+vDB88e4YQPQ7ZWKHx0TH2S9oMF51MMw
9ZnfYBSd4rzGN1O/BCBURCMAww80y3jElFp0cGgfS5VOCOt30XTNFQKXR7O0oa7KMJN3+c0ptMLw
pnJEAOBjtOi59Q6zb9VpR2szRuqu+phjKtRINyExO/iHVtvgp/9BOKrJ3OBXyp09Ip5LUxdMVT5y
bmXxWxRcWA+eaTkQDKyTyJCLcdPvAwraUWmq4Qx4I3k1YOd5D8RPDbTi+HOnTIfjm/29F1Ewwx1C
bZl5HEOzK6wMIon8WhTIhp/EVRNSfSoc29YuuJGjHckXOgb1rrTD/8dUI/EoRmfnfsJLAuKkEQzj
CtPopdxafVEVr0FKZG/GhypaDEAcpbtCtUadqOwtXsj1LnCVImIcqsWaZ2t0xYmusO/qu+u7IWOX
VKUpwGXhGqt06xFbdfoIKZ7oxeR5WGBMKhjPcqs1bhoxREau941kuS7MJ3n9+hOiM1O7tNcHYFWs
qE7hjE170a9nXOhkpapD/Yi0LEN4imYzg+HeG7MqGanSvKcfyjcC/1GfCjPxW+ANnatJErCPUbdP
4m8ngBVXV8yAS255YwVZpN1AVZ0w6JQIrgY9FCKqK0wzu3cJGPEyWm0r3LARDCz5xOlCN3ji28Il
hjisSs4nEx/qAmKP2HK9GpXnPQix++5mzJeEeH72SYHsWG9M9yaVwKtH8KcXTSXkf6sVsyE/C0wO
Opz8x3uoWAiX+XmqeobDeH/VZ/w5MPWbxTQPAVubRpkGfHGOl8rOBVxZ91pPDzuFsp7nI0adAF9X
ae+Rrbej2Yg+4XktbE4obhS5fY++ZRlNogt1CeGPOM90+bqOUlwpu02o+u/1hibnPgjLyc79BZft
2u2BRHcYiRSJ2pkQuksbayvqBQEu57/cjj2wkMz+UHoAiEzKh/A/7PRSVQP/dpJxHnEXEN6oVp1u
2Y0wynz+9UHAMgCMz6z9M0nb5XSuqrIL7Y9qEIcRRmKNFBJEZLl8vnb2TsF8QwnvdH576bsWqxO4
j3rDnDW6RBynlh4FV7DAF4z8tSL4ArC1ei0FJvWmeodtHdTWu2yrurv10PVQRcmNmCv9wVJ1Wvfu
XghaFWwlyf5MZjZ3HN5C9gBQRFTp97X8Y18IJIirereH3p1VJ2FTZAzgIFz2CgfHGlCx3D6Z1zWH
lZdzxevYGuBo94rwl8J1p2c2OJ1EWeWIbwYocvEJpMX4Xk4BatqGnmQ0o0JxZbPQgXmUlOft1NPA
JnaY5NtSK0eS0Sn1ry6vvRE1HU+TnIqdt40aYsfxTvZC4bgP0ryfan78Eia1nx4DMmGAG9VIW2NK
nPJVMASLSB3BsCobxZUDyUX25aXuoqrV6vV5k4Tk2wxrKYXnOEMEnHvGTwE5olkZ+BWDLeDfrjPA
YNsG0TCuA7Il/HWGcAnQGWXNhgwA+3TkMtcdTnVIwELv3/Cca7iDSaW/+NPtTRTyyuxMJNrWWjLv
CF0wiWjGX7hK0NdIIHqJgONxoYs2Lq/jIZoKfKIPepTRTiSUingdiRc2Csi5Ud6viQydUwe9nN1m
4jRbG7R9rSaArJXOg2FX5rIxNMMptVPM8+Sgq3P1oixdHcKELSb4SdwSsp0/OnajVVyaikr65gIJ
M/5buyLxHoSN0UxYwrWXbFmqrSNNSzZDDCglpf7/6m3doxka/NO8qYU9toTyVVdQCUwNpzyuCPij
DBZacbpAHMLm1Zq4r1DTJwBCucfXPAMWKAZjd8/JRsMgI+fRCdg0VtD5wiHYQNOFCVaXMWeTHYYL
c7a1mfYBVkJRz9eZ2y19f5AwWeKGb3MxE8soCM5sGFi+lpUJbgldtdOEkeXJ3iC+K9mGvwtYgKkY
1nT0jZ92bubafAVYPW5tFSf2/2Bb3xFFUgGOWl/IqgLjIxXHGIdUOJMzJV4t272rxwhtftNbbLMu
r80f6RT+xT9dpp3ou2uBXtWqtYdUJJRvzP+pADWIr6Dk7EbQPwdal7sdUiwbY2rJu+nO6QV5O+7o
JoKU0kFmpwaQHdSlOU0uweS21iY5I0hUMBbLnBdVH56HE5xnaydw4DJh+zmvBOe1VFRmpmTtoewx
/N47SX1xhAXKwimpFIMOQ6o0C6T68sBKqUzmoxyUsEVddVvV7IBIjEfIfuEC99VPNPbDPmf9yLb+
ADx/G4fscjl4cp59Lny6eHiA0w9Tr/SANql90HYDUGDfN0f0gZl1g8hJFJxS+MsdCC7/z7iimQfk
hso+vezPZ1vWZx2bxgfzpo8zIUSHXlzL+ta5m0NOem7c3GrsPCZcd2KaPZZLf+UTLeFkGIvqr7BN
/2xy677wegzFdmRR5fQbXdR3dU4pDQV3TbRDtr37krbazJvYtsgyORsKi60kEC0DeWyW41QIjdsS
6IlTG04VfE4ZL3MCuHWRL+hbMJ97jT+w162f7WrPyLcqOq1TXiJnYIzPrYqsXyIuQpS4I654P9NM
csmcuXkMWcR6HqDUO2ZMRwa+sowoBL6tqN+wObhvgj5Dn13p3yNEQy2hF924DY3eUXkBfE9Lz2Rd
Y9J4Hcz7v2wbY53HEMW9I5E0m2nnVac14yFVUoY/xOYyshNHft3AvfFVuXX2sFvOGcK+4nUym6Sp
w1MBHGJoQDGk34aPwbH10APohJ9B6J7yl3XFneynzlv1TKS4xRnSfNmHWoCGMcyDRPt3fLyCRhx6
QpRdNrF4+y1WdfXsFlB125uDgAS09AU2k6N0RK5+QWbBbAfS+CO/QURV+k884uqiRpzuOKeanrvF
7evvhLMg77xyHlTJrQ2eSUs72ceYE7r/lhH2g41/MBETI6zWlj/4vcpQSWWaBdX63YTrh91DdJUr
OHU7W/coAlFGjeIuHQJ1v1V3v/IQ3JT3dGLr61O4UdqtlF7ytVj16n3+gdRDDKoY85NoPAbG+YlX
7WR9iTprfFKHvzlacrSTjrA9zoMLD7lYOETcTx41+hWL5tV05qyQmKtHdHENiEDzp++HKCA4UtE3
7RTA84vSNHQgYIMRfZgY3xhOicm87dj9EZGV8VYuR5gl6bvWSXhw4yyimoaRWMaqFJoN4cYtUfpa
EWJtix1SqHqRTgHRiN2mDWJplt3iuagPhBo6prpbg99kYo6gJaUCL6oxzMuqMQHHwEf5WopjqxyX
Dxa9XVjKq/qtGL7moj50B/4CFG0RTbh0mfcu79oGM9T+d8osQTHqCmQIuAEN/wTWcSpdklBXgpvB
otaXkTPUxuzIIe7Kx5mQcVDPUTz/F6WxD3K00paSiQrVQEzCVtzbGTxdwhizsdubv3nLpjoPnWKp
/NQIF/DIlisBZJ/o94gym/1mK/vKiBR3iHaoPGSS5ns34Mm1F4LOS7KFzUPg/ZGsZsDeOd+VFUxH
qsc8iLg9ETAerDKxPCLMzvDQP8KGbK/mjEpQNynlfoJqRbwbY7UviIg/GT5DSXvmU3GT3mW8vSin
6krCsHOmEje1AoLUVluj9KLHRZ5hbVBWaShXi/9kmpl49hyFwDVnDIC5BMAEyZVf3+XDwr+WbHoH
HNlhbdYhRDD+qU2pURdzbuIHegLQDv2A2h4AFTnpg4OXnFx3ZPD/dXRzEW88VNVTEPWNrnuxlM/V
poyaVr++JAJJbatmgqKjnL46rvfP9AkP01eJJ9niw30NBaUx3O+rhX67zWhWqYw2/jieSwHccezl
zwZYPEvAwlBIjKd03ovJ3ajy6x8AdaTtklKfb/HTTuoXuhqAav+fhGcD0UOpqTAGDS3gHojwfvpE
1tGvFZWeBgUNkJPwLQ7jmTFwCnXlcYxiGQ4YiVMFG1DBOiJ2VmY6Qb3fYBdE5rjyOgW0j9R68E8/
VzJD2D951DPh17qT6LTop3+rs9Km+z3OosCKkWTf4menrLwxpxYqKH6X22eS8DaIyo7ra6DD9aIm
U9+vp+cTr8jxgpxIrzPavbwkR+55wVfYwp2BMssYP8OAs7W1kW1h6KPFUKDtA9WT+41MBgo3p0IU
rlOgEQIvc3xt8HSL1md/cgNx8zjIR3Ws4R94LI/b7gm7kBNlonfYPLY3eJLHgL0Py78rGUpIqTT3
0Ef/AxdovFeYNJ5sfGcH25X/Y6n5WyCWT+sSWM+6lgPx2zgC697yomerTlTFkLySOxcKWQCOAJUS
0YHQWjVe/UZ1/UEVDX29Cu/3CK96NmUZMbfcABu7uuN3QnezyfCxrtzH3Eb17Lw8CIIldcwG+CaM
VZkilVMT2JNncRdUl6kGNP3iZ/gWgAo9y5ewNSu3pZHxKLHvnTtPLygvAgSZbTw5cNj+DJHDscl5
8/R173PjrbcvaQ8dJLXp+9JTnQmh8ykXqv9cBXlfuEd7rntAXEKxKjAn682/wIrhB2j7p6knmm9x
B60bttdlQEz/WXfb8YL0D/90dH23XsPSVFYoIPegaB00wfJc7KnV42k7ueuwSZGB36R8qqbOFIGF
x0T60/ATqKfGxYpW1UrX5thmhH3dwlaKAuJeJKcagsCtpBx4LkVNI8K86LLJ7rP4yrd6U+nCehk2
5CCjNlQGBJmn4mevupiYrtcr26nMTd568aQ0gJPQkpUCXaA7RHc3HZedAAxC7ROlx9bfjPLtfLAX
dMrBF+X2ILdKKSZizHZpHtm6N3kh+VuntdKAEx1offvd6bF9ENb5rFv8OVrRt5IayXCXep5mRlha
1/ovOcjX6C9V/yLuoUtH16flbGDA3O1BP5DmTfBtKa5IIi3Uj3cuADrJjDBQ8K4hrM18O4fAzliO
MTgJ9pA0AwOqYxXm1BDKNb39Z2eavNi0+U3jAU9EVmDSYURbnniewXKJu0j9n1d4NMxq0IlA2VSH
zT2cb8fQfECtW5AMIRDqXp2gc/O0BwRp7aKA9lv11xhV1qdaqLgDxR5gE17tP1GWiTMM7eanLT5B
lqrvt3qNhP1yZ0p5UsnvaraXGDD/5bb+edFjjSm/jO7ZmuP06Opbh1VY6OqEFhOdCMwnJP9Pyx57
vAbIOdpJuDO8HgfKddjI9LIiL/zhFEFrvbq21eSNnb684ZraApctH8aiGGsZAASSQHji1n8u6XLL
rDXNQYdmYStA3C7aqL1v9IMsROlm/oMbxZ6lwIlF8UJ7CTDpJq38jUYeQkpigbqymiXDFwqaFEmp
T7Ik+ISkqytGTen+ITyKAAvJkLsuTf2AmEriFTMHJlp1CSAq7r3+hoO/HtlnDGh/6Omq7Z2jqDlF
sTgN2h8pRwSO6prnT+ejFixxS/9LsMTx0OrYk6IKvAUCNXLEzEE7JxJR0pjeh7dUrRKdeXQj2t8a
lFDRZECuBaQTxsJSXlAQwfsuga0iLIY2bjKtYCH8kSfrAolnsWvPgj9+haF/xX3nBRG1zKS9LWW4
iaQGT7664BFb4FYy/UUMKKJWIZHUQiHOxTODXM9YyFJZMEY+22cnh01WHK6UDBcWt8Nbg5EpIDJN
//wVYErckzuyUf0YVveYmNIs/aefA6E/FwpAv3dAFWuT2wI26pkq4rHDreIgoz0fsROaxkkloE25
PpZW/R29DU2H71Xgi09f7MfkUvYQz5nTI8l/4cARraPrF5lhK5qiXE8PnQOn9irvGiJQbJQITO76
PSoTJADoMOwpiHqQHBGSw6Wx+udGLh7mwJdk8Q//6hnyw9oCQgES7m0J4GHaTjfyjW9pt6IiZO1m
EjexPuiRS8Xj6NztxKftmBMvfFqxP6V+hMh+/I/QRh+gQKX7nG7DQfyJOGCUM4dBWSbvuy6mdrls
oGPRzgmNudIbmU7rl3NO3aa/ycGN41Q/9igLOgp9BLlBXyIQETH30bPuXwvIFLm7DQTxG5W4CCS/
0Apj8rl6MhjoCvu7UM/1X6bpZmY329IlfIHspYzZz6cAbT3WH01I66lcK06ut52A+5A+/gC5NHwZ
IPu1reeojpEaxhHP3S5dxQoWOvXO/JftcLrssqo1E6YVbcpiqM7b75tyV64TsDkTWwiv7gWRd/x9
DvUmHSDzLeUmguHgzvqyCUPHXLuY2FaXRcv7kH5+6/ABZBP5FkzdB9RpldnCYPcNIfqUZZFc7j7V
Tlmo8+3qTOgOCBoND/zcSIFSsbceV+3pS8xEbDGlsS7B/2nztW8ON49JHUixSkLnd++kiQ0ZvXNB
vfHFylAo5S7qt1p7DmWQ3V6lCz3E1JQDFBsMHRG5AhukOYCxCsBq4aw5o5/Qdqxo+/SX8reOLnGp
mGldrANA+6/7S90vDB9KgEpUJat4TPxwiRW18vmwTiDv7JrvzQF2ypMPH3iPhHdAzG45Lx78NwCN
noDiBHFkcvi6sve/33M81V6taigqpsvL2sRUfbk0CzuEWwZk4vP8sEhtnOyrURbjirONMOlHU/Fh
S87fo4hUeWFdErpxzAbC9u4n3KwkGXymAbAwfdd1Cuxx2/+f1szIwJlr51j0KAkFewRR6CJTUGzw
bhh5YcvazrZaTbgS1u7x+NxCoxrxppSUG188Bv2oamqutVS7lRbfzyJLXLIsXzQ44I1scmbmgQxx
JrEMyHH8CN3NlgPtHyt8RCWBn/OeuuQcI1aB+qg0FlpDr47GoBiNEdkP7oU5dWDMWbX9yjx0x/aG
HN3Vaf73KY8SyBTpFJF6zJy1LGFeo5NjjGjQKRnMjDb/dtzFLB1pC2HFGTr6y9qAGUJ7gRLTtdFw
6HIoyFN8inNJnsxFnLP5jDwK5buYja4kCwSvLhbJwM82Rxaa7/YZzBIR83vPFpma6A5QVTEEwxph
0sKiq2AzY9kbUCnFAbBe+qa067tEvNsXC82Iv95iWyGvHp3XvbTvfz+VPyDV1JOuw5elTn6P1dlj
wdrFA2ff1UJn0EZvyghD37+l1AQiH1E5BMtEf1RIedJu5nb1hsuNXu5oT0C0K8PzPWiX1oimRKDM
471AMA3xc7418cXI8jGsIrBIjrR3/Ny3i4+qTxdeCdi5rQLVo1rAIHOEKspg2VF46O/0dYZ5eoeC
rOcEyq/oylFK9cLzFOwWF/eYMB40R1NHSDH+0ebznQCAVO9UV5uxY5MGJLWUPC/fgqbPXgdL1HhP
qbbUyNm8Anjm0x9FoJcuQzRHQV+90oZ/tXHAW6F9HFdkEoTdaxacjbUjosAnuuuR5FhQCKEF8fz4
d5UlxNYGJCDgLj39yeZZAMGpATwjjSFaRu7z/Zmzgo62IQ2qZQjtZbJvTLe6F0QF2/hYB6ifkMNL
E5WmAwu1kGVMfqd4Mw4sD4P23FxuCRHOGfEThD9PGRY+BK7wc/taOut3mbIa9y/438Qx5FScaGMz
412LIoVcq6qXtwWfvFkpDvTeazifFy0ua7KJuge9YQK4kPxtMzcSvfH92K544ek/xLY/9h0MYRqE
dBwSGeSJR5xwJgEGGhykISP37xF7QXSL5NUtrOj5mo1puc1prpwGTZhZfsTrYKFT7fzvbaXlaq1Y
Oqmn/DjTdqXBsB/YDjSWCDyXbnjiqcXrXmQaqp/VrI22TfUjPRsObHZwfj7AGYfgg5VwVIsiP+1H
M+Pp52nRD7SjcBelD5PZJdtqXxHlH/h1a1v92+FAhq3vwHEnFn2CLe2xdnX36MuBKfqURF4Lkm7S
P2HsOLi0wVeOQEVe/eJYDFcIwF6AmHtRDdaM3UXl/B6q2jWuLsx9qu2R02+xmPq72ETuyazzih6v
xBxBVmH7FJAU3+o3x+EA7I3Y+iwJlL7J2278EICU4Vo4tIvkw82l4uh+zcVTs30daBE+XsOzXEzi
stCK0YUGKWzzNyaY+ESlZT4Wjh92OQ0Fnh+CNn6Ld5NDRJMPkI0jzpNZTQmMbu2JdATLGpOlbLsr
sqx28hoOp+JneZSPzc9o6sw9qX/7Y7Z7gH//RyQxS6P2dwN2wwC+G7w/yjOvRGv/b24RI5mdK0UB
nNhq3Z6Q9KZXof0caIsFEDesiAW/811kZK0F14fsk3eV1nZFkmvISFvwmrOmj14nySLh7JElEDP1
/AMIglI9PRK9jedaoWMHJvmyUOir7MEGPsJHMFn00/Q1Pj6JHidgzLkHUINR0KAP+wlSlFDykTuI
Z8YfIstj3/b4HJufrTMht62rWq5J/Bsm2RI55BMUJaQOmHnb/ts1ScECo0VR5mSmRLVcuxM1x0Gs
ME9Qgyi/A/a+0G95FbXOtRKt4d7MmIn9AztmLcBhQevdOtJCAhr7b1AerliKOmVViK1YDSOLluf6
9+4Rd3CJRfcNvWDNcqsol2wR3lRxMOqeESwOgofA0RqMuBNUgKk+KdkHwMTwMrDb3Z6TwuiHiMbh
NrYpH1aEqrCXcW9QCVf5PMkxDB+ZoWqIEBq0wxXIlopgRca9xifAFcNYMDg6Hf9kvgoGwfD99If+
NbqMo1TWsf3f/H3TXfxofWHZbav9xzbwYUUYJohbToYWnigALe1sDyBCjH74unsDAVu5w6/E0uhW
fFZ5p9V+XIF7UWSmJl2hY+aOAWIlRdDu2RMSARKHmiMVB6+LB4ylt/XM3ikD+w5pOjZW/lqT/aVw
mKUUYNtY1g+qRaPfytX8Tavymhnuj5b9friSqMtOsJ/CUp37gU1YI0t9H+2QFY9/xZp/y1oyFoaJ
34Turl+SyHEqSLLp9PyoRjQAJzxfuYU5im2tVRFCsn9eorlhvo1Zgdg/WZplRP8aSEl/lD6vxM7O
kRARgBwDkNju6JKjG2rdKS/rmysYpIiyd6n53qIDYS29o/M458xOcyePTiip20gDM51DpaLDET7z
t3D8gxPWJJgRIo9yGt0FjBGreQB8QvB9DdkKEcjSTJ2P1ka8Wtvh5kD0Z5tpakeSeJ1+HQ6C9TZd
YUsSOWCZo/DpcBGQinHGgEXOblenGOqcXn+Uf7Algah429ty7lulv3rtk273FNM2NdJX4pMDsN+v
MKmsLwIvsSDAFanlyWDD6v6ENRb8G1uWFNv0LXb9DD9oGcHE9nxc4PeAsp20FocSCU3zr49NQz19
4l91BNwL92afGbgt5FmzhEwg/1Mqoh0eRA+MP58V4nBv/Ewat+Go5cdRFx2yjmT13uODkKXsUPQ2
uWUnGhlujSh7kLKVpc+b8YDbMJTId0+b1WCsP20Choa0pwb0I2QY6tQ14FVtguBUVFhMOg==
`protect end_protected

