

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ltvgyxLpfrd4CQIHx0i9yQRXWiWZKhyPIfPNAj8P4yUJEIwQ3SV/uvzt95X4UU6lqyC0DAwi340L
2tCOWMS6Jg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
T/ROy7I6+qrn90f/0VSFHATpTV/qSb4bOyDEvcFa/qIhfsNYeFqmPT1KffwuaURYYgZ+yDiLlUFI
4Z7nAU9FJk1GXym1zzfe8JukaEgRaYHwwgZ4issR7Ap/zYN+siEKRfemE5E5PUDBM7KPK7Tli/bA
gKHmoKYRFF2Uoli4Reo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kOD1AhfEB4MquvYQJaA5HyJ8eBHHXt9/F7U96GXIseGJqtjDpuJ+DOtLDP8/sjEbGhYXKKTFNOTQ
NNFMgeGiRlDeD9ZwOsodea4SmjEFks3wprFqGkyVGav9pK4dHfsK6WuXQKw5zXZaqRxK4f7u48sH
il0gJcoXmVhIJUDOGdf83ijpGz2SRgAbq9CncVgG4/WA8OrmPdqkWR2thQ4n7j4x0F8PrQVhUDXh
yXwRcmtYrX71FIvN7er9gtP/8mFL4XaIHJ535Qww71ITnS4SQmHYGr2tq41qfmofJZNMpJ4te1qu
edvC+kzK6Q+aMLN2vjHgTOstd4CX6ZpQMczvVA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wBt6RbjVFYZ9f1ocMvROAqtIqaxq1U5+W0Z+17vSBdx0TloEa9FdsxNfGWME0UnJu2Ww45HcBbRH
UxQ9r2iJKHQzqAnxqMqjum8PdXonJmIfDPFnmMiB1xmwOFgkKOVnjX1LYq5IjGe8nEwVXstSy/6J
o/r1mwB8IoWh9fCbQ3o=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lJwnyOWWv/v0sCf8I36Espi0gwPCo8wHG9LJ83oCkAVVGQ7f0zVbhcYTkm83iBK6l4C8uqAvxqmg
vB/q88T086S2K106Z7ne9/jH2w+Ukn//2naEOufSMjEdNmJhrECLRZSlMC2fCss3ZxX3PJYSxlyB
QZlbCtFVVT9x+mpuutBS/0IBrR+H57TQE0kgFE45W6f9vPLN4Qz8JthwGd/QoqwWQXwoamPg75Mv
j7G7MJtP15XzBsP+1f2gsKixeGMP+pkZ7GKhBZvXCXIskrT4kOBht+Nx+RUOOzu/Yi2omnCuU0oe
DFufeyUE4lCB2Ld8cBl7uF2A3/bBPxl79zjunw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4704)
`protect data_block
e0Wg8mTjVLvMAd2cIAtJGNjbGDY61km72V/O7wexmvB4kL77Ak13R/QAALXyA6ivVhuKzNl/Dbr4
yBrnb3Y+rT9oaUhhLMYfduri3Oo+t0xbUon68nnDncNquDvZonjxRXwEYE3OI/L6dMLsR6rY1GO2
/jfqDTARl3YIVDy/TR93EFPsmfDGW1xh8teFt59IMhgLIzh9u3sOc3eOnW012c/gJatzK01NMBad
zK2a9OFteq3g0qELkFueelmwLX+X6Mfggwjdw2oEIexdBQImY7/Z/Y30z9pPSIJy10j9rtTDwVcv
EqJfseQ+O9DicMHW2AQkLQxtFOShrREYDIE21W67E1G/ZXKcgJOQ41Y0evllr59SjH1JaOiYzy3y
FdmH+0Q0JFQjvTfHgmTZbbTJhu6sRPnpKcCf4vSdsovR4MDHeNo2WeZ5N3DVZHpJ9ZwPh6sI2ed/
aYMYhlz4+5aHUm9sQcUYzYLxJV7vjSzWTT4fFk1+yqd+XKi8ibqxNy5EHamGxv5lnt0y+oZ34fwG
HweCIscFZbQWsSJU3OKpIQlxRTUQ4wjsUbRgCNhMKZhxM8T0emN50Vl4pe3cFp0a+s1PRzaY/tX9
d37heWeNdMoKTul40PHRj+0Tj7wnDQU4+GYeAlcxLzqBkVl7V1jeAqu7EFK56kXX4sIHHZEZKxDJ
lrxIx78omfw5PaO0KE7AGQiUz66jRq4i2y8LRvuUN2734FQhIu728bR+gkRrO2rvbUrpIMd/7KVn
Etgqjnj342RYueOOK+VGR3aGrKo47SVk11WFnB0/bX4i/19AvWDch/lC6kQEneLhnezqc6RwhymG
yvNiX0tcCJwM1iuWqpDARP32xF+7N20S1jtQeJVMyeCMY9QUP69rOvThA/5TtFUFrqLanEoIwduq
cxGQ0loGIWyqoqmGMy5uzA5vTEOKeD0/mt4nA+Hacih33dHUQzNdtVdPuBVBsEne9dao1IGSHaet
VV7mpU/G9bNp5LF0YU5/trsFJ0Y84n0IEWAh+jj7n8CpitaOz8R6sg4yLAYTM6STKpeON1WpqhAs
1uF/hQ9wocMDJg8pHL8cUbjLYEsH1jUL5KHfRxHavYNEq1rhNV3mLrWlgoY3tQO36YQdVo8ZLxBh
YXimIzxRUi4OVe4gGQoOwIGQtQ+8CGj9w5xwQMtBOnk5tqKIKuQmYipNbWQJcjdhMSAl6t/p+CPt
CskFDH89mV4FeMiiKlf+J0xbTpALu++jbp0Kdn2elmWGttkb9/u/3UFpuWfwuDlP1L+xcfqZ6Oru
VUFUWzLPedNQ0qy99M8O/1hZtwTFCh2LjoEdbyWgNZxL7kJBKG3jTsnP9WQnUDVVf1LwhwoJUy0T
c7Zap4fWO/+2ckBzqxpK+pHRFCy1JuoZQYhpc5hS1Y8J526XpbweSPcwNavWuykAMiR8KCqwL3Fd
OwJUl7x45tTmO1z3m5/WU5qSZuJJrLJF3P8DFauWDrj1ri8rLoJUV4shuxoApEp0C75gFRothRh0
/pheTg1ZWWCsYMh5arPWysC+zSVzmKfgdC2LFUg40bBmetVWPE158c9QpOSzBrThzTPW54kRD4RD
+KT/pcQp59FrVlV3I6uQPR6l4AKaOyp1ebUh4BDUKGk946wLmYXVS/DKnDwsbwH1JffMweafsjBK
5YxyKpP2BTRHKaRvU0q2OsPOF3/3RqV4c6J0zsZEOHPPAXMZ527Q0dg3lex7KLTHN2RkPNpoTsas
TKEvt+XE9YgPeIX8JA2zroH4nK2pGjea4i0uBNFSxy/vCcYHky/bbNc/U2qAleijED7GWEug3QQZ
H6Qt0QCuqj1GqOI5T17A7buvOTYQ+vK4Q7AM5L7TIn2YESgyWFSUcNFVEfoNjwpAHBilCU0gPFF4
ctbDSWlUgknVSltNdTEV2KjSq310UjxT1jKISPAS1vw509iKV4ym7DEoXOxmW/HCbhfjTziZXYAd
n6I+oMPgAMPbxZK6dL+laJxXxtoX8YdTs/V1q2Mp80T86M3L8i9bZlmmxZ9jxIrJtg3nAO8ZlDKT
A6N2/DOXAhYumW6EBbG8zmKqiR17Tb3zsJ4k7/8v0QVaZF6UNJJcUZCzFeAS2LPkMxUCDjERZxMN
qOLMw74VOZ1W5R3zkmgRBDsq/1X/gwfir4KAE7c8awMaG8VkcWixRmU7nHTpe2WuYPvPWUiMZUcV
t5WZ6+a7hgMLxoqWY+jqH76HlhpGeJatkj3jvjhxwjAf//BjM4gc0QVenkf05SkmGfIlcG0BIdO6
XFwrkZCcwGDgpvYa6egcduOdnMJpouPd3i3A51y0OBHoiwKGv9fkmnJIKL8dbHzJwKXghp9xlLjH
ggrFguYTXNPhfEQjycGMwCkRTjtnY0blBZWdsIcPlJeOrDvhHSxw0mrU5uY1QOqtVjqPf9H7Ne/D
9gatRspKap9wQX33Yv+8GHjKiZebslR5PGi3zAfuv6El5up8WMjgI0RSUYWuz2cFtQYUifrrm04g
hatagusYm1esVkZIW3hzX3IVb0HDfmq1mVMIrdijY4UJNufzJa/ms7jSbRkq+lJk0wMh/C6t7h24
UiqG+Dky7ELhv/EbR4KpKSC37qDHSgQYIMmNeXFBa9ityGxQE3FpOFAgUqQuAbCYYFa0YG1+iEvP
6IGs2v+ybrqeWsoeqrSBEypsnAU8D7KSQuLVfFBtqsf//0UT+5YvLAbEp10wATXGlpklkE3nycQ+
qhEjMN9bChA5vtYlPfzphRv90nVlUE2wYC05huK5ggX0Zst7KAtwjWI0OuZSp+Y96qhLiI9L1BqE
TTgDcFOtvSNtmxpLFuY4o3HtLGq2HYay1xrD1i7MBc13dCz8ma/quk8V0tFo01CQLNq00An9ovUJ
qFvTb7cBY/OciGyvLSlo45JRI8nrdjZixpxSPp4ypG1eReF6vWA59yAV81huNBLhRnn0aM4yOoM7
+xWcB1bPW1DjzU3Wf9YiPmQmFfK12ybkAiXtdyLjFxcvFo08FxvjqebBePLhzBRzLTKS5CPmlGer
n26w1ifBjmP2a1R6N2BEPnCJXHWxmuBpm9cpWYUOo8sqVU/2S/Fmh0acVEr+HwdoD/UyxFhPCgq2
EUy5B1feGTCILEPqbJ3Lj49W0tvT1/5pB8e790lTYriwlYqyktlCl6+NNXQu6piCQSNhM48w8sZO
qLpVqlTfrQ9DRGPq/uasX1UkCoKtL8zd0LvDcNaWFqmA5bWX4cTCSIQGzYXj8Nwm2Xduo5P7l2i5
N5aI8FfSGSY7V8YlrxxgWTnHqIYi6Nk4SYnu+h42tYlyo/9mohlYBJTJX50K567RyFyBxbBpnF/p
QVXsPZdcyqm4Tg6dG4HgqFq9PcTHPlmWL24k4NGAb1XRIYFnBcGRDKTruPtghKrmupftK7NV5ynz
13M/swz9+To2w1XKNlRlSvIM5xDjlAVl+H6FCpjO+Qor65Jj4b0MIn06cWvIcTknB7c2tPoiFbAR
FAtSL1KKAPUfK2Lj1tC0d+/pqA+0RoJrVa8SRp3Cn4oei+p2yBYuzHDZOomfaTEcVKhgSKHWmxZA
YOapa4keY9nOpr2jbVXgeihHmUgwpD3AsYeWyVIi9F/U0dIlyWIXzQy3RlK8OWCwY/B3Du5BiTv0
CfSjHXxj3Zxc8vNkJ+XycZmfISvHf0pMxDxZHZ7MFEnfsCWsPOJ/qVzBO3o/BiRHuf7E/psdpLUh
KgAO1mBhgRpmNsfkubKZTreeuvVo1zui2fGl/X7CQZLQBDHsotlXdFXwmgACP2zpzWpG1xLJ7ZLb
AWRuBBAQ2JCCBEi7C4WmAW589BkRZH6o7icLPq7+Lsz5FwRxoKPx5bU7x9R+C62EUNU0FJ9Dz1S8
w/6PGlKwGKzms6AjuIUTYDHRTjMv/7+IasqbiouXoa6vsXMiIPrU9xQGf7WE5z0QOH4pZPCemzH6
pUOqO0bmF5eKT7bNfdflM5J52VN+vIzHCw5bMKs41u8IRJ56x2L3/mQoncAha054uo7ozgrpxKtc
O+Y9bXrR78BMzvSRWYHNNg7i9JUWm8//T5hI/tBgxYi09P3F/3qmOoUO8i1iqxfXnNvQyCjwcS8u
qaFKuOPkstumW+/yZSGRGLk4S+ukJvZlb+s4fOHIfjat/IDB4+09mE+e7u3vazGBe2uq4s/sCQtc
9+vs/dwB1+MXCSuhAarKvNrNUQPruh67wZaIHjxUG5TNeOUBwEHsASKmbsI/c4k+qg1NITdXsl0J
x2xBhQgxih1kqxy7g5a9RZDXCWTpRpZWlE7phodSpYkv81HMUl/FAwF2tFYXA/dd/dVtRnXUNXvd
XJVULTHUJ4bejTXB8DkoC8/ftbe3coe+FkND/76NBj4+0W03EtHLbIGkOxUICpZTJwWS5RhZheGO
6+za7abcoo5dHcM/MqR5l1DqprlfsNvvMdMdMx3Oy32o+SWPzC7HaNjITFGT1BADCnE8REXTLC6X
VPsx8Gq625Q/uLk62Tl6ONrM1pd7P/cb9xX02X6klV5sHW1/vDgPOoTQP+Dct24/nl9roz0Hq7II
0q/rznAVEXBJ74WjffOKYzMgCq6qws9uSb+RJxe7jZA9MTYFa+fH4uB+0jj4qJiEAjiVSzZtqABQ
dO2CsFXq6u7cW/bcagg8q6XanMObOM56zBELWZNwL1skQ7edV3i30RFieuPe1ZQMaZ+rpGsRCJqs
TpPVA8U3EFvZ9VAmPL7tMYIDYfvtsXJJgT1SwHCYshzlJh9w1Ffvbj/0bkn5KLQq3w0fla4YQs8v
HGwfF8Zx9lJsVie7rfB4O051uE4b2z5x3t2ZDYxfRGZi4Oq9QzW0HhgMlmSKTOsr8UsDrYTNHlgw
SDjVMjbOXksknYSTMvGIcP37XceoHxB7dTyMTtppis9niCMbFvd4GmnpKS8AmSzqlGZ8gOceetBw
ZlHgowHNna2XgUsWxLIIF/9TKQBSSjaXFATpjJVOF/NAW9bHUJKLTmbgGX8tMgRxsCRPaFCr1q2K
HSJm0UoJNLgUgSwU4ElTn3vEr3/0D1edtBqQEHeMwbkxdpQ6Pld8OrpGNzb8t6nTG9HThh5GvXhH
cXzKWt5aHnR22Xox2f9Uujrrk0Dilm86yz+7HtSbTR7W9i4IDCNYtExbEn+mgTtPTmvkL44ufimk
6YeugnzzEtfeJdTpXdkvB/jOya9H2fWu7IuCm4huAl2OAqLLXn0kROndABEzSFM8G8B+gMElI3XO
vcMcZXI/ZTVPQGYp7JYfYUl+xICab9lx0Xgs74CSqwpjXYpGPjcETqam5StYIAJbsKgbUNCZ2PCk
AWgWSj+kcfJVSXTNMPk0O49DRRNsA7wkwQVY7zM6CXetoEDljuyluOD9ujLO52zlDccjekmq7k3Q
27NBIp1kvqWDSab4505sqrkvvxAey45uOj3f0kNWtXlBld/SP//Sb8AjoTfRPfreZ7t4W1fn0Vgx
qWCe2L3V4SBShTaepk9lbaU9CXdOaVyOjyQ7dJ+cA+zgITJaLyB2pzadf68L1c10Qj6GWo8wmXHa
rQEe90T9NDi9m8+eJz+oADl6EMCjyos8apOB57o1iGHM79vU0Qb7gIRFPJDhNYju4VSCI5m12ZMe
GXR1KLmPKVFDF0yefl4Yt07LYtKFsYJXEQGcJX7N/QpmvkvOHBHcaWyWaSmkQX/othqv2T0uqTDM
ww1Xwi/4Fm0iHFCm62t1HyQZ3ejfbZtr2xUsieF5Q8TVSCFxx4mTSLSQ7P2Ek2R/bKO4Fd1yL79G
0jkAepl7Qwn+mP2TkwfdNesz07i+beaqX+8xINMDe0CojXIa6gQieiDR2RGp2wd4wsYswfJKqukT
lN45zn38HHTCKgnp6ufv4o8Ikx88cX+THsWGgWwnxhHpRkDkRRkSQ8qVj7R05GqQLsDlVjuev6Te
sk0auGXMktgiQZs/FXCsvVSd+zYV1jduYXCnvEZOTqsSIqXVo3GPUj/RQhcwdQvPaDS4y0KszYLy
hnRptpdwGuFI7okiN/eJfNLCK/1I0G9LItOoFdKbuhC8iDCQRZbAK04/XfqRdR7LsJtai1yA9V7v
RmQKlwju/M+dBX3QwC70ZECNu5RvaUfUo3x6VcdGQSTUJHnN6le4Xh8K+8icme7xaCvIo6m3hETO
p5huBPiclCszlWe+yQn7pB5A5j/V/DNnZsrAl2j4aeRylxcBoTOIN5W0aV2KV2CZZVFCxKuimupn
nM/iU3Hj7qAVJMAeJRMOJNUYxP9wXdUsuHR1f+Cs
`protect end_protected

