

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GGz53Ico+oqWPVynCPL37qIEBfwCVjBweLtHTDYGXIB9pbDfpitk0gu6seoQjNO+tEFN106aIQS2
buWW+EJmGA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f+ecyr/exlgL6N9a90krQ/aCzXXwwTmKhdFcMalb2xa5LYisNSByaSZdXVxmefjOEtdMtzdMchMa
SawS2X5S4Qa7p12st7+J3f03r5Ed/0B0XszRaMG4JzCm6Okfmfbb2tHANIHAMIlxC0T3UpfBAtcD
RU7Ky2JYdulbOvMF9us=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OtY/tIZGcVNATR5zSgwUoVZcp3fChVKOEgUVdP0Thi8povX3bA/amikgZFNjTCMN8BonoudWuJ5T
8+POwlXGzkLyiiHwMWxoo909Ct7a/cJofJRPCmCoZU8nlq/OVDhnmZsuuhezUdvy2lblJQZAWOj5
+P1tTtL6HSBS/4+43uo5PYWmqvZv93iNJoF0NPUVrxdCTHGYnUcVhVLRSpIzXabR4ONfwICDBOwF
hl3SYiGjuCzx2WVsn0LYz9N/7kggU55MtLR2XDCIuAwqeIm8902cUPNpXDGREi6rtI4hWZHhjAlL
Pq90waxJb7/VveYNCoiuWe9F+vGcKK/soF0v9w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ke0TW9U+p7qFbXIbzO0Ht8QzYplvZoq8R+SxzYIaL9hBjS0wX1p8ArICuWb1Bie3E6mlz6lsDO7s
Oj2xJ12tkGFSOBGb5VGMUYiScOwdzpH3irdJ7P7BhVflL71LYIJcwqihpBdrPB+qINjwUrf2Uj4Q
aAc/fiGDGb6k4uPMRcU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aC5vnzxPkc8pQ6nt2rD95lZvdKhLnumEt10eT9h0Z+/5Rudgfav/L4n1JybCrPCBCIsG/SXMLtrk
BzI8DTuvNo5qpY2i5i3oaiJlgsNOS1NmHvygfg5eQz02QhYi66R7Raz5NyO/jaBQ6bUEW3B07VHz
pK7oiauJ3itb+Q65tv3lMkzr0prtl34cxRJyoWyOdf2sn9XLPq0+KJSlOdbpDeZvtjARBqW8F5dK
sLQYy1GHPNxMKus8QhfjiVcBy20thp2b7MSJm0wRqbdeGwjaTM0SBvmQLdatsDDY+jJzwGW2p/qy
Q42+2Kj9/Xmagc8R+8p5/MF0If40PbjOLnfdgA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jmDkMhZqF5kxsn1I0MzTsBhLjHYTe55KbszLon1eFWxROOpc41jrG01CufB/cmYM1IMr/JhinOuZ
02wlq0whuPptPE9ZbiIuSeNL3L+Tck1j8ah4Mz8Y659pEHOMVCF4oLzGoL3vYdi2vOBxYs/UpC5e
bG7sb+RPS4GO/mf+QShhovywptHScIZ/tOm3ooYhgk7Vy+zSDaYe5SRd3f+sS/LbmS2R6m9VdZgk
VIkwP39p7xYZ3hjzGcpizT+E7FR5XWv4RQ3pfcM2biCVEs7HcuEXajDGVMqF+NRDC/uVcI7hNTM8
N0mdcuKKMs4XtO9nCWaqnwNn65o5ZfrhEoycZg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504432)
`protect data_block
DIfHB+OHB+ue/VSHJWTaJqy0X7y22ODMq2Lf0wADdAgpFMZ9A8cENUDJ1BnFf6S7CebLHsmPs1o1
FwcATjLzdMlz07U38kJ0QYyYgl9Etp4oUuo2+05OjELQ+GyoXDHla2oMnITXrQek6KTkQDVJsdf7
OLY8IRHb5AoAcjfl4ZNjWvySH/5qk6k7czrgTABs/cRJTE7/jRlKcWxMTP3LvKL7krnO1S6EmBAd
rb0bnflFSXAq11aHuW6MFxmC8vIum+uzYpgPICWKMn4o2H/DBCTwq5IKSnJ/xysF49VHoWyJiqlO
xDK5NU6eD1SxgEH2vJXp6qNi+TNXz8EvU4LQzeVgslBfQHp8egL/r8RDZNGO5XUynZkiPCQAf8ij
KnVX+33FCYCsGXBEMIE3r3TQToUlCX7V9eYHtOSoikZUDidlTc1jNAIerP1EVqagLLjYoCz9YJe4
S0qn2aMdJtAb1zOD0b6MkV+G9SdBn64QrinexULzxzs/j2U/chTQJR2AQfsNEqjIQUz9CZpaAc0r
fuSrtPh8d3Y2mc9PMr7w4FxKOSWj/Kxng1hlGKkvmT57FF6282iEDWi4V1LYhNXzlOKpdGkWxUT+
v7XmA6/B3bfAm+wFiRSe/74+A73EKAqViExIgHr09+1+Ieyilmb0WzWV82WqqntEWyUbFMZ442J2
A+wtNpfugwp1j5vpTO96bknU+Y4lY/2U6xq9Id2bqVWn9eY5YU1l3tpLCIYIoj6oxbbVP996ysm6
5ww0ex+VV3lSBd50nDudbMcb76TQRuAkSwrAodsJTGRUNe741pwNOD/5xEG8FVp8DamoKJk2Vt8d
23zZx4SklQBEUTYLfbzniA8ZmrJ9jw2E9bFPVxwFdYQHIoGUQKHDn7q5n3ks/ccOM9WGLMEK9Dq/
T8dJaDcgb3in4vTQQ82rOXHGrVrzpKpCOAcSKETtYG7IQnAOcHOj85wgnIuLqJGfJZZFTrz6cDSn
19nEEAgjaE8khgda6qR+mwfkl1CM+9MoaEOfT6P7V5hWafQe2HUAXu16sj1sfSMgZbeyC62Khx4b
Yx6Tpb7KjUR1FIDigvZ2N1bH8ZiPE3fPctz3z5J+AtJAzrVI5pGXdFC2/GXqyqEH3MEaCHPepYIa
MMRtSN20Rd1Tws+KxS+lzxMyRjY0HrdxzE5B+zP3ZARr4LaLD18SgjW04AedaGqdvean81q5jm8z
awUWC5VSUdgf3l7bdHNkQaJoP8lGiSrZtosPRirSxT+lZnMtHavGO0PEbFw7ZxgNzMJNojTkCOZ7
rLK6ogPYLGDt88Vtw847RhYjaGu3HzS+wbQWbiIY7hQ0SydEM398YHWYZTvFnLW+i4Di9fzNI9qy
S8ZlTvarrgTBCuF0kGrkOeTgE5YNzv4L6ICBhCW1qpvo6Ro766RbEfctzsZu71umIrpnO1bQDqF4
0LAwbg1f4kBPWVgDZHn3TWwIuf6rlkUDCOkoQGOpS4U4Uuh4pqvGkbYyNHXrbGkH+0TuiwXGICpK
oY0Dw9wfLvr+aNsXzAKthgybvAdLD/S/T6mXl/3X/P8l04LL0fLEDzCEYCgukd4szhLMiolM2prT
5cp0Eo1qraD+lUOMF2FtVcXbI3CVWJBl8RK0r/94z42igihGYQBok7DyjsMEsy0VRJ121A75zzAu
IVGOEqA0whA/cJxbOKYia3pX0FIu1pw4VaLk0ZHgE/l7uI+epoKPPvHF9YEXyD0EmgTY4k4I1uTD
UfC7PaOZzhosxuDmwbAAp168r+2rbXUVf5g9h/4x0mSQTFnLBGOWKSZTu5asg5isbHUhP+0y3s3p
j3N0YGu6EE/33K8/g4JXWLu/M+hsP+4fa+1e87oV/f/hlavZ3DoQ+ii6n518Dniy1QjgGjIYDkF2
B7JSK+w8exPzHFu4BS95Q8aKGSBwppgXH5gECWjm/kyemcPTozH4WxHxyKst4yGbTB3Oxj05WqsU
SbryGDTnEXuLI4I4LHxQLJPHFA5O9+Wbitb+0xpNufkQNUcH+h2BtCxX0tWhk1XMW8gpDr8YakuP
i2DPZqnGFVz98UsUw5xPpalr0YujXweOc19G+oJC/gDSNcXy5fVCt7S/ttXEvrkOVCEbZOKkklVE
5kqcVC4mPBhgej28TwTITvn46ll+svZMkM6TPbzPwjvcA2KgBamN7oFOzitcCC8RhFaXFYdY7Agl
PMhhuSRIP1AhiD90sFUFR94CAam85whBc0oMjU1NZQeYseGDwQJLd1NalFFimzbj6dfA0pGGWX01
dOHINbLoDEH4C7ffEcfRU2Snxb9XMc9jkHrhs/s+02e8Pvpb3x5tptrXYUFijTZY17IatsbCVqw9
qvUV7rKgs7b4WftO2NYJaHnvYaND1r74NDe1EULryjvRq2SxnZSB09eCDok4C1P/c0yE7YbEEBVK
wjWLJa0dJLyLTBGScC2RzUZZfyAP4Hzg+JHvKpoLbs5BdIr1esRxZJlmqQSjUcvapKrymHB5Irg1
91gfPxvUzMNFw7jlqTSMqrqoyj3c6Tmkylt8uTetLMy+oGQWNL3bZlCokvbezV7nfDApYHZC0M/f
Ce7hnBc/R7myP/yHV5vsQrTyO3B2faUq2itUS9vPmIl0ShDM0K/NgCWldT7UF5Vatb7frmUDQR1e
1dyUk+EVIiZb85CN5bBm336Bb9LmGSv32B0TgwrgJygO+8qpoiOWplHnwJJlBq+CrlGOiadyzTJH
PUHzhlnidKKl3d0rkNknxHu99z8t97CcTG1ThRVwzGK7HMtacKGDkSLHNH2WDPe+pkghWUwG+YHz
lSSTtu6yZYVnZvMSwWNAfzTdtrGT5JBO8JCh9IggTd5ApHEkjSRwaDnbb017VZXv2b4TXIP373ky
zKgT8jUTBLjlzQHpdW/hVjUdnmx4FHBbQmDHwR6uPuLDY3ey7YiRIH+Xjl3/8hPINJIB6/09v3b/
1hIO4FcsIbXRwqFMjQ8VbHU9hpViT0YI1hRKbLGBcZ0KRiDDs+0vL4R8CG71fVIm/FJTBTQrzVsg
2qb7sjnJpOMmVWHMKGE7Y91+zh+oxNzTU/CftgcoxOJ4MCa4XFXHQy6w+DR4CAHbntIlOPG+F0tH
EkuSF3orStPESdbsquLWsMgFxpuYNzOuJr+8E1sIpVDILn+c247LFCFJkrvZUaXUVdZGptUg3zSb
hrQq583K6JDqS3LLKpvzHpY/su8g5D3mJ+sg8KWY7PymrSueuCZ06BH/FJOy8TZD6Ap2UI4wRmbT
WQM42oJfbgI4IlTX3EWqkBiZt0t/JasXsLmweEojStd//VMScv9Wq+xhoDjZ7RhQK0RNx01Ccjrm
vQfwqgFslvaS+EhlV/PUv5DV1t8BS/EZXriEQrQE4pQkhWv0aQGwbRbNUUWdfnyp9rxV1alipWeM
7toD9msE8TOjM9njUtAF4Dl5JceGJK/Wzb5cYbTzRe46ixVQhq1PZ5mfNNQlhs2b/v5wqe4U8r6w
guOxYGNeMv9pN/GtwJ7gY2iPnI00zlSEANuCz16HRNpbDpF46O0crYfvtPFRFppzvSe7FUyiai9v
mluXY+scGmStmOwIesfHAdhKCQUeVHjXvhl68K/W2piLlH11/YiwGp0VJNDKr6ouExt9XuG17IaT
eyjAm3WLjYHTz2do4q+dXUd9HVo4hzjZafpJfypzJcFWFxjsk5UxvezXAviKl11uko2+PsJOupz8
WE5u2BoEZDgTCEAKEa4ibe0MTP962NyFzy/DZ8/+Tm0Dl5Mb+3EDNITnONykimlXUrP6WPWW5LQn
qNzYWLpTu74TVcY3QXhSBPSAfRXs07sfSEh3kEkECK1TkN1hPXe0qD/sn9SpPabazZrCvPCraFu+
qpc75f42JFGodPFlGCSkwqaPKhAx9tAdwn46mNmPJxDuO8w2PfFWIS30gzzzVZI/0N4Cz0m+gD4B
YybmoBkU9Yw79hTlOzowkd1jxJ8gqS6LulCXanI3XnDM5YCY9hK0YP6/ezZ2X13cjhhmlG2RRUNp
3SWFMXubkM6CL942PUqmom4LWjZoSUNMuLIapMyPR648acDt0vtOl1SBCYop0DlViyuvaD9sxclN
wHzKJealeT4NLCcwookPZSZ9Y0IY/dGZ9GvnvKlo9HNs8+Y+aHjvwIOZI9iPha3b/bugdz0mjJcn
ZdvQsl+byWmFvJTtKNa7D4HW6MWY5fMkqFopJQooW8+iejFlxJZcYnx5XYXkIUo05dR8GBVk0Tad
kLTNV5AbVil0N5ah8Fi2zWUvjWPVyGCxERNp36hVSzq0smOLJoqruLr74+VVcJqOEHbpjzNec9pD
S4RXHC1JOlzh95PlPuCyKBk2tmcO3fFRSxxkI4/p1GkBgDfJ1QIOQ+iOvLlac8+o6yUYPNW/dZqI
uYlAADC6nLgZR1zH5a3hOMh4JQkqO2zQMLIRIFLVakuMsrVOMVOSg+7JGui22cUiv48ydNeMa/s/
FwAL3qIzHIyVGLpIBXAcVbygnHam4tGkIUAxwW6IwLOnf1/ICPB4yRNeCJLvYw43Ax/jNWtF9Ko9
0uvhe8XBmz8w8ZJQCOyOkht862TpfXzxDXqWjVzghUA1eA/t/aEQPLk35nXcdfRirdM2w1/p9fLm
D7gwPXc8MgfIMQosV1R6Aice3Z7EAhlARPB6ZM5/Aznx2v63HlgjnpAG/9xJoeAoudBK1LGJ9WBI
vGaG1NVqDMeGANjBHaziDddCrNa4aeEY16aeJ9lzei2cb9k9vR8M6vc4k3PEDNlJlRZHmEx3nWID
nWC9495L2zPuKndrX/Pa3YHhEFD8nEzjUEmyHdym2JcN5uKtNTTbuqxvIGgTXPkNjEFyDA5TLloO
sIgiNtuCn5NnNHX0stcC9n1UXLYgp01Z4GB2Z3JeQFdr/uS5+MzoZtCTHKBOseeCQwOSZU4R1yAB
OaBRliu7/M33Ky3o/YU/lBh7/9gYGxPphFF1VHotzKuLSlM1DoYDryyCnIXTbTIELI2k5UECLSaL
QlcuhIAP2CwlCchwm2JvfyOzNyZL3lnJQZfeCZKhjnRYPuGvKAsTPH7x4vFSoT+EEEsaohPPDPaR
SsSY4oPdekk2WIIF4HV8pq2N4UNxsubzl+rc4sYrnCVZjxHqzqGdbW/8IfmpiPheKtDSqBGEUs7I
PpzQB6R/gol2hn9EGJMFferIC82jnPPxrBj8+oVqyR4SFNPgZCd0VSM5SWvVtWlsoS941GGsYGF0
30bFJJDcbGS+qwYgeAnzLHfbfMO6cGD+t2wHwGn2XXH/PzBnuYl8THNH03r0JxwXaLxKyrfwGLEF
wAftdZdF4p/9atRBsLffxmVUWGX6Bzgkjx9Qlx3bKjBJkOHIV8xf5ey4rMGbg8IAOXLNG2Xtszdo
eOb29uFt3mVTFIwLhY1hdHmP36xRlSOmLgYVCuIKA4MTjmKrMGIfJBqMxbgm8jb8EEmqJypAXPGS
5db/v/ikKAzfVKBWB5kHchV6ULyEWJ4GquVp8laWuYCtCXS3qh/YxHjzr44umA0LVWcZpy0w3vZb
VngjUjDG3hHaRXLotSpE9fnOuAIXbxDN6943Dbjmb2tT+XcNcwkdcxxlYEjOI7r8i6awm7qij3MM
/V2UFwEbdUS6wtmadKdRYfg/DDepm3sVwzaU+Vu0WBnWqUkxs1ljJr7qv14PPNCJQrg3soFKuLqx
ntw0ojkrymc8BrkfXLJolRAuGXV5Wk574gHMNmdZIzJQUH1YxaQNbPi3leWVfwAKGTydOIKMI729
6Nt04orP/ef/CPLktqyZ8BRkTYpjmURaC3dQjjGY4l9tn1Y2x0yDF+L+Vnw32elEL9jHHhty6WcK
hdBBfcEkBK0J7yD7gkQgkmv1W7+VZPvr6Iqo/jlXKEU1kA0qZ8Uq371TEbySSfnVsKyqffQto2cS
8hvcJngD2cSCESAWNjjzzSsHD841nTY46ibz1OIJsrOGd50u+iaygM/vTOTjT9+d8fkVqjKEE1X+
H9EEEzHAsUFQ1ozJU2wWJ3oVw4DF7gxSCygqgsw9nnnoS0UC5by1jUNx3lC9j/uuCL0nO6GmvSg8
HoNpnah1yh3fURixF255Jb3fvGjVHkwitUvI49cvd2ha3PMIklOB/IuLXrUie+x4WtP65C8WTx/n
25/Gzmc32E+Yd7DYM2UbZavqQTJ9O8mFDEPDL44II+6AxdFjMNCyL1vuUT4bgpchH108lLZQb01C
U1JjA75sUcnpWQ83rxAifRakWdgrKxhoMLfZebYSGjhLTv4U0rEPLK50hZrsnpmi8MLaPOUpYbhc
tDaVvxe9dUpYsa7qGdN4yVl1oCVO/esqyuK7AKFgcgiSzYbjgMele0Jqbblifak/MVUlVhcSUAoy
rmb3uSfxlNRTMpYQVLoXtYP04JLm9b38PLtvwEFwqVLzNs7FkTkdN++czq+W5vKtRGryhiGNKl2+
mxzIoYhLgvc3dHN3k3tkMiHt3OC9BWMggGRbb7Kou8OZs41w2thRAWAGeEUlb6evu2uINsiypZRn
ART2eUqj/y1Zntkj93xVsYW95zPcADccLeSvehf4+UHE/fAiOURFrya+NBSnLcDe8aMq7dtNrrWD
DKrvcuk8J007CVwjiP7PmZPRTTZQ8v97tEeMzFGKcxzisYgdEcl4qYZ9/fKPGmwmYu6ZPiNICFJv
i0QMrzxlJf+SgRAV2bLnWCi8U5kqSgF+KcHR+LF2TxPEzx8gsyupB3pArIn53DKjOBjus+C0cuBl
32OvaqjMsD2VuTcuE7TIf95GB1htYBwOmCKj24n4GPkfDF9v+BVcGsnF6MmUfF66N/AI7UCrxv9O
NsnHgGsTnPJPB8QDorZ+uNzvP8zr0KChgKSPAFWA3qEajwobGpHLS/TJsSa0QewguPC+7Cod9eVx
MDIUYTm/AIFlLV1NFmkRo9TCTZvVO7lwo01cWXY0FgyqWekLOr2ld56OYpgB3nJM9gC2GCMmnY+w
d2XQr6nUCR+su9uZ19NNUAHJyFaZ9fC44FdNDa1e/fvJS0KdBVniK/ZraDd9Zq39T/wV0mPrZzA6
VvEKsZSrw4aNytf+7Q1X49J1g45WYT9JIoNXwolL+MsBLuZrzI/yF/T4XVYZmkx8Kp4BVwpjuazE
luBtYpXDMNnDRgrt62IoNSLqiiznxAGPJA5LaMeMod3Ri8fC+qJN29zH62loB4e45oqgQTgiTV20
ADZwZF/dCzOlIST07DJrLR7NT8gqSe/8NB40EKWw3jKyGV9SnazzH5WcaWWJdp0IUbU197PZvzc8
urHc6WIO5TXrh7sWp6J4dc8fDdmCtJLB9pwq1Vrmh8cNsd7rZ0rRYc5cxFxRTxjM2k9Oju+Aezpi
3gFgai5mthHkz1T7TKRHBWXUI8IyHXDuJocKbIcKeZNcjUIbPzgQPBTlplUTiHSEj9qa7VBVAW9G
btmXhgxWZs+Mj+8aw8b2axZ+wPu9RmbbTT7wJ6qh0M9hahYNX2CjaCOi08C7sPHPLp62tO3ysJFh
qoUf3T61b/SRO70eBW10yLoLds4KIwGZdd2sf+A1ft7dlU4iRXMnWKP6dqgOQ7bkQylFJO9nrw4K
5PgxXvt2+1RMAuYSQHCyltT65qxPXpDqiFMx9PNC4bniBT+a4IPM6V3B7RPGgV/aiLdXwXXyUi08
TCTcl3aOLmOU3gOIJDDb01pePbKuA2bmBdNt7D0gq8JB50p5cqhyFcjO5nnd/CaU1g/Gk3Sg0BjC
kOC4s0m92LvNWrZKI6mTlUuZ1rYDC4wPeY1GEMGpJtOXfM9X9T+4ka6IJjomBObmfDu6+t7rc4n0
f8eo9sG1v5XSzEmciiCqU9vZLnAq0IHSQOFqIpPp1mM2t+AV7coty38NNOVujY2HHoZKWs4gbSmw
p3e/YjvDEnridpZvBcPCRmt3/ZzM8Fl1kkHiEPs17jmjpVPL2R/FJoSin0CyN/O/qdDMRhBR19qS
RM/bQiMirQcYCh6poZ9Mb3Gi9jGH5fLYWPXRK2NyRQTVFYfGzKim/Um+ZXsZZeL/BJCnhsDRpoVX
S7LSroxHp5fl9zdlZCDDFY+yYtrJF+5XiKWH1IGcUjdxeBJgmYve/NMGFrMMzPj9YsICEGxgTG0e
ary+y0IfRwkBXoBZS7fLkKffKpnT3/OmxvCZGJAR0r9X0WssDc9Wghj9zWLpF4LiR14O23uPpcWd
fRz8+f3zQtjF1m0NGoQPY0uyWml2IJYBQcnCTvZgJx/1DxCEGPgjyCqK/EhffgEygJ+JrNXQZPIk
2TBq+MsEiE3U+N3UWR1GttjZbr72jSElLWbqD17234Wd3sttweQKS6X5ms+2fINoaXsRl3OW2gZB
oonlZYBl4/RdUuSvs0t+CRtrR6vtwj+1kN1UdgV5KAbXeqMzXWh9PunrnSNoBL23XLMm3bDuMJiv
OV2kzJW9tyn6IlSWvrb+JHAXJl3NsJXmIPmm/yccIynbyhHZs0wPvOXkVx1iE5HiYIGhSefsGC6j
J/mZbxoZ29+HF62o5vTtwO2fNunbtxsWEfrn9wPO2YfJ5IC95QGwaBohC5NIsK+aM+mpirDYs2My
hHZyf8zy/t+PJ7Jt1uxuvctzqLCrw3eyyBx/IGHtN1OoabGLKlcIydsNKSfXuVRcrrP71cWeC/OZ
Edfx5xSZCCY8qR1sAy3aJlc9CQSxwNkfDVoQombya5BNB2C/Not1cgRbEQ+zaWB6F1X8EdxHmR/X
uPR49cezHezRs813vMtGeIPcHx05inqdOy3eUi0DtaDsCG2AxEhUPYngtWSxFpPev1mMmMOMJ2vG
8pYvOoUReavzyYu6GRgmiJK3L/9ClQkstaH40kkU8EzbJrSj8oq4HIfK+AlQ7WWLSPYcIcjG6C8/
0CK2or8w+ewBfRuGahTxHbP8ZL5f1N7v675+OUqOg6fE/x8nGCG8Mi8HmH4nTg8nesNUscHvnRXE
qpJTjU5rTdmG00OoSboLpR8KIzPSMtrQ5BQwuRQJhIOsDAytbzbV7CUspfvuDjWQBFem/yDPMAep
iDDGd8pNXF117Vou52gzGwSjjKMlvVbBBRo2UPFuBXQw+dwYINf4CwYJ0Q94dwjbgB4bkILsblFn
0SZjw2vVt+wnMorOxx9ijrFLqOwxVdS8ZeIiWweCo0kAl+KqqBe+6BTcUj94zE0MvRm0VIotQuv9
rSffGpuNXsAh1eLsFcq0MRQiryA3ztBaIWJWiqdfM9NxN1gdK59yOQfhAO5apZenUbaD0ZTHKGIm
35phZw2pyP2bsQEE1mpyWTr/fyquD8QNMOK6b8V8iv428OIQwxmmqh0yPZNfhS5P9UkgApWCqA+7
WEC9+uSmGy0eqYy+BnE/JSmM8Vk8d29ylaS3znfLG6lVtzYH/ahbJ6LSeqqtoAoX5Rv6QvNhaGZy
y3YNhKNLNiWFVSHAm73phqRtwpSUS+jj8umGgCw+ZKyVGRBClTqIwmWgAoJPfTE4vgGi1bjQlG8F
suzzNeVKVfXYHU78M/XwwHzhIB7G9nKDfx5NnploJTNYX8gJATS9Bc5CmCUiOtxq78Oec8qTShWP
wrUtT1hqCZkO7X1Rm8O/wYKuwbZQtysi8cz4Gm8381/gkTXRBqhT79R4oH18Wub5XrOBWuDjrPou
KZg7WARa+yi7SkdxFSRCICv80Zi2a9ZNp1ZkTWFeHTr2I1eGspKroE8AFy4deU6Kim9HVIzSTltV
P9ShAhKAAmS4KAa2zi0NE6tJ4VASuP+ymyUmFMRaj99LmQIry17WPfSVdJJ29eo3xXTGV/clGJhs
o69UH3l28xlO/8uBgFz7M/whg0xtC8mrJ1nvtZ2UzbpFDHq+ewj68aTBzVZLZjDnts5Jtmd2k+pw
/l8qIqNIowbtLV9oXvRHs+3/m4jJBpEJQXbRa/P+YEbiJ+lS+K+qbeRyz93XUGzsjguL7w7ureYs
ov3qPoV0hE96Bu7/KF2t6y9BBUAtn/2FvkNfyiHu1AubAxbJHbtlVO300kUyo1AC21mmI57h4JN8
YWHPZG28GiLWmzvRebyyKvpfVE04bYQovV2PCVSiGpS8emal+WbUFY03pMSijfImHz0Z8uLKmTxC
9Ra3xEIs3WHJhhSKk+oWFDyn1CAVROCeYfOBAQPpZWW6NC9qw4g0KpL4zus5n1Qikm9CKfM3WFEb
jb0Dvz7HlmsGCBO8C3flwK8O59KfC7iALlEruSCNQmJ276EzzLclhm9aKj5ATs8qngumDafUkJnE
fQbXrvbtJAqVfffUBwXIgy+24WUOphkEKQ/CLntU21RW7a2z9GS8pFjQw2MJ2ZLXoywyZw+LKXIk
gcd6qNpIe157sp7u8NthpmL1cAbA0KohLjpPCS+R3C7IFZER55iYxbgmTyEGrTeli4cPAi91Osfn
y6mtUfCThfQbJsbZ7k6eTvPIE74glofFbflvXGBw6rDljo6JOe69XFAA7cmMECmyga+zsn3j5mGD
Qx7o+BKswYylK64fNMH1EtTyNt7b6mic1ghqTyLAGu52hA7qLiFhvd+KZxzfVElQUfilDShregUm
XtWH/QB0ThysFkBH/KdE4t8sWUomVYL+0H1sKO26ZDGullT/NvFUhSrn0BHWenMC915mcZSY/Ije
a+yqUU6gDBPkVGKDUNZiue08C6d0cjBYjc/hrMIJXZTXHB6NTEzjcnVLSz2IeNY7X0Ijn6Mcd4m/
yxRd+CEUxiebTBVVAMeUBDJ9TP0hnjlsWYRZUTxmeyO/IxNNriZYV14xXI3uzhcQieLRBH3GMeWL
rurlyHjHE7VIJfnMAizLTZkb8SWZh9PuDU6pXrasyY6U3K/I1REwoIFIMJLmLMuFGbw0eZN6Lg/V
G8YP3UMS9rH+0TwZo8uclifHOmv1mMCcOrum035pD3tJb3NyTl3c52u1/1ndQC0BLDGofW1ahl2i
JfaufQaYTDQyX7MtIMmXsYSdDfcqGzKEw9Vg1Je5cfdyXAx562JiLTNPEL7Wn38SpCZ0mOkxVOj9
XTcB54JxAWPB3L0h7RcqFHdfHH2W9Z7FSVoam/h0gxtq+osKkNW61AQvwuv+WiagePLNEZ0D1PDp
6iOqWkIIKxmcaIC0fxZVJk1Ku7uPbzd81UFOy2uzou4h+LxnLzqBkUtls7qFhF1ixY589iAwYLuy
/hxiWusW3UixQflmoTYvAOqc28DkCDxKtnRg/rwInT7lDkPWnUsuJo12hqkBMvEHYTGwz9jiVxWh
3D9Mhdgve2e0DvJNWOjuzt6YBbM55KSSVoeg4bo6nMv0yXqQuipTbaDgRpNE6JXRtdD2vp+zhYkv
4vaZ+43l9chQHKgmn+v6FQ3x6ypmjGByuGc0MfHmCEBy7zoRSoQBN6KBryxhG4USDa4er6CA3vYT
RPh5ArBWxxWO1/N+2uD6BUz21XpTC05lNQVkmajCqJIzL6b2AfesSK901MFpyAKbTNFKZuXJsocE
mDc4wMQdKAYAgXmSABHJzmE2G0ggIZYptAGmhoBftaqoy8+dNe/RWPFboP0ikpxu7g/WMmHUrpZk
3lJYE9BEs57TkJYZbyJRlYYpEcfKfJHx7C+b/bW2Y3k9He8lxCuQftsWx5HJbkVkFNTZzDNQA6c5
UOX1K+P6nrtMFXXvb/g5ZnoP2w0zmDs3khtoI5ojV5cQ05Of2B3IPXp7Eilvxh6nvlnZIMLkElHU
8YXQJJ3XnrOzA+VEn3WlYsAUT0kOjjEt+dA72hp1T6//MTimMdrZzfQtd0ViuIJzoa2CsWN/KiJQ
ahFnR7oBT47VBrBldESxS4FaHrX2Y3Mtyfq3z8JSZ1Ma4ZmcyOG35jF8E0rFyngcmLCAbnmo+kI/
kIM+TVGKunfFRlPSBfabXLs+rLhhRL8P7OMHry0UHFIgthD/+/lZ6POFsEltAwNM+1iQ3ib5p7eH
SH+vv/9nLlOKMJg0FGqBIJD9bprVYXECzWM8jpCmXcVUt16DVWGIl91eehWJ1B3Z0U+H/iZVorau
WwLLhAapvE3BkGqCvjjVOCmFGV7lX8sidqh3iITKXsu0QoiOI78Vqg0nx1AQz8Q2N2TGy09Oznmp
PfjvnLqaoirXP3YAwxFz0MkOIPeswj5sUdHqJmsQ9zA8PeuzemiYxhNlCSiN9M62zUj49A8Ve8gZ
m3WmTVpYL4uzBN4k+2duqSLxzGDBvYlXEyjAz82w76ROldbvijnNYVarEb+GwZubosG6dILAJDIg
jGEaIOMYLQZGgC6/95Z4vRFuyoOs6rVbC3/Hk0yeIAqMaiAzkCM8cFoe/Y0hsfMoZP7n9eDHBFZB
FPVhZJTPDR7qgKIIyztFkmvxjcWypJMqHk8CdGwXX0EbYVvJWFNQQqqCv0659Ous6OwuY+robbqt
jUQNm0rNhHiT7D2hk20EPH9BtBOuXn/RaRPuakMbp/3lu6/LAz8615RrTAjxJVatLUWfw5bTAAwR
jw9/r1ycnv1+iO2vvlslFy+PuO+886r1H93lGIbxQ7ZxgnenReL1ZOYzq9fmlbjDvUfbBtFBawbe
/OjxXFoWhS6NklY6ivHEVqj+lvib/e0X/0cRXa/3F34/NBV/I/oltHm9Wr5sN2kEbfThq30HxjAU
jZMc4iYCFF80NO12T9fADGzgu3KtfZTPdRc/lRFkuh1wc2w7fMk0UkEjjA+/G1z8nqjgWjKxXHJd
VJmJ4Mp07l7LtyqqIOx9YuxVrjgaLEAO6JaA4IpfKQplQH6ZHcR4M+g6QUasO93S9982blCRv0pr
xj0hzHEA2vATcRGlUz7w1MHFsMQX7OML/o8y1PWMnacnLLdXefF/+iZspVCUHOoQa6D8xn5Kr2i+
55e2V2rKvK075dq54kResMPJweUV+9i5XHygUj1rlHcyyfRey5Bsty6FRoirwpJ3EH87iG1v+tRi
0/Uiceze3zsod+7OehVh/Yv4I0NtYyKDLD1u5SUQRjnlyIcU8PoN0VW1o6tJBVU2RQ5Po/Ns8CL+
hzQhrrYgLstBwWcyyYCgkXh3TRO7VnEinLUNBw3b48ERDJoevVA9vXQpCxrCYc6siICgTly/AEcg
CKmovhPFWqyd6Pge/hvG20ed18uB+O/fMlXueqB8qaSpP9r654Y9MgFe3GNeHKjQC2lkzIwV0BUp
UBNSXcMeghRKwiWrqPq8OfmIDwiNWZVrI+m7HjFYKs67B3/Tll4wnqHuN62mEza7Ip0oXQ1uvhy0
8Lgl6Tdcf3hP2oaS+810Ttw6oqAnKIoLf4Dr2QECY9GereREFd/DVAtSSopJ+1NNQGq81o+h1kkE
50IIp05SUpnMoSrjGzo0qKHZYW89Uek5/3vO3bQl6OXWcvbyR3nOEYqcw258AtYX0/+5uh/zgnAd
nUWE5H9uhVDTxr/oNrJX+vefkMF8BW5zPAgoaPO0kuQ7DO1yV5njYOytimvaHASkshRg2tm/sH2O
nCsJ0BlQ/eonb7cdE5M1/6KNS9RAK8Uf/oQO+zinuCpO65PBPATDH6qYY0IkBDnim1Pw7axzbH5i
R03+egpdY7i7xrUD74ggX6VylJkJOLB9kHqo87IzTY1LQNpCrAg3sAt0PF1DF2TNsgNsCubiQeIf
M22nQ1V3C5/WcVxj8Rs+gcZAnNHThtgtG4wQSkDqKgv00/+S/kKLtPHft1AJehAG8+rfF16otmuN
EGGJVp0OzJ2PxITNubyfmaYD2BB1HD4o1C7VYOKRBQAv2We4BZ/5EQhHw0vD5SRh9O2wPckCgDuT
j8rhZuPXlGS2+L19SpAgHeCW6q7GTW5SMmNayu0xOullh029wAlJR8fjGn+YGhwxDsJ+QaQ4QCL+
Su1LjiQwiPsEbNrXaTVN+Zb0tQpxd9AhTPthzkeJQCFMEpeG4FackeGPDRLyqVhzx4f/DjsoHVaI
CKLU4Dgn25Y43ssftsEx9CCt2jRkMDA7y4QHoX/RLqgtOmPexQzZ775H2/paOBl1J80taRQXBsGb
8tM0SXJlrpYJSSgLGunu1Dd/xVPMlt4lPBU9XroFg/23hYqiQAzpJIQkJWUu8poantNUZZ476Xtc
noncZC+e64czwaaThMxf1TSjSKSIyezB7XjsJJexAVAipDOl0mAoNVxOPkq3OE+LUOVCNNP4ibU3
IjzNXPfOXAbEE43kKnzU8TYbOt0j8oDtPPuL8uJLySELk20fbAdzbC8tVtEE57KqUzy+AWFv6i4f
5Taqa+8cissnND8Zsxlx7LTvzVjVIIpsnhDqfCthzkCDwxRQV0v5qpuDvFfoyup+mIhO4pNM7L3G
86d6kB20EaAj7cZXXhWSKWoP6dVUqpyN8bbs4jZucA2RhVOnPe4Xm7gmASgHG0TsqXDd87XOKk+U
Ic+I+1OOwluhrzYKww0XBTWxufUbwJoynrWSDDXZq1mysWSlbrfpCaOhSIqWPOpWBe7QzQGMetKr
gcT+fdXZMRPLVEZTA40F5AH9g4X097nCs+i4graIOJtJ/YphJTeRJMaMMpp8UHEAcioFW8VIHuZY
KbyD5Dha/Yw7SR0djWnGemaiwKlgIRo05ynYaVLBVZ/v2Sz4O3DD/UMnTaZgWWsPTZRhuxlUGPVR
mqHsmH2nwjpIJAcs1ckUxePGIDmiHZ4MpTLVAYFjUHLmMFGeohdGii5KpN4wnUJC3kd3JLW8E/i6
oYzmbWeeVTFZg5I8RKRr0TbLtGfobvq34JrIioT+wXytXKpwx1+Bb1A8+yvA6NvOxYbO/U3xkbiJ
8xaZrB36XgOkPUguLbu/zFIXZ0emW9NaJWeNfg8wl0wgbl4Osdy1mpVimcFDV+Mi05OTknuuypFu
NpNnlvdy8aqose4bwSAWvtP7/THQ5fh9mxQArVeq4uh9VjmMTegkThkL5U6u8AIrBWnrAVM0J/Ps
PywOba/gvtL8GoRcNKf8SgirEwaNzdMKPL8YhIhvLY+5jrLifhCSdBI/TmAZsy2iYNFb/uMqBCaF
lIxnIeAvFpIivAJtLwsm4O3kLZRosi/Z3Fn1IW1SD+LJDnT5tZnogKB52BiboktFaGzaBbrGvgHh
NVagQ/8tDEj+nuCXaFyvzO36jZYwA8QhGb70WUWNGgwimQXk36zMmkq6+R86jJVWxtzTgdxs8vay
aVQWuSqJNeaI4sdKmcHON5LLWaOY/CSAemBhiMqYF+u7J7/ottzBxexdu+mYJ6LBTbSHgDyd+okE
zvELqrMWMAB2q2nkaGJNTMq4bcRN8Joca/72TyT797S5IJujKSnHf/fsf4chUHEkBvI9dzkz0/SZ
lFlweEQS2cxkFeLhdmOANfSAZ823wh0bcRuXmxrAnm+YYJwj0XrHXqmCesFRhcZ1/IKx8z8iQ50p
lHmzuHrcjsbF1KVdlPRX5XY/wJ/pNeshs/plYbm4O+muUYUR7rQYHDvDWKfC5W8Hkz13Octzns3Y
bIa+Ip5IEqvfYv8slBWukeQo+u1nns2tW9lPS3uql1uGgRt3Q2by0uxuEvpHQpMEIGYxfpG63Lrw
4ylQ21IxpvlEt6vf2qy5mZDgbSuLw6/0icR1tJuZfHBrkyr60abl4JgUor0BeVPrU7mGV/Kza6UQ
4jgDElxzR7HswHtInsNYuTSsSNIAhu+/V/x222H2S/8vObVD3sEN+Ec6YMnIOFGY7y1V0og7N5s7
JaClBOIGgI9rbgUEG6sul+NDzkrFNIyT27HRSksOfXG5FMdX59LoXx/zTzEMdGVbjhCDP3cbCQD5
bHmVCcyjSeaMPxrYYm4QvWh71T3rtNgFpSY+t4MZS2fLYzwx1sVhCU4XQ2R5QaZXhjWPER1TEA5J
fmqkxoMPbNvOY19nhhTM2K/36nzu8YKMrGI5izrv0F9uXfCPe6muPt/Mjh7/7y/+OEUvbwWmZZgn
O04AZQzJXjHboWFjP1JDFdCsLhSQy411GlVISDq4AHodMwXN2gB/G7SjUCBdYvuyVnTMusoofDth
Jqd2MuyrahX4dq8gTgGpaHyTOFkZmSCajJWOMm8ZKoi6AUtpsJaz6h/jnYsJZhs4WHtfSaqENIoi
ich9NyoG0RDneGw1uw45NkuY7gNXhMqhwgJEDP/XP1ErwqSnTp9fseosphSoSk3EOQbsbIsoXFxe
wd6n+ED60ITwMx9Qa/KP1aDqh3o7Q3K8Ja6c+Of7Pce0MGs+taQzsc0NjcoxeDIznGjhjYnoC8cV
QDZhsOUisz8jh7NgmCqBjB6Us2vVbSu3CpIL3EkJBO6KUasTJZYdTfn0V5afldJnoN6gvJ5uCFVB
QNLDh92PHOxoGP3uCqmdXyQ/bmxESpTCghCvg8I0S+9J53+cf2FCNKCxn+SgQHi1ONL1zbaBZZD3
VT11jJbAlzKMy/svazTPW1f2WmH+K2lSxX75jULrJ0+2kRgoKtCDlRC/lbqLKLEboBuh3z1/asto
1a93rDC1dLPZU3aS3uWaVjat6SpHs+9nvERfE/HHVA6E1suPo2iq/wrqcCoVLcDc9V6iAQTK8/s1
qnhoBudlHiK50VDu9bVMUYeWZdHeY2ZLH5KY0Wm0kn7nt2Q18rPOv9XT8CGyWj62yIsEAcnDgvJB
jV73jLGwCJBmm4h/+iVVXRbzaBY5zGD/MK7wjQZFOlcg8i21sJu33W3u8a/SZcpuaLg4+F9s8dsg
H93dxx0PggjBg4RViOnZcYWdH5GWiKvkOcryjdY+5J9FItiWyKWVQ4Z4DInpSU2ki8t0sFXvSycX
kpm1181CpdvzMB0TonNqLLLK+UBO56GpPO7EXtj7C0xN6pu0widEjNctCY78LCrUR8M//F5u4MpK
8YT4j8EtzGsVkr9ZyHJoeVaIoLznW4TdZU3bLWR9AydLXf8W74l5pAUN2GZYx2OMjGRlaH+aEmrY
RYeSuw2HGmdRg8JB2SJpL5gW1U5C/Ry4nSDD1L+0aesx4jI3wOGRG+9DOVibKGa37OeTExX713v1
zYxy0NIJjCYN7hR8Ai9OufI6uf4OxjYfGK6772VKc8KlllS2b3P+4ebKoxe6uNFI1p/om85HMdiS
Ykea45F+uslKDS4KQXwguOk2CjWwHU7rmxvhSFabGTvyQpqNO0ZCItfA3cVMU1L90JYCBpG515K7
xMwCz/Zbk7hgaKM6WtI8Y09M4J18qY0vtgvpPmLaGmSMWSAW+75yZ6ByL7wf8P/hj1x04FXlCLps
BBZx4TWvmy/xR0My3ceX+4tfrcsf+hNZyVr0v5eizBGu7rsxcNQuduCq5DAC8GOgUazEtnaOFCKS
NEvvPhjhD0kvR0K3uvGZCVLejnsJIxBDZxtBpGKvHBAe1ioG/B1r48NM0woy2W7IE5a3h+lv3RdY
vj+uzjyG6SfFL4nXGs2ZKbRhj3E+r4RWYoNu50n181qQH4qar/6W4jamzRPAAEnlxSk5Bqp2BzOy
jA3L1bIwAKYSdhRd/cqxVpOit/urvlCdmzAEKxDwRLcuyjMxaGfGD0btYdU4OM9tOYsRQ251jQwW
esSz2pna168HB8Ty+I6cG0srMDz8tIBaRqnfBjj1QTRZylpilJ441tgg6WePixDcnprZImI4pcQm
6UtDg9s6ph519yh3M7ygC5YoHoBaIJajUg+SLtViuOJe0s3oy98KjiWHCqnJqkDzwrvT8//wIykT
QvP+DwLOa2rP1Nib7kNzYsdaarS6TSOjSk8+YjCCXAst4a1oCuODu4ktSJz1ke7qEqbguU7eGyf6
a1py/js5g3qgEvz/+TJJtwMCHYCr+idqgsW/fnWRQN6Ah7kABMFSBknPupNApmQLPHrUEz7cGpaU
ggJNTDZdfIbRgji99BiLn2+NdS9hzdNFjiTXL9EY4nnkofDkCiky+MGpOIf43/lFnQhJNmsER5FD
BmRZBaBEsqj19Zho0hhHLOBl5pSFAbsc4tCuHcihnD8YTQS/O213/wkk5x/gD4JjcP+FUBA8elUy
QMCkq2mA3Mx+fyBZQTX+0LoNmMnKlen+iXePTyc6tU9flIRZswkVDrNMKW72/TAYbS75OqdrYx8x
/DAxGqsrsSS7EfRp7++qg+pxxe8G/A7i17rKf/OMyrmGFPs3mqvk6/QOVxJ23bfg8F7TejTBvfs9
Bpxa2Cz9zPXd5SqyS7rOSzlicYoU2H0eO2V3OCrFqCZUXgz21bLbbzvhSPjabquWVdDBbU+QFUmf
U608soFZ8g70H+hvMFlfpHXRE30uWyxDR6S+IGDcIbtqrP2wbDmVOCHSLhcnqmabfiJVJZ+oKdZN
EggT4OhQSZ/Yy275mYehWEyVO8pxnz1by630owsxD5CWw+nUljNtJJ+1xT57T11CiVPy8Hrp/EbP
QbiEqZHhe7k8s6Un+wdWN0N7Xjr8UAM+85dvw65AjwE1fMJWTgxiN6+w7lZ4F4qG/2hZYY3oJQyM
ZU1z1UejHOJcq3B0u/wMnBd15cAhW264iwLVrvfWv/w1F0TUdNbE9GIqPpLtdi82jkCaY3YHlELS
cr6a553O+H0idJ28E6jsP3MYGiSaHjpvqHgI4FAQ+tqmr530gcW/BIzN8EJ+svrf3fYhF+nxlNuJ
/iHjbL99/BFpNcbWJ4dMEcgbcUGAOcDoNv81qOgRGSnB11qaT+CEYzS3dbZ5jAuh2MKUwmIhbp/M
J0fOU37RYUfkHwpkm/Zzoor4l0tmPOdbiag7/rmo2TilxI835Qvh5fPTphK9oI4TtA1YCgl7SVxh
PVakzhDguCFGpvuC+YWEiSr1/kFgl9/NbVJcxcYw8eLHIvsctvpN0l7fOkrE03HJ6mGGIrlg6rdJ
T9NlykSvb/e6iO7YCkxmOGRF5IkbU1IeRgTlJYC5LsCU2UnEcNofNfVX6gAJAKr2iO+d99RckUYJ
tvYaIO9QvsT0ssqOD/hudk99yvyDL/aCvY5pztcF93JmAujna4AYRAULFurMqCgkjsZ0PcJbm6Ew
bQqgJF8Ops+JI8rMTx3zx9CJP82fTjNe3dGUmCpySrrS68q9HOawH/GY9To8l8YYQSAK6d3GUwwh
glyqoV5SkXab/q4jDcPf9LgojNuR8zhkdLWo3etfXi1T76TkKrC4Tk4qF/rPN148fsKZtMxYM8/6
dqnRa0oX6CkrVV/px5opdtAiA9p0dUNdwFTcBvX1pcWBJLlkLVg4NVejKTEzhhAyF6N6tTEX0H41
4Ja3d8RmC5Vqbxivq1WzRoMw0UqVI04/NTNjWJnGa+i6NDGwznocAh/qzP9zPaijVnQZToVVl4DR
vNnP2Ua8MvqYcfQNclMnAQce/6soL8fJhG8Zcg1bBtX7rpDtt49HUxCny9vHzWq8T+AuOVGRdkyB
xgQWH5OC4CY7IDb7BzVS3+QgO1K2ol/LsDL6ywBvHZUWgMNscKk70IndFhbbgdHHmjI82f9IqsZX
mBnWFkkyPYH/AqyKPyHaWvXd4ueNKh9hrqgKiB2WBhbUnQaJvpkKS4wnpkZgR1n7aNVVoQ8N+GDn
HitJZA/C3/vwJ+grmn4Xnzzmo3lJ2x4cSsju4GJ/9YSXw5LcTp2L7804/CZNQ5DbPcVQehmnl66Q
8ArxJe4gSqR/kpaU1wIOVG/8JbvZ1xHgTlUtAqEg5r1fIwQC/5SGc8hz7K7dQhL5v60F9eincMW8
CqMfeByfh11RSneb/K/VKCpr8xou4PzI2NAcZ9bC10VBpVJj9bx1ChLQHiRAMEQspNFueo2oUUbQ
pGzo2lfnY+uJiPYNSkSU/Ikv2KtxC9x4nsomSlGVa6qvwAnZzhRnEdy8jUqjQq/ZmG6xT+XyX+DC
bd6b0E3lfvmfT83IDV9b3Wjvt6DbBH181INwo/qXyDAY5i7Yiippvh4Rzd0jfR6z3VYwzi2TNq6L
e4BR7urnBLpl2MGTOUn2VVazHZMOeMMsrFRPq8Xs8qnACG8AIMK0Fa3tQMNHJd1Xb3FBMzzrY/Hj
VGu/qk42HbqFD8UmJjzEkZTC0tvOOqArgAqijyP1WZFliTWH3VR4e/D1jpTkv/FphaJMj1IssAlY
fb2Fl0K55HB0WkR2dzaqDor41ajSRwsn3xqVMbaraL+F4iPtXHQWcDzLiPga4Urdsu6cIvMvP2CG
c7yq/Ehx8MrMrqRFViYjQPGEzsgD9oaHovz4UKX/xo3nFkCMh1JGXSW3kP3wyYYq1e50nJ1Wehkf
4TNzarXEhFbog2/6795q2onDJ2eAQK6K2CWFKwNWHfwVquyuXwYgHv6eCkiuV9BsRmg+Zi1z0e4/
haT9FtEaMAkU0Gwlx/GFh7jQXcfmVrm6dmSMZVMov4TLo+DZhEM0msJsTg7HfIcp//WG14NE0pCW
kULcp4a1PNm5ydhTT5R+rIp+uHbqFN/5SJHCLyeA0NsnoxmN0BTLPiDsD/ZxZnvXNN5CS8ehi5mE
dYVF6KLht/Prg57QnE+NCJPlI8mFzReuwrYxA5KOnlhAtXW5GBJSXPbiWn2oWlyoqGD4ZVsJuv+n
GariD/3uL9R8iaLfYZrGykl5/vr/XH/IO2Z1XHw7U4bN5MCOlKzoIZpXbOueLO4OcJX+KKCzWrE8
Vhqtu/Hqva1nhcHoar3oiEfss1PzzIJOzQvKlsAJssmufrEnyahyCzlVS9ZXpxeMPWhk58DYQyyT
N5BduUrDGg4xrD5LAWX0ZAud4zGVA1tb5XOMjwRiLdufPIQBBAIv6aQ7SRkvAlhiqkfnP3PjJCOO
chbGoB4zQbrkqcaUAOLbayhxBmSwYgDJUW7K5XVgV+IjfNF0XndC72aRoYe+3gCUB2sEWTo766RB
gleV1oRWjedTXX6zr+Bu3YyydAx6RMhq6B+ripCSdirWZVxJv83stKpI/USxzJAgukQl+Qkjp+9q
3uyd9q8ytK441CX7ridAHGDotd3b0wlDN4GHG+doW/KZTdfdEsR0M4vMIBVgPAqY6Qt/Em6yTfH9
Dnqg5Ccc1TosdZW5KufZrPlNU6walKDZghQp3elh0FxU87mYMVeTwudWvO8//2HxmPqtuk1cIglT
/Rujbc3+dyaPVJKHkgVi6RO4H7Mp7ddBZRO4MRLT26fFkJFd6Yb1ni/ExoJRPYAckASIzdvq3jNZ
TRmz6abwyYazO2DQEkNCb+VWs/UoCVNR++g+bcDw8TC4HQV61VVkGZlY4nQXZ6u1gWiqBSSSXkbN
MpQ23BRHT/bsnfhU0P2S2Z08hbP1VHYQdpwYjeP4rTvvvqq9QH88OZ56cJXi984fRi81os4LVBW1
sqGnAZKQZhvJnz4D/3IKxB67gWv2qkiz+EOA4rIOZaDQH2Yvf6inHiTgJ/6H24M+tZPE5MKzAuOD
Ktkme5C/UYQB7Xrut8v5yvjZtvSLSQF923K1MbYGx95J/s3oGl4+VMOm9E5sg/2DvTSmkSGE8uKQ
SO09y48QPd/gl5HdYIS/gHo9hBMWCJ5hpBggSmDuG7sqm+HxWf2gf765h/Y+Gk9LIbO5/vtfQU50
SdM4VWJYvHXOmWcQZ6Q+Pebwd6osgxuoWrYw+WKZ0RGka18U2nWASLr6RhvtjNQWg47Vd89Bn1dc
TpXAM3muEFAbGPKQlcDfgTiEBOAukzOtToePU9OMaa4PvYN3e2KmcQc5Tgm7VOH+v3HMPsDZoTBh
dO1rhtAWFQbogFxe4CVA51Itn18EWu+/bK/gZTEwUrVDn/SvqMIfPsBdL6EoAV4d/5bkkbeYcJJE
biQ1/kfJAatDfMd6B2N5AgxkmanzIzStr6Swx2lvhDId84yvzUtwh/4Krc8tttRDDDhxXIMSjtQI
yGVJ6+0PU7mOHMRH9O4AzGR/ucvvmwI3nwbf9WkCM0IKZnnRl26NdQocxnhdWnpoKIRXivwpx+rf
nPUFKRr/M41RtaF16SmXAa931w6UHrstVxQfIZv7GL4BUP7WIK30Wqc5TCaaYDA69BiMpeuYA0Oe
+n/zygYg6pRLEqGhZODUyZyKgrcRHOcUMNc9yJy7Ftxk8eyhECtmiDYWY6l54GwOzdybS397UPQm
6B43TNDZ+g5wFy+ePUWGxlUhsOFFY8duoAF5K6yL5PMUznS0FefiNJTYv2WNglPqKcFb5eqawWEg
IOSKkk8pDvvD24VeSU/ODYcvTAXC8mGq05CNUn5QXiQ1tctFgOKFmfe2HjddQVlL4pcXYqgmsxKu
wK/wlDCYfouNf8SSMZPZ4cR0ACeTmLoCeyrUbtsACY+kNVRfiEBlYCvfazGIUQZkglJij/zInMld
HBNPglxrpywyXGsL5rqKzV2qa5uYvBMLVKTjba5eSCc7sfm1/T9aoTLenWiQOTxUQJedcvt3HOiq
8SBslbwHTOF6Uhc1RAmM6fL7APwTPcqFTWrrRiOQzeiyKYEDBNltR72G1GtUNek45gwUiEmH4crl
RaYrGw+6dy+I+PXIlg9wCK2j0r6+7/wLobUXFYIrJdOve5nkufCW8EshmFQIcQyvsAKNr3YJ4jdE
JSd6Q6GziWAJRRw/lnD++0Vu/KRRXdtTxk3IoCp1Uktj1CJyXmr6lAl6Ddi7XfLctsgw3WtVST8a
BMQU+vrmcASiHwh53zawCreZNZAwwOY4+YLks6mKOBux2NSjxOV3JrJeDhpvBziT5JK/A2qKHlRw
zkSNFotVq11xX04sCATFuZsXn6jaus13E9+QN2K7n4coB2d4978QrP05yGD9jRW52kMI5Gol+50i
SnntjCdgBb1KDlKiyJ1v99BtfyBZ9eTUYaz3NyiWvMLnbQa2URStyuK9U/rgrMMToXF9NvlBhVEf
lzXC8ZkuZHWYy8gtEKGlAYRW1AT0oVInpg/6LledWHC29+g2uDa2yEq/zbcGqpsvpatnT05U9vg7
N4L/HiPBwGpfzekMC2Btu3gJd+CVokOpUABCQs7mcrbFcoGttggBcx3vkM4hGcxBdG8pwkFOB0Hp
yxW30yGDsDYV0xHfx2CZlqz7Kqficd8XjN9inhb358zJ5PgN8cbDDwnsL1O1R3hzGc3NV7tXQvtW
qV53V1xeygDahJEb83ywsffl9PhPS+3PlrCuRo0C4PhMYDZXQ72NHbfxMODCCX6tfgNT0dR1kXBC
LGaZaDh9FKLOOXjcxHTmrTXGSPJgK162rmlntteYVUbLDzYQJMyEfqU7PSifYFb1pwJb8RDBqTA1
96ttd18JcJrr/z9k/AQAqGQSXOcmaaSTyKFOypAnzzIZwsZbzlimudnb9wdXi28pE76+hxoMFucs
A+sBqfCjUlsSJzWaNThY9Z+jQcvzr+aKwXwzSBobA5Mf6S4S0oy3j7DdgiRQETOTXiIRG/qu5Ict
/MtQBGidTspMypLLpiodtyD4s0iEZT7Smz8u9BQmgJhifN2DGFG0WAFQYYhDzPoG3L8CWmNNOQVa
tUQBulBcWQ93u3Cnz+GJL4rkGR2ouXcKRPxwCCmOr2MLk0pPtOOvTodGUqGCEt28X8r9VQ0k6i2K
a4NlIgE4t1XJ89cZSE9FgB+MhNMV57tZBispIG0mV534nSQvt7TIltRIsZDSyKdx/0TPdLfqsZ45
FXkYhmacLo0pPmkiCW3oaF65bW2+XBP0rdZgBrt0oj4k8u2ywewFNhAPejwJNU79QdNSeK6eDzb1
YvhWN7eGalNYnEWO/qrsZ4MsjXusq8ws892zX/iq5KJ5MPYlSoD58FGuq2SxLj7U/mh4aZgPRys0
MYU2wZprvN//y/YG+326gXj8y8WvtC0yI8vPi5qAtXWrKZWixmaDd0myEonVUhdkNwQsqK93ra40
y0oYsG1ZcIS4q2DF0TmJ41Trlu+Wo0qe3FzFRKQAfenUGmE0lu/yeaUK20e9fi43OZPGMAWOIqN9
cGeymrQ+FBzsRIQhdar1uC6gzywRfaKf4SOzlF02Mai8DzDjrZ7VzFsYGDn2R620+tNKY9Q/IuN3
OSVDpiJsUx2qjdArVOL7VeTN+GGInOk4rwmgg7cRwZMhYG8xyuizpUiZtzTN6aIKqzOtYnmKVNQ3
T22ellxcv9joASumTPoknC4WBJVAXwMFDPoKvBoGeNIs2phH2UMqUnPf7M3ZnJmHxU7nRJ6IFYxc
wOhROgRa2RzCRTj6SqIjrOM+7bj7+6TwjwH8NcDGlfs6J0TveYpJoG5YLi2tpaCLLK+nlk+GYAyk
Nxb9F1YD+zdauXMo2+5FSWeZn3vpBIL/XfcyMEn6jdq1LoDQ4DlWwmDMXUwOBIstQBTOESDpjlin
2Hlod0jQliCqBKePG9A9TJIMdEqyCi2+dS1vzLbmf6tD6ghtGrYocJt+GtXIfnGhdMpwidapp21v
LUw3XfEWy+emjFIyQsjADtdpxedQ3+YcNA7EE9iloPGh1noO07Yic7vAT5Ve4qYsYY9Slqjeu7Wb
lRE3VqGiFKRDmpMwrCO3OwhIodY2BFkmenw2S4h5hYAyqDFSAIu8k0cA8EaiOaWzBEg02qNwEZWH
UwCZpqoj7twkb2SaUFY/wuZorskcpQHk1YUNByVuMXAfjPyJ26vDDPxOHVt989AAln4TlfyPE+Te
Y+V4c2n1XqzbRTdv951oWRe9Gl2SdM0bJ96D9mWtD97NSMtM5GdmG6v/Ku8qqdaQStne8sH54x7U
4aNIEO5ZPHvO6Ze0wUdEyghTSLFtO287w9Qrlx9c2gytgo+o10OS2nB/pvNRM5YrACTp+S4jBYTg
9/fEVCioUj1+d5FFJbv8EcN8plNvytOeOOw4GVeM5ZErfE6LlaJegzGuPamMzi5beFJk1yxI8pud
tlWTJT3LSuj4iz1UoeB17lveE3nAzYgLJNtC+zDUZERXNcx3Zp8f5GXrRt+b5C0f6ljpjhTRGduC
7o6WqrGxSwEFtTQ1KZ1PRrvZ7EEbeTaAuhLrDy2IZu/NiBeY9hRLR2vesn13+k46DkbNl1o5kVYQ
ki1+ZqQPxtsIy5heyk1jmS6WMGCfOVwnAC7CI61rJTcx0/WLEFrAmcbb6kDBRme7c7Sm9EBYyUQl
2yXhIlRz9qMrLBGi5OxQSsp7boghzxZ2aOISYXHvELH+EcRHHFuTsAnY2dNpg1+0r08c7xiGOWpv
w9P1qkMLJ6yhD0sdWLCkeJQSJRekWL5SD+B/amjx3FZWZQRRbPIna3EAB+Gdcqw0+24niuolB9Jb
rBqHVbs3o6ad/xr0ogm2xqzgq59ZFwzLhqZOtfPSqoeBGnOf4heVrk3k3a8rnj2uhqIXUbr2NJOG
g0yT+PP5XeVlMZ3ZoQw2M6eCz276aI6gBtC2Y/44Ue1jb/JD5jhJYPuVnrtNuLQfdMxNHocnmCu+
aNEVWt7QXvL4vEGfuM46poUt8e5gelDKMqTfG6Yc6yM7+MdJLXXQKjkVrA2MAS/HyldhaDRKRYvd
BOUWrtHyuUciLu0hu8y3B2xeldzew61Hdzlu4Ajf8yVhwcS28aj7vNGfGEMw/uNMOerHTJeaYUn9
qmQFhET0K31Y+CXxmEUZ5UJlo7eL0xVv5X3Z3j9dCS6ZGv+5qnXrd4+rApFl++U4bK+ufiYNDxpD
tL0xSEAfk+3mxsZvJfMF2pTbhsyTEIXvs7RuwmOShKdOspdIUlOqkPkmU2B6YuhBxHZwTHULsUuH
Ne3XfFNPRUwYgx56UcYGKOiZxI6mMhJ+57j7J/Cl9k4mzZBKOiyeP7OvVyjt75JA5vYk/rFZ8KIV
ZT+02vYFyNlckz95rf6lTAlFemHd0awhNPVi0XcFesuR3ZQ0WJNJBma3BR3lMKDbIGAVs9bbaSBk
8kP5kbQWaeDmK8EHIJUCcQBl6QcudJMOuxic1AbaBJxSRqw/lQGY/RxhYglJMxpuES7v75gQMjvj
QfsZN+zAoVB3Fi3UlQlcix1bLUJtlkaXqjfn4l5XFacHWVgn52mnjoWd8zRpn+WHMBoef26ncxG5
/ejjATYX9j5wb0In+mnP68Z0oQ6Ii8KeBU50K5JYh+WN+O9+Q5+NC+zuf37T5sEgO7FA7elj+Tbm
1sMPvHu6AY2UdvL7n8sjxmVJ/cWa73vhPwZETxhUpm7Mtwd9ZL6ymOcA7dDjDkXLy9Kal1+Ptjbi
Gw/L6roP+sXCyW5Bo+5MYSYxlgqm6PRJy4Kx2XfbHoQbSc4zik/un61DHPp6gYSELguRNc7TtyqS
6TG73Da65rBVTyMERFTrqvateESdO5moCbnm9Bc51m5k8jm8OBblLHBtJ77yM2MWVASh0EkkKMY7
jb7Yd6ME7FoSsZyt5FUfLyx4z1602ksh9cmPTP7qU8gv02XuzCrJiBJ6FaUS9YbylhMM19s+gjJN
NuzCgxHOdJcth/3TCh0rIi55eZIqRI3CxrAOMchqAPraPCd5PLH5JZO46Xtk94IlHhOWEmqaf5fR
iuvHxnPZa6rMXILxdvj7OTt+3c0w13b/Ru3umavowP3BkFlkvwNFxaz+yVv9QIowcX1N6Mya+A0m
VdfQ6FuE7fNzpxniG/mexlukVHUTYmtakMkckCqhYEMn5igs9U1+IJYIPAVYPHvqD8k/rUVBnurf
aB4Q8ytI6pCeQyHR3ggYwdgyq8/3qcJrFRiroCiqWTJAH/MstSzB+uRxurzJYDJevYWnGkDgloSA
gfUE6NvkrhfBk9Yktw4XFMo+U2cVnJNa057bepWe++pUReahH6gtf/aW1K5xXE8UZBrZ/FM/vysR
b1kPed/RIl3GBkRiVLvzuJEg7WHuHVqnJAI9POv1Qj6Y4GO5SzqXHC6fJVnAq/lS0RMRu0uu3kE6
nwrq/zKPCNRA2aqO1sfsE0b4yDsc0iknvI5PbjHZlO+rquely8zS1hiLA1keaiZ4N6lGZegU3vYK
2qcL3jADMUpQZirm3SvEb8NDyx8kz4lOKD9Nh9w8AWPvyvTsKFPEgwzJVEVDyEp7pTjo9J5MNqLR
M90+slOttEiTfzTCUP0gSanU69GFkjSWs0XFFzwjXdNVK3T2T/B+KeA6kHzCnJd58qWblhSrquE8
FfHKaJtjr7lHGkAmi6eUytOOZSKYLVon893LBSFypz8IPKmfs9AknP/MTY6SdcFNGZoKr6B6UHs+
P9J4XdNmThsBF2SR5ww+RzysYwYuoY4qr7Zdo6hZhA+16EC5jF8WYg4BTwVA1WQV/oAGU64cHWUK
+bxOkA0IeWUWaNbj4OFkC0LlJAFTlf2cbXP+d4QnrOIJzh6aqYRTLoD4T1MtNtO4XpKh0UStoskR
egwuGVPV8fsFZrtuwcP8zC6bk0OVk0ZWNNWfdQ22NbsW/4WSGHLAvHML05opFy27/WGvUiHBYlSh
ix1MK0JI3ceJh3Qepan5awlIwN2zodNKDLXCHx9zijbIB2Eo6WoFmpVEiWFVtCVkg3G9DXoLX5US
AbUeEmsjg1UCQ9IfPaRGS9D6Xorf6zHF51PiSpvI0PrYhAyaQe6vymaIV8Czt8dAwkCQbQdUeren
ncEYGD6nEXM9cFwSy/c2KKsD13LIUjGKs1jVWnWlBeuwLt0/WiLul/XLgF7WYBBEFRIPkfqutP4j
jhEwHwdVUbWGyUJ0maWD9U2052L3o4GejpNyFSUZipvBQ5tr5C7Xyy/8y3MXfehEvQD8e5WFsymf
pkAz2OgdLEHbI5NV0TtPcLu+5lOaF/UHdS5Qs9KpqenjANzyCrPPu3z+vFHyjhAamSLxFDeBjy1o
boySLGmVuD+aORHkcz+wOj5y16LXycaLv98C9Z2W9em19LKpJXiBYE3GTiQISAuhFBJCaSp4V+04
gC/zl2xafBqlL/VlDSevXlbX2N4og9JFca04KpP6pkLnWlMlUoi1U7Cp+ED/GuVqNe6Vh3TAzCNB
5lsy+6SlRDpFIY6/IJd5JoUSV7u4bPM7Cg269GsVUpPclWOTT9oifYU6Y4baDi5oBFt1FyWOV5G4
XzOfCM6/PFjiPNJKdjE/rOBZdIzm7zqFvoUQ5wDvtrZB2yp/GYRREFhhS3iftmNGtpd684tftWRm
Gp9XIPNffgElTx9Kmha29z48/qVGJIOHSJneOykkIO4iS607dEXv/PWPX22cLaGhqbbSrzdaxazV
O2rlxJ801oFzBqOhLvoLDGuvEp7++CL5uUKPb9/pAUsFIy7+nJm1PVD5TV7zOBw7mvNizxBpmnf5
lvKJJ8PhPHdS1f0Od5wO4J9Gq2S1+it0pcJIqs/EvQb0bGFpFwbgG6rT3FABAuWj1/I2pDmbqcv1
vA5IGBV6vWDzq7QPryFkF7HqhDzgAAjjhcbYZiS+nl7hMC39nml4qC9Unzhn83vPXxB1Ei1ZG2KH
l1Wuz9FNWFCI8PgcBGbjeiI272fGumVvcjbIZ7B5ruWpfiRXLFcNikOSxtTvmGm0qkevYIQRN/lo
SLwjBMs0TL345N35gz/V8wnKBZHOUv6JC3ZFHL5yzjPA1nu994iEuk7zHsID0FtcXIiLwj9iOyTX
qfE7A//n+SYWSPuFpVHPkg+FOgMn79ASMb/wcVHP4MeV+qFZpHf8Uzpiyv3catFCQPD+z3fK7jIs
5YhSfAePaGLTcEO6uqAi3b8JyIoCxyWLgq8KOUPQGgVOe5QyalBOqhMS5Th0hHi+YSizJOJG1ac3
XJeeVcfUiIp4Trti+rUtsi/kqqqoOYtzFegQCYHkfwzUr7EUyzV9AJ7cI2+6cnoLC7f1x/X3azQU
lKEMrsun9ZXE0y9hzIonNIgVNjNmSV4z12fJCSJbt0mLY3EcEotGQcf4nscEINg41TdfIhiFGajA
ppnho0D8c2JYfrtpqoYioJR5lq8zQDCKT+FE7xX467EaH7ymEHs/Y6nO5Lk7UHUhPxISHaT0r1Ya
LJzGr3Z42uQG+knxvCHds77NmS/IyrCu4rKQcxW+Vs+hDJ4CBWeSe//ORfsaUocUl2b8v5qtvl+Q
Tk6SsjjbO5lLBcZN40VRc67fMKAfgyJxx8dczsT0qI4KbrZBNW5KKIONxH0iG6sTKBdXBF57Jswf
hIV32qlPyNiPtGAryqkII9jbqN5riMDUPXnKpunsVSkoHBVH4vfKKQz2Edsl4G6kb9LttU7lzurU
0AL+jeCf5PdzLWCHw/zUPK5IP6tPav/XmSbZKDObZxjJlARopvfTt7ljk8xyNVbmv2qcoFMDAyvr
Ej5xgJ4qklpDTa2GExTzJpC5buZmuJdGJa80yeS8AuCaua2MrY5jU2hE0LLx41aqTM/modpxoSMD
LTwJIpOZrwDCYLOWzaA+KLvh6+LH4KPQaZ5tMl8pMMKjcILXxz9kEX8Ah2F3lASwSbcT0FShL/Iu
mB5/zd1xyIi7Vhhjk75Ee0ilpZmfepu3WOuIgcup7iaYgQ4OT+60Q8x/Ij+o3TKDweD/EPK66wsr
CVEXyzZXrDT+8gLHkzuysBhSvxEU66/YTVHVb+wDvn0B/SYYJhdaBPkrsVy4FkzvHqcmedivhN6Y
jNgS4X96GYbtawtPRzKY3bcJoYTuwpbvM1+t/m9Vb2Zhg4xIzzbTTGvqKu76YW5+Cw0QU7/LVWhA
UkbZ+r4KwtOA1v0s8dFSHwRZoQGENIAR+/xZSGrnQ/1Vew5RUfMAA/6hiPJUSre3H5iyDODyY7Kw
XyCHieff7aZZMojpkgJY2UwbAc7mXmnjq/ny763bhyvmEIFphSFkKtQGKED8FmpzSoHcAeDbd/U1
Jx/qdJb2YNW4JUWiBYwy6lcO/N9t4+/rMsuIROVMX3L50KPcL/syUwbQDckL/0wqjPybyHUQx8yA
Qd9naTsO30FaiV6f4e8ieSpIl5vrD5QzrMGRFjOaAp8aIMCLB2EEBjuSrl7fI/Ku6/zt8yKSVy4O
BVvgQcoTDWQKELpEj8rqVBASk9VakPlLukGCZAKxIhDJBpJBmErDKEyzfGS9g0O5pol2ZFCcKmR+
Yqk1fmJ16vyRfqi0VKsJ77i/XCeaLx/T4H6OAKviaQ52k+tVD6ZgX+lIusPXQkhZJ2l7B5I8E5ST
HOQGzl88BwJgCzskiIfeuYdyQ4Xtqu9Y0AzmWjuLGpNvQP2YXgnSnFCoc+PZwOXcRei2+51dCsCo
hVamVKTlRw0pk4lj5NoDUYG5pbx/kDBxJhaYAjfkHzHjWJyXepHzHdMw/5fmX0fxPF6Nt5jLPaZl
p+QAGJYjcrzbGVJqvd2ycU6P2wBo5oTrEXqgn2GeSUSrvL9/Ma8RtiOKBCKcwnJqPyn12ISZOsHX
kqJcE8znnFY8dEBMM1YBP16jTa9y8tElrvyGAUZD4/he0tK+IbvxsXiggCaPqvyKcxkyE3QIPOhR
hIkeaTYGomE3GWwwepJfB3DTL/ybti5TU7xtgwGOKvHafRL9ldG4QT57OjFmkfjAuox0Mw/dVeie
7fqKSMURPW7F3vQgBjmI2a1Svy1PIqWHWsZsw0iFt7JjMv+1IErMOtDABJmgmow6Z/wLxqZ65YvR
eX84oTHJHfpCblD8WgnNSoRzfAgLB3TJF2owqEU5U5zFiGlImgHH4RnLrsppPLhzqJgFaTwj4rI5
imjYHUFei9Yj86c4kzHR0pHPLVmX1hTcXbtITcPOxr3BloxucAlzwt0SS4o93mpgyegwdCY+MWMi
RIiVKnVB30I9PGm+6mbOqqJqek1UPh4YQIRhMkS0gmIk6rdIy1qbA/Naxs46U6GEl3OSDTrMfo7I
MMOU5S+gBO7T+/4uxjoY+As7aS7iOy77UYNo4y6atFjcB3cAjSbSYi/yOJheQAmEAyhupb59WUqj
UCbAUUWjK8RDCdARb2eiAtq7g5uZprBZyCrJ/pEBAvOppVbDurUvlk9XsLslLyxzz9taxDgcUfle
PfKP49KzCig808KkHcN9X6+vc6z41XQzW6wbH3Jl0VTV8NVNvg27LLTR24opFEyJhfJ7iEZzqShG
Wa+H85CB0gtEslKXCqcmGLyx/2YnHiza0q3RhD7H9BT7h0J+6QrxLvrdrxKSqUL4HjSh9BO8L3Ih
HjlxnPHMgS+twI5kPdnmnRAF7BNDdgAZOgEHICTmYu6SlSl5Dw1LJaZIiIA7RJUCoXf06DVht8dG
v0tzt3t1QV1hLzfWJKGuyLYjtn6QVpmLeZl35+VaKyNetdQgUaEWUVUGFBaQCIYvQ8IoHUaO+iqY
OMBYKxyw+lCo/v6Q/D+W1EAX1c4suNvo5cCi4KHR7yJz3WDtrhB7W0s5QIdxs7fZuc4g/F2U7M3w
wh8wd7AUAPvsdsH5xImYIu4+DypYq0oPj3JfkrT3QlDlQuOCJwfR27yvA3f2JqwdnZF+0iwx9A8+
Am9E+yA0giKxkGBDXLBKwk9pTSobSbHSa7KV7KVEncS3InRXgcmmBRIiWSnAzuKO0bw9j9Bb3A2G
UhzVNRwmRklsNl5sh6vFf1w8SghgSL8xxkmNy+TQoYNOpGZFe7RVhnJJ1vx2eKF0yHD7J8iB6oLA
5Cer16sQbUuWIYmT2Kq+dD5CmImvxFye3LbGqffzzGjHEjFESZGIc4dc398bNcGAWjR7KU7+OVJO
S+axHsSSMEEa7TLXT/Xv0otwW8yoImNS23nzeud0jNZB5GtHwi7g0B3W4eAGcwxxpEWIlV/KV5tZ
+1FNTk52i7yE/h8mjwuCbnRziIvHdIE27xXpPlwSk7bzsQY35ZDH8LxPI7AmbM3GnulSCR5hjBYj
knjlOfZTCr1ZV4L8BdLeZ5vEMrQgMwuVIUuhk06wKbvh/0xWKh/j5npwv4e4J6o/hTcMDQOLjvEq
wWvyeihJmiFhC5jQj7Vg7QrkpsAsne3zves1EmiKZEGSfTgYBHgmfVTJs46o/6/luoSmo377Gbt0
Qkdc9cj76oiWJOtWHdPocjFcSkTeDbCUBv0NiAX9pAf4Q4sJt4s8obeXglMzdSHGDd0LFUV4EzP2
MC8sYsUzVKwxonooFd5SO+mx7eqSajxhKaEzggIY+/LWuCy6nFdDBpMN4jpqbKSGzLQNmOldNyH7
mMdu9xyr2AXWD7uk9vhEJHIsfdfoIIh71rcjjgQUU6fp7Bc7P8PmJfen5h2ql3RYO8d3kDZp1UEu
LWNgFkC589X5tcchgUAe//MCRp0V6bnfbKMU5r0dEWOLGYSrEGC4NyhwES+p2LZjpBLlEM70TaLA
ezLn5Sx9f14Bs4nq9rR1ighTpnWPPTKQsQVS8K7XgZ+/V1kaiQPr2RbNzt7446IoT+SKnTzZLY4a
NebVCP2C6+2e+U8+vwz615d4wkTEksNveTFxBoW9VRpFQFOJ/5kjkH4L6fxFeJoT2GXS0RrYOrzz
HGe55ZB9kQk0TKg6yYmmqeKene58bzSHcpnqVzH27jfjbKNTzHU82atgCFGTgtmVAY5n1u9HfW34
dTnSTqAklIASVlIVSOnPBhyxUQIIxMvY+yz7r6uB1tm7xwH6knVaxnf2cRo2vag2Zxi/hLGU0tbU
SazwqpQHuwSZVd/+l/fTXagr3YOVUmxdnp4CbsJasjHtCdmBnRPnkiLCnj3uEWV/ShENkCv0v1K5
I5JoAbkpsAeDTZg9Hge30/qTac0n5XdebCEDF1Z0iCPl/3eMwXN75HchA8HvNDwmz2+tE+96upRS
QEYfzN7vScasVmLgs+UmzdwuzNTkWg+UHZwo+CNSVDLr7zLKiaQp6NGGuvTU7lhGEXcUXao5uTBb
44rNh1YA7/JnR4GjsM62oi4Q4jx1KadFBTF3Fhpb7ketr3xB54+CnxCP+tVxqCPz3C1ox5POQhvV
vQWKWweZ5nu60VMZiIIqzrkjfc9dgmiGJuk2i/Vtpc1CETpGmae7AsKS9pJttFvQZI0gIHgdQmDw
d10ulfhGClMFwULE1k761+16DSMXEExmh82BIw7cilxYXnqUMjpt7xE7on+8g8rDCS2nQ8tWll7l
JBhpqcC2bP84t8Gpl3ATydTgxJEtW3klZZLfw6OfXddIgz5YrFf2182sRBBCGjw+en+z8y30STDn
NQN1sBgapEpjt0sD9YkR2fbp/zdu6ocQPY68v5TW/R5i8h2hnG6I6P5dj29CFJU0fTRvfXsYcHzM
iylykxqjf8+FvGMppIbL5CPlYFGHro3gnkGMBuCUIIUAVwzL5YwX0x2gY8Bp6fhGXFOIVbTkEU+t
qE070diXkWiQnOZdRLpe+A4tCkIY4sBkBrZo7BNe2o7N/FVTryqkAqfhJVCQxKJHnXFf3DAbDcQz
Kunt3BgT596RZO9ewLNiGmzdKt0hyENtYRdqVa65v2LjG4x/4C8m5yAG5+JncAzpxXOfY6KOuifq
GU7KSLR+V4D915/N7f5Gl2ROvyo29jFq6kCz4XFuPNC6qI23SSXo51FOe7J6staKBdJglIu0Tox8
RjFrClRJ0P5BECmtDnOgMO3noy6KxqsogtZo4o55WtNXLD0NV0YSbibS5FnuJEZSlVltKHC4XgFN
GwjTjvUhb6O4ml2nMF4Vgjry4N+WjD+u2hCtTnmDlf8Eic2YyK9qXHEG9qAKEJP/q9823XK4Ar3I
jwGQPSzg6ATHLAJ+pFD3X8FmEz9LS7E5+zTMVh6hr3xFvfzPR6TgyJi799+s+expaGHvdBrhKxhz
kOEv9ZP5/W4gXLy966vYpZJPHNCom9oGUnn00OpbArljWtfbBu6aZr7jJI47vW3zyDI8jxPth1hf
efvUhRe5mSkgC2VG89O9L0nLYZaLgrP6JCpeFDSHbvNFZM6lN1kHY34+74rXXGJ0QpJ1jB+ZbDSr
aD2CfzzgJoFyKeb+nsUKzRfU8PiVhucx3LTXHuTxhbEHHPwi/K3pgBIqD0AxZEGtrbDD4BXEd4V1
LpL7AeUGZrKnAgSIi5i8Vvv2AjxpS7bzNH+I74KoTjPidZw3DkFFrIBEndspDaw+BIS/VLQLsMxZ
Om7ePp9Q/71XB3cuyIE6BUIJ/bu5Ujd4KaS6O9Gor1JeweoASVo7tyMr3HHumyrN+vOrHNu2Z1L7
K3QdJfePGXa21Jr/qdvHOZRqptt+lopHLyOEwvmrczk9n74LVlP+IkMa25SaC1X6WhlVT/bsS6VM
mxAPXtP6BRCi4FTyHdpxZ5M/K7m7Y1/QF54o0CW/BArinU/WSTcAglqdsVbmya3loIWDL0kAPrMC
mVlsa3ZCglG4PV0zQ28xfD+FsaZmon+jkZW6fA/nWCeUqJK4u9wTc8ZO0SnlsgQ8DXLqJDzToUTq
A5wuGX6zI1xdU8dwTpGnKXfvZ/rpQxI/tqkkBt7A3b+34nJXBbg9dGDvR+7Uh83BgJOfkpW7GDUx
KaCZk9xUQtnGzlz/lP/YgGbIEkGrJ4UuinICvEugmmpQ3lrp0hsQw/16giuHeWezPOKP2kyF3XPK
n3u389x9yvQDj2zjbxs+RMU6KjBk1Qelgs+1LqFAxzrU7I8/InDGA7/eSyVZINoISC9tw4oaxPk+
NMsv+jdsuPFgLzleTsIu+uOgUZ5lSq0M62hXEgfLPzze+0QygB6zpkG+3ahvMTEKcvgBxlv8M1iM
ue4YXsd+/rQvu+s7lCS7cGhc4mg3zWOAeWZmt9mBgCBOxU78DUOuD22Ha2FLKjFjYnecY5zwbS2d
vQixMsdYrG4rEuHzky+ljYuOEVVhlYMPGQ1BxOJqoR4GacFO6DY+Hs+oU74sITR36mqm7MG3k5BT
MvXtenHmuNXpoVFjEouVVqiykh+o3I+biBWyxVyF21AfiPhb+uelqqjmvYVacy2jStANjCFeSLnE
F8aG8yCEN+ep+teJF0SNPcLd/henFrHEZsj2/Rl4JVlYrwGyvKHe/FFYVToCSAuxABQemv2nOjXP
tUbtknUZCtkCcP18tlP+MYdo5mZexu9tPyAG9z4pFjOYtzFhEpzGCcq9jxb8h/ezbLxrS8ENvkbX
wkuPGGiehYLxrxloVCi//7VZOh416hXaqNmfKRsVbM2b782DWBEy4D5PfiyvARJATitJd9kbasbS
x3d57OruWEhiI9RgUjlX/5eAr7FReKq4iUbS1qXZm3bLra3XKwufuUJ6rSEuvWYnLa6J6E6dPlqt
kjadxXQeL1HPoC8cwNl7i8zzG3bakRnLnc6/1YuxT9WIBg4opK5TMXilL9W8ckfcMGdjkq6mDDDn
WfCSA94iHUWOE1UqNXGg6NoJqBjSzTuwkIVmB2V9Xhr/mQVWvNY4MJnHkb9LabtA4/da6/1NTS2Z
aeFgUrCeu9ZrAbtyoQWGv7ZEnK8EWjw13uhnRZlzGnofdkk39l+lvL7dsRHdQSOPWcO3LXs3LQz7
W/Mb4nuEdNeDmhfi3YqYx/98sHvjaHc7CgfuxQzlXRMHJHbPEFgOKHTeBGA8fuhNKHcGQZ9mK0bF
ZRH3uqcKLp/DF3pAFMSih5qfrDeYmHQAMXb+fXR8477jDkHg1PC0iDqyOpl815+g1zYuq1t29DIm
A+Vk+nn0X7KKD0UFj9RCSJnQbA2zb2t4tJmWN3l0ZVYJ3LLqPK8XgElt1eaO7HrmAKeD5o88l94U
XgRxPTgQvCheE2HMdsDO2HtQi662S5b/EP7BP5dVa+7Lu9jvVo+bXJC8vJRRKlmc8f8I2uxBYF4O
N4orxPMPx0wyMShthCk+a+4YHFJZZiWJJpHfjs+LTX23XnvBT4CsSEtEHtpNS+bDRK+8Rx1CCa1p
4jh5wziWCxee6Hx5p127p2h2n1RUIrcuu+8+KaMzkbYfsGho1QiQjWV4q9fFkfYxWit5ATIl+xe4
UddBZ7eu82aPVABViHCBIOqUsmgx9QrB2qpTJktUVb4f6x/kd/a3gRXta8V127fz0gy72Fg2M3tA
BOwuCU3domcDDhyOaYBNL2uE+zq+xd98AuLWChLkobMli+2E3Ky82uWsa+vLxuGrwuZoG+CG2+wG
0Fjsj7gCtwsIKDZUHwl92fF1J3qntZgdqquF0fAA4l4COZRJM71OlDD6JDrsQe/KIvHCYiy4Q/JD
4+/iui2xrmlfIH6gR9lRTnVIZnkaErsIafTPu46kcjzLX6BZ/hctlaaGElWjLTJFCofFOXh4zdMV
vQxc91OZ+aH95oHIadfAMogou2ojrMbnK1pblossR6aJ9CkDxBVhBRtYlDBA0Eh1vJK/Xx7CrxCv
N7y4dMc0FJFdU6uVXBBI3D+alZUV/LArkFc6SPyyJpVP6BaJWkKerDOGVmrIboleRwRqafEHVciL
3ZO/mWz42GPDu0BX6WXb+GRmZ4Jm+ud1zeUZC9pcBo6HtXwzD2KmrUhm1u+SknPpqDH+Ah9D6Agu
az73AWh0XiVHPgjHby3Pa6KmvBoXve43Lplx181Iy012XFVF1/aavthJlNXuFTfwBGJM1EAdCgSr
1oBZ/sv0KrIeByyXJJdSPElOAXJn7oduEqFuiIkoK049ZiEPu4AfVVskefZHFkzoOsZkD1EWeEDm
F16vng/CfX7ZDqKYo04SfRAW6wgE5aN/RF5MEF8Tkf4dvNWUP3SpIq1NAdkghbctkvNavPazAQGh
yMYErAfh4b3JpwCL/bxKyGBaZ8W9jbbCHLtbLPPCilm3prd+erDpBFGsIXIcv0SVnEcD6qcU10xr
gxtR5A1xSquM/gcvwarTC/6EkTvsWfCNaKHAdagWLNCN1ebcP4b6DPwUJdB9dlYsMLFDbIZEfFCW
6JjXllu1PllXlE33o5gjI0oGUVHq7FAP13qwX5Q4UbXmLy6nyLh7eTgeTBDaazkyLkH9rPWkW3ar
SVxoJp1k5RusynGBsqYfeXcBadBobwzEo98s6eenVNUJ2viH0ZW4+KH0DpFlBXi+TtZyk/xsF9iP
8/nKQtN0hfPLKPl0mmPJxLBKs7Z/HnUOJ6R7Nm1oL+dPhfw01He93sgrba4ZVb4F4Oc79ezGcyeg
fw81VH4G3W+1jBAuhWHBIxxawJaw6ZmarettzqriFTf/eBWRaWQPmcHzPr7HTb1NmR5Ad6PJIkAy
LZoeFLKPknD3gZ3EmWgnSUSFpQ0gEUSRjDT1g/Wf9dJw6k1BKpi5ue/zcWjk+fxh2tqKxxp3qtS6
dhGjVe/ndoWTYCkIzHFOT5UZAQ/K0Vk05QvVuJc6d0OGUMCnA/qqH6tFi5uOw8+TD8+oBoY8t6+1
YhtjVjS0rSmifusUKIAUQP0DOF9IhZXxSrEb1F/WvrgD5YNDw/FI0DyZJcm31UNYiRp+clz/6qBT
4//Vv2TLD4b9BmIr2MQNoNNB+kKU472v7C36G2fzJsuWbRu+d3I4rXi3AIXIgYnWcNMWilIY7IhV
bfT0aoDU2WiNkqEPNDyqxpc8QIgYbXemzwh+jIMVpSXlER6awmDOWTcvniJ2zscBdovwwUpNVsQL
eGadIVTwqhelLqS3v5bPAoULGQKfn1sV1yPLkUPOhhbd+CaMJNiQQlCETw7smQUEPziGN/D4I4IJ
uyCedzdQS6WHnBdCaxFYUg7EzVq0SjHN+FoSIkGVUzXOb2YqumwKqq9L49LvAe8umt2qimdOm5P9
Nf+aQZObgrJZsFzkpG7V1x1x4TE+f4Lv1DD0VTV484rJYsZwGYVIVA/4FFI6X6smlzAimaDwwZcx
Ti1bBBMxH3rHIra3OBKO/fghcPMeSnKR8gYcsJ8lWOmpMKl04KiB/4Q6oBscAXI1XF6c7MAK2FE1
2ZtVfLLgvE+5ixobGdCcKkqWhkq1o8L2X2GlOtkEl9XyHKBNp1BdB+b8bQ2CFjV1gK/8eCgUvYjR
7rI9h03Usa9nBk5fMHKDKYU56QmjwE5DiA9GvF5xLXqS94/8ljJsyW7xQ+cR8k9BRbcKV7ccZaX5
IcPtUabp1xIV4mv0cCJVkkwRE60DTB5fl0rPu/IVcA9SEsw28l5dh/3q6SoiSbAYMCiBaX5jSz4f
o9efyqT9zIQ1+TjqnkWuTApXUh87QMFPS56lcY2cwdaU22fRpSzLdAhfr5k+iSauiZsdofvEAHQ/
54t0PfQDWq7azcka4PYNcUhEdXd7kJrcWyknx8T5zPxPf+2FLpn/vmXuEqLRBazXWyjxUF3AzLLQ
UQYTK+T9/EJGHuqwRhG5t4PIxPiQdzaO81XvOxrXkKwVgGoo46JTbQHEzfYUtGQMI4eMRw6ytlM+
bEjCGDQXn8+6JlhrMipRsTkAexHkuvRrbKkmWtMimuqbLWC1ARxXiJtqe3bySWNEFAtsIUo3DXd9
rYW6wNepdPw2/hZBhsRWJ6ZnUcSj34GFX0XyaUxLD19vg2kNcjac0FHBWJeC8FjEqSxOUnCucoOT
VsQqFESfrPCOMPCsyxncigmsud42twa1qrb6S6FKs/UVlCizi9j18CU04yx0R3PvhM4Jg4P0l6JH
qJ8p28N+FkWdEd6rJlkn36Z4C5p9yjx35WFkN5zalS8KT6WteDB9syLKlBWHwSs9ToNfHIv3AyAo
tPDUFr2zADlMcQpBPvENpVjs/J9wmOV3hFSdzYwF5NNoSqL4Sypa+UVMppy+yMVGWRfAmoOs/IHz
ONNnRRMLn0b2Ri0lve11UdAtiNBtsrZhd3S7eviXXxi7KpS6cyQd0uiKi2DgcMx9JPLKPyeIqCZA
XFSyAHctt3mw0rFjCobJC5Y5OYN/lF7pw6FeHyuxWGDq9FvGMG4WWLoqHE1ud1rEN3X/pqJOiMiD
Q2Gp/0B9o8wXtIj65zaOiDt+zc/rmTKkHcJ4J4pXMzrHwudHZv3/V2HpdeTDxdBH2nwDYlX8AXwl
iOzpVdBLH/pkIjlu4V5WqlYj5zcbasVb8H/t8luyVk0gFp1a3RYU370sKBtODMZvfvOkow0NdJHZ
PiDfq4x3L+PuuyRSnhL2hHo+9ye00e8QRuVa6ThVHSE9UWF1fEFP4c2c3fM68fSotJ/n8O7zIFHu
kJHsSPNQmNmTDa2Oxs6MWcVr7WTwcFb63ixYltaRFOfjuSXl+SoDPJOZsS1rRudSjbmSz+cSb4sM
WxZw7fIx2TL6idy0TDglX0KlEH2tzO5cav7G6qDf3gR0RGh9XH5Thv/JUDZkZcVwsKstF72T5zUF
4RcFPJ3JC428PgWqR+yhg6Wt2lCqlDuw7beWX5eSmXoWFYpygBEKOvIVgqWK8S9bTaDgs4CML+wF
7gco0R9N4fEZ6FtTqEMSBYYu/cCOVgD5hoTNmBICfK0Xw6kH529sZN2d59UBoBMNMuoGsSFTxkow
Y2LAM0eg8IsW9D2GnGs5WarXpe6uqohgom7U8golD6Cvj6SYtuMNlajXCHmLV9EHXPG4Sf09dlB9
Ef2T2eWgQ5vDNZfd7u1n48do78PSjpOYPZVEte4TvFkWkbHTzvsh8btXAOWZVtHjpl2XdKacxlvS
EhgofQaAowhXqqT+sl1SUO60x8M7kuML/y1bbmGQIWN5h+OCGzYxiVLN25nIsuzdp/DE1skbnYQX
4s3EB3BMqwb5u+6s1ILNuYaEnV+Kttj0HQtbep8G8eAFiBZwxFQtPh5yuOZNUzmoGxKCarOjXxUJ
/+8RkGPxr9ICd6oJbMOdlSffGeI6jYo3k3YGMWg0aSAbHvA3mQmpEJLZ/OAPZcaVuuBn2jfR7sfw
kKesJ1RDDgeFy1v0+i/t//HgZKsXZrDj4yatNt0zu8lyxlYS+UugeAv4ktepy804eMxndOxIVPHh
4T00YL/1DVZO8S8hcblbEmVpjr+auSaCqC/TUGftXjMslZUK37zmkuMpEGU/YBpmXE2BEWQBXSlj
Wv/AWvx6R8EkKF9+sO7dpLAr+FR2AatJoTgFR4UQKiTYNZLWVpTOcdBTFqSFKnwOU717eHE53HmI
XhSPovmykXJZ1/pRLookJNdM2XEzKzL76DQhsiWrWOuNlaDCdeRcW4UX0PsbIzzVOP0RlVp1S3+Y
4CHDUZou9mPiFQXmK3hBLJs5VFlGzksegXdng6sUKYODYpQNkxoo1T2GZDLPe86PVMhyeN2MnI5j
OwkmN+AYV5xao7UH5HNFdENEe1uQQWZYE8HOQUr0Ai3Yzxab0CVbWdWbPCHGFiwCU2tPeF7/U52a
CtQvVyPLRL1KaaBFwmvYNcwCeXDxcSQWZmkJ242C8owRT6OAo4Zm7YX8D4aUs+5vcsX5J9xn0buT
s0IocecZoG2grkhENGg5XXjYYsfAGusUjmtDk6ZpFDQbz7Bf6qtG/Z/rdNjQAyLWLCLY3gLAobYL
QLDr9aW/BfTV9K2/di2BeyezCwCCvAn53Y14XTKvkTwF8gi5MbzEbTtJFSckjLpY0qdPyAWJc1QV
jJYJ55AMakletrgdGwkxxhDV0Y5rskgkLqa71FWLOs4I2tdXrsMYD/zC7f1e6j3dN5GW114XDr1c
EKHADidW0T90hg249x432ZaEFW3UYj/yzrH57ZTnQdZzhMycYsEuEj7REovZA/D32tEDqgkdFaJr
7piTYutvlVv75Ks/XDr3ajResqJIziz+yY1jqLjCqTNBBSN6VjYQAMB/Qf+FBWKlwhtkcz2gp3xe
HmyLPuGWEOYjZ9YtK3YYFAo+oByGrb861/3ye8gpQc9+7FkKdxbbkMr8YP9j89piPFJIF1DQIhos
SZ8fN4bbqI1gSv0lB+Vx1/tcr5y7+zkZ9PDrsht/DogJbFpfhFDbYCCLk55YnP1JwQQc10rc4JTo
ald1F1dEy0utkqZObgmI8pGyZp8EA47c2YyGTUxAauhR5sshNVHt2SuDfzWEpFPCNKZe2or6RgYF
yKwQvzooXw6WZXzIVygBjNomO7lpQjLesTqOPdgErH3OysILcBZW3hY9APGZMj/kq2F3hNR6R3g+
TUxJcNgcYx9edNkzdeoiPhY5TPrsU3dY0BV7dURCofO2NG0J4WMjH1DCFv43t9/e7GgD2RjcPcXW
NP5obdLZyVJC1eHKJzogK2gH5iyfGlI7iN0WXsFbXLcrX0nAc0WNB0jWqRRQ4xwSV4Z3FBkO3Wu8
cen8pVSBbx8jaIbzIicPldep1DCMLAAF9yq/3jBC8OU98szvphb50ypztxqAtQtCsUo3r9GguYX6
B5j2NSQjheAeldCeRXObRgvwOfuvW264LUq33GTLMywM8df83+ua7yqCnAq7gZHd8OIljnI8Ft6R
3No+fgkQzR625aWKDRjyoRewfEkbNk8Kx8qMpCDso8awyrRq13TkcWveTGTap4wQkCEqASUGXdfn
q6Yu1oshxebkemGjXsKcBDtcX73e4KUHpj7tNoPTvsXlQJ8k9ZHnSS499Mwzrex2025VotfzBCTE
0WPMzmEE4p9s6B4kDL4SDhXqyML9eLBO/MYv73rY9lREgOucQPQSh67m0X21D3TwzougJxSCv3Gn
TPKdhBkE/bE5auCUraF58LRwJuoTIfCt+1hfe8XFh7OXoiPE585IH7LOBV504E2d/rvgFXvPKoLs
0MUVrUQkOAcH9SnGLI+C4H1zXO20TwPRVJYfvmK5XaQj5x5MlBjapdaaoS/C3KrtBuIcCXAO1DAX
EFw7OOiAajmKfOX5ES7Baqn3WDdswk2r4mSz9C1uAzcqoYGEr+r0mbpDcem6K9znxokIRI18O/kS
rkkGLK8wQEBakRf/pOCKm1wmOLxSFpqclcc1Ef4muCSv6Hev/vEuUlcY2Usz/FQ3MdOgCt21uBux
nOT/dGz1dH8FSyOTV3kaqGHSV9bh9NYTnnnwWUrZTnOEc9FIY01DnISyYHZjs8/hO2WkthJkOIoG
mxECpNRiMkG7f5ZIp948/6InfHJ5BgLYqKDxxK7nuXLD/s5RSa2BxjbgxHHSkH+BlE3jBOqRbQJj
72v/lH3eshWdl9H21D+OzZ5a9gvlHPfCMFRxtGHs+Mw6djfT7E3AI+SwmMwD6YQLEOGhOBm6o6b8
bEW9XX3IHvfv8GT6vfJj7QCwzIpam89TmYHvS2CIYHHaMZKof3jKB9xhM846oXDbSrP78YWekdiM
OvY0OI32N6zVtzkr4Y0eDxYllGTX+8sLRPkZFgtM+2l9stG2dk9bE+qvmmqEzPnzJgKXRYhkz/i5
Mw+JW2Ik7JhUc8zH28xNdqcFjfglHXUWSeCe4y3jOtPZWqY5HiF6gXhWioc88tp5LQ245edWNP5P
IrGMABIHoDK9KtgvGgKKG9A4A91a2oRuEDqmlRYCYT56TXUCpJlbVtUVYi85QGgN8qiGzqd0xbGw
Wd0GCTZowmUsVrU5PhwMcp8dOoU+MFnkz25nSl+6futS3YL5wuDB3ADuyUm+OIOq+Ca0JazjwbcC
xXBcglPv5AD5erU2X/oHF62rXtI4vxLCEAZp2l5xco6NbuGSbHepqky21w59jbPT1AD8HINVLWNU
G3Si21ofNg+ZJoaVSZreLIHONcaEr+2wV9V0L2722jUEYq1RJ3ILQH23J8iAim5scRQf11Ok7xXd
paKOcqp5EaKAq3SQGjsOi546zJGkmET4mk5/IWO4d0Kxl6Q8ZkWfceBtUf6pvK8iC8GNmWiyCsk0
HoQzfpNUKi4lJuHYCZOnQmWmmrry1HxwmjBxFqMkotDPi0s5xvf8d3UrODWz9IQrfYsWDmrZvTxs
4XiA717YoX0JuKuRm+9buAadEKEgXFIW4bqU8KPZ/idWkkhO0hQuDdxMOtxhE9rhKEJY11T6WDuj
Z39UDn1MK4b1LTEv0oRpz4SPXyV/eAJqpVm77Otx5Vd0RAS1SfvLusV91qRBxqeCm1qydDluopDJ
X/mHVilpuM8PaO8Kd17KzX6NvLcV6amVPazkt9ykO+oZKegtg0oyESM6JU7UCyAQ00Cm1HGIixDI
1oEmcHAXBASb6TPuXbqZL5fmM34c5ESVZ2/awwZVTJmclAQGg1aws11dp4Chksc2ebxm7k7AOOYC
z1YE4LRAPsD/Z2e5oWgNbqFvoFjkWpSqrerGgLBerwn346a3xSbSBfvJblcEMqcO9OnRCRmkyTql
tp2YCaZi1+4+lQNb1DSF/YLO4mCI55DWBKXAsmuMOy7IkhhrNqPVHXDHXxKH9ZhZQi5+htbJH/3P
vepYSUtpJn164v5u9DLItHvNg9bnK/KjCbHCN57x9JgtxscC+hgY4Upu915xF+TSQ1q6Z4jGQzdD
9HTnExJK4ibvN4GQuDnejT5wwuURZnMWK8tgeGFCr2KyaxAgBSsWYjw2r4S9qnbKg/orPI81Azgw
MX9iaQtQLsZEDXD3jMI2RVGThyvCk9hvE9zYQ16OcClv25ThAFORk4EdyX1K4GsT/SKmJV8N9GDY
QCReUCVTtfZ2oFjaWqgIJkX1UTbT0westbnuHFH5zhANZKuvEPEOaefx2pUqHBDXcmHIuu/bGB4f
nhf/IsDG6arYB5g84dunCJN13K3gSddZtAz9o0L6Rb5naSxtkEJPQDw9XhGDULazzT+/xLw81OAw
VZyxBTWd8hIQnMk+KWj2obz0cKmRuD0adeQukRoSnLn4yIE+iRnqoM7uC5VnfB3nelxkbV4mSym9
Ztn/OuQckvBFCqFMDtyl2iwBLRaHO4TTz3EsnOQivs7WzAyWtwnYKibWZwgNfYQU1BujQ47HKv8v
/d9dzibYyEFGwTVHpXvkld+DvM0/ZJZfLtGrSr1hZgOEF3oKkyoUlNNPp3t7SJTvC34im21Crwxe
UeA3DomUPVgyrHQRSF8OSGjuiRmjlKTUv2bVTXaN1jvcwD8IR/bnsRZxX6t65ue9LQENOT/ZtNxh
eezoJwesK60PqFIfnJhoLN7bSV50jvsIPHD2vurYhKnQS9kB3G4Sr5O5R8P+dQkuX5QUoWxN2wX6
7KhAyZFZtJi+Bfly+A/evVUGQqom2vmeXBPHZ0pE+vc0Md8Ya0mP8AaNR828e6pOk6A9s1nahmAP
5OMJe4IEjoAoUPKlOCeeqXCZw5c1/2cX7iz8IHH4/Q+gqgunHnD8DDlQWLkXPUcPq8YhguW+miJE
fAD6Y0hTPvB8GivALjojXSNcf2GWPOjAkeJvXsb7zLgQl/U31gdERRkWSKusakE6qf4W43mYVDAX
oCGoPdTCbQ23/LZ72ZozxmFz+ed2dHOC2DdUePOIG/w6vH6hyZByhdATywmOqcxXnevhnwIMVIUz
ZOi3mWAdKVYwfmpfahXlAAvozmN3NVivI6ZOR0gaj5Z2C0+1x/wiuuqb5GrlyWYy6LEYpd2GZy6e
DAKPUo382If8fBiqCKtnR/93lttgTVLS6AdGmER5CYE447EnPT9882+JUpcyyAurTEiAbhj8HKf9
mFjeYaJ7SzROVBb3tkuEID/I6UDU9eod5Q1FbCamSrjWiOBxSAGpneAldN+mHp+FKjPwy+mTgn7y
Czu2VpF301V1Nu77tTDmd4ovZYRUAA1Z19Ng52Uvg6iH7e0mZnXopSZRfrnlmkxRIEf6YH5C0DV5
X0w7vu377/Gl1KzlWX68J1NnRwgZQAiUUeJa5vmPqLaLAb1009MZNxPYpS9m8/8gQvRE5XBpFd5W
UUA6StjqwwhDi9/QmaiSDAkZz4+T710IL3q2ctcC7jTPp63U+azsrd/E9OAx5FuaiJ86859k+hAK
+BxFf4jmy84UuUz4cIZoqJtGyHlTK9G+n8LuBFPG8S7k1SjbBogCFa8D1EdQoeCseNuXriA8gMxk
qkXQgZ7lBCUL3PYbl3hUoW9ZBd5jeVmme7o2jr5ZgDcyxEQMl/g3OVTHTYhmrrWmLghfjkx23Pcw
mia4+aVaujqmEu25oqaHm6+wHfc7lsnSD44c6BqXshGApQiZYUrb0E1YgUCrZQNHuGA2YlgirV5e
c4IsFQYWFXNtVXD0Q5x1aJPiogpSL4eGfFKzkpaes6UmCvYHO3p8jA5nKtgl60FmbmzreLfRDlru
6FmshfndDKAUGV4P+KkDqcS2bSEPEXKAyHFaQEtmhKaUt3c2PXwTiagm10YfHz9vOrGuMQqRp+4D
Kq5/Q+V2/7ZzX6hjnPTgs3tljUjzRSvuFwHXCxXiksmBBMkCF1OSVOyRWaYpSi97PNmJNC06L+6K
URkxfEv9/ApuFEALGDyYJHq9QP390JAgciX4Vcv3OIhaAge3WYtzxLTl/EEM6xaucAkb6QEXF7Bp
d1WfYexmpigylo4IcGp4FOfZAsUWbrhkcGsIXr53FixbL2yZPXm9ImTznEe1pDSDj72671CP5BXn
WkXVKTOPXX/nWuhe4040Z8diWgzgXu8MqGF+e8nPTBayyaesexuSZoAlhNPHbNAnNCfjmAVQAsnd
VP6xs2p7JT1z+P5+vRRFkIY6JTuRE/xCrBGRwBTsWHH53kpJUwddYOFImqKbep+p7B2qr3ZaSiKX
qRpJbcKiLcQaD1AAojqlwp+XsbwGm/5vJJALPMlFD31q9V/+092q+8zJdVsnNWWYvelGLyfFSdca
V0Lf0+T63/Z/q/wAFvcoGf+2okw49RXl9pCDP1jKoAWM8i2XKUJsWqUC/BREYvmnVoNbly8xQIUB
sJurrrWsL60gWRT2rMD4/7LkQ/4M8bwl8IHXwYftWszz5Y5sO7FajyHdvT3levRlq5mfY5Xxy8mo
3IiwmBT2dqTG8XiWC228hcEHtEvYHrvrVWVkgpvAUhrCw130Zn3nQqB7JdOa72peYlY0WEkJyZYP
NS4hUFAKEbQUb1xwTC+rxNZ/nBUKfL+2rpl4dm4arfN9XgwuYusfBwC5QmVEWDxx1wGUdhsfw9Ji
LZXNEpZEMUIQ7NCoxF2dPSIRjbQxEsZT6ap0IKKQSmTxtQZqobkp7o3xI8eLg5ZG2jKbxW3iuTOP
A0UR57Y3xlXjD83gSJR61Ndo3WNDxpA+uZNqKdm7Fkx8BrHCEHi/oNT46OzLtPMfwIl0QIiGP8NS
p/tbUxqM76TI54PsaPO/NGhuVn8PDlOGk0DwslfsLJrKXuggDeLoFOCJZbVkpyM0YsYqmRHycum1
CpyUg+Szn8AYIVLz2Lhc541hNoISlx/mCLCpWlV0GPOV9dlCOeOwr8mPCtIdE2Slr8wZqo7hVS3c
sBoFMZiviax+z4oHcDU5+M2vs8+2tO/Dl2WIWAikjI+TW2xaBi4RxlWtXFPizoGHO9hlWYuPkFvW
6m0NMXrJpUF0FcY60NXtNToTiFjlp/sfU5dY9OMpOftVeOtAuJcIs4PAm509SAMvzOmSlzhPZkJh
P+QochoRtgcWQMy683/4QjECG1FSBoUwg3z9O88WE4P02mRPXlZ7YM78T+InmFXZV8oyBpUFkSZX
BRF4knjKLr3Zyw350NlI6XxzYS+nBivpmwFH6ZUf2JuZfQZh4wKd0PkSYddwYIoHCru+FUDx/jT6
1efVQ5h8+zimIFBDOCuR8V1S+Ie4V1JFrOpgJ6idBs6amJRSU3S75oRooV6dANoqwZq3leijDEIC
jb7HpHrJn8/DbGAbmWJFPo8s69xxwqwoesGR2RKgnS7k0R/94BP32kgD/UymLAHo8v6Tg8Ci6wef
8zJ00BeQGoDYb7ntOudOJmF4N5ceManfN2jFR4Le5EJ2cMw9Pv29h6VVATJ5Y8akq/I8VcP2uxO/
8EifWGGqWvmv5XptYx0YKAjk9Nvtr+4qUn8vA2stMVSAwiLaFhGJpBih9m2zEg9wrHIdv7mk6OoY
y8Zv/nKzZxGTZSX3+6SgLhxr9+osR6qcREdUzdR6a7vNszubu9CSW9DLzrgBQa3RDCtnMOBlAcRE
ExBqya95Fo1WGtGIgmSaPaxm3eTzwjknuqDEPbPHwCF1RsAo8X/UtNwGKnn50VhUP9fdatm+3Pet
h3gvDPDp1HMDKOub37E/17Ik3VtQ/gTxRasC393cV9PHCeNPydc00Cj1RZfVaJiNNt4U5F76lKuh
nBVPGIvjf7MlkKZ4jBWa3K55IWOR7xADpSn+0+V2APPa8LDBmMGgcWNiMU8BjzV3JLzdPBkkdISS
c5A03VqAqCp4e6lpWrcZC6yzZ72yZh+/k6ziJ3OB15vQaBHg2/UrSM866gQdqjFZAZozB+q4kzQl
/laFVM+FVtnCSInXg8GTcaZmqKk00ZkRvJxtHReWnX2l7N8UqeEzz68vYWLCTkctByUzh6pK9xUm
EflF6aeD3GR+HEbqPWAcBK+R8ej1ycL2uSB9Tgb+tK1t3X6Nlos60ewEQPqRpKsMH7S7u9+k1faA
40BGvzFdLSGd7Ccer1QwLJ7oOR+KISaRx8CLh76hj8lZZv6s/FlBRx1FhukRnOuJYuLiugAKGYob
NkmU8cZ3/oUSVxvHOUiky+w6Rx21S+4lDrRuswHHjyG3Tgkd50aWUNpom/VrZ6TLPSG3JnBeo/aX
Ob/YRXiXPyfq0zpKaUoq/AWYhOF3fXHsHP0+Km/5xu6nwmy90QhQ9KmFLtnhidq8x6w6LCcA00Zf
z8sjLzuDZzbbmTZBLcxYMi3wtzg250FAcqeW3MD1+Yd1S9DTPxegSvJNTKDR9nUWxq7fdM/OiJZ3
Z3D1eoo6oOi/BjF+/WpMGd8Q3/Nj0UMTnCoLnLMAHe1iOB2uN1yfE7gxxnF1kXip//Vo/g+3Bjlw
h1GlyVxEn4RT0BkZyD1AQSVtIcQQ5cpbv8jP7nqCfOUFARuw3W/mrLYJFEE6O+OuRAwWjZI+gxjr
mBctrgRA1yhw5E4uiYZ+aTK1yF2loIjOirBXzV36s+eJrvKlFMmS6QTdl6Z6KPsuT2mXUSulOFh2
BpAXWxXmx5J8SFBLXaDBW40IZe0AGZd8//T9YGNH87NcJqpTayPalfOZ5czlULx0rD0leGu1LXpf
xasTpgJ6GStLjW7u7XXd5XD4mrBlkGEVbzirrJyWFgfFQPUCcYv5wQEIt+7izPOIAT+tzQCvjByN
OjgEjRpNijbTKvW3wpVRKm+HZQSqkMfMhFizm/jG6KSmRcoSkWkIbgvuP+riQ+VajFo8RHknca1O
vmQTj1d6zhjRJn+Q+7hd8XxfYA8SrT2Uc72Lkb6eS85THpicXx/JWBVB6NX1k9de6eGSU5GMldp/
8kdHhHX0OsOhfY0CORYOgNeznN3ujf1/jsifc7+8KD8JdqetGu++IRx1OivGfHXFC947C0clIm9s
9HeXTYizqlMWs4nYddCMNcYiLQWM7bQ0d/tT1lBYAkMqfOcfy8HbxcATzHYgEPtIaAEUNnxixcCQ
pOGl/KlipZWo0MKWHoqFImOwmBqQBVe4JDlQISS2ualW9EsbvNqtRmRCS+TbdLjGSQS6N7fqTx25
i4nnuxtqpp64pigwPmSeZG3OoiJVS7DDGqovMA6ZvzHnbmPU1V31370YqEMzpHdvNN3HGDwkY5es
L1oijU7nAkjPLpN7OZW+u8XHo1/8NT+0cnj1mUypzuLW0bX9TbLxmjPLl5C8mzDHBYgB7tpTcpTG
8xDJWfRayM+pVe7hFD2z9IA4bX653H/BVl89xckuJIq7XjQN4uDdS8ASTT3GeMdySwt7Dw4hWQCk
CDUnZhgcVre0IkMxkp6qKGuuD7BE/a53pyNyHK8+Wp8hGOq+4QSqDwPOMX7VXKHHaIUpT1zMv9Rz
GlGF7mEucrqV30iCrpXE0i/03fmDvJaIdGwE5SgGP3xj8CrpEG8nuysW7Rkp5/Avdn3hEAxgQwa4
9/S5L5nIr7a8IK8lRBUIXNzMgp/xxGnKmeRyqnQF1/pEOoOyAzi1lylXtqcC59hQnIgEHIf43cuw
M/lwpRF1d7iD9dmIZ6eVS8bmRwKmVStDHECkJfCW1ijXMjb+2mtz7s7TiXE9Pd25gxM7ABLvJze5
suzvOFIqMRH7xKGsSaAhoKjKsS1RXVemGnjHc6GcJ8KoRPY988KrF+iHMTcHP6PDbvj5oNmiGVb9
iTZOFlJW1FY8u4I5raZFwhG6CM9ETdHuMhtIYEO8J1QWLFCVUOlnSpng11xCzXsqhQwoXEh5X5Jw
M3nFrAqI11PxY3EykZt08reYqa01XGDmusPIxPczo+s/wxGHltIeqaUwcru/jwJaV6LmaLviSK8J
QXOxVTX9oGyPs29XltC/L65ovfMK0rdAgGMwKmzUz8NkL9a62k67svql1hxA/TLy/PifNTt8Kh+G
auyqIzS4FX5VmCB8P0jGxgoRxL5800dkVkT+HTWiQBkesEol1rc6ep/mMSAvNLwGm1jZ7XlViHdo
GtkD58qZGhLy/eo0CB85l7WqAYBZXXwa5ugTmOCxdGcdmEjBvJuP42qhV2M2bCZ6Zx9Wc7Y9+2x/
glRUhV3MKW4vkhsMMuHmKWJm1FMcdRGehAHuvE/G2Brdy6oWX87a/9N1gxAAX/0iEKtChEImwy4I
oiJ13QTnnatqYNqQ3V1OzYYpbKCdvIACvkffyjPtKfpOJs6giM/fVmri/gY2MSsb9deiplXV5uvH
na3o9EGTDPkXSteDwIv3xparPW7O66PQmfXn/RUxUj1Sxo4JikUGW1Ax1PoA7THWlKT9PWpYj3tB
RFK0bVkgFh9yydk2o9RKqG558Aw50ZgpYHkWhXgyP4Eb6QRB0qrxoLjIAZx8+GexwVD1gPt9p8/G
vL4ZAFe7mt/LlbBFRwSi4DX9Dr6xlon0bVBqjYjm4DS/pui/VJlNP9/5I7cogl1NTDUk0OZPqWAS
bdK4TdmDxds02fiHGphXVAvq9637pdM+eO2EjUEZuCIBpeSi95wIpQt8O57Q5A9WXWGOBbHL37Iq
e+sVNNU+vDIHpB6dWRcY0X4qwXAEdP0XIwQchnWqaGAlkddqFAVBOd5L+c0hykEnfSwimb3aX1d6
AjxIvAGXS4C2pgiIoZPn2wiwRdLhcQHYI0A8ZyYQBSJXj4r60gr1ooNjaC2AmrAoXy+FNfe9L8rP
eyJX/l5CCSiZeiv4krgl11TAZU6TwIQOvkCNZam48ohptsclCAAok9iPGPQsFOVK5SY9sdDqOu46
5YVcwnz/VvxDlKHExWsqVNe5CW4Y0ev+T3olg6kIJHIiYBt/4jVyeqDucDl3Y+SKqPuMIDc1Iznm
07V472sKQVXKxXHEXtZC8z4WXXUVzmXJDkgKfjXiuLfW4ajGl1nMv9tnhw79p5RL/TGq0wruqKR3
vUwgHk8OISIc6Poouj5QrNPMwNR7Q1xVoJNhUKegMNRWKhzgf/yEoWYD7DYeZZssDmGSH4wAcuAR
sm2zm/rm02lJrAtIad2Elff7LJMlPZGt2IuIrLnfsj1yyHBzFIA2/dCSbh7IsEvPbU8O8UbXLREU
cuZ2fGMZA1x6hoIXVgplqAyQBMsiMWHe64b9I+EBgmoShDwW82Qx2+f9TEjd8TqEkV+nPht/XGI2
oM8FkV5+UnJwEj8IXmQr09O4gng5n5zifUcgdcqqQ+oZgXzrb8lNvZAZaahkiKjxwa5S0Cai7cX3
TXCBEH2302XTf7+KPdUnHeOvACn7iL05ZAF4RX/MUxmdaK85rzrcgey7ZNQZ1oJTdRW5dsn4jidc
d+VK97geeYZY8cQuq9xiJfqb4uWa5IdE0WRRF3CpjnxZCr7CaI2XqBHKeUhhHcfZyHJVcV91IT/v
cqyKJNapONNIGuAzqtRyPAk4qltPSM6YibYwG8r5WtBAcxn1IGyKhV73GbaMswR3XiVuQ867zTt5
C+HIR2RVdWcDc2K/eaKQ3u1zI5/LS2go5x6gNGD5144ZqMjPKkBeerHLIqZ8KKyl7+i3GdYnnvRo
7TslvUmrtqhmwjAB15ETM3Tf0kk0InFhiS0eww4QwThWuYnCDdF39Uh2DlrRHKVRwLdwFeC21gE4
GWafssW8eGpElgcJAwNIHXRtaHvS/BwclgJTR2wXmWXVjfwP7AGEHDO5GdoWnVarRd/tnUZJachL
NTpOdvrP9dxTbt+DrzjzRx7k2z96bLZ40nZdMLIuBGTxamVEXxK/pQ+uNvyCZXOvjI/v+wQ9W4eS
rUnRA3tlhnBKGx6iE9x3XZEivV3Doao4ZPfs90N/maRFRrPMcKdXLw2RXPFHtC6tOMD75Z7XcROh
emQIwASDTPk/5MX8760gp4NTNIal+U6sWIN5mG+Tc7vxlr9QFPpcqdCgS0xxC4KzI6c/oBu7DYSt
h2PrAbDPGGaZZGecDfZXLhqWDkVLy5/XaVmPJvgVpUFJWPvoMcmzwrx00uiyAgjOH+wdkGSd7nmB
e5jCs5TX7bhSwmrJtYwqcQDqPZIK0EivLEP/7MZM4dq9eVu+h3t3YQpqYHo5QHfI3zq/b7ngEI/g
6BU1Wrfn8T/EFNAEuSQr4hzAN58X3UKcvuH35dfOd/sj0Wzhl4u6FMmvN7KzTDp/WY/G3XLJ99MK
LIOjkuVMaC3Me2Jda0wKjWc051DZhQGKrUST2aXoyo/jnlmJov9vkCPy7zQZ9gvhzGj3pCSSo8+L
tDj2Q2T3tPPIF+Zm1IybPa1ZLuRPiwhtSvRNo1LD65D9v2ExYPRxadDWP49iivjJEBlBeRtlOWb8
nb80bc1AYFc6d/ggE6k9QN3aYLH/shRgXzf9hnkmR+J9Rg53AkDwE0jVpTy1MAo5kR3fqCtrgWCX
B9EXEt9D/U17yxCg9XZDfytPdNk97zfXMqFBLNREpMI9COqo7PIQgBrxAAkhgGJG/GsG660DyrRZ
tIRf5lJOtSeYpYhyLYfaOmvF1KHLuDyzc6/bIwJ5Y1KBD2q53fbIXrJFxaeyer3leGtqetdKxZcT
9x7hoHkCze+EoJ+NvKvbyiGZ4HjzUIJq7YhyHvbj4Z+v6bJ6r3iu813L7cEuwlbGF/rik0E+eeSQ
6l+zkEbEDfAE5QOwM0BectLJRPgly9j4t27fsnb7GMjxYOHZ8MPGA28mYUKkPY/0b/mRRG+WoF3w
my8XBt20NWw3a1J/mzOnBAfl6MPsaJsb1v3YBxYUJ4WtmkqNp7JKus5W01TLQoUzLvJa4W51Jzee
VQXlgrYxZIBNW3gcEhm4XKO/EAZbSM5oLoKhMRDxSCxjUoWfHz0uPupYHiVwZfSugh+1jalKDKS9
0/n/Y1//99G8wgzCnHEcVo2Gg06UrYRkzypj+CUXTm6q3HbcXQUB451Y/KKc7AliHcYnaBEei6W0
+LQIN1cmjL6cPb3GJcknTTXkDzRsqw/YyIGJA0xiUF5H/HuZlkIP8IpNyDm0swcFYlaetJw7NQ9L
4G9wyOEGB+17OFry1Kck/PZP9OjTGL3ZWFSMbh39thPM8nQhwQHZtzdKcz0iqeFLNTl0Ll/xQf7N
uNnz7Ki/FMVuKtC1eUlCLKmxLIYLbBFKiJdUnStkxKsittoeqlf+5HQWbBR15K/Wghcx+gnxMX+A
REr54hRjVehgBxAY0rcM2LCICnEG676C1nLCAnky+IW4pi+HNrhUuimmMxAZsur3ylQer5hO5ycf
LCtNshsv7pNHF+ObF2IwCIVo+Ab9UU4oV7uluS4mWdknD2cWmS0EraViWp3g6UQ/ws97JnFQeU9h
OUktCkxkab28icsL969HMIKplo1Qi9X1JKGtYmFpLrxugJPhayGk/W5J054nNiiDdEk9yC45ta+8
2cQvmLj/d6x4E4PJ4YElqT8A/8Ozpm/oWWzz+cH4f4GiFiAFsRqTHsLnlKv5Z9X8ZjldEjRJZurK
6r4c29CBU8vkUh3a/ku5iSrwDMjmlaqe80AZw0xjMiM3XSU5BmERDZZQce79AolSTc7poTbeScic
wpNfvZz+xI/64yCgzezvvaSm4UsUpgwsTiyaIPDR7055SyF3XbxVdstWqIjUY7I+7lnukGF/DqoD
4/YVCzj5zYQEU1B1X9AbzjIYp4kK8xb79USzpgQeoJbu8Jl9Y1T1+/z1PqZzVq6kSDfJvbX//9GZ
XfAfv0ZXyk5YHQ/+s8L40g2aPNJkFry7okWXfbzY+isKjlbznfZySFA5xQVq64wKOPfucL2oId3J
JBM5bq3KFkYo+CV8Mz929Rhen9hpPJ+3VbWQYMG2t+uCGer3mxiCNCPNoVZUCIyXysf8Qa5+MUQS
+/IlGit+uuLLccnrf1BxS2pLAJj2vAlfNUL2dbd5kfWbdScXPNp1FjjF0PqRdjPzzjwbYHcEgyBX
fZI5mqaI7omV0NG6QOGuWa6VNdYpH2/cKewtHR0GyvbbrL15iDUd9ogFEoy30IP3k47Kmoyd220v
y/ztG/deTIpF8ioHeDPOMGlZdNtAuaWSwYw2VaWsIRCrikgUZo3ZWbsAOshQcqS/aINY4ztvaN6D
kURAiM4+vwFZd1WElEZgGQjH/GYoFL2BlNZH3HeGiX94MlaEK5HDu/EQyYiJLxfReKghuOSBLOlS
7fYDBn+0Pdq1XUSZxk6y/WcdGdB9i9xzOQ3Va49dmnAxazpjqyBnXxGJvTCcxaDCxtrtEGZRNEL9
0eMmLAQd3b8dLnKmIzTI4V5hUb2KRvoW0+FPjvwAycStTJv30oC0fWTKwlKAMuNHQHIIOk1DjKQv
UgBB4HD6OTMY8zMT+/RPbVr1f5/Yk683TF5opbDNfUAXzymsTpx/VgCgPn//iaRSKlpJQ5/uO58Z
ASUjgg1Gel1ogamJKgFooV6xj0+eViBeHLAuAleZWy6arFQ4zXta6lU3JYiiirBr3W2Q1/ZB/a+k
pYcFaZAAz1zVfu5/c260zLTVNWsfOzQ0p2OEriauFY/L6HnONWnFkCH0kzCzdemlwyAPNLqYumR/
ArfvuBj2aCIEH74BU3bWVVBz5+y5QqZyhHkt0Rs6lQ2/PT0vlFN87og0imtruhCxojnvPVuJXdqP
9bTjf4eDT010xtrnDe/PrDJmZ8KbWcJV8+Idk+e4iSrW7hv+C2BMJnoYi4PsnlW12EOG41UWlSde
uUw52RKOaBz0bpretCClVt6oY96VMJ3PAfMw45vLRvLkp6m4PkG33y3buKU5rQhmukhkJp408sFU
VLLW0plwE/lMjiPKm+fqQ3JoKgPTJz8v9VOuP3sRsVyG5wIT3ahSjSjTKiacjwUJX05OTdnfXGqC
A4jWD8hyD0JZKAR/gz3+6/7hmgqVnjaGW55OB2kA0/FHLcgqgPbYMnERnuUXDMFqd6qRZN3O0niN
TG8f0uPWCelWZa8WUXeLa+Pio7qP7iUGFE3i67Gx5q0f3YdzqhZwDrR1OeaL5arOI1wvbXti0s4v
+2x5gmPjyTselR7+AiwJ4Lo3ERxbSL+jfdUScJhv76+gDT/DfJO30QwlPDlouSzDLa9powUg3W/Y
y6wNsgr2q+GRdqCE2irHEYKln6eCh1FLahKO2jmpl8g4MuAEEE0+DbLHW4598KZ3aMhQIoeRef7w
z/vzSNeahZK0TGB6hmoQrVrcf2CaDYUzAG/mtCMAuz42WchX7R1J6ybDvhpim2a6BCLev6AhzdQE
Hr8dOvFqPLt9qW8AOXq6i/TkSnlUUHSzAVLC3DZKMZmWCC4N5Fy611kOHLTK1lx3fNpaswXATGxG
TxmGu4Vq/RqDAY0kVPP4wAtIR4QcMuStkUawKPgRWZhMDiYtMuwSDktpU+eKkEl04bBYsG+WT2tW
2CqvjjFzQVdYIlMYXzaQ2V1TUUGoQKVoj17iEp9A93XmQOMRUnE/KUXS3OYvRFFsvKeEO4XU9eHn
ceeX3nv0Hq3c1KDFa+/XrbGE9zxRvh5pRXXrabUsJb1WsPARp2LZJkrV//87cQxN4YjCvWU/xvJg
MRNNvm/pQ7H8vUptq4vc5xuA7AAthDWT66+iIvghi8bfD258wYnT03ZZPtQbDya20eYYQTuKIg8/
tl6Et92Q6rC1qbnftK9eBGzCo9jw/d7jMWOaG32ZozpYN98JlQciN9h6zdAFd0XD3+jvtqC9BSBX
i+4PreIGCJrv4pLMq/wheNCs+54fziOzRMCJpDYzJSXOsO+LoNAUAAmuTj0mrMikGYzNOYX2Ecwu
7tWHWzWthykDGWzNn0vzkF/XkjBRyxGfxPxWB0cRAqTmUSkKaRKgdN5GV1YqcrZ0eP0z9UZ/DbUc
q6qGz98xtt5n4Z6p79CMR+HcASV+57Dfv7AfEsvMrFUJsOI07JC+vCxKSLSlM8/o4YKImqBIshH1
1B6BZB/Kz5eMFLL0b8T9jCzfD5nzBowS6o5AkdGLPqCihfMTbWBfWwwhdCmXnqr8fedG01GIZ5R6
P+u+mPVUlFQ3PBPEbh4sxe0W7lq9Wyznj/4D9SyyY9foY2R+ONODyQd8KeELUfrUs6jFgfde3fT2
ENNPa0ER9MWcuOBK/03fDV64QOuO2O+5ygrBLqmvRcgaV45jE87Tq/sPVna4bn4WpKbK5h+kc8O6
y2GNwwQDm2eq6+Bs+4iot9huY4zN4wAUBUt4HfNFTWcyIXBclhNDYZgQOcxcqb9mQzDNjyqiD/NO
uYK4yCFoIGXl65LHjdKDAy7QojNh6fCRYuZI1CQ8rVe+bSx4PpKqcPMZSsbbja724VdiWSlNGQHQ
vDpdXvSzIv7RVYvzsjGEwGHR4F3na2VXNaA4DrHgDViY242+cr+r/V8sc316dcqj9Bzfuo+TIWQf
bvzvYbRPSoQQRlqOl334GNBPQYinPPM4el/B6BUouv9cXoP8V0ekQ89m3Wpnb9Ed0ypfQblF2Mzw
tmho/VM738drf1AuqQ/5iNSA1qa/G3tydV5TQhyjV0d6NOImsIij95zyL90zy0RUKEHbNIt3iCAk
LD7eSHA9iYoh4oohfgsZkenWcwTtZ6HNSqLUHMMH/G0x8a0YL85RU4WsRYqvrC5ReBI9V2XEMMAm
/fzogpsSsVWu+XoaiXJfZWOOuS7zOO9fW5h98/UXwsGVdPjoR5bMByrxJcQnSlHhHx7UZ5sZ2SFT
P6TdE2uc+gxD7VcfDj0BGyfUKS6vMaf4uQAqM5S3Bq9R5UWwbGbpSNqNZOJzloFufnGQcVSicom8
X5qB+gooLhE0JYQp7FtOPyz+gMHInz5xA1XCcMtaOUPkxJPbUVNkc+cRqORC+wDESySQV4Wt1a2V
zPO+0o62BiqiHKZnf24RnU/1mVJuTtH66NfVo0uOSz9IImrpO6fxBSulckZloIVdUdLL7nygndG0
5/Xg/uGWoyqSwP+VMEducjVoQgcoDEvMxbsehdBpSt0rrB7gsAIoj2k81UfaLPlGhAa9A5uPmZk0
sYpouHppq46NeRGxEZpPe8iGO6BlJKUyK+H5lLuuAKTKeb2UZGVSJQhQQ48ibLZN0+t+h5206Du1
MGWsYjKKM+28YZmaECh0pTJaAjzJ2dcGlvivu4YXQ469nnJJ1AtO0uRE6/E/EAUu7Xzs2Xb8xPAQ
028uYTlLPQ1iUrU5K6r+Z0+DsqtkDbevgY0Cx45TbGyY2xAAu2ICjC0FmDxhGSBKwVEVxh3OEhdH
38o+ZLaACxBRgpqd5xWzK2S7ppPrFTVZd7mD+s3xPUNs+z7c9U4MhrMBjcrVhWK5uZPdDM20ksvC
CqllSwDelgG7yiTTyF+L+PHrSUTUQ7O6zJhkmpj5ZTsvUwDTPF10WVGME/Cz51lABVjr991e1KnJ
CdSY15ew0GpewX27fnwpWxSNt4Yq5FovbDz7Xkm9Sphw+2t/YUUCvmMEgLHIDZDObemIElucgBIc
6HiO0h64iHeMxeDWvipumxtPGYhlyyMV/Y0wu8Mcm7DK9Ef5MiOziuhLy+aeuU+GVlZC+2Etjqrz
lt/6Kur40L35/FzucOvqTvoIMqGSWSKrGDu1T3s9nhevfNcRkNwIt7cIydMJ5v8pW+0Nb6OX8Ezr
3xdEDw1dvyyFzM6aK7fx0QP7CiN1ocCCQqIJGoeL8yQ1JMX7klTbkLZXUH88Zv63+And4dqywh0k
kZPVU/5ITAhP8zO4ur4GawQsMF1xbQKV79kNSziRH0tpuFqaPT9pqkUGq+d7Wu0eyMRWQTzdp3yw
w2twZ8HrHicA3uLyot61C6vFdhXSwZS0MIVYDCZ5LRZ1ZxI7Umt4go2Bp1EnwtlZT6BNr2Myyid3
WK3tf5IvnBE4vpa/N5RawJFnrsSwdRUdI0gEsYM+RKNEuKQZ/AZqwXSARhFn3VQGi2WKtKmUEVsq
NPmPizR2MWOG/Du7SvofyiJ7WfJMSXiNDffxVYE4kncz/motODjKYGlKLrJIVblvKnPIy77VfoWG
hvgOwXNSAJ4oftRc0TGk/LnbWl+dGS+DJ9Gq2ItfKUuXO9B5Pe5KtRW2H8D4Vr8uWHYJno1w/5FA
mqvtKzVKzkLtDCiR1TxKrAfoefJn99zsWcOIFQP28mcOQfHs1vsmI+/nzU4KSas0WHC38LxNaPOr
TRgonbzTx7ObuWsyb6rAsOYuX8J48Qvr7zdutVvcK2bZT7DvB0S6wOgY2LO7Vb9HDm1NEXXiOXMk
amyJaWGOnnB2I3iHO8eHN4r81vDPUNrGLJzqZpuHo8UtrY12nDhD5WLR6G8wVi4xgUjneFMLqbKP
/jFBozfTw2SCDlZY10LFEP5RkzHgkGqyzoPi24XulqR4u3kaalFsis9U2Ip1McvkA/nnhgH4jOoL
ON0N9Nn0dn00vxXavkb/+lo2qGoo/uOh/OnozyEywwmDFbBeJ4vU/fmm9jUT21JxNbO0p7hXSUE2
ZYNsoYO9suI0hdiVRaa8uiwm81ZrY5opMm3B9p3Sy3Fce3IpEIZsxNzUWRyjSelIkw69KjqnadOe
qlo6G/N+Pb901x9lwYWC2chjwXkR6KVz8TKJPNpsLXidJfvf+AbeV+A4kxeDR+68ccgxej0FgIVC
K6y071dFy15jaOlZvhxJmUbKsXgFx+CPipkcUVWi46iOkiy28MOJj6II3HfNoBJF3uzGryzodYML
mcuTSytvajxlEhU/VHlRgadmfu96mKOJ7O5fyS2h7ry8gupM6Op0wZOVWOK/uphlsOOPxsSvcagv
6pus47eCBvnzE9WPr7kiE06Fxtq5g+fn8dSc/1ZX10l6Nfln470zJwMGOKDsmzQyYih92zObqZzv
ytAuCN9ykm7P4A5XrXj89KoocuUNEECtuTUjtRIPQOJlS5y4I3IEx9rcDFtOyuSHKFeHwiJIg/5n
aA6EJNHunw7qgTGrltrYphP1GYeJ/HIF3iNhTSXcurSbI+8Z4r4rWerExco0lWxhafJAt9fXXgdB
XUVucuwx9C5vMs5I8ZfxPCYzp5qhMSHyfTpR2KN+dPoYbqmpX673cwq8Y81kllq3DS0PnjW9HQAi
tZIMeGVOj1PrT7koA6W1Jn3KrKNHOfMgOnQK5LSPATojDc/JowSbRVpvY29Dv32atOpPg3i0N6ce
YLUTaOSppZsTui/igNHYzQmglHkvh9BZvZU7fw39TPB5ZVTxl/DmCFODelvGY5qXrncIhPIxdXqF
/OHdSbf/E+VxLJSds346aHjXr0n45hM944JDWS96ETk7s4rS0L88xH55qlK6IPq5IgHort+qYaAo
O5mHewyYE/MUuIKrYEwlYd3lVPjBBKrSXtNdNKAi7JGQ9lkTVke66rftv8K1+ayedchoTeL8kDyW
IeBh0rWAa2pvbLLKH0YaKyXDRxWIExEW90RTyI+smpKK0ZgWXtOszTjqkeFCC4OXPimB/H7yN1RC
8dPjMx2YAfUMxByGe0AgB6d9BvtujBRh9X9D+4sxOvK8byLAOgaSTcAOw/bdetgY1+8e9XCNUkk7
PWS4tSRQ1J6w1AT9XuHsLJq+iwMzrjuAcnP/tH+VAIg0wdnORT8NiLvOW/IA1cJpbvJiVp8JhKPE
vQkMsjzu0T5JbMFoW4GfOc/zAS3M0abacw0zsqSac5SlsPjTp/kN+NtYbzw6WQes8T3KRPwTEFMr
N6/oTNQVmMfINkA7ufWzbwC/OX28MzcdKXtZev+B/pyoN4TcrCMW1HNESi/aZrLHvSxVZwQs5MgW
Jy9LNep0Ux2ngjNSBk9svlzRhzKAAB+v74NbpMtQuyTikJDq2OKBAD09GFT/HkACP33J4pmxBQXR
1FJkbH8S5y7RHZGB/wMkb9+55GILRu51Q2t7sFpn1CK/lkVdg8uRjmgoThpbmdPKMZzf7ZJc+TA8
16Z4XQf7kG30XCm7KgJeqIlL5rG3SpRn1sOY10Lnra9fHHjLAbqX2yuBO0wMY2ROZwJYyrGZ53Mn
dqn3gx9Ewc5IId/hAexfeycH7AaKjqAbA0i/v9ohQiia+L7ayETXXSe3o9WtGe6hgAJzOwVtghZE
Oa2ydMVdaYTlnZzwMOenfeeh2Tt9f0yYyHNPuIC0lZVDpmavR3u3s6QEGIWULkunDMr27gvwXBcR
wnAGtd0o44lvd9/+QSTpDPkOr3jk3cjjCFj591Gwp3J5obnCnXep2UOGrFqVuPMK1gfjJeYI8Q6w
rFofdLMWh4+6ljySSBvU2zw8JXhcNYy5suu+uZ34Qm6xT/809kuo/pvpQcRat3wOrcJ789E7sXUo
3vOxAT+3svpJaTVw2XosB1HKQFKUoDagfBziXK19YRelATWnNPxK3Jmix2IfNduCTI3+CbfNor6K
d3J+NF2Dpmo4zV9DAsns9aC5Nf0vjaYJP+QjkBbpJsDIrb1NZFQbNh+GniAZJ8ntC06Xhq66IR5P
NXlJAXVhkgoZ8Vj/XWNABF060GG+y8pzxUGa4Ymkb4I5QXjB4wzXOeHVzwebVRK8cGTcOyLYGNrb
k1keXohPEJNTh8FEM3NP/2sHl4osQzB46oO1YHWZplJNH0fAwZdpEe3hUbVwpE1a3we7JMhI4K8u
Xe5qRrNMMmJHCXfXHdqKIT3CLBAyB+XbNncGzLk2dRNCE/AGgMKEgcRf3XRl5EgID4Z/7ND/gh3I
I1JpQt/42mSyn9BpK03F9yu+BWw2TsrL9jXVWZw/3d1xeWG8TpEjSz0uPuXBIZTyvkn/o/5nxFOg
sNktjU2TLMNB1zPxTAqJMre5RxD/Gu0i3esOSKWp6DNYCEzX6R3AFDPAr9hgw5kxUPHT5FNMDTAO
OHFfutqA9yXyq6xjVWiVyAZTXRAZo9YyHb+7iqAxsXXdoHFQuwcxVaWzt1c8yl//2SJF1b7wVe9a
tCrkznvMdn1eKp0qPxcykBbt5p5MS8OIrclv8RrE6K6aJX114HFBbv12UyF25qay1HnbeZ8byBpk
LUL+m339xlOIaSAt8CQCkHHnqom/bdwYBzJ3r4RNlBuRWgVSO7Ut4fy5Ggp0Sfpb+nUj5Yma9UV6
OoEww+Eg4pVfXkS0E/L8U7NIgYvsaNsej5rCPwSePDCLRv8i7Mbtmlgu9lo4p4L4pc8Ndl0zVyf2
gwQ6UTUtUqgwvFt5D5jqALhw80+Tjew0LCUFwt/OUXafisEHXOCFvNl7s/DWniwXvQkERMc7iTPj
X3Cf1H+t5yCbp0yRTQp0KzGHQphCOItAVHEyGvsDAaGbS7402t355AKgoo+LgMtkrD1Wg5VcaTtd
N1vs6HOWMf5cfx4aVys3Sg5RGoy485es0sOLvAcdcHOWGFgHXxvPATNGH/yJpoCEc4D00FuhxiaX
3JvOplHEg/auCzLZUUY+gWrnslNoOtqsN6YwHe+5zRTMjxe1Hcty0PcsEqAVf7Dc3buGOf1GNgwd
fL2HHAY4hQHoxNN5oeWp4+HwQWgQhFBBrRl7PxlF27NvVbepNIwKov5SfSjh1k2a2eVSH2sj3gIN
6l8MM3U0BNiQllXFy5C4EZmCSJ9/vvURxc6Ba1fTY4Uhok9aMHbDApYyIyTNdbJteshnqUqNjpgb
CartKoXoRhKBTakkxMA1uvaLUL3xBG3ZP5wHpC81zYKcQZyzagiyJjpMNZ0Lbz0/Kp2IZZHX9aAJ
lA/gTCNL1zPB+xwj7kvsNXuIP1NYPnxOaOOHkRo8onFtEEdtRQJsvrNbuMO4UrdU3+FgL1hVwIf+
k5oxvwAh6a9v92NIRhlT/CWneREowk7UXM58lWjLEOe6rLd9/6H4Vt6KecYt3lpNW60j77IMfqcZ
1EUuZseP6C82rjr2TLR0EMjf0PH2DKBGINNwXK1GAXeaKXNp+8BHjRpxwKllS+OUi9LfhZo0WWvd
E29t5JyKVypcqB58//hb63AAI4ecoijVjjKg56guSQr1z1qGDLtnHdKW6C3L7/zWUScDTl5fbLGj
PDI6UAT6dRi2pho5R4y9pjtXEJcHKJr9do0ZM5f6X3icCZHcX2jcMunplbBgk8xifEIwI1qNz78l
EmYs873dEfMF8AeCIXqnR49HsN68UIasdBO1OivEDkiuNgo06oRUd/Mju142uWJlnxIDBKA1y0aO
qbxF8ODxMZPyVIqBhwgjCtMyZZx8F7JD/rH5965AIfwcyD7zLE/O0mBGxvkcm0SihvBqFtweRAlg
gVLa2iZNJUMoSpboEB3LvBEvA4Ix7lY8n4xZQKrM8dytoex7NiJysz5aNOT7JdIH9lwWFx2e/x+H
EZn8nGh4z1SGBRUQrATI9++g2h/dY8jE4YiP732oq1THus3xeiXq9Th4b03Frjid3dAgz0nhbKEk
at+7iF8ULKc4EYpBTBZlsIvbdJ2kI7vQmEZahfidzkBRCdFLow3b4/WpQ14VMuQoDiSWaQHGK6rK
804Xy6azotNQ8jl1bsBn9wSEmOOGZgGQtdwWYYAw4kIV7dq00CHvdKaSWOzG3Av8xav6m/TyCB+r
AeFJruFX02rZyxVeGVd+ZkoQobXzD0U3gA/Ho6PPRYZ5xj917OJowscTsW6niYHooKO83RdgmwFl
3iThEEHPr/WrwPtnjwceyc8cyxldtF8b0Feq4LjXbXo4ZlPSZLDv6f4XwZAFD2tdUbqGLI1b/Odb
MgoZdsGmENOsKQGLW+xCJYJwnjcoy15n+yDVk22zY+Sl3J3Jnh/jGzDLmTTKUCFM2p7Eh8WhLrgS
oiPzdLrQ05XAzOLtW+EUMlpMZN0gQSFC0besfJCfsxqHhTyinRvMUmKaW/GLPUxyNrnoe4o1D7Hp
xdnmqcjW5eW/7hC3+E27LMr1GckEnobYXVrL+xp8Xol+vA16bD5WW0EY7BBFQ5R+9O2LJtAxwpeY
TuIzaIIadD8bQghHZKnqyMsr+HPkn4vXqMpHG/mh9/YNU4MEDFXQ/IOyJbF53QRseus2YEE3tapX
WZ2ElHe0eYRJs/VePhsAeI7XVUARkLOCJHy587gHDHBRf2VYrPZJwYmbRmHBzLup96qraKEYVnUJ
DnA4+aguL/XYJGotMsiUUVIDNbi0Gr6SkI6V4T5HzEPMog7p6tdL6NUacApoREO5VvZQ/L8rFlej
LVmygaxd2PeNHXqp8imNHecHel/9nbYLE3xt9SnZ4Hppc1vOTKOTBRf10KEYpMky6TUjwBkAVWyu
ExbPqgsNKzv0GYLXe1/60MkKfF5+jNlm8zn6e37cAWobf8piYQzJZl7mJbws8nu/BZvnFvo9lL6v
ZlZJHcSxzkOi2CZq10Xv05g5+kJfBBhgbbjobWjbOINTV5OaUdDKAl9WI9K5aL0A/IkLk0RYmHBf
MQjtPxcnxk+LOScVYZhy5mhCfDJId+zoaK72SaFO6k1MHPBFNH5rmu7OZAQhq31Kzhd5nmIUeewF
7JHt7o8kXrnI7h7QqxVwuGTkxEYZLwT9r8VtEBEbBCXC9ZGZ6VNwnDynvHiJ3ubWmdqjm3qipfPr
M0W40oFPm8RqzetG15Q+DodK+1g4y7zQnbQkqZt0ogOA9+SzjJpMQWNT+a+VfYLwcBrzJl/z13y/
N/LGt1PWvopuwwr5YYx7NnDuZb68lJhW1mjwjbY1+RD/hZsio0DAwEnJUlpxLKGsbreLaylDQwtS
QQzzLC2e/aYEnGxIKgEc/caWbO8DuhDmLJsPCzNEp1Po2w366Mc0Vqdl8C2qp26zTpIJyfo76NER
PCcunhQnAasjq6WBHtzHNm21QbWFNL8kDdd/efQPm7iVpl2MR/63OrjVR6g9wr0h86sjH/nNDAUb
TYr3jBofo8lcwxSgT0RQ141QAYzvIBKCj/jX69j6qb1LdkMUwKR93LgjPrNrswbooJFgsZv4oe98
eylZ/juFVTunmiZ+vygaM8fS6Z+2VBwDIcscB79hJsG36UrLwpJ0ezND+EZybODvsLM9vmC7e5io
a55tghkvFcS3WwrTODmHV82OxBUbYRVQNqjvxhzLAlDAsQ11Ecite6JEjG3a4tq5FZirzUx44/vc
FrUuGrvJntaWQA2JPtopENepCxD07s4mDCOSuWGTSjHupLHjHpRx25/4m+nS2fMJ7FswmhfD7VGx
iNjifbKNqKybLQKNoPfLpfZ/XP59WRqSgqEVTUpkaLWsblwy4EuQJ5EXtpDW+bsut4+P70MHpztV
uQz2SSWnvCvsWMh4L02mvGQTcx+g6ZtQLnKePu/InRB8iAIotJC+qEajFTrZu9hyXzPEcDy2nWI8
Y9EraLRGcdXExVG4g/Bttu4Qy0YByDhVjJBYa/q5pivMN+RNbD+/I4KLqyXNahDLdHlKOeoPVcqo
1KNVWSJaz7SW6M0CLV/zSWCmHpWdwGFRvxEbjQcYbP6syOv8TL7uUozLRUkxD61AlOPINXkqjk17
qYofD6PY1K/Whqa5IjFJtU5QXanxh4pMZVJoKMyn9JbK6OfjIhMvdGf1LpJZd0zTp6kxEtoZAu6S
g2yvoaSE5RDAT8kZHj1j6pTsCfwhrUKZ5xfI21na7lCW/LgzMhSR0JRqTRjZiEIya1VlI0GYtGAm
gvTzPqi1VN0Vmy0t3lFf5VoeG8lZtV2fc7RQsdR2eUjOwzcqmJQXZyjw7W6pkilfsvVy4g7wYrYZ
NrRlFxMtH6Z8x6I7PVHUUxiN8nllyalAqKsJ4TGeGPwA4KAZvL6ej5Lbk+Oxd7qC/wZCGEA/WkiQ
mVNZDMim1H6wo4TKRvGjw0a+HTS0TYemGd0u/PcN+MZeuhrR6n8TTDFBVBrHaCY/eieLaStKs0Tn
FKSuTouJwknL+gngBC5VmPUcrvyJTjwIG0/s1Rfq1pU1IFq5oGKoT1bk6WQfDII9oqYiTKkzz7hR
MF1lVOCQpPpoUCD9jgu3mj8lUjqDRKiHhRelEgyr+6ZPiPT2u3h1qqvea3BrWVt+Vd805ridzFhU
xwiUph5MqFRTJcuDfRVsEcHMOQuLwFARYCsGaOQUrxJGDp+03Q47pStmoMN8VeX7Lv1tolUJe4a4
isEbN86Q8IX3ERF2sw2AvwJ8qq2vNNv0AZPZN165snu2MTBMBv9ymb3GVmdwWO3rSx09UzeFgfLt
dGhW89ubvdiYiOKOwkEm/wuisK8vKOZ+MdnJJ9xJz/BZCO5G5IjYmS4vEbyDmxYCWojUIXVFh2oZ
lW+SRBFNWzqWRkQ+sGxsv8meMUhqbt0e+XDqWkKJByvK91RNiSa4EHpkAp6l0pjCzAkAhfKMkRof
+0OkxUzJpQlXpu0rF6DX5FaXutYFYfnZbCnQs3RewtWz29oa10wTgVEpo3gEXA2aLRNrs0DKRdeu
fQlAfCZmqzC5O/oN7qz5Il0qH7Y83AULRX8ezMhkLdomjQGJj0P9cl0L7cSkSkfysnVeH6dvKfpH
NNW0PW8p/eRErmArxWNZkIbaQxpL6acVGWzMsqD5/XuwENu8DRfJlqbSz8Tb3dlRS2RqWxOYGdzD
kvlueQiKeYGqcPfkVEOtDMEvjtHhXfFFkjHvUt/6x7jdft9KbrXDbHZp9QatHO0+e2IVdj8AbMZs
62cB3a58cDq7to9m6S9PqRQIFP3pN58uDay+Ezj9ms9MphICQE7eX14LIQNd3g7vtXEeSP2WaNPk
Wqgs69pEJOVWL23QTfnkQr99SL2HpybEtqTn2ZrbQYlfHKF0vEqelf5dW4iZpzvU3ryn8uD+QEIw
2+T9hbbmsSAw+cSQbPdX+zAbdQ+u/6wz0YId8H9AeCSqUrx+TJXOq8Pmg4SkscaM3aWYn8GNeeio
+PfljMjNa+5lw0wWL66PUQRe/goZmxQGCvwvf6Q1LYDoffzFJBdMteVkaIjvMGmLetOh2n6AF4bx
zePZgk1Y0nIMe1i4DOO/jT42o9BAG0u4Hh6ySXilFvNd6e7VY2OmNZ1Hv3CsLFaOH6snd4czdXsd
HHOq9cQfOIzuwPjPErmBgVcBm9Ennnr+Awdny7PK91AbvNHfunP39uyqUfBIVbOyC4bW6giP+vj4
ytDER30ezZN6R7lV0IsPTXtMK00aJpMOjBayKX29MtP5nw+iDHZSmVDe8oHXa7LZIuyGIigGGJsU
ByBZ0oYRrZrfpDPCj0WnGEAtcNKq2gvuMCZ5UwcgTrRWflClxl7il8C68Ww6Xm+jKnwXAldbmKJH
TNhRF1aQksmaI9Gu0DMD6IKKICvY0wKPScgpsMGeMo/4eTIAMr4r82a9b18pOF8dzQMyXavDAWuy
w/UMNgdkpzVbMKHM4O+8fe9H77Ccj8NfzOchH4sKR6U3RnLo5dxUO8YM0Oxidx4Z23yuGAtjM8f6
7whNG9nnOZhgUXsJc47ZuJjJHVPO0zpr8lJvoCsVfBQvpNqB0iHgDfTPSccecHF/HXO9/goFCuZ8
KVDsfXgMBXNAyuIGOHO3SNv9xPMyRpLNA0SBPWhAm9IAsKEKQtIuXUWGfguZjmuXnPtyPLXVonaX
wzM3+wfVm0ObAf2gmcG1Acbo3w7yqz/Kfp7yDwncJKUQIRyDdAk0tOAzUpqZ9QMA4UN7U4PVpEaZ
16oDqLGCwwBrqlz0kFIRXuB/kZovaqwWzAr8AmwcAxxTMWWCIktfBpZzJDhWZVZXaHrtLk7EB9fO
HJJda+R8gOyDnNBsIwxKJRp9JqCEFX8s/QdxcUX9MAQfj8PR5rcIusB/rhaV/e+G9Xe0MT9PiwRd
K9x13OfneIgQ7W91NixUwgKURHTLGmSuUJYF5yKCan4HdK3WDR+mdqea3vXbjjWaMwPzp8kkJlka
pw6LuZCjQtFQwQUO6R89DNMYefTVww5uXt59rRZPhm7w3CTWfAXqfP/PdZVydq70duBRszH/L714
A3TO5SWaLnTjmeg6Av2NuqCuvlAsgxadVlU08YO3NRAilupB+nBN7JyFkeHpZZpkVPnvRTf2GkrJ
C5H2VlDHEPVjZ39mCwte7URvnhmbffrBN1nQis2C9fjOg2PMeuPx1dNYkb1mhX5s0N3X5/E/XpR9
5NNI3P6D8Z8mjDUJq3I60V6Qb3rDxBrZL0boi262xbdSc5EEEsZr/J8nMwXjPtWAyHT80t3+6Wxm
A0Xiktz7RD86K8vzg6xIJF6oDXyanH0OjErTS9epKvb1+zm2JVhgrBtbSrBwMV7Mbdk+J09cDnW/
JpRzb5YKV4XtiMPQ0yReDFv7gGTnIce+7hjDtTgXMIT7zj00cqIHVfbviF+br3qwNZbdjfbMNhgM
lGnz+88TUx2CzF47uSxiWzKhkboAM1ygfCN7VN9oU1tzgZBPXsc71AIziKCQO7B8RBOLHBpGZTr5
kMpS5QozWFsz8nEZ6edrLXE4g6aK9bhAcn+aUzZ+ZVJiS7XzkVBRwnz24rKah9pT8MMIZ8u4eVlb
C07ujIG5AFoJetOuELYpZjYVg5/Fg4mDvg8NJDhpNHFQbf4zKXKztGVFPcACuhT8nZ23OK4/Rtw/
//HymPbxoDwSOnYfccItb2kePekP5jypQeJdN0WBKLaD+z7U90p5hNZtZq8fI6wI/yVeOZPczeKu
fxKYo/De3cdfFzBz5j9ZjGaEt1s42DP+FhHEvSAgX9jV9hP+gjt9O8qKNb4NRvoUk8qAkVganq2l
wDOYLKRZTa5fRvtlzx1Xs+EzijhjBk9rxyqO/jSKJ7JFwqjfM2N+2ObYVHtRb2PczaxzKVd1iXCS
tuRO3K+mIq7l2Y+h8jy4KfDUQrhqoJVqnMIsLe8ShBRRwrM+Qi5B9qT1kiOVtulRTMKbNC9d/AQr
gV9NhZA4gy8e4xg1HSrvG2YrwEpjJv1pFGsZzI+xK0BElvFta6hMSZfjQ3dOrjDdzLvyb+nm5NLy
b1u/EUxz73+GxsE27j8sp71RVcr0TNzla6h69n6PSL9unNdVQODGaPSi3/PCEreS2WBSjcKUNawQ
CzijOy+FRsOtY24Nns97iR7L2LqTAeIJEQWNdWDd8ipX08yc7ZbYT/nb/It8mRRcL1Pio31ZQaRl
9N+wZjFdYtfHzWXNF1wtpCYynn7PAwgQmAy2AjIboLcZttxKrAFf91X3o57Sfh258/rsW/vIcGd2
oLo/hjuDoBl0iDQjn7l+cPEonX9UkO58/1DtUqMXn6QhOvK5nR90hDVxhCuuqnCMgQdf94VY8t2Z
tUwCcjjtHUogItgGqttXOl3GYUUGMMvft8duv4W0NAjha3HOikwVvUkApxlawW7o+0Ft2jpSM0Tp
00lTpulb6rWny00o8X9JNJdgr9n7zQ9qKG4oK1QF5FEI+mnYkm3t6a1cUDjLKvMu5+yEU1jRr68S
+ql9Ugqcncj7Ds/jsoqXnL1+VdbVjeIAECHtSqWnon5BhsihRAznyzeuRfiIgVi3amN1x3aHzhYE
xL24F4/p+M+eKY7rDs5psPgZ7aWzegpMxyA0sKI7E7RRgJaYAQ1ZeHjRTSbPUD19SpdLfppiZ6aL
AKLvs3W73y4ED+QfT933hce24S7Sgpf2L0iq41P0aW6lOdeg3n6F00lP6f9BSdSHHFruZGtGeU3y
xT5UH+p69iYP1L4dFq0KPgxp/D4+Xmo09FzTeakgFkUrKNz6l/4FVR8RqcyUKlrTp7Nla6bH3FSp
g+D9I+jdu5CChhAqryd19OvBN5F5SkgJStr7WJyPzrr1MVYPiPETGrUUfooFd64gPgkdLixgZa25
N1sWXxRVt6G+v+R3+mEQ+OETlWFF7Lj8ta1JxQ9IYA0ahwtNRehb2vIl/zED37JyU4l/s20QQQKe
fbadWoul4oMUXgXFeu1IoKIfmGJeyS2jhTtqOEzDwnr2l5yNtQ+ZilBMoNS60LDWnCqeO+DEOi1M
Oy5S9yDK/RqeguLgeDagBvljrLt8D9JF3SucBL/yml03tpUuD88mqH8M97YAWoCPmMFEKUerCgNo
bVmydUcSox3Fmn+LtqeG0PVHOygWLvEZ7s5uz6OPl1vnWr3W9tMdf+HmeXdnk4bmjoIJHmZoIPfW
ORv8n2XGo0k6mNfUHgvF+r14qNgCUA3n5ninZ4F65CgEDJj3c0oDNxCgmOF8J0Y+i7kovodDLJR7
/KFPGTVuFgQKS12k7ANPY1TTl+bKX73DSyqGk3cAf3KETM1xXaWpqCvE3IjReRoSF/lfWksvKOi1
qRKkc+vf6qYCVwHkbd1iM/Y68/htU0wX4RI5Sk2EPWPeAQchKje3WfU3VW59TP8JglnkZp9XR1NB
RCsBLWDIiu+CgvxkmBzY13iHj+57dO4u4zXDl6Sj0lCqH5IkaYrbBlpQrUJXN0LoG3Zf0WWPsUyF
Fh0blWRJhT+n+pco64Z+PXj0K1AOQEU9G5brKad13ghh06Uy6skr7y7XWT6O5Jidcdm/TAdHmmy9
LrlwoJV/G9knGDB8NtO4BtKdJ4RhUbLHHMRUveQ4d/+8xXKoQT59g6FW3ZIKeBmFVsSzdlAiQ/jZ
vNMj13hdOhCa0aXsvGzWzv3USsHwQFp/UJpFcOAzkM/jS9RHfVKQWBB2Q19dkdCvBqPMeCaHlMCn
pgLflOlZH7/rhdNoonJ836361aohfSfwiEfOUYx+uYdIcN6HKxOoPu86VVnqGiPnZX83QeMwKvyE
FnXfpGviaBYc4lAlrC1mZC7R6bnTGAgpBvSit2im8UUJeGmRVTdby0YnnvPychL/GSV+tFuFMEXP
UKseKB+42PGLwYpEvvH2QvQRDiPm7oaQyVQ4Nd4dLHge0VNM6nFidh2oZyQiQZ8o/JCfOT3TewQp
aoyHkVaSvAYsCPcCiyKEMoyO+8XVNiHUcXNWrHorHF34tDKitUEgr/EwlSkJvM+o32DI30UiwDU7
Omyo5QRWiNZn9xvJq20n6njH0rt+6KVxY/bLKn5MFBmCV/VkNvTyLiQxUnVurbLZF27l33x4eboN
Rjqp5DJICtUJGQ13nwbSQug+f+yXRFuNxJ6Z83JOliO+fQiNLCg1oyZnfs9AeijR1gFhD/6TtLxf
xuO906xDco3Xy0+gtN7ts5vLoPSGz34CZotpIL8GV1jAWuSguuY5P36F9VRLAmyon6Fsj+DLKPvb
oKxCbWgOH0aZpUgCdalTGBzDvMRRPjxALxdO5o1X6Ds6Y/R7K0nOHiZwmMcl92n52fEuidVx+gKL
Wwb4psy31rjWaoh/5oRYnvwPZDIRzHesouprsW3O3tnIto8r9dEiTuZGrSUTgojnr9QJ4N6ZEo1p
YEDafQECO73xQLCKBCXQJkhcs0J6kW4z89BgcjWDca3kiupITWvMXvHFMgcy0b2yN2VIISuE6VMU
cccfhU7osvhp8qByB7P/BoGo4BpYp2vsVgKz9XT1YidHlyS3f3n4m3Q+D+71OMLAPxlAXbURbYK7
O/cWS5NGaug3L1GcWBsb7rYbR81b/atz23mTnV03cANxOwGHfZBkO5pvkgjqa/Qc8HbCI3+rcqig
6hP0Vf57Z589A6cQ4W5FEzYUrSiEc22IrJjvw22r0EuwqxjG/fRySIeF2O8EgRYcwhe/ZLVyvW35
b5suTEM6Fdvj0JVjIiE+6W17ZxXzzB4tCdPrB58O+w7jvuW2ssFck6J7G4y6GEOxYKAxp9nrF80/
TYcyfoZVPPSUzAt6yYXo9ABIokDXMIEg50NAtO49sOxLLB+QFYfTlTQifC/31Zn9li0CDboR2ujx
7Ql02MMjHmLLBW10UKIT+1RM3QOxxDticlk6hJQbeZXKH5A7jl38c+sBuj9lvoX71MN2No61UkYH
LJsHTBfYEnhMUIgC8O1P6v+B8EafF6OdxPcgmBlGS6ns0QT+vgEilE8zQ93boViWb3xzY9qNB4Wo
ZMc1n+njus9mXyC5q3CGezLJApCBWQJ9jOgMy6FXzNjEvSxzHWR1lKqNxy6CKjOoR934AhP/MZei
sPk/9c9JGuX6uuP4gorcwuwD0zJfZlVpStyA3o3iZ/BlTIEmrenvqjZ4t/V+OtqHlC4ZwCaSPXvv
nliflWkM+OaHKR0hh1GdVm1doeJew8SSLo0k0RITNOKWytc7OsHUzHiBn8dOEPiZQVkMBirGbCtF
mIhdCPiPwYjdwFv3+/9vGuMJAMxEspDEO+zqs/cKPUtLLVyn/tBuCTKMnhA3UuB3wqG7zQAp/9ui
OtKb3Ot5G140H+v3LRX+zwCPDcR2FV7M1jC+OVEIRhrrecdFCAiZ1vNN2GfnioNGglpsfmeHKI2u
Qfc6MiB/p0vgf1URcVfqLEa2COOxqkvuraYl8jhKWPgaslI0kiZOMv/u9tvmeqsaoLTSuRH8TbZH
woXJyot327yMiT6KdZezgIewGgxS4DTDGgsrq6yoeOOS06dFCiMIn+3IXfx4GxAgyEhkz7T03txN
W/dUbAue3WnUr/5wlF196Uvxk+OhybSqosNaXkpwpwz9VC/rNkFFgLG494WZ7U3nms6e4fQQkpfz
NJCcr5f7JEXWzfx2odwk1grSiTMBPv3RDpaXif2IvysgTPaqhrVljY/LEx+h1rbPwRGWlbiAWlRR
wSFuzEulIeBjPEwLzwE15QMHkFUeDi3/0CQckMlcZmz+DwAR67G8XoxMV2X3Dz1mEh1sbq7GtKq4
Jpi3nHs4qt7O0BVYi8sSzZWi/+SHNPcknzUmcPF7nBSzSDtNYr9pq9YzFbiXn0IsSnCEycbjKclw
Bh8DIPs0X1k8vmtOgK7bARO6q+B1Hdqr4+SkAI5bS/vt9gfUfPtf5Uvi5IDxhOqIbZwh/5btpWQR
x/P82dmz1QYakeMwLYpNAhVVSmMrhuh2vxw8ryIQpRnw93xOxu/Wiy2fyKpIu7PzEkpZ4z6DzJNF
Zo+5prGeW0VdShQfdClbMx8/Lm50q/fTUI0Msh98asoCbXx9atlYKzMt+VU3u86Iwtz7wM/2Xyuk
W1z932b/M3NKgyJMOoFRmPzbh6aRZ3+u9DTwgCG1kVEyRxCT6oVQ8UKGQTN6OOPathOSDCogG0Xu
xvnR7h+oRE1cOji7lkMAdMgyMMcuTqrjymZWTDoeZtHsLQnJSlnzp6sKuwmIQtprrk9dp9oGNijP
eHKIcxn5ILu3P29bUeYMmxeohg1NRzspxQYLkmLMMKPwCNXVn8E5+qKa5MLgPPHEb8xeRr3/JmkS
hLo3JG/ebXhIiQfKq/SNQUVI03lospjYStePGgwYzhFyPYe+6WO906YrQVWnCUBmlGL7bVQSZt3+
utjUmvyI5kbnAt3u5YtqJKZZlnNwNcZFXO+JM/lydVYVSNCoUXt4AB3DMJAW77sgbZxwwfpzLSRT
Myo07PfAyyEIhNjfMW47C6fjO8bwBUJnZqmJ22FKKl3yOYPUT2W9fnaTZoJhnVqGqNfy+TDk/3na
Aey1zF6xUS2zW4q5fAV6m5O4lP5f5KijsE+/3aiOhSf/xmBgGLQx9jziP+ZYp5MnxQEZVmD7YLJl
MaPk6RF0WcQfuP7DtF94107aoi4Dq+K88TpEXmVlL/xudf5tbD6WzfdpLXAUB/MA0JzZ2RRqTN8A
n6E256DGy+806TICIaLjtR0T5JVZhYbjLit1lWTzm7UVj5j0m0/tloJUKcBCqjDt5MTo2LrzR3Qb
vSBvYFDeWxkcEaDi0TrIVWQ/JvUQsaVugdyIlxAz+IvYOuamdNum64n9d+Hz02QgANpS2cpxpEqp
o9fxT0Iyodp+Be3fK4YW7RUg2Uxl2F5UrZErSC0+SU+ha4RyPAyzt+64jtDKFTfLlR1jOFWoZ/VF
4n+03Y9eD0jK8mCACDZ/AWGtlsmtg4jRA6c1zsVEtKxAKFOxSAFIPBwCPnV2F/9J84GWetgBC4lL
3EBmtfgDKjyFWM4iEx43LekLaMYs2PrWX9wVCDpjFJHYpRaffB9wHfImt9/gV5I4G27STpa/ifky
brCR5j3A8mZSVrVd27brjvbeXpU/BmFhDyvQVCHmgzwBf2KFYcDGcxMsDrlr2xDu6gjZWYZ2OM9L
gjh2lK8MTEfZ2ChrtBy20nrB/46tuiFK+EyK3fxMH1BEFgJvKqCMMY0m8qMY9eKnfzU8+pTdKI2F
x6jgg04xGPNCvsYEsmX4ilJx9VY4bU3j93H1gj+kuRwRVJmjyVf/GTe7hSN9LIhlLmHgxUSgXzCp
P8AonFPy4ypLLuU3e6SVfOJqaqiQRVRhgnDRUrGK058Q6Nv4Zw1TwyA2etHY7gCZ7I7E2HX0VJYH
INvw9+rt+A5i4ifCSkCtVa0z+M6Pda7y6JLXUCDA0+VFC6tPiwS66RCsTcKTuBrsKjwmBRkD+di5
AHY1XzVSsI6gvGNAOoYFlAc+Wmti9IMBNq4VSMOMDMwZpme1/iohcuyzPbUfwWEMqpF/uwcqWf5j
bp4mjCiuGJ/oT6tU5/UKFgVv9REWha97q5AEMy3BwYYCGzxzI7EbcNGT4Py31gZJTPRCqlRZ4otX
MT1cha14hyKa0Zkd2YyTCHubtoSHNNvHX+q2RnsZFYECIhiA8Dr6mB21iKH2I/RP5NmPg8oHHdYQ
vmHOULb7ioYbR32VAj3LNvK1mhmqjOFWooKrGLECbbo4OBzX/isbjvZXFaPCxi2KO1g6c1R/GGdr
MhsrCenbIDdXPauDNqyxGD+IpvW6l04GJzMq2hF6CnmzLzqYPeeZgLGqldF10rGDY/anJf3/7U70
0ROnCfJRsgeI1sNJW4K6uOIedKy8frEXPamGIRDpRPj8Bt1xyb012G6xdVI0x3ZuF5lKum2b66s4
VDwRkoGkCfgBKAMgK1wueEI+vgJK+MMmJKMr5u46bQhpQL07PH3s5rzhRKq6gWE3grUSDJAOrQZa
eyWwarEN6vuZO9i3C/rrMFJwr1xmt+ter28W9J0/VDxN+K13ujys2z8K8jx1dNSmWaUVgpWNbRPZ
6S++B9s+a1PpG0MduPxq+3T4wSO2LLHSxDbJF/qnKwwywSM2oT7pDivgKslFVAx316M/l5bqZ7n/
wROSGRZnHEnwwECmiz6Q2+z22MF00esq5DPq12homGeiWJGer6Y02kjJCGYJu/TIYrAWGfrKZk6v
RKvbFRl8eu7Q1cqndsGaPGziEwGAqsnzdMqTdx4SwLue1/40FmK1Is0cv08U38S25pzHMDlh2aYA
hGXw74aoa4Ze8SSre7n79mC6le5IHUFQiCGFfNr9TcEnFYx+Rhtg/cpq2yw15qthXMNkPgXGK5z5
S1vvmpoWxFeO7NYnu7Bn1Tiw32Dkz7eFxwVchPeu+Jg3FGXuwf4jZYHHq9bOCPVzMmAokuDfUt9t
tre+1sfZNcUSJuMqIaiRA0/Rdrg36+RumH5fcUVxcyGDaQ4lmDGsQmDCyMnm3a9q7nYscyXsbCRP
6R+ZRwXMSatQWtl+asUn28s2I4gtJWzFHUbwOIAP+uC9FTSwGnOPVvFr0/rige/a4swYKHcaMjFJ
bQQB9acClP9QvrnF6+TZ+379fW/vavgJvR295mlhomz36BAO3UuToKdjWXfGzRHqWbvsrA//Jw/j
8ODWlIiHutO59OSs5F2ybIhksA/X08W+mj6na83XvRjRUNEIZhJpRix7kL/0w/61IZUQxgl0oG0q
iry0A3Ba2VOAmDstqTZxcpdjyC5ePjyi+P6C6NKHQVaS24d21dSA7G2/HWVc2GTsbdPdrfGJbeEe
7ysctQRZub8VNe9UEw60fCtHhd80erZ+fUtJmSW+O9RURWy9BkOSOGdpJlnIN84CDP7r3YRy7dpI
dKbclYBMNjMvDLk3tO7XYKTeYkcw8/yGw8V9GfodKWdpK3pMIsAb730z9bjEESlYJHuHa+YBnUhA
3EfexPUx+wOJyndnU+6C46xvTz40HZ0XRQxB5Fz1qEJWlCSjYYAO/EwiQveEueJEfe786ubazVl/
NmZlr8X/KHAJVbioczJDvlVG98npwy9dajLKnUIh9hJZZLz9U5kTx0UmDeBbXHpFnht6aQVqmUq6
ihXyV6ruTRpqIMdi5RAQW/XcilzLHIJApNF29OQMAVbOK2/kFTO0Cdcz/NH8AG2xpfuqq4imoCBi
BcZV40YcrmDQZimC9qJFdcB3a20skTP4kSlsTGYTOeydGDrekeowZzJgXlBGkAmG3r+PVT992w7Y
E/IJPGymKi4LDrwBCspImndF0/PkBjt7ERGiBZ7+Euk+iVJwc2ASUoYcVboUckh1fMLGIWm0tMlT
/zbtSpGe4bm4yxLqEaUGC3kJ1dVoYrCtHoe/bERYnxw6aFcIwf4XiUfhHUZfg1GVX0hwXLjeQkzQ
qN9/uWm/jSmkAaR+SlYgJeQzZW7+WazrlbvlXl+2EFIGzxa3XN8yFVM6mXuXLwwLuJNPQqO0VvPx
U1fCro8gM6GBkALQ0uaPMoC8wgstb5vmp1kR9u68JMBMwezq+cZUoauzkCrTU0fZkBk7Prr96id3
8WLq93afkks49P8M4ElnEIPLWlh2iffAt1rePib4Y4xCRvfnKt2JRASbexlacatjcPfkpN7dhOF+
iujVvBIg9ZX6T3ic94mxOmEs9i8olG04/RCeRoaKCC0ME+khZFCjsbH4u+S8nMOAYoROf0GLM4yw
xqhHohCUlwtE6fps/W5SQRf6Fd7TfC00YnjHW+KqqWbForvnKzbn/iBgp3WCMetq0r+YCWUk8qN8
1KTjC2lqtYpMOCCgYNP13rVbdC5KkPpsq30oE4RmiW7EvPGY5Id8kEfOK02saeUAFsZbMvo5PIVR
lto9XwSpu2oPs0LvHiLKMaHEtpopGne6TQnymkAwkkLw2IjWg+YqyCKXJvR+rXMDhxMVnV8Ygr1m
u0XPwXb/rdIW54F8dzaZYFCrHfpEG///VqbH2y/IQUes8IgYgbIL9+NXgYL4RJnhakxZLl8qwD0S
29F331qmY53sC1y+HV+Iix4tJmcR2pwLrpmLsN7CZoDq2CAafrM2FAlXFUvSTjirEgd/JgjXtNy0
L5rI8B2O8HfNlP+dRs5hOC0SH9H0vkNIT/b8Vw+rkm0xLLQG4bq3PdaMqJZYVvZdKj/tDWe34MI1
pbcf9niBla8ila4CvFIRl1QZZKPxo/1dQUrhzJuU4rtYs1sVCV+ZHnaM7wu5PXUvYDBtO6x3vc9b
gecl5EGsxiQVXP8ceGdfeOZSk678Hh9CgxiaGZHFtlw6dumISmZV4bitKVAwXfWFp1sp2vMVtzPg
zQxyytRlspT1FWd4xv69Qi5pXTpTdnu5hW876dG1TO7huTDZDvFjbJ2vgvgv+VfqvbRIGtt80Tki
aJS8k/57Pnitq78jx3IP0wmFqCR1PxMHyxscd05bzODnw/AwAebhXY5UqafOiAu6JSjB3ElTk5jf
NC0icD2X9Xc1j66bZZB4hm2gWh0WCBsd+MaiJMQpTbLrWsOWsvwuYRwnscQmqxfzOYLLGyRqkjkK
YBondfepoq9VWvKmzS+WhkAUeFZRSwmZWRbppWJm9zBbbq77FZNyiDKbgLLRigHI0LvW+hE2JlBR
jTj3iVBlnxlcoHFAhjcyW3FKbO1ieCO1ejkkHmYnLLDyKfNGa/XhCG52eg8xpX4Q/H7qXQohCphz
gD0MIY45pH8FSybXzMwiEnyzOnIphBYXHypa5b6QVWtTo6Ctf095mRz5znIqpCr7V76HZOsPXQPK
H1Z8NQmUWGPYBwGO/14RMiWpxGKFRRxo8q0GnwfD5kdOqROhTfTzfLzinvOtoAcmZsv9bkhzf1wm
g4MOFESzfQcjbkRF5yy+t2HKOlvwFOYS5FVPTYhbBmD+Mw3xu+Ay+C47yKKBzS9g22CkuCbmoAP+
HzDEzW+1pHrgQt5BHbj50DcHIzbxvV620scqFlP/oyG4vAxUVyubMg2FlxMIjyzTy6rhMekYUnuc
KXI02mnhzw85gs6BwxNxv+hUfe5MTNc9j1w5v3CmUhrH3tJX5xPSe+JuRPWx7g/jn9IBk5Cwx7zO
YTliS5GK0bP8zh5FLBDC/YRaXNzLOf4mc+1FOg63JIZsFfKkrDeJ675LWD1wAYaKHE7moa/DWwUA
euvZ9LBesirwDzo9Woo/aJzaHFRC7htXDsbhLq6JrL4qFa8Xz3BZJVmCKhpO9NuxVcrOQ8KQWXE2
rHZOUA0XCC8T2gtoVeW/hWI0hIgOWnOFA/WxWQRXSWFiyoMBu2ELKg6u1L/QxuryfAWRUH9peM8D
3hwdoiLUlwyMdi/q/XcmgauIiIjO61zD77rWVPmSlKRjkjKU5dp6hEjv/8vdy/E5hV8eWPMWN80t
ZzxB/cYu2q7hQiKBym6tDlYNtk1Z16TKQwU0PBLZ22K0aEOgMxLCWzpD8slKAsYF8NlywQHrsyUb
AV9FXMypj1SsXnLagT8HDxBQTutXQn25v359WFjXebNAmtlFPd/5uqWclQs5ZC/jGBZ0JVVaijNt
KNm2kjCYmaHsaXqrucz9zUCFcfJffr0BqdD2uqbtLQqHA/br8xYzF7i4BGdR+8KlN2fuQzLtObGk
sbien/2HM9VcdBIZJIQNoU1aktI0g/FXHFM89aQoAt0wl7PyB47NMLlM4/L49M4CEBlpAJKN9MSJ
Gk4N8JBuGGQz8vJDYpOD9qCSVXQlgmOyjwBGRpbfpKiTzeupJF4AOaV+gdccoNMZHjx8fu5t/uxy
FJ8gcaIAqJDuPbHQNhhovud3H8KKHlCdEDQOZFhmOnbt6Qk5jpEmDH0eVuBeWZfa26+eYMZ1XGPT
8PlpPMo5A1w51zjhOYiVbl7J+mn+GED7o4mKsKNkW0kzf5osS1HUxz7LHsRSLdtSaVMs8jom9m+q
6KzzmjRtru3+hiSM7UgowZzc3HM95CNfWkDZlra1pZvTO7vVKiZCKDJ+vrUHoxMDm93zr5m2qsQZ
qsVVI+MVa7SGMe6B1lqo1sex9xhuunGbL41rSkQKoe6fYcTLDIgdYEU6OJ/RhWqvEEjtspvJRmZy
+RMO2opqrtTWxJaz38lYpHxuWU8RTo0P4ZaegkXMMKtJ7+OLeCOu+u9kRjIc0E99hqjj/uH49gVG
X2yAS6AxnyQuT5/Vo7tg3zuu/KPjH7y8hO8f5yeFYIg/ngcvwcCEiV68C5PYZ39ztA6JgMSKyFjS
iyE6qviHxB/QTk9T7iCf5FCVXjYAkFRna03KS1cgDUBdOWsM16pOvUoHMaCoALtiCPwBsuk43XSc
CDvABw8Jy5tkDNdWnvTR6TBtjK/OSr+lzQVfdhTXblbA828D1YUCgYy2rguyt+fPad1V73w9yDKp
h8iJimRsJQgH7xhC0Wd/iBmyMMYzfBxJHQdAh6TmauI5Mb6+hUqvQZMl9MxCmZq65fMbs2slrHLA
IKtWCeTDr1eEL54f0JHfawOamm3bTsB1H6dERRg7FE/N7KyxkrhgHLAEuqaReVwkg4bFuwEIBNne
xEygbO3bFQVc6cbzaJ5AYQxRiNVQDYY+YPbaIJ0Nio29dkfflwcSlJ3OBUAuipXWJ2iPxkjFjpkk
zkj+ot1vbK070Z2WdPpgdGFNUg76UfwCOsXGQe1ZZMsTgA03B4kHJFaeMNwZAA7bkQ5bJpuZX1dF
sFpulew+SVNLPDuHUWg1N22jogOr+U8ytxkhzHgNEco+iddcJ6rtBgA3QXTxIILHD53r1n66QtV6
EjJ/nbEq+W5isPSM7XD8bYOMebAm4W0ixwgzX3eMRMYL7sIGsLHJjbwi3iWCP+9LV3wgGcpZsq/+
Ue9uVTEGGjk2CotDPFG6CC3CknF2c8M7/FuW/uXcrTWa4z9lQb72qk8kDWQYgx8GpdhYXFQEE9DO
/glRNaXuS0aBmAwwuebnKxrc8IiwZMIuu3vAtIkoCue5177ZyYmh0RJ/vU0KDyJlRbRVlaBb87kQ
+yJi22AhvMenN87DgFC8RnhgfYF6zqyYwAK1Mxh+Q3zgo8FTFIjEctNwD27FAZWqBNo0k9SYRwEL
hmlczVl/fuWzpiDIId1LJ6iI4OVsfNxbzdZLxxZ7lAUyG7VqIgx1da5YBf6ep200YAUPSzFeGHRX
KYshk1wmbfHWsHwPkxdBZbjo3V4LRD5/Thb3DXxRe3zupRbEAGfaNfsAUkJjTcwqAmf+DzNCuxHj
KMw/+jII0XoIA1Q+l6AEqnb3JPpAhUQhV3PodasSA/PlWewLggMTIxi0xXUKYKxDfneXMit6Rkd5
Zynj+Ao3GzUsq10avM0bef0qgT71DEEMwzNi/2IpAuTGCVyfUQwVYNRhPQeYfS89sUiBKR0HkPH3
mB6GhbphB3NEOseASTCJI+y93nsPCHDBHvZ4379JqFfvEENb9kx/mMNRx5FIblNq/tT1b/wb7oKG
3wIGfIGKQNaqm4lx2oSUU0MH3bhdaAQkRJeHXDDiqRnRLQTnhosckvZpG9TiuV0aX1GUMVKT1ci/
Z5UUcldMAr2ZMAnnwUTszsvHylI1bIwgdlXiOjFiV9rzC27WY8AzxWbFEFIqhZOTVt4gblzzbK4H
02p5sOqHfm9rE3Srpnfdcoa9fa7NMYmYMtE8aBQ4GN4M8++qjaMWECJNMRuSCLdi4uT/ptFHKbCt
kKft/0srf1Sf+YREoBr4gh02W3fQD3GOZi4mMt6uXnVQqgcZNP7J6pWA+6uYgdz8TbX6zIPO6q/X
1yJdw8BPTOvQuih8Rgy/czDeX+ToGFjLvdxm7fdwnEFpaExOprcBU+SvLWF+qi6aU7t6noK281f5
/WjB4e9HaAktF+FX0vL+Tieyw/cGFpsi8Qwi4jNQRjZeB8J0+yONEZjV/BEbowzfitSRCnqR8IIq
L4Sph7/tKDikgHJES0LgugTcyLpjBJWkvWtAGWbk0AewgHqBzSEXDIHs9FgcpnFbyEyQz/4k8fgq
oh568xXYad3WaZhSCgJr8GKm6YY+7yKsgPDt7PKexC7nRsCnpndxQJu9/3mzMXAWzF+MLjZNt9Yv
AsBBG8oGXY/nnb5Pzgpb4//ZMJHlLC94X7TGgn6ImWOw564ICXcn3ub9PrqWq+ECREkUchGFBptf
M04CMaEBHM+tn7gwYevXIh/tfBFdPGy7mwjAohivHU0QIau5MM7dXmjed8OjlzHbDkq3OvczXcHm
8NqiisSwynjRSFTliAFPWMFvcM2404nh7yVp5oP8GeflnNg0kAu+bTf63bIlT/TkAFOJ70DNd1EP
F8fAa09/iC8JEynvEbapPN2cOckdyiwmfYWeWiSL3WX/yPjvd3zAnz3Lvq8p3xmXMZnJuS+mJZAl
OGTZ2KdTZOAT6f+atLrdlXvmk+vlw8R49kuH7bjKKcnidTwia94ViZivcHqjFQZWNmEnOaQLOXKx
rUYgPcfyjb0PS6cyji2hMA4QTtk9JnhpXtx7SeJEXKCxM6Z/1SO7fljg8bDDJd14XirCdeO2AMq6
FJuhZvejpI6ExPaB2zhkQhxzQP2+E1+vHdPrPoquq3/bVlH2NwhHMjjRRI/aOaRJLC+6Ae8Gt3ZT
8NnAjb47R4q8x78SpAMIU+braH75rE5RVhtX/lOAbvfLmiJwWOzlo2N45IFG2/ZLrlcZ8zmHaUG6
ru4R+MXjg+RGhFA5m3lMfSZKwP3mHOv3xpWm88km0Jcce2GTqwKExp09UgnfA+IWYoRsk/cXXcg3
DryZAEfeECCt4S0pFMfiBEmyc4LUbMidgN/dy1sQ3xLC9zh/qmfZqSLgndm/vZruSEplylcRWjW9
IbJ5yzbFgIyyDs9+v/rFemtvbO2mwbtVsKwcvtZgGFjZTYkl9JM1dy7jknaZPSyMUpK1Zw14vLNO
yH7TIZi9xGqCGxuKLf8Y9u2HZm2tXRVMF9CC+rv7HPwA1yhTEjD75wHhTgNFg5XjK4GxdAOC7dgd
KOUEGFQKN7encrjhhVMvr553udzTh+ki/kGmpZlEpJA88bnTBDA9gubml8VJP2P4GQtEkttwen0d
jUWNI20KySbx+1GBnixEcJ7BViyGxAI7rxPF2wPcixgCtdlHafvG+MDYoYgo8hDbHlc+UQVW0z3s
1+C+azAsB5UyLYtJaOTfClPlXqzUw5Gdlu0URiusRBU0xXFLsCJTxeA8NKUyBY9EXfCUTAP66m5q
NSUlm8XyqAap2gPTHcicLNaMeT4hAhb/QszDhfaTQmCxgo0wb6i8pCMtfwrXmMWZClQUgbQjn2Vu
OU4UO5Z4lHnrS9qdoz9gthhbM3Pynio81F/qOtsZFNwJ08+UptViIOYv6DTItkiP4PBSniK7BDqp
cgpFkKemPhMcqy7awzxq2uEIFH7GbqYTo2HEEdbQpET6RkBQDYa1A4Pste56J7jLwn0tGjalYwWN
IRbrd1OF+jMPMgilXx+MzRZUf3aEp5qAjpkcut6gfzUQjpe/DNtW5JDocpU1IEgloKYnBnoRwx2g
xEyGNMIXM6wQsZA1unYhL/+InDWPvovZg/8GvA1ngtWt6K1RiYMN2IhxpgHnvREMpuXytJOSWDWh
lqfyaR1eqvwo7PU/wFITH6dD/wPypD/7hBgPGrZbUtPg6G04Sa2A7eI4L7P9Td+nLzvnVCjKAunz
T1e9h1VJbsfEvIbsrXZLc4xZECOZbmC5zfNB/K8fdl4TxZEqyi37YmV+ecovqda78h/vEpoQp55G
c4STs7WaIVZHhUUzPYmOZAZPvxZHOxvjf+WIAu0FnFoKZq7RbUPgvuI7hMRIn+vn4dBI8uYQQpMd
rPRl6jsEmOfmYz609mvtoYvzSzU4/gCxQ27BM9E07FUfixyqvBmZYrQZLTtEEmIaNEGELxbi9Ce0
ij2AxVMGPEl93aLKN2wkhlPf/zlHsT6eIuHdBnsXxgo/GZ7WfwBanhPiRwt4h6sNoQX8ftO/u7E/
VqZQBiGEewyAImrF0Z8ZqVu22YZXQqSi2q82ZrDO3zT+2KmQpdv8w4IlEcYHmlGG4JGwJCz6pS/L
m7CtsEgV6yfwPc0nflnygilFNGw12Meu8XkJZOh/zixM5NAuHB13EkZnjNyDEpki6yEiuImbyN/D
huKoGRJoykf6E1lKOUEScJFYRJGy/SYmV6I6aKvmPiO6Sj5AycPwsS3g0Adg2Ef04Sb/YFG3UiNI
Ye7126X63FkFuoiWiEnKYqyyq/6KdZaV0zYC4Frn0z1ZQSubacUblThPzgWnoFsOrIlbKDQQhBzE
CDHGrk/2wxgGsBZ3rsCFiPYj8wWG1YeZfb3zRbwJLnThFiOFZ/YPsvZZb+ZY2kxAPOMNKPjHmbye
KS9+ezpC9v4VA6GYEN4jyOuono+U6nKSxZy3VxBWDGoGd72MPS+XnL3zb0HHiTIi8CcFE/KuMYOG
490AgYMaM9f0RGEhSE7hNPc0YgceypwpD2eaIziHq5y0EMnhynKObVmg9ROHtcGD+X0tRQX57wFR
mBfT5nrUUT9HTjrAWaZCGW/vZT/OdUOaqhUSVRLkqHerzUBjeyHFvmYj7L9lARKiksn7HNm+h58f
6jlPh6r5HCu0NRRlf5IN7MSIUnJePPKjVKkvDXfvz1OdBIg85wLjpWMBEsl8BwhH2dzZBakd3Ds4
+M0XaFBzmQpelEWZLXnJwuAEDgqcc1GtQ7FKhj9fV/heu3YOLRgc3MfeNH4x0wdduOio8t+kc/8T
1ctE4dBWmSK2PxB7G/e7W1OL2gePrM7wf+4/SYs0pXQXktPCv2qgPqG2SbXPyDkDjaZVdUii+0XX
PvqcSNVJC8VlZw3T5QRddIz6sdx2VSP4gyGnjF8FridN00fnaBMIhfrJ+VMVIQaRNQOpTjbBGK4F
lqUEhyv+cIbj7hQrFMFbbH1ZpdIqrlajh4x/Sgl8fSPWHSeie0opGTy3GHwx+d7dos/54QESX5AN
yzyM4pWNNYKuWQpt0WNBtSuVovU7vu/X3seY0WCBP+MjLcdB754oWMVICSDzhnge9o8aQ6Dx4TW0
CucXiKGnl7ou6YGjuuPb9D4+K5IIcSsAx3tXGiv0taAXth5PKp1/AgMC2dYMADaEKebwBuR+knSR
EwtgNaGoefOj83TEKD6qnCeuJ/4/af/v1YZV62rSjfOIGdm3ZNLsBbBlSMNp5z8q1fwuKRIPSpsT
oN533/AyepohtwyjLD9TOBIrUfJVNaNKxd6SXnB88drLci5PrUSpZDYN76WxGGZsQWwcTh0h7TbG
1YieMSIw59m6dEWOdi/6v8ZXRpPiXavW1bwtnHLdH700Cw1vDaT6uAR8KmO435Aw36C2JKDXrJfe
acxXOOs96XetzMncwio0ZBY+POlNKpF9Wr1ILOUnp8xNa42LnZDnDBjWzCOgffxxlnIPpiptnHtp
m9RyBHK8oKDjoT8eAX8NVFJFIDPUSbnsO/J3/4VmqDqTlmgXqh5qQGr42qntCwF4U4bnzCE7cIyQ
9RN/HNhD6gA10XuiRzEK3MmGm5uDGWpi0nAHM4I8juw36r+tVzGqCIlfIWUW9YYgU60ajJTmMep1
1sIP6kjj6epTUE80lPzuxDgs9/ngpOMRi7i8OkHZAJCoXnbhSKtpPb/DtA9Gduw37L9br5khJcmK
NdFkQlByjnsfTZJFUEpTPXTxLwVvJKxSe5Lq05lGL48+MW7hPKzQNdFz2H6pvhOs9qanLq2GLCgF
Lyx3b8B2KpW8DUTOOJq5hW+qYMPmzOi5Mxtmg+cGZnuJpqmicxPbazyZw0Z1LZKYikB+fXntrlIH
bb6G5NWrW0d53Sfz0ESxaQk4Xfo1bk+v8cJlje37potGoOrYUQUrIFpMgYlZkRmsPTwLlFidERiU
8HM4jyp1ou9pIh5QiFfXW1guo8heVaGKRHXJx9hqA1HRW8soQzekjCfYZe7XeS46g3Bxy9wVzBAB
FYOow4G8fvaH7NQ/O0Gn2ujjWWn011uPRHME3ZufBps6jsVbDOgsS2RimBZGN7/xJOT4TR0GDOMX
zO4o9R7qQC6+ikZ/WI5d4+dukZUlrLZYXYugEyn0miXTE+apbahcfOnKUbmRlVPczcl1QlLCKUuZ
NsuR2wwYPRYjUdm9eV/NpZux+52SGCrrYUm7zu7+gVh4M+6NplaYSxMXsbYHlmLkrHyd8DoRtBna
NASsUGJPs5mwJxBPDbvU4bhz1yGyVi017d+dbxSjKRk6mVRucut1isSwGPdlMDuFNs1uywwNHLle
P/yDR/W12L/lI7Xfn7k4xJEZlLvsMqyRD/qURzqNnIzJizPGRrxjNY5LVXBnM0FnrYgly/kCqfaX
37mKLxbr499x3+tAVoqVlADTWs97lLGljwphr4AXMPe3Nf1L0MRskOn9Jx7+iJbVt7ErYER+tV1Y
QEro1bHpcgO30KJDGXZdvYcARwpDIwaqEsOvd3FrroOQe5UiBhiEFiBxyvUmKsWZ54LVfJXr92DJ
5Fyf2u6NdcBR76Xrv/ubZoj1vZq7v+dOz7nR9WJ8XZQ+yCGzNBfNd3KDYIr/ASXiBi0vp/aSr6tI
ra3IsuX37KAGRE4I8yRL8biT/q0r0A9mNsPw/Z40hAsFDaB5zzv12Qh7l/1fnHkFEbMkQfW6MRaM
pM3Kv9U9hmFriJ0USfOcWBlaU4WwfHQAySJ5lA1abGcX5fStvAuvyBSLSlguwY3ZgKNlQsgGHC4T
me5fpe66qj8qnMtTpEM18AuHOZmqxhsKQ2VvrI+B0r8wMlSLWH2jZtSBkfBY9Fsl1jN8G0IvAeLX
6LKA2B7+QmFnYn7dqtG7XTnIv/uZfGBBjWi5bvSAvUHMBHvLUkkCYcAl/CIEWS7HvKnIi9wbolHp
he1w0F6UMRs5/MeEGH1Zm4TrWDd7LIsZXk36qhHLIU4FoTQAj+TmyrCKngL0KZuscsCRXWwKQI+L
2Ckp40ugR6vL8ND+OT0uipTrjiY2+1ATpmoXGsJo7SXM5YeH1fCqaa8LYgCfiQHZnJp7FFV5AvyF
npgANk3jMUALJSLDU1P5rB9w722Bp07Qndh2Fqo9lnoCZVgAEVdWTODc3d/scZzZLLHQcOsfRecg
Sgx5d0hWGS4GOQZ2u+ntkKE1s3YH9tfcrUhc9NO+2c13SccObBk3zwUrnrNRkS3pfQvdq4/PSvGH
QtdjGkJQ+FROkn7xRdkms2VE46yBDATa0xNMu6A/5nWtjxxDuhriS7IZ9anytNoNgkDewYFxqaWc
TtTbBj+RlihHz6Zh1zSigzFlUtFhiIBh3djB7pFKsVgoE8zuBX8QLlzI7sfwDynhInHYUsouPLni
fWLmqFHJ9D+SR+c4tHRlQVlPYC9+UUtHnbUHujAyBfNWoP/oqtPefwUfJlcKQdY1xwcKLiML/aN+
HtJmJrrb0gduw6QCXkcRdpy35GSjYuCx+z1vfFFqO4D4Hn1QMki9VwENWHFTi8b/oL+qJE2NbBx8
5bCLlUzmTgNTKZWWwW3omy6k08eRu7o1ATkCeLIduCQxjmJSkkdqt255VQ785zZRVjb6AOR7xcai
tyBrKT8GfmO5Y9i/z8kjz7ID4inHfbw9Z/x7MBvLkrdpPe30xFjLKBCjqBM4ihoaUED14IiUelm6
ZGRD3r65NSyrCBp/aXDoa0VmOGlVdTDSSSdSNfcx0l7bfPKXaOGutsnZkuN41AmLyciVbOKWLd5j
EsJj+BdBG08GiSdjD0PzsrPLTv1moN2+7gMwnW7GEAs1vI9q01JvkqXos4fZeZD5E5oJpRgowSVY
1XlAcwXA88AvNxrO946mrA1kPDasX1mO+2szPjGAbfYVv2FRnt8M5PjJd+ar69i9+QhRn+j3p//t
t5AZuHQtWNHT6v3V+a6QulilQqG2+3hn4rtR4EoRFKTMZl1JTjCFVGErJIY165AqmKRG7Xas3V65
3+XnRsqcusEVjT403gleXgrXAKN14B8fzz6yrg7PL8KN5tlYzMvAL6SMkKsFdoHm+71/HZ9cdha8
uI9V5D6RSkahCOxjwZHERWuwC7JUK3FzsZj2ORdGA/y6NrsfeeaSkL1JbXD1PGHmWwIEm/jQ+mGW
eYYut/nWiAoDvOVm/9oJ1h/PaPH+XpQOturM/hQ32UaL3iqlO09FvxJ5Cy4D+jd3DxmoPXaIFPGg
9X7gSMI+o5L1OiTYcEEjRX1YA+iG1O1FSlzwPPWpJSAkRlENcyxIwp/+rLQbPKxdGm1G9u3lzVJP
vr5jNI3cxjiDSRq0sY6SbdBNykL53wPK/sardl4Wnk/6htszlLlna7tQIDD0f+Pbfda8GYgXpIwm
BLNiJyVUMpFuGpZQ5RPaASm4adR0etH7gK9c7nAD21UvU317A6qqr2yOWwF2md6W3zNCQYummYQs
yhmOgVyEve76zgezOmPbXZo/pvHedtxNm+TaY/RHMoUaCMqM0JTqQeMILZoznYzJx7uwHXqaULn8
tFT8m2A3LcRqEasq6IHLVZU5Nq01Ht4VPExy0izzFU3rWKUeqWgoBJRsjRwznE39V5B5pM8okDzu
il4/fY8bTfbZUoslWKGgVoKfv8NGYSaPj3VhWk/Bay47qgV6MVEhQJ4GfoOGKRcbAMuXDhuHOtyo
b2133vwnjbyhK8L+e7rELnvPwmfPMktoxnKE9zxQ7YSV7729yySkzRNnpE3vfLm1uhpqHhQALAX6
aDz9hrmQAJeAWCiSdFshDuR2mkSDDpfJtOtX8VwbpA7li9x8ex1g0D26UBZ2NtI7vjjfVMvwXj9p
/AlAbTfN16PmZIATxcHlWTbKWO0aywCqmIziJVDXYZF5UwsrvJ52Iym88IK0zIu5oiLS01Q69fRX
sslZu1nwnwRnKESBNJaTRatAp4CAl3Rha3rNftl6djWFuR6xVt34f4gU/dZ+1z30mrqiCDyoZRdd
RU93hPzIVldqQ1RsIvPZzkflqON9fgn7Yyg4nPnZGEVKa+ecOY06qCyOR6p4p0mf8+nrH9qZgDSx
2gw5oHRCFy0ymQgb2FpgFi6zSibOkNi9X1osuhnPe1vZJYtEkaH1c0BnXowRf8wz0BIe/ak4h7/7
HoOXhvsj414RZb32BY0t3IhxO6wjzNl44WO/FCsfeQdecBNc09QRo5juNdBDPYXK6ocxMyb7Nfr1
w4iFoVCWr8hhiUDS+9cl/Q4YBhu8EMLmLsl8JxECqCvVKunyaCIHCHmrIGFSv+BJ237mqKrOXUBe
ZVrjEUN9rW+mzwm/GwnvIGNNDAUVqSsrsXhJ4pSzICI78NKZ7gdgEyL+QYQIUrBzF3/NvCdXKmXq
efds6EnwlUN2Yi7GU5lEy0yBJi2DbVOsjLl0IsYFd4jmQ+ZmlXpQU4zFYpOSERNxVZsyOWzM0zoM
gKtOleW5/DkNepXEONX7ILxZe14aaGTw5ziaoOzmz6fa8wnykO49uiMwPZDbPmXPdhSpxf6W3uEh
ZeDGaFENVQlO9FkhxZaxBCuClK3hbycumPAMLMFNKRVi4WYq2orwjIegt/WE87Xq5qcVOMQHxQ17
uFEStX0XC+oBsKGxAB18jmvNZP0IaM80/PiSs6nq4jU5zfAQ0rku3TsjoTtK2ASCTEx3GV+OyBUX
AwoUvSRU07h7HRa0fbiX0daUpL8J+7/rxaBxAcvXHcMKlE09leR/dj0YmDBk5UGYuKiz/17TIEko
GtOzWoBp7gwAL+9dGVpEZ9WDM7AAjVpKrQ4wrEIJUxtZWLtr6I+7wWU8dhJTk9iRkpgtsUGAjuOE
LUl9oG1HKIFHuSWCNxE0cCccqeixx1ccpDMRnb33uOGLV5yNwHB8820iPN7AQmOEl4qE1e2o3aOO
FzUiDaHwEmdeuy6qiEUfHZBpKLlHWwFEAbPK0ce3g5Nr3uarm1roghX/GwRJhbPY2Nd1uK2g5FYF
XKoznZZ+3Mjqi80BrTgZW+b1nnfBUdHkB09SIy+RUqVhD562Eh2Clx080J7mIBNrQGveh4im418d
HnMe6WxamrcixOFyYtWj4Qdsh19fqm+bjV9YZwDEcr1b93XSebaGyFAQzR7yrT9tdP3eMZ6hMLNn
a17sSNy4Rbqai9HicS/vjpggLtBmvgMenAFonmLPSp6xgd8gTXggsRaiyyTkYCaaPyBI63ruWc8m
7+acHj2Kz4u1t/BdalAFuuz1afOcnwuHluLRdjy9fObrpYVzZLdIiA0tkDE2MV22J0V0yPqbq04M
MTh1r9vO0YKUpvWB7GFDkOj9zfp4yJOnCjBqTnxCBRC3q3BJq5VKuQGf5UiR7T3+cUFiZQbfx4I8
oRrgouS+V3Ikzeg74u4ZxUs5JDUYT09A+lM/PVqR78qjlg1lDCm/nRawTZiE/VwJVEZz9bwSKzy3
uydfXuOhdxjZapQMOWDRkODThp0/hRMh0OljQRxA/lXqB+SPeh9ddsnIkNIQi1pwFGSReq+bUo82
MHaWtPbRusRNC2fYqk+GqCWTI8sorBXajdezzoJnxCrMQPrlgiRo4fs6GKVjiFwPUXVxuprT+DQu
sAC+21Fslfj0468f9yBOV6D8GHIjAPhj9U5/rIZOj0Rhv9DN1nsS3DAWfk8LvFp3a0eB0Fk+ip0m
ejV8DY9IbmkHQQrnNPdGYieFwiQOQxOo+1bBVQcjbYUnwnfv5/5CwHajLvOKI4dtQCUt+MZBhisG
GAB2XXOTyH1Q/vk4Y8jO1I8qM7ItKsPKANF6se7r6QVDfZI+zxXO+GqzZubbhX45+Z+/fozw7OMa
CJu7ePtwUorkVtcFdqG9SuweR+HcQLXwJOynqQ6c+O0Op3SyrFj1LyRVxjKpfOVZkfjObQj0eX4j
f5iaz6t2dy2RHFnZJz63XQ0AzhFHbtkapbYaBRYeypcEqX0PLdObNt64Qlntu6/FjB4W9+qXDcfh
YoPvCz5Sq57SHp2vjv0AgajBIvpGuX4SsMxN5IupnP1BemaR/dhnVsdzBuw8xkujbcxGazuWKhvO
KQYh+QuEJXc8krS1Yw7xeFsa5lrxlrO0Iqz2cjTLJKwxzlfgXoDueAnmpE1vnlc/AA34JcrV4BQM
hw1Xe9arIyAjzomNbT+OfnoRhzEQbZISPmpX/YSxgiXbm9pWtbwJvN6ot6pjua+lyCUQ4WO/mvHZ
9hycwrgBRO+XzuqZ4MvVTIOkb21SVV/cmuIpBsRzdIL6CN+Jv/hX4BoEAm6w0EHTu4kFMup7+N7U
ihC9WwX3ILPcbbNl8wHEINsC3Zz12ZJcFXEPPBBEHo+Ut2lSWI+iA8V5F8p4LMWEzLRR6OC1coHL
Iq36a3y2aXNDEYDg+xz8wtLHp2Uhki1if4ouIcooIGQZmPaHSaIWoCnsPuE3uen4WilYn48kF5Q4
idyOYovi29GDvm5xhujZDEtC903iVha6IlRMug3+zpJPpfq12jtOrhJPvRFpMRsQQklHp99BG1tH
t9w9rlAvxqua+wQt2IlyZNbFU8qt57cNtJdScAvahHTYABi0DR/JWCcR3NZFNvAE2hK5nNZI93OB
ANEi50C/H3DiK5Fo9gUz7FewTUTjsjzyDgPAI9aHkSwxmMi1pDk5apQfMBFEINeskofnbWbDanaS
F7D+YiEr6rEP3kjwoZsUgFD8N14py9MP5YPs4sRg3YBDdCzJZEGjkSB8Dze9KHgDGNlYT5C9NJ0U
kCuVoz8qCuBSEMA+Wi5sEBptRCky5MlWYjH4vpxOmckuHqWF+cz8G7dnyTn3b3pDShb28RwUvshI
vmyH2XqlKXPdiG4z64nfYbGhzBhQBx1EHw+zX3pxnoy940IB4PXO7nlFxT6u6bBgnoBUdofxiIk6
JYJgTsJaT92oQjuxjSvwWQUhciRL6EqOsn31cquKd2oJw7xEmbfHyFt8V6LAARmPsJMzj5R2h3k1
ehwF7PtSSdgBszkmoVz/N9TyfCXfouEsZqkjT6XaCI99fuXUMP5aAL3g9q42fHzid5dCy70p+k97
Npd6VJjrWHI0eQYF7YWMGFil1bW9ND0N1WVCQZkChewq7P0lDUzOzODd4BJp9e36fpJ2HYSO4axe
JQZl0BQXcF+6cqbPdydfIPA+yuwyC1CyNnt4/AYXdVGiLlZeunfxFxDmAcuGYIdJeG2FpAZ2Fd84
OMltxo86pVWzSB0I22x/92mhzJs8PJcFlvn4QMnuan8o+Rjm25Q0+BRXmslB8mOCgdaKW3jUyF7Q
Y8LZx1Ad7XLyQAl1rLsi3NffLLczCsSSQ/bA5ThIWvB3hv951wbb53cnvHRt8sCxWc/RO3Z4apIr
jALVwzDqXA2pOn5y1TTfG3JI8MJI1pv1vNQl4yVpT6WF3BoVg25rhyTem75JOeoUs9x3zhjq013x
yymrKY4H3zKPZL43cSVDEAny5ndgIGUGbye8Yyi7JglFLodNAHHxhanCgJ8fNK546/j4ZjaZ/4Co
SPQBCf1AYVdSEEUc6a4PBNoAhN7COsBEM9l+d+ewP245wW4Av1PBwB516+mf9PqVsnTOTLzf5LeG
gom9eVpk1rbDHRcO/js3WKY5VKlhDsvwn3ppmwDciVJZhWXkqRxsBvdWgX7aO2oQ0gxGdavNAFIK
NjrI2vdZ6wv35QSAslRcZOjh+9QtCMoRq2A29PCaBI96RFTx+UEJQ2iVYikDlZ9OCUtRfXxx6FF7
8qN5diWXOFhri+lqGFJG3cS36aZwSiUyasR1S8W1jOUqa5+DoxqjLm8ht+9ke/0xjxY0peF8MeXF
6XsihYBMzrAr4bEUdsQGfM+fveqYh8wJ/m62amEpHG5WBz180viFUYDxxM5FxN6AASvdn6R/aIi0
1BWm6vHG07OCwUwqmr+nIxbBLZ82l2DHRQDf0aIVysQDApkGUe6qgaRVqF/WdRAwJoZlnbKnMovu
UZvK8Ab70VCro3++MfFw1EdjVLv3qJWtHSzH3dxTG/FM9T9Ota3dEIa0GF0cmXtmrLefKn4S54OU
ibne7+lNoCKpqQB5Q6fsMtSnmqpwgPmuBMrH5SgdlRFKJjtnr2mgRkzN+vAmvEKvNV2rPZNlhk3U
w5EOv231a0V/ZgNUr9krIjGX7PM8hHK1IqHKuSvIzINNuZRXgaeHNMsAF5uCYjzS6nZSv0cVrbgi
hkJTqc50u00FnUdRQ1EB+WU4ksT3n9moOtZaZBpI9gXlIM1zZUfgnY2Ym+ixeKKCppBBoGwK4Q8o
SgNd79KTe+7pVjOa3GXIULWMTLf4sCUnmfVcxAewvlgb6G6/5p4XzU8PEpATLUc6QN7gG0fDil0c
7/1PYJ3QA9EksRmkxLUDJLtfyBgUnDflWEImrMaxBzahNth5h4KhZaZxryFxhbmzSharzKG3yUYe
hKgmULYylg2mVVyktghzJUoBNnQ/N1RwOD5pVZ4YuZo8JOsLml8SBq/FoDJLOdlzKjlPd/EBb4Sc
ZitWzr/tL+b7SoPiq525b0jVWoAUpZIdcsj16iWn1n4u3kOKKX5QWJYF/1FmbOsmcgdvCW0DQIIf
ySp7O7+HxJHpuux6fY3V4RP1yzca9h3aueq2GjcgSOcPMpsbxqvK1X6O4uc++CRkbcAJ6mfDqpuG
DzO5QjbePWJAJlB60pDO5/acghhEEI/PniZ+5SNJdKGe4++mjngpa5AiuaitP0jfgDjGEYXDvUNj
3gS+Q2gkSgWblR/6piBS1pruZmzMfrar1Id0a1xW8QsQU76pT2noGmaboqTtC9CBgrqoTX5y+U3a
EfENgfYq5IOVZV2lRAqXWkLbMobYpZEHygz49/v98W2b05Orqator1Bc2t2Zas0KXXxSt2rFKS4Z
awminuJFDZN1VJlkHL0yhvCz+8P82LPrXGI48sqZqJL4W6K+3VUCjU5/cLd7oRnE88/6V+UOQwOv
DkOD/sMgXD5HxnZzd6th+LIsGchPro5eRbb9iYMf4RVfs1gPXE1muq8F4lqxkdSVVDidBHTgf0F9
OKrAO6UxwPPJkfPMLm4qQM8AmmDgJWEq7DU+exLSq3ObOcDU/nkuIEPfJcQde5sZ4Ddp+R9KHhKt
1Vc0ldIhe2o8Er6gUkxHa73wfiFaf+ra1W3dq8yoFegjtNQzzPigOgIZfKgCIvd9kGeyVpY4riIZ
53eestFyQTtzw8HD5H/A3A+L1LxCWJ0Po0NuAXurqrDk/8l+yU/q9XLzl+C88vavZyxqtrNI1E9W
1mZMrXdKCaPqvf0wFcb1fhUsV8kNxsoLqK06h3sISPk42G9ZW05YGscHHInYNfrBCGkE8CV+nTKo
sXbO2gBAZLVxHK+C6V1c3WZlHTyk+iyjqk5oJe1K4XgA047vkbJNgCvSXqJqiKQzULNT1wcBFbdr
3j0N2LFfXLVPe+03SI4K5j77p2cmvRvHtxmzxCLblZqK1X/TpSDyw29UcfcPcKRIxvrkk9WyK8Cj
6BMLQrjpBpolg31vdSDE+Ka9fDmmKny5aO9sMVnX0PVysDpe9g7okUbYBS08WvmMQ7NtMGEfc+GF
4NBt7YHlDWe3Dz+IxHU+X03HhWcW2c7taIzziN3Q7n8iUJcbFGlxMijKqPeebxbxV73dsFuRYob0
bJOOs1jDg3ZtD/+S55UsCVONGitkSjd8jfw9aM7aq0wZDPzpSh6ybTEL5b4++8C1s7rAjP+KyNCq
oXS1ooEGQZr+LyvMP4IkX89eT/n1XW8pyerryXsZXIgkWmN/zQIDPz2SB9YjPW4ktj4G7gUer/Db
aywXxiJxLuUHAMb45PcTlby08UuYBkrMKyEYCQqxqfipQEzh7DHE9jzZmfQhIaSGuB+r4K9VtkFC
H8qprn2vA7A1TuR45uMqZZkqwHOkWnmGI2uJewbr1thdrYZB4ZiS6d/nqa68Vtz3KGWABU2ePlSW
N82BfPiTwuL8VfGPgLV1w7Y+qWpAF/RXixDqaujdBxBdt1FCBMJghEa1iu3KiJqPi3gpDzCFIuR3
IYvl9dOm7p7qGQLEWkKOFdyg8Lxbte07FXNFl7b3zAQHiedRbwlWKxxyZBQdU0GkZI2dYOnW+Ibr
YaROR/+b1irP3QMYoyeFhg+PEH2UQ3QajxVI7koWq7JzfHH3IUficJy4Yg2CWcTMM1Qngrca6SBR
RXBQp8KEUq+Nzzb+1Yl5Xc5bhrEOQLAvI0dwarnwtxE2GOTspoZyyJ6tpkA2c9WdDOdMvNCcTzTF
zoLtjU+cRBGNb3TK4fwXVFtMG2vidKVBrGxljWZhVKQcWbiX7UG6+F784ZydKhOJxhcUGXwbcSkk
Sukvf98bNHoEaB0OOzDaFy2/DpqetiWn3R4f0FAYCoY9gqpUpkIKAoqVhel2idkcTz8G1Le2n6fz
BfpFUszgMAENPZ4kn1xj27Kgk6mKuN1+mLk5esJumjDbW9gztDsTC9tghcd2I6Ad2vmQNlW0Ritb
HIwe43plTDpHCrZ/92qgNzZ0wsN85cG+iqCm91LN9h2Hd8kEItLHxas/8DNa5sdX2AXpzkBEDOAw
lshbYMGLthGXvfzBr0vonyqYLTI2lqyWXh8UOkf06rZCl67HBmlTZR3RFfvpUHyw0dgxyJWCei99
FQFjapDvwRsjxYFrEkKYJ4j7NYNxsnVHScprv8VMRYwSWVzpiUCt9UeAFFtvhhgLyAhEnEVw9lxR
yr/iZ2AOKDSkBwV6YOReal2a0n1z9QPPbuAUbheKycoolWDt8XcKAl88bq4lCD7/MwCmQKvBpdzf
XMU+49ISF0hKi8vYejjNEP6xQ8DAv/EnRcMrMb2Bagm+KmibO+rQYNjbnl8VkgqF/8QHkACpT927
a8dfAk4qCfoXZgb3HiEtXYgYxkkU9lGGBqJz+r5KzzYr/gDiOsQRymHK2rNLz2+ajkIWHnY+PbjQ
GIl9gqP+tuMsmj4klnUGE14D68Z09ImKC4qezalbI9CRJRTiD0Eb9pG8OkZlFt62E9J6b7CapZTb
RZbnoyXffNpCCN0qmfO2cNRICKqrF/IcPm2K+IOn3tPwfjhySCDdYtNTRe2wTYXZA10fP/FyJqBM
0Kiq705mFX17dPG4m+8YFsq88oZ82e+Vjjt1xRuzvU/fmfehKoLtB38aDJ73VLaTrv4YRBTh6vss
tIXGWP3eNhlCHg38L43A5ZvMCA02SzSbc8mTUEcdDKawBbQ0HDoIqv7KEKXFlqo9p4Yrvu9ZkqqX
jQKIa4vkqoVPkruXItvJghDPJhOM5f7v31OB14jZLBbFHJKg2GtGFxh7mtl1MWau8g09zGDbZhci
h6bGcbaIsBKT9x3zo9oqNgGjWR+Wa9ScDkWn7QVTg0Cot4Dz2Rg8YVE8IHONB9M4NPjY0Ce89mJ1
BDIzim20FnnoLfmH+yeTyNqkQRG0TpjZ8Mc6O2N4QUOxInoo9FB7yWN29R0YYik5lijQNyvP8bUz
3+jL8YEzD1h7MhAlsTB4njImdsx+jExk0PPVakXMu+E5lfvh3UeMMKQn2ZKsXdM9OSH8QKWjqPwp
YwQPO6I3agK9GZ0IxTgDn+RdQtS1OPjUtL4WkVbziyV2MJH42qAnnOA+VnoJFdK83j48TIENpGtt
mVNDWE0Ry1qZ5mp1OvkmCgM4kYwcgRT5RHp8M/q4mCWC/EnlUq+GXhysXY4di6BlUPtYkvFTupGI
TT4uHyOdniXzRHQ3RCzBsbvKjI0jGS+l+1oOv8wQcdlzc8BJ7CYvF1Rfb4ztczC4TDRAx+43p8En
oeosPrTW2ZLhaywbprBN1MbHv1qKfhDyDdWvWMvdraraT6q5YcZe1/nwTa9MlAXsoD+UZGXNAhSd
fJawEhpGnJWhH77ayA/W39rDGaiN+TZEdUJan/KtBhmwO7b2YjlFroUUs/7EhAmdRe1aWHp+Gt26
eS5C80zKOKCBkcR5aX8OoVwEzCO1BUy0UWdjIKVzQPqu57FFmUlX7Hv3HvI8efv9qN0qmox22lo/
nsneGoadoDkoRKOWsSN0ISa8H521KD9BkOVc6tV81+4V6pZfYc/2rCPOw5wi0T40JqUZga5LmfLE
5IaFI4Jl1Ro6rKKbhzupGwmOD47Zb+/i2fefe6t8HyKHokEZoysEKkhjIvpsuvM3EeAglE5iK49E
snnV5rC58XPkIKVF0LNF+wLqJJvmdKpYp06uZFJfh1dyiNGV5StKd/Aeaptc2mkpFbKT4x6NYlO0
Vs3u+kyqsCWdiKtKxGTXy1oddCh9T6Z0RKiew+dPi5KzN3JBFa08IWicHjRAgA7OaRHV7oJQibmZ
5EFFr4aXtwKWOEmKXOeazkKbh1Wq/TaBqy1YoSIyktYFH560NpgpxP9xn0d4Qv0cngc+GmaWf6DW
/SY3XhnLpnooyQr3lwF0ozibzryFtzTGi1xR0FB74lh4ba1gJLfqkev3BcyPEb+SVxzVBASJSQZI
S+zWFgCmZHrlInioo9z3IlPcU5J+g15EZ0kRO4hkblW+x57u9jYX21evrnM8Y/ov31BfJYyHeL0X
CTqOguGTMQR9/yVl7Okh/8PSduCKXf+vvX0NCQJuvCafFw5SAI/iTywIF/R/oEo0iam2z8lPQCXw
GpdGXphh4ukA3bQ9wL/mIR7nniIRUBUVEOAAjvMGnyg+DV5hhqRzWg/JvJooYJlzIXVVokOeZ3kp
LP00ZMLtRvZqT6ZP3Qt8ngRwnjF6prrZziZagv/1btqxr8xyxcn/A1GAkRs8M/NQ4OWU1S4+ne8+
mJUqdVm6jJUYTC0lwrBgnSHUYL/BnEmQK5DugQlRPQcA8TXHJ6rwKq132pUIDbnIvOwfFgyYRvR6
5TmIK0HRJZDgnohRP8LD36EsSZTpIWKasuKnmz7R76HizzoL5GxefwkgHUsXKzMNNl9zjBkX0xIs
j/8XwL4//Le9FL7PuQoWqhOYxqtQcMuoA54Bgf2bqFCiZL/MgQZwRegcXhlsNR1Zw34a0w+SVdoU
+Hv7lLmdG4R7tsQ6iejhtC+jateECH8bP8lE804nfUEtTlTZqeRpVh6XXQ7X4/F0DT8ixMk+Q+h9
i/j7TJ+lHp+kLvY7QI/Zb0ry89SeD0fVV7qLo82rTrRB+z5padq3J35vxvgy5YDP7d8ol58vwy3V
aF3TXm+EOzdSuqa+e/byuttlA8e8y4ectfCsxAdByXIQHl9ZNgj4p03zwNtdcspwGOuZwSL2JjKm
Lya7kYFmCudZxrs9GqTQRXTsGBNqbuixtvhMsMGIGZBBwiGJPbJ+3vwt/O2d7k1iGgZ9ntUbEO5r
Uji9/Tre6l2yCjpGi3JrYf5G3hUwrfo6w59VERE1xwtKxm/ixb87WL4cPUQZCBKLCXug0LpnqvH+
W+GQEGH1dWZ3RNSrs7qrT38slmH6LqBaTxTWxJecnokYWApwATiCzcpKfziL7KDY1M0Wy6j2h6lW
xI2KiFn9QwddhyEbvxu0wGC2CohLzfS1/NgZ5TTLTodzFhqisK3VKxMzdJHDgbgsOboE6XjL8+jM
1eL5qpHfOzBx74j5+whg0TrYLfxa88nymkHYXM5hZtqbya1UQO+s0BKGxm2uUlM7bu5naxGCNRyA
KWqKRKGt3EIaQotHKwa3vV7vjDCoEIklsBxhBEyNmv40h+s1AZEd3d91n9IMZ6X3YqFqeakwlaPu
ZMi+OvKDXoimkcx/h6DGH1CcEptqJGux9lmHJUTxec4cvUrAEoOGEhJruKnSMkxuP26qBvYMAgFD
Ax7NNfuHmEhyquqDE063l7ZgdISTY9/CFpWlwSqWanjGiDPns9A1tL7Q49U1xfgDWCQ4oODUm9qo
kGMuNFK4yj9aqSd4bK2T6aZD02VoAF+uKbhuusk280/Ngki72liCBAe5K8UZs1Syx6y8YXOt2UXH
Cb+Hxtwi1pLyly3vDUea3Jd9lKd8wNQlQlmZQnireWG1LWTk7/eusAMpvK12p2D8M0V0VczaaBfu
oPjJVO83S8BcuNa8YcpoItZc1wHNsVtdXVMNuUSxk8vtg1avE+r3MQGN7//B4Zwvzgmk3erf1CM7
fjeHTpzMPNhp8iKXIpmPUJp02b2u7HL53TMioFIUNesX44GfhB/YOfsiwhns02K3FFIkS91ckuoX
8r/TTdIg5EvLzC5AR228/1rHHbk+uXc8/vQI+6LxQjcjEybDWboNFf3EvmpuF5pZWDRvis6Bx0IZ
mkDsASj2RjlH33KprjtjT+wHKUb/tlbhQFuwYIn8ujdM8KJVK0gjKM9h3a/sm+1J1cEeEtgbphI9
TJ/OgT9tnqN6yKngncxLDhPHTAN/5rTtRt84WNc3xA/L9b0HwDY3UhE90QDv4AlZw8zUCuOTYZ8A
JeJdaFEG5vpSugRiUO8DtZ+c0/sWoTi+8KchDvQeV3G6GGjtwdGS4ne/lN9gRodH4Zt9ItexV+iM
Sj+iqITKR2UWpXlN2WQflowZDdEchJBVdSiXe4WPCPq7b93NSF/Sp8LVsTwBh8PQLqOBU7rW30j5
oyM7t4mticD8A1FcB7E+Xgnl6WVRBq7q6U52G9qNv93j6v1DhQpRncIWv5CocQIAPhTcFZ1wesuT
4pczmgtyVfnTGxk5t7eAm8EyiRUT3Xs8PKsD7Tm2n8rfXoD3d+eCuisODbyMaB+Qw2fVRSWGDlf3
5K3WZjaqUBiBYeuKqpYC5JUb0olKITWs1SW/zCJ0/1u70mRane/Prs/t7R1N+aD/9bA18e+Y5RCF
+/w5HzMGLPXA+lLYdECKXmAWkBRLnNaV0fj0YA9bzyJTN8M6X+3vc3pcNlFHPkojAHE4x41+StfX
Bx7XHkpvqIUU95T/WbfcL+OZF625+F16SoTvKg3tWv65bTy/Kfcn/CRI78DIDahlLKWQnEzMwr48
9b1+qlfyn1HH2g7iDSAOK0Y414/rH5z4NDO6KfmM5NZBEvCR9ntYVQ5pz3fxsCV0KoNFax42vuAT
2gkrrGkRABqyODIOy/a+StZ++8I8d0wTeA/Vsn57rL89BEf7cgewxS+vb04hkvu0hK7yN7ijIXYz
5+rBWUDIIJZez0V569LX+vugCd7Afw1M5PSm0efVAjVvzKabtbIOiVudcd6MxcSQYTuPHYTViLrN
cjPrc9cHn9tCcW0RMxVC94iO157E7NWngKvD5ATv3V/OMaFrPH2byvJPGAbIhXRN/GuO2yeCBEQM
fzqNGsutllrL2NOM6/Z7iclk2ikgmTd8HV7Jh/c5UOOsuocENCpiBuODoUkSawufTKjYomobA7Zx
gsHGpNtUw5DYMXh9WBqLhO6GW/fXlncKY2FjR8E3HgcS3lMUgRiNL69LYTzykPl9iLckMGLrZ5XC
vl7VADBQ5BWQ9agaA9Kb06I/J+mu4AbuP1Rzo0j3x4WtZ8is9zOcRzYjTsfs9NJQ16Ugq1LN6p7P
K6mUM3pEkI9AkC21AaoHJ63LxlDMjigxfeJJvzSgL/9B4YrtypjbsTJ9gI1UtKA2+dKSTjjzkCke
AwmyuhuGa+TTfdwlmVo+vD4tPWa0+GeA62eIp+h4T/1JQX8u7ryhIwQ7Ymrl7hy/WUv5tBw1pDQE
U2jSEZ7axf0xGb6o44dsKop5qsWljB76lkM4A2YvDNmOkOO1T1r5q2hhtc0BZlp3v7FnMb6h2xFW
JWURGvh1ZlQ1aEEpzHJx0YXrxM8sqozgzqZtZyVeQSdVnIPX6XzKUf2/TFLnqcetgYBqWWaHxgra
q3AZeyTGT567yMSM4UTi17RQwnVZUlfdzaw65qHCyBQyIojIpkhg+rp4wPO7xZs73YgKbbBzaFN9
fdBZkyacsJwOWNkGAbvqr2cKAu3qgpD5Waf1XpqUPZVnMU64nQt06Hy6/WwjkyJtNj7VYm7p3yfI
Fbz1HJfQoVL3xCSYJNjjtnqOzi21l7d4TXoZZD4cMbAEBSQemCNoWUcLNgGKmJ/elix63GZYpcNd
hWbxgDh0Oc99DclYeq4DIMqgZ+5JYbcTvrbDXzRHzLy4EoDBhMF4wjShzUckkvijSewrNB2BSgX2
FLjMIaUMC5s0I35ocy6tlSiH4yvRS9wp5Legu+QbwG8UpSTvutIGcFdGlXceHrj0o9sTCrr+fvLJ
Gegk3cBl6msw9zMfrJRs+POx3mh8WFGlp1oAxmMpLWc4RYz33bJs6c0i6gGwzY54P6mRZPGgog8r
K0SaigzdhhCXs3L+HBxzzKHolqVojhG0c72V0OXIbhZkp6btXhG7nT7zb45vfDTP6l3Cxv8hS0ct
YA/7YVezWMdm4+48UQMRgDGwJii5iadfyV9Y+st0yL644AoRb7nTot505wZ6cCYoQ1geNkzAWcy6
C4mVbDe+qkaXrHbS695uGQ4xdFe1uEXEXnO1pKxMHTMnupKl7G+lvIPI81MewtL6AUbGMar6lMH+
hxuM+gandsvI3ypZt1WuGcGfNyBiXU2hrfXIAhuaFQE8iQRYJaQ5NGFyYCSj8vPjarYTPP0lIPR1
2QqHN6SmpxjLNShFbcY0GvNxPWPlwdrl1UA4ut6flgGJIaWIJRnQAJK9N8QGuikdfdbkCOcgvn6R
BwECAkq534NuSbquSIXEfYsy6FHpV5/cB8/UtaWwYD+wCOHyUQ48EVwPsxY8RnzUSl3jalWhtcYf
EYGmF52Bxqllkc0+eiYeJoRP/JayW62hhmqaEbrXYF5jbPbykKHbwzRjd3seNgYSwrX0V71l72wL
kVizAQgjzW/1Ce3V6X2BmwJcG2GCZC3Hxson/fH277hQU+JfGuNk4iKilVtq4AP1xwPSFIy3PRjI
3y09slLgWw/Zo08ljDxU3Ghvzf7eONGbn09boIzXiBuswmDe3WGf/cjpaVaeehq9Mi4hNq7lYYjc
Ed6614idIfVt4u/5iBdwvTBk+5Qx1+PpKHVv/V5hSLuEEmhdwMMbQ6ZXbYgEJ9LGCL9usVxDu+EB
jXsBJIL+znu5k5CD9ZGben8pklrpG3EtJ7h6bBZxlPHhvz9/PjCjvmnA7uxuYLp7OVjAP6xsXOMT
RWkVdL0FUHaxgQtG8hFX26oCAV1yclbjcUAfzNGFlVKEDQeH38xiemw+tUxw6z8QB3fW42Ho1AvG
Nwczsd6ZqOmk/wjz7L8psbJ+YFCDEgxXHqP5I1qhcMkaGTw0orNWdqT52hIvatKhzzB6znwxCA2w
tFBNLs/dVGB+u88VCXsW9sLj1Lp6RpRK0p7bfn/pPX3zrlduR2/9D9YNh9hVb44cyyxSIvqhuxbB
ilSTL7buaXTwjYc5WvDpuC2TDu6jL6jglCZgWnFHrEjzI+jRaaN5OEzEypOUh8i4lp/fx6jWd+W1
7qC3swLdMA8Nd+n+pknBYDNONptvz859cHs4mlDw3BPbF6GBbOSueY5L1nb9YXd7vGW4fYBEbuUw
ZFOokzdrXLsVVW5Upr2sfUtrPqsEM0ti/rhO5EA3YeQy78wrDPJYKLO3r2+5hzv6ZpHcm6gQ7WNr
gvuDEm59QSdqMoc7IJ1mbR+huQazvG4NJr6CMwsg4WBf+EMF78vai6ipEfxiYZwCOJ4bHFtSFWd8
hcO/+zLnX3c3H/OiTa1mxhJZZmZEvQURgYWQzrlJgyiLsmlIeLtzGrwfhfo4CHcpm9THlVZBjWg8
F0gMS69eP3sZVqmBp/tmB7eIvhQp62VZLENG0rIkvoeb5dzK/ZL4EUm35MWY2J3iG6JrS85PzuGL
q0kLSbjx5JlBFLG2k+3CJ9LherYrMCbfNy/e0Sv9z6keeiukVGNBDYiZOxvcFwHwV4viIlvLfcbB
L0M2BMdgYqtIZ4k7oVaeFwv5/K5R1/Z5qMPEJwPC39bVYdzamerSo6gqPi0uvjxVpaksZMRlTddR
Y0UL4ZGWuUIbdzlke5GkJMIj5UmhaERJg74JjNorj7NkjzOFrkEo8lCE+rsWnKGrCY98O+w84EwI
bHK0C9VcAEdkyRZInTmqaw2IA3R3j7g52MRfkrDG+l9gK5JLuqP8Hr08xnTjGTwK7FXoqGk583q8
FQA+apfeeiAUSQ+f3MSpKBNTAa4W0wejr8X1Hw3RHG4m2rZm+0AbpRpw7jydXe/qZjfSbwlUGJvj
tnhZM2L4Tld3Gl266HB+vK9VP4XKSGrD3q/6y5mZ7HOlkb/DGtKw5HWqpXhkXpClUheA+c4L6suM
EZyhs9LAvB2DQO4uPZXihoEyp/BgieXGLo5cjv2XcfT3al5TzC7udjA1OOR5Lizux76sm78CxVAE
Zwwk+LzRBTPcxhARZEmFb+78jrgnxer6m4cgtlm7/s+cSJpCkDh6t4cMlNdPbo46No2kDHWx3EpJ
lG7qlQ6ecpsJOUxqs7B+EUU3ZL1gI0RbX4TS4JPy4THTVD7fS4pB+1rm/7wzawoLdyZAi9DPd+h4
FydqeaOFC/8Ukzpy7gMokWrvNl28SNGYdcK08lSKwWeWLH6wFPqRwH3c25ExEN7kAVHM1UxxqKJK
JD5tmCZkYyixG4LjKAXBf48EpBbQYqBB50YF0GnafTPJzaUeYjp6RKHvtZyRYL6VKamCDLZXMyC4
QUkV8JLMRHtQrY+9IawhWjpNE80bTtoHK8xa7IkIEejE4SzWueB4p9t0cEbZc8VNiH0HmTxRYIgQ
LCfXcf/fDAHbTvr0LHos0liTx24xBLKwWmDIcY+2YHOOMZ2hXn+jL+KY4Ri+98mN3q25rRd+vZIl
ujGCHiG4ZLwp1WrvpASy1zinIHQNIilhVXCFxbd5RpHr2YJFOxGjysL1IlNMsqawELYTzFpNyH+8
ibUrk/ykm6DCpFMUyo9HnPvJTHDohZxGRIVBc8VzUXtDiOEUCCjIl1wVAMDisbqXdzG5yU623Dkj
ftgksp3QFX1/UetD5EQ5byGcIyxcOR+2O2LqIzGufZpb+wVL+5Vnf4Ch/AjWbiNZaTpE91xJUwsJ
Y/j/7eGdF8JSw9Wfsa5GLBs2yrCTJxkjx1hOjyZvHrqaGUCZ0hJCY7In6LrQsAaCwjYHE56yZ29L
en7QWCDCBrwGzMavRlSO/lYTb0bVZQEake7A4Hrdn42tIVx8NVnyhUOn81tsMpu9rJhxp+PEyK9z
Z/5NU5Px50LLM/RgI4dmt/gQ72xpArl1YLho6dXefjm2KcSum7uP5XjShruB3tEjyDXpJ3wSbkEs
uXqPOwRLajaIc+Q1ii15SY+r803mp/chs+egwL/meNGiJvBo9YP8QcfcGF/7kTPzW6hZoDojxOnN
F38gITCMPjWYXZWHmgXIwgwLPfLecHN8HHjIU6ke0uxsNrIq/Odz4U8mq4cVemYt/YzzyBprFbq7
YQeg6wVJIVcUVDqICxi4uJtbPHUXyN2wTArBYBIvdNXhGjPv6kp7NMQiVXcsQUSKc45heIrqVNOQ
nLnbXyRM03hLdtrXxQaJctlXflcg/kgu8CbR0TQrH3euIKDxSA6HSIrK7H9C53qHKkVOfvdy09ah
Ar9IuaD01iU0drJVZKEl48xBHwJD/bE4TmrYr+fY/ISm8O+fQ/svsxXkUF5815/8ozSTjOSNLwtM
csBHhNt6BvgOOhkP4F4M7jSwam6NbjJ4+LmDHYD88ETmeSdx6wqWfVTz0IUVy3W6wurAKqyLPm5y
iEerEspUZLVxhoLGBTG81HiqhyeMj/ISbGzDKC9gRlqpwJwTq3MxSMIKiqNBuJbgKg7zI790ydoJ
/iCYwj2AtS8uIt/CElRdZ0qxeFW/yvCVUjsmGqbBARGgg2fF5wVAzdZNfRpiBepLjQj/cPEzsrES
0uwjciZADLgkqkIz8VlqyH8l4+C8mUKcCrCEB/wIh/Aw/QVKDN1qwJP0xGhdOgcpOckNUSoMrQI6
qcR3UPEHQ6iy3L9W+j87b6qlqNeYiPDZvEcmFzFuH4w9UA/KnYhUHAHLn7FZ/SSBhZSSK5K5IAV3
jA0R6kSFfZgZl53QEL5N2dbioqTWIWM/aRhqYzqwNm4C8y+/+IJQwudThgLF0UZDm12Ff1nBaezE
Pp06unK/cGpV8yIVmAoyvH3bRSAJMsUpPpiBs/pT1EKr6EuWMhyPT/+MaiSQJyDJVBWmhZnDdKMZ
rMCO7V2SRu+gQU8Pwprpnzguk6/0XOSU5SE/y+j90seEldK/f38MX6/caTNNS/Ju3t7ZgpDFqQ8F
l62OOPSTGw/ZBnfYe0R7EQlMRhEK/nELW9uPUb9DCx7WLzFpEk9vT8+s9EzEHRyrCKmvG1aTbPv/
5/HakgCI4qtYRBvuIZh0EQ/wPfn0yxT9unVRWX437oZUxGMvedjfNYb2JB62JMhK2SPQDNEyVqig
F/oJxWOAMJOoa9U5lzHq37DSmtnIbtneXD9nqKoHOWh4RMHLMFZdprzOwJDHCRk8Jq4T6GgDjXB1
7xmrZYPbInaKg1xg6anlQTyqJUFm47JKT5h30MHdMtu3TuDqJYVV/ulLcY86kzpQ6YHHVrZUlngu
VGG1+Iw/LzlLwI/dnnMQNUZ9yp69dFiI/gFKqv5DosaXCDPItKkUM5hVsoTa0vozQIyxs7nJNs94
h1YhPHZpT5mSsEyoLc5HigeXiLWghwza/9lHgDM6oEcgemIcBNSKmY6C970DpTy/Td5lmPlVlZTb
De2+E0VHYXicN2GJpLM+prUt7Z6NcK1zNBpN97mrglHHTdYQ143vqNU8KaUrGXkAJvk2zElHd0R6
yjmeKHF8RFNdyI3NP7kQ/mRE8I9pX7/X8zhoBpSx23ZaOjQaeus2u45M3a6K0I8D0tYwXXjbE5ds
kcmQXTkvmW8AAmhZgiRnT/KwcwuVQRRHJ++XpEgMNrIdG4VjfGyQRC5DBXw8pj1IrCbT6Q/dHJ0R
t66u5SF9gaEGOQmwIMwHAv9SP5JNxzuncob6MM/GtAPuxCiPVHWF6ZQzBz1GdltjrU6EzoygRukk
sVbuDiasteDOozpboSXk5OptO8D4lOfRMaYLErDt8cYQf5XXHVCHldzQFTpdbARdZptt7Nbi9ehT
wP1d1rtDurYcY42J3ezUSo+y7Ogo8hNi5/NTdykk+DMTtS0qTxfKwMUWN0KrNTOfF7MNLYLp4AyB
5LWNmIupeyAJ/VL/FnlrrpupZhHxvQ24mYbNyBL4nW1AnJ4LzytA2e4KC1zmvNzic3hr5quHYux2
2RkmHD4w+r31i/4G1+xqgbbvpGw1jpORA6PfNPvtKCVwJj2EE29pJTlfoYVyqo+QwbU5mpidYfPa
WPpQ8qPB3dkAQnKcCJtnABfm3A079dN+EqmglS02qanyAY+YeBtA3bcXc3zNR7ssBI46g1577VPc
EXn9wxSWIZHE/rHKFuRzIslBxFL4hfZUj2GKFKKDWqRX72U0tYgVDEcNPMyAAmcEAvId5dCmmT/A
cJJC1V0xaddHSBklhasv8Uc9czkcaS+tPDZBP7VRXbhY6rmS2OEGdQVQpxSJXEHwEiLy3KJqfOgx
9H+PgT6xyDLblC1YhYkFG0ht2cKyMXaOKqikH0wDQIFwedAZoZUSzFdr+Qri7HFH4w+M7AOFjywf
ITYSvM9lf89qk1gB+Pg/J9COBHjjqtp25+EUsWzhyEJhPvztvU/+VXiJyptCKwb9V1DEnFrbstKT
LxuQLCSdRZSj8jKzwlBlFsFKYO1uovqVvWALWY0v9kVg9EdVfgS20qbqmW0DZtXsiNwLkh6DLV0V
hdHGW8M7CtNYUpuFOTHd3WFlC+ltu8JpgT0i8OGll/F2mprR7tWPe6NpPbZG7pQllcyeMP6g4C92
GeRUf/vUC+KHfCof5W8YZgMZeZRgY+E+vOl7nPnoM+1wtosfspahXf3r3QTidKjSGlnMfGTo7+IO
qtQPtjoLacG6n96q2yf3j4JYdqX94TgAtpckJ3MvzxuzqKrNTrLsSsNmdv08ZSTsICFXs3PebZr4
mYVG/zmpfX+Jv9SA+yb0fYrX10Lqu4sEdFRZc3Sphl1fXAQUvBwpX+afZ5wkKJeJ9Dkio3ZZyV/w
iuZdRuEWmyLT7BxVsWsYQ9RGakmowxHguT060XF1QZ5tehJKgqrDwYZTR8kLI+OhxRs1XXfTEbUq
ERiCtGfMbBLsZo5TM9l71Sl4ywc18WFxl9nfeqPlvlFPvmUUyg4jlDPzKCR35tKtRtPI9z9BSAvh
57Q/vWpXCMgvKCMiV7PV87C4aapuVSjz7xzYuItpKR7+1xAq024sO8M10S4e8g0ECSXSS96cEhtU
NXzap8Tnym8iIM2m76ujLJIfnDF1cO1mOZZRhGd1/De+0iIWx4naSdFJhdK5Je+GyY0OjGyx3+QI
y1V1jtdc8n2bZIpvgqS9M0Nlcxvn/Tk6gSiOOR9h7K6btWS3grBdfPLmFeTx72CTPNWI2jsQ+TuH
SyGzfnnVxSuQfmIUxkiy4I6c0BZ7i09RVi6rZyr7/Iktfm/Xv7tq4w+xAUFQ36bCF50cqZ72w4QE
143fbePKz1nE3BSeAEc6AOWXMt2zsoh6O3+d5hr8Camv1OvMJEnhHlPeGUMVgGKlrpTzTSY8S6x/
7HbRZaul4vKHEx/2pugSXjtdLeCMwpfjpNk7NcqbGb1dyXiqaCZsZcO5xOGy/dWej4RP2f8sJwmX
w5zInTAiGBcsOu4GPyad0laWdpRa5sqvHcEALrwkyb9B7JLyScd8pPzlqfeTuuS0PRd2GwJXfvHn
K80g14jcJ8DwToL9WX0fmTJhnErGggE7c1t41QgkMHQULYUauZScQCM2VwpkXe56EH+RJ4VGU+Ij
7EpwF2z1agBTMfPY8VPqeBhcrrQBUzrS/jFaPaJ+CyvuRPwmyHbAIcYtCVtseQcwU6TsycjWwVfV
jPb+tkqZkMtEeFx9xBpZRqhnBaWwYDhlfR2ew9JVdsMHhe5ZHSFEOPnu0HBSlwNF8eutvMjRup/g
isDpOzsnCq4PWRxZpxizKiyM82/E7kcOK7Fi/8gQxwfqPyPzH+32JqZ996R2Y1/O0KS/FKmMtne7
sKEHNkSy8ur4AaElp6EfFKFBGOUF5ZgnEuMIX5/AhZDB33oxNU5SPzay5W5p6JZkOOOglXa3RHOo
fQzv8kQY61kebjlWdmitZHU9g/bERs4g8YFd1ID6u47Zmnod487lGGpV+iTX9HubgrSQzkGpo/kN
cbpCenYlTSToSQ8f43Qu82DcHa6oM5yH8WcWVQ18J2ts6jMgn1seBdqFnGalRpC/gMXlAXQEfIgO
aljfWx3tdFVdePDmxrWpZs/JVMDoLOjWsz1QhAubGpHSl4tyD/IH/7jxErZ0qt8WOGQGf7SwAaFs
02T/oF9xY+jpC0shSzLIuyh75Q98YF5D8pNTOx8JOcL/4GO3NPQgKnhpmPzuDMMRjvsZ1LsjZOny
mBkvUIde5DdolupzACB/YhIQDTH/wifTZFB6z4hDd8LLtqPfxDQsq5442NGWbec9Yb6yQofo11XI
A1qkZ4qrj82M6iOqCfQE2kdMWQbZ6JivuWMldwbcbzD501uDp+5moA+GSG71Hw6LcTcS+Qxro+9P
jOrpO3rbs0tfqbiWGTm+sU1ZqGbkMRH1WDNwumVUquiMh7Zhp5EUIck03ZEQNxZmAmy1pvQF+i2+
b6Mz2qAGSxEd1rPksdHcwYVXPtv9ocXULU/6DRP0vNv5N8I83GzIdJomaKoLL8EMfNbOBWN8XB2C
7yHLUSzNdA45lrtnPW02BxB1SXVDOCKjBniwRzoKnOeErRY/Mg+973iBXTPePiOFThox28mBIekt
0tsRF2X7+yN8wgqYMOLo1lXOyalNGlxQ8zkL5gfL9mYO+psj5zw/PqV9Z4tiqI2gFwcabxS1RwLG
OIc0/U3DIy4pAYCHpSSBWJ74XxnvrmpskI9lEh0QlqoSkLscUAhP4ln3zOeae0y3j3ZbS13VPSjx
G8s0wVK+snLLY0DRbsg6ABxUiXQ6cTfW4UxMSWR6m9Z6y4RyXnxlvKUgdeXLwNwqX8dSYNbgTYeX
Vu8WxtEm8f8xnhjZibChjooY/HCrvd8eIWHv+nmEfquf8DY8wgOIfy6LfpC8x8Bj/hwxqiyGMIqc
U4xQL7YCQ397uunl85vB4pxw4lB4AIKb7jAZ1K34nh29mqxXyLdoGDxV3HCRcUHMSX0AY7oTwr2h
YlRK8knEo/efUQ6mZS1zh6mt0qFojQ8ipiSoiFz2nIcxObnX2oy+jOWVzwnqOBZSterQ7EkAw5mG
boPaFMRkpf8ww8iFcLpKGG6DjJzJK5oDh4ILu1wWozLvTcX/ZUkAP5Vt74QeTuSnYzSDhWG6ZTcH
LGdvC0rxUCI2JwI2b46C3KJzb6CmsYXKS34l887kfFpI2Wgguuk7QwlJdW2l8dja+ZwwjhMfm8qU
mEpIOc2d1k+LY9XNoA8OZOWTvHVzYWHUcckY2v01bN+Ss47Yc70ZRIGLxzYDffLpT6GRJghNLPGq
nAyCsnErJQ6W10mYLK+w3QYXLBmRtITDdiCJbTgWlVm30obqqImUrnBnVooad2Jl3oX9UqCxsMxn
ZTCpOF226iGfgX6ciojdC3oVS5XsO6g0WYrS65mi6CsZDoD5pbc2EB5VaeaW8pGYezL/rZ63lTSi
2myev7oJG8rNWxOCzlIB8tgHkwGJz8H+aaRkcCOcuaPNoP/yFUJwY6nY3ZNpuud1/taYzPuvR0Hk
xm/AaxTE1EcI9pA2LnwKKRnEOl6qXTfH6G3mqHlZ3hERomQUJT6wh5ZW0jZrQ2wgpMXA2mUWoInS
Vrb4BJXh/SXyiR5zzq0oqutZ/wClMuE/gtHuiWvEQcb7r++sUiggXb4sexKvt7DYYAkQ/pRQXYW/
+lDTk217SYS3WH/sWALNdokbCcztN9QuP/cBKKIGO/4L4jEvw8J8MVeZQsN0Oo06hg+8EjSz9moz
d9YH24YJsfPxKF4R7K+fJXFOE4bLyK6KJA9UkwWWpZ1deOWnW2pVF1XBt9MfVVLEdOONfDzzV9Lo
fcaXiz1Q9eaaUCqhOskBUHU1cdi8+QniAiN8NjS0EIN2thzJ41De3PZ24Jb0U64pWcFm7LuMcs1P
RNhgXxtfnThI1HSdmApyob2LDFQNvaHcvMTtMXuNFHhIuGlT2+wZ7eaD/t5QDhXjMSGImEVg83Uk
0LTsoqm9pf5k/pOHgXRasHt7WTSAVADlIRsjGCEa4OUPSpESk6IQ7IA6hySlqRLdzaUI6UJMkfOK
uvrZCVfb/Q8grDaakvsFgqlHGVTR0Zp/L3L09n8Wp6z+ge8D83DoIbM6+uZ9F/l0kIpSc8W21dEE
AIyQXPAvpEOLIXjWNU5LJIoN0PRaIZADlt2GM7Gu/952vP8VFTMwHTTb//0Stg+hgqFnxC1soSKJ
NIjup+Em531Ot6e0Zd7+OMpaSjVMfzd4mNWLVIrQMu953hDKe4z4LEVtKvQHZuKrPT6cqFqQlLBP
ewkxA9/RCCnVcVSUl5IUIeiMqDYE1ihttQ1IHS6TQzDbvyM0me6Cmypseh6aZe2EZtE0IEz46U0V
UqT5EeqsQ6M+98Il9tV9NiU39a5iabYn8PBkCH4TJ+gJyo7lf426Z512iobJnaubJ8mGMDdE6Yg8
ohAwlyY4sQqLGdBcC8IPyrbZ5QHuFOGfyYdsw5gDhTj22D2epaIn2INi/KHfp28EXfQ9ozEpw5LS
MTeJ0E8iGpo7sETHYxSsV6hzbK6QLqoWfJsKiX6dMNfS5cyh3vbTb/HaeVXWgXjiak3hqMHHgjFJ
EZ18tM7dmC1ObFW9Ge6kZ+NilUYNgXVmFM700BjyGYJHh1PJd10EBJO516NIxjKAzrz+vM7SaAP8
zmB3ywZhxsBuI5ZYXWRRwzfPPPiKNj77ISyTaxlWqCljxTUJ8Igp6MM6TsEEcYKcAJi5gL/oFLzR
vmyNfQY+lSagiu7Ejgsu36dWsFtjABaelP5KE8AgWOl0fbrp2iVehUi2yGAan9okMCYXwK17hsUk
JQgNIILX2R0g+n0neDMw3PumYC9TGNKNR4DdGw9UlTCNO8woMyoa5p7d7esitjEZBvHqThIyIveY
42emvYpNBJMDxAG7TFk5aN1eS4irItrqgJcR60CTOtvoCSTXPI8sIFnhf/LrLeh12mhuRpNAJFrX
xn4I3jmxoK9KUe57b4fpqvSVJdRpcmSElpdJ0O/5Aubacl+kphDz/rbxrLN03tpQ/niAYLl+5hXB
hDmrMqCjeddsPMTaJQXWqTsuzAAZbUR2EjuojkDktJgJaFqS5wfoQUY/qSnsroqtDB2FqHkpmlpB
az4J5RC+JSFdZVgMufO51AWsyYcpWN4Ams3uPipCEbgHYLCI7op4n3/9cyjFvsRRwPS7066eBLd8
pC9+9m6TB2wAo/tWNLI6O4O2P0woILtYcWl6Epilefacru25xPIW8c5u+8ipUlbqOJidoEvPkLZs
dyDOIfue/N4QWzICF5vH/Qw4uX3ilUz0fB7E+pZracXipnyXfBgr63u0jl7Y9P7fI6RnS4OB6M1i
YptcOkqc6whqUUFYgeKlCa4I3eCVmIc9w4aoSDSPeGdGO1rbsDmm8Loe0vJOUNOq9U1mGJZpRU/N
0nunCBOSqs1nHYNoLUxQ0S0pgPrbJCO3M6OPuPLGghJFawSl1wh2eJduxqP5hDIMnR8jG6BUWi0b
IKbITHLm0iK7rCK9D4dNeQP+RU5z2YkKqN4+Hso85FoWr2dj9vmY+Mjbnh8Yy4e8eIcRxgpbpXsE
8TGgOcGR7WdcTzmzW05ly06qzMk6lTR4c9ywZIrxKXyFq3g50arWE5ozq7+LZsuXQROLR9mY7RP+
9hVRZGPy9ykvuWuaRbzl7b3NqzeBEnaYLS/k0BANzij99uyHZq5D1Pb2rhlNMCR96TJLZINOAtBx
TpbYFktx42P+y20EaVEnRAqN3537AGcyp5JeMWZOs795QZTVCJwuKg70lDKCVXnMFsqR/QmnIEyr
4kECIpeIloONXYU2iA6rFkvsi251rP53l8Eu7M30cQcr5bpy+7t5rTMu6rrHEJTGbH4xUBkl5c8j
999SRuB7p5UsX4QeD0GnrerqLPWiBA5oKOTM42QEhjuALdnqnCzxoUP+KZtCSfV7vxvYvzr/XkVw
xy81YHXPoWpsJkqImgE8z6sS+sVPjvmRvGna44DCbsXfPvrnthy77dMzT9aAZ3hVa/K5R6N22Y+J
DmvmRl6kBLFqlAYyEr4I6B5Ei18GTuEoukL2YQgvhNWI64zlMDRsrZ9m7qXbcGRwpM0KDwolXkjQ
VA8PfeiwbbU7B4I1CESjE+/H95L7vYAoqDTD/xOEmyJ3J086Jf0pIG5G+OGgEEVsN1RHdN2GvYqW
e03sSUwvOB38yGI7wdeKJgm6Jf+6qWH6yp4vqUss+JfRd0PQmTJ3C7t5ROVJaWFEYix2cSt53OBm
leFcynEEZttrLRFyT9nKcCXy5vYuBTCTVa/p6K+bIxrGR2PWuZnfgzvp7qJgeAy8LckkRBoUo7CR
shqpyHMea+QPoZXxJPWaRIgjT4i71uL57/+dlZ6YzVTJPvN5e9dXJn6OKuM3rA+I9/yQqgpGYsbC
esb4KC4a9b7lPib+Feg588vZTxEXisSKWRcKZjh9b+shsQc15smBnWaQtZhLM2UnTxckLN6ZNFPG
9OCk/ohYGjxHjqdOFKs1TmyKile6f8vrxaLw9UAhX1pTMUuQ1YPKGQl+0A7V21+wdvuaUNDoroUc
Y5j67pg3FNiLIa/SZ1wRs3eA7OMpaEtCg6/qSipCVZuDWJxPuamGV8onXDBQBbvQZrbKmuivnWto
IMOGW/eju9EhgbKv1T6KwmmYjVdhCT/097SZvJb6ULD3qQs+8kHWFG7xCEWmuz79Jy5rFaPa6L/z
rtW1wKiTccsGX5quHR9Nk+HnAYjRLRFpbYaYXK12LOani1pT+RyQMzMAyn9WxQHQNeA+VC5vudCS
qOD1FVzl1ZmsOAYOjf82MnS383SLEc8glp8ckdZV3TJ4Pp6AC5q37zRRIJI+wJzKY9XlXfmq7lu7
9NAO9tEpywfEtc+qy5IighF/waMQMhLWfjNyeN3X3uRACdmDvMAk2qJo3dD+nKIHY110/kwIY2nQ
KZ2KHo8kQy2V1BTizy16oWnTWuBKwa/WZ0yKLFVsqUmG26wX1ax6cQdw+MMYPnBpMCa/uCSPultE
XXI7nyadbx1X7Y7ZOxphAzYSJ+kTbmNbsrsbFlZpDKxof2mvblSgVze88OdadHTkPgiihUOo50Ir
m4jx/hSP+6ZcaAt7fu86YZP3tUEyzRURj610YcnItPZSv+2zRx12FY905wy2CX0LMDSJu8tlBwNs
0JaVu+sNvTUToGYDVp3K0HetbTqRXPsLWSmqiw275d+TFxev9KcqSXXWD8SqH/PVcI/seFDS7Kw6
RtytNkla0QJL7tMceB8Vtx28eC315Xx9QxzsBi5/yf+GEjiyxBHLTvhRM/DQNtUNH/751duTlb0t
ILPrG4yXgoRSfD33lEPBdxFKZIyfV7CIXt6yi8zGpvW1znuug/AVgDydMX2qHN0RSkFNo/b2qpvF
8U3JkjKnXqtyYixbWCDhnQ/d/nhtQiNO+dhhX52DQPJgfNZswUn8Wxcu+KEfmb0x7J6F2FQDbihR
3AEGxR9LstH1Ideh15fIq0xCxOnvd2TvWZc5py8rn0NNZqNPh4arAhsdzT7xSY7vV3YY0oG9jk3F
7grYVGIeYVyhRyXVzAKJFJx4o0AlHb/EgLV01g6xqbF3nj+lDxb4w5Fc79X7+TM3uDkxOEo3J+Js
RPhmPaFZyI4pw8AKRDcVrT8RTvgGXbCgk5xW8jrHhUpoVbxZ2n1T4MH3eDZmoT4YSGo3p1zoURN7
qtSl7c0GPCWnxo/o7MhypejmPAgcXv8nGAtJM7l610DSRLMWAIuxIOXWzSnSOgKE5aPhMLXTiBmC
OYRxuO4sMkYeF5/HlHk3pOo+2Hw6dKYqZ+9OZiRKEyTQJl12eh2xR8gwfQD+RpQhPFwgkuea+6cb
LtHi9mopkTAcf/qNypTIT9nkiSXlwFT7hF/swZN427vhVfgKkeOyi3Q/1GPEXJuRWv+kzttpARf7
pO5oUOYL/94D99O90717jFafEwi5QXNMcII5iqNcxwrQmHouGWnWyWZ76JDAZr0USNb4W6/3JZFi
c6IgpGCvf+hHybGIg4DHHwESbtWckptwzc0Gznc67Fr62dEiJuiIrhYQQ6N17XFC6bPDVB26Ka4Z
oWo1lgB6Be6/113C8g+rV/00wQWF6ax1GtaAFvLTp/BmXsJHeVEpsEu1b7FA5ozRmgcXgNTxZjyC
ovwbrhhYD2HcRo0EEv5nEiqgbe8l64FV+gaK9ZkG7lSgvWgfatSJnKIvaYXQ68ZSKRadmG8c+YJP
k3VHUVV6uE3ZwpjIpA/sf/tU6At1V4BgF+fRF2CgiM2mLsLfhFalVHI12O85Hyk6w6lf8Z3dOzIo
1E8mrd8iiwE0bscJGx9PW2zk9rMzA9UHq8/eeJAQGAU2wM3/xQBY+2m7prj0gqJX2tsEyKxErUHh
SG/mu1BP/dLMcWq5wtGTEAFFWvVO9HsThu4IkDK6Bi3ey/61xSZu0RPhbbG1mXVZK8u5F0PPGgmj
B+4CU79cZPomV4+zOKUQ9k5otNaCTzpQMsVEDwSrPZyaco99Uy+vSvFXWS6tSavlOYmolgj4lunI
P1perKLIc7E9onqja964/CPMInSPlYxkCiVzBEDIy+xUWAXpvUTdK4WRq6wa6dxlkaxfskzgKd3v
9uvjVhVzCHmbRciSnke+89p5U8d3h9gSo3Y0sLx1bZbpy9aui1doL5oILXFkKrZaTmy40/LCU6z4
VQHPH2K+/wXaj+ltHuiJu++XcsvcsjZgo2FH/wTA04Iuz02B5D8AZO61YFCdlbrCKjJWqKgfA7Li
65tHaCz06qlZLbU276BoMbMwSgxOjEH7qpQCDctXqicKXTfJ6aQXhScqzT8wpKd7baXr2ejGRwdL
pUI7stSQBq112j5IhG/kCb+5jgTnax9OVC629wECFpAkEqLaqwAU+rgCuLpXK+m+wduZUQpRqmJc
h6+kUg0WbuGykL+0Zx9/keTNNyl/0vNSrL7IOCF2BhHFVSFXMr30RJqMRqkP7ZUJwEJ4CvmURXvX
X6UgzqehnAtjwto358/RVmjSNntLEhj7LO8yXOJY7QXVhinrzGwxmgIE/9W+2rLv80aXzJTRztjL
xwgRl/T+ie4V5vcrb/Hv/R3kUPksV75VtOzCbN+UNnacdOADbCktNMxp+/3O/wgsDALYzoDOEdV8
8b3i8u7Zakdyyky7Rfjs3C69ArusNHFvyBiDVsYCbKBgWlf4lNRynKm6PIOU0fBAJPSy7dAcsSjN
nJNvKsdVEUyJt1y0TCfz6snkx1cC1dVtY/GzcPXupkcDXTNj2ERs0aF2lnXakPD8okqtNcFXjheb
SJ3WEO1ZAfwjOOtKGL9GnY/YNxhQRzWFpUibMgi/gBaIiQ6qmmuPJ9SWHqlHjFQthBCk6cc/Qtzk
iejjC1rJMCOzhwh8vOjO8tGtZ1GWwd1w3E9okMWEuKyihnLBTrG/cj+/2QKCKdc8Ef3P5npK8jzg
PcRMNuTJWkU7uNULRRbCjd9OaqwOJIe5aehzWc3Y6EWgTmsB1FIgYHZ6r1b1/+rBLiqixdc8ivfJ
uDb+tDyavrlbXlm1fNlo4A2sI5U6Be+vTUeZ+7Kgk8+1by9nyh5y7cR/ppyGmlg23Qk3wYmsvWaw
Fp+JZiLwqz4P32rJxiDYo/+FW8VtSRVATh68ehmpL+VxkK0Fq404A8TGEsDaQNXhGCo58n7HTesE
qgWUEhVbAx00rjVzWH4E1I4+jzh2dwdbirhCIIW1nKO91ryUJQNwDf5Vbmu7DHet6HlWyLk4RoIM
dXmMEL/KUDnccawFLHPWPaIZuI71M8bNBgI2U3nfkLS3BuM2GcX4ikCHomaAjHAIFokSnPey8vKd
6FXDWKVjMiEMfofXyDZoOEXw2sS0nILnO4IZZsC5FafQ/Z0ostKvjwfmHlvw6+9jAinJKfkO9cpI
GT7029++nmuQXQwlLxKTnGuJRN46RDcKbI8PMGG4WkJ4T7qg7ePbesM6M+hnOjcK2mBv+rAJvi14
5ZUof07z44LsrrAigYdP+Qoci8naZwLO8uxOboZ8hqOH5uU8d3S8Yu53wX8i4FbWYgz9koJJsCey
/XGaYGP5+n6jkUrnDvARdRBHMbc8kNhaYq3yfT56KWOb5j97XUX7hJyzT5+5LF99gWdWQUVDuvEI
tf/A4hvD7rlpXUBjA+46963CY4NSZHB9aNhLVk/6+U3rxYgTZmJfBFM7U9loCSiHwG2LxKi0wZxl
bqpBw4cZ9xJ/GAle0gbxMqfXn6+RHjywR8/e+wH3kSmKoXshiK4zU3wwBZ7bVeTYZVDK9ZR5Mkug
7cY61PNRFDgXJYZ9tfnJObSvpd8HTyyi9PdNgg6oJ51XqFBVA/BKa7ZwT8waKazgZMbJLbnlH8V+
STRRS2NiSr5czkKE1z8Ob3jcoLvReczmCyB79vxPyTwbufaU+mQBtF8PFDI6qT4ImH2VExGjRZZp
CsLtgquy4H8muJ1DHHDPAjkN4Gx2EBXPLO4yNLYfn7cl72jm6spr84mtWHrgFAE4OYZ0hTTZ7Fh3
jDg6IEAf5FaBHXzaSuLBuTHf2e/3KUuH9RxZGjcT8qqTTsFO3p+Xx7FuGBVlsSwlqH9zbyjz5yZE
+pSnY0ntD6qoYplprZdYeHxRklIzeygBBta0A7T8sPg0xfpGHOvz0ty853Py/bp3gnLB/JhG/9HJ
R1juzn527RQZ6sqWMBduUOYueAMzETwH22dvggRhQo9jbSIUm2CqTGqtX5MAEUatO3nXG9rRhkw2
q7QsgbkQiSx9Z31u9+pfuOzrb4tjB5UXQNOCJS41KMAROt5Yo73W3Gec3Ep+uipO3QwHnMAGexg9
xTlXYdf9kG+72CLmN01Flv4jO1N5CSo22f3qiY5EJlFhK5U5PmJnUYrSJj3/oxDqp8a5HbqaSDcG
GTgfDS8SM6zGMn2EKbYE8KoKtWH8fPCDIf5TKDhS9AdbrwemrjQsFhHgYUnXGkG4Cuq8suMDiqGC
ig764CwpTrYbX2KvNo5f9n7v2WKu2rIj6O1TFtYvis+IwL3qzG5Uc6+nJC6UerL3E6ueF8i25TtK
q6Rfad1/sbqCAEj7MWykUULna44NVWjqXT+bKWDGImSlfa3CDrsIbY94wMVvX0So43G+UWWrH67V
y0wS6RG4RiZpv6m6l0PCXNywpry1XK7V3jk2ohxck4wNGNp9Qj7XxFPcxOeT7ZKJpblINMI4iOAt
hfl+yTidAWZoEuhPT5e7BXH6CzE4oZJPhPeeyvk+R1JAWr66jirIvm0iG0Q6E75gqFwJ7KYcXE6T
MvA+nwT3tpWCewpjqMwSbbCW9kw+6ks9NawdmTMAZGL2s56fT31CmfdJc9EaB/VH+h8h0QSKbT2b
AQTX8KJWkpwvDBIog1dxVNPSNc8pGX8AXudxz7t3UfU8o8G8XGOAnaSVHO9P8PCEMNsiIa3JInLG
agVLCB1MbraXUX0wNxNuqZOjLa14kUhQRnQWKY/6uW7pD/d7+Izm/YA9ULNMCpCMQNs+9bh0+ODh
E1TzAGZjDyiKwzyDaW77VnEaVYo6M1KPwmS6HKm0CdO98NNNL2+C/bWmdx67vnyD2DpW189f5QBI
ePzqMvKDKklOgPyYM5jK6bYNwDReNh2QmZKTwV79VOrKpyrs0YbC4DSCYHe1iTfalCEBGP0bNjYJ
4IphKS/NoTOg3QI28eAzKdOUW3UDMVcnm0BkhyCHx4p0drtJQPcTNYcLGK4yyuhEVky2LLSUYV/C
eZekUpmb51UonoLIEScCKgWvC9CnFQgpss/z9hG+nP3t9+Doe+VeS6Va9sJC03i5X4nqowinSKyJ
Lt5ySYETGWR6NdgdhJgApXYlU+8fM6+j+ujlXAG/5OVKYi6FP42QQ1y4oOiecYuKSF2Fq4uouWK4
DXaqGq7bZJl09c2O6Dv2VjHXYeeW+2DImyv/xTYxfP1TjPyuUqpIpJ/HA0mUJe9VAGgCpwA6MKNz
+XwH1tbttwrcz1uwolN+26lIFPkorFNK/GUOWM08shEFc1HGsJ/nz7L+VH02xuobk/BTzI0dyG1K
wyyMTnt6k1ZTPNZrIck5dBxHcc6DsXKDJ4cBqaWoz8PoYyb/D16I9yJ14dR0eiT4Ccgg42NycB6E
6yZcS58hpKtphEi8dxvv0PzC0Tnnw/kIeTcOUBxVSEFqneoGJ3col9zB3wEIzpyT8BnepmkEXx16
vW2txqp2jnWIDlweDVEdO7TaR/w2gByzn1Dnp8fzOEkI3FeucuK4x6Y8h0qYdUmnJjz0u+WjaRWY
9fGQhxTlv8PieC8Kd4/9hj8HgTTxXCHZADz68efeEtaggdHt7cTxKp0TSwa8DxZ9X+1/OY1CUBQ+
OP5+5efXrcV4WKsrct2KmCR0rfAvDCEqq0+SSSZhSRE+ZnufHbCiY+f6O9NoxPkiHG47k7+7QziM
Pne2vPSHSSDdjEgzyCnwcawwYDdcdLobIKCsedVDX/dEMrVySXnpz74bgjecM23RArlHOMmvwUfA
ryROKvypgDgZqXSvsgBvzo+muNqE0PvC+g4oCBsu34dulfmNJwaAofdtQAplOozeGm271QKwY+fj
lQeS4eWKkRCdMc3WfrlVmCWMxXCxHQr51PBbK18WmoQNnKruz+2CvaipzrRlZu6f6HrsEKZhwaDa
jozS9NVBDJb8FK/uqalhBzuES3HFw5S9lm37Jm8tmHurqnv0ywLAtby+5xngSQJDpUhXofZw8FC4
8B5KdFvUdVKQFVbkar8e1cksGF6qUfHzK9idwaSyWijygVbJioJlGmCBlYaNt0p0EScPbYQxVhoJ
KdDK51gnSOeYVZGmYaLjnVhh2nK5pkVTj0ET3potyZQxtZCic19dIJHcXaFsmL5zqXq9IHnk0SdO
rFYC0/ncLlRLWmu6lpQBFIOvZlE/p17pt4N9LKg5iN2ZvUC1Ug4qOZba8CO4OE1x/8jJR3c8D0Nd
ApnO9dUNbYxkTwQjLbwJbej6N5onP2Szs+T24jhVswffd+6LjvM2jJoF3Aa7n6wckG/SaBtK/dDD
HxEUOf7JQqmM9c2z2We9+9Jx+H/vC6MT70MEk+k128tQqyFbdoA+bsNTYc4EXDa1hbRPvwNUXukF
bTz5cay/1or57zew2jk1XAaJG9kCynUo2Ew6qHFCs0FP/PoOaW3j1PblwHyHLBSobART25F3k/lK
ZYh3TJzk16XTlRS5UpJAq+FBN5MY5jKfe62uKccRxm3WJvo7yoRKeu4vc1Gclv6gnRihzf1MhTAs
WoNaeHSls6bMFm9UCgJcqp04XqCnjTaH3eKnMfDO5QjwOUa/e/BnlSxWReuNbqBPelM9VoBsD4eG
LXqV0XFgsvttB9n9L9GN322/XLCIRoN9xuFI6lLZ801IFqiVlKHkl6urBKuTPYPbJLAOgFuYzwdA
i3ZmQov3RpRPKFceWAOHaBCQmkTtF1iY+y6A3vC9voXgvguRWAGb2H8aT1bNRpYWdjQNKureJ1Fs
4tafBa6n5VtzG7KLnvsD0JQ3RZo28zCyVWiGrPbapKyU8c7u+e4l05fqHziSP11Z72nXW1rpmbZZ
hsJn+fcm5HGDAgEYKfMdF3tZjyDxj7k6xN7Sv+bJNLSONMqtJ2zesX7H9uO8z40CqB9K4Zh1aSUC
fTCnRCb702VHNeF6V0AG+Ar8/C/DAD+AmquGqGBrlXx5vvZvE8b3eOW97TdjEknfKy/iEdWHfn7c
V/g0WmZAGkihl9QbvIXOhPb5JrUGuwj4xB7T2pqqEzBifeZrrRQb4wMgaAr4w9nZ+fBSB4mBDnXq
E1b1poj6NzeLUs2VUYUbyhSp9azGMCqW0Mc41akQn6C1jpQ1Ch3Dkml8ynCXecYihRrOcsum3g7J
b+UHBz5Tf7t3HlDBmlUDbUUe65cSiywdlM8W8vXVPrIWj1mLyCOeELu+a9ytF0JVx7TGYAXLDfvj
9d/tZVaYlLKRxifLphH718jujSxDKcl2uDH6my1NXwoaBLLvmnigIqovzLoxq5f144EIx4Ax38Je
OgLOY8j/6iGKC1XUOWDbgEROrynrwX7U8iiT3EkQP14Dwn4ZuTpB+jJgixzkj1feYQOa1RnIChgg
8Pl9a8jQwuGMrRG9bsuZ0x+4HOIjj6deMRBsNsVkCZkIiCHXOc6cb9DaDveo/BFML0oFd+kVkHRt
2nD4LnAqpzdFKCXI60fMpX391KW8mWWXfzA9/NlnWtflGm7i8L5R/9hRAkRtj11DRiLKKaf6xN2s
DkLGBnj3U9QN40VmrHWbZ7Jvazn17pggVTL/B8e//sMbqIVa92SbfoET7goBhdNmv+23S+EiRRzj
qQovvWcS84mk5GzPCRr4SigQYUfXWrFb0h2R7LFsWMua4MyGRYOscHt7Gj74C0mvUG+6/m4Zky6T
5PQSojX1U/84ADGIsclYDX4913BmeN0/pIAoY3j2uCxbI6VMj4+EbYoX5AS3tyOOaz4G7nAo5hT2
YEUOPN8PW5JnSJXDqJNpHyXbTFYblGyCUi3bialfdITYYiLFA10Biv5i0EH7WOZ1KNep3N7pl7wt
tHPXwpHVJU09Y1uQECKQnKDrqGqFyJhF+m23p4j1MBdbFa/Iur03d29QVaJGyqhVnAJ/Vm8Us8sk
0fAszeVmMRu2ZR5q08UtJLTtCTD5/4wIQIbS+pf16p36xO8vy6uEOWtd1yJ9d3k4dE7MPyyq0191
2ZFeWYgEC8KI3SmMsAxkXmkQaSGqher54UgQNnMqKbL2iwcm8AOmabKtJe7YeLumhI92oKA5AJam
AyxtAeZJakkcO4og4chrwtReLLpSUpmRw3xDYBoRilFp8kBWqudNnVDYgdD6ftfvk8ZobiMWrg3C
XA3zXuK/oICvq6DEXQ+hYWaS0fWv0jnt8R1qcwzOXeumuURoZJ5WL6Nwsr3WwNAEM/GbBRj6QQDr
iI18m5r/m7c51+39k96R8NLNzJVvqnZLJnxU8PTCJ5/SHY0RyZjdWv4F+Q2kfgIAt09FF2wty7Pl
oa6dJO5DNUc2w63z/Nb3CKgpTBkToVNVAGuCckOtPzjaFwmHeXZIYaaP8C7eQd420ct02hOltq7u
Cjw64rsRODmTCWuHUuLp2SV8/FDNELnGrpc84s/T7ZG86H+jxniHz9Jkw3/4rzEgxhJQE15xdRan
2HlfvzkdSQ6CaTDYFuIyMRLCreVuaIJvPWeT4MI9Nfgpu8JqgwmeM30xojHcMaCtu3UF3Wre34N4
hKwryOJfYM7ddO/7B7qaAELg1hNKR7yEhuC4KTQP3mZvRV/AN4nqB9RJnA1F7tKOigj3pHHuMOdl
NXmnB0m/jMtXhNmoMhVIxHi34iL52+TYiCwj2n6iPutg4BhO3l0dyubPcTYYlzZReRPeEpHz/rsI
5etzo7zcE3bhNclca5XygeRfCXyIuoGNIuJ9w1D2RIs4cB/HFqFpwpcBeSONq6eOez72JcemKIS3
TyYvCRh1CtmmsL1ly2cYV/l/Kl19aTCyEQPTXOLEicyQnorjzs0WUkbukn9xWamBHwjXR3wvGhxw
FoUNRGh9SNZ9dO1OMtuk3seyVVVHxOxJsNuI4FzN34LVK6FruYWbflc97QJN0RI7mpuwD8bjeRKh
T6VFItIqopkJmIe7Tyxi2hLMULed34kq/A17czo5bDx4aZeEMe8THzBX4SMPQJtIgrvaIbjreQzh
vz+Q4n6aqGGTtbPRCrIhgPL4bOVNppVtMoVforXMuUry2pAwwd/VEd+bWsxVAKw6iRjoV6NSr0Ey
8R5h+lgvHODXWaOc2YkaNBAuH6HgHrjsapDFN0C26eW0/meflCGBeUjP/jK6I6qqdTqAyZmkBKfT
L+EPmdAOc2mGTOkbEG9HDdj3uTw5joRb75dIIbGJD2eF1W9fARofvZBUPIake7tsWx8L41c93vVn
LE1mgYL5zwMkm0rgzhT1FdkvMpqO5T1ygXb5v4jmAJeMiETOG+RvgPvKwotQ5SId6mn0ySoGhInO
8tpfdUQJVD9gKYNhmt4J0fTnQmW6CUvFuUosimw6aCFa968H9tLwI/ZOMQwUpZCSLCm4bW7GldHJ
5Fri97uYbbRpROWk2APcgAyHbJY+2KaoJM6BrQIqFBKBG9WK3h18txSDMATij31YhNV+HDit4Ga/
Nw4g9dSEHUV3IhBHIh6Int+MwM1Jka9Nl7Hd97NgV4lSjR2Gi9ur4P5EOKxQU50XNqAza9w/R/by
XHyXA01tKSRUD+lBsPKRx8Y4DKxKdhlKBc/POaxCV7qlJOiPdTYnyj7McuIL673KfAEc+5vXqAUP
i+YiRyzQR+X+wDcnjdVganZyvDcb9ebiGNbg9b5fEGdaYcFnw2n5CJdFzDv+ofL143vcJWhOaF0n
9gYI3egrzcbxFbcIU78kSQVi33/pUFY1p3NiC9pM/0lbB5SN+Fk+JcJ6U7BfwLvWbCJbLjM+B6Pu
OVgWBdDoG//QEoNFKC9z11GAFGBkjgf0FJbEHrll6lc2fT55aETDY5T5bITEXz1Tjlnm3qdR40Uj
aHTnifgZ2hValF8BAn0wL2bHKcIacgcKBmMId54/Ch+HRzFzsTy9KJccLLWtL+fS27VzP/i/dkYf
qgYykxXyUOd+iDcVhhrk6eJI/M0ykoPJ4erbvgBy+K05F77tqllVOCKN/7clPSWultYfOJT2Qyy3
7SrZl83MMbWLS1J0zruGo4m3Kfd1JQfiNCxFGCuYBVBVfUEOwXQ8o1ixHiQQuLZ86LQjbprF8975
gvdh0xKApMpA9AIqJ/e8+Qo/HoAhXsjNwlZHutB45uvZ8fXb7nInKKOJSvqUtrd/kP1K+XUUZpV5
L0nScXu/f5M2hqytowHUfRXhQODUGeSmIn91N01YWpyXODbGZ+LUclRD7jVOzJXVmkuSYJ9L0hYF
TCAfLOwo6A0yPmm3BDUs2K/BeQtB4qBoUjO8+dT4ER7Lz/FEAHBDbOumNeEOYzxIzZCpWO019R9x
bRbx01X4OWXt0B+aPPNHJAa7rtyxZjJvyocPwK5zDYvKyQsLeHbBh/VHbm38LFW7rbfMfeE+AQ+v
EZXstXlKasX8wvpGoiq60JdDc6uwwaFoO9harN2jDHX5zBy/i5KhPbfbpmGL7piJyC8PDGFOvvIO
0U+0YFqZRLw5hZu4Fa/GphP1NoMGhgYs6kdx6Cs8QUuzJ3XWS1jEI5SlJWch3+pmfeXblXhZaxe9
T+zo3IEXQiMoeJNygkHwzk0IS3o5WcctcOlLbUEX3iQ057Z15Jy02QHOBd60znIs362m0McjdMmn
MqbJ1ZiKQBUC53Scf75zZeTSBdDWAeSww0ESQCEESogb6IcFmQ5CHBcMowlu2Vc2vwF4Z0y+b3/r
TaiSgdxVBWUR4DfJXcTTT9NC5ZbxjVRuffIiFmCKHBI5hw3AzvJUZtY3CRLOp/G1yoeGnlYv7oMK
eEjKXytWEcu07qfA2LzwzdHzV+IwwUHxDoZfEk8ZpNrBH/cZrSywwUUUUnmBGajuOJV7QwY203H+
3ctpP75E/r22hvSpbckVj0no/7y9aMXj//XOaEaUBQP7wYqM+lkO/NVAG9mzJTwJdYLoEER//2Nz
QKrq9fifUKS3RM51+D5aDuHbjj3WwZTRgObDyHJpBnynYgWFlKOZ20yEij5qZH7RmmA1qhK09nac
kyhXdHI2l0qNS+dTulAM1ci+HpZayiHzHQrOqGf9a12s5YEK4RsiDppilZ47m0qf58/pgfSnM/XX
mu2OUj8+JcR5Q+HYais94AoKoudAlNOCtazIDcgUfImdYLD3t1o9+M7qjqLQxSn8e9UaN5E9qMAr
XvYcMKiOSwLClMwioNUq88WZHGyHppH4Z1iu9IVqijRZFsfnQ+o/rN0MUiNSZZPHgnMrm/JKCL7q
NfJIflIzUAXLTrRW+q6HlHYzaR1YXbbpPhHCSX28D0cLAdxZwFBCXZvaqx6W+6iIRwjYe0J37bEN
nSUnEgiQC+AyZxG4W4Dzt53JlDayUbg1vRBJDRKFAIrnL7KBYV+clNy1M1dOoxGFIX2LM2cKsdgB
AYRZ+EEI4g7zIUfhHOy4psuVO/K0EP37PVEK/8Tf3VX8HllP1BbOU/kfmp0i9dUwPf1KAc5b6rvJ
GKMngbT4Bb2PFslke78e8GNwIuE2TJSbaptlT0UpE113Hfdn0gBf/3OJ/wCozOiRooE2j2x7izUt
49Vy0eO2TVXf3pkygyLkLzKq6AiPx2ECZNoH9bmyqkj0sHngQ39W8ALvlz7SsO+1RCvGDygOAVyV
Abysu04wuRz+RtP/L4ppqMMmp85kQiW4lwiOG1PZm234FsOnAmMOz6SX32gArsFHnkqY0iEitLVy
Lnq3KPoTPw9Ca4d3amwaTCifDgbyLAxMokVvlERggQQEsVmsQHXNrk1Javqi3WLvtaWZPnmP+LTv
JFoGwOiXF40AurCpA8IC49eLD39527SNrn57NndSVARRlroMVI5aVgwEwiYhZwBxMu3RzR5A00yP
LXaDUI1jWNlRwGH0BzQnQDeC/Yh6TLPf2Qu61GBmo5ldliDenlTHf2KBvxv3uEK9RCmDyjHq/p4c
MSQd5/h6Unc/Hvdku5C6VJZuB+jaXbO2k5TXxhIYeJVM2boc8IHPkr+NN6r6izXcnS/is1XWfjus
m8mFVHTcAqxAkHeW6yZ4hLl3Y9IVi0E+PmMASSYY7Lk5wlV7qICON9mc5z1e+aN50wT/bnVbqHI6
LwnvseHbx9aKOwewtmJ89WiEmFD3X0IsmzfzB9ilYaqBLCBrxkqIH7VEiM+v8czNkce498axuxEa
K4kOYnufrxSjJrCS1b8PxSTn4ilbQaxmd4rTwpwfHmLsDeXQbkt5vXLTZmpq+Mu64I8Q2xZIMsUp
7i0NDR3clAIJ1PhWiias4WaR6XfK4jm8n6nuuuEUM0wT/SH5cU/pqXemRzsm7JpGifWrp25lCwJF
FOhxfhRGo2cLXTUpyxPA36RHIcziXx2+RpWVeRBuBVg6dRcFKvgbwGBlXMr70yheIBPiQ8EdrDKE
UWxEQwGBwgW8xMldqGXQa5IZJ37XCalwBeYjUXRNx/kUohC3qcqrPCls13zG0MUOR3UaGbaXehMz
A5KxglxFqvAu68e3JGUlLZ8sPNRzuidgFndj1XwldFH0iVj2MhYQSsfiPl+MMISX/18RS0oJ5Y31
YD/vE/okQ92r2ZNaE7XgBvduj1KD7GNDPinC531LrLegWCcp6JRu7V1gA+3xYd4BrgSYdoy+2yhZ
ibKUquhOpGcVaG3cmioPni0Fam28hJSZ3rSvzYT2VTAh/2pmNeCZVPVoQeUkiYufC+eRLbl63pi4
JS1XAYVEWusV1IyvXQqZkwzB7aGv/6OeVaLZUjX+5aOJwFU8N4JNo5n8guFIOHVpeyv6eU7teiW3
u22R8Du5kL2BOR9INjOGdKshD8qwjhK+od58MTc/5j7c7Py40Uc1cIYavOYrxL/OT7WenJemvLhi
hUoV0JZZKCFOqzzpnIRU/xxlIwK9RzPl/dpAIA6IJQb7HHR6qDpZ2SCMHV3EREODECzu8G75769b
xD7pVP0Eji1qGTMq7Ilv/wwiuQb9P5u2a1weaSnWnf1oqnQhgDruurLtSMzLeBXr0BbFVhN53It/
ny0r+lMe01agbU7YPDffOijh6uNXSRbpSst2PL+4s1b3EOdMXsWq65Z84C6HeLkjx9ENTZkHfzFk
kEFyIOfu8tpR9A1/surajtoR6s6hyGh4p4iy6plAmuOpo/UWLSsjzoa+RSHSxBYvz6GV8KewFA8K
Zioy7LDCRHFVz628Yya8kFvcpbs5iikVtMUZaArSflpROWJT1x61gUf7As/rre/pGLWsdJhRV6QE
s3fwgefE7mjGrkBA3YJK/YB1Nzt1pptWvFL5Lk4xIb8EcMXlLVXLPqC8mQtj0H5fGNlFBemOlC7P
eexHtkTQK4nCw3BImBM0zLSg7pn67bA6V+xp9zPXpJRz91++eWQ6YV80m5Yku48mNgBuB4zyrPPZ
yO4nM1GtWrdKvA9nNyD48u3EaxqAhRd1eJ+sdNL5eBt50wXBneDBZs2TtcT/G6UDGA7BvGSPGuaC
s/sJn7jo/+83DgxhKqyWSsWn79cRsZjrBv5pXBcZMot3XB8XSBRl+cHRzR5L8OqQ/VKpk6FDHrIB
yw1YaplKIOe21UB33KBeQfGMz1+cN002sigl8O8EUVDCGuhe6XsOGXDvPIhCEnWDzTrlK74hb9+d
f+adE05JQGhaLxXoV5C1b4EWE7twF3qoyY81+3B6Rly3xBTmVECpddAzm1xpBFKrnx5M8D/5fsRu
rvpzMa9A1Ysusy1lZLoq0uus1czQHLv3Impgj1tE+opJPPixHX7Oy6e6a/la5Z4bMTWn4iu9dnbN
ZtBEU6ajC9zhzDdhmQKIIzHVRTnqAnZEL74SbmgruL77CXZkMusbiEeFndEjjz6TYsfOnxKFkMWa
/fixlvyswmHVL/+xxSrxwZWNc64JJwZKxdvt7uiNk68jb6sOb35wkve+ddBTPGk1dg+R7Hg5VHGH
+YnxCqK9O0bWtYKwv/Cy44Z1tLTHWfTsanQr6YijkWDxYK5T2NnVCs3pXNls0TOFIaJLjduDk6k0
IoHFFUQAmRy3Zf/9G6NT+y+oCO4AxW+gMpGFMKFO3hyk0OuJ+ROM2CJrRAYpNXCm6UaPJL6ZRLw3
Te05Wc0jCXg7JtCMcMGhZhO+JF/VFsOLU6aR92+0LCHLXa0OK5KUZyMQUnpY4CX1tagx7kY+RCCh
IB1hxhkxHCIIwDc2w3LJLLnKSSaEnU6GD9nrgwQC5HCxizsi1S/bwjXU0UacOWhohJEesRvmTPLG
5ArrNf7YUWNhufTaoQW3+pfMIeYMmK4ZGLBpTIYfGQ2WOr5B5ucvZBPXRb2hkkSIovOR+EWVskW1
+IfA3mMqKqppFGP4xAaUlYl4IH+CHdt5Fz7PRFqViRIZWraSdsA21GhPMV3512sblZ9VobpSiP4G
1sOsB/+TOlmqp0REpd9cKBUQ9bUMjAR6Yx/COAXDgOEOhqd2/w/Zt2ImA/ucJqzQkFWZyVspXNc0
YwkfkwGaJqWsWn2hEWfUYfZq5vt6RMwf+U+CQARhRgRG+SKmag8pAawsatBeAFB/PoDdUzX4/y10
YUOAIpk74TA+ubzeXqAnHd8/MZ1NQ7AkVu3/b838Fp02Y1rDG/U9l2WXDp1uKgqq1h5ZYr0tsc+2
hpBPY+QjNBSrG4atWB5dn3FnNufvy5hP8Ibj7cgghAs7FXSASf8Zd1+G9qvhaUuKWPZZyppoIady
cWrbSxMB/EXdwMvP33RU2OI3sDUhaN1OOhyTQ1FaocN0jM5AP/yeY7sgKVTQ50s2Q7XEWCdt1e4g
v3RUWbnpQx8/nc2507Qv8HOsf9RjyTOB2KPfaa/KPX/p5pq+g+aWFswGRnbIi/LF+zrB8JQ0VBys
7jSBaFvMsu7hCyhuSLAkgkRCTlJF5oIOS//Pxr9vGESW2K2/OnuacUP3OC15Hzo0QzVxsVUzv7Ab
OJi1ipARH4uKiBYW2XzImxJtCbMlBssoFOIQ3YcHwMwx2g6FEfKm/F9QkhHpARKARu8OiB2lYeRi
e9lhau7qIkfw10Jn28fKNbhm+fZTsdIvoqP/UCs5DWqRza+/p0Z6ZtN8a6orAl9GB35pPU4nYzZQ
bRcjBId81gsxI4O7cXpH6iCP4mc1peu2hTNuzlvwqbBNdmG5uO9sz0fUIoLvvF+ay+Mvz5vftRhD
amQNM2QcvbYZNeRH0G5m8qRv7e83RM0w4ES7YL7efzQca6p8BZhUOT30LMaO3Mbf/fxNvdrhvzse
m7I2Ewvdv6u2A7MoUloNirbbyu0ySI7YgOexMEpOP2aBBtLXpBbBPX0ld0AmUNs0jFoPHhf+b+D7
WFlRz1UETTGUKNdLMa4yQbhSfyAcz+nNRaMLAeoWLfj5eTFdGNMnUcRCVVVK250VA4Q9znscXJTl
7xY0irSoogXNJd+T2p4oxokcJ9dgLxaki4MIH73J4p+P6x7UpfZce0d5mziLp++Fvvq6fECsMFbs
rpkVJziYM4rIzxfrgMEDR2ZwYQBXKvVgopRsurcFAd4DVC4DfHvRA4ZqB1cjrZfbgkK7+EO56J75
8owNgcChHUWex4cjK6W8yO2hhcPALtJHeKJC0SX4t2uPyo5whJseug9qyW9ZNpOV0bEboP61lKoH
j24PwLjkpl3sgURGuugBsBtkAWxxK0/coHxNNhiyP3Mu950XgjHcOjHjNP3VQCPSsEkCnct1NPfd
vUQALNinI5cKDBfdRb6n0DEul0mTqdHQyjvAW6tHUqPx4TrSPlnva0hbNNsu2q7NvVrwi6ZB7EtY
eZRMxN42dcG1LIgkI4E7tcY0+JpocGWqTC76fLctPCfSMAchdmJy8YRSyyTvaeVZxCqHoHPgO8gK
xY32HAVZWjkggMvBOlavDaTE32povV3hJTxi4yj89auV0GggC7GpMvfIhWvjY15TS27nbt1uzDaa
h0l0pv7J7IY/RSjkKabvDvlzvamHfo8OvIjew2F3kh/mHA3TSR8goTnUknWT3vw1u8Q/hiEspmoN
9db8hARGaHCfSEM67BAG/RdHJmDwwtvGdplMCspgIEtK9tXV71FXkVmMqqfSFXKXtxeBUDaFeCHN
0rjxGFyWWTlE8qfyiXJvcORFILcMYMVI38rHgAnIlzcP9gJWYxpJPA2V4Az+YU4lrnw31MAbqmg8
g6SE2RJxk6qsy78IUF8R1KuXWtaNqqe/gISjb1l1A8g8acSsESXx+xKL+clbXuFZnAVJSdHSZr+k
vzoXNuWiW8rxd/PnuIjLSzjC3xTumM3iYKUMfPfDH9ZnescIEqynSWz2F5poUvalS3+l/6O5Nr/Q
CtNwWPyrZa5JydYhK4JfY1m/ImvbOqt0yN3jvS/0ybRz9+NCOOBMOXBJ1zwnlZ/CqTKmlBkPLNwS
LzsSD4hR4hpOx0X7q7h1Tj5jn8zyO8ueb3nWXBGN4cLlNRZ5/0AfxgfBDK8MZkY0nraCMFbRPdDX
lHROgZq3ebMvt5i+beYe+MwxMxbYZymrxcFA2uzP/OQ+cttqmhk51aN7J5FOVWRrUIvmzxs2I89r
uNEjyp4GrEw70ZtKE4et1vPvEF+bQLL3gEvskoWSFlHQvXZyEI12DDOT+9ClR/xrmEwVLmOJk58g
Ixh9kajXughp01jipOpxTkOVw+nxJ4YhhomofL9ovWRkgUuGhlVrZCnd3ij0C3LahpOOVUwcTTpQ
glwjm2m6EKMgaJV+8ZpZCPnhdOzpccUOYGFh1uFYVPOMOPQ23+4pHCtMWcGhfoF+EXUWkhev1CTr
kSFbwsNKD2wkCIHI+d5yYgP62hHxtdJpTObGvBRaRAuK1wZgDYBv7I/6shGI4w9CWkFH9MvejO7k
+8MefY1G90g5T8oKTjhRnU+X9q1xTgPutyjD01RZrCVXaIsBqgw/BK0aAJ/ncQB/BVQQyYax3kig
yZv9Un856aUk6iMJ40mrnKvx8dlqRMSezoO5H80adiBX2bOMD4Ru3NUZGBxneLRzDIbcC4+ygyS1
irlsF13AAy9cUa9pS9DO5QK6qReir/8QpEd+fXeK9M21IBbq9kNHd+ekXB9H7KYmbfVuRgC41RjO
eKe/a9Zjpt9oCQ0Cy+kF8wEB2UP6+s0i8P4bEKGEYNj00ZH3nKtSxKgCDz7RusdBtaIRsk2WG2lQ
prjiiTzN1I9BCMT6BlRSHKA1SLHwBFd+yCdggRR8aJjLrbxN0fbMufB5v3UTzo9tAqgokJtRR4HO
+o/Hae+K03aFGjhCssRqYZc7TmYI24dhnmxeLJjrxy1LJjqL09Hths+jSmgajKEFbMRWnjE11TDL
6HfMTMvczAqEE/xPqhYgcS2vx0QSICpG2kwxSgIMjPUhpfVg5lXeUAySmZKPmu8uf+kVHw+jjS9g
tvxX4NZDN9tAcONcoVEqRddrzN9XOe9AitbqjITVvSJyeOB4+eunfgIPV8AcxMtuaQkBMAqyy5VN
KFEp4ssPhaCQl96lCqCyQ0N7E6431iWb0jo2nh/Q1AVLaGNF/0rCuqMpBPc+9NQKxHXA8ANDcYc3
Xdu7iOhaOjC56Qd9OGBQcdsv2m8xEh3SAuGuOGPWhjFlmPfROaxDgpIief/Xn+Zo5lPbq5lFJh9G
Dy//CRN/uBqgJW/jaMeo9RBxKQw8F2E8S2EMU4biGz34pdIzac6ZVSyxiPD/pXHJLuNcqCAn8s8e
nARS5jGdUiFbP2VKAFTh/raF9jg7WRSkOmLBWq8dXgiNeOoCQ0k8DOTaBMSR52kHQcr+eYFKe/Ky
6diegQg/cVpKWSMtC040uIFRuX7VzD5t5e3g6iBPDyzkUGdO7J1t5IZOgWK1b7pcZjZWGf6mRyWA
8Q7xVXTnnqlGUj9BMSRPA2G3Iek4k+km5Der9x88qXjZdD3i+338dxh/e1KfLxm98PErCuuhPw3a
/8A+xsbPnH0fzHyz+DnOnef8f/reIpiYRkRIVV5PNZwufFN60vdAnXi6MOoIDwlaVuydvY2fWmY2
Q7S3LVPJXmxZUvd7KwRWDea8iuzN9xh+e75BjOHVQmu+MLCpxEjZI9SK0sl4K03iLNnoj5YUZV0n
Ks9Z0HUgj5nsTzu8xPz4Ks/V9lvZiSszQM+63IL+btqhReSLpHe3S2MVZqX0eZp+8l4XPQck+MtH
9Bq4oylkKpyi9BcncahW5/UATwgzW6w2XRFo8rUTR1ZZBIzM1IMWeyZQLRSXK1KL3nyY95Ke3Y7P
H9ZXTntiH/L8NoO/YivuSh7D/K7Hd4d/OGxH0vdgknqSQOuzvuEkNOSIXneBOrPqMgvd5TWck7E5
X7WsBSaCz6f58K/8nth/iRkz5a0GlKitJgWVXjoiFIbfvRDbXw1MQkDImmUm87dijFYFYMIicpds
b/GIYZMkFDKPM/0Zg/BhDCcePgHk1dNf6K7EE6LaO/Xnf9Eh9xZ//RHxq7rMWrppVI4/+jCZnlYC
hg7O/Y5AkdV/eiNCGwQA85K/VVO0TyyWeCwg92txFCNjGzsJte3MurADPu3kUfxO86Kco3zFJpt4
XH0rmspWiS7o8OVO+DnCaW98L0IcUtuoGZ/mYjubL50zUmCNrF/d6oKF0pgyTkrj/gWNCU/L/MNQ
2Cb2HuQnWDfzPPQ7r1Gi1T/D3VZYKI4RpsXbmTc9OatHAD1Fuu+YaUAAAw2AueXDjBKGqdAgmrpp
4ftRL9RxJVdM0+dl5kgsEHpW/w2RzqzudhpwPRXWQWxCv2TZh3dcS+TuK6QIp9S4AsEogWymRLlY
uLmDebpwDzOIvO46ofdnwp2+ItgMOZn0DZ2eQi7DEszZEzhG6R1wCyngmCnxTLB3i4hhOLysdiUL
mrkTjvcqM4fFtL3+tjsiwOCsYHAXRn3O2eqNSvr6KOe44i2E9+2TczZKp+NngrF+MAU5x5s4RCPm
rV9nmGUS9i8yUtiOqak2ZpZ7JjFTsTrEK/b6OvC6rHzhqmmtIZbXDYoZrCt5LlUkcFu31tKeVgpo
Yzc9Lnxbzo0AfiDoQlLNr852CoDpa5OXYEOMXac+QOippkJcQH4q7PQFt1bDVEO5CE5C7QJq4vvg
xYFILY+an0wBbgXLCctyVTEAQksBNtHXrUJUXnMGCcz9oCpysggj7tNPPS7hFv0IW5Q9hWn3WHAz
JJYxctwax4xrECkIFBUUbKj2vntTUGJEXGoDiQmRlNSAWtgi5P8BlGdZ/Scb6EcfLd9NxT96MiOH
ONhmbX5CRRTU3scUIBzbkZQBT148nXzyLJtXo72XFEuRuh6SsPNsEvSxgQ4xBBfZCbw6k5uFziz0
pMtZHN/zTk2vj717ZGVC8fc2c5j7Lq2vPYDhQ4uonDc3H5NdB/MefW8wVxGOtnz7hV9CQeThH8E3
TAPX47j7Kz+xWK352E6dFaWrqXyYWXf2CMQRq5NwjeYpKBcu1dtkyVOV2OV/8OQ/pbOO35H0mMIG
bNWD41M4MwYv9wlZNiM3pjm+X03pA+HZcg2E7YXditfIYV/MnZ1sBvnsstNThyeE52rPZKokcEOU
pdFq/ekUAcoA052Bw2aXo8kBDimWVtRQKAUujBk6cAuiK0xDvRqhvqhYgoidbCuFSAEidEn5vKOt
RLL/9jiiWhgNfG9O1DE2FZLcKp/GkNPDdNvCO7ly7VzqbSRsdiQBi3bqz/Usa4MMmWiD3rLYKvZd
4UaNzWzua0681RcK13eRM/o/JBqb4gGeSnhSNF9U6XaxYf7WxT7rnNCl90tpPuGgOZYwx1XI5973
iZwuz8ccyFvrTWq3wXBHqK3r1/aHr7hBvDC0xUOwb+o3wkcWLccQLkWaZFXLJPCmtxdyqwG6kmeO
mYnpyQRWD07YNi5o9epbExamU2qjyx16soG5QW8x0fvXadtbTMAKOW3blAjvEmqm+8jPZjzjAtTi
PrxwMI1rDERC+hKbnD5Lyx2Y6iOpZ8FU7JGrxiKwiRCGA3hjJ/Shwi9PV5mXoV+P6GmhBssElreC
Z0925r4/0tfeSwlElfMEzoycjMCGdK2qHmvvK6PM3UsvEspolylmxq1KN8sLz1U6P2atOg6WR2B5
3vh0iEbMmQsxGeWuxFHjkNDErD6t6FC1WVISIjQcObJSsIKWc3X0uVkpHw5EttsVMvpbYvnv0Gwa
Ildh6+ANIAp7skt7EpJvhw+6mbo+yi7ykPfkX9raPlL5gUtCOjTU0Exb+Tip2GqyYr+nKwlt9mDl
BIsVa5l9/T4/cABeuKoX7JG0L95pNBxC3P23mPzUkdVcXGHOJG+F6a0f8Q0ydSsWuDVbFw5m+FXw
9n9cYplA2W+UbXSRd4ZnP96HEaoNxJgfpuojrAlKyNCarv/f0naSbBOYA0to02nl+jGAW4OGWb++
tfCJGj4wRTyd2bpmtf2+5M63/PhNQa20UlRRsS6BGwRDi+uQsGEJq08x5wivuHK6RNGrl54ZMbto
8+38lOguQEFQB7vtZGfHelQiDDLhjfpey+2l4xMgyhO1fBbNKx0GT/urNE/B8kOT1KUz1fZBfqfl
CvlHv/7w7YdF9Rqprztqnsibh9Co2AEgwTOyw+DlvkQQi01puSIw9GiG9x86708QTcVRLK/s022K
n0V6fJsceV5ZCgMTIFutmruWRhpQxWdXCIW8lJdv6I7DJLz5HoHXgvnVocgiXz+tG0P905JbpNTc
t3emvynwGL1GYr/1ZrjrVx1kSJvovy+QmQ1m7QyYcgNrl+jyvZLB1OwdrebJcEd+KApkTJMrwT2Z
oUJFDxm65pkie5Rhx/IF/HCUFBXHlh8Ugd/hyXQ4ko4RT0gFWrr5Mqb4JSSkQe3TZsVxML0r3ANq
h9bnCMcX5+MnE45C7nD9OiVMN4DdvhQvgRTMRVn9KvSvBMEY2v6eC/6sh2PGk4y9HEyXZZ06/Wcx
8X4WKceHQqbCNr05vBEGbN6DcnY/muK+SBbaOwdlwaY1ivhpMD0YHnjB+f33tT7JKO43K7JJSQKN
sbDpt1dMNGe3vIFKY32Ql1TyhZx+tUHqzn3XtWycOZnr9rEZnahq9Ifq9Fl66YRx8fCib99WFSdM
ieKNXEWovyFUrkUIkCKwPY+C1Pz4WUFD4L5vcsVAe1SXxtshbui76SKHPEqttwHEglNg6eMZdcm9
7I2nSXF1k9tODNo2FxO+YJoglmJPJW6f6PgmIPGISSBeQT0KjGRe7WspocjGd+rhwRu0sN9iJo0b
U07GWjszfUPx3HHpoHzABs6jTmN6KX99k7skfZ7LtyC1fw8oJB00vDdHfCoNbM3fxN3X/NXtB4Uy
j0xZh3HSD03mz6o+2pnEuLC7SQdsxalEm+WFKNjg2wHmBHr1fckv8sGJuTLaLFa9hvS+JxpaWqNA
eJrV/Dm7caKYO81a19RP6S51vvWN7DPSRKrA/h1/+BO76hri5hhIsqrZflkWKRT0O3ozuSO1Y7mw
u4kxpKXbPr+78/4no4RLo+t9FP6MfDwkHm5q5iTLRry9fE2peOTRaKHgS6ZitB0QUn+nSwzghw3D
FSHD1UEkrur/12ifUh+pz8rAlPnABVgGoxhcnltD7FHTSEgIx+TCkWmAh8G4fJhFVcLrMrJfK7MS
p+KXNLOg5ib/CyOlZ/nsYrlUvExI4vym0++5V39jz/DiAIhEvvx6UNEohop2FUsrFF9gLnayVX3P
SlElfBWLzumZgtBsiqYWD6o4okzFszLt8H6IDpaG6+fxXRypZAZ5MwlEjQ7QI/Y6oKRtIEgHMmpO
nYSNjUld5dXTNET3XGZ0CNzP8+C4S+IPu5br0qMK1YhfP9vD2d7w38nWTA9FWFCkEnpUJXHpEMfZ
5FGAsnefe1uSpA7sMPFcpPQ0lNgpa9WUotTwTtD4XdQEajkfib3PO7Cr+MkgS3glqhsZGLDSKbTB
4pr/evWI0wDabrBzd0Czc3HydLHnbFEbdJAxvyWFG5JgXkcyBBenSgLMF//Vwj75M3tiTyp+N4Hz
ZrpJE3/0Ow+HZRtiTHlC6nxT3S2EjylWb48/YTShSZsQXVAcqadcCBzy34C3XzrWmM6It2s23tki
M+VicePY5uCSlAdNABkmGelC6CZ3jheS5HXFCLlmIwKTCv4GwJeFIvqJJjQ//9Ax5yMnGyIY1MV5
lLZ/ZZ/7ZVmRuhRyEpzF0iZ+pgY/EzBOXc5oeyqz+31SdtKoO9xRUqoYxVB6Efdd0Dio36UtlaCn
I0LjmUAaAO++SXv5a7CGlOfo6VLfLAQqLNZl/Zx8vChDep12riWs2NCNk3O8V8V+rbGKcLL4+6OJ
LnscW4DPaNvr76SfiOBbiLDm02zez7hBXrdm40UHOEQqp7KEmoHOYbF8E07Jv5Zrh7h5zn6LqP8f
gBCn5i7mssPcUiseps9cOhqSKNgRUvSgX4PSRkK8jxvnQ5U1sNvwHRs1YgzFGn0B+ort14MWA9sL
06rjmpz3V1LjHJZVp86Wis8P1Jk5wkGD8Aexl8Dak3wti/YGv8Q4Te4ePAesAmbSfkw+okLJfXoM
jpQQMYrlzpREFUbRgo9oT/Rowl7O4zj92/NW6MUzpK7Szv7YowxXYM+LKdLA7ifD4/VsJrkHw47g
oRhXcnPdjrhY++H6EJAgTXLrwxv+ATcnLADFc6NTNvPDu5DRzzZmemXxj1g+2PC1/4DZCxW/NCd0
hSwjGCHXaYZbzsmdYF3hvu8E57auAT1wTsKJPOq+w+1wooVnA7c4gLprX9j6yDeL4wV0kk0cucGE
fiQnUlwsD0GBjjr9FmbLSqd1rdohmVQFPGfNmrhOr25mMObYH54QOL7xW2j6voehP02QUeZb6frw
9OS//8MYKurta8VSUiABcrHa9Gc1Guv86Ib6qJOCEHfA4m88bV7POk8UX7MAQ21wiDc8xCMvg5ne
FkqxzJ4aq8hf8GHcNDPAIqWUcmrEhpWEfdl+xIkM/dAbz0KJvg3nuPicqtgGYtOxOIGBjlOayakC
sinWWvBfumtEG5i4aomCxDDAhxyt3YiIJRGF2DdIXyXzBlrMxhH7O9QtNOHfQDeEzozzxmZfhsij
DTf6yxXc0DX7dLkUyloCbgKYvCmb686x78agPxw5PccQAwjc0zuCSEtB64SZ6qicffn3+zhVGHCK
QmTWa/2oQrwxKyTYp6KyccYWlM11m6LusYdqkSw1Nu/OyWQn0O9jHPMl5pRt0JrkEJ+GhyMNu4QF
D4hcThJddoXm21esVZ2YIpH4Tw4JIsBZDtB/LNX+gDs+J/8chZy2p4vh2sPRtIxKVbS2hrOpSj3k
+zxNQzwn2A4cY+ZMhWcSfhnGFOzh/z13KAleTwMwgeTbxegzidaYKVVmplE1pdeQMk+X1kHeGt8n
NFB16tNZtZp6oaDo/5FNS7F7H2i4lgN3m5GeJmDZK67TutO0R66Ei5aFDolxePo3KchKFPtbzLp/
evSJF/n/xAJFbY1B4v6esSF60KAvBJP9MJNgjakQ8T37aeBTkycGQpEt/rz80JQ5PCp12EMv7zw0
hc/gHIHd8K9czNKCaI4BCbpsutGgOcLCQ0WrpKq15SMgYvZXn0NaUtBd7YX0B1lMXFyzIu61CjwA
WC2UdZ1nZcy1hc9XP+rpNXlIIsSdmX3O3KfT8i9Hi+ybiuNJq5myHudtmKHy39p/TxnwOrl2djei
Aj1uHcTVJo4iO4nXyDP4D+4toqlel0cG4eIQN5vBv2oxTlaLnhIKm3Me0FHLOUyjnX/h0UqX+9O/
DeQw3UqRdTtOoOyLnjqJ8+BVmaPhHOD/iCbNn4AQ2cr1T4l71q+NjajayUYJxsWXKVRAhYdLvggK
nBAzpRqfp00Tdz4KWhhblMJWoCisxsMbUY+bDG3C4gvY/08u3q1CIQ2QsKLNDTDBDcQZt2W1TiSi
PeSUpKHSUPCLndInye9KRz/SU9ZuDJXzH7CPHEDHOnLJoCJHP9JElS4D+TAZ18pNsuZGGiM4OR+n
xa+ldNk5vFG6Qe4E6Yxbq6RZOewtsdxCFWTvtTuKd3CMf4FhfOHdFelh5iB1hSsYsT3fhwlyz/ZA
w5pW3uONQ+XKW2mqFQwJ2iCMFpVQ69yqxf7Ty0WANHdX7d+acGFqJIJ/DF+q/rHo/22Mfjr8RNaB
BZUotYbCO/3qbMa6mJ5TCDzn/REjH3jgyzzb7v3ooEAIWuCy7ahiiUO7PtVs/T4ylkTBZiVdcwTJ
tJa3343ZppmDbmF8gG2xW+o0tR0pUYxirY8Xi/SKKdAfluKahN5i5hK+yy8+4D+gaO4c+IEkYAkV
RCj802Y1sl07rVNQNlakhoX16vmyf46yn04XIECJf+jgIkavafHFGTFcU0dKAWo/EtoAHCSmKg6f
gDmHHHwqPCQHYrc1ohTrC9orpJPMSRwg3MQKJfoTwdpZboRMCnPwm21SZ61W+GqKmRQugkO9Evi2
M8tRkRAhtOI3bHWDN8OS/RyatmXMMybi2vhV1x+EvQk27PPJXuNEO9y/YJlYvILyxLTEvPJtzBEm
K2lrpCLOq1/03Qlq5yVm0Zgw5gkmuqNmeJ5nXtSHs0KNzMixFT6+nO6ulGtOhPJZN6+i9ORvmewi
QbYpmjq6P2cVsj8LAbHo8FwG1wYrUJJxcvljWvhoJYxIrftjh28N593LqwKiOrIPMduZkB/tjkbX
/vMkVJZf2O/04cGi+G3IDrZMvgGTxPM5idMtKUqoa16RPZmiIQ5/8DQRScKJu/I6u7bh+kejJkGE
7i1dMV7GXvI1XBHGrYXn0AgKgGGBr5q48cYbo92xeqMbBAJd+AOg5dNEf0jKJZdQbZc1ymg9hvQu
guNEvpnni1YmHU6DdwpZUJlT1K9wnYJhMCIBtNQ/AubnC5iLzLF1mc4l8/k7NPcZmc/rMQ+8238k
sfe3i0lakvwgfC5h59Rt6Lc7GBU8Fph/tgalNXRy5ZkX+fONGAAlJX0I3SZZEWCYeXSN9mvfKdto
HAJNNlg/YTLoyxmKoQst+360aUsPz8TwbXz4I+9QbRpAPaBa7abfcNOGCZRtAwL/OF+MPYheCg+b
WlX6TF8YAL/4hSNFdGk1Dl9iGR//mtLGWM9Pq8oBW2GjWbh2rgJ/hnmoPScDuPls1P8W2HTOMgSl
Y2FtVtvAASXGjtQ7HKwQH4L9jRLClj58DdBCy/Pk1y+lj9iVegbFdjcgbBRr55mGArtahs7dUX1v
8pq2iP6nc+B1pUDRBaC1A6t7w/ZwP/tNOzjEiQI2mFfW4iI+xPmGAMinVk9BS68QAWlrjuiXiupm
3nw5o5nYBSSiS2WM3t4k4WlqInGbyLPMVmJpLlfmBGSpQyN78dklfjG9lZ0l1rbXQwAb0aMYBFVA
KP3UlEPKQsNhjv2GzxHTF3aYkeqdCGGoc7yT61p8MqZ2Hyh7Om3IuQ5XPQ6UoNe5MUk88ikqpB8A
dM893WZpz20njXUHU8dcq10DU+ByRYPnehvFOKH7L8Q2hPa1FXKBHMvRcb4xYGW2ldCqs727q4xj
OvnK0vcGuAUUna3iCYxqpXueTaRGB/cwKzLpWussnLXgo44JYF7Hn6RqY3LOeo/TdcrHF6dYmEHW
KNiI/GYadZDejbYPZvQqqiDdDlEdyIwF7wUJJs2GHFXbHU8uU8l+1TK9bnp/cxYYM+YhzQmiWYKY
mMY0OQaI+br+tM2b/1svSCK8eefL3S9SsIC16OW7jz50S7gMzdKz9aEAztwdygcZeOfT8x55dMzw
2Y+rfb0qHYQR6KlCXR8o/pWCuA2KsFm5+2UcCLkZ65NCFWshJYxM2P4rYorEQy5EVtm1DkZG+GoD
i5/TuyJUQtni/KcTMUZ+7oAiwtoH3/lRvLPmqbHxvZns6v3+tHuLxBgr5FZOfApceZf13FJP5xKj
EiBr917alPQt4ukkmYP/YeLefoHyzIOeqNnYS1YNqeLLeLCXQCB/kImWqG/zWTGAfTjAEOvCrby5
OsTiW26/Yk9niuIUsQoj1UQYxqr3RbqRXcxvHhBciiyfaBEpNcOIlO6DKh9Etrr5dxP7aSpyT7ta
ja+OvzE+pCQRS7LXZ2TCLhxCI6sifleKkxHjQLtQe1gQKQB8rvrVU4n2xVFCc8VqyJNIb1sq/kHR
AJQ+yH+KH1q2PRr9Se6Fv+v+mAxWN5OyObIqZMZM2WWzzXxS31ZcIlHwprQkh2U1WqbMuH+8cop/
wBIJtTyb4WpB1Q8aRyzyX0thXTGtwbj9MUgXQsJhkhwhWlqbloPWsUHSFWynMIbpO40DqdAkdvvz
b5zuAQBFFp0meerDSA2kRVFMKc93vHx4wSavHOjMtW3se4siCkIJVv6ZXpYtM/rjxyPE687ggG2A
nf6XgdhdLBxmPtv9HoIFMlzGZIUhPQ6bB1zXfjQOScRidWYx4vdBpPb2Rvr+P0Zu1o4il2jo2k1A
xGcwXwkHbGUJQNjy2/CAP4i0wIIQxTNKlS9fOpro/GbbGoVGTiRVc1lb+DMofheXvwhcdtl/n0Gd
ki50mIlM7wvYLxfTCw4B1KhJh4WHiY3OjIrEeu3JxvwyUfmAPlbZ2Ut3eQpQWTphBcT1m2j6TGzU
qWjYuEuaaz2YED6fOqD7zxjVCRPNIFIoLc020cV3R+8nUXcdNlN8kA3/AOqbbYB6rV1Cj0zOCone
Tg9s6cdJ4JcK7Kemxd220Bnv2eReUGtxxcCz9KBIU4EaZrt9P/ZukDmCFT+0TEpkXYa2UBMhFpyM
Ij9engnuDUJvXG7ZhMxf3957sqsWMQgZ/F84B5hXUNSUR1/6aG+qtC7dLbzbwwu8/LbsfmlTtdfu
c2D5ekJRT3i6Ql4ezBH+Jh/XObvUvdDoEtk3Xh8osQXkOPrpDM+DEvA0rOKe9boyJZkdGNoAG19V
LPRSvgywk9yMVB6PO+IPz8jwPqA6ONk+0Kp2H4Eq3uzlAS0CST1fe0eAke21513LwkaDVEmyv9+0
vCtUyzQ3is1tW5BJhuckaL4JiKEzB+/a/bVOZFSRroKD/KAEY0Sw0L4QVBzLQnY8ga6QODLbNm4k
UFnmVjflsl6piJjB6IK+aICiN47uRNT2LSlAKE/9/Yb7sae+YzzQIbJ8VWMsUWEgjDOTDTwy7+eX
xCaO50aSYda8zn6xtJzv4nV24avNcz00mh5ExZYN4alz/re2Pl1y0JCAyylONV4Ll43uG1tOAWt7
jdRy96BbhOYE9fg9EwAzCR773vXP3g8Hf/VWf35C+WzDy5YDQg4kaYOwHrVlno40pN7+aILPdb3U
CE+x6F/itvA9YWR+gUXtvf985C3R5sxS5YeFDGWyVTedF1hSuwtdjCkjoQqcgTi8zKlQCChW9RLL
8ElQ1TohqcRL+1C6LVr8NA4ihEL1MdokZMfla2qn2lX7RLVRRH98RURXOvLwrfQTqvRtJKhdDLLf
uL/Y6WpWhpTczHJnU46/CabTDookbegFiZSUmFFnTQH2+qUUAAtYyauOM6eAmzBWepaYQmQEppc/
W9zX9TJASSa2wwAZd5Ej05rfY7aJTWf8piEvNlZV/uCDH2iGAzRpTVZD3QnjiwCuMbbRFUqGyuBF
XOJN65OWha+o7VwjxJFTUlhTcJXmm0/8+zeN4u8V9krSXNIhz07M8XHccOVN6pOcSoke252iRvCk
qW8NuV2CieEFNdIVQTVgd5GLTTlj/1DiftyjL4G/d5HsY5JVM8VDMcOm2Gxsz21Xu3abJjUjyfIa
D0bKfluwlSR8eQ/zqTObq4iqz/Nm6oKGSRnqt3jmawbS1t3ofrg3BZZrl1C9ftlEGvgRoc+0yyON
18Y3pbG33mfB+RfNsPmKBWfoi2JDqSg9jt+/koVo8MoLeC5ZWi5VQt/3cJNCMIOMEzHBj7No7RIL
v8LZLSIVLYGJdAb7/3prBOv3DrdtZggRh0+fddddaAY/nKTD317dLHpL5+iVBoYkgVGLmnAjAvWJ
bDmIYMS0dvcuaBr2K3ySeuIyzy6kd7WqBfpwG+6YwWHbEmwealrFHZU+7bHVjiCT4+zt5J5rZTxw
ZFF+HZ+2SU3DUzO+ho55coRUSgx7PysHtBhrG8occb7bAf9uwS+QnBZltZw+FJXSmcQS2DX4G34U
1n40cr/DNNXekOUHhLsySNfM5jxL2QSnD0ddP5dj1gGrQas/e1BxRosGp1SMiA56jsyrFzBK5I+s
naWJNE62ZRPx+xpWyfITh8nBUHpMbNG5tb0/nLhulGgdoqqx6CsX8A/stbewkw7wsKGU8a6dkYNC
P0JSko+dsdq8q9ocHAycMVBV0t9qH5bEc4jI+lr4F0Y/QWi90IkMKe4XG+YN0D2BW7wh3BxJ64ck
SYmlJIeojEuGHtRC0jfBnyd/vceWZunvOPsW8FSDYvG6z+263OVLvs6OvMsL/iwMbh2mEYWFyCEJ
Hn5cUkJ+NeRlP6uxzX4KgHh+yyPtybxXak7TdSa3QUzYopogmRb1riKN0KWiScHA7ZUjB0VrDuf6
F/EAHa2SVcgoZn9ms+CDQeA3unGkJWdiA2HQL47P2RY2m00nDGJdD9ZTEV8862fmJ+3X5fCKTyC5
vxCHZdvIVs+13pUQPTDlqjNlsDrndFbmexrf/IN1/h4ePgLPxGqbC2d+aaNtgmpiGn+uCXHECrSn
eRqu0AYvBXK8YZqW+eLGLDbLmca1oRmQO5Dqs1V+EDYjw6+1lYDlpuFFlVEuBoWEcTikDJgW1MD7
offhDQ0p1TEAVn1sQhtzmgiIlUMF6uY+g9ATWbwtRTHPK8S+zocOc5NbhhbQqnH4x+HwWSsHJQsI
ScJLnpqH6yP+NTss6CvgQrOa0nlXLeaj7vBWqCDGB02SjGPJd5g70TNyc9IKxWwtRl1Uj0p9zMA+
lBGWWlT/tKnkmw7OyCd3zvvyivlag3K1CiujJXgy6KS0OewgyEWElvo7slDKjqL/MPC51sWufiSF
dBioTdHjis4Iii4hbWoNQeJl9iHKSYZH5Fsu7y9+7Uaugoc/A5Qv0JlnVhpiSjoLdl+ZI4g7xzTp
xtolcxq1sRwsVZQZy2OI0qr5CONmjoQd4qJZ8ifqoqlLJvDHgjK/wqCBpdFkqdqGsdj6SX5nnUJm
l98D2sNjAc7m33UryyzZ8G4nRmr3VHrH45+e9PXjAILp9f4z8ksCTu4dhmYQf6f/bMh6+EIQJOnM
2nMMG0z4QHHrf4RxSlXHzN+lFeeXjnpcoeOQ4IlLU5dwqrByR/KBbKih1R20IZ2pjOXEdEoc/QbF
CsiWVmBNL9wnlXbjUpSimIgkGsRzwmwjLmrlTfPTbCfKa1iv2hFzDRnYwC0x0OwzF2jmm5KHAyR1
M7sBOz4cG0Cg3zemrXtbRyEbKX1kArKNJiFVNvqfsB7YXAqpgav/n9PyNKx63sMHaAFIstc+vuF6
V+LPud++32WP+YA+hy0SRAuNzwzV27QMiCYyROxhl1JCCfhaZMmQDUZ4WCJBIv7SJPXqEZdoXhtp
KW5gKe1xDnhEQU4AktP2zwRA9El4PnzxpUlsKHR79UbpbmpmBjl/9YPhaVK8ryIsorO1fbNc/6fd
CBfrU4+xv8S5a3a7W5z5VaIWxk1RLcK+tQCI/wXag44C3Gr5eWtLgLdhJUy6HDrF3pkCVXJUbFMI
teNM1vETcuAi0igom8fn83rFssKKtnVcBkO/AcCphZwBhujiG/Cg2XKDDy2djhkOrYXPDqxv8kyI
T8SNiDS2Uf8fL4VjVKWTWvws7cHEoC5S1EHeaOUR/i/qezWOlwLhV+ZN/IPQKnM22zufURlAxAZm
5yZmvquZSKPkpofxo3f27UBQr6l+OwOBjRPPHp+71P6k0ABQ0XysZMKm5m4356R2yE1I5YY9c5XE
RX5dFWH//q5PQEYwBqCX4LgdwqG4pHPMGUw4KhESHzAE1JInbnxzUIa3PWM60GIyRVKfE3Z1AwrE
Fr3AaZl3bmmkeJ4+10f6iyhlYjUumsPaQdKDQUaiYdqCaCSKJsTvnzXS4VxkTm7BOCmbtli3RoYF
BOWZYHfOLh333e+q+IlDBaCMXL+9qQ5Ipww5UP4+pAgsaE3oFieXuVe+kONJ2rRKUmnJLH5Qa7L9
mMPkjlFpYsS4HE5ByBr2ftKjhq961Xv6V6w/tBO9vujkQrIZDPbMqljk71nwg5QfdefFY1aS/peZ
zK4CVqorl/DR8c3Xms2MsmXMgkNRVICxPK/IpqjpqsTT6qBqY1Tvm/0xXLErX0mudQHc+LrHcxX2
04v/pwtPY9B5fQ3dfqHWqNUkKGvg8e9UJmRQwkpZ+KL8rdpnj5Ear4ISMfHuS/qlpQBa3Sg8fTuN
m0o/vayT3tJCuZsBF5Dar+l/jh8naMfciOVl/QIVZzke84bhpzEpiMj5mS100SA9/5flSBHXcN1M
q5EjRXWMixyzdEHRSih0cFvbXgruckLqKeHW9ENarflAwSs3kLn5G5lj6kytEYI34vfBI9kUm0Tj
qj69sLa7ymOXh6Jh4bmHthiP4DPIPubqgMmsO9sbgPNhJuB+kZiIQk61L9fIdryq/lYIEjr9oT/r
nKbohO5y+x9WMRw9AawxT03A1BaToKx803LCpjt6b7y8EBH5RYELir5lgPeB3tOViWz89oQH8D9C
LZuDoj+MMBBzikRcY1VGC0n4VPPOaVADz73W6k5cDItGsNm6mbgBllqysxEdKIq/8ggzmPZyoOhg
/k+T2JIsFTkG/p42EF6IHn7uRBX+kMqVwrtxbnPO0o1juYoLUphS49Sa3TAwMbBYpHcKtl8sUZte
OjRM52ZrUrqf8+pPUXZ8xMVaCb/fMgPSv9WkEhXyLJYkltVsdFhqFsEkd0tLR3UvjmnR4zMAjlmc
W1ympPlMdwzAJqR2neWcqCb53prJ4tLhfOMh+39QYoIOqA7qQSCRDSRb5bSxcfN0kS8ZlWtXIH2l
sgN4xrXZNBzgMcVbsfBpQ6KNF2e70AaTQumDwqjMEz/7lIATUZkOGnhbO7WMYDaMFUxCYzfPesin
kq8NJUhWFC1AQwtRpm17jqb2ROQCrd5d+ipciupR7KYbPcefokoOWJN9TFKx9s/0OzbHEgY+KpSN
dGEjfnP5v8/axiKmut+F4R/52F0VH9FDgA4rYoWq3Wz7wU7kHCrtNuH7euxxOoGAb9QNeiRnS90s
FDdR2vv9CuC7FH5Gw0wweK1Pq3opDpd+euV70ZCGlMXpXvLkVvhtE6HbG6iJXbuUPDLduj5cwdzA
Tp4Ff/Zl23wI1ktv2sM5scYGbmuCT4EWVebSC3JJSPDNoQMH/ugDbTrl8MzG9/GPuy3ivH2tY4ul
aoMpQ87pi53+6xPELoMx+wGQw2dV3pnMwCRlr34XRtRls9pTCXfPUm0K1HqPuo1aZnmoDOq7ou+B
QSAaL4a603IBobIHikgwXmtwvPm8T6XEKu8urN4B4Gl5+wj5a3l3spLZtxvQjGe/F97rdueMdjvW
3bhpMWPVDm1DC8/J/zfMVmHT/cqxnXdBCHnpgwJfTsBNl82O6uoYZs4BJPqs9GPcPrgZ3BgJ5yBv
WCwiJKGdmEhKVfCHxmio2BX0+cEtKd7r2WNetT5o3hLZYrGDnmvfBzn0sS3ZTHo5AVNH0ofBfKjP
Z3B+QYYw098njZODFBUbzYNDCTi09BAKY1lptbrV0FeKX4nBj921AR3H2cVwTzDyhEyo3FQ+8ZHm
5kSfh9akja8539ydQigy+B3mWeE8f9XyiIYmYYgFxdk7p2KBrSd41KzskV6wrEYIC35y6vBmBr8z
h/oEWtknWZvHA87QymtsQ6eEXkJxnI4nKJVk3K/6LVN0OcUgOinf4GAJpc/hnrkOdwOj0oNA69jO
nFTxhExzrteK5Zfx4uRG9SZsAP4Y/2kKnPHxfpFxN50qlyAMTV445yz7Mgc/cJHZAAl86FTPBKVz
UyNCckhuPgUybao2BG+YkpYju4dCox0GbDMEpIzzaE+dlZOJUDCfLWtlYQHF/MU/QLnw2tCkUexU
dJm9GAyXrYwMfrgAQFZqk9d6zzTyCvymYXZlmJJFjnEuWJse41btfTiZUHlE2TbIgLfcFiGfyZG5
LkegDxbUs6lzPLsJ2RQz4vqKOjzoIjHjwFfvR1yAUKWMJXvlLmNdOg9RcX9ktIuIxBy4fpcEgfbv
hLRs2SEURkq1J8oCotqmFBsTzGZX+/GmlEHghGhYV6nGvB5nLEoZTbNUe2anIBmwUOlCdJlcto60
ZLkFO1DlLwZeEoGQpO+V10SlVEtNt4V25lwqWHx6x2pisMbd4Bk+5foYWqqUuw0rBn/dY8q4pR/R
Z2EUoSlMYKpjBykRj9JZSF2wkgszkyHpTZEhQA2qpDi8kN53+M0L6Yx2zrJB06yIRkHGOLXd67eH
Vs0CsWm7rgOI3S8LKvJymJO9dDVGv3nR+MaKl3qrkVhDm7z69mPitASpUBFRej53TLUERosscq25
gDlGQoQT6DkzyakI1+a2zuE5lT+uWC/jZoVNG6ORtAu9y2zEOxxC9OqRLVPosF3qDpdtmkJeXmP3
T3LSv7MwHSeo1tqASs7oyr41H6MUcA1rIHMn6F3Z2C3Xe6XBhRHUrfYQcqRO/I79+CnlXmoRzt6G
AukS8Sjcf5iAe+yKWM4s0bK4Qv+JCnbBv6w8ghpDvfGaw7Zi0uSmkhoZ4SQ2+5c6LpvTMOKxT4ne
zhha5gHsTMefYGYa093IjAuxqu8VHRPFLjtY9CtKT1WwRJU0c0ftuYjEFDbIojx6T/wCdAgOt+9r
LHWqnrG+QDxdp9TqQ5J1k7MPD3NNE6qsTGwdq5vsAi521M6Rcuu0a01j0VENJvIDRsBiNsfnZeHv
Bu4pGWWn0eci5+S2toWQwQljQtusvWiSBa62Xh85aib/PTyu77InkHDrW2/aNTqUiJjRQmsMwFTr
lP+R5UM7ZVm5KftkCzQqMhDuzzm0PgOm1NLgwzxSd7U/2hmvFiefKmyxLIRVY+tizuRiykjsYR3c
2dCG2JTB+eoMqyPCTiW6V4b856BcgL0eVZkXjEJqI48JhegKqB8ubUGusLriD8al8bTXWn+elgAx
VodSf6hn3MssQeSoJh61QG4C84zxllMKhCKQC3sG+cfOM+5xPTWlRo/sA7QGeGkY1yRZbglpdIFx
Yxs15zfeiatPLrc5v+jjrso8j5gkjBTEPKywKtG/rlwZmEiRermBA2EqfZjVrpcMevZuOHeCQ7uP
qI+mWR15Ynao1Yx1vfaWWJjnfni6DSbiqXbxgk+Og2TBrOnfw9e1gxfuQoJcwPrfwSvQrb9uOj1N
7ja6s5KDHgA311CvgUk+TY4Lr6ccxwSGpUbfcyGF/YSmcNB8r6SE1Dwb780YiSFtHkBtCTJHdCkY
ghaS7YtHjvG4u0cp5KTt9rXOt7IK12727KC4KC8JK0ovKSELZMOseUKINyoZmjRkcX5YOKBAW30n
dnzKVNCazMkvyISLVhaQsfKNMovUeR8Uvq0W4jHRQ375zVtiBM2xfsZQI1u8fKtBEcI/cZXyOhAf
l93RQ+MyX/M19JNbBQPdgcsXIbiIV10j3Hc5saYd5jHbspAFXcc+NVIAJ2L94tr4nSNLMa6iKhVK
+4wjwEjEcyaUjwISIw+uvP5CeATyXXX/6VVSB6RY8czsREh0mTdz3c5hu1uhg8T7SmjlBQNcXc76
sEziTgAIN05iH7rNd8Z12LImQVS1PTGEBxFTmnNFyaQhgciI3ZoHoYuYTraRmX6YHR0JnWNHkh29
6qacRHQUpwgM0wuUXDH0+BuOBOC4X8CqU60fw706Z+jh2++JwlP9cVtDxpVEBNWBnrtzYS+gCoMP
4XBrcrkytRNUed9uo6RPccBqdq9weDwhfkBkFbm1dLzmg08FrLWQmwxaNT72TNZTmafnbOVqLNmt
FJTsVv6d5du+ZK6xK39xzFuwN3qHHhA3aL/hC5NFS5nE5jkrl3dmoWwB6YuIP4Ku6+zmhY8yrAWT
vydAfPuHmifXMvxa7mqt6VDllag03NrwVeVLVeWwV7kNDGnMVp2G49ifIdeAKm0E5MuX/ksvqf31
1oXZL8nARqT9i/nWCIIaUhrvpIzvYdYAHMq/Mp2SVU5vZ7H7WPKPknjFzZowarXDf/I9EY9OXn6o
VGaRWsQG72c6ZOypzNu5s3Rkt15g/6GbHp76iWUxKJo+ljItMzMIwDxOtoAAxUEGfBYHw9bwclFQ
1dwdOYjno3y/J+415xjPF07SnR2LaHgXBxtmcbQaD/2nOroFYIx5cIntBsp1lUOyzolhffaZf9Cq
HA6LL/hqfpYf2rY5xnWlMHQPJ9bJbmmU/k3IIKgw58lGkHugNKMzdWOrnaJjbrVVazKLUa17RRxL
DnyOqieXYiDKwfOCGDh3U5+cosHm1KSH9HMr5RLbitY882GsEhYUCo3M6cSavpaGpAWsmBneqvgB
qmR00m8Lv5MUflcnZUTwvXlLrbMsfJjs/D6+yaGwx835aq7yrc1MHWlvUE9nuHqhSPKOyVmzis0b
MrA1lDO5gqY4ze1L99oE+7D8zQFdhItcvCI9sYq4+p8t+3vI4yRROldc0Gkke+fEghr9ccwl6ODC
OgKgtWOcM57Wh3/qYo3AgdrGK0/9eTMXfqVojXzecETOLq3j+Q0P/UC1yPQoPUSCAFyU7I+NfiHQ
IEwKR2sNXiimGcPmKdY5lGalHgFcwZYRP3aB1d9cV29d7oKD3yU0C1LIN+wwz4y8S5oZQMyV4OJ7
2R0Hls2WZ8ET2cMQbgtJ+FJAZP3dURohF4X/RFDdOkaRKESf6kca3NEBe8SvIf/DMXD4LLByOnDh
+ArwD5rF6UMkUMffV3VX/UlDD5xASe57dtYl4crauD9tjnIrTKB9FK1N7AP8pgGlWalluqBBtlv+
PixeRPz4jh+acWpeDalG61ikJxq+IjH9/o3Txxm4pzx9MIMJVl/EfqfhgOKE4HSY1aGnE1QBQ6FF
OavUcKvzheoAbQGjcEoC7ufRy0GfLCreHSZE3nLgBS/dKssm0gAmdo1CVnw5YBin8CBGQ2v3pumi
9rlfVHSY0K1tlmoQEWONgQ2bsZ8/3UyOhP6D965sB1rIAhL56V1fAq5+MsGVQdbv41nvhhXF/daF
7MhZB30+DuaRNkF3tSxyetmHCSLc1uUK/Gna+dVIFOohyvD/yuu1M3loUU9snvmNjEi3DITewgQx
5sNUifBhMg9o1MHiU/CU75NnM9pIJEhrBqrFnDBdCHIbGOc1aejL29QoRnT48slJG/mf0QUTTBwf
qS0rm3Z9UfA6VVoWiSqCBVqT1/F/yoUm+lXlMyklHSFDNUUUUD0+sMZOY8gIefskOsjgF/8CPSzz
uwaiqy8jcgJu0wmR8MPRJZMYHtuCBJjisA4eQTxhx/Z45pnn4wLkg0IFvHWy5BgiIg1xyUJ+twZs
6mmE9Z6rV32p0eHqM+GbRCrYGF3ioYg7im+fUas3omGmEHEsz5732btjJ8Ct5gK7Dys/MMgdebuU
ukSns7vyBaOcIy5wemOHrzBVywAoweni0xR3j+I4hQfniRh4ZwK02rUQ4aI6iEI0hYglsk1CXGu5
OhFbaEIZN/1q3rkKGk6nJoEIxsQePpfh2EBiePOSwgQ7zpfEgYdOohEOEmbvoXtbyateAHtml23O
AH3KSAoQAxR+75OeTbnle1LCS4L3etPPElbPSNGDMdbmcdriGp5uMQvWQQvEB8zL2ZRShLpONlum
DVva97WWQJ4pvY4hY/lkbeoyZRu+FvXEk3qQic4yPU4zKTNrW1eODLss8j+TmtGhEDJ8oZ8KOEj5
PI7kWTSr3nLd/kvYmreXm8PJcymnjvPvrBczyRa2hjQ6fA88PWncohYkctzvtxOPF07XtjIfODea
BdoxLvZ1ztSM5cVwUtG2cCZuNIDhbJskxzVNcvU6lmkqA6r7TKMDd99sm067llYLro9fMnBEv0a6
oNTsR0movhn6VmYFdCn3sf7TqM376WjmBbdNZI4tPwJ3WheFo7Ia7pFCgsks2VDRA/yDCN9FOFBn
TevjyreaHoY4ebCiBhNxK2qU26lB5T01/ZbvOEW+ZyjDMD/y3DWIQ2b3FmjxqnfGgkz218P5FmDl
RuaCeC5AXr2uzlD+dL6hNhSpQdXKrPKYtHAh9PgxFObv8d5LS7vFCTUrBA48YH0T2PEmEGNB8oRi
ZnklCVasCWbqt0SH9rJyaECkfcUNHoJ7uicQO/dsYKTkM5rYVT7maMcV/oMBLub5/p4hvB9R66ga
4LPysjjh/ZWRUin0HBEtVXkLNctEa/kucdj+cn4+4x0aIvJZTSinDoBZlVCkt1C/bO2+imx9t5Vv
RauALtAXynQNuF9IQEamvf9+tBspjuExzQkO/pe4S5j34iJJg2Kyojp6iCCKPglmkRf2KHlUdnvO
aWfHjSjH/2wONsVkjvIBsMSuMAdkmrIdSmavfAsRtxphkAmlpfknv55SxKRGwVC63niNKCWF/8DV
Q9m9Hlz4SyjpQoV4cF1t14oQIT3Yy6rjeYGSY29bJ3irMCMXIIKO4IBkj6TRrAWk/HkHuihbF13s
zkQvL4mxpQZn+nBrGKYOv05DM13Ixs8d5RqdVwFysgoM0iBJVwy9XtBkhNpoHlQEIQpxtjM6wzYE
roYnfaEGOI+lsd3lEnm2DcfIb4GvzKYfrcyk29o64oBGW/B/zKC1PXixZDscJp0aOM+wjJ7mDnKh
6KaCqubh+RVSTdAnHwFSrFxoZEFYHJWvhIK8iOS/oheGUKHROjFP5Posbyfg7x4lT0Vjpk8e+mUy
XxvmgvfmmuHQV+VxttXfO3gSkb/c7J7sqpYfjbuViP94tKxhMH1sSpMyo1HI2IwOuvwlR3ECHNAL
2UDnG1agtrAhVOdZzpV7CZn1R+hcoUI+UM/fbhBvtw/ryvku/6LCt2jKPbmNEZ5/L66mrZy+HkcN
/hauwy5z0iC2+VkFdHwEMzPRbJDqZR6o7uGg2fyW9bg08rtZbaleRbq+rnEsk6yZgfik+oF06rTN
Fys5zms1yI31D3PJS3wTZdoZ9eRd4U4oLBxzN+nk7/n8PRrr1Zs9qkJq7mTnqIH92bZ9Llwqrfke
kPcAE4TaLOLHguwflR3wKoL4ZLPbt1g/B3rhp91S+dT2RZ5H/HtM7uq7DbAQkgw6DxK24W15fnoE
LhpP8JBtwYFWFe5V+iNz+40yuQxUp7+JR6Tx3oyHr1iU6eACThRzd/10kVgwQHVboKLkO/H53vhi
slbUBRmfuuenwv2yHOcytM0j4LhvljghrtOWwYCEb70dab9begMYgHygsC57uBPgKESmqZNS9vZj
OYF8pWoMm/Y4G4ytJz4hurr5hxOLOYjUsHb8mtoXfa0CQLjpQ5SAttHh/yqPjq2sbxe1XkXyBFkY
M3X5aiCVqyMFa8B4I7dM32FrntpzhfWwtbX7Q/Fddg4TgROjJAWnxydip0y66PE3jms+8vFX71uu
ycDYbWrtbYcCEmrHr+iltWZdYVNJtg5oKoqkCr/ZqXZV6ApFtGXU3aHm80ht9OvsTW07lN+Jt5rE
xqZvFB3QzBYIRDIub2iY1YXGMgM2xMfIVTCmUuBgLxDo3NkRAjPDw47RAGTEqR9d9M93mlM67gXX
WDy7mSxvmHtPZQ05A9iOzj2Ur0TqYjJW2mJ/j+Mj+KwIgnbqg1wDJKm6x24WnvfOgcC/qfsodjoD
8FEr+TQi0HsSpcFk7mRrYvzo9LIp0XDg42zdcLCJLGgpACbLbWbFLL4sHYxVtcCvHw/+xLR4S/kl
dJSpwXiNXqFjY8hVhYHBKjIfFQBIiHAobIpite2lNtREBeuBC9sKUCHT9gu6UgAfjge1TOfcIv+o
d04a2ACRJmkBY9ZmwQ06Q6jCRDzQdlfoo2AL+hVVrKSdf+A0XS2yZE1q/SkEcXpbmKwb5qEsPKW+
LJToDWpfLn6FYnkcxzYo3x82AnO5NpJaXZyNP7WcGWTxOkdu5hcDU3Thzqejzt3Le5EUZ4BipmtH
kBR7oS+TXnrIvp7ETG+mmN9ZR32hqvCwwG6NapeIXxIaSjcPrqDlYZvBsjwjeorOKwL2jQ/AA+Gh
nB2+0iAVX6BcY3W0ge99JL0pah93zqp+RonrrFqK0OsPHk6ByV+xIrLjg+SFuBGVyy8H4BmAK0bg
QkWx/zx1Ag3XHxqFvvEYnJi1GIjKbh5jCvG6wuGsjzIX56awi6nmX1ncDBREYH+k/X/LrhvK3HhC
O7N7HXiuz4pKxvsUaySOP2VvJQ+J88pDjOwnJzGyEDCNX2lXlKwQxgW3Sg27VM332UNOyEkds/6+
u49VGa2urnvOqiBy9QNguOQx1SHnf4ww9GBmaJ/Cfz50AM94UUHnGIqFS0plCgov3lcICgDc7sV7
jIcICd4VRamGtpX1veAE2x4G2kz96lRUFaIGMhNRWAV0sXlrKLsDjUivBnkDKsxQsYfk0e6Q8XR8
9v7On8fVdyQugZJFXv/jZpxZytLGCD/rE4tXjjxvgwT1zroyVigH8vuLMHvLdF6ZLeK0Tf7yj96r
bWXW8eg79ZjCT6cLOgEwUR3hPadDk4HQ0RQ83Oc83au6OHKXLiiPVcBvM0RnrtzDO2GNiJmJWKEq
PNZTiXQQNViVaN0M0J86GcIsvrI2YejVToyf9q+yAWfiBmLGzSoyVKBV6X5/rwBle+TPmrF6FW+b
GEjrYszW7UOcBa8xs9banMtCUm6SNULFURRE8m4hpMN9GUHFaqWxJo+Xp/plkyX4we1cpVn43KW3
x6wo+jotLUgpY+IbbNOLW2wDeEBKKEV3SBBL2+1n06l4TmzwY/XKmkgbyjwYHxe3bq6UhC9fG2Lm
rRNY0neIJZfLqfbd7QNrpwFdTc59WoKXHq/T9hYKA3QUrARQDlEALu+ASVG6A4KYB0eSAFfCA2Gb
OLUDL1mj838jJW/QnyOaAkmhlU9NO9N74tzEd44jrIohSM5mnvBsb00WiRYTEmh+/T59A9vbut86
ti4HdDewx1A+T2JELRGMfkoqy4g+ZlhVyuEvgAodBDSLHaEvFKFTcc2sB0P8xRlWJ8Q8TWYociiL
OV4jLTEfIw/smzU/Wp0SI4zgTvAGuOuPRSxkJuqmvsdS5tvvLTyv8jkDdkGJATOwSx2RbJJyqJr8
cR9ji51PfeUkPBofSbYYdxGfEDy8FOLG4E5wc+gwhq6UggZnsCD7+g6BRx22tCeIMbd8PxWpiykS
knhGJk3dgAhBBRNyll0YbVJTGeKy308ZkTRW9TrNbqCQ6jzzhxlqfzdVFflEvHmxaybZCT1y0L/P
J7tTQqtx7424iTp4s+5cYeEHEO79hIoNnuk3hCRFMWTF7CKhMb8IDj6efgCf72EbCbJcLCHKUApz
18WKG2ppG3MvDztxhjjEtpdBZ+66OaohcKBK4q8xWdW/5xiRudnroRqCXNalAGFjDxpKW5HiVgJd
bTDaaByzAPVjpBCfF3GP8j2dZquj/K6hqWNDwDYOd7vy41B+LrZ3WgDc4WWJtGbINqyhhNNVSXtk
j9T33YSuPpmsdgDiFWU93lKGn4iElx3m858D7rpG2SqRV4e7i3TQCSAOoyLKt4kxwHHIZsHSNafV
ET4ZJgYOYsuHPkanG0LbW7Q0cmz0Q2mUB8Q4ww4UYgQ6N+DDwAtv1Oh8smePqIR2lVGkjLqD2BOo
zWjLWJBMae/97f8S5caCElyH9n2Tr3lf10VLZcRJjVWj0HAMJo/c0C8HUqshB/fBO/gPqUkLiyny
vlxC8lVyvLJagW1f4TOqW0aLrLGW1BQnDxtsyd01y+HvwpNbGCcP179FCCjryMloRRbkZW91pRt5
2h22cHlbf+5w8aZbnsltNhbadWXpihXKqLNwrgFxirX2yhi5gYwK9GYWjCXSidFJen5LqkLd5UVw
iVVw1WDJzJcWzFQ1XcvU6kb+GuD4lXIN/1ZDxTTwlNoVoRhhnZ6AVMMLRvr3yEd33Jb+zbCQ4MO0
jtq1gK6s3z6VoF3idGqlNN3euStPhWaca16OsH6Mj1O0ynurKg0MJds1H8RUrnb1aTE2CLQpM1j+
pKkJqyOLaVcbJP1O4K75kzmwjmEGVYoa3rO6KG8A8m5IVyBLqq1YxEjRrOLndV+rgQ4n9HMNI+jW
IInFuttBw07R/ZhQfo1ys1CM+8BU36FGWN8XOqF3ybA/T0PzgArMIBqlIOqb32g9r2U3pskShima
YLr8aKwJHyLTJVBsdxaWxrMY0qWvAikSACN3BbOeh4V/qRjpH/YH/T8xk8k8f/iTAzvx1E+ainiw
4ZbV6+iuYLvziOBQSUySCwCHBqSi4a9vAXNxUz4fsHGGsSGUvLx0K0x/jOBysqItEdM1Ueb8i0/O
UL8/urtUW8XlKizh4wt9kXiy/s7uwloM+VV+YAF/oSyrzkd/gPiQb3QnGJp+g2un6ZyT7r0+ly30
LZINvACpwKjNF1FNkYi1XM1a4+ejePCc4MPFenayLeNCGssl23wXzVWEEfXdvJG0q6q2dl0vHQKj
AKqlgEkh3RbYkSaTw9tj+2xU2J3fRtHlVSON9cV4hyLX9wfcMXeXvTvmDjCem3QaKNetlhNRa2nx
OaYOOP8iE3qmnn1bRVDueGOFqrlIOp5UaD4nZpsBQNJcWcN+znNZOS9t1JNf5CP3Krh50HUeR7o9
W1tgzcgqz1J314SH+eKnsLefGa9CAL/WIm/ePJfxGfSa6+jNdrsHUAXJ0vqqAZLWAiTGBEaQ05gP
je+U/FOGkliYbw7BjT+kBmBPlMS84SrIfqutE7qy1H6FaPcZZodY09iTBOHMxh/s1MqQ1kOo6S61
GupYasQtOSFcKCZejM5Wre84auZzXVOsVALKBqeIso5WhyHpO0DbBUCFM4KwB9hKmhnJZpI0cc5D
WDjVWorExzsrdLX/WZbDLeL8LDdRMymRSHdVoAM/7JeDQ2FB9N39pICOPonK94NrOikvp4C9mva6
StNrS4nMGlFhrTfcUWx2cEMoR1ZoJAPlRHJec1ulApX4UnDuhiTaimzhClfG8aSJzd0DzrMvZhtq
i/5ohMl4Q4B8f5+aY6wG1wpSRPHSIIlRfMCVapkg9VgC1D4EtAMquum2ouMRJT/qFGVFgUyJCZL1
N3TBFGveHf3zThjxXW3GkFJpuznr6k5ipM1JFuLasbGr7Fhle7ABDbILmjQJjTDz72hBjgOaTG4I
4GkAz+4aNY0k26KXPMvCVqbCWR7Ia+36qUwyi4h0o+3f2NFhDuv3sFcAO/wXmOZ+abclR31kM0c2
2rKYGUxaKMdRELkPd4gfoBsFB12MQBbc1CvyTqF7ZVrfXY/1pzc4GaRhy1pgu7c9amdzV4QSY3bX
WxOeu6vr3v9p6jXXZw2aLBhdv50LAQDctO0BrfId3BtGUURjSqxWOowH7emiziqdjcMqcQcAUPLA
+rIP9xB7wXkUoAWtmxLazTF7168Lw93WoK/tFjvnQ42yWc3QkttcmwNkUtz+5WfAeI5l3LaTbIPM
pyV3C6FxtMeeRQkE1zXCqraALyFiXLimdUO0gMd991GyK5uSftYsdNgUIFF+hlEMvtma64czIaSg
VjZk+En3N+mTyo5gjU7P7PoQ7/pJxSaaH5LuMQQBH70T52HRVbbUNZyfx4WMuP90C3sYy7x2ThpR
stZxMHkFGtTDzabeNCX9TkQJCDS2f9eszUMtb/07nNWQOMZz3WcLlxoEJqiX2KNYyd3FK8S2knJQ
cEVLpKy9D43AxoNxuI4xIn2xufK/duG1sjIRrRCVOdmA9VskQRhJbwoecSCn6CpsoxN+RAYzRMFf
BU/JFyM3Aym9Annak9QgRjpurm11bp2NokUN+2eUyNNo9m3a6tsVpWqu8CkPkZOgmg+ZBkzjVpbj
2qasb0f/FV4p42+MhB0HnGI2v4ZOuM2wayfOkE1Pe6usQI/1+GEVjbyAQHCg8mAkLPZ6o/jWzWVY
ffNp0S1PRAAuasEMyRVu2bVRacdcg4896IYG9ObllLpmK3ZfTaWlC4dxTGfMrC+OIWpkSHY0Ebsd
vFek/IGnLW40klehkK+/07k2NOZcpsoEVG/fIyszwpwGGi6ejVBtOVs7F8MlFLGkRyB5rQDgVEp0
qxAkvyh0uaPw3Osw754TO4nBZLieBFHxIvP18xhptu1OZby2dxk2KUJihPh8EM1lPo+bzfq4w+GS
xAqiNl3XMsMMo64Xd4nUxe2JqidtWZF2GgE5IN/r6eeTxITGts7t5hSASdJG5uqOZ8j6UXnl28rF
aazDj1Ow5ghJ8NZI5QxqSJFPZdyNafK28tEhV3XA+Vyv2e07y22AFuVB47pJ/ftxGlazzb2m1JEI
dlokcXIKHWWgYpD94nAnYHol/aikfK3o9p+++50xbSwOdMcUryPlRYjl1NflKq7wdyyix4LOUpX7
gXTOCN1Qq1FFsBLPU4RSzOnd79UIIDCmyoC6ZVnV27mEGT7wnd2OOuKuPJwRnZOS92Lp+yhtABfF
KdETj6ZxIpgdU8Z7jbr2aGykqXmbY+qSgfLqpphRhmmFkhuQI5bEQxRMVqQ2A6tP8a4ITiS+UTE5
k8i6K7CQ9P/PD1dW4IFCg+i7AHBOgbFjGou7lFJOAzYLS66f56x2v/vLdwox6rB56BimQCiPYdrC
9+XmGHezjX8bo6efXKJKy/98XGU7cvSkgiQTBpD1JTSB7lgs1foaQqL94McpF+hVLCtLnPUSzK0J
OBLfU0J0NJuKuv72vr6igE25WsiLkWYOTuCofuAq59fhetVUysQvR9fXR/SZ4pKW2fkfnnLUzVuS
ydtC5Vzje0eYylNlZi17lifLk3mJnTOgYXVzcJe/fL0I0r9GYGu7gE5TEcCw35AcTpkICACeFGWI
zFX4fbiOMRfCkochBrGdCjoTACBI5X4+zOgT982wydRUMiHNuizHMBgBbj/HqGlBx7M2vqiKKmpd
Zbr3WFuJinvP8wuadK8g12LvHssjClT2ESkx8YPTUFNmITdA/xqdVGJvbPgSkvblSNB5IORKHZUg
5GY1pS6z74DeFDoMpQSqojDVfHq6D8jqIox3A7ouZoEK3elT8C7/UJVdKXOgBZPrmAw4jPCSjBe6
3+4cBjP3ELk5QNLa0WCkvLqyciFbPbk/omTeKungxTt2s0Ry4Utn0+JV50ZgkoA3C/bh/csQfuXS
3F26f3jVuZQp5Zv3PWfEcdjfPcq+wGhFogBdSAb+JqrejsuGlsN1Me3GZkVNpgMyZrwWyQC27dcK
eNcjDGouiLo9TGtZxgbARBnLI/CEgrkJH75lXsFIOf7v6uNXzABN6dt+IOoXD5fC0okGwAhJqYJ0
CtToQO7jWGm7MxMYRlCQC52TOPv8WRCx8ACL/dwmbXh8qhj5vRRdQ/dUL/PCwyBnVO8QQOxRvePp
oLEccO9hm0ae0ekGJKFeVWb453Qna6ZL5+MgFCuuHJC8FOQRdqKMy51zISkH8rBJy+5PDh7VGo9j
WSKkcLj0IMzmOjDtM6J+hw1rt9KKRZ+8Ga3xhENNxjXQhituL7g4i8HZwB8RRu/x95Y04a/dOXO2
2yeZPlVO6aFteTduWIs3H2UW1/0sdlsqJ5W4utASxj0LQ2KqgziM7goAknQyDHArkLt1JQx5U/L1
g7rB8dTXesg41Sdy0Y8+3wAiwiL7JMHsFsRES6i8IHlEY7oFKC7iw3FWyXEFVNhWO+G7Nj1qE20l
oIe33Blq7l1DobgHX98LYF2VJWYVvIcV7MBoEHKqFFvjzz0zdomCwreGFLbNEZQOilE7sATc3GB6
ftmfa6UftVrJbhfXEnrmXa24VFbNPdjRIMGZwHEMwjZoTgEM4g9UNrmyvNkCsCdaJ+79D/K0TXO+
E/JnaJR8xyxEZUhLhgW1xURGfA27wscf/twJl7/ELjt4NZpVjWahuVLWRUI98qRJ2+2FyEcTcgCl
hzq9a0/SKd/rT/yZXn4h9+TV+KKFQDS8B6K1EwJzAYMI4bMV35YDyyC7bfDj9I1OO8zXpkxxVrn4
1u9CnRr28yCTnDB0ZHzh1hriagr0O1D2RW27f4gtt2MMgV0wtn5UCMKXfmWynyopt/xy3vndrGoU
wEUAHo2+INI+E5E2S4/zQTcGi0GGpbLuDBWi02wR0Y7GlWt3kMkACiHtDIzHjCnhHT5fqo76et4c
SYGGeantUaHIKXbqzmKVv6exLQUsuC3QLr066l61tBKAd0QDau+11MuRANcVjZulEHFL7P8u7/9x
153HcMrJbasOm/Su+BBAV8+KlDvCSCUfVfCZpFoobNQcJWl8kr4tkynq81MED/5+xNFXPvX+u/3e
hv4ujB8zxos8aY5XJ+hB2Uq35liqLmBcRE+4AmkVPvztYsozkRL6pYzlb86aaeMb/ok3JeQ0wfIw
CyId3ZMRx7yH0guV2jVFOBvH1RSl7kq/CujjJh/10+5Vbnda6YWGHeqN6vcYJac8i4Qljcr/py68
yQ/p0/c6JPpdU0B47jQ0RpXxYJ5N9Eqw5lOw49NCtiS6wI60UFLj8UpT4uZoXJFPyk9mbP8BgNov
DxhG69UknazyEC1Aj7d4tU7wX4EOHfbREarHGStRRqb9KQYnRfucZOGV8Y589y6sIKkogDbTvH/P
jSd257qbP76kNJjQeEbRYV1NxdQDKp8eCFadKPyqTRrF52RtOaVNNUjwhm9foRL6PdWPTJjUjhWX
+ATWhsvE0KRsm8FL3fheDHxtxVcTqO5mxrrYLOdTELS70A9072ZzlEBrF58vshQxi0CComO5UpDc
NzK7hve6O54ugEGpTkg2Xm+e3SGWQ4U9wm1SqvGlT9mIk1ns+M6rVKralW9u1LPCIH3KSW8YCxLb
6UWCjIk9MBisrsi69m2OKvYdZpvWdvN4XadhYfuRHNN+gMGPZYYIZYZp5hAfXXWY9GJXCpYdxn7x
7+7QP2BKpZltFFiGCYQNtS4Nvgfi5tVue1v7nOs2ifHhJY/uTlch2dx9x2XCatFah7jW3xqM+GTa
xRwv/vALePCxxFGDGhjhRAnz9NhhB288dB40RurSoBNL9wEE2dk1bDF6aOZZDuoAnciRj05d1Iy7
gd+coy0sp0aWzi6t7+vT2zTzl4fdEJVViUeEcQZrY86+TfPIHnem7TDDkc+iBa1wZmJ0WcaSS9Yp
N/E4gzSbKWnO/Ua7JKxRvZjqFCX3q00huyztOx15ReLaYYpB2ytK+WTAil+SLMDNhnh4eBm05dfo
r0I30hzeOqZGDyKPKjRhtOHqzChFEeOZWz6TVz/dIERDFLVB65hWf4DY4o4CBPwIwnxb1rbIK0yy
oLWDAzNY+DJUPYgl+CQZ3H8Qy1+fcoA5i7J2RSlTc3pV8W68PM7d/mYYN46DDpyHaQxLPr9BPxIe
OajNeiZEPCqi+RmyKQdfI2BkxVr7vCx1KHYtLLUXWn5QsqGHJpDnHq67pk+jTLAGm7EHvzQ1A3zi
7PwV0tNEeu4l3xCTknG1zESDEQ3CACNUxH4mavKz3/NKuQ+C/k+4TvwjDD0INfqjcN5xtlScc70v
UeS8qBf3bxNq+c0rKxJbnoTKMBRqaSIdK8IoDCTCPYncbE7utyAZtfdC7uQtnMRCCeqZ1QvzvR+O
HEsq88HcLQcDkjgUJGx+idlIDEqAl74zPzzvEqTyTf3ShzyjWm/Cr0UEV2ZUUymzw8mzXexvB0Np
GR5NRLhgeMzubmYkUrqG2r08eLK+CkzO8lJYJqWCc+mS+//JmhZmVqrphBjsC5cY6055u1zq4oGN
xy4qC+uawMybh5zucQUgERRpGBXMonKaoZ/0OoPLz4Zt5C1+9nNV4EeRe3K6aUp4xRAz+32GpihC
rCzqSJjIALU8+2gRjGNIFXVIsH60BHdYorDpQmQS4llZwANRqO9oj94A1mFQ5g58c8UHpNy1O2/t
KCIKXgOX46JzC7Cd0ONrrPCQzo7+UAfpwcDM1xWQ5KzZnvxKLu6y5vCfd1fqeVdqD25bMqnPnYDC
k8r63ioYXWUlJt//ftBkx4hISnGT9VxOTpeTDVLldCYmNFcaG0evQPVP5z0WP23++B8leWoIFfFR
luTPtTC6vZEkkinA9SQBPZ0FCkUXDDwt/OXV8iNPX4ONjmPHxIBUcMXKnSmpz7qO+/sRH+3cMocS
4a6hLUUIow1w9Xe/lbF7sQpoXE1MVwsjCWBxS06kVuqph9p8BJkL/ld/DdT0YhCR6ymNIk8j4RI9
ZGEQ/XpgEPVAE3UNzglDQZr0FBoDTdmIxXKslgb8X0FQJpA3ijYetqjY1Y+lnn0c9edWeibos6ta
hqdSERMt3JrUBD8akt0dQvt8iCRX74eGr+DhO2EtI2OzLZgqI2TeSKek0Dz1SWfRyggowu0V8GwQ
m5zbM/cm1Z6cRSGc0Me9Cwj6dMn+fk/xCLrzRM1uMwOvDGrUv7tAkBBcVfd7Frxuzvw8JzpWroAV
DAK8pOLyESo/bT+IY+yYPjlMIKeKrvjoii96tRmRfvIO624jPvL52doZs1tVrM3zCN6NZm2eLB4t
BZ0/l55usiGKwg+kN152em42KoErqoJ8Hl306mVbBNa/+KM0omfjSESndzBexugy7LX5DvYcKGol
z4gjb1m7YB6StbVlZciGzDgH9Lb62Z05D5GEqewtf0iZIEZGVJjqx8ow/MaSoFejE1GcF3XGJ9jl
/DoISxFFpeKdcAup4ARiKt3sSwRTO3Eb3MZW0IkJlXfzelPWHBdAYgCzRzxJFzoAcrj0N6gPSwNs
cYMldxIaZpgQyE7ipy7OEhNKa2/OU0G4mi15CZCwHbMPkA/gzYoSTBxiz0sdqx6njdibN3Ftr53f
d0l2Bdl/0jAIriv/MCzthIhaGBw6hk5DeYghFJYwPEnAEsEzIBTA80duRRjQdUcnLhzKtwRaGDrt
FLc0Te9nCz32K6guSakV4c5XeP3EAeOoFUWZbrSL4IaqsE9GUIJB94ViYGhqjfUDh2Q9N1oqQIrN
RKYQFI1KwsQgM02wgOP0B0L4QibJcjb817v8IQgaf3K/Ecn+zVNaBhADUdRCnUXLwcNybjhop8oX
IHPRQOO2q/Yx/32p0GqoQ/vav6JzIwBlYsf7magkI0q5IGnAjXuAMoH0xh31bvuCjUfEa3mLZWCP
Nmxf296EJx1VjyARg7LL0VPWxM99+DU0Q3elmaoS3WM9cIWIvG0J4E0pEFp9tvzBUmW0thyr2uiv
1uFyMaxzfvhmFWWhTp6ZiohW8Z6Y9q7fjrjrHIH8X9NWtXLqZguacixtWLJLMRqFZSbEe45Pvpd9
FbCp/NxP2bZw9eR5vweH8i5scFAYOx8vP2Mwpqz7DyXSllQUDYSBIkEKHPG/DlWmTISXiHzEsEtU
Fob1oTUfSvfpJGNLHhnDlWQ0U3eygwQcjxvHOR0EtSzfQQnzNojyXfxhSStD4ZZXxtIg5HdYPUUo
6Hnsmrqboi3PHOZ6RTeJXPLGgf/10UHmpjtsyoxSiLDL5QkfpKVAfvqbuUL+4swDsTTum9UNJsaE
FsKKYhtaM6ewuVCB4rkD7T6c0U4DLSXY+KRZAo0rT15LIQq20jEBErOV2vzpxSrKo6pdR3vkFFBU
0YgRT5IrP/4V+38TpkjsQezUbJygDFXUZpt/haiZPtIWgBdp2TenXPWcj7QgmuEe97k6pndPWLQT
0nqaWF8XlXGgFc1SR07T6qNoPeDA+FNGKXzlC9iI6FdtOXmpIgpZUQxx4IjU53vA/dijmfwF28pv
Hn9tm/jDL/qpidtkgnk9M2hOduYoEl6itoHtv6Owcdwh2euTTJnV+woLvoNnMqxY2eC7P3I9UXsa
g248ETOigM5K4JoLCzJc6eU9SzBYpu0v07fb0YZrw/tj8myp+x5ULnUhrB8+5v7/QW1+ZxS9o1qO
V3wSaNeUR1k5K+cJPkXQIuspmpK6L3ifhX68aIqyOfT7sV4vnK4CijJxmdUHvZeWYx+yfLVCWu8Z
N22IeD86X+5OsY5rsXMWE5/7zRnpOWWBseGlWNIX3gdsIfUXM5pLGrqzQsf03YlaFyJEUtFWnrMx
DCDPfRJqYH1TJsyTMJRa0PSkr14PbelawGAcRAUz67Lnk7isVD30ZtIQW5+O/XlEQUclyxSYB39v
tZ4wvVFE8MpAWIHCWsv6F56MC7wIGSoGClo326F51cKvL2dkhN9QdjPz0R97NF5lAkpsMZz9scC8
Qh9CznGlstcvrVRiyLs0n+EFICwCJGbH2UuztCXYjomvi+HdwdjT261+5AJMVcagVQKZ1vLqYHh0
xcHvCA6Y2PiaKOKnhcMySmcQCH1VyVdUkJGL2MxemvWwSxYcFnc49Sps8zB0X8KbSHNuuANirgu5
fPf5LHTMJafZ4ly2l0oK1tyqPYhBSa4vEXNYurXm7EIjnuqVlT9HDpO9QUltvES/hZQxfTDH1qbg
GxAxeFTKMiqPhhE3XztyvzL7OraCaBaUci7HBLqMnhpUYafQuW61vN5KaaDg2EwzC+h0Aw0c4btU
ix+4cddZKNAHyT0o3hC5/7KjVAo7XkaOCZIOlnCSinXgON9FeLv95y7+BQY01yL5YkDH0nC/quFu
/+LHaq70jWSq162cii5NJWTmTTGnFqxj6FKwEnJcQiq3BK9LXsj1V7F0YarQfe9eSGhny6YzRRsD
UO7E3cKbXBpZdnXlneEFT2Ybc4DnA3P+JY+nFofvtxnxyRQi3mDDfQ1PAaJ7+u1ndG447MLTuTRM
XczWOgxopBc9eEGjIphbFnJb6AhNLcgtgZJNWWeOCngMRx8e7H1JvLJr15YM6G4tpNn0nbxEmAxM
Gdib/s0XcwcR6CmYwhkFRYAQqMT/YeWRDJwxETYwz5CMt98W1cm+/KXu2eqeG4B1Fn4SDqYBOdAq
kCDmZ0IMIxCZIBVVJ+6HyYi12NCI5NMtV2O6aPC0C37vS2xMH70h3W7a+AK6RtrxuboufQHCTgae
JkUJ1StfpOGHR4/1AaArcVoAreoWMuexDDEuYxvPXbtmlChXCQQBdINt9P+mDowYexr1Sn6BvRd7
nIJDiNOoDfoo5AFRJir1ixZXOm6vBuWFQrAA9kKxDjJYO3gQy7LXVPSzi7uIlpxCnmIuiZZbtIHP
eDLPRNOqmuvF1QtMcknPVWh/2bDbYLWBgnaBe7Jb4/GD1WFuhWJW/9QMq4Gnmi/1PPxqD3Iz4r9q
omA5XGN9AyOF04A86cdeRq5YG3+O3PgZ1LpLMZdtH6KDanontaRGdSwNOShRhF+ExCEmr72TjpdG
Kl/WMvR3bYQzRehsXdFXOqzZBb1oAKWTtxEH264oxCf8AIcV03UI9EwpxFMTPTCB64N0Ws/d2rDy
FgmpA0ZkK3Lufd31Mn7awd564+Tjif3iExc8Kv5xbMeTVm208EX3jAlm6UbJkqAanncWOEnN+yf2
YBFfvHEjokOVgUVtiu4dYIVx1RHXbeKyreIJc1v577EX+ho5RxTsir8nNKpSdjYRKf6cj/Xkjc/y
PlqIedieRDAQdvHzww5qip1eZb1Gb1fdSpG7Of2PTQFZgFBgK+5bwNh8mYC4Vpd+8A4AqwNtDl3F
c7lHr3OId9cU4Mx9P/1BGqd8/+P425zLxboucQ3t8He/YNd+LYtNy1nJ8E2Vkb03HRRTAtALb9Ko
S69j9L5WB2YTvAeEfi9OkRSVwQXfMuJ4HfCMB6CCjC21OxmF248h8fVRTZfkKtlmHtPTxuFkFSGd
5YB8y5rZKJYr6ritTev5R696cMfrRfbqepcRXW2jcoN9qFxWoobTZI22PbBELODgncl/mCQi20Ak
9kJyYjxVGpbZGilA/0YYdK+FRL1TzrfDf4wUD4izxxc7hE+qkNM+7FFu/6uzi6Q2Fq4/c75I9dnA
LTLqlntYbPVRcvSU17H6PCkZ//iqn0OzipoNTCTPRuDVPrHdloZeXZJDJP+kU2mFx0vNZgCQHiDx
JlB60UIX5qnM/h1czHrLbjO9y4VG91iVcA5jVFZmukJxnFnGHvOP6phip9B6k//Qv7h3uRxn+9PJ
pO5YEKA0fKJxeukLcoWc1twj7MLAl7Tsvz7ROvlvRBqHnNGSK3t+/nFfT2vtmpqhTXoskwb0jbg/
Vvxq2Tp1Bihe5PI2WLKvYs9CDdqmuisLkI1lTyMQJWjRWFynekqbW3u2/QFPKCY7qInWN2S6A8lK
8IqMvVEdcvoSM+cBJZRwZMbRZIVrXPTUko4QyOhmQHTXh+xbuIBRwEkuAGsOO85HUcZPP3s717qf
5SlhpSus831rBn1dm6+fT8HTLgDOkR0x5WQZsli/zO/PNn68CBzKCv+F0qaDlV4RRv3Shw28X6LN
UwvgSAlKe2/lXBB4h80qB/zz5kyyaDlu1AzAaQ6kAAhzdHY6GKoXefmF75FJLZTuad/M7KXYxZO/
n1QBChfp9TzZoLsoDt81GEaQOqlIGmAE9+JMdyNrbIYEICRqyxGzYF7cNRgbKoHuQcei+hFqH5X5
92k7QxkIY6yi1CkE5ItbsAPXT0F0rpz7Z6cSCiieGJYAK/YQgdqCWOhBqBO0kzaVY/Wa+NnWx2qf
IO1zt9Nba9SHq1iOLfo/SJb0M88t29cFq7XCCjNoqWOEr4zZFFxqKIByZUaZ9eUWQX8QJ79I4vnG
v2DMSBRBmp8qx27mg73wAQNHrEm2KaLPFUZtaH2nKjsXiej12QSD/RvwgW1IaeKV8/SUE0dVPGdy
R6fYRE6SGEPx93IxlsdnnNUq76vqf2KvaR3WD0dkhydSosjQWHMF2R09KrYwVSJyvLRbNXkedTPJ
o0ifQPACMo8un/cnyPz8NEVfhyyFYkWGB3LsQ3dD4T2G8Aln5+DI/z6zQOioHZAKRAzwbKC1z97t
yM9VJIfXuqxD4yen6j1RximJqe+jBhDWe73aoJp505fDBdxuD0yGCxslLbpWnYjGgWOgL8XYYb5x
oiA78EguGr6QG5i1pRJBeq8BeJiUddgkrfofKkB36NsQLdCCBlQbKNVSB9m5Qiw4aHSzH/CprK32
QxuJZ/o46AXK3fo2r77iDVjvobieCN1THOzKMymxeikH7gMr+PC2XNktGiLgqlE0wWfnfdt/d8aS
tNheZGTdYWSvlkl80gZKZM+gLYFtmi9d/BE5j75pZFj98EWHZo4YTytuUsvKgenrE/VFN07xk1OL
Krz9jCq+r3hI7NaSTLN/buU3hWMPHrlC1/k3x3ad7rivsl+EPTbYQN++3dtozJfGilHtbOSsP5mM
NveY6Gj1RWaYhGTBMOcsz/eCw3FFdAoKq1MvWsIzWlvxxVpWtXrzZa8F8zbLKfrivgzSre4TZ/VW
kG2IoDBOx1Noesjyd/FPn489GctrIna/wyhPRwwB0Ie2yQ50q/KnixdGOREIas4wwZ/Epe0VEOEl
0UMQo1NLxY4RCR61GDZJbOWCIarykg7wm/fwcFNO3/KRr424g7behnA2/N6/uWRVIovYGFJuap2P
SNBIqBirXX/0Z7paOuKOC6EopEBLHYVQQ/o1DbK//kl64u44F1nH4Ph+gUAjCG+SSkfllHQ4dK/3
IOCygf/L20Ij9jj5IUKBCEpzw2iF2WOC3Bjwb4e5eJ5beE8d+rxFpoVwSQziP+1JFXX68YvIcDRT
FyN2JepxXORAms2h1kxEM8aAdXotCVBiTS07T9a4KPcCqAyzJ7fw7oPCDE5n2ZuWsLgJnp/n2O1b
WnW0LNHSmvxYQvB5BWKeT/TJISn+C3lZEQA/FKbNFRN4BLpb0rRA7VCm4dy83EcL89s1VN3NTKPU
k5UZ7M1NSL3ZUUDNvF2CMm7Ul2Li55ra3FDlkIKUecKIbC9O/xIo+F0KTtA/YvJxfs4VJkkg6b0K
W9G4wNwSkubSrGlthIkiAEntEXjP2jJNIrfFVyFBr/kcGzth954mYU0sF7GNYMrVIgkundtxg4nL
RWAqYZXvlVUpUODwutubuUKllU1EitaefBjlYOaVGHadro9pXUsKXlZBJZZxtxkWFEJyEKPW8H/q
dHfnRBUZGPORCdP/nYweujFU1vGMLJsxMTM99vLtOu/ddGGkoyBpyqK1lrhrA2C3EoCCNZxv2iLg
g7p4Aiffvh8ldldp4F5oKKB81yL4SCRz5pgv5R5CvVnURM2jdVHDzkAKrImKaZ9UHMgoFii9eixk
6hrVmEQBuhm+oil1poZRflhDejF8ZFrs8iacCOQM2UftMS6PQ943HOdaQcShWluO4tGoxCS2Tc10
n1WXmypfac6oHtJkOr7QetzgtLpJ4jlxoLnti/mo+PDC9y9SwSBMtTf2M8ujJD+U+2+el2iF5aJ1
gv9Oy0ZYxumu1hE3tPMrvE9MpTyE5/HQ9HFNoAluuyPuW9QHUnKXh5qTHxqrEDtiCztcVn5PNpKd
LUzW2ZVHiniZbgwnWu3kPZ2ovUzLurXm7u0Gkoc3Gytq8NtzMabmpJ79RELR+Wni1yEp+mvdWZEV
2rEkn47TUZ/iJ4oeftLGdlfl3h/ifDTnafkGgRiGA8cIcyixUpqRgoos7rtBeOogPldanPcOQdBV
UcgiMt8rL6TKDvoMZhZ8Of37vqKgoA/oZRmxMEiop9JOXtPwmcsd1cqAabbGh7E4WC08hy0RJ7nf
LsGBObMarqE3tdkeWq6E8LipV79Rbzlz1IsWLXE+9pXdYj6Lsn04USXO8oPEPa/lG3/uMy/Txtgg
bZz9XLPXatIZX2k64j/j3nigwIvOHzPyJqOuzAbewPgJHFtW73bZocnhQlOTHROSl5huRCZlTQx8
pQta1Ea4m22ZYUNE9BhMwL5178IaTJc5HZe8gQY0X2E2/bJks7Ezuibg2fSrvXOTAq7Ruo1wag/a
9Y5zOk8i22yIf0/+H7ER/PpFj3Y2A414dNdALnx3GXlCD4e8p3C2EVBDwHqjCjaNapx2jqHtMjI1
CDRY04hioEEFQlOz1it1pZyPH/lYY3TkAulypj7FqOSOpn7xI4oCNagXlWVEi93NoTORBUtMZl7p
1kvLDKastlx9L8nj1STTB7FAgHBfzTkF2D+KAhX2DfmYcWSYbq+7nohP6VJ1m8Ha0nFKLm/rzslP
H8/qLyyxQaVrkG1+7njrjdWLpHDN77JmAt8s6YJi1WIL2oe8eY/jyh83BANrXvYcoUU1lZ4r5RPZ
KyAUjN6ssqQSneLmJjZEJ4wTHwan0YSYbDwOrO4tmaETPYh1Kt/j6etq2O0oI3OPugJBVesE72Wq
4thwMNUpmbT8QFSSWvfy7HCBv/0s227wQGAb+Cd6yep1Mwy9aTnNL152X33ugqaCGK2H14PN5K4U
S5Xg2x8MH3nd5moU3vkQMRIP11XCrDeFmwDQseBE9sp/5Cl+TqDkMlaWPGT+0DfoCHIAkouowgUm
yuEUM6hzFKN3tXcRtwA3EKaN2gLVb9KvtUoCOsiZNxrZs3+x0aydCf6LDSuRDL+63jsYR/Zuln9K
18zURoizAbXIPX33ClU6hFeA0N3l02pxGR/coNssmZ8kGHiuEG36YKOsxGQG+uAWVRvvSz6ztMq8
eNj1NFFerZ7hrXKAST+sW8MBw9TDglJ/XA9J8CiF9QyaAX9S5pSfY0msmJklLEemGPj1yBDljIUT
oRU2INndBy9TsDLWcez4PPJLkykdI5eXyY90XE9QqUaPviYtx6JmsnSRMbLZOAgklcnG8KyFZ7Nv
Md8wgh5EY0Jj1yOS5Fdov2t3gg/moaK/IC2rlJUBG39yipbedTZAxsj3qL0R+jBxjCQkeUWiIok3
FVs3UstetEfsHRJ2jDmNaadIWOdEYOk4FxKN5LNHFdAVXAQjhjZ9VbtIGOnqCvXcirTZ24kPq2EF
ZXa0K7ttgdyYuF0laPMXrWBTBcS9awsfNpHHF0EL3WxkK6XjfjnCTwFPrnc1LBru3Ejp0PJNAhfY
NlUltT19FF8HExKb7lqH4BU7B2Q/kTp1g00/05g0IwTzsR3jdASb3jwZFZjaJOqsFxGz4u7MBYLJ
d/SSmxuKXRqHYnaVFyY+bpTc/byUGRj4JSFWXloNsfwTiMhew7WQqhah80xbV1BZErJIBuKfSr1w
BFic2wre/KqAQi0BnIWak+a9uWW7lPD/cgqoAL8C6ypznzKWBq5+uGIJ+p0SujXQeRH8M2FYdnrX
6xFJExgOK1pHvIUBBK/p1OtU7CXV4vjaA2XYGr1YBjmXV563AlBFcADfVSJfBjdB9RqwOoC591Ht
9J2Ov74Q43jVgPE+4GjXZ7OERJpFdYNmZ6MvSzmW0focwvAl65umxrypIfwsd02qy2yHOiB1VzC5
J13JPI3+YY0C605lM3rS4nZeiEMZEffBsj3MsuBfdf9f4xZOmkW9LgpYXDjWU8ZrMkRAbU7vRtfu
Y/XUkZiGBFN8jnOMzL90nObwtq5o173Cq259NqnHaaNByVRA1R+EGwl3ZI+rzW4gXiAQbfUPuN8d
f4srlEt65c03nluNYBWXX+3UtE8iyJItPlwTmlI3epNSTJ0tDoguhzZvWfQDJPF9rE5RoYq8xoux
yj9rDJThFfIR3HnXqB4NeMe+EsMq7mHOy2GbagGc0M81e1e+dpt3WAhF4+oAlKJuoVcuJzne1zCC
m6JTlBEyCD//8FARS34QeCxexNkUiPAttQXpKizH7jYxqx4I0fpDko/AOGfFbBgKK6UieREFND4Q
CZuU1k7X9VH203FMchkjj16c0whgJi1G0T5eRa9EKBtWFeUkh5FrOcQK8M5yQEKobBFmkBXmIYY2
zIoAR0SXxEvNtGNdLDKoc55cUlxxfzyDa6yifZSteP5SU7I0ih9OFrXnbHxTepUeA6xE3TQXOS5c
3pgXWPQnA+wxMva4jr9qVogEcYRXON8BRXAJjJMYA3jTyDqPQIsRS5amuczwYlh479qS1B28wnDO
lrQPBON6CgYcdWbFv39fTLiB/ssUE+X45O0cpSnGLgrIjt0l6G0ceZfECg6X0Z6/RTn6h8xvRUWh
pBOJ6pQ+zfUdIqSVl9CjlvObgjutE+IS5xihm9AtAoIn+FiUWzTLvPTtqnKE7vuBZR2KQjKKIv7l
AI1AvvXXEYA7M4BSmh+A2DRoRIeH4QCcjDHvsBCnL/ouDgw0Is2aTV3lJXvImSFj06IwGvVLhw2Z
rJwLkX15qPzxfsdAxIbPcg+ljCq0+1q6hVIg4j5rknfMEckZnejIlhCVwm8H9u06AH4/QQ+y8uxV
2k+hNsV2ZiGYIGcxnW6qrAPW4hIECIUvQocwRrWm0V9zoYpQOEStYokhD9i9ms5dW1mL3ZNPMcYr
UkvCoRR7ca7+sqilP/SEisYfDly6W4gRDFzS8GVEOAB2eUuNyU+PH2C/EujUJVFtTn8GUThMk0v/
DUffytVMUl6rB6lzvvRO2Q/xOokG7Ki7DD6e/EuFE7/R03Q0n4bmudGUEzNahagNyc9RE3ipJMrU
JhO18bqpVLCbL6jUNILWTvLq0zxUyvYfk6mzVz1tAt6kZzNiy7LIzRqjhEUnRq8exJp754hquh3Z
xPwv/w/JhIPmevTPvp9tU73lwZnz/9hxfXFpqQm4J1S1tNYsittnvQaSShD0vWW63k9dP/GJOk6t
FKL5uEm8S9RweQ0aJlNhGqLAr6uDGILiG18AiFNg6kHU3Ns2dmI005P8QVAYnSUmQ0U+5sz5tjUM
O9vwVKnkXg3Xy996C8e40sAyXUfx1RFzcnIEpruYglwyINcmRTcxt8RkgrfQmSYzyPew6Zhfb0Yd
gZboDNO5dATmfS1MCNiDLEfWxRRVi9GhQe6AZQm1pisqWm1ab+h2JBWJ8oKYZ2FV0IwYOlRGaR3f
ynt4e8vEI9Re84M9BtOru6d7PgJwQJwoqjOLBv8Dg3lqLAPzYXF6hf2wz4kCEqyVyecMiz9wwM18
jPxQ0i6PQ7ygHIEHblrnjahAGEed35Xats0k5+N7cBgAIIZ3/Y+cvI85Z5oTso7TETBAZTNoALEZ
3q5GUFvzh90s3PDXUnq76MWs+LxRRwp9UO1TdjB8SKm/OVkIggsY0Oy0A3De1+nppzOYk7L0il6C
sRl5QMQOKHjmqb14n9Dca9mRaf/QHJRHCTztuQ66/DSgM10gGf6GsDhUNaSL+NzqVWoKQkwTJsvZ
nNUlE1GKYrcbt/sEIFpOh3QjF399qak5NcXM/Qmwq6SWm99BoNL5b/ZxtESJM/FFdFwvYlBPA9lG
Z5J+fz6tOOB45xSy/LJrOLiqTUPw/tr/3KIKV5ndW3rECQbNWPilTJfjJpKdEKCyemcMLisCNskW
EWW/WhA7t7e2rAmlbCEk0iOtS0twN3nQGkzB4mVlt3/Q9oVf0MIyUyvqGLqp2TdH588hq+wZU6zL
RzZJ3mOWppGOQGz0324UgBPFBf3OP6vEb4U69wh8j7veWY3YrW31JN9V44MrU/csMkfs4X4hd5uQ
Q0v/SYahFqG46dHK0jo4mvXZdMI0kG0v5QweQW76ZzXx/d5tmEyBpnyxXNQgjANKexMGh/90RebG
tYjRzUy721b+I5wmngQwckXkU2vAJte3ILIpprVjcLi/kqAXiifQcSX4aAs5Z9b6tfkUFZk9pMqS
p7Ii9U9RfjiHUyB+XXnV6DFsm9FNb5Ih8alnOnvNXB6diBYK3T8J/loyJA7BNky+QrvHyrJnkm5j
QQlAJ6ijwyRJCb/vdOKhTeagU8Uzws5UdRAdl8vB1RySwCghAg5Mk/2IC/QEkRuW06isyojc7HBj
ud1bccKjZgGJmNZ41JiI/nt/sLbJLZ1fc6ilqjwXNeoiqTYw17ET75Vv0IAV1AcL6PPHl/T+IWE9
+MPBKJa/E9RHMZZbQI6WEN+zemc4oCefJpvDYr1+heZrNpYACDGtdyeQGi474H/T0wBd48LVTVQx
y0fJuKX/97mDsFrYo7b0+2jdjXPIkmwfO7bb3vHpdekoyyJk2rlcDgXxIg6xuL6o7QoKsix2USin
oK40u5/eoYGY2htv7n6octK3DQjKMAxilQShuQmSQ2tgtPurJM3fr9EBEx/flMDMOCNA0NS/YorG
wpmLfVKYEWfkQnNJ/acBJ0z7Dl/G+4ekR7T+4+b18kBclJY6KcyNB6tabedOxHnZQIP5lMRjhE/K
KJCb5kFC+N0xHyBbiYk/Y3AICdnE4fclq2ajEnEyJ6b4RdwfRtiu26ZN2c3rqMamOOdqNNdXxgrE
F9oQ2G9ApSHPK6OarU+/OYTQqRbVX8T6DjjitHlrKS0U35J9E8IL3JjwcbsLfXKgKLwjWVJQLQJq
GnyAnBcFtesK+m8WxNvtsJXYJeU66KZW8oCXFOqxos7rMwxbIOTvcugSunY2eA58QFA3jRGviAy/
MKLqOgo0iJG3sHBuPvSDCs9hIaqlK9Uiu6EteDgp8SVf+8Kz7Uq8FcGkzzLLjTFO6yBczsrdAqGy
vdR80Bhm8ZZ921PFt9ed6hIW4a+v/DCEgz27GJjhNh57vBZmwZO9GkbQV0Zs/iZ4HoF5UsHcphGE
D1VUUUHgC/ytf37uKrng78fYK/5HS5XNjgnBday+9bQVQ7euYq/o2eD1+onC6s34r8a8nguO/f9J
Gbr8PpD5aqwEcWb4eEQs77Nyylnsde9SXZJAqNPH891CJCZeGtf/n3XTTBULm5RCtFw4ybYfLDsl
6PmNJ1eMaFGn9a0Bm4iDkUtwVcZEKFfOdpKbY227VYyMCwcQOS7ZyGsQvQb3UM7Azx2KYrWOsIgo
p6Za2i9gCOZ8fpHbAl/vP529LWSfh9BqvNFY4dQ2G+amNhZm/PsWKYGezKp/lBsAwqD14fTC6vd2
1WoNliYy0hOF0Sp7JUfUeBWi6kW/srI9qk5OE1LA/G1nDgNpnks7pIoQXPv9Tanifz+gcJayIgat
MyQ8eorsUoIcba3YvI0LPXSzUtd5z2KeXTDcpu+Ie6hG8eAF0tOYESUqOETRXv0JsPvrqVnmUKYI
kuAYQs5PXDoqCYkxQ3hw66/GWNRS70pXDwa0wbnuW4/H7jNTG0kQergAfhfmQ0+VNH0X3INdjvta
5YfxObvl09utkv0RczlWOIkHXx7AIO4ujo1KpL6zEwswJBl/XVDSwTe81qphKcX0KWBJZmz1geUg
O8SJloIbrCg3CFvNMnZDW74c9O9bA96rDEE3Os5G4zGBN8yrwkexdsPSxv6YdQpCj+BLdiFeNUB3
lF7nJQ/blC2TI3KvrbEB6nEQ9X2t2arTlcTfVh9V+SQm+nNP4b4jbroHYpPokt7Yz8+F1gvwuSwJ
VkgfSGJ2zU3lfFpR7XuUiIov06dRUHw0QHpwRWrO7NJGbmAKKxvAkfy87tMd6T1CNH5IZURmuY29
TZDLrUDD+7paYrc/2IvDI994f09hX5xfTUeyjPmyjcfhKT7WUPQkoM1XHOZMO2w/mlGoFSlcVwyf
AU477Ayh9vC4nyrEePMrgeZNXwygzMxbOoZo/LtorTq+q5CnoiDMlKXhsQz7rAUEooG6JD9/Xo8J
yGEhd8A4DrW/uE1a3gzRI9GOj8spRPU+wCPpGn03nBfgd4NFy7g+9qbuDBnpQdkfcTM8DQaQB+OX
QuF5htyiHAeFYM1Smde6jguV3RIrC/jzLRbonjLmq1XzY3pFLrpOpo3EhI4zYaV9XE+hIa1VItu+
zRVRBHez72M0NsHbzdqelUMMwj9g60uft6h8aaMZd1vhheGxFzMVteLnPWG/YdAOULdSxAYl/E8X
bNeEfzhhqY4csQCj7/PHhO0LlA2/n0s3syCpK03LOzkQ6Bxf2dq9ux2PatBcjDSxNQh+Yaer9LgL
iipb/3ym3baFr+RTEFUE6R12viPzQh6NmuIlPL3p/+iyJ+fMKiIznWZFpWu2ksTzw19cI5QrLugv
5dIsDZrbTzWcOPsPNPMw4AP7h1s1FSuBKRpWs4To7BRMr5lcexA6pbD5w5GnDm67hKLkkIjHkBf8
wwzJCcjzQTxIv77LRBleY0lJwPJMAEKDbSiVM1qKKbHUkC8j/5jHBqZ8u0bOoCmAS14VFHMquW1w
vgvmkhiHHHB3E48WVBHaUxeekFNh7krulBFS4+YtJgnr5bxJI/5gRO1M8TlQdcnV6STPWzsLvOwA
2GoKzPPkRxqhauIZ9mYjOlx2FgSqM3G5ht0idFQJazqY/+fWxgZWK6blgs1cB4Zd/bnfPq0XT7wK
CfqBXeF0rR8KjNOSEZi6nxNgWpzB5xxgncSgHGdD8HvH5gJtPKGdx5jqQzxJPPTxO78npLQVilxK
lCm5ra9gbGS9pyetb6wOeOHkyOhGlvgyDac4htzFJeD61WU5O0G76YInCytqHtq+6oJWEHFPippF
zi9kAkv0o4c2ixp24X8qjOboTUFyZfNV7X65mGnMSGIeqdjNu4PtzsCTin5kaxrYcJNk5aTCqEFA
H4BZxga7+8oWpNBvVRA2LZJlIHdRGbQPxWg6jqIqLMlqMHW4h5mmIJxkaqQd7Av9Lv54TvSh3W8n
8cgElmvC+d34kiCd2ULBrnnnlN+/9uIPye4k5DYP2jSMDFjk0PMFdbFV69zJFdFMx0wt0Z9S+mto
MnVntQ2H6z+/flKlmkVb8cVA1fwK79VwnyaFzh1dJlQj9uOKe4C0ld/CPpRDDWebM2dqmYEbV1Vb
OCxt5+gHoJAdm8nFecKFSRymaLJ52SMMolmz3Cjh0kV8Pei5G04jPRBJlrXAYDOhjUffh0uqwE2g
NyE6c0mFnq3E+sP/vUfa7/4uj1jk9JW6kZ59G/qISdG2XR6n4nwvBu9HWLcBYc2IWAyixzWAPghN
NpEQPUv3JQogc0ZUb2lea0TD4JsN3KqZKF1il7kU9nO8rlOjWS+buaFcEzSANba1qDX00ya9YjoT
3iUfLJRZrCIq4BQpwewTArhbBuzm/nOiDbt0fN28tYzMWJNIgCEBNS7D6hMCOIzb1BmUuU2dcC6R
FtnuFI7lOQXuk6iQScYnUmAyNNXUrhCufYTVly0+zA1Od7zg5gm9DDUbJYTmY6oSDIOWD5Lz38se
3V/krwMl0DHR9IgScQ5S9zgAqzET0SxLW8CuVNRA58w8hmJKXqlXCThyRe+1v+zXQXre97CkoKVS
JmMGndqeIJx3ucEBlrlwnFjOyEo/INa594TJeiuYf48h6ggtGgp3FF9BnPs4fhddr6bPdLqILe/L
eaq5zVG2cRK0D25lPm23SaLfEkbbwCThZvPyHXaLVkLAUt+0vWke5WftotnqyK9s+c2D209Mm9J1
oGC4CnWQIxGUs17CNBxxXYX8A+KoBDXmwdPAKsRUYolAHmQwiR3Rg2ozMdzOU2nmqLdD3nzcfC5N
voHrgI22JqhGo3gwsRlfA8WFDEl7ntKCBdlQX0ZyxtEmRMjorenD9JQ0KUB9OXf5X78OWOMvfslS
YUs+pf+mMqefrCraVG1COKBbjjSH7Ez+9+FatjDQVNKiMCcjlBvDgH2t+Ho2ZAk9YZ8cZ27ubzEB
uHaGsPgWFu5P9PkhwoRj/CB0O0UPdhnHGpSbTMLUB2MdOWaj4BPnlaLC76R2eAcIiqgDDxm2oCXK
l3MfCMSEd/6gior03elqB8bdvX7VNbOZiM0uXKSalR1EPeMpVI2mBgKbTG8/KzfR5cO/YabjFvz2
sONSemwRqB7+BPQL89HGcFJnqDOJXcL15ervEe6+Cc1AxV18nnYsz7gX5TrCnzJPJJ3VT59r041R
pGiLESMlV3nk6KO2LhdG+zkDCZ2n3dr71nIw6r6mM9Seoe10i1VHcEChbAihPC/bJYRtuGfXfVAb
QCeE0CMkLeEirFeIvCjYdG1qpoI+kef6ipTwFUm8GobvuNkBsKgMkYrRmCQoVdzLu7BP+LCsBiPh
SeYWCc6mqGJaaKVG0cmLW/M2B5Att9D6wyOZCAkSVflENCWlgxnBVCiCZ1NSTNM5REDRSM4koBLQ
auFB14F8296O7UV8MN6Gzmdr45zDWeov5Jx/ZFQKuvy4JG8wj0p2lHLmp0E5xhB47lEGxUTuIXAO
SHK79Z2sC+wULKtrgvyO1J21D64jcwzATml0qsSbCbvlIg++s0cibRhESNuPOLM0NBkWHwwE3GoU
mc4UIZmId1mfg9fDglIV3g4xWN9AujgdMyB9KjH7T8JqlMLrvttNBhBwULzCjtAppNl1avQgo/FG
yE4ubGgi0XNUppZmEUTsV3cQoEt8xRieB4PGwpUdl/xGHO5SXTLG6Bkt3YVctKuwv567SOOsbPYQ
pXCTDIgzFAlCqjLy/ULgFe4blx7Ks2Q5KBUu+dLdZDTyHBNz1Pvgy7Mnb9NSJt2RODylcQXXm3mc
Fszi90QS6oAVoTwDc5AUXrffLecTadzH3r2Aa1J7S/mU650NmZY5Cg0r4AE/OxiDFvps4nhOwUDv
F3Hch7pc2s/Aymd0eudwYG9vLjQv3xLlMdwHzWlSMAxPQX7IKrXh5Zx0Q3auk/7X8/M1JVc0S9Xa
D/54OHS3y+eguqB7H4V1MUV8c1bI2RFs3tfvtoKhrcpHJK+R1W5mrwEOtIdp6Jd/EIqSAbaNb55t
NdqX7soTlu/suqflHUfD6cResQ2atHX4fNQZv8B8jTrxyIBLAAgr8HiCVIpxHDMFvl+8/ouyN+Vc
+oPEvNH5vuur0VysF8PgvWbAzNTcMx7UoB31mUkhjCy722o5X+rHJwi4b7GMzpdBZIewEyvlKHFJ
djMt8Cub7Q8FWHoinRqEG8boi8/+L/3la2mWk7BGBidhYZAdebEkmbvmLdQU29JzBtcsLGI4Er4z
+iuupev+hkNvbMXkSFvAQiZQWVLq/8zlepK75A2DWN5diu9YXrIB+li8mPJ8zvzTu72CamNNNP6d
mzJ79C6ADJjJIVenwZb5bQKs11Dkia9pMPieklfv+Z/QVP9DgkCkBV04I2Qcm/yrJIio6SME1eWz
NQNljwS0C8q5m3ygzX3kvZwFwlHT7vXWI93mqiSxKnxli6/GH5BV2n92I8vQkWy5WeMTr/iJE0qC
q0+ZITWccgFnutcbm77cWItmMm4lus73d/kh836g+xkUfgevo/ooZ2oCZz+TH7KFPL2dFWLt5ILQ
i4sFA/sXagBsLEZjOERZ0JNMDD1BrqwcRcxZvIv61z7u2CyhEWvQPQHQ5fTDrtqFY/qkBqZeTEnr
/8W1NPU8zqv6yBPe+DiVCnvfGAdGm9S6lGKJX9OuoBd/E8CIP5ZCUOxxQhnKvVLxL06yaksIko2W
e/b8V0VRwIlepeiSnGJurMTNp+22cTcfMXJljbXP1YUhP+FjBXAKRntYMctSCQ7zNdXCYpQ9GeGq
gJlP3jKZvI9+lexGtmbZNwOJF6CbEmP/Uy0ppIDUHfnJ/6X4U5+E1vmVAJLZRzeg8Ekw8XAVmTn+
+s6MlPfJ3KIiQAELp0mOvDCx3v+2Hkj6XF5CRBkziOF2hv2ArcNflyTPoykpbf12rnBiisJJSwIu
YtowMI9EyrTRrVYrJM3h1gyiLVcizHh82pH9o/tN/T6o1VvuoetyEb4E7HiN8ME+GKNv/BfMVyW2
F4kqKu4ln/NWNyCcbHaq8SJvfnPKfml3gKb/TqSCmEJCMv32/ZzTziXSghzRExM2+sDgukdtVAss
+u00cadM1qYdIHzeTJPzo/Acfs9hrr3dn1SEq7S85MYtaoB6k+UfGS79BoJOf+7NuX1+rfYBH8Oh
lE6iZDIfEgnwpaa0Z5Nn++NqYnmoRyMgTm1hzyRCaMSbu5ilaj+mxh9Tgo4CcJ7LiH2zM2khIvWK
C1mjL781e92fBUzpcmC6sHTrvFYjpVqnUyUwIBqhRXjpjsjTS08ZoBBkOUkODikAHNf54ln+9HHD
Ta0hWyfKH3ReztRBuca/J3hFQM+TbPYKfUGKaT1Ix/0jdD3E4rOVPegcYmZkM8yZSfcA8PWW+b7R
RdoTgMNu+fz18egWuUCfoOMRk0IefOcDejq47hKRGSTLU5Ty3aVtUOnUI/ZHAT6iYBCj7w1WUfOO
ydg8/Na/GeAIWm0WpoGA39G2T/X835vh1R614co8HEqNg4y5McaJ9OGZ7JUP1mtByHJ0hgsydzT1
5Zzk4T6cP7Jveq4I2TPHzpBxJPi1MkPcfSoUWqtqw/cdJzAekpjgz8B1HtyaLyWuOtIXOUVM1JbP
zgzxDArcCloirsUvktfMJ4GOMyb5ypyOenB9yX4GP3lQwyGS5TZZAjDT9FFvnDJIqWQZzp6safVD
NpeoSSv01xZwYhwadTFFm6+NhhVwK5OJSvAxP0sTFn9k/FSdN6u+mm0pFXWQnElvR+RN56nc1kH+
VwD3QLLGA8n7BSBBCLcUYxrKf0Oav7D43lMtRCm/g4JfTCaKoewoOG+EdFZ4pZ51tzZSdoPtMgRL
aAJ1k1dXxOYy5AzQGPRwN6BkOClYtK/Os5NfQshHzUyDfhBaePgLQvyO6QzErP6Y7G7moHBNnNlD
b/1k/LFCUDVBfl121nb7cDIC25t0ZfEF3VWvcbV3ni5AbiU4uHCoAXHio19kwNKWNAu/lTECYO8+
ph0KObko1xiIRN4ujFhOrzy1vWNKwLlxbAv8ZuTfdwDV1uVTi+YB0u9poYcgrsUzGHVCIjFt0S+L
bY/rBKUNQmQ/sEa7LdNcdEYVeLwqFxSY3ckSHSg9Y9EHcluchB26JloK+Cv4v5mtBNLv3GtL80yW
ANQciHWHSoUTzQC7c6RdSTU1Nqrbt7e6koruesHFbxDzzThQqtWsxpAiY/Ld2bB/RswKlTGvnN3j
hGw8DqXCDYrPkYNSTt8xv1iqPxxB6unuu1W36gqcx12/fR0vYxD+aut8ARPx68rgnr+2bWS/4TeB
ZMqO1hyu51fcO7ZTBBLwvBD9GMWdTRvRXEOV5HYTXfitLE9VF7WnbPMCcfYURk6eF3oqBk1SWSv3
khNRJMeap+5jKgh7a0Ol7kqNBueebLpN4kHQO6bq90va38HMAuE+sRVpabYiTawdZzX7QiP0pugY
WG1T6niT05zfyJAO8zf3F0ybODijLq52p8a79Dj7/Kp/nUFS/JoL8iBnN2jeggebNYAur3BozRBX
REHWZuGgXN0seoTfOrwwwDPwItEfns2TOeDe3+fTVAunWnmIlln9waSQft2P6lZ+9EiMDDGLnm5D
YUUvpU57zDd+GXKHeCAP6hmMQEBRDAFxa0zwcgyRMFGwHEy7O7J7bbr/r0+yDlNR1/Qa1AavinH9
PqIx/gNtXNhwwKghD405/qrTB8jhlrTwMJ9hXCYZYGIXsnFxZa/DvcLzrTWj8geYGUUaaL5lLW3b
MWzjLfI7pGKmy2MFeFtgOXq43C9g3HIoxZ0NHwg0QSjKoO4xDL6Kewzgb7tsglGaGgS5lu1f8un6
nYzEtSbI28/5lP3FZBojT2u4i3J7NOj2pfGnpFBPV++Yww6nhIOGLVr0mKx2ngYJH64HHcEqIbNb
zTCEDV0fvkS+MfKg/oF3vCe17KGVFW2nTabreRfwPY6djYtNNTdzlAJgGur72lJ4Pnsesy/zCfkx
bAJqzZuEp8qWBVBDCqoMhkJY9E2Kda2YfPTv0RIbMzhOQblrUKsPbwpTBkosgUq3L82z1yar0iLx
Gbh9mAnszaAPPgoiFp+RvEgOxEwIx4hydO/AkXSA8V1il3uiOceYYd8IdX/BoDL9G5a2B28APcoT
+7NoZteJCr1DXDRxBrjA0AWj7pnMDAGI9LQVgJCmAy6PIPBfmSFUyykPy93hZS0wZZ8KIB44TXLR
UCZZzJ64gCHMJ5LCItUfkpkC6Opp1OSHLSVYQh2rh8xJWitam4cEJi4WBbfySHJ1Fm3QV1+i9AVd
CbtMO9V1iWpLS2qRya138p63IAsmMUSwuFAMrrfKXVFVsDDn2NflmyypmGCX+cOGLC3ABwrRDaPm
58fTrcI3ysFGopWQsDmy1Z617ey1FIbNe5pMziJjQl0p9NcSi5XGky6i9pevSSIf3buiNYSr1p8P
JnEWDEgrKBaiO9HDC4L2lCfV8yT4Q/hpvVudMjfpwomAlocUDg9cJ8MQkTAN/nlwUnqu2cx5dwj1
0zEUXKXVO44mETmeibwuKAN9pzVM4SrulK6LAupRNjMnxjUU+4tcEAMsY54iOaE32lt9vJj/UAww
miVHfRnKwhxFPHCh+qJjkznnxkjEkUdIE6Dejf13QMqePVq5UaSOwapDO6syGxOgP/c0b9DDJtcd
XeXCzcIx8bCkPrqFHuRtxHHuCoSLhO5Z+NkpWi5bI3YjNvCu7ffI4gDnxAenBYWDoUAISf2yZbOg
GlqhjfjcfoVc2QoLCiqJF/sfW4M8x3InTrVHc8tbCnaMGQ7NV0Numn4e1xZVn/+0k11ZvEy8xQ7f
bnTVxplV9FSwUo2xQiHdENJYDujJYnDyMS5ETvb+oz4fgXpzFi/aBGpZ2R0w5P37LdEI7AQFwOdh
wagopnUaBNc+SZE2dKS6I6x0Cgeu6A36rn7bGFkNXi8mifVTAr3VjXkTujqq82ExCd7mXUjEy9pT
3P+lTQdBYqMD3ie94DMzlhYf2GvdoDz4ENfzscFOBIH5h8eSftCbYcTDYlgO9u2dLlGmuOdkkrWz
MuVcFg1bgkl92phyxYvBaiFT7GXLyXRAISY485C+RjiUuRcXBTE1TeReEkb3Vj/2BDmou0VbyJxb
7Pt4WBLzBs8kDJKluLC/i7NLkBdeCcoauUr/73rubuAKrYt1AdtK2QDDIJCR4IhD/7suYTUG2N/V
A0NuQBsEzP/vzCxHxki6MFkHw2IS+SUGSOy+cy7m8nEJSE6hebnjqYXm1HS7kgeuB9X3xKB2oizV
Pj7r8hT2lw/CETK6OwzsscrqWRRAwtx0GHpiMFb6/FMw3ikKTo5x9eLfRzsQZig0TmHR8v5lCVRH
Ja9nWmNsnr4z6sgxD+waVXpq7xLhk552tSYf46wbRYMcttcIy996xWlVmhGcfWRf9jM7bnVSnpCV
BGAJhldfwZjvW6gkhoiyhAAfMrTTjfoc00oD6Hl4bkMxmhi44wyTvLSHHPKsNL/FaTAMB0zGpMk8
HqkTwL6UdRKsoIrNYaUpIZ7nIEDoyyOIywu+dTR896mSGRm5pzoylSM+IeaJrE6jkdQ9vFv15pmk
51U1wzjt4wz0+KYhj/RjOG4U0fwQnyADBVKMab/HsO4FVE7bLhdGuj37lCiA8Bi/xvXl4Aq6GEdL
2ks7fRxkzmnZ88rSrshcpRoZlaUk0ZqjEFLckeDOnnKupSUZy2NPUNEZkaYD3Yf6/cg8/UMZwZBf
Y+qpHopmN+IjMpKzNObA3Fz1XDzUPCZxHq5xnXE7BD/NdqVj9B2TaRHJu9stJaDZcZRLYq9yCsCm
MKqQcBgn5iUfRfjdZ8ulqyHpyEv7p6KBr8kvagYP5ucDTsU2aK+NWhPwfMH07OnzUNS7bcjcQyXC
rf3rGv1/ksJGZvYA1iOFSfK36HZsIDyEHtY7aGex/9tZz2UiSiuAtCyGb83Z1gjw9WK9s9DaqG9i
tDvnBWGLNHeEwVhKhebXGlwdKZjcaNMz9PlvoBzzkSFtZArqTzbbvtLHeTiOy1d45vwbLv7lD665
MIRD/F/TK4Wzcy39pumJ6+alq0qz84UnxL5C+6j+EN2vpXkqk/s2Obelj+TtDgLi41SZabzOH0l5
unLqCu2bsphIT51HbRTVmu9SEPDZAG9u6kANOKAZOq6g1bSinlTgjSeW20z68JmKtC0s4Y0jv6VY
/QQ1B3XamE7iF/dE5c6VFqBxktrYksYXf/Zi/IlSQL+0BMPwxRJ/6aIor9gJwKcBQo1hY2+y88Ff
oUpnYXeBP+U58CcfNSOO2yCbp4V1ar5lWyX1oeC84rmAYkkUKcyGvxdTE+fuf+BiYN/i9SL2psfV
/p9FSFBpa/pbgz3M/O7DIO9+MGxwZIXcVabtdompiq982vAp+AvN5ppAT+jeqoMeSyC7pRzcDGoN
dNH7O6bi/Nf7wVhLCqnhKPG0yIKsVWtO9h9+C14W+ZE7bvBePF+60STefBnwlD6P6GEG2d6GSMpm
RSSZnxvO8dbmiu6aj9YHMi0jIwrn9ccxkQTlI3niwlt2YSoh5jMPMEZpW83cVAx+5qim21WsNW+0
+NjzleY7CowEyAqx/nWLrWfQrGgBMPkVjv3T6SeEysonaoySwB4xBny9Wpx/agkejCV8dV+q9Xod
2n+/xsx1OKUSHDqEz19w5mbaw+7QGHGamICb+4Aa6oTSmnNW73FNy/zXAFkGe7C5I5D33bQ76gfJ
L07qi8Ncn4Wfw5qKEx4cExEsn9D6xSnSncMnls/i+cYibi4tRi3ocd5zBFCMbKq+qbP/yEn+uI8b
T/nf/KUBom2SYQJPuKP/HZMqGnssPs1VuMrAOoEX6FS4gzOOEZ/eCNHeG1qpFrlwLXXzuTpkzRt/
BnqDegBtFav02J93IkxKeJd/UiJ4MtIhxaX27CbyXO6516eg30kZQayvEWLRbrherhYiZ/d8Xg4p
rgtaEUGLyKtRiUjD4SJxYddO1RgcoD+FAWcm27og5mKM7+kftidIzFhWvB09dPtFJNapYC+amqeT
euv7RzURNztPxGaEd5V9uHSnChGs08Yh+xglQB8MHPjCrSbtryfOUuMFT3qTpJ+2vZJP/ZSNrmYV
aHMVcevyxfOp2vhoKt5n9VGqrQxzwS/nPbcz2XMFd08YIb0vz9pyKCnAwl6wnjkcrxRyMYs0zWUY
Ne9pxltEX8HRvG6QW7fGxUoKnroXGps7eicLJGWLM9ZFsRXERj+GMdYDhxro+4hX+ougq4mpj7Cz
iIkaYnmAMgHeNYSSmRt4m8dJSoVymVjaOVGKtiZ736ZXgEXXnh2Omcqv2aqWLjvIVar7kx/21Nz9
3xMtCdaP/+Au1dLfX1vRy+pJcGgvhoUS/9sGrCW1I4qFySN/atqqvNKQpOwCHtP3zeToE/RJnvLq
vYYJ5ggD/C78jJWEvLAwWQpNLFmVkBDIRwhlgr+Q0EY7e+dhA6H8jE2O/muIZqr8Qo2fYpekw3Xd
dLh7YDn8AOR1VLaaT8iqcCtjVIgit0yxiD9IgR8T+j2ss+9e4l9RSu4Enw8OOEcAK/3JtM6vhUPB
thaHX1bbdTKGs8sQlg+zKPhivjCD+nv6HFIxe+Q8MpTT+0a+OK+b0U14qdacvBlrKOCGU64fS2AI
RbscwLT6p3Az58e9pNfkhf4pBCMjTzh8nf1/FITiRh9udndCI0shabr4jkCqtV9VgusX4MzfXMZ/
JtWqb+hoioirZeNN99xZHy2htNrNIeMPTHPVkuEhS7NcyfsI2TGpKwkvKcS60lpQfQcVUNqyXUTs
v+hHaLONNqRmCXXBTmfIKMKBdvjN+7e/YECL4mgxG9ONIbVyFgk5BENo26gr6YaaHiE18pRwYqtP
9kFBWCANyek741QLT7XGhFX5lH/TXq06XsrrCzi9xjL4mPhMh82X43OjcVwxHt9iHilfAV3Ye3ou
QewARDZtltpMJAV99pxhRf1V7luhXC4wxXXjxioeA3MFu+hGDEvaf67bwxkYHxhWwDRZSZ31xwsc
fJfBeRsmVVl0qspvsZiK+IRRBWObplZbO6gH/kml37E2cYFaCr8CDDo7wDGgLOVDjpf5le/t+KJr
h0N+DuDo10d16uBvqdLrM3BYXJPbjyod8z6vdT8oqjrrNvTk2wTMvb5kXWc3MNXjMscx2qfgU2NY
8bmmgPmrJ80pT634EkDkDMpVk+F3Tl+8+uV5PbUTVk6BfEY/bo1ofLBIssODe+IWEsG4YaPdByOM
1+iEHNHcbRh5ecUaO2bNYr0PikGEKgcSuAVM3hs0y3G5OcaEnsWtYwtwYTxMfw4CjYU9kBV5KNaL
tQjUy3N8+xoGA3qB+N0NYH4ORYS2RB5HdGZDHp/8uRPEGzkP8wesTdn6IqM7O/3x+WMapRhSL/eo
c26CRvTQIHsn07/q5RNehPEfqy6ViGKxqM1JOOYwcKr82Y6B1Y9xrWC7uIBeFNFvm4+If3cc4gj0
UN2LcIzspBMii5fCyVFlOlAv5Y48lCNvlICt3bIpXwY77HdWJUpKLNUNAPkimZDVgDWxpieN+Izv
/ftho2Wx+jo6NTJRlGEsfXMIWGJpNYa+L5ny+Eu1GZacyNjMOO8iU8nP1GEM29VMqyLv+fbzU2dS
LWRNBqELy4QtJOh4ijL2M0Y1LpFMFIWSaBo9ykWKkq/hYFm3EptZNdZnSXHDakKnUqSYBJvlbYdc
GlwL93wP43+r68ZHF/1M4KApUeyFOBuodmymyR6bAy7/Y2ZYrz6WW/YLMtBmi32Ol1cyidFuuFwy
AdogFHnchG8iTAPkHFSEFdX1eYYmuESL+fNUOp3XkBvEeTc1tZvXNVn2Cue3NKTwJABlYp1zLom2
6++TTTQ0KixEW8+OThp6V8atnqlSw7qjsIcyucpUFpQp+iDXCwPGe8GeGNkXN4cGzLll6FrtOBq7
OEy03C9dcJHiJRqdnKd4hP4vQensRp7CFJ4IEca/luBz4T6KHg3k/f7WcAdpbiMSjoqU2oYQKCB9
WtCxmOJUZS5xZaiEC7nCY2d52ELWrx4v6CJYM5iSOAsXqxa+rWjkVK53M18LUdPXhuy8/k9BlZ1h
N/RpiMRF9MRHgSF6n061oaMM4/pyeR3E8pEIGI294o/+a4znd/1d1dYGSuHkjGy5Q5wTBDFRw8Sd
uVhy9HQnCqjV/WWt9l54TZBLcbUqf7zXdxUlXzlmYivelQzP7V8AARw+NzjNIY9vN1VFyaehC3Dn
M3C083mjq0nPAnuNS7gUHH50/y/Wdj7ivrVE2Cn0PWIflxICN7ZRRFID/6ff5aDoldGdAEtpWI1y
lPHJ2kJZN7h4uaxVvsy/RafYGjSa9UgaurPeHstXhr0UZV+L93BRpCX7u/bMojnASW53la9lq51F
s5We4ovqrmZcm0jvA1lothTi8a9ySPsiHvXbE5N/MDsMCdy+kTFWQ+fGyCHUoI8tnL+LjyDVaXUw
lu1pe+Z/GL6AQCitGE/CJLu86Ej9sateWUF5pSRkdfzfQnFtH+zJMvQiP4O5wn1f5IK+QaQEG/Sh
f5WSI3YlUA63hkXZ2ivNcKFJcBdesoCuffSm2JxhyPMcEl9lN2WSnWvBn9W7gFr/oh3eq2XbJFcX
uQ/qRx2/4orTZiQhaL70Lnz+KSw8BK3xNoZwG6aqBUPV9AtV0rPwueWfHX/MkUl5haWo7TMsLWNg
ZU3yhKpXELtvPRg8spkyaTo4m+D8GKEY8aqldkMnBoZIe8BfS89JJ/3q8gmmbAisnfR63cbJFPJ1
1WYO3fqjxLd9pUp1kBR8y96fp1IZ1bh21t9PhDdBFsZL2G0t0rYhGTKfHcFnH6Wciiji/7Y3zHSk
37br/DiVhNUwFGjNBgmMQS5QtU9DnqLue1XtkxPCS5SJpU6MMTbOC7i6BixMkC0ERUxowyXlXLGb
Z9pGuaGFLXKoLNvmf0AjagFFHkIOWzoiunTecdYdUBimj1vTu8LGEDA1mwYHLdcHr75FcTVsasgq
lCGrsEQk4tpldVELwxQcIA2kWL1MbofCR/1vJsEEe2SIyDnUoFIMNi4cdpmPd0f5djmDjlSAGM+h
q6LImvpo+NmNiA04un54gin0M9qNQO4Za2V29GoEqCJu5R83iLobsJCzEJBpeL3UvWONLkgai2py
b/cY9DNVUHHmG56BC/fThr0g84GhtYxoAIxpsyoq53T/bsR2jZYTGE+a+h8sJw8bhZs+Z7OutzQ6
uwrmOUKqzcmJlJTOpCOO6X2/y0ZMsOT1Df7a/DXB0zveeMgwkGVm72FVrHgNuJtNi5GoCKlEZ6lB
17VgxFEqZpLbJ9PC4KCb8NpPEgVkAgzC9RxokydZB41uA0ky2hXCW38pZjE/6VdPfKwbLayhh6tt
W48p9pIwTqCiUdvQB7yif0bg87PGfsKFqZjQKWNFapW1fwMPMcOwCoTfMQgg9M6RXbRlGVXJzSmf
bqVIMbpWnOZVGg6Hy01wR0cCG0CcyaIQrJHVlFz0txYKr3jaDBzZpG19xs0vWPM47LyvXZTORj4w
SQPY784OvwWW3H1ftFlY9O4rxocQhpW4e2uA5fD0tVQjqWs1+agDb8zyp7MIPuq6G7mbWMUOUDXY
fPJXdAhx07QQi9r/DlO7rqM49Q0hpZQ9bbFoi3BO8vZJ3iCDyq3AJ/TYl3Ou8tDR8wAuvEW/VF6y
L16XdXHk/RRSnTDpMpnaWVbv3F8ozHQwSq/M8KQ65fvdLRypkpYxmPjUKUon+rTbEJDvcwXQE64X
TnhjkxBs3oRT0LHOy/BsHi1sLFMVHIvK3WtRvAWf4rlL3IDHSm+iHgtgGIIQSKOkbl1uatMrAAgi
YgKUc/bpOEgQQ4Gpl36Rj+U4ow1EfwIrPK5B/F1ntobdOfizmmFHHp71wtvsCzFoI+TvlkdBX+IP
m8pzCC6KIgJbTpq+IhcCEjbbh5jlmXsCddwc2NvDRSavKynV4rG44xhbZ0sXS9NVZ7MbBMG+4e+G
uSVTifu/UGpIVnGrich1ZnJ9UIwSTouiMhi0zi5qR8YbsVCR2mpQj8o6ZvbeaCHIxMeHM20qdlSa
QuPwXwk8cC35J7wC35OYUIOruCFXUyB9KqdmB7qNqofwDaIeSTgraBVoH7Y81jsN5kwqKgLDawFp
ysfC3Z2j+vPnDYkEq0M6BOnDNUcv+VqS6z6jd3AIjkVNIRlyFIGV86Oe34ToKgk+AGKuqTgxjpsI
wM05GpKFye9XEqrY9SWgP8xgGhGs9SfX5O61S0tIt1X6e5ET+tr1/7DwT2203/8AYpVD61VG11ZD
kHvXJiScleIE8eK3rH+cMnBRIS8YiFjOW1o5jA2EcJXvAP1NeNfDNAxzrOI7VuvkDdtQcr8dZqrP
8nMCfSW1v4EOIMsbhQlRKnIj73lnk5kS+eNCkcqn0Al5t/PzkSBYZJjNKWrjMafqbayQhyK7uxuo
ca6Ih0aC9hbH2f6qiVAJZP/wYc6EwPmGdr2z02HKPHi1kCCHveBNIxrrpyuDLuFq/r1+143tUxIT
IEhxP/u9equjikRsAkor4J9T7bjHjNXtiF8EJOUbwHgsNpEk9sztwdqqz1OSP2Y8f0plpoFrB1KV
TRmN6lBS8fhjLPAuv04JaINazx7UALAyMCXC9eWvmeOXHknqJleKzEQkBxvyai249033lKE62xuR
VcKqzRhrdVFH0jwbmGxUeMi4/GRdslS5W4/ANpW+sMog8fUPmoA4+Y49vRlUMAVmXDRuw42oinNp
ilUKDr1/ncv3sbKBxt7lTVeTlyESw5zULgqoUoOHOqAyItk9xyi3Y2ECBE5XlimzZ5/godSAAUfn
yXov2QFpE1ROrJbGenSymuag04rJW4l8FRR6MdvBom5JH5bWzi9WNWDvuhRNlIOd6Q2xIm7uNkZf
hX/uJwFytRQIPX9V8lWmOTvEGWpILMjQpSAqg2qjMEzqSGRsd9qCCcsSzJ83/AcPmyAyPMYN35sj
kndakD2bC5MhLgv2aOYNnPBLmatW8XMyX/qtoVctSuERjSWai80o2Qyq+JbiB76LJ1H0Zkv80bjU
MBVpcrN19e11HaUQwV6sBJQa/Pebu5a8PiusEqbwwmH8gSsPQB7R3Pm5VrAjtV5qpv8uOt7BfLWl
U+iJPjS3h/5KwFSOE99Y4EJWpYzPgi9AV1kOJODpcSygyBVtd/CG4hTQYyPjRsTXQKs1XKS4R25h
UBCZnEZGCXi1+uLAm4z6f295t0TZOtIcJ2rcSA8a3BBj0n1zFol65sbB31tS+Yu71/7WDyMtioKA
IGxzBlBz5To6Idc+96Pww9XGqkJYLB0zMojP/KRKVqTsJWGS8jhxysd3KQh/eFleorPymkIWvHFu
Ifu5VfZnonYvKWiXE3uu90yR/m1iqdpMWBRUcfc6O/uIVUjmnRrxvB64n/Cl4LgytVD/GnXbiVFT
QRsHvajTVDsQJkGT60c7njV2NyYK886MOLhiGKAx+6fQt5aAWbiuDz8CiZSl9Xeuw1xCnTpqxfvl
AARmuIGzNK6oqT5MGlKMT7KHx0bDeTXNSG4G8AcdBlmDyxeXDPV1rO/AWt4CV5H/+SGn+HRJ0fbm
snipYbYUSfYWoZqx0yczN3zvvirQnuCFZbs0snH4UwUkZPBQyKaGL1+CXDeDqMZt7D/6R+mWgGa4
i5fFY1OMko8P0HE7zt70AVxb4nXP9JE+cU0Ij6DN+PanAX2/eL15JEDMG9/BL1uX+eOwfkqv/lxB
xVTbu5DRETcU11biMdt3xAteaSftdgeI2QmlJrgVRakKlrr3g9f3CQUP9YMfpDunlyoObj6Kxco9
XgvCPic9MsSkNlipnmwCsaaFz9zKfJE5e/liVMcDEje+fGEbGFNkATCyLy+YvaxAtg7LWjqqX1Vm
TDEIX+zKJm0ocLFmEHMfXTHMfSwly1nQ70kJjp1bGIC6apeHlTkkKVFlwX4WDzmxFmOLdQZWhOGY
GSAzhmQP+fcTkm5BX66g6llSY460y6726OPEANnbRRmd1GtmWW3URIXcggrxKWrkgc5fXFjMGAZQ
6xRm3yVtONr9pZp+Jt5O5j4uKm1gNm/fk7lW0/0oqHvWgBzDxhXPbqM4j1wOQzzzR1heqG+7SQa9
wJ/0hCpGxl6nfRNkLakdi3iOuSevUwy8uDaGs2zTEbQHEWffdBrdGl3HkKWoVMPUZm+GKwLm4Uia
GHoz+SbOBablttxGxtIaLFmYaTK6VKLC/W/dfwndfJmf1Ls+XW17qO1A89VyiLY21gD9fwQu2oo4
v6bzJq3yyPBmhp0SQQGTPzFOY55k9PFyAhoCR04T8maUyqMtBJ0LyR6EQ6mV3IKPbkfpSFxwyOCa
7D0IdtxC4aA84IEd6wpbDXO85VOsmwboelrbfKe/qdZpkrlXByojNa5BBVz1WWxswJCW78nPFv8m
Vgd+DwEmN+/7ka57Wzpr0NdHFvUPLf0OAWSsgrtHTXGGkyLZAo8Z3QieRZjtDv5IZAIKf0SIuX3o
QuD1yLURd4IOqXJ4QVYihW0hpy9gnzlK58EX51/u8skDlXsXSQY+JeA4LTt1GhPBb4F6q9jofoem
WBVVHuW8t1At++e6msIZZQe6jYou3tcLoz+aYKsFi/JsoBTYeIA1CQgya0I0lrzO0aMrpqlpG6V9
2CKBV4o0rCMFKAP1LTDQJKV3dPfkSXanbVvPp/22tMUcGO7thv9GiSZymNi6nXm81Kx0CAA9ggFU
ZOHIdbI2iDQ9PeZ1gnww7Yqn/wkzKaNeqA7jIcZQtRNEBviWabDfxUu1VRd3pPJE7KeyfeNtkcFa
97GUnJP0pgTc6PjRPffWETtm8Lv7AUhUDfugNS2ofclwz9FfMlz91HVlzP/b9qAenslGdhHxwN5x
W8H1oDcxBBxYZ59Ehcy4zyPUiKh9LE9yyKfguUUwh31JAceLFbKgCka4KUowrQbDYYTwZPtwhljt
Rf8aPoofh5x3iCUj4hehn62rwQsz0VlhkXm7KMIKrGcnHjM1wYFg+L+lx3L5dLthtiKQYDxlNh0S
eZ+4ir7SBK8xjQAQxb36ZeC3yOXCmq4XwgCkRFKU5Leo+0ZohuFvlTCK6nN4SiIEGtWTY6/1lYUp
qEej+bnVcCAxW4uyZTEaTVeKEmRHCgT8GcrN/8m2Z1yB+YBpzIC8iwLq6Hm4ueGSq22HE235wMX4
GTVv2K7+JI0fMeaMR2D2zXg/+mlqEow4WIYDWzmIcIZbOSvmhCAVGjAJfAY4Wz/YDYOiA0GVkzk8
0keVM7fp50FHWCk4lf71Z5DQLSXQD0Im8I2YjaB6SuZU0V1XK16IYDtdU6ytE7fLFWdWgYXlEmMR
X721DKXaFqzGLda8yHZ5FpiMtBdY1oS5SF8FrvYP4fbb1FfqDfno6mhDA7Nzt8uuulOvmMrvisTa
AlaVD5UKv0cGqtx4QT6BsjCcp/zZaySW3Jp0fCZ9HPKoXUATlacK760kJ8rqmjCsh5Q5Z8o6uF2o
teEuV+/Tjf5H1DJvYIOWg6HLi7IFNfCJqMVsTfGjz15Ejzm1kUluco6qNWqDInUa/lOUaOVAgfPw
+NtnCD1OGTfVq/70E2A0M8/z8YXgTjV6ETgCnMoLtwuziutkFMfZe50rFf3VldQStVow108Y1QKD
dfJJD69PAdwbdNOjhAyMF55pMtesal9yNDU4bDaO13+vnngWazz7xvm1SlY/Q0W7t6Gh5d25j2Pz
rjrdMbY/86ATSr+j+GYNzsW25957GUvXcLauYn5y2hkwzjYhIJjfmc9ssMRKOMNj6msXZ29NBWdl
dxlDw7vhvHGaYaG8ReFIL7RTlIWm917IMwmtBgBl7zWHOnOeyvwsaAZZY6AxRCxMBlTtOcAmOMo1
GRrpQdMqZ6HOs5bnnGh2LNqAGO87ipi3NxvBNfGR7thjEbA1vq7IYcVzvUy2Z7RgdjWbP3DzSOxG
vtpvRqYO7u77U91Bn+fY0Rzx5oIPUU/ICW6VDvdrcj+Dj+yl9tRErxAsi1eNd6km6oC8aZr3Na8v
+GnQmxOVYwH8GEMir8xWHMR4uTY1rYZmRR+AmfJ5r6aQ6H7CLAowPSXuSkqRpoAEqWu5NBOpeV+0
ma1zgOnQCN9rVppr8/IAvwz8qWFLyUIt++3Fk+kgX3PEpNsX1jn732o2+xCaV1ESOIuY1Zsl3fNT
foNfXu35lzf4JVFRpWUpPibxgJuaMWnQgmZWXTJwxGI6oK94/PARQgVEigGlderRtcoLhz7JxhCU
8SrAX9tZKK60KV9iqoQ5UruVoGOGxc+KH2gldzLOd4lxzx6X01Opd1a8jOpMSwMREKifmyt3K/YY
kyo+anx1GOza6i78xQYo77X4KtbwsygFJfgQJP5bVBgGhSUnOG9XwYuzBO5eA4y6vFmEz2KjDOgh
u+I3zJVQBelDOlcUwmOxZJVm2yhynJkrHkmYp2cNmlqGZOzz5hxIsiCevW1O2UQH2Aav8rIzy11C
9bB3O8YDksso31zh67pnw2CY5swZ2loegy9sFhczRevcC6/MWY8wTy5xfOmvEf7/IhabDvA+oRm2
x7tkfw8eTjFuOM8QjkNRHVXPy9+huWGj4p/71+V2/yiJXVvWWNuTZxkzxuIoQIwQN4x3r9ylmHV6
Ll10c/+663PF89XtgJ2ZBHk3GOWa/e5YgOdOgUh7AkWttIWL6PvhO06Pq7exXPu6EU+CDiBX2VtN
N965pFIm5l6AzcYZjxN8arwf+lLq4KnSTcUulMgEYeNETMy0NaLVqhvoc15AWOsAK0Ir2ozkgx+j
VD5vCgtpr3a4QL3J3xkG/cbCApAL3oF39to8y6NvJMME3cpe9xL5L+fYN5tuagNo4F8ipdFoEPCp
40nO1PAYqVe/uDEvh9kQD2yApoxrEkgFIATdCzoNH3EdYBKTxC/8ni9NKcuqtdRVgjCcG7PsXOlp
57QrSkMn6VjqyEUhgwhmX7cQcujiuKI4UODGga1yx0EzADNH+A+BWUP32q04hPbNChXaHdGlbZe6
W1QuhHX+/VY6iYL4JzQmegCz/rtobEzsyRIBvBqsfY8zZkG7ZFuXGP/zpZng4tfyPKBk+RIiXVLc
dt98IA8I48zAFscCzd9HCa9+D6b5ooMIJKC2XP8g/ojtVSVYprLQfZdtl+AiqEucMbpwKBunXjXl
12lBIXqo+q4a10nZ8WRpie728hkmYwdrLJW7ihF6dmChmmKpeWOnDGAMStZodzLr1R8J9EoVRj0V
XNnVhJo5xb2b5cv7zHE0XxFBYwmAg02+ZPZ2+OGVwvHOq31dxwXdxH7GAGO64WNOY20QgBumZHir
njL7pBlkAnixGZlfcWq4ipCkhoJ8p0KDQckHzVUMuRWpXR8GNQ2cLZLvcUxqU6fVu8vP33yFA48w
qcttEbkr+ThEk6lla/hM21aLVPaB9Icfm3neZQ57/LDy5O5kn4j16HQl6OZvU5e2AoUBjRAKIc+A
Ys72HwXLLJaTjXEak+8juS7xT2wQokqF9QAsOn7pPn+QHaHdfGS7eTwJ8lV7iX9F8g6EUq/h97Nl
ZCVg1PRAf3LRh8FfCCcg/pG956+DmxFQCUn2zATBuW7a/ZKVLUPlnXzB3MhvL0w1+OGA4znakdGj
PLeBOvSCuMXGvMs0lbHMHAFTsnmCVqewShWcX00j+fKBC6ZnrtoGLHLMDjStyl9G0RCou0qEbapP
8C2sUVXRakNNJX4Sbw4/6daoPe/WYX+mCTS7ohnPJfGQrQYsT5On/9ERazxAYW0yDPETXnsgE+qN
Sb27s9J+UssImTd94x9JETNmWOQAYC8J3SECAllP1LtRw2pvcGYfx9vhQvY43R9y8CO6NLhM4xZV
UsCI1Gt+6FRmSWBWikeROdWirVb3OQGIJgIvLSJ03rAERoFBmKZiay3q/eXxgREtXaP4dMaoathc
nx6P/5cPHq528+MpOeKy8osZNTAExSmmsxnp1Ah4tmT7Jc2XO1MvAh/R0hYPfvMmpeqmws5O/SRR
VFj4r7Br2KMpDGgS1kGaplBeZiRIDr7jiA3VbRrNcY4wZ/asJ8o8VvMvuwzbPHg7WoNOJgQy4T7Q
2EcNxm2lXbWtyaN6dMFiLjVh7/ptUm+9wmFbP1X8YxvWNqJ2NO/xXi2tca6J0eOss1j+6J7mPtC+
uwuFiYzOsPfbgP+f09SUmWEGCp9vkcy2WA5FQooA5fCiL+EgLW8VrsVdmXiG+ZpX4UE6unomIl0H
Xth3JH9uSnf46IBZvca+FyXpIfGF6StbtwtfqdUXADMyEHBC1m/QddDI6qzVBRvDBuphSMTOUakt
B+4TXxupyvPLvdrvEFLgy6EeM8k+LzPkte6tsx+MDATYAaf24NQz3cFtVy8M5ltUtvwsgEpKBkXr
w7emzbxH0tSN4s8aUY14yLH9zoamAFhXngn4PLbnGXFRK32yt1+53tUBpw8NP8bO/GV3NMYQIM/F
csPB7YsjtI4QxvvnnBAlzusAbirUda6UmOCyearmnPjRZv35ZLaUAz8CUNA0GcHFXvbZFTU+klYA
jhNaoIM7H8HjGbPJh3UHbzw04sSp2ec8LC4NYrdExEcePYayxtzY+PtT+Em/4s2vXeDWu8Tfa4UE
sMTHifDlCB/EiotqnxzZsRp8wF9gpngbGzkmB1CH9LNCTgTcUn9hq6Ff9bO/WBtq7fSQX2FSvjjY
DqUs4bmAaB7M5G2jz6G67VimLV4veWPvMckMsnP7erScPDIyCWu+dqiyZRZ3FQozpBd+2DE+2guE
3HxG3VtKtamx5w1ivbcQdHaCD+zgG/KOwwcOu02KxFPcKIi6shl6TQd16KlNHQ4n91WnSB3fwKom
DDZA3aW8CaxrXgtsASgn0g0cDKy4Z5HlUSzj4nrV4XR2+sIKc4YCXdCbL8B2dzzwkWOpVk9qDBWJ
DMETN1e71DzsotsexpQoo6Z5BdPSlrY3j5UpxvGfWhcPsLnGMPZ/VzqJOddNHGOS82VX9qmo87vc
5dEIwtkkIogt4DqEaVVeGhE77eUjfBdchR/rR0svZ3kzX7Ge7Ec0xKvgWe7msFbDubp2C1X5rz3f
vd8hzLNMwZ6g/fkASCQj6e7VEkW8q9rVbbzaFLBfET6xTY+DWyVXf/rZXadAIG27wrE92Q0CdDJR
ThX8WZTlS4CmvAurcgQ5Z6VVdFgBgM+aUD3c1qqFYHddKyosWvjmbrannN8kAatekK8Ezb+Vm0el
VYSxZk8PiK/tnMg0NGq4MbwcP6g3ZwAgxvhl+C/Etmd1y6Ikc8goWRkpyRVl1qAS0WyEovfF3lOu
FzCpO7BdPfqVqI9zSOvyUtL8oO9o4KUeq3FKtA3jc98Y1aRjvMUf/Zf50AcxvbabjOVaplknHTnc
ra15q6f2nyHCVhJ8sF0mVXcEdwIvHE5c8qjEAOHmeJrf9rrpCpFkzSK6nAprnbkcZTLg29wbwjTM
L+CttdzVg9mMQ/Y87ndRC8Red2E+fy2yF9f0q5nV+hNIeYOn+gp+StDFugeCyUXLCCSFGQ8qxFYy
YpVqvozp/ZxQA7HqJ32RqAT0LWFLw/r0hzx/Y+sWKo1vZWICOI9ew7mPQtstIyNiaaelX/Ud1gJ0
LCpQZSSCGrPMZhNLaiy8p/rUlSo4s4Q2eypmu+23YKyOtmw9I4O5e49ruT5B6dLQwbknyd7edLcL
kmFIR+odpkiKhM/LOrtGeYMpKPpnC9T7mGD29AeFez/GdqXbl/kqjb5ZYlq4WLAsxLK7bMiEyind
wB0qRiMuH4qCsP2bwpJIJkLt+RtAtrLKtAjAYzilToEdS9V5p0ZYg5WDzCip+qFTJ2korp7F8YcY
sDo6RQHiJdwWqTjoUjLV9iivrB/BtNUspVkJpUjQBVPQPeHEY2p3WXJOZDDmpHa1UvbYLtw/QW9I
SIagEWGCxXqKTdU/JtB0oYj5UyNOfcNOVX5uo/Cf4C7kK9uI1bEAOG+H+rxCXHYOsI2ItJ2qEOrd
QtbM+Hy4UK++aq26dOGY72rWMc665bimP24p9YCbYNR+h9y0P+ayMPvpP3f+OwFuxNTCSGVu7q4s
GpOdZR33gbJ8ZxQv3FJuRQtWD+4hAPKXUDvGod3d05K4VcsQQcJZIUm1+6yABSJP4/u008ZLImsM
p/FqVNnTWob1WkAad87bZD+ptgr9fXNi8AMVdue47nI0MU9rreUaWf8vrLD/ulVeQdD/j7XLzg0X
0tE/NaczCkgZ8PasgjxswXSHfBWeW+EEeut05Copja+2nvIKomRVuCNQu7KZ/h9hpbMp9AZ11fVp
mw4EYO/M52CpsgcM9CMdclxrE5yTeip7VyiHsx8EUzk/gCjl4nZjYeDDxlXW1IVP37N+THLs6x4b
Xg4OUqZMeGdrPMYie0LXWhB5v3l4PWWPZN6w1hAfEmhuwy0clwwtAYM2Cr8Srm2zEYY9E52om23s
GrWiQpx/W/IJkLy+hYKKZIvxiRdavol5Exmv1Jzk6FgcB8r51yHco+N1m3tN89pM5rjF2xtp9MXK
VACgiUJmtoGCQaRMxas/VmwSr6V0aDYg2BGzZARxndIdRH7rhqQnRm19D0+zeqYaaISssqwT+pcO
NmwrNEcFln9Q3uaSyyh+LNLuQwcGZ+CP3v2YoM5JqnOJg5a6KJrB5O1wrgveWuZK21WLJjkEJbQ+
bxrmpUDUlocGH9oImfb/t7VElir6m3EO+T80ZocNmuc38gNwrPh0YfKlOOGmM84+7gIER/glQ3Gc
mG6U4xVB8sr8Vu/XSm1qHO353xgZAfKAx4hZwspVy1D3yqbDZ/EULPM67W1Mn1/BlT9CEgLpIjRU
Y6LwZEjP99fKL/wlvvivwxO9RIEN3awFdTErgTLtwzT8dh2qw+NyfOkvF48Jk51+sQZwkoXgWrH1
PIYIa7DJDUZb6jjs8U84i8ko0IQwGOZY4lzflf0YLSSPYC98gUhzOAN4P+7n/xtT5JXAG1SzIbKX
BXYwKYtJ5Jr9U8ylbRTK6urWQMJsLEdy0NO4b16rOY3TRGd94EZGqFZKfLK2rmXTtnKYr8gH05gC
YlPTmJp4I89gqWYz2yjr5edJrlPYgh84pNl0KTfPyiQ1UQotvIqNZo4VgYOpiSrHesPAKGxeCDv8
plcktG5nVJKhDcOCspFv0LApmCcbkkUP61uQXkeBztOxHZLAFocLmUbpyybB2e/gtLtKWcn5ti/R
NrXYtCFz/OfqY1BqsewZAy9KDUIm9q84e+dZEvQZnd4jGVbl1VoNZ/rSVqAKjEOsnr8Br2649Wec
ys7tbxUmB/mY0SdcgHbCBoGEO84tgAdjzWwtZu0Qiv6MsvN//OS2A2O8OA+woVhrAzBuLy/xyf0i
Q7g9WwAtakXMld39oIytkrJIoUMTswAn7lUJQx8qBVH8W7Y2FeoY/jKtP65qrPhU2+P9h0X32dNf
r+6lC291pOb4EEZfP4XksQi8jojZ5RLPPYqHIA7Ndn91+lfd6gr6iY/cpsu/Fcy8CnreC1cyrS4Q
jSoeZxuRzl9lL3nY+k/qU+ug0Np37Z6C44gFDYLf5Kh9e3pVRnB6A1INMHnt17CmK7XS4Oduw+aQ
p2pvDPdGss633gzHMlDWYxRdd4vnEpob84RkwkOh0Vdj+hBZW17sftcSwnDSwncbAFq6V6cQfY2J
OGULOxsDyrtNMHxtUTIq9eYzeYfzhC5wF9K4WbcD3hz3I1NzGA7md9zrJhkr0NWSo2AnsxHNbxGz
oceAyBpPfahiEwIYt5SDXM+W5n+bQmkWODE7bXqz2LcOwEQjXGUuIgOXnylgD8Ti1ExF+3sSkFtp
kT3vxA9/VW8ZkJ/0mK0Z1OPWWL7Fta9Udq58E9IZ/hg9H+H5y6eDJnkoRpU7y96+KM8KZIljKJUx
lCjBdG2T4ZGZdsd+olc5KMbMaSAvovSPh4vvOVaEct5GsbT7h9ayZ/Cynr/TM15d2sKQzlZCyICW
AKuXFfPakAe5+sO7wyHgKg4CqH/dlhErgHJK3EJDYFu7rP3YTC6AS7ADNWm7dor2X3y3CrvPEtG7
pTnir77r1Wk3JCHDXhBdAi6Nu5aiG2Ysqif8Naei8PJujaDMLVi6idAi/8P7SlS68BPTFt5ZEQJy
pNKn3ujafyLERQA+xG+Su8yROKRWaiGXhSUZCmrrp0umAni6FV173Rt4hfwwWuJW8c6g1tEBrrtM
tKOLWpYqsTRCSNkTmb4lQ7WAQHUjwDzwG4orWGJp+QV0Xc1+rNYuymBa600D7Y14SkNJoIU7AZRv
heXdAzJjDVeDFH/uP46gjxdSEZSOf4uUC7cWljdcSQpxrd4AtxejMwCfzmGMhbyiACtBjxKyoJq/
R5mAPrg02dj3udFz8+QLANx4+Mw+R+78cGPhDv0l692gAWWTgDSoyTl1O3QC4Wb+xj99BvrnZycj
Kk1gmLKG6zlL/aYQXlK0Ww1WpqOGwbH/PU3CzA9bjTBBFxXVguV7QmFwMTytWIFyiIselOgcEuBR
bY26Ccn3ST2itcJbpcW75aoC+VybwMTE0U6dFaLqLYl4jxbwRXdsuph0H4OLCVBEsKXpZo7mxcBQ
eyLyjcrtxHp4Fz785DAl6q3vi5btFQSUhBaz1bpyJ/vicmydPx87D0H98N8zvoFPnLO12sjUsQ48
vUdTitVI6OfMQv4YzctAAd3JQrYscen1O21/tMsXGotuQeg9A5ukrr4+qQPk2gNbM7jP0vUqecYU
i+h+TSbYHxVjU3auGHm22l2cDaVo38EDANkMqFTiAs/koII4RkrD2wO4gk3WRa+JvIKU0NFlDxfn
xI6frRfzib7vw725BjXd0pPqOJOlFr8BodPaPRTjhpOQsONtcUPdiewaxw8pshz/xtTBZynrVQmz
xFTWFSuKXrmOYHl2Z3gOpCvv+BWKneJAOt6ajeZdmQN+8DSXwyFZ2z3uz8MKU1SL+yQoB2oLWRnQ
CzIq4/M1mAXpCykt1MATG2aMFkysbGraiwwSrvX9AICDJapmkFRSxis/f507kubWaA4U6jUBJmol
MG63UORxjmUUOileWGSqhmriucCd8dIImoudYdgmooZhgyEHHu1R+p6J/7fYiHyQZFN3HRazi5Q6
4fxeP6OOSYm+IP0o6cKt4u4TlgKS0NoqSP00t2n7AYODw75QSB+MzPab14zgM+arxc+jPA2mUCQi
54P0qXC52+ObglkJmSmmS57Ny7VCe1OAYXpGBcu4Iy32y7fEKphvvzD480lGKpuSpTulCGZwt2CN
Fea5PuHwX0Frz9vcRxgovECtuEjN+Pm1ytXnH9CKpPd7Zr2NhV7E6hjIzTDBz8+grUarSNu6/NY8
c3tKaxoZJ25DT3YA8L0uczgaz8iW4/xtt905kJ2k/g32Vf55783S80rkAzL13yUNTQUZsHWR9saT
9ktvbNE3PvB49rEJjb3fDx8mt3U5qyomFGIeKcN5B119SZ37t8c6w0nKtSzoKPYLXcDJIKp96dt+
2fjnNitEPZgGXu0DsQciMKYqc6/XekfD29sLengvEXMeYQyOSWFMe8oEYb80Pgzd6qF1TUMyHp8Z
0YT9LGlBvbq1pr4HwDQLXXLSovJN4KmzMFND8WaRtwkP1TTOHi7JhlRFc2qsmZEeV3Buk+8b+/W/
zhrpBgDzjv8N48RLE3SWz/+q6bTWs+NI7sgORha2akw64ausDTglEV+rt890r1dxNKeYH5F6Vk7M
jgrrA74Hf43aFG352WG3aRttmARU6HFhZbnBEMRHN8r7VydKqF5OtNScMrPIcKA8fF7vIoF4aUDg
wsSpSnzul7lUZ3MPgupyavUXPq/siulz8wKiHs7Sy6uYUpoJgW1EDSzbajMVa2d1LVRSjBl/xHiH
5dYozQpVx7LFoM6t5J19VWECx+/8j8Gbz6qhP5jGbA7t5/1jctSY/v7yH0tyf9HY8MsSVSLeewNK
e6zf/m59F/9YU6hTDRRLQ2wXsLqVPl7tyv0hDie9IMKDxSHFPT4E0tR7Qhf0pWH0aYpEfbc5ffwz
DOPUPNKJT6WP+zyuW2lOI4nQBaPdFg8wg4tc9Vdffv3iG0l+gcRrXtAMUpl2RABqnoN6lqxDZpUx
Fg2/akbC2JN5C6010gau5OmwjKRX7RvXlco+mA6K3WkHuEVDCjM5AT7fn6M3PtWt80g5skENJ9lW
u1kMcn7clRvisWEZuooR5LV9NLvKu6A+3NLihrXx714cp7C94aONw2j38FwdIZ1ylcnqOqJIvyat
ZiEtFkdzddOHCYgQr2Wxua8zb9VnnqkIcKBLfBwkE+rdn42qLmIhgmHHLLgLvTVApr3Gjx08w1gR
3qAYI4NEZTQZgCFItT58h/Q9H72+0BGOLdFiYSxGMfPiARbKFePBdrIEwa6xpuzoA6fskYPdlT3q
YTNwKN00Pf7sfM/kknUkhWNBoVacKAKMwsPQgx07wYasz75N6sJHAoFWNAdkaCJGTlfpwuWYE0QD
dQvVfy+Cnq1rLI6QYnsd6G32QdMQMfAgWcfQ8I/KXAjmEFiDIruqxCDi20py1jgoHcB2qH86DLZY
/KH3AXHhEeAqy75Ygo7wzqwkowAvqk6S/ivbzHsPbFudZTvxdpps84qoSl0OyRR8pxDGlwkxVam0
NM6VZeK/hR4TUdlBbpxAjnxMcHS1yMUTUyM2YBrxciyXJhJ/S5d4mE3ffSEo0bxN6qBEouB8l8Cm
rPNbdMZzgX1azMRe3vJu2pXXB+Abg3sRGfpNibK29+7doUs7p5KsWjSrlB0E1eqllBkCc0/Hp7bn
NeUHIr/ODMvkX0iJ5a/3yo/LriEVwqsAiXPNSCKlKsi7RbVh4Qd8QGqpMDXIv4S+npZnpFwEANIL
K21e3IXMzSTkbwCtVF5sQDO85QqkFzaz8PDU0tWbu+wD5oCryVZspppPqqwHEdiG10Cts2XchdD/
ywqkb1YnsvrzJuvYgdpd0KYBWNHS04kJmCB/4gYc9YC7HVsXQmIqA4fxBpcdLMzPSXZSEk0pRF/f
IoOgdjMPn/UfctQH9U7JTS8mMUcwp/FAKF6M71FMXGeGv+3eM1vxsGJZDbMnyCpPmSsk0rnMX8cU
xjcRLT215mFo1K6mH3GLq2MEuzpdDb+zmKVN/LTFAvBI4nK+bMkUUDmjVchD2qTujcIEzEaNsQRf
my7CQr/JPIuQ7P6fdlVdpWb6dPYEJfURKe2cS2b5mlT1052K+bqTny1deLrwoypAXsVCSX5ylSzB
0H4DBDxebMynXUqP0/Kr6kyAs5JPv+LOQAS2QIhEdq0GaaAfd1I0u1H4lzcMiC3QuR/HBWM4NARH
SlowOViMMVTlDmR4qe9PRc9nXjwSoYw8e9MER8mxV+FVMxOFf4w6pBvWW8wBahND95WMNL8xZ1tv
kgESOzpWklSlfqtM9OKjO8SyhoiQ4DYYACDizM1NRl6I/4QXpVcPz09P6SNZfQiR8b1hOVbza7dU
zuRNNp0g51llWRiSToGZatIKirOG3Wu0HsmJLOQQ5Oc7VrXhl3ekg1l4xXDdWKtoE24rRemfaBni
afJij7th+N5nlMf609mV0CjAcDbz32BF8L/xW6J5l963J91s4fUVK1U49IBGfHxHlHv7jc3js2z4
nfkLjFV1gW5Mu68M1d0QzygQtcqCIknaJMx96T7tzfAAMnGW47AHFWCzMqoHoCJqek57YrhdLGY3
CSxDeKKPPMKzJCplFgByrGljgAFwz9FYKpvPzvrYhIC+DsSLL5iVRkDrJC+rKPDaha+efpSlHHhJ
b5gTCpw3yYp9JSjUdn85dDUkqKLr8W4329VMvZ4PkegexO0pUxsNVi+3Z0ov3cA2tODz2f9k0dqU
komxSSiBFAW8evU31s7VDdP69jmgbu+5m+HlrhLeGFHbYFqKzZ+b2Aqd8NF40DNL7m+Gfi8U1iTR
yatjbSGagMFMOWRRzpgQHZIgqKaYXvs1DpxHHc8lqkqn0m024qck3IiYHwh3TV8UZhci8UJMG9Nj
PDJdxMiNEVMHxnlgoTVN6LGXsLFrdXSwl4i+sh1N9nIzM7mnIsbmWWxK2/2bhmPAnt1g+zbzzII1
jk2wwyw6Rv32/L8b4ldxBgkb+f76IlwtpI09uLcT2h3zZMunseswN2+/+hKuIoyizlwk9Cgr5RyT
EhfYm/0TFGWtasssh4Ua6u7voczpgkQaayR0X04rpxpQtMzUBJS3LxavaLLQXYYuATiqa9UDqXxP
9ylt50afxs6M1LsjfqseZSjrwlDNb1aLip1HK1yU+X1vkw5Q0BKV+sdqgXgrhrqzWKTnR6k0sPUD
jkrFxRhN61OS+/GYu1G2CrpcLi5ceNF3cz96N5kq0LCCCcvZo37AeEjN2yHTrLTKZ/b8R11V8scq
enBaQvzQkUmuCs9ozQqmYE2AIP+d+oD1F45UwjpwUooU8o98fBS7my+25PM6ZHZqppM+w6Sl36Bq
FhDr2Pa9ZVF64bIIUY0dj0EvGUm2xWj6jAR5arcXq3cYZmtnI2M21fqxiMC+DD6yUyu9w2gR95iF
DjNzMUF6o+LD65ENbm/mDes763ew8LfLVjQKbO/fbCf0M8Vb/KrUkiOvUfwLdGesd/iUSTyGD4LK
ta/KUq1WyE3ym/Pmqs29MPbbub/EncKeOJZVqM/bAmEC5PQ5TXr9VNmKJAPLCzY05acDvNeIVGeo
55RJ96z9mJi2+nLoM+IyL0XH0TDsWifUCJUd+rgb74m5MuBQTO68HnGA/Sq2eLGlT+yOrg7Tkt/P
CrvxfTfGX5hCIxL4lTIFGQYP38DXxbXJrnXwbnNpeYR1U/1lOUaI8VZOow5I6YFGBB+ec3m2Fu0t
qZ42eCbvtDi+OQ7rEIqDIrLG8K+QTcuvLqZXWoBUzx9Tv7Mr17tAc7u7viHsRHlxi5fqnTTc8+Ke
FMJIefEqwQNetPQL7eGzBtDX2/JlmSDxIJEBGofLiwpzi7yClQV/OA37OFc8MNaBaYI913ulnmHb
thk0hduqoIzsF9gZKZF4eh8BzQnUltiZDcXJTE+FETfdb/tHtbTjmi+sXgWb1rtboISc9sjIf4dV
7+We+gW23XMslLqJLRT3WKFbl70vTsVpDMxb9HjERY11u4GsMutGCf+9iOY34Wf4/9aTqSZmxEYp
yLHRHYCxMhgkU5XFGAaHWVk7QGLG1/aRzvBlKB0OicbwfPm0bMu6sAhvGXPw2tQYw+ToY3uamCA9
arlkpWjUg0VurZytW0atQcK5f+nzW5SS/rGPNNhuJ/phoaJ6ykP8Lp2ari7Bhc0cbMQrhq1vFP+u
Bng62DBjyDR0Lz8sRaVSe4GmbqMIxEBFzSaHSJd2YJ4LBp2q0xXm4ht4x2HYnZlxi1klxg/kqZ6X
q6HYEE3gfeJFRmtMgyMwUE5lZK9xjy+a+IPdUxbb5zlxNPsECoq00grE+yUrpuuEp8zdAe3NRA9i
BeMWfF1Y5i0LD8zKoXRpK4XZS+c7K00zSdO2LqWB2E+Us/xnm+sx3D20qmc/5nhiUI++5YdQUUJR
wYI0O7x477Fv7q9DnEbLPfY4FMe85j6GG3KVblbXqReBGNVnE39AGE1UbC63AXM7MUV8rj/PFch1
DfP3jnr5N75nZ51iqUe37sqZwJ1dY0AsgFkaiIdILJQ0KwvFt4bonpxwdYHNBOgQ7MeYpUTyYO9S
RWbdPId5SncRZzTmTRIy+wAwKOhvJ+MAElwIrokfjMUSHoYLZ1Zs9MwQPUI+llcQ7KiKyrsYNlP2
hO6sAWU4jtR9IKRME8YEnHWfDIMWMsh/oHm05raaeJP+MdwZN3gtkA9VJ21iIJBjXNc4FXAOrhY/
vhu4ScuM4maRAftrak3bHRwMIFqqRbAjub+p9jMmeFcY/05pUNCVNayUZz7NawBHbMjZBODKcQzN
ZhaRG2aiFOjTfFv5Ql+JP8ukjbyr9LLu7tBilzrgIoh/lLVzbJcNVDgCzwHzVV0opl0IxuByriYg
xxjsgxngcAtmm0Ya+wzcdTNWE+8WQ237WYZD+RA9Yyi90P2ekoPsBC71kYbLM3dAGBluHg5O/neR
vDRLxx4VzYMEC1pCr1rcBLlq3lFtMu1+zPIBs5raAD4qKhIgmaYE+GTEQJRmoCeonwOQkvRJLCXw
g3m2R1ulT11FpkWXuDbLp11Cz2khVhgEBaq8jJPSokAlsFYzQKy7MX0oPSiaVnVKFSJ+Mio3zNAc
b8rkbAiLyAIUn5J/6vSGzoXDM7RURie3BjNnQLMln+6dctWF/k2yE3NUEptSc1YOPjO0BOIcIECj
Gz6bYkcqgkXv93cY8uO+8MrNKp9C0NEYLcsZMaBEREomBorFP9na8Bw4zweEdwOK0qK6675XHlYE
FFdg5DyCZ4eMD4HJNdEcwN6X9T8vNLYVYDkL58MpzEM1o2YKl5mLqu9/PzhMoA5pj7PXOzB3CF2i
G5wRW94s7aVyyGj7wKfFlw9gvH7TSKdBLY/8qOc6HQNixDYaDHtBTzLr89xTYYYWyDyII7O7dv52
1hT1fetQDzdJnNatBpQolx1tQm3Xd7oHflDbsym26uXLmX6fIZ1ZRqK/hyZTOScbi/682tRfbEqG
36R1HZY4/7r83hXmMNM1QwEA4sFeP80ANS6ynjltffvjD/vF8KmhjSBsD+rAq+i1AyECsuqDa30e
sSLEsOgb8TywMo8sKFNsVtt9ym2X9izny7Q7Msusa2PBbbkXI7fS77ccXVn6uQy54liPAnBYlGcI
xn7KZGAyX6n++aU2OHMlimVqbkE/Yc2q2///U730lIZWqEp/YEqhtTL7XJ1+unK84tRH/1FSbDb2
YwIGD3U4fLVB82hzu7GeBHgDWCKfYeoMWWsCP7VhmpCxLDKCKkvPyLSIMMM2RCglFn40viUUU42f
VzMprMC7+OaB6bCcNO2PZI4CaZPe0av6uk5VRRspUdYDQNa+8xQyx/g45BJmDg87qCTawGE8UJNq
KKXtTxma3zhogWHkRI8w4Qclq87LGx6wtyWTf8da/FJuy8Hf7S2iJX/Yp7+vI9IOir1phWAklf90
mPZID2V4u+ByQ/PDtXnPnnJEayG2D8fovyZ1repoczjPlUk5SBsMEIV+xZlnec1dR5GXW6/fv7VX
HXRyJcKMhYoU60sGIJsoLT3uUIu6USkiHZSbY4ztJFcrRzKkOg18yqz8HMcsL4uZDo5mjY6cAWL7
Y80iG7v1zzZjXPAZ2qGhtlLgGXJIRnE+hlAlG1lN6vnb7IUITRUOC81jsbN3xTiStt8wdmZX4tt/
h32On0VOsCBIdZdEVtAh21GrAOOXE/bnxDk+9CxBr+hRbUHAtkUGc//RUV51SSzWrMHMFe6ui41O
5rlJr4L0IGboTwwqiqTRJrSriiAm/haCPCRhNac5SFWYbKt3+z3v72TETXLQ35TeU+5xNkD0m5uw
yjBRMX3SOAtM52Bu0tDMr1dP7dgOACs+NKbtKS8u8kEqr15LGmZfITozUHA+LB6ig+gJJ3GBiMHJ
lJzRGq1/jmRUBiIaWLhRHC0G/xlJhq/1SZSgGtZg8E0ufMIa+2O3BhbuSMzSE7uLkUyGODguR4TX
RLUy6sbqoizAfmI2NgdeOiLIDLqhnrI5TLrC+hvJK55YhQ81awxU0YQlrRyNSPu/aEkkreQ7VFF/
tsompAU5BIQb6fkrzGsTeDIh6ZUlWRazM8qSufTpLFvicgoZxclHCfGtGnDqX/p8/KA+Ty3feELt
izYLvzVHYnJOmPaQtSrYDWfkzGTLBokdpI7nKKKUjzl8hD8+S+h1LyyV1vOehvJrLrw39Z0ISzQd
WN58Z3ASP7nvu47xPIEDx1dlvUnWhWsCzswnTy+Y4ZxRQYmHzMok571C6hGW5QPNUrsiQiTQTc6d
aiJlsz8yhNEL20zIug/6d9YcAZ61ZXOhYYeGi/EYafB92p1orcBbW0lC6Bzl6EXLWzvkFMxW5dL3
C+ruv7jzCEZgFCqhZfyfV/SQ34kOxvHXgGA0m8gdHbiem5hpYO0YOxXJeNaCHGCJOBBxKW0bP0ID
KW1pv9PDSKWBrAWHlF+WNa1GuAWfM6mgFWI+ULLxa11yZNVDJ/bdlWNwsczHbRwfrCZa5MFgk3sg
m7aFwQWnvndXI57Rk1sGerQqQ7ueYe8h6yJX53vRWQCI+I+8bgMnzJmaN51TPQRR3eKAZRExHcDT
gWAODbcxaj3HYEQ/gA7noln/eSNzAxdWYTT7ZT///62NT6brQ8RXau0ZLsVtQmzzz11Z86pM39k2
IPU1dNhPrzZ2DoGVtINMdjPsncbtWaFtEiXXtIwydIHyL5c7bdWCmAiojPqtaB46RcfB6lUc8ytX
J3qewb889jJ635MrP/iQ2gdCggxPO3CZnYPzA9haKbYR+pyJaJvtDPCO3reRamOmNQcG8bULbkUD
ZQJYnL4YtevEas6DY1wDWvATdgm1fLjtLSUfTaGEBVXxdjRTMF/WRv2KHNn6r+KbUyRhttgzk9ci
jixQsKysHfx7sC0pS5EOXg9rrrz24XHiTJ1+s0isJ5apDuKPmzsG47PQng23ApL8R3TsDrptxUZ7
c6um1AtQ2PfMtQLFtziYj20Kk6U8MCZn4UInhMQLtmNAj7jHfyMeUAmSEaWkY8LpcpfZ/hi15uGG
kI1bM0CMxqHztLzHy/+m1jTuagkV+r+qBwWTU/p0kKiZi4aHPyaFGVrMiA0/IgM4hMGiPbyNwdBX
DNsvTRzEKypi+h8cwb2nbUMyoOWfmP7EYnte7euA3oX9FG0RmsgoMNb61SIZ7nviQMFQIK0+b+sx
SnWp1Kt9n7gZgBZ7mR/BgByCGIl4w1KE1DXqDHCIn1xL+j3a2NuqnPQdeTCuEQRTSPSsvyev6UmF
H1ZZ/z/+UEszDvI6XaOn+m2HS43sqeSNCUtz5Vz4qPbTcXdV9/0OcP8fuGlE6BnfsoEeKIx8kbmk
fkFFZVGlvZRocXYWFb6K1PX+d45AmAQg+md6an2PodYy639ssMhW7Sym0lxAZbCNicqhDKuMeOX6
kRNhubTpgtQDMjBkLeK21XoLIvGZwGHQyfjlxOa/xX7Lmmpk7xANLhgVhOaLoMr6ePPDDnJnocnm
0NuyCNsa1X2U1pynKELWA99QR41XP2SIfTCmM68UILr5gERsvA9gNzdVDXYqA3Bfteuh1HiaeCHg
1ABdIMjdlRy9v02rTbzWwnZjvn7EuQYlx3lv1Q1EdMzneigDEunJiIbTAzjzl27BfGM5Ut//2bjx
jceavvH5whf7Ah/E4z0QbKSk3ABva7uEzklrAX6Wi7jkAgvp+QOYhIHKYiBovxVCc6CRKIHV+SjY
1btOsD4kFcZ5nQY8w5e+TOw1nQD8UvzKMP7dMzMxznBDBMfnW5+H+vjpOAbaYep0b8LPt/tD2UIm
Yi9/E+b/2+3ABG8szRbPxgBnKqBwqD2VdHsvMg2+GDEV0pBL1A6MwHSoV9CU8tL07lMVaB9DIPZ4
KS8jmSjG4m7pw5iV1IFPknm0PJHQsLC+0oATOk+OZKSEI4PBNexfH8ax7/rxMbfONMRz+ql1P5zw
p1kqK0YQQ7IlEPX52JeDl5TJ1Gix4zTmdq0pHE55lkpy6O8DVwvgeIb3BVJJI7EAGp6DOAVA50qg
qQxHK0bg3c1VCEWFiSHw1TmxP7M9voyZ2janZmhqsCnKU0KkPqQAL5puV0+63Vu2DMxFIRufwG1V
2DnlNCfmcbouD9i+Pp4JdSdCYfyfC4FSroAUB6Gw/EhoUUgsuY76iLdeIOhf5sIaPnOLDKiA9hqQ
Yq/ZnkxKPpalR2/Nw+MgJaDfQjauQcf+zwQbkJUkbWWYt3kSBHVaGL8TbY0J+Dv6U3KyHBRX7ypF
l3G0dfbPbNcyxGsY1gBdprvIWAxksoU6BzEUuM1clELhHC0SV9FWqlDHkNLgS/0Wd4j0HrZwr0AP
U6JZeZrGe1TI8K3+2QHF19OFAp1U0tMEl0biFsHDkJ1nyNjEoYPkDm/rfmfMentR8Cneh0cQoi8V
45u0GMcJwd94yLdNLRGWnHMZmZ8m3K7fA3RwrcVFgUWqfUlZjyfgVZQE8dJ6pgQuggow8MUK4yqf
L/peXJTFPZWCeEz2sHgYZYcV1Q0ZNnJ9i5gQFSCLad3Q7T6CSwQw2xDbbGacYdnpkDu3qJMG3s7Z
6glGljsC52hi+FCRYPV/tA5M1bncsGidWnBQbzEo43xtUod6mbjoeUv0xsZ36dTWEjZQjjjp+Qys
m4/5vXTw+n16Nn/lZKv8B5WSIzVcRN7jaoJ3/c/Dy1E7wA7DmLEEk0v0ri3rBqUr50KNbEly7+KU
NL2farTC9y4sXkOwYlopmfrz9CqauA636DWKPysEH7okzuASMoh1hpInZ8d+iUiGtziQ+LehLmHx
q+w7Bq7oiq7cjm4y7GtxSLp+topG2jGmiOq9XrN4ZOrq/Ig6bz7J1DqhShbRvw0NeEJroX2zVsOo
AOPtT1ua+alAxoRU5Z7vRYuWIcgPjhzhHu25joi9UOfvk3JbQzRBM6KE0rZA2BjHbBwyPSbh0liJ
c4eetfGrxa7wzdrmHCjy4pyr95VHWR3UNSfdKxauYYQjhSbiyTyb/ZgsuqU3OWqZkVPK2/cXGGEw
A2RTzBsodPmnup40n8eVUxgE/nEj8YK2H7CGb90r3sGHe8UVWw7nE8OFghWrJAD6kDKFli+6SLcB
vSKh3vNWVqUIQAIZA1EaYVAxgdhWlmBBJ1xYciSx1Aim+v/2gLF+sUzUsBIEeCm5z6ksNDt1ODAp
zxX2SJm3IZq4/IUlUDRzI4YGcmfNxXY0QbU6pGjQTWsENzt7RI1mxjDfxOJHYWvoUVY+qHOXdATl
Uo/DQDH2I8PbdJh+FPm/Xcj8V/+P6hOyFjH7DZFtPinyhrZnSWnMAiGd5kx4McF0dlAVSfy8iztU
FO/OpsXvalVHU1cAhWxnK+HnHTYsbhJkKAFvFprmm3SSYUV+U+XY0ZjKOilECuNPOPmoe/pUIr9F
1dGUbauRYCdWmkUOHUIppjbzyXOE7+Y5fnqMU+7lcQZFsfItDqwTLobv7BazxtF6/d13M7hTwRkl
L4YdIVWJtwYiSEe34PP6UxY1ea1Qf8WcjojCfaQc2VGGWs3ZnobWO1KfhPAg9yzzqvH6el2EngNG
8/bGvP28+m39T1cGLjCKF0Unv1EvqiD7ZbpfkrBb95BgfJl6cqiZV3jc4Po8cCNLJ+zeILzLfS6U
NP5SPdYQy2GiyFaQ6m4UojKwJssiND3jsmwj9kZrk97/LBuvtdWqaguVjbuRZbrfwDMngApAsJSQ
IYtRjyDQ6Ws98KeX9r1TcNLJOp10ggaK7sedkn4ap/gkpVRQRa75iQ6fiaheH2RhIEBG9DN6I6xt
MO4ZO+3LiE2oJKW3qs6Ari1ajxm7sZV4fdflRTlBQ0a0LJiWE17Mcq+2Y3X33UI/VI52qLEY1p3l
fneBxfekzZsYsCbxDjVASy8wRBBCIjGNh2Hjyssz8PdD7BEeIkjFIcAovINWmxFwoMtp+czITI6y
/U4fpb28qX7X/nKrxhwt6Lgpv5nC0Lpr8/iFmbs/ZXLeBJHkyUJGh07h1yPFM4RBOtA99iLgbYkC
pe36L3KHQb70gnopVJNAQlEHEolknv8aZ7kyi24pSRIxB2KBwYZ4IBDubWq4iT1JBxrl7tgUCleN
wUrnOrX6M+jXtcE+WkZJfW+S3r6QYl7MDKiBt7aG6dxI4cAAOauhqx/zXdmJUH5Dh+HOxpthv+zL
f0GhNCV/gdvaxl/IpBpn9Sqhqw8E7GrMaTgd4tW8icPmUdxHf0+f/kPtZmW+KL0bZFWx2RxBpW4S
SYQqGsF+nobfyqowMeLo9EKvXaSuoacOuHROosgb39LIaAdDHBplGG5boE3iALXObu24e/KUJFbT
S0wczSTrL9ZcuWLX1jnybFbfswScnVBFswzoGFgfSSD1iqm0AhH5Cydv3jJmVc/3hZo/ryJKeUN2
kHspNWehXd9Fze2NW9A+Vai5mnWmhBQ2/jregptijR0czQ0y5aFh77gkCGVzK29oBWDAWzjxnI9+
U56Ke2Z8VMe8T30af/HpIhdvKTI6/iCfKRtpl5TUJLTsObC7XNEf2RsCiIFm+q9PcAEPbfjhLUgQ
liA/ibeez6ObWuWJL1XEnMKEHYQpS8MaAWFt2x3NneEjZOPs3p326gwfx1T1VVOXlStGGUlXyz8B
yUYFQWuR8yL4UNoMWZQnD7A5dJ1BGiZp5QI7VKvo8c2Er4Ru2lnlqk/gBr9rf5cjQJ3e5eVIBbJ3
QyrsQeUbneNRFLCTrFRamRKoHsCvdP1ZTrjfR3I2YLCvMfj0b0Ubvp5VDvKvn7X9STo588BnH77S
Syqi3GKAjR8B8L/Kc64YF61Pr72QdLVoMKqx01bJLHZYN7IA+V8UiGniL1mO0WrjBTlieYZlMEtu
H9KsVvddKoWFF0uHLEvQxhPWfeU6IaHxy+5R2wDxe4dsRG0KA24dfpDADDESNZEhPFhYjHFLIdz0
660iGOlyQVHbIhrqchDcpNLZEsk/Y/aUFRZnoMZAxNw+e6eJ967FFWmXqd7etXAEJxihd992ymzt
/pFDrJftNGIZ+Yc/GLeWbmo2EYdmVVQfx5lsvV1JrzNcvuVm8s8buk/NB5HmLOHmTsKrv11cH3C8
lDdsNnSDRSAdsPpbxzvk5txFfWGt+R1Mr3NKouRw9l1oRnm0idebi5q8DNFzgeafEXsaw81QQMG3
zg+atlSKPiLIuKypfytpxdvTUhGDbZhC1YiRFCwSDmc2KHGQLcAaCiCbnyd51e91RbvKncHzgaFk
N/UIgcL156f3XMbKmJZ+K419TqwEXYu5DLBkwlZJ2JUveuhFgLAWgkUyrXAEWzqeBs0dDOqABitQ
Z5z0xOxrztLMGC7rfY6XcpYyY+kQgYTALkaW5J7DmBsZqI1cLsaI81ZBysmtYERrXYs4THNV3F9R
r1+Ov/qT7YsJzoyjY02xZtscFX9Ixn35YeAyeisXThJe3X6RPRE0HoFXu7xZaEjwcKk+0L8bfELD
/UkS1NWOz8/yiQcGkpzeFzdcEf46wBIIQqvHzyx5bE/Z9F3M+OKBrp2tc/6lnRuA5tF8hCOPOkTm
Hey2VFHikHwID0Z9gIbDPL/dR/wyQN+AxV0ODaLMS/SNg6FrYVu3iLgeSV9q3DCRbUyqJK3vWKEy
qUBLyiG4cmqqrvS0q3jpEWc2+TkEspW16v9fMl0y0wpfBi3ZWju+pWBr1cgVdXY9bSfKIVeNPmsM
7hZb5rW/i5Ec6wGKbKBtbSH8+WeXQpLBd2RPqkwxtcAbZash6qgIxwWM1KTGemsrBRBGExn+kM28
P5lOxZOj3/UayjXaW1HQI38vsmjezfM/jZ7iaJuNA7glW9N7KjFU4919WJxJYlaUtlreb2uas+Bh
LVFQzHw2//pPV6/z0tD+fkpDjETvk8Y+r+gU/PHhy5bitDtywKb6iaBHCI3UncmUGdnIa08QDGxe
yCCQlbNyYL3t+7YMZdrOLKC6K9vjcTGiI2Qczyr4ccRVlouVWUhomS3fHGbeiSEPrt35/Wne1wMT
MVYBt8/ygF0Uo9RLPzapAbbYx7AisFYoEfpu+/rjlIfOgNIBJH+NQyV5F/Xt7ADbVFndp8cFXaaU
Obx8M5hAb8S+TDLemFZoL00P49LXSGonYn19+WlSi+JQ0pqcWqUu5DuVY/zXYApi/3p1VFQbWc3s
fwCK7E5VcDKge83MRxvWYkN/H5hXVXmm9jzJ0eHRBKrSdMX+1IGumkE8XiUylFECDCvTdBaVZUjn
L5QpNnh/RacdcARFxtKKfDLMOu9xWqqUyUx70kN895WJ8EwUiu4Z55svTxoY30B+Fk6W4dX4kFq9
ObmN8csGQCZbGMIAwbViAi6/ClSI+5elNST/TJR4AxydcZUSqPJfiqvOFETBQVamgw18nqLEC+4O
k1aRKc7vR+i29FYEKMcm/bm8zY16n6MaTu4ycNj6RHdUYmLG5rbEXG1BHUCnoaObxsIbnIDKHQKX
57d+/ZonffUdbp6kBl0FxmBtvBqr9fAbzts8DGkZ1V5FzZUeZVrZEekHkPnFg5dNQN1ovAPMiOo+
sDz03lhRoq8s2nm0OSUOknJk0gACEUjypBfec/WD9qLWcUOEGMg6e/vOZl3rbJHFSLyc70ilX0zS
QnZMGx3F5QYwL63Zwc2w7irQmXVJSEwuV8pfGwNYnDRzB4JvMXHaGSazGZzenafr3wJ8pHlHT8rr
g2fGMgJGYGbgu5MnPD51ZdLZ8qW7YwV0qgbv5MVntyt11+tR4o3g6c6KuAIHX3MUfm26fxpsSG53
QSgIRUfuIvsNQ9kNpVZ4RGxPiumQdR+TajfXvdOwPnZStN+RuCJ9kATJIcJR4I4FxYgGKaBs9gkI
+UppAoJYuGELjMZDlIrQFKE07thBvUwF8JxtdlTygaoqdCfUk5NwFGm/0QyhqC+0YbuSwjR5PEqj
PVHr/bZ8G7g/rJ3JhnzWUxXTOA7Kl7t8FiGV1o9/6Ax5qVGa6RLUinBkHSNYMRQ2qZSEhI1Z2rUT
GyWKCOLMXYibHTSzeM4KTj46kzipqRztDt3Nyx+URM1bdDvNZUiW+JtriSkdo91maGj/5AHCRrRU
Hy7eoQyAeoUQFevpgtT+INFOH1HVB7dort/PpnalJkJZak98/ezQaLWloF2SMsA66f9RrJT8a2qT
q80Uv/UEIENpSQouaba8MdcCykgoJ7wFchoT8qaTat2LS8ZXC1XTEXl1GnSXQw9ph9uQvZlTKjjJ
nTBwrlfqFACnF0carw8BLz0mw5zOzv8jS+GDy/WwXUe+l06fngcRnfvrwH7Xp2dbYnbdoLQQnvAK
sYwUEToEdM2RH3cK+le4xM29kxqWBuR0wdcZfMzzsann7F9KD78dbMOjjYvSamQc5NoA3FUIuZr4
uG3udMgx/Ah8TXRP80aqWiIZ0qHzWJ26r7DTewqMMKpu+jCKr9VkXXItg1pB6X8I0D5sLdDkbF7A
JGMD5s2BD7QksdXr73KrRIefF4TFBZEitKTHpZWCC8CXAAmg3FCu9qGQ1+OeDLN8Gr3qqlNHLXNf
mn7pCaPhGIHfHJyz5csKQNf0RXtNoAmNWU/+U5eeK6zlUDEQ9yopI2qyaySUh/Ziyxvw3afBfKD1
BOHn432HzqnbJNWnW4kAg+7mjuqT+kJyCsZSCjhFPO1L9InzJorLJJcX5/ZCLkdU/bymeDEvnqFk
3QcS72wT9uoLyLTY4RxYH5a0uDRNnpnWJs8ynCTbCuoekKSDyYNT2d2DP80UvFNhY6/kayKncT9R
+k77OfqNhws3Kd9MivJTlwkwSpYWDnjiZltl20Waz+6dLS0ovmgOXjtZDxpI+POcxTEO0KnVOOOf
ts7cjAdwnVz9o7IuO6YDtpNyI05x7bS0T38P080K+p8zIpzwyaORw2n4tYnJAY1GQPpmN2L1ciEu
MuWBS5yaB8qxx5FLxzLdW0kfP+uuuGTsV2mpPbGoZncL3OeDs9urntEGTkfzS/TTwpi8u1axJAkP
U1tuGqm2EpdM8DWD2bpJ28rmAmqa7137+bN/5wNDDfSP9yn7IpUA0HATTMjeJhExJvyih4VTRVyh
cut15LrVBpKaELYZas92/PRDWjvdBYiqYRSTfENEIHlNPlRyrZ9p1dWwh5X9rMIMOFOgwlAQFDdV
fDboKXanjtEoWaAPyd+KpMUht1CWfjkAoth5/H99aepNMIx4LxUfL2u/4k4oounR00tgo2lxGOua
+qIkhNy8VjVXfMzA6LlTsHKm+5BUO72Bouqk9Ayd5yrfZlIrwiMsKrZIEGbmqidubL1PcjsnC7IY
V56T5bN0CBEQ9C2Vsp2PW8eFTsfdoc2ob4Mw/i8sbKiGboD7hR5GvsVhI+26VAXeZyAxY9R0cj5a
JWhcE9LYmhfJhKm3JWXkOEwW5VAtVfxguXmUYRUCDfr/PrpNBIMZi77rN5jXo+PDBtQMr+JK6XnG
gSyumdt/zFr0H6PrNStWbUAO7sCC4KRDFGER57+qJvAj5I/Cop4ANjn8JYl+n1umDz6npuVnnneI
PE6MfnJjbXxjPfB1TNNBkWhmcQLVknDzOANOh0Or/j9RdFVQ2pajwgzjEO4Ryv4VelAAchNRLkBH
OA/+R7/b04V7P1wvx3FpLfiicSvrBD0LD2oXlx4cp9HMol6Izyr3ah1ToYGL6D7LTm1jTiAPBDmi
OssTNM/ls1ieyYEugBpi0LJsGAboSezePBPti3+LPEwZ5RXH0QtRUK0ORvvB4+sYs31fpTK0kXEZ
N8s0r2XncoYRoWYPTCeOitV4Asx9BALvBZOxXqrSY0WiZMAhpGldaKoy5PogZtM5c7ni5iWwVd2v
UrVtW0CpboUSqqg1BNgVtGimIrE5+nGPOQ4WGsrR4yPA01BzymrmYLGHt1EW65z9AOdrFCuxwYIL
YAgdYK45wQkq3FSVKeCqi24e4/1WvL8Vp1Nk6SLpMQX40jibpYDLGTs9JAHBfqxmYGudtUFJeBkR
nZB+JsftovjB3OvzpsjduBq5GGWByr3kg6EnISthx8yYSiJPVQXjF5ukSfX9Fc0qXBOSYPJ/03oa
d050Y/UVkcdJcQeuXgenpt96nJrErk6TcaKWVHx9hlK6RdsdDjh/gpioHY8ExEn1tD7vYcTZdiGu
4jhfS4eb00xSj6qscuTwQCdGg1ciN6ZIoLqRkJrfAd8fO30HcpPxE81iqGoyA3ljSYnHUi6UadCM
1m2dUJfg/R+CHhlr1dRzLIXzNuBZulv6HVugCKRnvX7sIwW7Z83RBXQUAyRpFZnymTBGUMl0eZnm
SHXIgeiFoxO4eDVTearmATITNwK0bi4mWO3E4GUjZLJ/3JkC737wJqYmwgH8tjncx1vtqf/x6ciF
H/h/3vqXLhmSXO0GKqfn4w0+8cEDsgrmqZI5Un0Hehyhb7wb3supAraaFUq5BHBIX7+f342uSVfm
2zBhEaRPKbDZzU9RRhIpKCeaydecVRx/xl0oLOs1/sKaPzbkWsPARqLTv+DFWRAbjCJ3c4ZCW9vX
OqlVQy98QaASrp72h01A9R5M8NwGXxd1ilW0gnlhAvC4aHWLf6fz7ymIEfdZhjeB6FPQ4pIR2ONG
JvV6UI+Wbe2f3P5Ef08kt0MPNClD6w/czCxCnyUyhvgisKub9iKObnNfYX3QMSZtGI6lOqbdlLjO
OUWtzCoH+ZTr7mcAqVP0SnTRXSpNi3Za31CgsdB2PADPJc9NbrnMvaX9vv9o55xixvkPM4Fkjkn1
wp1ZrXP8iKP1zLn9tuvJTlr6qSrs5I/GtTv1tnHGIIlhMBDoxovKPFhhO2j7b9WYLkfIoXqAirQR
i/FAfpC+PO0lQ0NknU2+UVrdYbBwCKGTyroQaJsP8fz6hNS6QqZ0xbsmcsA38xMe+JaBkJ5T6Cok
+yHlwoxdx4O6eQbtp7PQ20012/CbNnHLfPFxVwHTTS3iv6N4tpK8b3Gs3QS7gxOpiPif2LhRt+Un
q9CQFBcG/ky5w5OraFT6vvhF5/WfHZqwGr+k/n1ou9fSojZkgXUJE75AP/H7r7IZyLGjPjmvE9JC
UmauKNTrO12sO/0H0FZaPtqOWCo/+rl8/zHrUpUf2qXfOhGCDDLij2G8Q5Rw7/SBgT17VOz6/4aN
r25SJucUke69xEmrStekGYuJ0xwfaqQ+2uhZWnsSMbSfkxnyBZiBt8jrmFOBMAJRMAN7yMeMwvUo
OmaBQs++FOyqSUajrHvIInaOAE2T7He73KiwRR8jmRKkekMjD0AJRL8oUmFfSLQ35NCs6qOR6y7U
gV/uOVaCOvH8Wc6pC6+6g+q/+caenXgBMTcl4JpGcL31RC/Z82xV4Y/vAFplsz+3S0STIePwh91m
6vZ/WI7DouIEoKRap98DVYRBJKERBFx1oFsGpBYxlyb3YEL3bK1ByjktTGxI0TFKUjj9pdTe4jvN
ThevV3cQAQFfkwNQZolo0Ugv3shhWbF+Habd/Je3EfPhEsF43vrGzMLD/2wO01uuXgM06Pvd8ynn
/S9+a9kbHg8om2jQNrQmGFUkrHN+utal6FxPTb6spDDl3KSCVzdtB+iZz0ol7rIgq3vbAl7dCdLC
3W8eOKla7Ga5v+K8G7wG7P/jD9uflUatdypzgz0Mcj6I+wKv4deBqJDCyRyOVJPAsWvEUSR238NK
zcUlaF0bpxYlSI/F8RVnBLezbfcBI/CysHnBi3f6M5Ypg8xFVNmulxJHgkV968hDwD05LmTA01+w
7gLu6Orr0SjDYeD8vWMRLdexBBoYar5V/8sdg94eW2FiSmRtNSx4bSsGYH0KVVd4YdDO5Dlmori9
hzaFy8wNZBpK6kzCdyALXVJoZt2/MRLB0NAroMi0u6clqfb6/AJUBmrcr+dbSNbPJkvPei3xHMPw
ThLQpeHFCijl86RDGglPrfCdPn2FWnD/V0qCtr3PaSVZpDXrbmZNmxZIoMySlY28aj2JquLhssih
9DsxSZvBtrnGLc/orpQnX6St9kMMJRFW77vyP1IPhE9EF3r2QIl1BlpK5dSjIu21omHsGro677t+
ZjEE0aAhiRpbhvcS0ngKmq8goELEC+VHLedFFmDTqmcezAx9ZlXpSgML3GxPLb4+/nN0pY8twZ8m
uyVtGTCKQ7MgWIHAeXi6wMErbtdqXirtBXoseymmJsvmtT/ChYIrTQvVO0jbWsZRQr2ftrHQXUQr
uNWfqy1/MLRa1fqDXefDlbACTEHlUSFYItLda6tyOs2Q64VCHZjsCbc6ASSyFsbAAhOnkHUCfDQZ
pngTRmFUoKW0ce+lRnXN2to7MGDPqo536Xm2f3aoEnkVuKqmNoFl90jLl7vVSlW280C1LqbNDmNj
7QKkaKHutwQ26bctL1DuVNCojSURkUuyZicHed5jvZ6acw4VQOOHf35J6NQYEMpSKPTje7cdq9Bu
DM/bV0AevFPHjR2hrJqD43Nunj9eLNkF/ikgHUGydhYN3/zsxvDSiwCiUYqkL0plnzkdipJ+scKU
VQmQZLMguIQsZlV7WQG8SZ9RPxbngTZSupd42KD91+DghOu3nlfkBAit1fkKsS0gGnskdyoqvKPE
2QpFaOt4o0JnVnQMjrFMaiFcZ5qSwsToy3wp+gfHW3EptUPd38uHF4wis198lG5h02KZF6DnBkqV
mayqMDSg13gRlEwGz4Vzr56EmkA6wSBAUgFQGSJQ1SwKM3H8i+6DwOY7Afmb1DbvliepiGTbnQJ0
RWR5Gg8MIT8+hBs9UMpJwg7aWEsxZRjY6fFYi5vjEV3xhp+y3+mxVXE+5UzB7KMqWI4a/Ia2F1hN
1JhJ6F3tHVYBZvBimdOQXdSrstI5eX0pH+OM7N25I6Z1SXYVlw9k8u8FjMx/qdU89w77CJc88QbN
5aFJOSHADoRdFA6lV769rs+JftTNqHgEVZu9HpCiFwwjLR0lKMgS6pdWEayi8qN5TpGm3/zQA5+d
Zne/2fL4Wd7HYf5GHMDOuV+zQuJ2HQzPpqjHjq0d/l2lHq2Y+iVb67DXC9gZUdmWzZUVtOWd8PiP
Su2durS+7Xos+7B0DICva68p48BSE5HeeZli3oHm0raTP6s1TPbUCgkFSoG+SCXV1lMMbxzKZhdE
onmxBP86bPuvhmAIftS7Uz1GrYC9ZhTsLTFh6EkL4Xnv5q+dSmrudCqIZFDkvLf8BKku2mQ1s00l
YIJ+f4PmFDfs8joZrS+z70SoCyGmAhsveOkWHURTyh5domnajJz7J+CoEHDCSm8Et3vU9rXl0V+h
wYX3hZpUjazrVaN1d4uldhRgBFnoQwDwZe6mbUTkUYzW/qmLXnPFVt5Cx+m/F7m3GgkpV9vpb7du
iBr6ODzh7ZeyWMtw8t9P2ZYWh8t4KUCU3ajaC9ViIAYVFyxZM4aZtF1knudkNEowmsLm2A+h53JU
6CHiY0iMlK1h36GKKPT2dHJx/6KF7TmWYs2cfQB9UQsowwT8D1c9cqDb4BmVuBefJsgV6pOxwJYG
gEswDg5H3RDc4YzLMCFIIxHkSZWe/XEH47aebBtTqIBRHgqewO5k6w0JxhSTlH5+4hZGGF4NutRi
+zSApCW9NK2YZnkq1oFzaVjTwV9rZCZ9/fOTe7KSkEZ4yBjCz3bvryNzNPMPqT12TIIFkucfR2DF
6lQs1FaLI/rEClmZY+0imUmY0i69uTz/VRSFngEBLvc0tuCQA2PrnLMYMRyDKHB4icIHadgPOgAH
ayQB2OffiJwxaUQhtZCEIzxoaaksog1RpMf7F/ub8Hhyj8Laj1A6x5qeABZPgwUMDtZg898PPbwz
Jnb9POeAx7VoP5lTg0YVd22p2o0dChHPLM0I1mV6HnPohkVby6kwQwt5j65ttzHH3Sew2erDvw55
/Gjxo5wuSexT7EHDV9M5u7wbieNoqZ8SbmZEvde4gAbQSX3rML66BQUIDFDVnH+8GitslWB/Jr5p
cmDuQWE77uIRIkDaa9p0xWspFWOyk6DLB/g1tX6kIG09QS0xCSQc+CEkjJi1S4vWPArvidx9jrdZ
TWXHg1R7D2aauPv0XVyim1m70HPDdz/KHEo7O6GfEhjnvmZduig587fwXqV/K+Q7dkDexl3F+s3L
29GmxLplmENc+/kp2EbnGv/xXsQHv60FA670/jBePFxnohtaZ6KFgoaJG5qkvwJTAPUomEvbQDVq
KoRSHgwSMBDT3v2I84YFXg9cvZ4zitVebRwxRsLJctCXgnUqnMU30ZHAAcpHdfCApvkqHvgPOTAt
G4SkYMR5jJSAoTmLeRokXryx5Z3Mz3NmD8k+/KjqvcHTEJvWF4MKaiPnPcvmhd2nbFejmwl5gpQI
qqo3bgRuqgpQeGP6mJfLGvG8ssAKrqOHcKf/xhBee64DwrCxxzMwJ4wmghGurAChlflSxdnXzEzp
K/RN1tQ6IZJdZoIcxR3EQSji8qxCmNzIo+Qe4lk1eMelLENmhTQsLw/S43OsV0GUiEmdZGWZhtpv
uYSqe0HqY4b69OhYd6lPRnUJRoKwL3Z8KDFj6HM9Q2J9NKug2XCmSbW+Md0WaLj10ahv5vX64Jeg
bT6pPvvHWgGWWpbrxkw6f8dLlMDkj1niXPsa9MMfkOuodZgA2k7rwYD+rngvmxMRHy2sT8JjihJN
pnIafmleO2ZWpCpQrDjJfQgIKsGXHxkGigoKmQI+dgmjRomBA1RUeNlNXmUR5AugUa6i2sAwfyk7
vgnC31e6wEWOyYqBqq+DqTYvd2csHlKZYbMMUpcTNCofHnjmEgktrY77m8hV9LdTrwtlHDNP6JzN
1QilLKw9Bv2hWHrqzeqPrk6vIN0PRyaHfbN1JFRawHeP1yi5XCC5WOR3p+dnTTefl62CR7Y7gunP
TQbKKAleOYlXZadn06rSmnJNeI1BwGfflZtS57t/ctdrLIJgO1kVo6snXIRksIIKK0HRFis983PK
DQaelvxfXOoPbz1irrRSzGesiY8nz5KybOpnbzBrgU9QuSvmeTqlNxQo9gXY9SH3fhsYFniCzuzq
0zZ5RoE56qiPoA+GLwvEKcYEfO9iKxtplY4Lc0CFVTpvSyOm+uK7oXJvxPeoXWuzZcYfelC7rBI3
X3mPy9m5zQhvpR+5XPmoOrqCBwm1VF//5Y4JGq3vEMlV5sQdk9A9eYg7bXD2UPVxUjb5BmxmqEhS
T9+b9KUOlqikHavmmxoPvokBjLdVSmybs6ZLpYdo4hraCuCzPQtsCgetzq1UF7KrG9JhjzZ6tggz
IefpyketWdTW+YUzkMsh2YULHaSbnFM8Vm7Rc/RSeDP2GX56s8E8FlYK6Bo1xvtC2e0aUgEGeeEd
L/2CBqj8ZieDo7t6EWm1tDrAlaXu5Y2F4K9cUj9JPk1CDXijPrCOgfQU/DTwxO1b9y/AJcV7gwVQ
l5hzAICXqUPNYbDwxmajgEp/zsm/H+4ScdTlvhtR4JXknCEGSuO78GXVCGfNeXdNxn6SKuUxb9Mw
5J/mKR2r6fxL35RL33xS+A4B4lXa/fGcqQghNNcTJxf6+EhRzsOkXBIDmm5pzU/aK9jEjO3oXv2C
9mQEjjG4LiZOJYb+0/vh+SiQdsKD9XyrD7axKUyt9w/JJRAJWMmbtTOMlynjEecWp++rBHJzDUed
rRWjm1rcrywauAavE1I3QB/QOxJ68gLZzYamdBqrWxIjfnFmN4GDtLa6Fsw44LMUsipOokDd+PiQ
9atRiFe46tAk0HspB5xU17wuMuq5MRmAXere+M5QwfEg1/cRscWe3kopZe0LiqAI1XY97hmHjRe5
hFgiLekHnhzuW6VSspxO/Qk66WiiV58q6PekjetyV+GFINFj5alOxsnccjU0yFUW4dQ2E3zhIvfF
7Cia4th4O8KEies7QyQp7iswu6dymipNwQopU4wp1h37V8+417HuKXg3gjKUBwGyuR951lZ3GzJV
Qkut7y3DflbpRoNXj4NGy//mYRpTnDgkNgtFXAVQcWb9JXQ9MXNpO6xVlpWKnMqlT3SRQisQo8SM
orSeq+x2OEPjB98jCCmp/GRolU5LY0j6e167vJU+udq4ctpzPhahcZ+LkuxeI4Lo7FKhxpK9mX4y
8HULCMAjszofsrMK/dI2XmuH74jeb/NcmPYHTTplmF28U6ClT+Jso8R4NKdfmw/eCtiAOX7gQcy9
5qA4fUgaE2A5CBej7SIlA/IHCUpB8a5+FCr+pvCNBq0vx9Qv3jWVoUC9Y5WkYEX0lXVKGSU7o7E1
fPhaWCug6IQR8ez/d9XvSRLzmYDhLSmoSCg+ejs71G1xWBRwO552bivhREiAZ03unsDhD6grIjSw
uQJJjNsN9I6RceQ6zIElI22sXZ9ZKMZLarNZ7kHvAbw/Cpt+vUJDop+7HsNA/dUnymVeWYzdDT9C
rouPT7Ku+2yaOMBkxZrK9Z4YY3ifOuyqWiujb0hTnQlWyP0xbA2jakpJVu4f5lkHjZAa/hqO+f8P
dHL+Qnhf432wgd75Ka+2cRE7s1r5N4HAScQLLysk40ctsVn93/dPT8JY5wG8XGibsZOX94BM/x9P
F4L1bFVtuWSeQ5SPF6IWKVbCS/m0pk8shEsjLh0mhKPh9UBlsZP0DCbz9JDpC/mUte6q1SYgim2Q
AU99fAVKm7iIL/YSC3slGyzmTPntxEYkCvZUXS84bnJp9aEZtrAzvMziBqQRHTTkku59bdlMzTrx
3HDpeWXzFGI/x/fe4xFKs49Loj1CNv0Sa0qVuePt2gGZVfI0O3ZadKQ4KnZiS7UsuSs0NmdZxgID
bPTDDeTxuwXPMUM1TNUfCWJUSDyc8fnXzKmWnx2QDYyDk3k39VGsrtbfb0evzY2Us7L+XCCDiSqp
fwgyTsOCDmJ7VJ4KrFz1L4QZhRvpwViXn7sA+t9VBG+Mcr5amaTEcZjlr32odZCqE8Wj3SjBi93N
jyAQj/94GnftOfyw4sB359zXZspzntZmdtUqFJBya3g+kHKnZm/ebFm45L/JxD9UyDQnNRNnAXU7
D69/IA3yCxvVwhjOa9oOVJaG8MeOnu7FsDW/xDDne7y5PZJwnUJhaJrEMX7GT3occbpzxywMxmu8
j2/RsNWDfCuh18hEVocZBCN/OzzvHNiEuuKOhtCBna+dZeq3VamaiylRUIueXGSde9SFnCDIqiW5
I4OydgAskU62ZbHeI7axeQCfz1Mr7SQulKlyIMWE7Y+4QzETujucqsnYVaAy1MuuKJZk6JF9AHX8
+1mnnVzjkqgy8S1dPRSVKxxV3gt8TGgLOUt5+2vWtj8gwM7AGd1iHBIIPI5LhM9Uw3D9QybE+EFd
EvK0/jm4aT/mwpkbaEJ9D/0mHBMhS+9I4cqzyCPoAz2cXd6dCUa7y1hVNK5HxEnuY5qaXncZaDt0
p1dSfu7hU08t1RTfT/osmCisyOVMmVHIPiUz4BQk7VPw8TrIgm0ZZe64priKrkgSDsARnBnLrTQc
XP/aV79wAKEOaz/xfA6jKyF0osHgwf0pQ/TESj9NVAxXcrldn6PVf7BjrmjLBHgFzVxZaV56H2/m
nPjgA2YaPGf5siAlKK0+idRPaXW6SQnce5m87zC/0/87PXHaxONplt8CIu+R6Xz4OwZGZNK/ljMV
7Nd8Xcv8IcCy67WHkKhkpK2/kHz9Q/ZrPScmpWwdpLKenD0N2kTw290RYpgS/w0SF6s3NhaIvvlV
kxaWQK9P9TbLn56OiDxkLVKv4VfI/XKhoVTKPM39l96hd5tW0dyVoelwLfBZR779CNJIs3U0JRcK
76fWJwNJnCc7kVN8942579D2DEFKnuGZf0JguYiQHjZhNi9B8rUHMF5Lg4Xgs3gfanyzIlWYGsZg
dFL4iZSanO8ejyJ4dvSP6oFSArTylkXEt+91ER+NFg7j259cGt4cdsPf96UrHXEJjcB93XFIpIij
ndeIgNYBdlo3RFgVemnvJedpRoEuhoX4D3Xtc5guookvDq0jm9C91fH/DR2J0m6N+Jrv9eZbMnWf
Qgu2F1NWul6eOJs0efG6C5nuy0gy3sds50CM642UN59bt1C+xlzh2Ez3Ik1cbRR0Fv6Uo/1VpmhF
4NSkGhUpWXrFQa/zdFglWWoj1lFEaEnz7+2M+YfzwEkcNtiLAdLOCIVTF1SsWifXGyjZYAyH8YWq
vdGgvogwjYsQ90LbWa3/9yKmgY3NCxSycq4wsO9d+s5nCWvqNuRRfqTtWlHikj2pUUlhFQ6fopuv
K4vElbi980e1rEUtOQQQBIpwkzAW5E7upDiiVPRWlX0TX55gr3ymh3L8cDnIJu6Pfr0+vhcJCvTn
NK+bhidrZD1mzQ5l2dMtw4ACYqEGS9g9rl0V9fqawF89JRDNaek0CYehdENHmBj1bXDsd4sS3zM+
M2KQLHsyDeKg/k99db1TBWtJL/LT+ErkB2F1JQt2/VQXtPbk2ZeGlpLuDvKnIE0Ogf0R/Ml3XX8U
mh2lf3Y2960cD4gZ2D7qPL+oBGzV5kFO4NiCgaCOsv/bM/nu0QCyqHuxDdjcV+GZJK/x+4mkiD9L
j2uVmpeQxCeKPJlbOY820f1GB2de8nK5gwhI0Ck/5qcL0H/ZAYkRMMiJrnqRgU7cEkVfpuU6H6Ab
7mMwB3p5eIxgbWLR9kXf9lBlwsEwpFYkm7enfMB7ROXYjxff2EihceHBsNpJgbmfbaVhiN40H/x8
FrV+tW+fovv92IR3JXl8FwXl45F8M8cJWKas0m124yKUYy4lTNBu5pWql4ElE+zk0dy8VyRPyxfi
Iq8ghm8yqvHfPAIXm98q4ovWAQZlBcm8DoGROF4ZXq9SnTDDJU0FSvtinzYsAmo4NT3atvbXGTaX
zxG5fqaBoq119G1IsFfufPlD50CgH45IoLYjzvoLMyYvLY6parC+Wr0ImXobmDgMKFN7jUA97O0z
PDVJBqLYAVtbSqu7ulBexdJJ/ZRWCWK2kYWRmS1R+JZ0+nJi4iwqmwB4ru081NSTUYOTP94rv3Tr
R5grRSiqQerrKjMZTnwzN9g+fB0whike2AmTuRaoGiki9Bs7UQKN4lmChRjx+Z5zGsoF2M6JPGcW
Rq+fyAGJHuvtDyAPDhM9bSpWFOpx5Yku2sRoGL8OkULZOUuZhAag0dHDL+PdKvR1j23jGLEHhzw7
kkD7ffsXuiaNVAmkXvRsjZcDQfIOQpQxQMmJ/6KGyCCc/XQDFHNumzxpzP8dEH819KcD6ZHnwE6c
fxZstDgwmBKr6fnArllNdr1e88hWAg4MAlRR6UMJdw703SF8nkW/xUmxd2H91ZJ9dCyh67fzUjfH
pGiLTJ0kkXQVMrFMXYyi5kABOOQ7W6//gQQi332dqE7OK07eKaYYeV+xjKzXJ1aODdkP38roTYfq
+sCC/yPhAxGJ3giAiNESKtKYOl6E3Tc+EHS8vJpm7StshRF2XLLlaKwfOmJpgdBARL37vU9QLYe8
6fEZx+FhuXs5U+TdHE+YIOrD2ipgQE+1T3TF/p1B+5q/jDKBagSFAmwR2L0u+vKZm7auBvFHF7l3
3J75vsWZ8eQMFA4KI7ruYBuXd3+OzXzd7vjf09XRJThS/KUJHF8PBT9A1+IaavXrBN5S1doC1Gj2
K8rwh94p2mCYtT74piaaRWxm3cE60XlWwgCDX4jJ0bY4eaAE5v2GfTDDxtO3Vztw77IjPft3tAoU
XASGVXCCBcRaus1jGFVpFUWxqtjaPvGLvWqnfNgKQTMnNIwrALUyGcyJn6LL4mi1g7MuG3xETkmb
ZUtPcr/EnDksZbPuoY+a7k01rGfozVQ4ifLnyYv80xPgvsodQ5EstanwNJroim9ZuS/LruVo2Zlo
znqbz6JHvxb8HIIYlYOMLEIMO2YP4A/MxHRjMVLuxSMPcHpuMgd8gWARuUrqFBEfUaWPEMzfg9tW
jGzKzd9Vn7w7ZjqNxOtoEkhW4jEkoRT2TAnLeveEmCUJ4vr9Jsp5Er3SdMU1OuvzVx0AfquKgDgD
78fxt6duda0tGOJPij3qKNVlcLmItDOwZcBgu+FHkqN+8pnMAx/T/iKLwkV/UUKpGDNPV56i6AFg
G44LIUZQ3sFCwdpORjG12OA6DdGWAF1jfQz9BCBTDJH2IAUJDdo5F3ruqXx0+kSUD2iNFRVnLmGo
eoTFIj0aFNbNcsdmjwTm6VgZBJFDpyedjtFpLcOj9CuXWndKiqK8YPKvRjc0S3ilHrii9mAJGlRy
mJBMnsJfUV6/MOUDDAyT4UujGoa0IufWw/jXcrKqy79hINYCWOqQ+mhAXESB1r32ZVb0B7V4Prwx
anT6PbcBqwl3a9aKMD7iUW2lpidSWkCqKkTWAgYyj6ecCCq6ST1rC2qfbbHss1AhHWVh0laO3lE6
BNQY7AODwQDozKl77uEGcMziDYMX0bnSbhsoaXi0TkWq5MlsIiiTpITeVDld73yyfriO8S0GDapq
nERXwesB6FsClx99qGvSNGIrOcG2RwpPsiT/sn4i2LA6eWp7KSLnfE5J/wKuGwA8X17a5CzYj92f
kNbHovBp22gmMC4ikeFBTEPcNKL5Pngu2Za+LWhlZTcDgVYu/9aY6zEbvF8Em5WWzeHrKQ5u12gV
OQ8KYETM4n3/pQU0he1Qmsc9rtp+ykaRXEf8RJKbhNaGHlLqXTIHSttlfkTt/4q2CH2wUsgkKM+H
vf5pbmsS1pnqHE+AbGXsHu3lvcoVTkepkKbBY4HfkSiPyNBVpMKgBggZV/DWJnB3yGBNsSXRs+fz
KD1PbwWi+HUBrFBzK++gCG4m0Da0tiIoXbrinnCSwJmsfdIzRHYIGBcRTBUrSCR6moeTq7cBdKT+
fld85w6P/qwJMMec2IULledQPVxtHgoMX/WbXoEWnPyjrjRaItLeAs9Qia4EtPeE0ge5lCA6ptMX
Rya1N2dnBBkdDI6uxlOX+cTBCx02iXTJUCJHEgYvG5Fqe2A6OFBEIVK0X6oPjnE3gXhGkOb3asd4
kHdYrJAxJ+BUUeajWnp7310YWesQKkffTcq0LGgAYR5NL5iO51+ERo8ayXIkJABY7goEiBHb7zzH
Ph7UzsZssWYTxM0h7pS0VX7EsE+H+madcVcDFKy0h+DIwzQyhO/gJt6i0vWHtz9Rgj2kOk38jBk9
Gbmc6UHuAP9jYtZdVbBAX7d8cfCMZTrVNNxD1eU9W/zoyiROtykNFM6WIXZqnksa+fKfF/slonSG
tNajx1dQ0KhE4Q/RmVi21A1VoZUALOQEMvBeCGThGdGWk5rkw8XFHk7durQzzj1wMqNQY6KFIjdq
ihyIQOcb+EN7OEBc1KAi0rRW3eVWT/MohNlLGUoN0y/8pEOVjFUGU3LGxIDL+o0WjGiwAtOMmFlS
LG2fwA++V3rDxoQL7xi1+aHQP6vdmke5utwpEtg7SszPmz4ZWTabrdZMPP5sf4d4LK2kmYaLZiee
1oZNVkB3w1dF0+Q0GJMSPExJoBu+aOlgRsM1CC8GqulsCtE6+p5kCBeND0lIROsk/v6DBHD59DFL
1hZ9Z70moA4xZV6W1Nveg/KYBmrQekIM1XRCntbm+x46SKisbL0QUaWUTq5/kb+IGcPOnlV09sT9
JNJitweYmHZ1i81Ye83Z+QDNtDiSyZAFKcpBZrqcjodZu9dClPs4L0T2E8tIyi2ARRSLWuTRpeis
5WJNmE8pte3Bl1XWpsO52+bOEMcw1BMpk2W900ayfeaYSLTycfH5/g/eXhUSqDmqAJLkr8h5qCv/
XwaA63/hj8aEoQH6NN3RyHaHVTrbQIN3j0QEfW9x6UFJ13IapuuyTxbaA1c2mu/X2TjHksgg7tvh
xk7Eza2/UI8USoDXZorJ5Hpwq8EDQyaOryl+tt7lL8om+vA2Ri+w5J9Vl3KZMD1ddgqlg75tocSM
b7JWZT3VSF+F2d2XYayVmmUoWJDwnh/dLqbN1DhkWhe0PTO7V+e7xkqc3Zn7K+TULvD36dHNrvnC
L/o/TkpPCQMvuLolVw6i8ShzLFcNLj+/25XJ5RESAp2iKPzzFyEQn4kHPL+5eCLAQEspxCKl1aEz
aQNkpHTWN1h6GFzCjs2cK8AUo8n5L6AzKq32f0y1We0XbE5IyNRyxoxrelbzI3QPqE6UcmHfDAEA
AVu6ce3oCbJkYHtWXqQdsueQhqMVAU9GNnMzQJlmYedcrDDwOa+nf7u0ImZ778YNXw3X+AC4X7tH
lP0B/IZBmOO9+zwDON9TrDx3WUUTCtuAGgnwGaEn3nwbCvTQ25E4dH2HRAa1nnF+szsNfNqmsk/T
pCWU3B/tj2fm/Xn01HKbaPZUVRAOVaoA1/opGHgXHoj4v2DeP79FefxZ+KSI5w+hMCR/uzSl7Vcm
5jNSjSqVzPaRHz7xYkeaSGvZPfAhzaLH4pKVYiA+JSHeLfjqcf3VHE/tb29HYSS1vXockbsp5bqm
19rBq61AmHNux1hLuKtUWubO10yibH7ybsLPx01WUbfHZj1FrzyLd8qvC/JKRCd1Pe3iZtF85ELj
U/mRtdMQ/XjJQlF4wZJvYKOs7b112FDRKvnob9kDN27yWvOk5NhUtZTByGjCcyto00EgzrRh7U3K
pXkTBYSIH1k55kCRRLnwVCcmOmGAAzNLnWI+PwlJNaXh0sQAsPe0F8m+ONwrYqo2L3WGzZNyRzZF
eH8w+pCivGhsO6ShrmatC3aMMQlH8NwtnlItmUe/WfkGcLVpCEkubpKEmHY3EDT7zHo7YH4m6wOt
KmcbZwMe5cWuPIdS55FezbSG1UoJZ4Hc4agekCwzP9fCeQcgdSdEc3uMOH4qldkM123/H14BVnqF
0QU2hzRa3behHfgT5vcmqyqdiaz2/CwLZ6lUkgNlzHwGqEUI5toAaceNyQ2tRVGPU99cd/ohzGV1
VSJIcbyISI2a4kzw+FiIEeM3rlE4DVwcp75K0UFv1akQOfTA8DaPMgKwckXom9sOHvz16uhYoxB0
ybzgkq+WYz70Lzt+91hupiDG/Q4Y4tBJZerBnRxXoUn3yqQJsokjg34fi0X6zo30oZ/NFWpcGaat
MJLneMyEMGNPSaRYFzcMbtBrUvjb6L5ojnBVTpYw8Oui4cfZ6fb3eqhpzKt/qiYqiK+r9nEZ3jI7
tjTwCHukV/qZ08M4GRwEXO3m/XV9pnsTzwDQFiI3dAeX1PmrhhebB12FzTI+60VTYNUZUqa7522m
omd7T+T5AEWvOQkvmCO4QA8iooJV34G90mqWxHaPlyNtHlInnG6cg8jBvX4cbnVi0TJQu1l2nbPL
Z6X+jiLJmlmWKs5apoTUT5A9DKJCkWe1R4J6vux3if84WpMOqvN5n9Z+Qvi9rFtOMpZ3w55q0TTW
XXxoYXsHqVjjuHiS8+BZ7jd+NFBJWg8AY4LcdMVdnxfIWw6E0iBzTw4zZzW3PnEy+U7Yf4VNJdoC
dL0y9f+TNADR+bVoq2F/x1+NEb9x6g5x4/JBC1S4vfCoR2Kv8gR7jUtX+qQqbq02G7BofdIl3Qvs
8bK/GUJcbv1LjkP6pFKFMWBm07mfuGHuuZZv6PjNx49xKIfMSOxbtehe3ua85CxMAfALYUERb+K3
oMO8T2THHPSAv5Moj/fgIuTj1lKw+yS/TKCntZoG94/R5mIQWNCVm0FG9sFxkmbBkFVTWRsJ1oFu
kR1F7s017uFhW2mnxd6CoGI3c0UO80Bkhr7MLAIGNeAUtQzSSLxGugMmfgYSWLAZEW/JRqNec6tE
B3MdkYwgXcxVZ1SHkXBqMnYxJDXniKp59BXy7SulacjwvaoJz/ozlMbJuwwgenGxCP3qvOGgWKkE
z0bDeUwyhV4FsrH8gbf2eavaIAxFmC8exnhpzDSf08PxcKM0wat/9gt6GctahrzQiV6GtSeGj9Yo
xs7q6W7FqiwmdDzcaVSg1cRLNxqTexBVm9HOMC5S6cH0s5ZJpXCGhczjiYFvHTd800MOI1M98bVG
12FytcZdotxmRytA6pK1Wd12CogsjvIOVBm92PB04Z2HksUhPGvwgh5meI+6EQzyWcZ+io3YQoY+
xFLP25owcJi4uThzmlSMGwsXvO33ZlIfMC1mO1TJqlfY95ugu0Ne+lglds/RiZRoWKLlkpOCzA9T
uskhqXVFwVyzjSooaAEvHb3BekACYOu8iTA1wckXbxo81iUMEsZZiHpvTMCzD1r/KyOFoPR3EsFt
xJwud+kw7BLpundGp17Lf+XXKhJ7EgvFedp7t344GbHHmC8k32CnMPkHcsMG6zIDS2lXUGDGGju6
jekDlYoWGrdVyrPXe7EzLeMb2R9sq0wIDoII8DD86kRgWApi/6SCSRwEr9ikiKXg0N3PijA2wFOh
48f/Fhk7srJRXkVewsisLMObWSmgwadZXMWQyvgbJa+DSxLMb8hKBynSqV6pwJwKnj+kjxekHDrc
bmBcnK6uLK/7sy6SATcgPamwvYGL/IsC5FxhKv4Nt2/AQhsfsMulVffjeOTcnX028Ty/VjqS91eO
LW1+BwlkMnTziuetElmj5XFGXyIfO57lNkOPX/ma/VNxzWlcbLoCD6xrPSMhpB0x27bLUyuOrYeX
zuUYXqf7S1bKC+Ytc2nOY2vj4axvNQ6LZZhDkhQEv1l8jmJFX7AQsrelEICd96NrVYlaMacvqtuM
kd8RIV12Gsyu0LIWK4SaDdc9SquDb1mz+lURfrr9h0v23+X8m/q66E2QUr+PvN+PMLqV74bph2Av
iYz/dY/6/r9rl2Xbl71rEqfvGaxywj/z60Kr0r0+ZeTAfyYWFEbECANcHstKGMOImEsgeSDiFzrh
Q0piETRyFuY6MJ8DmB/9BUanwTAdqp9j7lgGQf1AJvW9q7UIuCpfvQP2AJ5QGcgNBxeoYxV38MAR
CpeMQ46J2zPErTAjj6KIPukaAhZamsaCgXbmekLyzmr8/x7EfJS6I0+nVO75xJgbWt1PWzGs5Zy/
yPq+/8g0XG8UVb70XOk/vSCjbbMy5J/ZeU4QFkkTF6cbdU965ATBUdA9zMbcfCB2sngaRYHOTLzR
Q8g9BO32bpqEXWU2njjDtyfOQ9D8vGyNERPtk452EvvXK852aaV/1WRIvoZsa2/7lb1PwEq1nTkB
qH5/yxhgv+Z4Y03gxtPD+UNGZogGVMXo7r6MealRyqDvaPwv53C2CA/kYXsw3d7KH9eYLt3/xea9
pgi5So/e42aupVWmUv/eXt+HK9GW45GScqep7tukCBQNehV02m1W9pM+WUk/NQPPtWDjwG6+zn+z
3gk1ai5YR+/THTUmk5S+CXmMHQsJ+gCPXwDDWHjr1vrT1RcO3eue2DV9kSz2IS0WNyNR8V5sqqzJ
PGy1bm/8QgL9ZAKkvjAUqmU9KsNW9TTI8XAwuc+Y5g3lmTOq0OAlMQBN3FTks0C51tfw6AQKvA83
/pYsLb9y5yQFL+DRDkP54NRvew+5gPCaTQYPguEdWN0jnQb9f+wWZsvaF0ODKspIqlhwe5gBlTTz
x9FnBTqad7ZVJQ54gK6B9wFMjOow6n0iAWUkRfsqEuWmEROs4qx9maPRIoUpFjIeld/5AMlb7vxF
jOAGrsTcaMlJkkQkPzFz2QhhT7DjrjSmBVMypHALG/9jKdcRsuC+MYppXpb812GQNjNp5968tneu
ZH9m/fULE4vogwgRxbyWe317OyqkOyhBmhhsPgzzy/ihGB54jlw0UdQnQsKngch3hhCcm/kZWh1M
6luHg7L1Q4ivfIBLBkqYTQ8YGjrooWeHPLxT/AtJldNYudcJddWayWP//HIha2fLt5DLX0oHNuJc
H37q1/8HoqIVwfP1EVtPe0AbuAb/gPM9CuaXJfijWg4ij8e/C6+T8cw7jtWzqsikmBfUq6wIp3gm
4HsNnGXg+h+vbDhoWA3n5vkK2MclFOCWYgUU+fllkyi8XTTRbs2yZhA1xFvhdPoaXurDSTYhD4Ri
Y62dp2EhjYoQm4D3g9pbwDSjEwnNHGCIurw7fM/dOneTh+Hnl8e35pSR+gdD473UCYW7GrE4F19l
523gcDwiWvUXv4hR9fFwZXUryJzPiyiLLcjIq4p1rT+LwA2lr60Bns73EdmiBtPxylA8RS4Qjl83
4Sktyspj7na1C3k0dS9qynmUApgC/Sd/2HoRvDsihPPW82gfMGhgwcYPyGCvZ4T8IJYWVFOtJJ5D
dpSYERhyi+PRniJ9mE/XOy3IbEF1c2npKxwSQIeSCLaA7LNxOOGKBCL48aINriZv+P+ISlMC8JKq
0HM1BimRuGQdzJcnQ1yA31t8XaXxtRZ5tsrwi1ImvrIZdCeJX5jRpjRL/5EGuDqH+Sjpvo7jy7xw
rsJQS7QaRv4lD042UJA2Ch9I5sT0ppSjH/6P/YUB0q7w6zc2UdSDkUAg3Z4kgqYXq37hQnqLxSWa
PnY07iGxWUCaB3jWhVpL76fba1pY4sDBxDEdxtAVUtrjqGczKe8e3K/b+WC33aD4MkzJCHGhCEmq
1I6MCXEmCrcev45xMpthZy/XSYlAsPup6mGIqm9hs7m66/bqN3o4VLsyI2Q/2NQuFSpWJHURv0Yp
SwDqpbTpM3efSKrfwMYrzwlCab2PF12eaQacw3UKlu05oJ9NJG3AEsUuiqtL2nUVWn06HetTg4Lv
8/a0+PmCWzwu4boo7D0qoDcUZsemnwFLHYYBDDl8X+nt+XH9pH4JZJgiKO7ttkQ5cJadNCeoZcnY
egamzU2AxgSqriboEx7zKWblcJM01qbZty1h8a1M3zLN8PRZdQvPgreF3DEhfATTplJyPfxXX8n7
OD6kCq2xClGEi11AoWu1atk9lD1YIYzL0k4W7B5fKSro1WNgymIWee22tJ2hPwsmKzevPRXDscpn
CFg6KplwMeCD5MFRzVhN3cNhQ7uY2lBh8BBJ4CzIH3deVukjW+uBZGhvfTasdHcL6j5tjeOeoWe0
jsMdHPG4vHq9F26r1tW0pOadOFUzGhf5QeDIM6ecTj+cueU3muYDjrbrNdjSl2yB/PtlRYpBm04g
OuYiWjozLM0f7EHaWkhlHJZFiK7IeeY9T39U+Gp/av6QwuS9bN51jXhJv/bIaoB5EQrw8jotNBbS
C1a5XsPD2zApx5awf/k+BQ8YbsUpc0NTIvHFVM9jirzIXjfazWfutnGBA3s8vaPYQn0baoyRAepa
Zb2iRfgjrD4f+PET7vqTqthzT+TP/R8uoIPpnLyxTc8vPYh3QyPYSywnM0aWpNZOM/+SZv0KFJeT
iUpysN+Ri76sAtEGje+ypONXam8EN2wLwwJi5HfHygRzytRRLEN7Zk9LqvWYpEvD5+bL6Qwn9/rq
u1jItMZ1Mmp0XuKzBVg/KENcQYGtN2bQCINXsbGaz8PGg5PWxvfDf2RyJeDmWMdHIJls3QW6BnHv
TxSHVYFpuGuAGfBpoH+YOXGhbWYroYZ8ElhwiVb/+xMUe3zu1WRoFJGOZ3kbLcuw8FPjs+bKurVc
tOY1zJ7K2rqH8sbBe7YbdC1xej2qFrV3SoEftmN5P+xR8ALqrEKneEkwqU9hejzt4CU8LwF8BKSg
MKVkMupuEkJ2ZynbeTpQRLMG+69gzi/h4TwOFRpoRd5pkyyW9Nshej+O4cUZjqIpa3XqMAJLYTSy
LCXPnXAavXRcvDc8X4maaW8BKbTl2SFWiU1zVhdPemvGky97XTFtzxYjV32PIrPwexYwZnoMeiSg
NLAvXwriGIdQG9/nRNvU1n2RhLNfH3RJNlgFk4uzfGqxaZYh/jWFnEKHCzJchjtWmckE2n5k5IUD
UB8hyNdTwdOhIKr2pZ7gVl+o6j+HIrcBJv/IbY+JA5A+y/0mgs3X3ljJDazX9z6dZI8ZCvkkSUIA
dl6bLbrSSCimGPlfCyUBClFbv9H2fVRh+dx4nQ9OdgoyT3h1jOihuhzkB5CCv/Bp6x8KwcshCZU5
8JV6Vt7+35HbSvl2jR38DKr8Hu4xz34tL3KpEoR668/IVfkssWkh2raEQX5capMkoOcRKlrVOCiQ
tOQlUXd/pSCzQogoJq0SM2Rac+I2dlgmn/OADhaqoeIce/srTiAPkIOyRHXZL32qJ6R/PAPaEBp5
UYrOnMuF2gnwY5A/rhRUERgfZX9xxyCZBnpBRIiWtMCXNie0/FR18BQauQYSNGsi6sPvZjIIF7pB
Z7O25xfw2BZj37OsK3au3C6iffVyfmry6kNvm8CgVjlR/IOz/0MSSEy4ph36cJkCJJQ6/tL6Bldn
VvB08MjN7bAfMxObkVTQ375s9pkPu/sHamNbMo3Wa/hhJ4lrE0h6Abj/rtY6Yg8FfZO/E7FhBJA/
SwPe92wEJhQmbCVoyRM4S8kYAsBS2vGGppjuoBoNPUj9btD+y8Z6/d3u+6MMx7aypEr7YIVVOVeT
8rZGB7eXV5Vwpk596HjIHVLHgknC8QTL+Lf5Z6KsQRhaNJM6z7jaEbaNAd9WK1R7QPu/1SwCvGYr
+pO7fPdMCc8GJQsKQNDfoxv5eaocF4BiLud0/buOjV6RB3yM5yUKz06808hUn9Iuyk759yvAAwDl
CWj5yTLweQGUIRa17NAkBmatzM7R8M2I6hh6oY6LWYYC7yfwqDWFcy6bbn34uF++0xqcFfvHXIQJ
cUF0h3SDjZi/iRUukAXia0tY8EkEXry7G2d5dWg9ufOCMA4qIeVCs/UEdW9S0h95bbmk/zhwTvh8
WcdyGUDNbsTEMg01BYBI+4mm4Y5K7r45fEzcXGiwUHCU4MX9Neb5r4WSxi3OmUvNe13MTvKGVDFu
yWtP+gGexNd4ohRWswQKsJCosAbjaNg/9ahhTLcME8Y+NnOLYmpu/UkS1BEIQnY9DnB3h+EHAGkz
HtZqqdZr/iL6E531eiUCOWDKz8NZdWjIe3HShdaP7vPo5R0PHkmHQVzXkJlUorXjTrkIIm5CDxVr
WCp/X5cXfJDao9q+DxJU03qgE69eUnqPNI+YaX14wxikqb5Ahnm/SFdAJ83EUApaP5MlneCbhbRP
dtLFHNGsu4COAnpddtzOkOsk1XGFMI+tqNCb+Kq3kkAG7qEoPGaF1elL9W5r9+Uavbf5QrOJOKPZ
YQsoJQKUvDPxjsVUmzCT0JRmJwZRzyZELc+NCi7F/LBxZ58VsENt5g1wRzmPwI8aDTIef1JR9RQH
Kj0r5ioCT+oZigPSXEvMafweP+5vPtF7heKcH2KmCZQbX/z9Xx2vG5ywbNAg3RNzfZ+61ANChDFJ
fgY1xRHtmshm+wRsLAKavyA2By+600UQGzL9PjnGQ5LrFqfR1AdWrzSmGVeoCwJYBmzAK7/aUMmy
UziQKgHB1q6ptQSkqSwIel5FTYizVrO1rvT0ItcAt4FTXk6ZCpgJw3ude+8iFB/00fN5Gb/PBmXl
EWCdfCGPi41CBaTNopMYPeVnxWKwhrO7eE7jf6rFcxw9TmCSDEAXkcLF/6Oh8vvQ69NWj7TpsrN/
ZY/oTEgODwxH1xPSiNNJHYGpp+49Gv/ldBY4WpuLdqrAz4SpEAHvsOn2ci7Iy1h4Fu0Uo978+WYr
thTicbaZRk/3dSlVrl1N+q3QuguNB1c0dQ83X9fi4NWAlNXHiIq7Xv5beRk5NV08yipt3Ai1F67C
8qNoX8eEuiuxoVJZBUWu8U+rwP2u/8hf8vK/w7inXG1MPnaD0yfK7wnTRWeiI8QZGDuUEQResBc0
osgeh2ygTrDR+kcbSXXvQaSPKHJYDOHGpgwZaVrDXW2P6t2OE1soi/Xt5ipTB3L+IzB5HWa2dTsx
1H31iLVOAnMVBMIPuIPJFE+UX/B7/xcUtTKtq4EpVvnusNUt4NqfM2x5IHP7oVIWsf8DiWBmYgDC
NMuI5+pwlu+hKXWpL450OMe67lt2YdZZCppCuhx2Jq61eSvaNJ+ccBIoKRfAQ4sYveFQpiVshInr
Ol1GHA72xKrIg423G/4vjBl5QCsPYlipwVdBkvuFBK4ZoREubxfJfK8w9Jhz4MBYtnN+sCoze9Gn
kBt/1ucfECRXRs0mZUBVKDSgTIl2u3kpSh+kQ0NDN2aPDB9GE7fyrGjKLmMmzJe4hwikLL2+SRUi
etdYcaqtVe5mIpXtffXUDPkDI0uAVW+KpdqwOoyuSOVMpyzHAHqs7W6ZOJFCX4dsBJ5CqetEcCi4
vpMEJPJZvlDjp5CTL8w6vqrY+XgMN3F/w0CdTgwP/DhdJxWj1fEJMuVoecKtMoX6zg7RgYuoPTl7
OOhu86dt/kBGPUp7zkesuxU2X0cbazI78gRzE+Zg2+1bjuRMUSRWNSXM2QkZbKlqDil7aIjvhVMa
NmHsK9ybdy9bV2zaj3ReXOlZE8k3IWYDf9vIt1M+J2HD//FoapSFZkQk8OGRTA7ehrSpBYpiWXje
iFmwkI0KPJ/35Yz0EqMWzipNkhbwHNlxO2DuA48d9lbA9Cg2EQprfemYOAFmeC2vUrguPL/u2mS4
0moeTuUz9yT+UdjXYEBCwKr3jCrLQyOB9bcXL/jv0wGNalRKvDPHok9zs52U1sx+PJOONPwBt6ED
Se6yppqYu7BBaig02QGsUa0A7gpAcH5gzW9rWUxkST9PfwN9YdIFMfC6Ekp2KjLg/yYFfXR/euJ+
F4WM0EwfvLXrP1IRo38sX9/eANo0MoMI1e+785dBOjnCfu8eAptXy5Z09qSe7DDJmQfEUHIP7ah7
bRhKzPr2d53gUq0N5PvhbEA6edq6xrvQMmm5Zw4iuBsXbC5TpeyIxRZ8pJSjgbFP0xIMroYXsZp6
OnmAcmEPlx0KaQjUilQVHvqwoAUdZd7TpDSL2aDcCQm8ua3FYGhnUsH6LVh3feh8zAl60S8L1B5O
ckUriEJCvjlEUrfrotcr+IOsjuQJqg49TEkcILU7V+BVC7/U6revXUx4o6m6BXw9g89YkWFT23VI
XN6n5kTSnLCnl6/8Ng5OgdMeoJcxgovOKwksH+VVwH0kakz9yq3CbqN/9CibCUG2lWkVDejBY0EJ
haXQp5oYWnI3kGjGQxikB5du2Z5s7hdjTveHrd04PLDp690oEDBDIHyXcyK1lfPaPbrdsSBTQZFL
vZ85NmFGfAAvhoB2zBHU4d+opBNaaiipd136nO8k/EwQIyt7DgM0qkXycl/SKWchu+nJL6GuwKiZ
lljhnDylOj0MBOoyHJUUOjiTtP3avHC6QR2V/KB430VrMWs3JOmMhYIPKaZKNEzev9+pmGdL9pS/
9aOGtp5pAM/mWeTY9uTJ5mcJbtcMkI9XQqardHv4x0JRSL+/9Xz/pUFVL3xcR+jsspNXS/lYguV3
9ydHEULEWRGmetwFTfl+lt3y7V7bHac/2kCfnIQPn+njduTR01SPNkzA2jn4r8YZlBMZtapXDo9X
7MCGUUnf2Q43SG37HQOwzRE36YXo2zCkpC7gA3TAEP/PU57AUuYUkC91zH6JKcKAfstd1kxzeW0s
vHFtwKVvPDnv4ICiRMU+80W75T14EXbUAeLNC/3Vk2VzUL6srp8l54nzHC9DEbjGq9czOzKkp2Dr
yE1B90Cbl12vSHWap67dwarzIpM7YH1oHVxFp4twOGVEQQU1XZYeW/uTOuQ/28M4woV+XvIxFc7E
SRr4NrILEo/6I6fAf5a0sCrRqcDm1PtRGMih/Fwl6JbQ+BgaHpVW+818M3//686kUtMK39f3wk9v
5CR/dKRF1iZHnELsHxcRkYXzaDkKtZ112XzPHiMPjDXziavHcRWOvUun3ad27Z7DaujHJ4noNbYm
mxJ9LBmBt4IRk+5p18LgkbmqCH+xA+EnPmukXetKV9YK5sdoJ9E9+XcvtGuaX+vklIMy3Zehnog5
w18RkAXsieAxKmRvBaGm5O5muIC5ZZaZUgL77YZw9vHHhw1gb4aVbqq5RsU+jQ6CzzWwWm39GgmC
os3xTUBsBf29ySjNSI7BmO1jS+Hrs1Law23wEwafxmi3dtkk2BGk8SI/jN1IJPO0GOf4dwkSyYCH
rPkaR3+hRPPdEWrAqjy0F9USq/x1RdR8cWNXVviTYtPY5s8gjLHj7gWUC5X16vOuIBkTxWlfHRJm
C60USCs2W6C2ibXAqtKtFbR92MarKHdGlFEpnbVw6pZFeF5hx/bEdOza5/JRN6pT1bXeR5jUO9Fq
wnXLpKrFJH4IOuo8DTSOxge+z2EMjHCt3D3xljTu20mtD7gk4ds3bBm6h9Utwp5tPxtvAsF5TIpo
Hx/S4G9vi3hxHXWttwF7xfRgDSffrpSyP46iu4r/YPwCYWBUKKriWgwxUESc0ivlNboehezDEOdR
xgZhkOR8FZxQyJH3Rlp4qbH0KVHs3Y4EKLnYEUUpA7z3w6jV8qtMmJG1AcGXwYOGno6n00oJmbdw
hAK7HLatlIOEFCUuUDt6lXrukSQsAHDR3t/unKR6TufLg5YyL4wV7zsxwNj4tQv92kfdPD66Gwja
7eiGsMgDgEFhGWCTI/ye865Vo/G9lw/3ekU1Wi5hOKIhJnYxNmazIs7Sz5RwYJXjZKLOYCgxkvav
Sxfyj9JSkTFlVhqE7kdmBdcollbXxYzh+V8ikBCBjYzma/NUmzEBO7nJ0tPXsnhjHlWer/msC5cG
l9bgt8PAjiQ4Nrf/Fx6r6OWjBegHwuMHaheKy0ewEYL3ZetwSOGLgnM0dMZH+dnjgmpppSBKyTbC
K3KSzAIO3mB0NxIR6py2K0QlHB0Rhlr4OWD42V0ekpSI9ek5MzOSSuRAW6OkMcm/HHtAX0Jg+uci
c9F/f+lNdZ4oDJtJyT/QwaRgp0LDFXrefGEKNdvxvAq4eFXTcgTcAYOSe6+gKQCtgSambvjsXnzJ
6D5MCni7TyhpsnIXGGK4GmLY5qR+3FXucL22UN//YMVwR6bv1PyTtB6FO9AnWYERKOoMKihXaHah
h9veg8FKh56PVRruC7l5R8FWKXBNtpGqf4fXbdVhqdqI4rjKseHB1E7TIlo0vCiCb5IP2/rrncsT
B63NsJhoZEliCNedVGlWDwgyfdWBCOEDSyVKqInlcs3TBTCxewLtgJr27i6Y3Bs0JwnU4x3kYnSY
LE3keIRriMeIwncuhA0kbxqf2woCgwswj85wUUNuDhhcLi0a9gQBFe6V6f+xxzsMyzEQOul7GrEJ
FcMS6O1+gFGZmilwlqcSHJUQ34cNzeR+8w4SPJMOtVNe/c7PG6ouEPZyTXJve4s5AhKkS+H1Wrox
pqpR4nDadaoBInDX4iyXahKhUG9o6LLHubGrV27irGCG1EPsIYzb0/1AUa3ASVS6lSQIGJsp95MZ
u1quUdBn6YXhgvVkpJbzOSy0bewELYL7GQxkEC0kMQ2S0RVqOz7apEMR6N+IsLhCov3/d842HM0f
1bXnqDUxvmPTrFPolw/AQhR9BPtll6u+/3txwpGIE0+Iy6rhK/iToae96fni59SJPchxAXzuxhql
CyN1+vfBbx3iJDd6ycpXko/6VD4xjA4mMqmiKrv5+S4lzzPtICFp6uU5uG1A3ldA23Ho55JzHHjo
+4C3yf1S5UkRvijrubem1fx7FahTgHDu+psBEKHGsQNZ5b9LN8YgY/DgUdU5ESCVcPiDmBC0ZdiD
Qy1/InAhiZIoXnUauS5UVMRordQOZ5Yodz87xbPb3zBFO1CumtVLp+5NH+2iYJujFvJWXgCRSpX7
b2uU6ct4Chc/kgj6gBxZM1aP7nskdnuvosVJmwv+qHAUQkS+CiDq6yUU2PsydQq83iQP1Uewi/vC
dSM3uXF26AQMwyBybN/qqTMEzJW5VvlrwoczWCjngbuK9U7B56ExEe8zs+aR362FzSvBOvZKlQIX
JWo6XpaYA+7F/Pev2SgRPTGt/DlsVngpj8m5/yOFXBRotBOlcch/ULCMfdXcsTDKktpVcikzyTh8
Y+BCjdnZMmTJrVDv4wfBXg3g0jMuxs5u9kGPxBX886mE3OGdLVOkCOsw6bkXB6rONuAMi+qhhn8r
xNbYaFyIPjIzbDiups7/KLyX1iblyL91Kzbvv0kzA5g7jDktLZSeOyG2a+QQjgKNjnGfnVPYQz6B
Cio2TRiLDp1aIHN5AyP10PM6W4ZujpGIhWe4UYt1wXlB92s32GMsrPh3xYTjMXY0zuwz3hbpT51A
tb5cDS5J92U5A73M3k7HALZeMGvTO+cHkZkPp2JCAfk9guUDPm18vc0iQ40hvTaJIg6GTMb1kIId
DH6MIjiMaXh41kYf29hWViNyfDvoBlN0atYpDSYKdz8VEONGxqjltJo3I2qwwDMZ9XSqPguRmJOT
6jD5XJ2QZ34Cbe2Kk4HdlfG1qsgKfkalsC54840Oa75SHhQHUPGKubQhI1XWZpWLOWO9cpuGmI+w
1pyybqRdSkttYqygaJoyATEjBGrTmnJXk5MMrsr4qsdB0lnkjad861TlkHe4s8tEmmEFv2ciNwh3
hPBs0eJqSyrCmXsBW2bGwgsLtzU8yWaLYJTPISQi2CvbumCTGwZHQBy3BQ3EiFbARNIoHId28JCp
67AHegwIDVYXeDM1So/7LIFegsB1/a17/6rr92cBXgKOBQe/lTHZFuiKHl7o1txChSCK3mm+Fn81
k81TqfOHbuYsFJCDc2kt+OLDNnlSRvbBXRBymygX7FxufZnyy3b+alFdhuzHG174rYncfEoOplqs
plfIPktXkDVUP3WGBAxdRRgX0TJ3NSLM3+IGe3L3ciRyQlnnwgU5RHnFIt+et2U8w2McnpRsvIHJ
ZorCOoJ32A4KkcX6gzN3MkFOcGUyUkTb9QTB7OvZyBLsw7Duq7QdiiGwZ/l8fZakWnHSj3BOuaiN
AvJd1mBGn838wD7J0+qrBgvsX0CvHJjL0C+3LWDLlj9MjP/1hxISzvA30RfnsfqXDZPaHa10D88K
+Onj/U1eDyBj7ZzKnnH0wb1PN1s+m6DS6WN/Y1o5QogEWh0aNDJwEryDi7U5aCFEve0/gcTMrmNl
5xNMP9n1AhPdk+PmPonvEfMUeLhanKMZJsUwMBmKinF823+bKgqEroDpS+4+i1Ubox7SBbhIFPXd
466oCdIw3Whfn+e3QQ1ov1bnTAZ3agopXe9I4RE3DMj1ZHHtFpEpXcWY+Uxhs5FkW03lk1lVwaD7
hr5ytAuGUJjkP+auIRhN5IexBPFoWbdLGABtuBhMTrpRUHxPUfYQOCtbAXmRmaHFKMdIlSMQj/Fv
x5xoa0vRt93ZVWH8zsFcRQ5e+DXph5s5pKoORvwEgm6mCBsTfSO2xT1rP6r9HgaPkOjEwQkEO+ik
burZa6QYWnFczPOaOf69NvQWPUzGZYoMBj3XrxdnAjo/SC0oNRWE5vycFp1tudTcbfoDVyMy1e5w
1+xjLFRUvy4nlmyNuVXYD9Axdpvpv9VPg20TIjiFwOLSawapW1KxpcLH7F0mZa/RGowomTtdSaTH
Qs1KfKIeYCxcV474afxsn5qN0WQ7wWz3MuLErN2loEMLRS+fXy4Dnl4zKaV2F0WKGLhCoBfX41FJ
ZkGtqsJ/8sfV+9fe7HS/Hje0A4eapAHYkOkqHG28lBUy/WWBR+PBMPDQVXG5QswKLcCjSzScd4bg
Dkj9YwpKouQC5Q28rAbq7QuTWbxNWh9xA+CoKau6XmePqdl62FZaLVMhZRCsOoJwo9TRxHyf821G
ASkcmmZaF9qXvg4U0kP7/yQEYqbpH/WwgIxYodz0F4wVyf8RvPVov6HvHk4bLYoYPBPPntc4LXpy
iQeWK0+aKQiVhnCYvrfa78nrZW+hjqtA9jYX+mbrRqZEPRIDSosSZEWKVxvFNI33BZYLJA4eyXS1
jvGTr7HwZlsxREe3fG39OZJMnILUQLKu80977CxjUANx2VLRBPYhIOwOBYHVQA9GrBLDV5QOthHd
LB2ciJQyOjJDkF97SRAuaIJeqiw7/s2XmttETlEPsksFD3SQLNPSKfyGIuyrHJEUH+o2Ryh6el2S
JYr6h8o2q2FobxA5o9BQc4vF8S5G/HzN/gWcLyQ0jNArcT5Myti6lVZIAob5+wy3K5p3TpU/1Mv6
4mkc5tKfo0vssBJwd0d5iTAkf/pga0E82p3gLYPOI4QasZ37e9EMWG6B/xV8Q784E4XwH/x0Xpcb
5cqrTqHnCpXgfdQsXyLif9SyNR4ohHOloDFWcGbLj5y6+V8hEu/m8K42MH//PCCjE6d0HjsMEM/F
RT3U6BEZndkdU78sKwDCwDsmvqC25uowwvkNyei6J+rkNhNMLDMq8OtiplvFv6wc7GKI9VNdLHEA
XGvE67XaQErqvcuxaYckLVBpSCiCa/xRk94GsChsev5ekaaMkjVx6SwXmuRMxQKA0vd9g+vKpFqV
owGT5vqZtXy5he6SpK8YZ8O3JAOryJ00sixrEP5fTYDQ5H2xxIBxg+TalVyXKmVSCTDUTfUIFJI4
8/oJxXruyy4rPuejBNSiDP5KgTS3V7/B3xz/359qOyBn+6+GMi+GjvNA2zCyZYlyvrc4+TG59M9Y
djii0dVO906A0BmeXr49QFKmjB/hz4d7W4RRK5dmDfu2SwrFaXp9scL2pEn930vq34Q3b5NLgvtZ
cNEEJj/uCfSLcjbFa5YaJ4kubyhdPn4UZDL2ODqhbemUCBfOAQ4yXN8lI0BMna/yOi71lpAziQ8E
BNxaLicF8JuRum4oxeCiVjAUrIbrgtWa7a+5O9PTliVRn2SbjJKS5VaqAfJLiTUmmHKNe80qA98m
mEwHBDVUhPeOymdWf0Ry6HVYvbSWsWC/ANANFbrOBuLISAgkEDg8sTgu3ZcmDIEXvpfbo44u5lpB
8afTs9KtB8zwkALzw+nq1HdOpEyCJc9+umx7SZGyyfYImxPAXkJWCNlVJEStFyWTObl2fxfhcrIk
4T9TLdI9gvMfid0mqIJ6xRxnsRkw50fzgpp+M1vv3FRjYBmEDdDhBeSo8+QJyCVGvG6+DnApiDbZ
A8QK7uFZ9urb0SLJmVAiMAwDb8F7hhYUydPx0LIYi3EYtdOFrY4tsHkpRdSQvXI1gNLBD+QXjoF3
o2zpJ/Hzx2J3fvC+DkvZs+Wd1u9Z7+aaxu2sPL2vX70uWc1EEkXdHsJQI4JSfPal8P2cQwRA/Wbk
lq0vq0mdQtMAgvdpLkL7J1NdYlpOKPMPC+Be7KnqV2NtpnGK0sOEBkwTdu0FlOVpCWKqI7Q553RU
qFOvB1c8Lh9GdvuRRI8PsxoIBGG+YwR8qvKFz/TSNVME10bmI7XbYYKVlejSMmwqJxkrd9nKdZQp
wd/Wi+x/M026mEQJlGEDHjojQIzXSGyD/0md89FyduanPE5jFuUDyOmc9Ue/guL1nYi3IlzSV0ng
7xTwNhQ23o1tZONKtE9jlvbWW00O4SKV+MHNWOY2Dbm20gbxxXgnRaIEHSrFIaz6ZcEaBIzXWIMD
QPXmpXBYu+RWX4KM0VAgsnrk69W5cPIpbzu/Ir+KO5DLPa6y+OgtsDOnTQh9m1wRZJ5mSikb5dSg
1I620F2w9p58eTdbfU8CtmFbVlQlT2TY5Tuh5x1ErDF8JIXWtf+S21SG7vMZS99TSzp/BBcnFEIc
lcGBQvYGFGYPDN23sjUXPXSzBIIBDIq6Kvhe4hUJMjjNo0EsQ7sfVXPs6mlFFakcSfXmWSyWZoUn
k662IwrMIl8yngUIJH7zvjtwfBJOG7V3Amo8JPTUW3TJjxzcSXYFk2X0iCyojlaF2GWZkIHkhNds
zE29af0Naccnf0wOPnACi281gWAQfmR0tda6dSwSrMjnXWpW1xq+mXtaPGo7YqOnKWAdUAyN87yb
qn9AZbaXmDEEh2cOJ8kYeN+CJgaSX1BVCmykc1YQsuHZDhiSiLIaiZtK65PZEP9vm42I5D9s/M1x
5rsPCh2sgDfxoWrmA3iW/aJ44vGRvSaeo9//xCzNKuwIFCvx3Rqr3waKcrsBhnDnQTtJvgoQfNjZ
AzXnAYMxUnKJiitLiqInfyb4tH0Io4viR6rqTP2iUNlToNwpj2DgxMP+94WvnEudRw3AS6xNtUrV
Z3IcNjMIV5OFHQI6etp1CrYUovlJn905yCJMsg0e5aszfrma6YTL908/5tSwtl+02W6pqBqzP80f
3O0MQkf+x8cJ261EeByEEe+lE4DSMXEpYf/bJMi7dDGQ8leDgSpsrkgKlhIjfU6BsjaZxatEfy4n
Nlt2LVDcqnA+pZxWY01HwoHINYyUFdEV4dTR+cCrYKevOQFVNDUpHxjZ2VxxeTk399N1f4fr4IYs
Ryzkq8f9oau7Uo8iWQlj4mRimUX9WKiWDMLr9PCFNNKBwP0d/olZqz74vqrLGpR0+gIGMkFkaea4
vuoHO6GOksTUVDUGC10r332n+NwkbxymdtqZNiZ7SuHU/MbmcaquCqdinWQBEkUacZbVZByW8msD
RBRBtT9J6Ga/MMtUbTmnHJrKK6G9OJBg4CX5Qhs3OsbR3nDABq7yJCbBnaQ5SuQdPDW1S0mBA3uN
xudv2iXOr+rr94y6MgICiTbhkxFp5IB1rnIcKPDraCRhoF3aSUEzmfFqOSDAQWnZRL0EfjkdUOn8
wIcC15rOoQE7vGTs18MfAqBF7MGfJG5otK/3uXzVo9Y9YN/ABU6a8rWttJyXmyLfF3HFJdBSD7vz
mtz4BlNx9XWM4One0hUEWLJkzirQp6K2u8T21Li1cd4XJkSPCcSmi6Vf15q2ABJBoFZ/9+iBcF00
l25QXtoqb6jJU8TNiwLSr7qbRNkYvpimjhhbDivwydtZN88qn9BZ0bqEFb5xK1Jb4sI6JoZbDjv1
NMa2fh5tIytNQ/RotPPkdwS9HLQ4zESGDjFpLVdhAt23qsqiV3htT74uOPv4G35AiLFwrhCE9T7f
xRiFypDJw7k4xS65ssXSNbIY7nwbmm1lSXIKO6qiS0mAeApSGe+VU4MTWCxEM2Hik21L7L4gpCz6
uhYJgNTgE2Wi1KxhW64Vk9T3wdvyewHqbn/hlitTh4+IoBO3zTivrIzi8pSII9GweSHGnJ4KpoCP
xOBz3i8HDZdeDyNIaDvQ3uvw7+AlvglpodSObW7Z8Lr+iDZ4Enh+gPN7vkqHfvg9VFFyoCnLCH1U
x/ImyUBbJOArZDP65bu/QeyU0gP+keUmtHg3Xexj9nx00MTMgojeV9paPYE2DQDK6icnrsTgV7pH
a3JhGv8igM/lbVdPJyj7qILGS8/QUYrqfQTiPK3dbQAd+uiVeS8Rq77lKfJKg9vBwj68etz7XWBc
uikGSuDqyc1cxASKCtooxuLiPJfGU7atPCTQLZjVGhvRXw8HsBLUC17FguuM0cAynMwK3gucAjjm
RozlgL3o+/mldzzcalPNp4NLlt2LWsnROAnKIEMf99kGzpUbNiO2hypKSBYeqvjHkK6LE05Wm0kQ
sspZMvZIC2U8Y/dDLP05v8CFdy9GLlsaWQSxNDBSFUTo5kCHHqkeyop0gjKhHq12XAqBa4AyGp2P
8pjCHlFu8WNlnfZnqrXQ+PvJVrHX9odOmCB8+KPQQBBqW0TzmTerQFat1p/a9f34INMAgA5weayV
UtkjzF2ZvXhCW2ftAFjAQaeNSPTe4+HC2VlH/lQtrm4tAEMI7eeyoJjNLE15B63P9YIvIrhAHgfy
LJYW51CjJgDtVicr2ze/xiz8HafLYlU+hhna9yT/kBA434WkB2IbbkJRVsnjZdwnxsgcktLtekHm
omI324CynRQmn2W6DNEoPoJyAYnYeagaoEpI4VYY8ljQZLo3hQTFEqb5OyJGRcqMlx29Zin+SHLl
Nlwj3Q/e5dcYdfvBdEZsXC5tip10kDLLDRVTX/AyhbvBHwDYPI+4HFrzszAI0i3fqN2+kseAKIYo
sH06vUmkrrVGNddUHcEQxkhWIf+ryUpANh2BS3fNGNzvbY73ccDX4C/PDJ4AUoZK2HTkj5vA2EeX
YXXeafjtO8fz82+uPPF8Pm1P5UHc4jWsvwNrwGe0paUCqUSmmS2pEhT8ombv+aqQtvXGXrf1fPUJ
8ErmTrjbkHVI34RJiPv7LnEZsXw9WrVu9BPKjK/uiDCr8Z6wkpIYM/D0zB4tNR9qtvlOefWXdIgX
GQx2LCe4bmg9ZYj4uJFWLtS8YDCsyKqXYcIRdG0nqvWACaIR9h/v/KFka5mT6ZacWsnn3Mmwg8/U
qRE9zN2Un9MSbH3sFlZm4FYoS+VlVtpDTIPHk3KIlDrCkaLFKpevQfqTiEVQ7N/6sxQY/uWS1dh8
23q8bgx1iTaEiOKkLpAvbtpILRlVCVrQwnMD4fZTz3Jx8r3Q40NTm/SfFw24TBHv30YDPw0E5BKh
wmMmHnj8jJ6vTv4hjymJ1KqBcnmJ5lndjbaq3BjAQGq/pToeIZSrEIhCRIyH3ZJNrmyezBa3j+yl
68z+cCNLmuyQyGSTC/rcUfS+S/f+fWnQo8U99rsL2FnmztstqjJv8+qr3Tn/3co7E9a2LX/N1fpg
fS3WKd3//VPOcQiFR5Yi6BQOScpidJptxDC2JKz941g16s8rAVC0kDj3gYaJjf7ydrJPwv6evKAG
MRDTc4BU4ogZpYCV3TEck4W2STYOH3PxTpsJLTs0ZTfvGstmJP67zGP7UPMvK8Q5V5n96ydie2te
QZwF2uLrfiGAAU0xDBsGLT4nxDjE96pVnq3kppCDl8Op7HUacHI6yk9y+h2HH2ReSv/QA5k3L58/
lUP6BDq0Rqw+bAykqCfImIHvTfKelA3xjt8nxw08pdI2l6km3igydwSfLf3W7YVcKJC39p32m9Da
ef9JgQgGK46T1c64uMEHnJKdoJxOsczvBGKpxX771PgowFrKinSVLgnZ7dlkEBnYdj0U0c+cFGlg
sGKqY6Hfawpm3BB8dtCAtISTFHdQzqQLueSoDdsOUi4h9LQYEnjdUvQ59lZ8WVYKdxQcps26Npcz
Vq+rsAoCZZ516GxnjENSBAigdFl2EbPrQdXFcuTEYg+jLIy8k8X6CP6PhzEXgutGJ59JLrLKYLdv
X4plf/xND7U3qTfIAObOzM7thDN4IadGDShV2Cd5KLrLBsCI2lJBXwgyLGYm8cfyb2ucLekOqitf
bX7TmMWQn+juuatUuLZYjiDQfQ/uEhmZg3ZkSZhK/IkZCRk2RHtI+j3/MKMCpKUsXz+5seNV9NkL
M3aaEpxFLOL+tY4Y+5Y/AerOciXkREpfRsC0oNXydm60bYJryUkERT5trV3JEgrSWmQRK6SxSWeU
WvrYOHMidglb7gDfZKE1aut41CKdBfaivKbtW9b0Ram8nZQzcISNt1iSTzHAiFBC8P9EycRrCeCW
K2GDOchhwLFtcXlUTwhepy53TQw9mKlYtN8Bz9YDLEE0lIj0GUmjdR4Jb1X62hMBClLnKPBiIETq
FgU2a7z3rw/WCyKHIenXEAnqc8/sEJzIiW4sgpxhszP/bBL41HLd4lMmy/8NrraMmFLRR+WugPVc
hxGSzB0r8uIq3UdaqxCUWb9LHpsQis7fP94pDbBPze37dtVxSK5RH4ga8Hl9Ht0yyssKbWWoSc0Z
n6Ieq2Vc2ExXZixav+75JzsW6suax8ZKCyyBFzEo2KglN7x2gf89s7tVUKrv9OjJxzb21aZxQBw/
PAfA2y5qvn5/cYB6gn2KVKKJwNMPbVFySRFA9bMzeku4BwCY8eB5ojKTrvTFUwPr+SXIEl/yFmVU
k1ZaoLe2Ngc5snj2KZTIG5UEZo0KpGXDx2Fp9yoGPosqpri7blrRcUkcNr/LRgXwoHhj4FilpmrO
9tTISXEIj8BhMIJpopADOz9V49iCE7l1l26z463MEQQOlWthSBNh3vKxXpRE7h8skFWNDP19qoz/
CkP77b1EX7MBBq4Q9CHiR/cpe/5uA5hUuqh/fFXL6ZOS7Uwn8lQEwkc3hcoCrBUMfEZ9qRQkZVui
k8myZUiA8NZDaWDLEJ6Mcr2Ph+HtyGtzoCxjNSY2FTKjy/NJqm2LUKkgbYB/JQbR0Azz8cjJrnCR
S2njuxgMjSEAdHal7Dc3lrPAa+dV88afN8uLe8xA1tQ5nrqSmn46iVabQuUFTGHii0wYSuxPjHct
wXXEc6vLWFYK4U4LJeQqd40+Nz9HtimLrhuwxtGgoI4beamcikzflvfdzNDNdi44u5ubYABFrDkc
FEHPejcK2G661fMcgVuNrO+W5NfzLCSbV8AR3NNNhrxfnHuLaMZE1W4tSEgLKaprSmNTeGc9sDvQ
SnB9PtJM0J020E/s905PdF2I5gghA+6hx0t2XBbcTePHJMQ5SJJfIQ00vPgV4fad89nr1gncBGqe
C7mlZgNBb4GkQEugq2YmVSpm1knflmRuWofmN6AKy94rVBrht83pf6yDS1q6SkUTvnXwQc/LEJXa
R50OBBsCm4vdP2NaDT/1V2eNGhqtKVsVvPkIYUBFp2smH9uPit9kUq+4tee7fLa6shq+uKu/bO4j
QDp44oOusXLzyLbkx3L9TthaUhbXKEOBpUKVghdnKf2xG8KAFf8vuo1qcxhpcveo6FCSWQNhQ/JF
gv1b2zdTRaCIewejfLYEcGMiTo5v+2VT+5o5Vo15Fu0g6wTSv7fLWABDgYBtRNREtiVcp1sC3ZxY
T9wrLOMpLdoSNPdaJRpOr3O0fHqQE5UB+56PDvzweASvkCksZMNhSzboCXQi0g9doWLpv8Drj+e0
JHyHTyeuWOZjdF9IpsM2Kbs+f6ZLu3ujZ/uRC0iOtT0g01PfpQDpdSyRyVIymIS4U2IqDythgnwV
FMdOF+ydVV+oOkrPc+1za4DPcz8K3CiF7xxT57KamUg6PsacIclwj4j/dNT7AYemA2FHx+w425bj
6sTFF2VFpWVczSqKVTwHr/dJLn3IJoc3ykDxRe570rEnIsC3nN1rGgLFY3mRiH9ZHZkb8BEnUHZr
qYg0C2LTZLvQZhgtRGYS5JloI9LHuxxPOkJIQSqMZ9f8v8CDWRB0FBcy/Wj1Zr9V9Wrn6BQ3OXrV
H4LHPXh1FO9LcEDEvQkCQwTAV3gRHIJRFn7Z+ruHaXVuMOc5aiQV+glmY17QQYlNhqhlj3oPY0Zp
ZoXsaXlxb2cAhF4g7J6rpcDxqdbMNS+ev8jbUMfA712//dAE/limMf6dDGfd/+KMDjvu07Xvd7H6
83fengNFDBzQLCMt2Guzc0OlZPtE0xnppu9mTp9Kcj9npiD+AaJhGjN0hHFbM/mRGAvR5OoAWcBz
t8MiO/KY8NpwMRAK8Pg6gyMJYvLLb+ZGDC6G/2kX1tOSwof8sL4Gk125ltgWVeXLIePJO79/iXuv
K3fQFYii5jkAVx1Zyi3FWWY0otsY/Ru6dRjf1PzfhtCNJO1FnzEr4db1tB1kUZT5hEPftz5ZNzZ8
jN4JxB2Pe+rCxAPyEOR/iZHBpwwdiIDxSkzludlMTaePjgWFeCjxgvWkTiRnP6d3CBP6+/ElLBM6
83inw9+GquKzaOThvkofHupvDGynzdNnDDfac70uhu64J8Zm6EljmLcKjhCP/cJLIkBykNNmSrbo
q9Uk3h0H+Ruog5kheDQvSmp0DuvfyLP5L/0M2fkAKlfm6y7HZK31P/cbsGmyFlxWJnxIlvInKLto
izam987L/mfJms8HN2f2Z1dnT3FZn60JUY/lXZoQwgNPRUZjGMlMFqMhUb/RQLdVRPG19epPehLn
dLcajkONF8MzElzbp2l/KQoj4emrW+1PFiO4vTYmU5SoqEFVFafBt0giDnu7SDaEwB3LkTJR/7E0
DXgTA9zyGhMWfVhgYmtBGXeBo3khC4yjAWeNvFXJIIZchCJ8Z+8TxVrVMURwiDflhzAzIu9V/Gbn
YlraDfYF4N+o8msTwQnnXsUO52qpseJo4BaQaRWub/4KF1ijhDLSB+b7ZkRhlh5LkgpEu6A4fPcw
ngC7IxAZcaKQ46YNd9xu2iU7iSszFq86iY32N7jzm8g8x9syQd1MpUg0k6prH9xSWjGBSfWqDrez
1rHsDsVRkxkYTlQXg0ssp32H2c7c3iGALoQeH8rBZjJ+hhP9Bv/m0DEB0w+pefyTfOyUatg8w+Mz
qNHM4E4qml6CPpQWjKQcmuIB58xSSs4qfi4H7syhKZ4/d3JmBY/g9ndMBeN95QU3w6EsVKpHc1Nb
2uwa6Yj64J6qvFXiGcMDts0ExGcv/uxKDkSmc5DGSENMiMav35f7qDmbug0p/VPNCQnIf9s3lKto
DMmymB2SdRuAO/TIuQggtMs0Mdtyxorb2RXKNGci7bsbhbyoGwoR9ROBuKS52PNiQbK0D5hvJO6p
AvY1VNquWYuHMPn15RjG+FwwPfUHtROBvqJT3elI4s/jtnKh4v3pUdB8U3f3bTiazbLMJT0e5q0F
7g12vzmZGeE+TZWhkIIxMmx7lSbRpVMDqXyaWFILxbdUFKhJB/1LvJ0hYwb9Rx/Vy2UF5Ypm0oQk
sfp0gjCCIIPU2Hu2zna0VnEI71lVv0YwRvBLY1UpGsOv23Hv7tAbcxE101yUzvX5k3VN/MIViP17
OTDDnxEzyLEqMOIwN5RBkm0HPvjLEl/0TWU+IRdsfjxT6Rosx0XpfMYtZpeuGMZGMRXusrSMuQTT
nPgtoCK3rliUN1quyVwC5vZJsmyX0u3BG2hOuXz1NXefiJ8+NnA+SbKhp/1UTM66SCl+fMc/+GjM
QmWBgpSGsZRKAFWslr2MFA5Hz51k6rqoNUfWJveEYsEfBJFPZPDFkI7ReVyeAnMFNPvlxyiaDgXk
MJpKxf+MDlpdbXRllDFoA+vXRPCWB2xjmX3nZ3q/D3tGDM25F+/ABpQXrocm5H8GKXNE3yI0QPio
bhIEwJ/7442JUcOxvIyH1P458FJQpWKInXxRXygqqOk9+SVdCgazllkMPxEm92DpBKVw6GPFqElt
AjzkLHxGjSLkYkYdc2Qj8WyIAV5z/HcGgdTxiP5bVWvpTldaqC+m4u2bDChobBdiLfx9fKoyiVs7
h8ZBvrq+b5aOrWPErbDaX6fh+KjU96TFJjGvAm+TqRimzYjNp6tgYs0rxGKnKkTAn2krhZLusjtc
jL8WajpdubooorLPqsnoC9tCw6wIe8AxiJyyCZM5ucvK3J7O0P9JCCh9PQmwKCSoGZqsTBHMVe9h
Q1yh+PfBldhaqcOwVAhAn3aM/PUi5SkDc9eEWpYuJ47Fqyf0eiQXQE8UPt9y6KSfSt1CTiMeqHMi
FD5o9LjFcddcdSeMleYCoGUvWMBy+0QgeAGEac1Q7xyMmA5vgC+ZaidM5M6FR7XsO0zxJl2dCYon
2fYPLNgdZW4gSIVFY/pEH5k3edCoRrvKpmQB5BznFFxdKc/i7C5DE0VPmoSKre9DmLsMOcoBOUxU
45QMSD/V3w7nECJl8SVmtQzlh+XtaCkKIR/8JwJ9Gu5g3Na7pAC3yk8gFU8spJQxmz2hPh65xonQ
IncMJZKpFPbNj4aKqfqKWzmtX3eqLUuS4Wa/5sBL44K+9XrWFyoD/ZnjaqnbyDiAQRYhS+pfO18a
xmnswqS34P4I37Igi3b/y6Apwyj/jOQksMVMDNjp/yyd/JheNiAB7lJrmR2kYd5ZdmZMVef7ya4v
WyTPOMKcVXDKAwEXIewmWdEzXeAR6xpQvAtEEsscExYQyniBj1T78JrKZz+h3+7gVrBIDCQ2fwAf
d+oPAqbOYU9cdwgnlWZaxk+C2b36P0agasNrbBNu4wGxwSWSj2wU7HQ3QtOFeXyDi+hbJ2N2AcE/
bJAwZEehrZPYCzH0DFHf5SNbJ/0q5jucpbLjIEXB4RQQS5TRKuCWAeIywY3yGnh7muQvX/lthG5e
50lr3qGPbeHKdt9QdtC6t9rbdj3sdHd2CedpQlkc0huX0MTlslnNpLycoj1paLC23XcL2TWvCTgC
FLFp2uZAo8SfIUIlfiM7LMjU6cvDNJ1jLF63n3lxUAKchzA9+Di4XzYcRlcGAjxrWfvc3PHkSJot
idf+aoB3SdvieCM0fCHtHSgUrO6RFTR+jUeA367kGkYHAmgRuLiKBojSgAwG3hNO+HGu+aMWJxk4
yvUUe09+i8r7cb4TXy/m4Eq7r3C+bpVEWBQg6xjeU44w8ohi28vAwsHveAvivkqbRz1aES3+gEhY
lCsfdJ0KanCwzd3WojHqpN182VwP3C7YmebzncwUqe74+rUW4FGnb7zPxU7essJVd86pm7l5XkIL
t1a9OxqUjfA9q4DBXSw0wNAcwnKa78fEGnLkbyrsuCp/4F1P0JXb3Ju3ypKPGh5cyVbdfsAUdA5X
ku58HjCn06Br9PTLlEpcQpJZnJWwcINfTraaTUabs5Wztb9gfv+DKbU/zUdR6W/F9SKISIL17KKM
npd6pQIdblv97pkhZL6A9oy0jjMfJmqjUzbulSSrc52KwE0wgbwz/RzZ5TuzD14sf/zVoPRuE0R6
Kj3Pi51C0e3fF0vxEwtQwi+pLcmdqzXmtE1esD2bikxyea3XZf6pe+fZyd4ys9nfWt/zqH1iYrcU
CRTld0Zdj743Xpg1XWyezv+o1TOuUkjkvzQJXVQsww/MKvbfvSwdTBbkkBv7q0es15SgDUDHi8g3
DRvam5bo4H5gVmAJvwxuRLJHkbmjoHRwAYuJJ0QO/mvemP15HCe4+AMF+b8qrDhm0Vcr1R9BRvDy
sFiQKA4PBFnqMeTmDKzMcbxl3p3VhcAUCdkAZuUe72sbVWGBBmnub7wf1aV20Bthl5Xbo+KrihYC
+zIzUFRGRUhYHrqBLaogpb6bDbkyH70usPdGQW2SEidcXi5Z1zzVgc2m6BW27TUibQ4Qt5crjdp1
YNtvTW25nPHChh6BO3rnRcL3wXUptvPFnHOOz6I0od8QuKekqNH5guJ6BQdhIjAQ3DcEdMTGlJbe
RRoSfrWWn3orV4tj8zg11xD5E1cy4Z4bNuufjdCZXeBs+0Ytfk2r4KWKhzeTjf5/qSy4pXbQS9Iv
4Bul4xPH4bUMHQ+IJyMGHtPsIIOxG5apAZxAoa3bkWv7NAi8MZEBt7n+SofUNSGD+KfWIIRMQo2A
YPBVZBljYodTGqBMfsncHmUttVzhW4x6CIdG8KCTcPUYfNgOmQmRtIN5i6bqsx7VxnIeYAFqNeyo
BSuRNEEZ34cgusdzwKF92wf0PehfGbWBfhlRQfNNmv12EDn135KkqQMWHegmaaoT6uuAKpltwIob
fzLGwm9q+yQI09q+rkQfvx0x8Q9BprQDMTZ2bhtTR/GhzSiCmMo0bhk4wO7vmMXE+ESY2nvklBcv
GL2hQo4f+VxU2pmVdSP27OWilbLYRnD23iqiDmOU64Bb/gmYDgf/GWToOdPVpRjlcxbNPZMV8f1O
m+jxHqrWCoXMFEafqt9NjBN0iG2ZsVDFmYvibv/wMevqzyRf+acevvdiWYTYT3V+lBqcwrkFgQAX
v1o7RGFsisLSyAiP/m7Hmjr29EzLx4brN4ZoX6s3fRPgYSdKbgilmJWHqZ0pY55dgVdRj2mlegRC
Y2QGZyAhKjZIeSvHO4MN3Dh7Vm6A+WgcWFnujtM9hJ+AKwLlYiezvW+AhkNYi5HS2XfNroVsz+eW
oZo+FvWDzRxr7ooV425skKh/7XGLPrfDUcmXEzGdSZ30shwxd6ZYrQXunND8plWt5iBsevsVfR1X
tA1e+DVVZzKp/P7obovDTPh1NIxge6TfhvVCahtv65bjYCy1rfXRtm9SkNQiZFt8ZGLj0gJLN5dQ
Gx8+ng72eTkp3hBJkm8wmcDAHHwdttRFnsXgWgGRshurKHyRAip4d1ymUuYm5N7Ce87LgvIqFX74
tSacRb0iQAinpuVKbzRoWkOaEzUC6a1FG66f8C5VMEP8AIu4zFgw5HkuwdZSty/r5dWwt9Xkc2CD
4Smdr9otAInn5rqdsKGX7sDJieS5E1es7RCXgExTFp+wzTTPxxTjzjU0xqscITofiudayFAauOHh
s5BMFocMGFEGPeP6Azz2vVz0KUAah0gDm01mVyz+UfN1hcDv0k0tRu6QE6F+M43qGmgMdWvzSW06
8wF0KyOC0NGPCgffmt/gUh2UubZPKW+8G5R8zL0t9/GxeF3c7SDE76ADxh6sx6tY9YWwDIylcJTQ
PyEpoIDbg3ZuhOwb9REU1UWALZPpYsyCxlROjE2YwCJV2x9NQazMCoMbU1YnVHJsv5Mt0KSmzoYr
WJPEVAklYWhxjChoI/pIaEEJijxvJ6y5B5GxeGoJ9+U6ffdJJW/3RR/2uIpupCah8z5dvxQ+ohRI
pUCQL0R5+Wuffxd7grtRjquQ8Hm58oBKze8aMt2gqPIAtdiy+0PRLXyCSW3w4IvrRO2xnnOIZxe6
yTyw18y+SXi89ZTJZDv8X9Rfwt+rAiaAOI/8LGHFcZG4c7rrnOYoFurRcm/cafiaf/mhxlOTi3jk
JPNgM+syBeZkiROl8CL9FV7nHeIZRq9U61lbqgqiBiHXheybFpNfxTBZC1cv0t86BcsrpDTNEpga
sf+CLRavQGO26OkUSB3RrZS86dmdOZo8hNDk/cA+L62tG9eQ6j1eP3AHJdYz+IR6x+H6tZoFaVGN
7JXuhtdoelt3fRvdq5Xcn7sjiRMRX+61OWRIaoRfduk1KeRpUlF6uVEMTDRW4oSTlSfckWAkI4O4
e0g7BJoXMTzhOX1QstRhQaGCo/0VlanHRBFEcUZ1YJ+oUmwumfcsG6ION8h4XJg0BcW9yGXOoud1
d2DAmooMLBcaXkONzijj1CIkjjr29tIzdntizjbNTo1KHyjWefWop1bbT+Ait3RUtx5zCCo9+KkK
d8Cz46d9z3ZqfKZXFt0OnwmyQ1Q4wxibqAeFmEmpbrYgOgW+dgk67raQk1B27+tNXSzEkkmueP2Y
ha+MmEHnlrSaWDu/8YyEaee3u4tsE3xOyLHcV4gpUjw5jefs/mMWYykpmoFXRKjDUIIDrMsenCVW
FFxehIXI5fxHvsK6Fl+tGv+FVyeYIqwxRWfzwppEcTK1nttY7dEtarrWf1tEU2jCSI1cy+LoAL5F
eXXdrdqQCr85GHljvxaon1y/idMaUoIou7H3Eq1Fzl09bQ4wPIL7LsbGE09rQNtaOfqmKU6oALkS
mUpFf+0NhhGHaIXGC4oJYM8LhyIGXDesOYG4vcYo/fyTW6Beo3cuWQ+FdwHc+7lVYmUSBFlKo3yH
IEbP9M+l28xr/zLftz6OcNNHu7tbqh0DwMfi+RmBrmJxmGU/1kx2AfG/F/30tKh/HljoNuiF3pyj
ZfAxGPIcD7FdtZuHaFQMh5vfjymG/8yX8oUrgvosHXuTsVFXCB0ZYWQQrz+Lu3u44ak9+m2ojepD
gUZpmAd0j83BDnzuXVHplF8HzUUqjob9xNe9zk8tx00p8zdy1Zg1BuRrPfM9q/GaaPkbi0Jvj8GI
TY4E2V8iW0yb1QY6cTIC3PSUBVS7m4vaqz6BI14yaLV1CSaJhR8VJsKF6lq2SIQhTQzSThOzNvA0
83ijWrx1xEwT6mFBQYn6vFuP60nJOM24q8fPEroKunaB5QxvwhgZ+tmFpUKh3JIhTe3wZ1r9SV01
tieRM4ADuptoENgYL31xlg7du4mw2QcS8ggEMw29KqKoaouJI27O9i5UQ4oOaYyUcGsJ5yJJzXoL
4uO+6uVs5iliW9z9s0UVLeqJBdvmG/APjb0/JmXoM0IHrj84LbQbCm9aKEKzqsGgH6pyOfkV2usd
CtH7r5VE9gL2JcQhDuEyyF8WI5vHCt4+Qg4qecYYk0U8PWj/I3bPiWMY0YIatZG+tktm/MGAcJdy
vD1UeIvS1OAjNsYpfY2eF2nDB+Xgk4hscOqvtB95jZM8SMSN2Nw5a4e7nWi6iZOPR/s8KUZJTSuV
T233/XHEbjiUt/ou487uE6KIyEsMmXc3iqscKagdIIAC72xoDgNwcbrrd2rQANbFdpNCgLHWExz6
WQ1vDa/zjJsY3iHWD0sjtwTh0LcYsM0nHLgiv3bsd9q3rRyne8dYUxBL12zB+UraEDyD3aVIyeQr
Qpx310R3tJvlT3IH9RbroLvj2HobNARmj0ahJm2E7Ixro1gs/WrWIE0N3sZnsSzTQj+UdiQ4aEHw
2eWB/k00xMtnc3Yg8GebZ1tRGxrtjRmizX/C2gn16mkJ+wiSsk5wwlWiKSjVT3Nq2Lubul4zbk1H
VO6GDooz6vP0OveZWHJiONe6zT4/6d5vBoGdUATjDW0BYiSS548+jQc6Q7QZE4ioxCDvxsET2jly
5ObHeXOS2pZNavjeeb6nshzX0HBZCWmRCnUFCCsCqFVYPvIRNBjau4yJb4Ei7+8fspOGxO3yfmoj
OZda9k5V+/IXgg9s8fZsUQNDcAZ/N8LzOtmNAw7Z9pw90QLUl+HyZ8k9kn0rtsBUpRRBDHqvIRV4
AGZHP8fi9kXlcTZshktQx3dBlT9aC9ehyvogYKaAKTEv6xNkmSQYSNm+ciEhsxbtJQ6oe+1fcM3T
YlgX4xTT9kgNn5BD4kcC0MrdnZD6L05dItE3jlqyvGrXjpws/CaMfhk0Q876hn+Eyccq4q38WciA
4NgsywZsG8xsrXiOg2sWLNjlFuZdqMIauxQHgo4XyQ8PAKZpLDKFYs5Denxc4AuIYEovFepbJq01
5SazlqiE/tvciVKUf7EfuvOA6NcVH8lUR/aIc+xT3aPOPENphO/VRwCbPCekVwTx9UduRIuYayvi
sCsz1XN37ZJxlnE3JQE/HjKPPUmCAZIPZ38dFAOrAZX7sQJnLMNoP9U9OHf8Alxkx0KyLtsF0soM
jTiPApHJn9XiBdemF6XLVmFklIs4z8yMtxDQP+jk3DHD++DiWfWNxOSYA2adEu5KqtmjwfSz6pNn
I5HZuKl4tUx0JFxL9lnuWFrlxZwV3xJF6UEii+H/0rrUxvCfwhfJrzRgWDvwssEM/ZPXo95UayMk
wPhq3AS034JMw0O/BwEDbgu0acNoIpJGnVDajLS/c9xaD5dbL2lLxZ3t7a5/+s83vvlt5TFHkh7o
CNhao4/fOVZ8JTY4LOozmpzfpSFmyIpYgSD7Hzrd2xxDArTYiyXDzeeOfR0eoak7gxTiXbQm9gSe
rZFwSbbwnTt8dohyiwvsbUDcRVeR5oGB5XUkSsPj2ZMHLtNNJ+4VCmCKNvdy/Njv+lCXr84PpVnu
qit/3EfElxafpaXV2OVWexzj3aEKnbWgKhvIUrEJl02YnvcBUqaFExK/0BuGxFiIrRRUtos+XMHu
MvmR6SpZL9vBVJpbPHO35zJG+9bzbLjCRwL/+/OcGhcCi+7L5Qo4MEhR4MllORrJJMa+hHW7cuxi
yp95zbmBf5EvJ1vsfvUTATVu5RUI24S6qMvK0Jm35FhmKdh0gROUOPfmCsyDGv2ZE/PnHXYeCcBj
uVWmYzGbHzCqRiKnT2znL8ws2zwnUCKjKxmzFv1mp0GG9ETyV01w+ADz9UbRcUO62/ABfM9R/hUj
CKdh3apt+2kWv794bYe5DS/HfcukecVjc2E1ZxGsxOQvw/mHy2wGrUmReb5WG7vv1sHw8ilPfZqA
ZpSL5P45ydTHdjJuzPIK1/IXKXmQT6a7ZezizjEnMehV5aEkY3T5VDJlbehJUpcgb/igAvtkU0oE
OOhpJ8p/R3Yrv1emqiffGq59ShxRqvjHY9J1HIKqfPBtgRlE4ZgotdvGI1WXuPwlLmjkUGsvLJLQ
++lmCfvzhnj6zLCMibzqexr+z+gZCfpG0ZtQJmJXxeIfbiz5yufik0rYZXJxriqlPZFnuS8ybNY0
2izS7l+L2Ak6eH95QSPg9zm7um4QPo+nhp4rH80nGvv8qO48SJBRYZGXGyh7XBNvhh0cKKyUrO1h
nWTYhpq3pn/jrKLkfXrZYhu5/VoiCaxT7EqCjkvWCLDoj+jPFVnod3a3KnBASm3ZwL90YK8MO2mo
Wt4WYgWw+FWHNjFLnGXYuOE31GvjVAmnJe+BGohbRClF6+id+TMMOGBq/Bd7QtTWwVWjL12eKjQy
zSAPz1hPhF8/vv6Mb45Jh+esg0MLpvWIEf4jVjwmZAXukWRHL9njYTb8qxejyO0+dZNweUWhFOzw
RqiiJvtpJz8SA5Gi5MfM1d4UqYTKDQys9+YzHiglQeVMqIykjCQdcf7Z/+qmrLYb92CvrX6pFxxk
V6TkmWBgNI1K0bQMzScARsxNXbCdnFmlnOOFYSDaw1pLVwqfaYIxtYUE2b5ZkoD/IJRaG6gzHdlo
FlS37OqVIay6PTMJza+rxxjOqICYcb6vOb+jkCq5DXLYhu7WogJ18gOe64+Ae5CLEyEsu1aeIBaQ
NzbN56f3eilLm7TVQUbkRvvM4nrENoIH265TFN0cuNRR/6j4ZQlIDLgHaOlqq3sQQHVmWm97A9Qg
BuRsvQXat7oFhFuRfwbLO7TRuIZbw1Zm9O6T2DkJdh9SUyqrTUoz6j4AOPvsh7GOPwG8sd5fXcwO
Jz5UPWxIzBQ0EJCHIEkJBSuOQgL+PR22dwLiFvL818FAdeNxW6c6kHHwMSrN/uqVXFSXEJAoRvJ+
slazbqwIWafCfWHROWB4GOwH5ooMCelRpjSm/l13gR+3f0RNMmacIkO8QV7X7wJqnXQP+cRpsPzo
kqxzsiF+Rk7sl4AzXGTyxfKnI+ZExphhkqw5jhLINgPWamptfrHS8+woSJA8uS3rtIkqHvxHosYY
TmTRiIjkMg7mSz09FC0GVZAb5wx60vCP/oGV2MQmNx1tZSna6np6dhej8O0Dt+AznV0F1O/u+WOU
f4gPltJHHSVvySYFB0XP+Ltjd/J9NRfEMOjVpIMg5T5DcHyPLK1U0rdld2py3xOEelUPhJMt8YQw
bowjo/fdd6MgYqz3efrTrqVS/4R6pBDPtDdz6LVwvoYppgnOwpby1v5XhsjbiwlqYHHn+V5I+c4r
sQQxg+ahypxU4RIPzKYMICkfetTIG+elw9RFwmf6rKMmNBWHROtcllDf94IN63ZZquqoTmLVOaC4
+qTrBEErueZDpf3YM5PlB7Yu6xGNEHXhfkbQEHZs3Z5IPtDytJ0kXL2MrY+ADDAA7svxeIGbYc10
ffi37FoTv2T1LYv+1z75dH/rcRaeD76W/F1RpleiGfyGG0eiLZR+IGy75/uLpAfea8ZNBjYz/UkU
yaKw5U3AyR4rd3vhOpciXh0QFkb0RgykR7R+vn1MsyvPkqGdF4x98Ze4Nhap2fiVOGoMF1D5q4Hq
HtVq0JqTPOjXlEJD+HM/W9arwTc4M48uitFta23MCOv+WQhHgaojFAIO0gBqvyxKp7t4chxyKfxb
uu5y7mFiXRtlUdbeepQU9LzHMexR2aOdUE/LuQZmqZiD/scZXvh74auHHG7c+4xqFdHj7BiqXlLJ
ArmrNaVn7D80NFJPmzmtjGKbFDGvvLjDBrUdZGRQp6ELXZaB645BXinzbsmweMRGy2L2pyllS3Lj
reaPPc7hcQ1Uyn8Z1iYBWEsSR1qI5OlDvB8ql1U7krq3VGSwn8BOqjC+FscH+KjeqCYxMCIIKvOo
BJgarXsV1k/zefV2pV0S4hCurRYWHkqxpsxMjy0ZMElV6hQA/xpUE2VtNMZI704OPd2DjvLHvXGo
SGdEshRkVlVPUrh4P7nySWm0ktKITglIiqUUtYGpFBPWLWogToFEoWWOTuXkrYbXoccPhRxFITpu
yak+G2AcBua0wUTNoHHwE3XtoEOwPEGp4AaxDPhkjBOAlpNMMa4VBDjmsvXY8rYonG4Yx3xAjnom
MlX3FzRbmATinlDAt7I1UM5pjfImfeflxKHVteiFkB4k0scFTlq12qH694YL6nsTTKIYTUFfD6N7
2DrlVoM3ENNXNwrKOvaqz9/j1hrW6kcDPQ6rmFkX7kRRlK1XZ3vbhUKIsz6SgaxHzCNsc1UC0txC
x92SVyOf+C4KCKK8Yd2rhl3COMnwubCsq4MySVXhlxthhhKQBYoDhCMYbQ+gly9fEfSZakZUKme6
8Y5pTYmhZEfcQScyo0tRP+1+Av/GS0rqPGMDpI0EXkgIPidxTpkZktP7OSfWKZTUElgw3RGoGBLy
MCno0Bub552GUlz1ZkJ5/CvmZ4cHvV6tcMowRNoEs71WlWaLqhBpj58shvxSFjdRFUIDs/tdEYcf
UpFTYuFYAyvCxSP9+eR3MOqEQB2R+M+PmDcjyuV+eXkgiLleRhFhU7XXveIckP+BCcXo3zuPNXhE
3i6OYTz9QPPH2lqbt2MEwSnELKdeOXlyRoQ3XABRdg/VrcLef1pLbaLWVIxeMCA1DHD5xpZrPQKd
zAynn1q1YzSFhnlEnh0OD+24O1+9CmnvXGMLiMbBJBDl2hjqm7sghjDNqbA+IzIQozXXFwR5gp0k
x1aJ/Txm5ZRHSAP4au6ngVMYr3gp2wNDSOi8cV9jNoUh4cSC9pKAjXA4af3BM3Z+76udMnRLJjOI
X0eXzv3TOmRm/8v/8npfMDk4Vpq8o6oV6BjrZeGkoP+dT1Vp4O2s7QhvDgpi89icsUEgtrc9M+mc
SoIB7LZpGsiYTjVyJeISuer9nIZFUzAB5Q/2g3gND+6NhFip/KerQ7hm2pgtaYFAD0Pd6wcvz9qx
ufZJROwV4E4rbM83g/VKr3H9lbRZYAw2cHhN0vV66Y0MusAmN0vIwmakYKlPrL9Mm7C5I+KtivGz
nOCmis/FjPpO5pSSiNYgJ/HJ/fvweF/rUZUUZPUNPSaAAyk8XnQDTzZGCGNdznJISW0aU5+rxGFh
mrRyanfSKsmwp04nVD3hMn7Xb8j5qMpygtOIY/QuAM+/K035CrWGFOXZHkYDvMgoJ0zY0u5IpGWZ
EPxMrJQC1hQKt9qsXx/eDCZir0SEVOO7B7fwqFUt91zouMX2ILj9ftBI01aNnApqGJHEBk1YyODO
ynAg+hGcI6uANlOhxttP37HPJ2DZqRDur9yQtw/vvEOrQXAAYeO63bj0K5jUykzEJUnNhv+568Zr
2hU0PyniSzutwE7/HBK+YBp3w6I9HhaFGT9krW5neA2g7nys+eDjl97oJhnYH99Y8JL8TgKqT0Ad
ej908l4xg7iA4WQits6/IBoT1vebJkgfUIUVpv7cHLwVsmyZKwBLfnSDIre0+ngErsDkcm+vEboq
OfOq7RHZtCmS8N1iMq+WQQBmqIjQ8cue2cMGCWkdmp7nkgKsFmBPXzMlGgLMIiLRu8bkUdAinEOM
AZWM/XArxFu5SbjaIyGVsQ43xwKzl6AKC+H7alZgmvWXe8vdS9DNs0f5oLuqlEnIDG9rbtJlPoDK
1jKBwI2a1zyLW4my5CQ397FoWTGGRGN0apc32pyp/lRpx3j/+Gmu1wAREQ92VqLPEAOhNFgtPR4t
nwSBQQN/HZ5DRGhKPD3hx2zwPJL2S5HUii/ABmPNSi/qaMV6msmAQaY/5m7BmpehGJhgOIJVpIV2
6ronaPGx4TUoy6BdA2dB15y5jpKQc0jo7N5bd4oLYXGqIHqEKI8TjY+NHh4c8bQyHlETdPAMAbb5
AAPMknhzkjSj0wq61/gjAuLoOx69phfDCcx2pAMhvXMd8ktj8/HA4i0Q9IaGU5jJyRmmWklMWbrJ
snhfkX3PlRNUrDQF83wHMs7oh4/SpydjZJoSm1Mta2vRSVGHIvCLGb2D0OSWhrNoypA14Fw96xvm
dUUiP0QoG0woqFO0WyUX5ENUCM2wfSEoSI/GmCnhUtooyVNgaTV5UICOWGou0h1JFq2zmWubSvCg
9b6sz1T1DGTiG4zHD0QmbFmNNB6RB5ko3y+KbsbMalVnZhJymFCY+6SNks7SUoqwNSQeE0BWx2mF
5/5iulQbH49QG+4O/ux+VJwDDHAzDgfVp8lqwLN3pM34dXG3D+MIGkNvmn14O7om/8cb9LWCqw7n
nbWtc1yLju0WMuqGMZJ8grig+J+8orvApA0sFF0281itYITPfxHUgjmWSwIG0XJ7ew9L7vwYroLO
WKiIeCnGYtHl37VmDQOcVhQ6pieFbmmTMytB04yfl8nHeB8rNRCmUA0lFAup60G4Z6iiOMMfN2Tp
cazcKcg9JHBnVkl18E4aMoVEm3NqKD5FaDGqtZE4PKWgZtFLeIFKcQYsnSO3LjjlTrk9gkq96/ll
bfwSbbLhSg388gDGlmBar7VsKQUM1SE11CEh8PQPMMPN9lxLn9L+3hn2KqoJ07WEp37/CQf2gQL+
tFWM/dcYr+MApm5Zb4mVbMFi+qVinjbaO0i8hjmRTLD+Xi6YYB+ZU+Jvgo5RxE4h5uDnF/gdnOHr
O5H6crxA1rPDxzffn/XR5R0Nu21xAENVKejQtIbODXrkHhKUjGeMmXyfnjjloCjY3SOkmbWoWrou
84P2m0Ap7X2YiFhJoiKXS7ITCHo4P+pxluvQ58syG93ETTO+sOthkxCeTU1BSXdd0TpYTYEcSBfO
eJsSU6L/K2Ryf3WBPtNnVVSyzddW6ycid1CK9LddPEtwz5UsascpKkt/o4nMEQOgDydOviBcZ252
TaV6+GOhQRJIw3eKLSQO+JaDlyEbaADZtSDSSDGZvgdwXNlbzyUvW2TzU+Im78woHO3ZjbMTfg47
gYltdYZYfZEzZuidj4oWlIS+SDvvdEqwGAZYammdN7hbrT99Xvsr2IsEyTzi0IiKkl+f6xqWCvJK
4wZbA0ikp77erdgRQQ/DDvyBezp6sTy+4ur9UoVrwQp9wAC/N+Ps4YtXh4CGjjIFkBdyggOVLTrX
sObm8QYuiuLwFiTOM1XpEiwYtrQtpl5atxwSS+BtZToM7aTMWBQSnWB5WoeR0irONUOR+CABNz95
KYTALY8bXBMLoDV2HDp0BOVwb700nF/if6nBoAnray8ffUqVlWoYer8jNCYmfSWaPJjxNNkoDq+t
Y7I97oayoeZeMv2X7qjZdJ3ULQ5c9674a3NttX5UOsC2VIbsTyjrZrbCeHIY41uG7jxjcKnr96Ft
a7PBJeXJj/A3mhL2LLzjWwu10aeu2Pim+rmggoTg6Exy7aP0cGaCMUMzw8O+desADxjHV5A+5Qyl
NFlxYN41POpjyRGC9DtBQR9MFhR3obbAVcF1kX+3ovDlXjTB5iw5tV+ilrT5cxuDLF8AoLdW2Sit
2dL3SDS5QOE3qwHe0EBY1HZLONs/0K5X29mEusOc89RzxcEeMmYgy4cIcvXTzVQ1bk3HGGzEPEu1
iXOIdD7VgACqyJqtgtSRYspdlk8VZHhwhBhjcYQTJOLELXHawXcd0AEidvvhaB6MR7Rb0+Ld0Ske
o24qFqaMD1agxYkXMp9g4WzuzhVCjO6awtjf7LT7VTDoDIrvfFQtstfqt9+Q2RrXdPq5CN3E3CRi
gJ8loxG6lakb+CG6ZJ8r/UPo0duz03LPyCEf1/sFB4L+bfol9rjEFDA1l3K1A14yh/gGV+JNukTv
lDPemUsUHuLGuUitlx8HYSwvSw2n4UQcT4QFXp2DqpPJFjo9YQaOVg61Yy0/Ie8LH8hDTjEfr/0v
O/vj7TvzfQeBRIVeFvGefnxl9zZDVMjAnsdZsy/Gbb54FpjYXMoCjhBPASAaZhzJTn0GPwDSs8JJ
n8Dv4cNP92tfxKLtBerPMF3oPDR/xDWwSJ0+oFctYPNdWDAO4h6We7rsm9CgaIsnyy7vBQbm34Ok
UVixJanZRszQgxYs7hzcqZCODAamgA21KxH2fEvMp2MMDhqxeFT/ASskLxFloVkxsw596N4pKrSU
quuyF3MnOLbnMn9B4+zXgBc07wNzwQzo2DvMg7vF/bWzS56JZL0N6L1lAQ5voHVxbo3wl1mOTu/A
UNQV7cYNGAFdimRA/6NCaaRiPQ3tHhWY2QoR41TVgsaJt5p1refa7nkL99LjsdaSVUden+Uw5JgY
axXXiyZYUqSbjcX9LQ6+vM4AX/8ZtKW3GoNEWxXDEGyGhPzf8uWYVCD6f0f9tDWbtxBPISJFwJYd
fNtIRt8BVplF8zQKHld582cKgp/R854W2GeWR1a9lVGNHiTwKrHlHXXo3rBGIKq2gO8K5f+91Han
mNnWlYzUfgdZLuPlbC6pvOMAt6Hf4Sd7LHC41RFe50N6fRI3SWEHGHeDMvV0I1ReNcbByMHUu40C
DW7jcBvt2/Kc1HS7RnMYQRKGYf6+h+TEP34tCleb7hpVq7TNArwePcRfl8uvz7InwhBFRg92so1N
XBfpGJw9arZuL2QUzU1MgejZgYuQbAovNNFgu+Wx+x5t8NWA2BAO3999zMR7GMeLuaGqSpwNx6Xt
KF1CrdKoA1M8OzTepOQY6fbOZvsWGajgWvqgJQwvWwra1Vcr3deU9Tf28/PBvCh5S6NO2xmC6Xud
QGm1baAgPxemXmlj9tHJCipN/leVu1MSzJexJpObY2pNpgQIDg/Qrsx5mKyGW0n9f45mTIsT+m47
g1dAAGxFZhDY4wNEvMaSi0KwiWEC5/TBwuUJ3rT2LsEtkesEdfx6VjWuyQxuBD3/2bwssbkadyCy
bV1dTjxfC5wdhnx3UQ/zxt/Cx8N35FifkSRvFLWmMPZp4B39JmmKCgJGGoNMx7ABXsh4sk4s39ed
aVfwlsQ11EJv8DU+VlD/YT/2M6YJ9tEfzA4ev0WccpnfxXJdVU2wnOgIUGd94nAwMIlN5bhcKFHt
XP8DAt80VNLQxFBw7je/Y1uGwk0xU+NnS/LeZPcqf9ukFihtpugj4SbqdHU2TEhJDSSU7z9NbS8J
UUZ+CGcuCPxJBBdN3UItVXeHGVkMl6oogmWcT7KVQ1oqftw4sHLPHmW8pcyiAtPqAZRkaOMzvcbD
3zFpxYX5WQLO+6AsMfB6j2nV+i6mzXNbZtgjjBIbIkRT07L4Xv7uFfd6d2OCbgTawXH8yza7TqP4
x14Jbc/LaabZdpUxTHQreaSXCohWssPE2WJrvGqOk7xMHysESQFfvEeKWSrP9GXUqeOfYDjMCVke
G+vKrmIgnXE+QCglkG9c/5tDeJRNdNIyB8OisUDOeAAB4vp8G0qXj/hptpUycgUd2xIpmjjJIUL6
AQZcmdVIukHB04EwIdf0M+864zF2GsSO/9TsOtwx3m1ZaWgVg0+j3aoCBBwdhAkC5ifCx8SyD6NH
+l+AlxJRqc0bIwK9RYtx3/u74rPeQu4pVCQ6KR9zHqXOlXJVOyzPcx0PWUVL57K5JE4isXRIeXkW
5iGZHbnXTXlfKPqnyAAHLHrY8j2FzXxJrCK/Uny+J4fBUDDD+1JytmPpr2JjWsTJXKeIQe4IGBDh
1XToORMAdWUQ2lk40YKQAtg4pq/zVMszBvjkOgLJ/l2wpdxGyLgCk+y/0WzppfjQ4pbpehL1i3yp
KJAPWfi0k2Urv3eGyOcy9B4brOizINQ61Y58zLQ4gEQ6otGxqImaqGcUjIxerSuWWk3TXDQ+CYLU
Swh7m/Dg0qlC1nkVwXc8Exb33DGtryWpT5F3sqWrnJFGpvE6h73ccNQq1A1zShrMAAiOWAuLIzc7
g3ZWC3ZVCnpNEuY9V5MUbdHzaw0B3i3H9RGwLE0i8j+Z5SWE0zrLNN20YRVxuxUn/9JjFWukiXZX
rChxs6BmJbVhuN6nb6WGb7gmqBm2JbElQaqk3KwYnB6clTGpDadEJ4Ri5+A9X6GT48lMI2xrS/kQ
HmtHK5lFjUX3Hyt2m2T5eqsfz4c0NRAmhgqBnhxXNKERhN+3G5VQ+n7zwvqZ8nH8S8+4WbXWxVJ1
kS6A5xqxPA2LxuNGewTp2RV+Dt6GlmpIaUbSB9qzsh3wIOQ3QYTUicW91K4MzUeCwgfk3z5fdWd3
tQlDC1LsmKx1kJwvGwqEZmWVI/Q8F5ZubeBQErgWGAFyixVTFVFiCf2JQrPzitC4UzU83SP5rSBY
4AynhguqTaQqRFf0zdMPedBt4NzmHfH2IawXqjjgJw4nNBtzLh8nI8jGvTu415WtRGiod+dtI0js
0QgB9Ba1WAO1NpWPS3YPGfuaPI/Ja5tDzNpp1zugmabazHksOj8m1wxO7uiboHlrSTp5Aoxl6emf
PXrvsjuGiMLSzsEGyy8S3nodWJfq7ybkHzKXhGXI1tQQ27T+4VIAMwWuAMPeFzGI7kFujD/DTAql
RCE0Eef/tYXzAATk7PPXGvfHmo5NcgqXbb9KapKyHFoz3qN17NStiFiuiIjPghLHmF1nSt1dltbZ
i0MictWHUCDUthtrbPNawFHeWorByMAb/XZVLI6b+cJrHzyd0CLyR3hR2JVDdB+fDCBiycBMBG65
k1gvfQH4l9kju8Xka0nbwAb9qXpVptUQVtjQRShH1GFAxePW0WiIj2UcPqtK1B8kNcmJ7RxKEvKZ
uznpRtiug3r2WB3BCHynoVPUemqns8ZZnP8lEv8ahO/gwzXc9nS6hCEppteQ/FuyLOn/XtkCtVOH
HyFbzrKGSuq+Tw6UW+v9EKRIu0bW6rnWWA/AtC1P6LZ9Re4kq2cYR1M0JxaC4HsXQGMZYhIxSU9n
Zhd2N3FayUoNf3SocVmwp6eLPQuj8Lo8ipIiGnmSrX+85OWRWlIsQpwvk8z2d0L805lNwDJzSu6M
3naZI7MN7mN10RuRoRVybKlqlkzssd1T7VndtGFpw/ktWVCYgsDekXXDt+og+eB6AfYCeWkelctq
7eBbrxiGcgQHj/4zZAfUnvfmV8xh0dUigNIGQHs0D7XyRpi73gq0WOuhx6CwFuUx9Hl5rvDytbBP
owrIlnUp+MIhlEKw7yGeWxxGafkZkWwO6NDVPbNiu+UyOCyxJJG7oWCC6LvVZ2KUiw+7ttBh52+1
CNeAkSPg0lhGvYTwEhLRh9IlsrOuHQ4zTkH1P9eQzpSKrih0NynCwBC94wf4sJukwma4/ifR0cjh
0ULMskP6RwGp6qu2DLZSPDfMRhWAY7cQCEqak5kMYg8dghMaOZAl6Ze+EGSZToPnJi/GonS1FJ3h
fogXssdPZFeyGWLQ2Q4IoRojbL4O6TJZowblDHXtAqlBBo9PU1BSeqN7EYjULJ5nVUhlgtEs1Vds
Zj9JrBI9i50EPwU7ns6Hr8Hu/2WUqdxOXesxvnvrVl7ti5FBO916UTFu3lLK1jECbIH/OcB9Sdtp
pLVu4ShoYwNJ1sPu7burG4/TtMho+I7qAjmgfpUEoW+0uz4LVY5KZ/a8idhUW5VEUJ4lR4Mz6r32
TMMIuUKsApEHdVWhCP+cSPGkFFTdCLksJ64BjsV0n6yuTG+H6nRnMIC1jRNZGnWvDtE7id3eCL/1
0+icJdioSB8WWm6wULI6SZcHHxYxZNaWGC371LWITHkPs5UqUSmYhJyk6tqWhfyT41rPX/SbvnkA
69+s/3NlLW1uf393b3p1q7gpt+PPixgwQOBqvQjz6B1Pd9ToHE/lnVfSTuM3e3QxyDfBe6vdHia8
RYc0uQNMM8iUd3gGvrQMFb5aGX8nH40SvetZ1aGZFUodSTkoSRRgDYGxmZM3/FiUWWV2cZoYoSpv
yKSey5MWd+g86s3bENIfvJuW+th19JgMhRMxoDP1vCx1bwsC8hmEZaoM7ti1BMryHtVLh3fIzjI7
16lly3NGTdg4FPIW2KmJSyINFXFcq3I/ASV3D5n864ZInSmzaoDX25sgHY4CZrltKrIXV4KW9GUV
44CGY8kXCzYpaqIpFIfLcuVndUtX76RU9Lf6RnutTHo5aaOEWXDhxL4L+TgDkccrnYCDrMEUulAN
2uV1li0FKZ/ViqbAg1AcsGd6X4SZiDCDWKj6biftxCRZ/pSGaQe8cuLF38nt0MF//XtWb/8H0nMf
kl3g4je1WAfxbwR2q5slFSBN+43XBJ5ry9wA/0TVnbI20reEsVOCptJ7jmRz/+yfsadbND1Kqtba
HafP9GAe0lgK/uuyec+sH1r3FLDByEQweNPrYs027iBS2eVCsRYRfWTMoVt4hIoeswb0GkbvqVSu
2UjA62vvpkIfeuV0vmqpfLQR8Lb/pe78RPP6qNwgJhuxycHHcBOy+9/lI9XjXcMpp+5GL0h16Ku0
mArM2IRhrY6EDPo/zQPKHqmAckEcy1oIdzeRtPpWwzqu62APBJ/INK5E+1Bq2dnpjD6WmMAMI5zw
KoO6VCGSPKqtlVTN0Q39ypjejDJaKV1t7OSaSbxapVxsV/VL/nxEYdLecBPQ9cJm47BFAj4zV0qD
f6sd3Lburiy7SPAeMq9iXBIRfpFr66P+4JYnLHlhxGpOUR/XxHe+pq+8lKWmhYfCcY18Hz9nfTyR
upPz4H/w7YJ+afWF7OLo3TQnvCJ9JI26r6IHxaqtlRea9114O1sqo+HT9fN0omiqeao/vh60jmY0
bdBi5Q9+t3hNW2msz5ZV0c0pzGs35EUWN2GOvu0AhQzaR0bLqsNnqOPJ5V6XEdAyL7b/cmOz4Jgb
lO+jOhAQkUdkkBUavGp54DE/0R6YVNyGS5dhWv+C7tmvxAlE8yYffFbEhGT9Ia3ZVkXilATWfEEf
YUSBw0Ssm4lNyEeRSd7nMXZbGPkX/BTSbNcrhpBCjdnRJtHkUW5iHO94FvgaMlCZa9M+/yqqmKBN
a0xrKA0lVybiAeM/4HrxyaFvmvIPogp2aqU9kuAjtNxOKHArK6niwin2U89dL+UU4vK0/zUP2X9n
MAON80qH2hd6eygjXnMTFI5A/3DOaDzE72Ys8cYgovka5pIKf5GOq//vVqBznqUQZJzziwPRPcMZ
5upzsfv+wntK36ckW+niERfnh2IzL+zWBmady3lJdc6Qwl1SlcUkvl9CN8+QddnbVH3CtbJE2eZx
CHtLlmVSxGYZj5tQMFi9NGYB8LnrfEfsfcBfkbmI8CGRhD6WlAa9Wxnygm7fcT7pKbOSYX+hF09L
Zlcak1pmF2ooDbQvCTQxjUnVLDrl6/FMMzI89F2WgaZdNr8gpx2ABnLhMRvS0/SCkGTU0jOPVUbw
cNQ1h++vcoEFpWg/Yfmt9G8Y2i2l5KpoFIwXvC9ZCLh21ncpjaoaX2++o2nJ8r/FkFDpJYjJNGTm
J8gOPAONZTsFcfXzMv/+w/NYHhVYJkfIoGQRKQtg15v5Dq9gUbsdP76f5Ugz7jRx6Ile/Q06tQNk
wTKZx0luRxDoCHL1mrse58n9e3wxN5dtdzQNatu2zAK7J6BMFiTPf0V+5grDS1x5agRPiuyZKx9S
LAF3WUBU6AH25TcOD82nT5OqvVSxY+g4kKHkWTpdI7J2mU73Fjc4F7MgWt1dGRboKK0X1AfaAvoI
2GVKyFk0L+4Tz4EEsTvnMU3s7ndmube8tlFw/9lm33nEWwjlgrTZB9QKsEw93Kmk58zv7E+wMott
7ZOJi74HrPSOv6fhm1GZNbYarOMRrEY4ARTS1UivcIzh3VOMDC9JHqbnFclmcsVM1pK+NO1dOOWo
sC1RsCh8Bogn1nRkZEvgAWtOrlUa61ibB+RAGGVJRyoHZ02V8BDdOSj/McliFGFtC+kYVJC3WhW3
NQ2Obp/YPgWXUCvqlPqW0i0Jopo5A6LWzxoPC6TuuJUMUjEOGP9Efvs8g9jTvYb+DwVrl5BuMsWu
AvLg24AHwraC+gN/1YA6YcpOYaX357REAA0JHyp6OW6o8UuyNWNAdTqoGRQQU++vQcJPK4Vf2zbl
6KBdw/r72vy3rKvqfsgbEl70L9rw1L0hBl2nfnpk7r6SceXB960wnxbsUcrQI78hmvz2W1mRt/R4
JUQFGGYhnmwp6RUz4lT6zuhml9ZK94Ho5JjSzkSFbJu6sAspOMkgvPQ8VPLYPqiUM5fwzuhbMt/X
WUvtBNLGCaXZ4C4rPae1hSDmM9H1HyvcJ721YdsUok6SxD+wDzTclEqbJPl0OmFA+py5lGMT+rKd
zqGSWHQt+lfFxxRMO+AOFiG71XUC2fL0r8ilKJh9H2uubyFeB4ATMAso16zQacjJ7T9qyQuxy4P8
RyiuRE6m/IRFv2+aQK7x5gCczUJbRh52n9MjzzA0wg50mBQUp0qv1ukcpvUxH/vnYTucVe4TknVJ
Xz0KDOt9RB73VbkhjvBN8UP1Fl/t+mwDGGxANce1i6Q4Bgb/y8fexstYOR+q1Aq45nSfCp5at1Yo
NgCixWnkHzb2GGUlg9O/QOVniclwoKnN0jgcJrJbxZFUUrQ9ugFEiji2yBBYTVlS0XZNWIb7l7Cn
9OmGPQzYO2jLcjRQ11a/nPY/dyJrv6ddOFfpUJ6KNSEYXIQ/259Oa/LsFB2Q4NJxlzbYtknTSQcu
Jbrml+BKiyFHrJeUK40HFIuoEJJR1Dwy7Gh8S/agJnGArnjTwNOOAGDKQhm/N9EMsG2APwxsC23b
ntTX1oRip8SCkilXLxmPRnOXCr2uzip+ozxTZ7JspwoY4Zig/ujALWRybUlOQQzfRZQCWn0EmO5H
bB47kRtIWWslLTBYDdHD+PP0I1kjavA1bCNRzMniprJepC0Jn5B/QUJlYAhb1ZA/Iphwzxmet91X
xvkurJ1SQ5IuZGIfeGNyA+9fj5E+N4WMSz+AIPY4FDnknOAVERhT3iKH0LtXS/Sc9ANBOvgu1I7g
LO658+4but0+i4x9bl1mUWXNHR3MZL0b9VUHU5SytmygVpZ1cJJEkau0THhVd2ovEGUg1JEljlJM
8gkWqY9Fw1MQ0RmMgv0Ne9nVmOzixdndQqFr+sbBWsKNl3YQ8sjbDiWjnseHgeEtjjYol6WCt6v/
6LiyXawNjG5K35EIUCBekosCNHUdUPnjKKpDd7CZm59bd++OOfGEDQez44EeyjbgWXt6suyw6Fp2
sBXX0pEQCj73iAzqvjHFBimPD9kpoM5cCLhhXJaEEs1fGv2d4Uhv1iIPmNcRMobQN21V4DXjpzgR
su0xO9bkYRseY0kpqS3lKnfC+XWrzoUrJ3zPz/mSbk9xGe0ThKMp+m0jBg1prYiyRS4qjIt7alnA
d5BQjclNkfjmtzlHcjsbdNS82xrZn8m+PUMBSJMUglcLaCmbOD6WX4GXdm54NSbiuvgExhdy3IPc
EU11N6TR7P9D/YEWAl5yVTFUSSPlGHOfsC30EydHW1JXUoKnkPN6YTd4RPry/wRmer0aF2tqaxeY
lVUL9NvB5QCFk1qb0ClQGekOqFJ0sFicLW1onNV+h738Z8ObPVNobA20avcV4TX5fpaPFM/i3Kqw
MJq6GDH4fJS4MQRDhsFrTfKnA7DQZWs4j0FW/Z+79mhgZ6VLWWGeKLW9GvJyueclDlGBOw8ZujVq
vRBRpDGe+slOLTyblR1z2+h8RNvlqJ3pPMOL1OVnWYJSzExkAtQrfKMNRLTtRucol2PQnfABFfrz
1Iwx1YwsuWKN+YqxmaMwYf+hhZmyIvaD5EllU/jKYsVgykCopmRqQMm5aOiifS0uvNoGCUa8ek5R
08qbdEbiImHVI29DQV764iJZwd4W5xHaRraUfS69rv/NCBDDVCLXPA/QDR+ybS5FP9ldCqKgZ60G
CNbI8NCsvSe3pTpxGmW9nK/GHGBcqepZCKTN6zRY1R7hrM6AwSUjy+2EQrBJMS/6g/ce1kmyAPP7
8mT673rk7cxo7hpgiSbE0S7Ia0nYnoZDlqgwPFI4oh6UycxyiOulk0jGsZzrdTt0UNLOUxbJy8TV
uHOlJKlGpfnb9uN5jM8THKXdnoJzBTeD55iWkZZYJIvgn4ux8SpV5S282FaIYYyoOPbxbXl8oPEF
ufrlQUDfuNmfWVYb1CL2O/FdsXq36UJFDyCoKY7Qyz2mhsvrBhCdSvbIJ2dAE3p29vl0Mdf078Lv
ub77XCjsfhYpz5I2uCFhw+Yi7BYfxSHw9unKO4JtnDY34xFaZgloVTL1Dfb7Wl8l9qnlkba2kEw5
OlMSZxnsjGCPTv2JCUiKNySXahnHRaRf5Y6G/hBFB4qR5hkLy96FvIbYE+1bw6OkAgSt4urrBbXi
ofhMOdQKFYbYOrg7vW9rvrzI++l7BPwgzXlkhg43F+c9amRba4WjR16QKudj/q5QeyxbikfzKmK9
lwiP6RS7Ja8B6Y6LEPPu1N7o2IPk2sbPcj6Nh3XwIM9wqPKaAm9bQeBMLbm/AmhbIkIDL9701Wp8
gxXpYgnscnRdK4d4xkf8M5PVNyxqQTDQlSLgs8zrg2sBA2jD99F+g2izwr9I2dIociB908j/O5mn
nYTJ006+lhP8gjHMh+SHZ0zi2iKIxV6/r7H2xKfnvCxt41u//HmIPikykuTpn63tXtvUvhe77dm0
S3xIFSxelHptwfYAI3CP8hFv6o2O94Hp/nP9rV6K15/DbUfXJQedI/A8ikr/5mPyMnTSH9973Xne
fztc9AcadRxAEhOkDHr5adVAohFy/R4OWotWlmb2FjRj7rEUIGg0T3dumk6HnzEtFpFoUbqhXtpI
dkdrBQ5NFjn27cM4XJKUiHo84JTdNM5MAg/Vm4LjVXz+Vn6YI/LhfqosRiFJ+XlTRnH03T6uFU+v
aBh5eQ5MDmby8BYvD8ha7FPlJVrb87Fnn1gA1yy3fjxoiHp8KooLwT6Bf8cX//XKUTbBxEwzw+Bw
o93gAQoHQ1WDbBLCrmcKkEqJYeHNbqsYFyoUVekBMT2DMn4T1RcafrWf+Z0FCFTKAI9eC4zfcsvc
QPfAsQFCLwsj550EhuTLPXTqaLgrXu8791RIjm0r6NK5HLvTeGCa6x48HtO4Gg1YKGkWAhNF5MLW
Syhfy0KW1szVDrUapOsF7gDDKofRgtaHFCrXmWKTDHtq0zMTREL20dw9RCHaCK16/IuqldlqGoLe
lOh8L8fNeGBldAT0/4XAl/zQLk9PkEjQ6+JAqUL2Z21BSq/DNFrACEAt8zFJXIsD03sajlNTilXe
tjJXsYNIPKnLAZrkDabko4FV5LtDJZvgw7ceZlHcTs1AHGPNHt4DkTqXXx9FQYwKqGEOoctcRVn5
bUndvtazeTtdIseFO12z+E9kEZfefanbV4BgXcbPpmHBvXC7VSKvNCYkP6WnpyCeaiy2UcR01HUn
Idnh7qiA5hWfygi46mO6lwIbyacUF333JN0FBK2PnXB7/dDpgdqkOjn8rxesrIbZfnz32FRIFEil
DEDnniqBcrjvYQvC1WUAf8OrmLbqq0lMUO8sEnPjJThxZzNTBushFD/WU/sQN0gjp0C8MVid7r6+
/YBeNs23sbfL2IfULMRviJN+Ga+J0Z1b17KkdUo95nnJxlXzLJuaaDVVsplYhDbOAdICGTvI1+0o
/19lsFhSQ6bieiwSWgOBMXplm2LvduiM1CQtfIoeXdS1Ex5kBVXa2GFfyjwPS/TVhO/ChirJyKMH
qebQAuboFVlwOfAf7Tpf4qTAVz0osY/+UwkPwVYqvrFND84a5fFdzhTmRvKJbm+JLVfQYtt/gWAz
DQL9uSECj/RLvIabTYC+obLQFK4xFF4R9HmX4CSiQ4tEIYxf52DPNifAYcGskfm1+iHKTuWzOC38
QTcDzJe3w50hDqL8VFxTdyRkm6x1EqX7a1p7i4E8m/TlKTbJIMBVs+Eza9HxT4dHtY9Hky+dEqiI
4BGNYaT+2j6nDbwgc0tA8Bu3JNGI2QO8Rp51T7z5TZ1oYqhGnqqUsjj1Mb0l678EvO8ZRHPqAlOn
fRfA0kxI1VERgi+1miY0k4hE6uJTEgkkTC7eZighQBhBdRsRamSrQ0iPnBa4y1RSAenrcmIlLqAs
rEFBngMcNPeL72W5h4dHj33ZBipWeCgPuK2HhBMuW69+vKZWwdRMPBH3EG7wYDJwITmt3eyJyztX
rGgdopDT+i/aDJ8QswLghxzXXKDTApuT3UXXk7SDYPPtSls9mPIiHVIPJlDmagCdFeNB7g79JJin
O3rsciu+oQmI8+KF+54XzWrG2qgtpk5BHEYw21q09z4OjaJRyh2ybP4woEaOiOC3H3FQsTRMkPb1
PQxKwkKpGyM9461GhW7B0zgoRYhHwZ7P9DXCF1tfYFNh5a7fQJ7Vr+CpLFTtNb+6xmvrn+7nbivS
Zj0vZsC8gDt4/JFWwHJOwTu9FaPCe4P8yHFYob1n8hdQV+hy4p/KFTrtSCR3KxR615w5y4vi6wME
Yql+aUUeXR6aOle1B+YBLMmJVmxFDWCfKxfpMItBJr+hcMZ3AK8g7a+ypOh76sMoPbH4CdWm9jVX
1oke+Y6SLBBDUk2yWey68qsFF1vN4KWSVin7dsuOe1Ne11WuUMGTES8e+Ya5Ic6uji0Ei1gFOnEk
AsJfs16Bk3g7nDsVpbSL2YIb39q2OCKAOmq/o+Elj5lVGO3I9YrXOSNJqICbwkSjnX14gIF2UfY1
FgB21fiwZQM+VDacR0tWmvTDPj3XCQzy5opGP4m/AR81YvSOkP8VJpWtXSYeGGwFtCBtAZpbirDV
NkaqzN5IEP26QfsRt5iBPTF3cLywTRqjCi9+YJURBt3YKw6k9K8mYAq/4SiiHh7MdmhjUZm1BewW
3+fMMv5yByXTucPzLIsOpvCoDmgjKla8V4shqMOs7LsHlfiayBGmWLCy55rU4vQZORICwFbf/Pdc
spKur+ijVL3HgMRydYgVw3oAO4zFkGGuj470b7k13ii4RhhrOW4MqKXPXmfvfqZi+V6RAWI/hGVJ
7hIsilkKWKug+53hfigfKd8v2N7m9d+i6ChMm473NfK4Zcuix/nzsCHiLC7sR6OQBGdnvvqfgaBx
PtvbebWNxIhl4WUr/rImIJrdXW9kfvCJKG5THRkzHYsp49MmDps/aHKuADC9HX5tqElFpjfjfZrj
Ay6kByMA8U8BxCEp2m36MfGlDVMP1m/gOsnu5pHBbrTI5x1Xx6J+966BmoPQYoVsBhESpCmzs3Mq
G/GWZroaFF0MajOch8bQr5Id0fehL94/mhn3I/JDwclqu/cPD7G+vzQO0a518G9gR9eiQXvwcVA+
1KzeJupnP14LLlWG6k+XN90pawH+S3aZ0LJE4ehQP0T8ZzQ6AmtClhv1rLQUbzMbHCDCZaDV2ztN
r5Pl8ZZMxJ3G+Xc4Vfd3kIkHW3RMXn3FFqiDFZJeFa5+qhQmz3WMYLUC7GxDQfIVwBgoeXQWjcxI
q5e6aQFhQQwS4VR8DX/Pyrywr3dp6vCTJsuUnYR7AkgVb06PHFfqrCpldoaT5GZuI5RTQMwGnyhk
m2u0hWtaZwQdC2C53D3nAglKYVQGkyCCnufkNzVfVtAxnRJVQBjqhjmLY5OKmNag1TRZ3o4E4K33
BtQkl69d+Nj8b5UXrPtQk0PO4owuZwjL8OGGhXkH18/eNbbMk1DRJnzW+x32Zsf77iAY5wUcOJWc
LqkeuYgcdhcgWmWPESxUsv/vFEVQLKPAr7xn+vV5VPFyXRMutbR6UZxcL+P1wI+OrKedFuodqmKc
DNXu8wXh8aQUBwItJD1nlaPT4wLGT9Yq2gvewAx3rU9kJrGUfDHubvhV23z+aQ7xiOJxuepqlEEt
fMz3F32IDO98HfDTPcXpdTzZOvNNJclBxL/KYOhAFMsFi+fkP9fR5c7E0qyR8eoRPSk2PIu+Cc5m
V9yYj7SrkV+FZrePBmqTN4Rf38aMft9Fd7aE1e8X3SSybI5mq9d9Mt3FjMq25UO04QGNLgDpMu/J
4rphdzrkkE3iwwH1cD2QsEdzBpogBdyLvrizlvS+vvzYy2RxZqQbZEOMAxVE/0R2BenMfkn6G3Hi
+PaY06HmnmaV9WhnrmjKNxdEzwWIxS1Yih78WAGTuUkE4BKkMrNcKjvGHLJHGwRv7N3PckR9JHkU
BUepwX4rj41RlLWBbW5ggfHSCVNmdXjlG+WFWSJ1fDZ2uqYSvgfzeKHFWhi9jRDIr1BppLuj8jpN
W0MCg7q8tCBqln5hSnr9oYsJtQR6JsZUcWYvFtQ2jFDVeIavC4psibdm3pxiPdOZOGZo3lyt68cR
uzre+49R8WOT0oJSs8pLg5qKQfDlfsDmsFmIPaGeF2A2OTJ/rumr2JjaOZSGXHYrcEUYMDnJf83j
SdTndfYf8jvX8LZH7lq+ekNareruqLGVqFpR5OHfx0lBEGkU3St6R4nVuTD6KeL5GU8qyqbHdbTj
ok19nYEQmGfLMO2pR8YopqeOvVQfQ5piO/dYcZNcIl7pYeODmMJ21AV01fGkD+w4tnAQCsm13OoS
Sgc4g+vZhpXWklVABKSnL1xUP9mRgFupZ7uE0fKkdcSgKh2yzkqxX/BMCVf3I6aDSz0k92+W8/lK
g+hE0ZH3KAU+LtCywsuqQd5HC6+vgR5cXR+L1CJGdvVnqT2qQccMk7F90pWhjHDxLtw2GzRSWEfs
2WVWs7j7EiW8pbXr30cPDrLyUL6WFeDIV2H9SCvitPuOgXGAlmzArpDxqOiJcGpo6rZUf0eClGoJ
y1uX4SvnFxEBUMrTeYCWrL0JmkJWuYUT3AcbiYId3D1rsy0V8zZQm5fzNq+E7kNY2gM6jPMbU0ny
PVtdaSCXUXYLiDSRJGjC/hyAUkt7kAHb/4Oi6qWS6+/nPaKXBKjI5xFLoTHPM1Z7hLNiHqOHKu0X
1IHPcbUn5dJBEsPL10UtVux40GTnxeuCXppiB/OQVJj7kyVIaBDdoAC6oYi+/yg9Lkz7x/D/hejR
E96wyPwc5LnrREIhWc4oBicJXhUfJEOybbvSQVUfoT/HzaTsbCXWF5Vz06vDTKQzmhoDqKLIXEkh
GiFvkCaYQ5gt51zFMARxmjGzzO5Hzb2Tx1pUK7MUIk0FYHrGtUkbnflC9NAOFUefpLe4sFQpmlYQ
8MRxILrvF+HXQWMh9LQmLONQIlzTyQ3+FphRT0PToEw6xS/f/pm2UJfXqpyT5w+QamW/WvgX5SLy
H2Sor6smeNR5r0bpgxaRJ134UNBGUcv7zCLX0X9Udw8K0vFnVTJRdyvwhftufSxfyaCfMlgiw8ik
SrsUveGXPF7sH4k1JTJYo4T4kgO6Zf39ApeFERY2VQYgdRMSSvZEyH2oLhppjehYjYLd4Nx1XRed
VCsFUiLYbNSAn9crJkGMFg8m5+JUW3ihewMI4ZyZGxSICqC41dcPIouLmLpoz8CaUpNLFAy465MY
4Lrr4sZNvaPbq8zWm++PmYUdokyi2NJuaQPljAywn1uwDYeEgrXbky6FdbuSvCzWnTZaoeBNxhYg
guQsl8+W7DYYjH2b1aIMSvGQb3W5aXz7JHAw9SRz4y849l2Vn0eN4q/2v5WQd4zIIleTEMjCfoKr
G2+ghNw14gcSKh8dJktC/jt7JPYd0Fm8ohnneaccfNWPf7ssQ74HvP+5CwD9T7WAAJOlVjMWNgL7
qC2J/8UuEStZ5P4YTd1GHIUOIIDOx2lAdLouYg0tcQJYqc2IcnNXnXTFdQq7s5KStqN22S5+YQEq
Eczdq5ep2Ko1WE+I/+KQFZnVB4NpovNPg7YerxYIXv5zIabvUMdd7trYkU0sWRA8BbBl8yfxYIed
TnL3jWia4bs+qzkWC+Y6wDFlGhIINBVB7Y/YL/dWN/k5cmje34YeCpfVpHj/CpmR5jhYjvUsafvs
NP2kI60B6kj7zoeB3gNjbp+bK2Sp7bMOmE7OxlKSpfyUEk5RJ5p9eAcH5xBzHXQiXoDhnqx7sm7+
LZw+E/dUQdFmDjqE9W3nkyXE6N8QWzwTRhbtGptZISvb75OpjCaTNtIUg60Cn467fLjDzx6W8/h1
/W6jucEWu8g50iC5VJhZvKFsIgH/ltk24XquJXHXVkEC4IV9xo0r1mhWwyaO9xET8+u+5wbBPUBA
j62RIu3ZJUUpPYkTFg4LO61gB16v7sifvGJhXVKQ4BIYz2QxIBmie31/5dpt3rjFP/heM4jAg+Ev
lzS/QHwavZsifDw9Jp4pm9aDpnRSZ1/7qH9bKeoMDPsmvYTDrHZg2BzgX4qvoz6opw7k13Jgys2g
Dl3PeCYckj1bzaVpa5zq5+uW5k0x+Juho7jEzBGI4oJBLSz12h8P631ToAuMc18TeIHg7ai01PMS
WwoC+qv+3L1S3D0hKDZPvlG6fi0ng4icq0CJgV3/iL6eGfbOaDb3+V/fPNrKbvHo1xAb7xYO3VSn
IqJjsL6EJ29HYm+DpreyytLetC9R+bhnHqrqD68akgkxi4bheA2kd8Nr3Qf24kyGtBhw6UEYW7s1
Qigj2m1fe1mnC3mkIQNkInV6ppbcsj+EnFFeeW3XIhvVe+2KoA/l+nLn5d9RulNsSH0L9XHUSeBV
cR8ABAU5Vczf0rFKlv1FOhPU068SW4pK8rZ3l0x0W56wPLS2D0J2jPqMBVAuYqfnXV6wyuAaf27D
Xni/94M/VE9pLOAgV+JeI/tISTykNMamSoGp9k5mlmqN2LUQqyC/2ytt0ehcdGkaCxd1Csz3Rglf
8yS46vwq7SL98BO26pPm0OY3PcNAWvPdwywSS7h+Qh0XD6gzSoGi40HWeJyvpuhtvwedO+G/YsXP
+9ps/iOvtfzoOSNwQ1g5FVAoaBLOoVnJy+/hF68tk02mUamblog6KCbI3nAu7VMdc4ULVm2wWcrl
gz7Qu8f2hjux3f3ndxzF91/iPqa56uOKAxIlvX6D8im+wIce7ope0F3c5XU0lCE4xAv3dNLtUip7
UP3Svx2epYK8NWwbzPijuLBdFBw//SkZ4780RcbFLsCb29z2nTTbau1Al7RciDi1SuCKo6ABwu59
VoNxBuFtTk16DGYF1XkH+TpFF8JF3lGqSE/vgCDYpmm3W7eyC7pfiSYO1bXxtY83OiXpRTEbmiIT
sfwqPeV/pqK3VNX7ST7zbPCFzRQw5cbJYjalG7Lh/O+5sVZfabqWES0HTiMK3/ATLU7685BC1Agq
JzaYr9ujSYK8BNyuYCffa1BhT5n3DZcDlKbY0ojG6RiRPaRdyvf9L5NTh88ett3pUUaWMh++EqNl
Z3hHNNAlmQW+oEvB2wlxvfVBNL9VJbnuwuS4S2/OqkeDFvWrq1q7xW8BM5aR1/NuJuonAASFnRQd
GAFGcDoOqWCi0eG3TFauSQRdvuWIb07+jWIbtNG25uwx94YovZICSD5H9k8zG+4rKCWWdyauu8lh
TsFFf5jXDuzQBhynb7Km2dj5ovxE19BhV5uO1wjJ2ruNrVr+ZizeDB1b6vNoIUjMGDQQNsm33ylq
Phj4kMa7dMyeA7L9Op1MXPQgbSa/6FhAQhsLWFQbaXcgTybciTSY4wiZNV1Y575KbHM2d9lWgHSz
EjKCL4q16BxgxifAxoXF0g+r5l9EWrd8P5eGhBEE+9AnhQOGKkdgWvctp77/xufg+W3THEFSc/JY
DT3SgMOwHHuMQpKCBACiQ0NuJHmYy7lgP0V4228umZuSHTJ1BEItVL3itxr8VCd8g8hZ51Wvwp1V
gOIErX2tJENP+CyaU+wFDl9rmOykXMOGnpuwJ1gBetXlQQ1j91tsNtc7PljQK1+z5HWVfLt9eHB4
0IbUDu1kzOfESN1gH5D/rEyZnhJ41ZE8BJBuPwTAyDkq5g18E3ZJNXxxdJx5wIpoTIa4h333Rhgo
ez3O1RSHZW1+fA0kGZ7SebDSiSNpZDk80UzktdHvqIwT1W0YyZpIk8aUuo8SYj3abHCyjx5GYFA8
2Nk3+zCRtpGdQgDEvaKC2ZhbtvGjF65sYe7eT9z8zjqVhNjcYXf5xv+djYCbYr3+UQS279Hjo6Zm
EfDPTO1nMqsh2jbX+W6Awmx8N+SONAq1oj0VOd0+0c/xVnekNBxdZ/lRFCTvkFIX4Kc1DiHHAdac
xIP9NADkDdiyXLo1iwmoKOL7UQ9cwBOvP2leus8VfJSO84cdkbEAQWhomwqoljQF9SUQ1Mr3uatJ
uVc/fxpZhtJmr6F6wp2xXPg2PrUoWLIf+Kfl86vOsDvlcTqJnrGLn1PgDJADGK/iEs4xEuoDQ/Lr
7JvTiJdbLTxPNeEqyUkaqG57XFl1/teGPEtPYfD55OZPyyrthhedTX13JaO2gl0nAkkrHX0QgBsB
8Rl+2pBMntdLNIxB2n976s8SfPmStpy0OqybTb2CknAZw90PlpP5sMuMBCr9Cu7Tkzq3CZANH+Se
7zsr9zZObls5yLJ2yxDhN2D7Sh/F4mrmThmOxE/FT2cLc2b839vOxOsTZV5a7Jq1IkhpHXk/gvoY
8MkTpgoPYLlPHtMubrTSFSn6jMzcZytesth9wzYBormiU7AhO5NSxyD0SXJjNjf4DByvHHZ0ViXt
5Aub9X6lMwauKc5wGe3SyDojV0/6cirBy8TXlZ5ND00Wp594w1Xan/2ndQfJat6NIOjZBtnOfAv1
UuRRRTTRWrjPOrKZ4HYKZimeBgzd6TxcpYEAfyLlNF9TeAi93TUe9lmUwFsqkOf2MmhLPePQnocw
ztr7dSqggay8FN/l1uFhmMZ268d1sbxZqaVKB9UzM2TXu5c1uwBGKgZ0Qz6fUGOAo1AMZnMzxGPg
d0fLD1F0AlRYgqL3OVBwyzvZau+j7z8WINi+BoBaIMRMb+tHuT0lkeMvMTC/qY7pjaMQZ/Jo8PDU
KNACuKIB4759FQFBu44A79pdcYKqtwDxJzRYPtf5yORw2XTr0/oLEEaogx50YU5SxysKwfCftvhC
F8ZoeNcu+0IphPBNMqfLsRb2d13nKcsPARhAaDPTJkQVlXDplDuq0XrrjSM9i5/3Q8u3x0uKHulm
wq3Qgml5s1I6lupHQT1omdDcxQ/6bbmklXdBY0Gym9+9ThrrDVJf9lijIZRikxLNGr/Zza6p1KeF
uTJVu2BVwaYHmgpDkdYT24yNyGaHjcqtpkEEqHgeGsyFDQ5Dzt0z7WV1HUs5zAZI1pBpkWXko9Jq
Gvn13u+ghmJZP2YvLKQ+FdbGzquvOwaYwNMhaLw98gHb39DLkgN1HqcXFWZ/8edn4F+k9xiLhep6
I7b2Zgiwo7KVUdBjFz1FJW5qpvifCd6DcBDCDZ9ytcAa5SZ+gJnwxz2e3Yo3XX9p2isj5VyT0zn+
DvPLK3JjXFURAiNwhhoyk5kRrWItWfaM/x+wqZga1fFeABE86XxxPoajWTJqF3Otjq3hwXxST1Pi
N9jlyrVH3xbYRMGS2MsU7I1Gda/WT6q462aMGwXKCqPckqDtbj5Tg81eW3CT0yeYNby+dzX0Oapb
897vSdml0GyNCQtsjs4XIVeT/lPa+vMLQ+qnvL7S4Kw+M03DX2dvFNXH1tIwOq9MHEVkneLpPXVv
eonTyQI7Cw5gGyQJHJoT+v8w7QyP4kMsvJqU2kHIP5GhmB4zzXUwRBUV6kLMwJN8YyGetCqrxwHG
20Q5Npx6RG1dKXXtlswFkymVKd817QStKfWm4SfKTL9RGxZo9z5gc2piR5ScFc3Ck9cp0CZiUuYR
TIUhZdBkkDJbFrAqEJOhBEff/Ez9xzJs8n/2YvlV8OPT3PPafQ2ti3Gr5ImxS9kald94WtzS0zQ+
tqz8mS7HNMM59ESwdq+I+D0U7elWsRhh9Gu9Fe0DAAecAScqDiyZ4AkbNWNnJil1lA3AtWrazdXa
9tdWvAAU3hjDSyDMVhg80lLPeJCzh+E42Llv6wECVS0rFj/wddbFoVLj8HIpFMJ8HWYNChZ5GV7m
UtaRzePQ4Q4A9OtN6xuna1COq2321J4/nVaEqnyLa7Ek6qmhSju62vtNmWF9WLwjCrsnrcMM4Ysq
xRIFBaALQvTAwzoY+CA3pzIS/k/LzWsdogyN08hCpnyKAQ1epI40pur1padOpCOVv8vFUbXCiVQl
/d34XHOXMeSlMChv3COipg7KGfVJDH18WERr/Nu8cygLbIYwpfIfzOhGmi5o4xC4OGQA4tB4ytt0
lBnASlmSuKSbkge9kQ9xSKzq2Ar1JsrVJCUcXuueZOLdtTyL0W4er07cnkTL9DNjtZGrOHLfCcOl
YiDwx0bGAI6IpYMBo3vyyU2/BXydfQW41nZs4CgQxe3GUyLyW39xlrAbHi03lgIFTSM4ZWuRxi9t
++WImZd4jM8WbM91S8TQ7akWAP3EhJeZVlz6Cu4/ksmwqy+sG7x5Z6//2QT2xFlY2Ivo1BTjwwI0
x47mQtFxZmbPnUrKc0MKWW7Xb+uniLT+rmPfksv6J4QUsPssc9DrONBtJe6qYkdfl2USP+hV+es0
Ti2uC8wVJfl2A9GYy+iHGay1KumKHEbYMI5WHno2p+TYgTaFlZFZou9TgS3yuDu9B2ed5Ax4i03l
ZK7Ri33qcsCxaZqnWIPtBtrMF6SFY3jqledqbYHu9+7lV0nOZXLtRVhCqD1ZjlcZZ7SF+kDeu70p
9c1HY9kvPfL+6rDxfv2tDOhD7RINMvydSeI6VhccfuXBSO/u8gcv3c9h7e8dEwrThHKuDjVBgEZu
rRdx3OWGS8vBltcSnnK8yZBq6pZ+xFa3u6yzn83xmXGykiZkDy+c7NGx3rXpkOGi+vfSWn/owsZm
dz3/QAqvacgKkvf2m/BdEPVsoaCMliSx9VKz0tSYdFgMyekxQ5vtr7jcMSmi5GoHUjk/9tIasPse
N/psVYVGhTBT9aCcbxff/tbaqEBNbAd9OXGeYXtEKSlVcVft0z6dvAEUnbcP7BvLR8LUJMMxe4tu
daOPKgjyTuT1tlHUn+oh31A037sYefSmv3GmimM5DIXrKg8TxP2D5XD7Qb8j58X3mpiUu+sg+rtN
ZY1AGGaI1ufA/uod0bvdVdrPoaE8lbVykQaiF8giBgPQHNRzOeHixsYUYcfGW5x5kLYaDjejaugh
Of5Tpyz8kFq7Uox/rCsa3SoT62zNtlrRfPrV34bwGivRLRoXG++ALVE/C1h2c6yPaUOWjJPCZHzW
Mor3mr3gWnqR92e6bDqHURedCJEaBvptX3N0YF4La+u4OU/Z9u+E8eU9wpRyixzDw4c27QmF9HQE
lquHDxfh5v/b5w6OubgIV4lVCM9oZZOyDuSiXWQqMaR7Hx/HBM+OdmX+UxNZYf39rHAHMmbtiOIr
ISGcLfORgu0jZCpAgxzLsP8EwMndid52y0EMqxoRDBbPz1uu7XWywGgCQwak6wsb9tBvq9zNYe9U
8ONkfrUVANUffQL6LTekamki0n5PyCLzkTgEWspCTF43mbYVDdunYQ49lVu+WrFYJbB5DKZjytd3
7irsV9cch6fJuF/TSGLey6KWJ3Af3Q3OgK/LjVrrBoMu013qJgw65r41QYuVvlbE0mQfgk1S2uIC
kOL8XI/47MvNh8LJAnXYUxTsoS5X6MPz3xZa2G368DkWR9LHVnHfXVKLHYerUtfay8vJJIOc6yt1
PR+CQBU020s+adJRga7JO1IRPPfLJPFAOpM78IC/DxmkdePAdQBrVAbBASkiuse4clENtRVmw4Fr
p/e6ZYhiqJAeVwZjpuZOV/eGM/eI42aSBiV671stjC/h8HAhdPIApJwDyz2HC4QEA33LBXTKL1dA
vMbarDZE/7N0OMSQPW5G7s0g12CHXO/R/3q+W7vgLtmTO/UMAFX7OmEV8cDG4N/BYtrzb6QUiNy0
IpzHJrENmvklbbYfmhoG/HemRWqC1n+2nBwp7ZYGYYjXMUrXQE+RuU0QG/gMr9vPPdDz0EVGPxjc
HfcMkBBeM02sKFq9IJkCa/jc2wI+2Bn2E9mKGnsQMu6z7qLfCehILZ1kxaRQ48GSHa3IQzc3Md07
2o04iG/+MU3ArRyBDdJFccApjFC3LHSEeWQjJomd1oueCAD8A+F56FBa8zgsB3GyOgyQJZoeW+6V
p63MdEE1c5gdCsx6QmFPkWg/un85HelK3rVfJ96Pg4SCj6wZYlTblviXcC9EjyOrhP3SyEGgQS+B
UQc7UdOTfn4hjWFBCkE+7dSxUZPc13F30KZioc9APvCpsjR1mN+13wNESksZTWqpoLFKeVK7XGa0
RstcmTwYA56CUoHP3FUHxmud/Rcl2AbN3GxlMpZIUeceQ1QCb5Si+fDmNvFItIl45nxJAnE05rXo
CiSpzUzjGgCX2Y3BVeIrtRkjVBFXUjrJEQ5LAr9ZYX31qZYKBdrWu41QxUQ0JDZVVDXiaS/9k0sq
fbzzngK6pZTIE2C3d1IzjQD/XzqQUpSnyVO8XCb0VQl/W3hyDSwQL5BhpZSjJA9aWAPTxUIjFC/q
6fAlPAO0GPslTNBK1z/ll5SI4QC+PIzHVWTjRaVDoA9mHqbbVg6NFk8m8dGFifMCrCOnCqo7jg/9
MzUbRTGqqAHh9ieSBeK5kXnHv2Pxd5SxHIDRc4kGy/FmXq38zjndC4Bd3j6qCNinnqDhu48rROBG
8pWxYYeKW/h/byoFLmTqEXLpXUJ6Bd27E1S4k1BvHHyVd5uD6uNVfq0jaZS4aSPFWHpuN0thwhbX
tFfZPdoz9rTzSMaTOUw30fZC2IpxPDjYPx2gVGWJz7HXP+aSbkDWax0k1ZqGU4tIDxpaeyII9v+U
xAonqkBptPAybyv0V+UgAesRVBxAKUp5MW5vKjLJfozU2QrZ/rdVXZ1XNTSH+ho4he+U4wwti1kq
HxECCqwO3Eiuk/ESrUMwHavtOndmBXWZe+J66UbA4bWdAACapLX9QBxyY10fKdbTKRSexaxkFYph
hmjzKz1ivklQi/7Zh84a/STqtbbWnMb62+RRj6nJ3qoy5CJGRpB2q/TWq7qQUqXzaPs85IQIjZVn
ofVkypL5kfgcOEm7tZ/LO82zfD/b56L+nunX1fGTAdMm/8nBftfnag9hJB9UQ2PZJbLDhq0SGBqz
DvwqfDWq80bwQi1DzDK026wPJxxJPGyvegF8sjeP6u5evZo/f2jqF8ZGY3DsGIiIbhIl90dHUxVY
TU6AFuJQnbgjn73fiA0RL/jLbH2vIEKpWJJrPNdJpoVjgIqit9GGrnNwSjfc9AMf5QkKmANPxqCC
ANjr1OPP8Z+ak6RCqhmTBOGwW1510fopwIABmGGElqfi7wn/kWqlONpS/9f/rz07mCZ8fL26Lxhy
1LJfoa3hwVnP16Z5YIjCMbOz+rNFY7zF5vfY7D3YqSsASc7I0DrIlkeWIOsIQK12m0uwGddA4hQR
UtmQnbbPTStQoixPxudirE9p0DuvuOFIjLwRw1Ke11TBxNXu1blnnkwVLYHbkLdcbbIplLDzfM1H
LJhIfhA28rovXjaLOpYmgk4En/dTUCD/azN9UuPB/nHRnf3gu3E58f0xEcd6XNiyQqKQ5EdkgyMW
eHyKV6vt5hoRsRw5AwJxErTAPxSk/dhf88mjkUCq0Fq6hZyXL1DTw9/DxBAs0tR0dudxC0/s0CKm
kbzejTQ+P4rkv9GH79WIcL3Jm1E5D/jRIgn1aVx4TrAUDqUvaKcfkhx8lLtSgyxezURSAGmlyPhq
pYm+X9ZwSzVDMkzbn1bttOJOFNG9trHZ2KJUaAFaZRTeYBg7n5+kv7GBnceDjCyaNFQgFlPUVmWo
ualiEQu4w4wwZrhnu3GJ/RUq6X9CqeecwyvjjC6FCVvNXO8c5obctQbbPX01lo51AcPLd6oqAz5n
H7VaBVFHmgtygzTjHXERfV8ZxW6qge7ri8jfGOth0pFnst9BdzpLX/CbbKLx7FEek5bOcD2Z7TY+
ffTHiTd6ktVU2Y9L6rX/nx9PFetzo5bV8E5eFEvA3E7Ghrsd6nf6TnCNFiHCA8uVAyyFDlksj8g+
bSCpWtqu8QISKnBRtV6OcOjRfEY4NbkU6A40ZEL96DUxI4CfgNWDVLjCmFpPvq0x4y82cF4bw/7F
M02oGXJbVDYnj4WFlQkWDmWZHzNXMpFI4RUuBvP0kgySzitNUEsy/ygxBICPfdiPtJXyu/dbaGm4
sWXUoJg4FUhMh8Q0eqF1kFUG6LS3Rq+qKZjpVF/RpI1+ceCitCdlgx8xNUDca9zLaxoXvkdDQw68
0AE8D5YbYSDjkxT0WYmupVl3zJdGRgIPFPsbRYMuW+jOQSQOMfkoAFMjy5iTQwdJQH2GaD8iZT5G
K5+Odtlp5+JdhjCDGqZylOpdOefzuEkIv1LMnSW8WfyKXto7YEVYRmoGaJ19g3ZkX1Ug+kPfCK5i
KUDrYXZcO59v5zmSHwUXKHtjmEVHjWjs8a5K4bzvOYxedr1VyXKbmG6JZEHL7FUpKlRI1OxEE5iD
YyqcyVI+3HNWjYgY8/wqWNA4thp5L0H/jikv1MwGZZsYuGtRKqlfSSqgypteUYxysyjiLu20cekG
EjAdDrjt0YKduc4POt89SwPNwfDyB6V6TKAGNgvofxc76AnHXItKWiZVEgZUeX67PlbBlSyQ3+VG
udev/+I3DNnEYIo71o/w74jENtKPKqbieA0yAtjsaSgI/1/kC6H7rGkOXfr6DwTEZfhAh/IVJfE1
P998ePQoc/6XwrtLCkrY0ZyL3YQj9urbxFZyXpnGbN11U4AnzG/pOGT70PVnxiNk7IsFEcCOfRRU
o4zYO30cCJMKWJ9B8x8N8is4LQKVAXvpfmIi0jjjMQJfIfSB6O+iB8fdKITqAdloaQGCU5HytuIm
/lx0u5dl40CuFOGxgRuyN6+Kj1ycCHcOy80B7FTgZENJysCqoQTWFMBgGGakgpBHGF9D832JJr8q
t9o4GXwPxNOMulkVNoDiUaCc5aSyhFV5sg4OX3663IOHK26H9dKIPWiWJyull4/7NNt5WDRsr/nJ
emVr+bibInv//qAM77uqwH5d6o7zNsOwRJVKa+KlBnQZj6tf4T68nv/94c1erjio+3npxFQPIcuo
1z+5qNdeOu0RrIZGe2UqEilF4lHDzO+2bPt5U02Ecr4ov3eY9bvvp9TtCPecg0igKqeQ0F3LqK4A
nYOXUxjX2D9/8InkD7VDcvdGRIf4XYAZoYui7QAgI96HhL/3BKuLpKsXAztz8UzjhQnJH9n1LdXh
JVIxJfUNDbjctDX3SbzkkmGnycTpQSDz+QDj+NPtxqwNEFuN0SqYIi8g4U8otMQyZ2VRwwdP1Wc1
YZSs3V7BcCGUhuXssrhvsZpqZv6ibskjv4gcMtBlckuvqszaceHqUt22HZ6OOp8eL0SVJpCvhQcn
JnwbQjWDbIvBk67VvJI03VIIOL3R8ukN7mQwfj9rWMMXdEIECnFHKMLMhE7l+U0hc1J7oynsQaov
m3OwxFi0LBHXa+ssCAWEuODFobkk6hhdvsovnkQvMFmjfMJZfdifTQSNom9wB+6NLykCrj4+Ubgc
KjjLKwSg/wqXZXzopgbDIA25cgZd2frYmYkVZG+RgctWR3hsgxr0JTz/zkwb6hegufIXK430ZfUM
iTFx0wwk8wLJ4ZjPLNtdYysYIo0KCFONWtw9nx+1OQQKsedqmDuPwogErt3wLY3HUQRmMn85ibXL
0G13IWVTiSL+WHj8RlVJ5SFiHmkc5wnEIzOtm7vhCZCoZ99vTgHJNVivvt6V7zSfLk9jasS5WUtr
8ITr2q0UdHqgmDZ25G7w075BkBluxt5dbTEHZr16jLng1qbPJ298lZ/wLV70B87ETmA83rWBgg1L
dYxJbAC06+k5R8jGefk9gjhJHHR0OxE3O0/GfAEjlHUHFHryxqZ6ZEhwb3gNcmU9+AfZBPRLKT7T
m4TPPVmuNxxFfuEhNx3N4w8cJFBx8bSwWpNb1+a7z2eIT7LujLEth9/XyO0ux3iFKhI1WZ+Caluw
aIxiGW3IslEi5vkIUHZ4ZRKh7wkXID9ixmWZ0pZueVZ+zstZsl0ivssR1pk4NJbvtukDcu1pOI+v
b4NUXnnRUDuG6KKxGwGwH59nFzAjutkWczga3K/pDs8sYpohw7v6AAFAvZVHRtpVrsg0EwWpgtsS
BEtmtZxW0BzA5a/NpATZVSi7PC1atsB6vOi9J/PIgbUyk09KMkp5nrmJyfgyaKU8ye+Op+eJQ6hL
sMkyVIY2XzvRYvw0Qje/5mhaseersCrHQuUF0fizYx4IPCBNxmTE+NuriZH1cXZwXyneXI7iyaKp
DvlpR7JBhlYnn2XBBC7LAn75fywg9aiTrbF3IX59cY9+ZlGj2Qysg+FzPqa8ykMglphprzKVLjRJ
JbUSnmgEIAivoqQUHvTVf1UI5zaYL7JSaCj+Un6q+X+Asj/4bSxDTXynqM4obqjdFJ5tfth+BvgA
WzK0yAlbNsulwusKHt2GhIyn+aN6/VAkddhkf71rGcAP2n3G7rMSs7LrbrGeZx2U4wxWoNhG+/wE
kXrVvFud7gtxPWlAauPXEzREE+4eZPm2VgYWLlq1A6kXnpNr9mGsiZeqWGpZOnvSdckgXKR/6aBQ
hDdzZ2Ok6baG/5vHNdpEZBeVkGlnN1kOQnKa3cAI0pk0BHbl7QbIXYgrTqquzDRfB5BebxaIsk5K
rYxt5621MDiBJ5sruFknlf+uZIfYl1io5oOs+/WxKDbHtrjtYBP0hu2Yz1oLZyHT+gIdG1ABAukN
djtlgQoY+U0ib2y+MvuOvMb8fzp9A+bm4Bhmp3BckauVxVd/5O6vjmBbtb7U1Z9Y+OffRWNFPbpx
rOYaqtc6mJQ1PpFUE/gLBPR87PJwApHC1eXDOjzieNOveG8C0daFO7P6zHJHzrE7Bq5JSF2RwQvv
Xq2MSDJgrjqOOoaxunlUCczQLQsxOxaR+5sORoDAmCleUZpxUJ8+7deYcIzfsEyqIBxgst+UXbss
ctfuiBZNNKZSVDieGKJCTFtkaoV8duWKx5CKDGIC51l76bvhSP7M1aFGWYkkFJavXVjYF5iQYWNI
T+W/ip1WofXt6JAoeCuLs3Hg5MTMOogUln0e1Xi4cJxOElU42Q1Yuh+HW1VrNUE/9Rk7zwwRF9Ib
8O0+8sUhpgERISStQxGbtKbmEzCODk4ZBaj2KLRLeWTUmQm6n0CTFpjSCf/0WmNUK9Nxa2084huX
zrsRe70VcWjRMxuOusyQ+fN+5IPdKJbpW6HE5UabVBGou9+P6j7M7T6OB5HrdGkV7Pa7NF56lI66
+H6XVZeQCiELJgwuXgZoT3rI3EplXSHpr/FZ8kvaod5Bv+47tj9GPWuYXFBn7HkWDbZeKR4TRebe
OGal131F8/FklTJzcKX0mz2sxVm0tnW21t3gv2wSKsMQjEIgr4I/yc6thzb3DtK/FvHxUUPryYJd
+w6z9HEn7r+XKra6D/TgdqqElQL6KnzNCMCa1gWDkLD8LJGWrYR3QZd+DLJNoByju3TzmRIvyweM
BJmobAgzNaEaZgnVJkhbznCk/OiNXQntUM2NvdOXRIHN/0l1mG3G9GfVBpDCKkmi1/WdgRZuzqad
mF318alToYEM8C7mdkLJyccYGAVo6Ysf19NkFkD17hPjCbi7pLSIDieNwDlGUoVDOUNFm0OugDoi
5OIYID3FeulwqZfvAylCXdcRvcltF/cc7fCOjfer+KvVjpgSYx+TnwteX+ksLyohifuywYzUlvYP
hzXr1aJR5QIioig6+G3nJteS75H1XQ4L9RiaeBvZHObDeQPG6ER1DWdbHzTFkVW7H76ZUxsDr7fB
XaJtXwQsWWoADHvx305eGAJpMd42Jt7IRByBgUwslMBvzJr5srv+coQWtEkbLNriU694hRODUSIV
BrIVBQQtLPVadA+Qdt4VZaJwLMNrOPvCeiz1hZE2rp8H5BAGUQWKZkp/3PZjRWC5kSd+umxDVPtP
pULEGDKtJK9fUiTlM9N0+IbRe5IomO+Jp/fcdj3CoI2ulGjqBxZRlGS0G6npB+aVOGnyJnCpvHQH
B18SADyK1t55tpKopkCnAieXrewdoQPYP/p1uRIiTDUZZfKF6Enhl19wqjpWV/1/pYGPpx+a5Aun
QM6hT3kWNii6O5UQQdtS+XuQN6qxk4FvWv0XLmA6uFXvoZD4LT6n/rJ7UBrew7NOnN5qzCyiqOEo
vWFAtjfjgwSVTkQfDbgpI113PbfasFxJn6au8KuRH3On8gwwrQZYbnIyLXZCjIvOP1Ox/UbCEs/9
nIJ2Kao8fIzl0RZV7gwQpCYxFJUOrfmgwD/Up6xDXuf1myJWuKPhjnA7FzVSphylTiGawjFvqEZ/
nhchJJUZskqkvWTJcDxOX63tjv7oZkBXvh64RHpZixxCMtsn9oQLItVEHA4SaC3xQw23lwEOMLDd
lBX+58TP4dsct5LMLJU7Fnbvh/WhnFdna2tI/pLXRUpfMJZmFFS61yJn8UyFmnNsMFnYyPYVTLd/
OGfljcXMtyp2axp2fSdpMKwN4pV2C5O9Lj3G8M8gd8o7seGnhA8XYyw/N3wSHPcrrnB/pKDgXwnm
yjB70cduMF1fNV+42VSMN4BWrPwBeiFyVn6feLzn/xIXfjNyE6SnDj7AG1P+35VNcweAdGq6z4ZY
fmGJUMPnuBfMreMh6xuuUjVCuF2itoeNAS+veh7SyEfGipzDeftagBwTJ9CcX2Kv5PW3KbF3lovF
CR6BHpiOyPsFSDCBN07ggP0xNif5x4yu4mCh1ibUYWZaINkxnGpa5L+s5CkiPZfbJHXjTkvMJA0f
VNGsxrs2sxeRAfjFX+2g9r8q49ZdhpsJfM131Td/toZbLKar2PddRXdWzZZPIER0rUVESunM0WJ8
Ctq2xgctlaTwiiTfSEG82pw3a1IopyTIIR1sB8hO+8ewQx86FWUDN+HUFxis8z9CA2KCRqmnpkiA
eme1isUss/d8gfYGZ6QGjDMS1i5GKtM5tojCZgKw6FCOPNmiXf6pirZ/Lq3KKrx1O8Ny61oc5ljX
rdFhvZOo+EBM/gDlwHcmztwaThyr/IBPTI9QtyDWmUJNLQOp0TgDonGs3nz8zWpUpqHm17T4mcfO
1grKoUw+JVXRmp8uUoxhZAbBi3zxcr0F4AeWIk6PpsXxV0ChN5m7Xlg6zm69+9XQZbH9ZK51V0yM
j3S4bjBQG1V9dQb6Q1Rj5IuSr24MSiMGZ3VVEzcjlr22gusGk3Y3xp1KisA59+aVnb//j2SnJzpq
OMUb47F0sDL+V+getrxnrxj4SdSJgle8MpH7RSwL03Y9RpBxvBJiYo4lmiBTaKt/xPITs6X8hRq8
Bx9y+2x9tFVaj5L7ni9iYvc33KaUk8r8x13OGr2NMG9QHvsWxyY8dLT0dBzfd3sQCR70Qe0+qzyg
PSFGyRFw4nTs7r3RUmhvjA6OwWd9QtipJAbkLfGT5WpesZiaOsWuiQCIsW99+YealvH35HALxkXS
2I2ci0itiJV5WJqc/yQU0ovfW7c3DgrhJbkL1XCkt759WfdZKiOPR13Eua8NFVd7UdwS+R9S7CbJ
D9V+D04u0ZBXUxRW1R01Ukdpywf/Lo47h5AwThn2VTRaBaQBafKn+qJEFr26PuP7ySlVhKo8vOAM
pqfOlZdbOO5aC5v2hqWQ71Rxc4NyzOO41dlXPUB5UtAYTOURaswlROQyU30gEk68jgoz+sityyMR
N8i2o8/0ESvkfsU0m3Q9ruTyvCofTyPJ+uZLtXWaHZxNmVYOhQlqsRX7gxHqUZvy226C/4C92EPe
frWz+xSewp+0Y4SCSHKnjxJ8wlHlIyx/M1H7y395VJQkx5uLB9wsN0Yuuob6v3GGk209WBzGe08U
DFBEh2695M6OeE8eo1QNTufnr03qMPFQ+aeZ21m5V9VAZGc+/FtzSMf4QuWPnSpS0H0MymDz6vG3
52X0LedLJ5nPr1oGdX3m4D8bny9pB0CL20XTEKK8IaMgWgVV0lS+KOBzH/XRaa5Fo1F0rcHtWjDp
9kUS4AKp2klZdaFKKEuIL1tZ40PnAxNo5Ij0RXJKetjZ0thRf/BF6xS/1YV90lcc6KC+CbzcE9Gv
wGhGTy/iOfpNgijxO9MEUnqEW71fGWKhlfiOuKLaJ/+YJgnLqlczH7MWlFyO2WdaD1dyWEdBK0Sm
T8lrvCICjVJmsWhReJURJf0huHyLp4CRa/Cjls0COxvgJZ0RFNIaQqwIFwywl19IcZlRZ/wOagdU
fWb4efdP2rpcKgNgAPd9hLDRbaomBGVLW1XPY2SB9pCBun+S5eo9AxRd7VjCrZN0IfeNXX8GVsXm
DMrw4793ADa5O+t5ae75OHmzKNvpQddVzVX2HqW6l3bzGJq1vh39R6e3QILYcJ6lnIA5Pp6GGSUQ
l11K9RHEgzhthYP02Vg3XnReHyrptIBjX7b7UbABljyDWp6RC8TwfsIchAxkSXNLMKMAI/Eu5OjB
HDfFEvcNvw03vjUu2T440t9lLgOSc8CqwxHY/Sifo1PIH/Gzaf0tXLNEVJSCRFyULCqXWwTk89MO
mctAJdqeshLLJ8MuMOEHisHxsTLN1qHcxunt95FppSSCwrofwx1BR0tlcEwgCR1N1Fs8fS5WS6m1
oS7CHhQHr32I1gFlArXppGEiZg/xkdoTDvDhgWsyzkx2RsABohpNS96JbVuZdcvn58cv1L1nyHNn
XTnWqmqC2c4tHmh+HWf5Xj9U6fyKUFC8Qz/KNT4tsDtbVFrZ1c1wNSrQ0+/05TW4B8ZRNeHGeTRt
eLkXGyYl1eb8E5wZbKMsf4wIqgWy49MttZbpWFxJdugs7RdqqTEDk9Po24UqAlZWZNkAA55OJA9e
xB3FxiAF74IwyPiX+483q/DeVpPUrmBPqOhrEEtwb1tBCgE9PiI0cG+IuJxspLI38QDEJRhNDiwv
zi4awLFpL2dJKSLb+5zcD3CQS3amnAadoBOl4esGP+Feop23EDHGUY8Gq+lItQ++bcjIb0v0di4J
CC5BKiF4f1e0TXB6HppR3SUb71mBgjMQ0B3iMXxopHGmCZhR0xc22HRImc8vjl2GQIe9rM0mcenr
nVIw+Fvc6Xb2+Etb083pS9t3UaRyhF3d0HZq8BBriMUCv7JxSkqxlbtO0VwVcVMesLQzjQTYOtg7
miD+FsEpvE3OaUXz3m+x2odiYOtZ7HiqsdH5EdY33YXSOtoQlMhVEzkUNEYBSMnM0T3OZwYI9TsV
Ezqnpy5JuKuvodmvsojKQCbzeI3Kjr4wb/vqWy8lLfuIZA2Z1H7rh5FLugyx1n8JJmXxWGZ06ug3
njYMZAxIbWIL4uDgA8a/IUnA6o+4V/iIeOFK5UPZlctv69imVg0SQ14k7EAp2wO5RfAiEgNfIEoi
4+g+tA3oOOPzRe+AypGlOUYfTN4mjwKjjST5KmVqZbkWn2UmK4zxtwfygcdiyDcBnEspRrDi2cpm
MFTHyVOboJxK1XCsjyj3sz5HFzAhee/JLgq6xitZFK5wUp9JcoGCA8aqcdR1aFWjm5ECx1QDQEI4
U6mEtelcOcH0fsu9qV/GLqSIuT/Qb8mb1KBJKNKedxmW6ADPh0Qtrk5AL4u37i/78WaPdFZbmChP
2pEKXhniPKtXgJU0KVhcRRtLpV5/Wov0Y62fENvCGDrYtO38RCCoKpML3Oy8gsPewG90aPS1TEnh
qLaNLpjelU/fg2zb6wotokwhTqRlCnrgfhUowHcJSWHXn9wUWNniTHOcZvZkqjNG8zydJectX8NA
G+JzmSPJKkCiNNIVucn1NT8x0ZCJr00eLn6J7DJ+034JPAOS0rOSgQLAK2aebsA2YE3YdEoCaitn
3BM5JCyv1ik5yuRTWiXrjG6v49pdArcsRaGQfb7eGacktXfF1jkIv2iOT0rDUM+J1dtqFmb0RdVH
c+63drArTk2WHwuT7e8NFofXKC8oZM5ySbUgwiimRE1sUYsdvdJX22H+W9l6et5Ud8PwPPyxqBo9
1/3go+19YBjAbPsKbllS++C4ua0I+tLFtVBjrLMoe/qNsUz/xHUxJ8CdQ21j6VijuReD+pM2tIn5
5kYgLnDQpXdePQLReReYatT7UG38YHgsbmPuDBTdz34PlsOmVqKezdmOLlNa2fTrRWy4BxOtsoaN
GDxyQy3zsyzBSjHoAr+KdtnmcGvtyQ6fJP9bLKD0YoRH6ilGXRtZ6P+3GocAwGqexZmVwtIiAiv1
tjWQZJrD6xQl5unA74PqRXFctACqeG3Xp2QrZHuJDGe///N6/Da0E+M1hCt4oLnrBnnGMc1Up+ZS
8M1jssDaC27iYeaAkenw4ivGB0etbS48Wls/TNv/Ytw1rrUd9XFZecyfZa74+hzDyYEojPxhTmdr
Td72br2+8niaUAMlNYNY8GrXKRQcZqPxGcvV8U73onOipIRse0G0rPwFTATAS4CV/3enaZ31xMQd
k0+DuO9jidPgSc34YlKXBKrWM/h9dQp7ox5jYAT7/sijQKcA7qs00iMxZClFfbgz0YNnS+Lg7+Sb
c01RjPqi9B/7XzJ65MQTrTC9mcnB8fUW7lS/bVNLfR5FOalNoEO6LkIsU6uahTuC/yK5f7TpzY1w
4iNEatYqM8owlRFMUTsuOyZqVvyWM3QvjmBR/X5PxK4MdICZvJEu2wQ5J2fBXart/U9ZWXWuWe6V
zHi5YJVFDr1V5a/GKBGPfoc3EqSbS7lZRth/htW3C3I+oGFuzZVFOU4sokG53lmpqr4Fgza+DZBk
5NvPz/matfmJRGpyuda4hekQizKy5b6tkEvPfYLJqvMpY1o4WsMJdZIE87da4pUGjPJVfqr888DV
NOavjINn+XrYaiwuuXMz506Ndk66jpQZr9/2aANzSKpyeKvym0WSBmCCLIWvv69pKlDrAOpSSlQ2
Tsa+5y9/E4TVbFQwV2vPQoY443uIE85so2jeyWxeyHTnlWTjce58T1QBvgQASmq0bacmfRP3K3ms
dsREtBx35z/jHZzMt4p/TwR61rWTSlZdo1FQHGK/o+f1SmK/YqoJNjq95Woh37t7zE/PAHr2JltS
OEmHut6VPcPXoJW1GPzSi6orAaZyHtbYqWrPX9NX7Ia8Vfn01CStzbOJA/60TsTEtfqc4iHyiQEa
4LHi3POenZCWbixHhq6RFnSKXtvrDLuPaCrGIA6Jb2zgwsERvyl+3ud03CynSDihT5DmMQ/CchEV
Exaue2XQ4DWMPCFFtElyPHlL9pexU3Nm/AEkCbWZfewqEEWWEfYo307mCJHukNXcmudxPvUX62yC
wSDRq4Z8dy2m8GTpc53WnfUQjFE5AeTGhjp/finHmkhQAPUcui1eehgROxEA3q6cTM2UrU44Ciru
OoeuCTjZcJ4Hbh3iz/rMJwb1P+xUohar9rZ7FHszoeKHHHsIE/zVFZ+O3MzoB8d3BWVF2Bba4ZVC
bLFb21BC996zp/63GbjBH4A8daNGaY/j0KNWgaHc6Xh+0vCrhsCrVKMvxXG0YAepureoRKutpYXA
XaED50CRJzA29T4YEddFJrhpNHv/7ytPB4lKw55nAhjvSt+I6Oxk8eNyv2LTja7RD9Oo7lZhekI2
VHUwRX4bv4cGxKfX3TGs+iUn/b+19d5SvoUYTeJ4FROCorABOO4g8XYpFFi3zJSRXeUU2KhYVZ94
oU8H5AC/9XRAk+4y5k+9fhCHxZg4wZsTKMn8O3TFArJE08wsJfKak1xqOP9aH+DlQIl9tuJRGiuB
rqXcScPuITMp8S6kn794hWvw3AIWaATDrM/M0gqILUavo6aHkJgNptKyZXHbWUAuFLIjCsYNvLWj
Aw4kgcDUCoXJEmT2sfm2xkrApoAt6X23D5e1WftRfr6eHrI9uGyUcW2gnCyVWvFqe68AoB6y12sy
vhivCGIJEr7nTYiXjt1kaOpGFhpTkusDKL/5SH8d3POCwkCFfYWxspItZk3wuUhhu/A8YN8kgNXi
OtE82hU1ii2ZLRhEIGk9OJTZvsWC+b1IGAQ5uXNbdvO8UNo2Pj0E1iAjvGFvXg4AbTXfPSnWvi4k
MCQWnPX4Tafgmc+npAeqjXW69NJPhDbEtZ/UtCjNk7YUmKt+S+DVbJAu2lFhC8jMPodCUB2W52RG
pWLXpJbAmdmBMlXcsjLkFk/Jk9XoKCBNVDFLb/ExXEJUgfH99h/UXuke1DRhYJ7MUNum5pcd+XvK
g3YxpDviJ6m6nEuAfwp92B/PjGpfYprsVuMmqP3GJMuSbRazxwxpYGDcm0nRzTPRwn38s/t2hftO
ylzkTQkJqH9orb3DgwacVsf9zLKtjue2Wc+fuzMnhOJkhUFBx13CRiVPl5tIGqGaBMT8mhmufxLM
Et/NVijFgcAcKCKyaztBflvyuR+7g6B5ioNwwt/2J8dfu2END2UDIssVLNAb4JRUHZWx40nJ/iki
sUhQrLnjVsbqhjpJlp3Ji1JhebCuGDCqH9XSMG04u7tYYQXXkCcYIHJR/G6KlG3VEHcvxfTzKHly
VBC9Uw47woQaEItSdwpS0L6P3hgvnWJbeZqWipvtSZxNiiMDpXs7jl4MVBoDwKZjLHtCPVy7WhE+
5cUXJ/qG556bSG0YKs0vRJ/OjvAQHSy2Cm+A+8m9GsTD15t/bQgdndKjIZsW7KUI7l9kX+GRI3UK
kg8djmTps8bpUEaj+nU9jwy0jHtVNFBoIbx6vVJIp1E3IHXFZgt9lxgFMTKnx+5rWruM0+jmPG/X
Qh7t6pPWOT8Z0N0XMhwewaouk7AFCIqIzWXfJmHakDu6u/DUSpSemYV2CZ5fDNvn5WwgkPRFL6O7
8vzXUbat6uRaGlfyFfcwa69GrargpZvUVmdyiBvde/YVo0Cr2C5a1BU8ITlfC7wDVSvYEVjTeI4M
2phorI5kLA0L3O2c9u/QW26pQOm2RL1iljAjxtgluBAB4BYD1BJn0D5wnOTfZb/7m4iQN97qAcC4
ZBYNPaZwj4ywuJNuL6ByQNtmzLDy21+oXt8YRl9dfljTbwdmKhu5xcxER+Wg/2wH6U/vT/X03JBj
slVmIYNxGGxoPrytOz7BQiLzdMz5rubLIDdjIiSdtFM4uco5EuuFR36o4CqrS+lICrtKf375pb5E
mnvEyr6PORtcXwVvCC3kT22vVjMus5i7LK2+r6ctmqBJbDly1ryJweGzytB96U2ZUYEhdERBAKo/
b1Sv9Yq26wxn608HRTMreL1lclqhgPEbL+DavIsbE4WjqJcT8XQx4XFOA1gsD+IQbYCqcbiIADij
7fGqsEtEsEdoAyZ7DV47zD5PrrEmbzL6ymFJtgsu3UdQdKmjMB+ufqCMGknvbKZJWpK06ql0ifis
i7SyYda/poVmcgwwmjVpXQDDfKHVPojN81mWFFJUy2zkg2FarSNQTsKtMPBZ4nQfmYshKNVuK8mu
68cM8FA6j78lLksuRFyut7BSyCRZLmwc90vOXK+F4hE9fkOGt8noxdWugsKkf8eR2NQ02qJa1L85
jm99X02gatGOlyG5dwGUYlAArWpS3HpMoDNMH+Fkx6iBClGkMQC/n2fI/1GAKHhbLHcwsAmz701I
S32CUKhnjNZEgzIXwwTpSo3SmSwkdxEDmljlMpuUZbumKpuqoR9YLZrvMPWAp40RK1VQyUIuO6P8
iyl3GQ7X53QZ23YxfuL2+FbgT8QmhxayjB+q1VF+uEuPEOvPaMVUo7bLu6RfHI4Z6g8cmbO7mVZV
Ncv9SWmCQDphhwxPG/P7vQVRxjaM+8BX7axQsXUaez+uJh7Ynst5lBfEmjmHm2r0cssEZzJnjr/x
WvCnNJ3/gBT73VCSlSzRCcbopydoM+9mQKnOY4I5tpX8TFV8dYUGgemqz77Mpo3T3+G6Ts8eYTFV
yuZX9Kf5UU7Wrd5D+Zj0I1P9tgmtDWYrW7om9G0h4J0dDwp/XIug4MCVa2m+zmlMlwj40KvXmT+8
aMgEPre/A2J4+3bHDF2z9PTzxUvtrqNgqph62xkCsIrtFFnqXJxt74gdA2OWceOIzYU8Kd8U9hg1
280UPcALTrquWTvchG5ayeJxkVPRR3vgjXTTjpnIvNgaK4DX2OqRTnFrPIRE/zwwsA6833XtFI6p
pzRBOQq+xpxk+f8z5EHoCJN+/rMCHKIY+FpmGtSwYtD7UsLm9kDoabYYtpfnWjjFaB4Ly1oo4XMM
raVnk22f3NVwR3P8nP5isfoYCOVqUxdbGU8b1FxzFFeWF/7MJy2HTQjgM7s5iKfcpAV4SACBS61Z
Xcp7mvTkeAlbSyebzake7IJvhu0jwafbVTgutM1q4qrR+yW8qX0VEOjksLadYb2T0M6g8KKDyTlT
j7Z//nQ2DtEwLnmS8VXm/pbbf5nWbzAdXNsxv7u+E7X9zlgK1qdbcT47feWqVr3mUGk2YpXSswEk
AbHGfHWJ5pFCbjTwPGl46kWbwSmTsS39O+ETfySIjTsQH+HnsIcEbpoNLWifXvZhuwYoRr2GADEi
rV8UvL+Hz0S/IgddBvIe+p51yC+PkZg0mJwnQJIscndkF1GR8yJ0etsBGxHluvReHm14ImcAmIlS
w5CAiXBlEkSKr2HX7r8NmK95iJU+yOpB1WzvPcGgaIYsL36AWjB3bzKQ8SnWE3QALa2CEF7mb0/v
jpOffpfQjlGXo4Yy4tpfuOlyGjL3HbWz7HzCm6rSrcyi3KVRTmsNmuSNzjcAZM/ia7MUGdERv0Js
qx8VJGQYUofhxS2zzcwT8zYCt2nqRdqc/xJ6mEf3wXGaUDRASDMT2/HinNK5m+aOUCemcJyP/5UL
DBzsEZJ5zu0Yq4cJDKlqhX3hNHj8x+fgiuOVi/0lEPeKkTEP0SLv0kS7pSASHI7r42DrT+/ls1jC
snFVWyOW/m5N7TN37InaqGTrg7HZ5vs61c49iSBKuh5lMgp5dBqxr92sr3w0WufFzdsRX6gEynIt
RnRbLKJa5bUG1CT64hfRcAiqLHyL+v0ZBTOPsjhjIpNgecPUJjmtd7lO7BLr59VWLBtwF5DPkXyN
zLu8zcHRoqNvtTg5CQi14lMX+SEonL/+Pqxis3lIpQlDldOA4/uKwbDrwVfOy8ea7rdImBGH2OKR
/1peteH6Rt0vcXb1VOAZPDomc4D8ll76wnqs4O3bk0UC1tlWRQkPAlCqb02H9mq+4h5QDiQ/osjR
R2hhmkNVMVjb6dGt1SxiN81jRgE94P7Xa35DUydSm903313tk+9bBTReBNoyWYRFe974Fpbd/kSB
zhWk7LhVI5IeqBvL/SZ4W2vEQUu1g8xu1VQJtn4DVw+z1hm7FhSpUM7en60i0Ozpcg+4Qp6xygtc
Mzi1AtqeOgmirOb2rNRBIWhLh5Jk9s8jGePpkgVDsgo5O5uqYHQ33znrvWw9Hhlt6niubrjYZ3F+
yRHlot16ldEo2pnlics7qkdtA2ODNsPH0ZjsTicqWiSNhbwUfEgh7A7Ik9+/9weXx0UqJVAXVjzR
8zk5aQfSz9PgKZRO+r3YHsC2gMhqcUyQh0O7625flVGMwQn82+ayAPZQbfIb/UcD7+xzpkNOlrEt
uHj18+pdHl7ZIQgxBf27PtwxWUQXPLG2DsNpbJQ82b3wn3Pev8TkarOFC/EmdLFYHojzWVlf6Mol
UK5H22CnLtwreIW7wOZM8YxGCcm0V4K/MvoE/5EwZEswIWM5buEaqV1H4MsQORP5cR5Di1lHwx3t
uy3fligDCog3uPD8LXgqsYN3u4Nf0AYlU0f077aZJlpAB/ZaTzpzw2vuOp6hlvdJmj/qPMXF6TdJ
mM9rj17oxMxYQeoO4FV7vG56lykzywM64vuWz5Jv43GVomrJSkTzr/mk/yU5TB3LdqLSXZS+xKYB
yBkJ4vwkm+a1yoV6/am3QhDlSexK0SQTZAk/SOChCPyKBHvBBnFIUZ2qE7AMh6rdjQY6p+F3pKSB
cqdaAkWoWVJ4a/751E6dz9bITRdw/gH5tSRwN1LBKQ1W2u+JVe2JAGNvtIJLD8JGmIUv5TDT27y0
DwEdZe61sfJ2pmGxyU4WEtfOLTCNpK3LdbFJ2NboCgS+e8fmXm10+TAztXvYNzXzOKANh3ZFnjZ6
wKlo38rfrIQErn2OhHUQUZcoTJgFHLW1rFIFHm08XpDBcqDyiFjt7CwDjnhmyHK0Zm/uU8h8q1X9
hcd/QnCtRSKrDzbIUXtuJAb6HCaU8VG+AOEepz8il073rxyg4TohtvTQNIQ7K+jccey3rrJHcxai
B3Qkfaf4DTFv83iTEgxsFWmrSAMjkybS/cd6eBnqSKNBdzB1I+OmWXJC1BlzqCgZtK6umhY6G7bs
rinGFVbjorr9Gaj4isZPHhyrXx38hOhIlMRlueylAnjDq+3zWXR7t+iiqI7pFe2k/gH7Xl/gEgB/
9BCRXEArnOwf9xi79bxqWYA9PECd0GAYjPWpQQ2GFrO+O/AZ/qb4YnaJYvHIYgBL3ShuMqRvJpK2
1x1w1nbVS+GWAi/MuUqGMF77eHmdk7LTOOwqjbJ6WrRZAgyR8FnnRtH+PCL0SemtBN/jnvztIaok
9e9/oh+jgPhXsToEku7sMYENQr5vocJnv3NiFxkiL//GPL3/FctI4YGqnN2AE+wsfUnM+L2gadyI
r6oBi+BGOnA+3/V+JhLtaM2oaJGz3x6GnTykrkBqdAFaGrS9/kwMvRGh1/wYLggygH2rg20Hpc0m
TBWOo9VGq1IGLPFf0aoMU2UOpxo1BcccozWXYPoLCra04v2WAq9abDtqaMLzXX2w7Mn5RxeAdzmZ
kLMl0Hr2yYGpOq8AT8keYf/Dxt+avcFnan2pL88xb9oPsEVe34H967yRGW7r3QAZaRUBYM+oheuh
gJXpoRxzoOCWwPqni92+FjmzrB+BC8mSGi5HHj1FBp+MmXnwrRr5rVmv38m7f2wW0o3Xxu1zqGOz
Tmd5XcqI+fb+LbCB2XbzHcMorSyI18y2u6rtAZBn4sn9uu/xXjmkWKlaRmpquHonW2SZObwC5oDd
u1qI1OA3pe6Ez+bZicOhNJBudhH/W06+oYZiB1VbYYt0aAJhu0zhNYAnwQNQoatl4k/ZdiN+iOQm
zl5bwba6f+EpXeTuC4A2gB/NLhYllhocNIGme4ShAvE/nJkcKmt3ZEb1/5bVCYPJ33NrHY4kLU3w
Khqcc9pDevoZFWYnI6R8lis6V1F5wooTyx5+DhRZ2QCAWP8WfbrXGUQDHovobwPJXwxj6sWETPdi
Eu6XGA+QU5Ix0b25xShzTegW7aCsQI7KxLtDhKNGS08fw8PqY07q0P+bUkwLgNkNZ+BflHC+aXsN
4SxgOintHXIAssJ+pnAzwnuLNaz384LquGEXR/nMqtvORNNJJMNLfX7qWtGFadxZ5NMefstZxoIj
wC5sQakFHJs2/mnHsO7P28ZdwAmnIs5sszGpIOy3myCcz3XZYb84XbswzE9xO5Y2RUoZ1G6hNu29
vYsDEowGMGS6blZxVrjusC56o+IbTy12R9GOLBAUzDZyeM/Gfw3t6fZLcwRE3EGST+rgqhlU4VaR
kW+avlM23cLJGkLvWb9BY8yRdUoDQlmSr6fedmSrdKuScIa4bGUCXPBGMPyxd0VxPQFueoNyzMrI
8nuZaWOwXTyGUlNJdFlnOirkqf/x/YAHxrcKI7gPvm5JBDwW7MGVcvQRHXro3GhAj+F8u3mVH+My
a78KBzQOy+B3JiX7LHqC721nvtX4lbB3ovLhPBoyWYOGxaIBOJfosr92MwGx5EvnX/OgiCulNzgE
K/To7iwoQS3RxxnLG91efTcUjBeriN55LQGe9Dsg5j5Fp1FWNEGwbbbAm4ilqjAOvW9txIsx9X07
Ef7S7QoYdCqGGYSzbL13of/E7g3ZY+/lq3zdgXPPMU2/Dw0sdWYwiXeBuR/I/r1INdRKuTFRr/au
BB2oEc2XrD25S0TP0H5zpvo3vQEXnDGCjfGCeikefmrkImMlu0dc0Ua5Pa3PiTntjUqNLnXrmncS
skps364ckXugosqciN4TCtYXJd3rnPrh/72rJvvXIxECv1mUDTz0/KGjfdiywIPpi6sfMGdaKZpm
xTm3WCeqAwaevnlG4xkx/0H9Ln1Cf/qmSiAkWsghIcgkhqrbEGAf5cFKv/ALkxT7UGea87nTMHOP
fBtwulJgxB/Wb1x5nhSGip4y60kwT/c7huPC2IyhwR7ZF4gOWtBLHw9UYssWvpNKUVAbWXpL4iFW
6Vi+w9qYp350HCmoiPHbxFbgbtT5XlKkqcbya9DKyp5oY2LgUTx/Zth/WTse+PCrUu7uPC1D6xTb
Z5oiiUIpMKtQapC+PYhILpbeXGYiKTp/JHMPXgp9ksBTz/zuLncUl1hbw16zVf42oXwierWUnK5b
EOBlsjW/n/2ekmCkGvFwpUZuJlk/F9j/Paw7fwIwwV27f9KMs1mtHyn9xKQRLES+vfEe/z2KawKe
+U8hPY4LiXFjv1VufU6PDEt+vlqHY6exDoYiqgSo54lxjFqsI3QP6+he6oEwTVLbPKFR2t2axFBf
CDFX/ZKBI6Njgh5E0FKRdBUosykw1cQh1v1oxBJkZ7SkstmkpzukuU2PcVOliQDwECg3oyYqt0Tl
jexozTimp2XDE6Mw+4EPoWZM1eUMinADTkz4RU5a8LJAATbZCvorLk/H69pTMAaMDeuGI8FbAbXQ
GC5azAnd0szTg3cqgENgKIWAmYqHpX4uwOdOtf/9Y5P2sQhHMbWvvK95zDySP1BQu6EEnp+oKEnH
df4QFA5EF/2wNh3/v4sIlQn7JiVghOBN3gqqXkSU0KxdOvBjYtla9waEccQtsp9btb3XEJw2HRbV
uCTHZH6htvWeqsX610yjXrzqgbXRCCtIl/D5ByeByGLTmAUINB3OHIzJT9TFlwRhxSlKcUdcQu89
7UtjS+PrPZJtXWxT4AaGl9sMTKzNn7ctb4zMXFA81KJfUTNNjJQV4ebt5Z+3UomNNByjs0Rau7Db
KALZbo1XbRY3NVaRzZQzFps3QA4Vm1rS/BhrgRClRiP+q/iKtjdxZ3bT9soxqPyrtot6fSvb9nO0
RQUwPmBE7uD8/1LEnfKF6LQCM55pP5RnQDuYwY/pWADmy8txOvWRZ2+VFxvNT5Sl7PcGxeuNcVZJ
PxxhnuFaf1hd6AyRuvw43tHSy9N2+DpABPT3jtfRlONvPShPZWDt4Z0jiEuFRbWWULIdX3ZEStAY
PuOX5ixahSlPLGpUglXsXwzn2liQZP8yq6FH7v+5JJ6gHvPCnacDmRgtQ7O/zNuy9dEIJk9MlzVj
vNq+tyh4q6itHq7Y/+1vYYf84K0SRUQYKMoOAGa2axN1PNZ7/ZFu0mz/JrIcPhmTa+oxdLHt1gdZ
JUrndKhQEKkt6UnO5X5Vm5D5p6lriG1fBJEBlrIzIfOH2m6+t22Q/48Nt7w8XHINF+0lhbXrJNlv
+IuNSNZt9TKKmNL6C30I5OifolYSXFxvNBRftbMPDXPyjO7WMdv3Z8hT8nh/qh+Dn/m1QmddSoIL
RiwDT8ZpizPC42qKjnZ00dyMJsach/CFoGJSpxtGRHfPxKAwmseE/ibkKBcfLG8YN3hNl0RVHNv/
EPKY01NAzC9mBvpIdG91Sn3C9lc/RQMU3rogxSOJZs98pEn5+mZwWoFOr8WGmqc1wHNnam8BvMyG
gEH8JiaeZzXZuGeaoUueGmwdNBVTo2QR9eOdaHS2TBya8CS1s1a6Uf+Ma5xCEs6JQlXt7T3AHmUh
8qZ3kB/S1nEKup/6YHacSqxxcI/02zCxdytcOETUGHDimP5Jluo/e5wWwjYcAxQBTGV8Lq27H/Ag
2tOitAMmfGm0mHsZfNaLx1dp7t+NpU3gST00D2OQWA2se0sW5Uw//f3VpO6sgSIQ2y9FgcwuRLbM
CGIv8ET/vN8SJILEJ1uJQTiGlX/E5d5b62t/GLkF0akZvcvPUkWPhFNGg+eoF4Btl73UYfUswy7t
gThWM/5iZm3ITW822V4jZ7IzFqUBjJxHEH66q7OTF4o3TD0agP8vHtMBJslLOacRLdXT5J9d5C4V
yS8HtreClCgnU4kfKKKCLAo4xrlUre05kg3uf/br0C6KmOxKsG7R1i+VwQ1+VUBYnL7MCOalOGdx
rLqoOFXKjUmio92Lr+qaesj7EjfvGjOeIxdA4Eh8NVmq4PVv4Ba8uI280pOp+O0JOOfJ4AOQRlof
S+vg4ffqXMwbg3a3MqlmmRKhtLA0CnEFcnRKFbBFcTNzTSNCNE801E3dC610KOeWhdaZBvaXch+D
2/6QdxWjXrKt7rpDzn+0d3SFoW/i7fs7ziJZr/gz6UED36B58ASf8hU50oRvUN48Uri7/kSQAEFX
jKGfGaPgs8ys11LSrpg94/9qHQZ0B+oqPAu5oJiQw7tNCcSVrhsORgWol5R0rkxcXyUVS6l20w+Q
MC0z5kHbrHWqAn8Jax5DH2d5bKCRX3M/GeqMUnor9PFY9CAcNYMU88XHfzqdF7ZcvTVAdU6lxTlM
bS0+v4WkMrNJnVs3DkbX5x/ejydwjPDA4XzSzv4SKhh732Pgg6+OuMNTezej3d4kSUw2q9hTUjNO
lrXK3eJZw/MOSDGGEEgXCP7yJ6nXJfzrK3Vfd7Tvhr3+EEmFB0UQ9CusEz6yEm64eaT+FBOwX0tU
Z9k7r34FeoUW1ds5wJZ//3vygIqD6NHKP4u32ZDW2Y5jbJKovQ9E1ilxkno+wY6tDVN85ulRtMeR
5Ei69ld3HdpfcGmn0zQ6T8Be/+2n/nuwUIHrUCKThrAnx0L5XkHuytnjFSj3mnjUyUE1Qen2xT/0
NMbof58RmJcZstmdRYWUM/dtLh/bJ3O5r5gNi4RQTQKexZB0j4P3V9A2VMFYaqE3YZFccQERChqU
nmEr5QUUYnifQBO53p9iv6XZcaQCdFB1LjsZK3ywG+Z4LCVtDDnmPNlqOGJB78UlQyvWIVJBSdPB
f8xwEXD/hzw4KcD8v9W3kiQEJQVfrXOYazwLJSM0gjNTHJPqmBy8cK9cWMEhAxam89K5Nk/bWPWh
vb4V22roFZ4zPzx3M9ao81EDpvMNTFW3JJiSQt5w+1GXseF3F3NV6JAjFvwUae0R1uRXi5lQlUD1
r47iFS9XmfFg9z6KKXoa7DtFY+Bqgv9oK7Ybf7yjilNqJvEH5Kd+Vdi5EFVFmiUJwfEwqmf/0HFE
V8gj/ymhQMFPrp366t4vLj/4CQrh+hawjIUXL7+qj6ePAQejkOi6vbBBGO2c9SQfigIWzEkyGUJI
JsCc2EVOHiXPPCgWyku/zJkymayqftAKFJHVMCkViKHLrjGkeFQTHf23DHput18hZwo3KMzjZ+aq
GD4195Fh3cEB78C79eOOga8vNOa9pbvbIIsuV6xAT+xR3yIceidyHIV8pKAbPB5tmCjplvosCXOD
ew34n5VGDHUUSwxCunWF6G82aPYOmmAmO3VuT3c5HGfgsAGcVrhyp7NaF3XrsyKGeuXJxtLniKUV
nnVXoEHRUQuduoV+z/LaE9AHyzc6mhyGLfno5GSCMuoCNfZRSLp2fwcWxLnco1mgrav0Zzu2jlwM
0zwoDpOTwFiP/b5ibcSyBprPYZcc45L0fM8onEMdixomrqFZk/Wcotmtw6eyGxZ6rIXzZuiEuXea
JMgCdiMJ172FKSdTkK2J/ecMbQOJTQnPUUz7ffaR9THXJDKQGFxgNU2jhFVI4FNp4Kh97J5Nap50
+EKinjEcETVO68RaDfkcgQ3/6/qLeFZHb95JT77bigFQqiRsKfNVn+Xuu5O5fa1lX/R21SF7mmyT
b4a+fYulC+hrtzsSZRH5HW/iavC12wbt7aqOckbQ9Gf86cM7dwhlAdiY70OOoTlaXZLm5UxyhlYl
s87k7sNegMb2aINsGI+0X4jNUb4maarJIM9UI9aidray1y718tXAFAg7UumwZ2SiZLsF41uYTkCQ
KgbmqxS5JtveT9qjwu2BMAOWoFFaRH9SMABpF6DAVagnouMWsT+S9HD0iKPuW9VgfkTNX3UApCqN
5OUqXwuWqXEK1FMgTz9loSgeS98/hmC+DVt8VQEf/lvT1jYhSdGc44/+uR9qrym1tf3994P+wac2
jorHZgqF6ra+QBmxlIRKZiz7zyL9/zXFzvApM8KnMZuXOIKEbRKOyMLU6qBq6hq8lmw2vfMjeJLq
oLWmDN0jixOY2T+Rj5xYHORDonByrl6+2VxA63jhyifMOnWo8RgOvZCq2U2aoOjA1wV5QCPk+Qc2
E6+8Sz47KW5gcGvGu7p/wRbB3sV45CUlEhRusIwZv8qX11gx5UTqe2WCPewpkbAmqORt8HNyuYv0
754k3cMO+y3ob0nNa7P/6Ny1Ahp2aAQqU9z3vSFiBBqCd5QFxc6CsXeeD30cDDhelmVP9S6H41As
ZJg+PpLRu9IROAVM7VA0tKJ+RxYYASNGZ/EHnca8LBGw7qzxMcoqSWEhF7bGeyKoeo+ME2x4e9GZ
6P65jKLOJehSRl84iGVBM05zEdt9jGNS/AU2j2tgFYxVVfnxj7XE6yvuVLIbaOAgXvoZRQryW/FS
TY+dOiF+TGLSKkVjSC4zIKqeiqdAVmy5WnChP4HKukmV9E3RE0PBVEwxiOqqrzAJA2Wp4FZbuCVD
P7YXXRir3XvIu819mTIYOGyeXvw6JsqNMibpzFtK8sFVCFiC18HLQpzO+quM5jyhoYT4ZsS08WuM
ywN0WDnyRmLB/Koj0OGZnXmO/YGKcmaCSK3On9BbXbX8VqN8edM0Ow7Ec1U7+zZ8jxuY6xb+FKmz
R9yKGTly4MzA+Vlf906Kzc2XL6ZHQ1AQeowEoRhqJG7+ttz3T5xXA6aYIRg5ftD2GE3sxylQ2MuP
Za931mDSY/IryPdZ3fXmvUBw5Lc1B3OzkvkrzRHzv7hGJc90SK6F+gjoNIK2NrvmUdzcz3IV0I6M
A9SMcOcsz7Gt36rqYutYQJc55/lFWkRfDIZzQkrxuYJf65fAf3vv2KHWsAivPwJLjYNU260GHFtM
tasVQrcB864rB5IFyZij8uCdW862wxGEyxBmP2hHsODTJwrjmpI06dSuaDLuJcvLTi+cOYyknDcp
RzdybvE0E0+FiMlH+VC648Z4dZeN6S4KfYFvQ0Wyb/VW3M0TxQFfvH8eS6f3s8c5EacSTddbFM1U
2Y+SNVEg9Kr/xnJGvVzwTdKR1r9kH5KPBTMHcjsrhziALXAPK+rZj7ebhiJDcpjGYJ2MTUcRbchX
WLwWrMIjoZpVT2nuWxnjOu2A3NKfn8DR/l8toGlenlI9LBTp8VJ8+YbkPefaaYxgG2ILYwfW3pFd
2vUz0JlD09/9/nX069CddtblCwNJMTb+FDebjtw3OLBvD9LFow6AX1tdqixGKSn0YDJRJ+Ajlz54
mvtnC8F9A0SBod4vNvVs9WSGkFNGtGf+7+uZj7Mm6yQqnYS8mDIbTg2WCxpaYgMI0lvf4kg72r3C
vO0V47+vRFkWJlH7lD7n4fLdN/7qr6vBTR0afFEHUtQhzGxXyBNNM7mSDsqCNR/vE4fCT8bByO/B
3ty3BnGfGoczwOT7GSpR3l6BtHD2H/EMR+xEmdSnTPF7Z1o+3DFilgUz2W8IogGj/EtzOQGqgr9M
dRqcG2JO3yNcRQv9qOVCavCHmWm2CS8TWTgu2+jVX0XgM7qlSnK8K4NJGu5VlFFCnAqpZLUfzRZb
LJ/mkTWR7Clv4m6M2+i6sDynBsyqt5WSCPBTN+1AdBqyAk027BCJxdR+C0Kyktrz35Vjl8kphrBn
ZPtKDsOJyGavmBwnhdDvnrPo/40OZMRpy0j3YVaoVVijk4goVP//pOTU3fIzAckYy3/FN5hCRP5i
FhidoE3ps1Pm0cTJdXy60lsDLUUFfChMYch2knomibBx6loEkClVkQrRbX0ZuMtc65yK0puyhfC/
DxzlLpTDdYCtc7D6X+jl/HiMTULhT1SRzrLFd9G+GAoxK6Qt6ogyO+Di/WBOXw3NgBpbPKGuorpT
6eB9aqy/LLlqvecBHk3ugOtLzx5E32frg98NnBibAHkmUH6+4loiZKyfdN3YWBWPoIcTmXxlwcQl
mFJAZOIoFB2cQfzFsbl+892bI8pn9Nw48WFdO4OfX3h/vhjEkTVYjJWvwpBxmQXPFMitKrOGalzV
a+RSEU4MerEvr3lI8FH1SbDj1LuuMjS9xxEZtke3BBmWSa+1iQ8GRmV+7RyZ0dkmok6s8eayR5VT
GuR2iOSFa27C2w1QuaF2BROO7EjcVpUUFpY9gg8vJHPaJwun1CDQ4In8ScaOV4bSQypZjtm1vFkq
J4j7MbHZUqDzCdFDyFhSojhM0b9zS+2mzEksPm+W9n2d43/HDHjJR/C/EdM5PsciKgdG3oWkFP+l
aX0yCkYELoRnaWyfNYaMYGRKpJO4trSEx4S/+8Z0pRFMSqcMtrLy3QPbyyaYbYPchiZlJIUqZJ1K
PVBlJsHJe/TH8Y8PBtZ2HktQFVsT4o+CHBoEtPZV8V3u0Bt4g6jdD2a/9T9m6WMKYUZQAr7xkka7
9et/k5zFHQh00eIRREfGSOYym9WX/KPKrZ/scC094emKoLGVACpoQJFVEFA2/cVlupxcDCE+0fxY
ezDmMXPGdjVDR826H36cetsbphj2vLNWVEyufz2kbfWT3QzLN1ob7ntGeB24MBY9pRWAPd5ssXr8
kKqXxSzxwqnvJpY093YNvi/bc0QDFoARglJS8p/GqMSmGV5ct5a777Wo7S5Av/yqZad+/Ggha6Zh
WKoBvYtXQvLu9EifcPo7DIZ07r0hXonlQcqhi0ZOdJnKNihfcNpTo/zswkeE4+/zMM17oGco2tc2
svZziGNLOmSJriw0oadczY0ok3YzPLSWSFGC1jFlUWOTHgqay4pKQULAB6V8nafI7BclfTQRCX/S
N5yqLZ+xcZ+18FPtcDWxkoIDs8M4WjEXAfXfYOdEi9aw78vrcR+jtwdgS+X84yJQhGaoTa+uZaBk
wuOpZtlqMQyualQDj89QbS7xogf9Mo7+XhRWxtz9cRFUB8oRH1rC2m5GFo3/IOKacE5303m/E2jo
uDAzjf7NmnWNGP8rFCLnn9bUTLYT5l49WDjgjUn/VOUBgoqZRZPfymto9fCmkrM9CD+g4RBgiYX4
17ytWD3TUcgNWSQ7MR/s/ibx8JfNA5VH+Jq+zxF4Sbs3IuoJrfUGypJW045Lcc+KGwwvtuNOdpi4
ZTtCzSSjlIwddISrkvzh8UqKVwEfTxw/C5nhznKy32cABSIIVLjCulHcU+mTwZsE26o8phyg7J1Y
i+1a/xpT4asQ7Iz9AoC+T23eQFJS+O5i1k/JdUdJfG/P5K6v641YqMSjHukP0g2/NpoNjRtRASlt
XeSRJ4Sl7/kKXU7EBwJBeIz8+NyfnjwaAGpp+C1jl+xxmmbfUj5WZwnslncIadiL/87WmIFMiVZ6
MqUJ55c2uQ6UBj6cIYHQqhQVkERe5VeDL7tL1Xx1MIRtEZFx0iy+vWR0H1RRemQ4WpZq4Gdvwm8/
JZS4a508O+SPmBaHeK60kczheP2+XEocDe6SIfb33ftMfHa+HcU/1nYNzPYbQ5aN4dAzbOtGC5lJ
vDf6htAU3Pr32dJK3QFNKnGnKKse6wKXjb1Pmsm0VpJ+JwgsEdRwMUVVcC0sHDnpDZK16Kw7+PLT
//d+yr9rh4QQW7mCEhy9nBCvlvwSKLsV0X9RAJa2E/ZlObScN8SAgc54+I85kQw5p/JItrdMeHeV
dh4qbIXLzhLuR4Ta7O4rnnZAcyAcJRJVKoVfhwviSsg5n1U6pPi34QyegbKb7wAe7lCB7p3rYHD+
xqUZ2ubx5MgAC60O7q5YG72uL64Yp/WSGwJVqNGRmlPW41rqyq4qDR/keoV3nQMQE87umxtQuZdi
yuKlABgY/nKyflA2YXX2O67JxJU76ebmelNlxOy4M35vh/lyqnDJ40FxCBYFIo5rmtCI3WWdZ0pA
RZxe4k49bzmwvqTIPHS7fsV9yC0q8zXIwwvoAAlaaSsS2zfdd4U91gzL/7oByWGtZuiAAmOIrIs/
1Guzae3u+ysAkJUhAeNttRB/2cCNb33EpvSNNyHcZkf7lHFK3esi7EpmJBI7p9XdwsJZZyYSuGF2
XsEV1S4IHCFUfHJkoIsELSHqv+isiPnz3eAAelulT4KnK1DOZWmvQ+WgBQjsIJbDLGAVvpeXrmvG
trJOqmQBBnD6pl4j9cis7+oh2oInS6TYAZp3ACkfmHzHgqKdj9jDILW2aL/ll6/ig167U8Rp2pXb
9CMF5/MK/E1O1sYuYPLB+HIQKYabqTiIOl3e2hxqgzG0nqBvUV76osuLk4x68IoBqW9eND1awbVr
fh+DEHsSV2Sy6AMHmNC4BQEYB7lh7B/AhWseXl0QW8W7iykZwsXDNXRD7EAbnVBlp5YxqArl+oXu
Xny3jKnGvoEWqa3XF4Q1xlIOIrz1GSzH0Bspoogmnd87fJzi/Y1Q77kQZmOrdGM3L4NNqUa/RGaL
clBdU4eht9K4mXlSzruF52VFxzYOmyoqHraVp1AuE1FejnKaxRaXST5g+pGB3ajGrOPkaQcyuq9s
xf2uPUlLYskxDjwypc4Gr+NtEHO7xSE0t5sBtEGAzTeaPAKzfkOsHoa9YCWhwYO2Etkz89jZt3Nq
YBUPKqr9mc6vbISfjnYhNcfmyPIXbj2gAKVpk9PpndZSYUjTEfXFHYS5oiGuMFXagPtR3fIgnVDg
/EnpNK/aSmlWWnx/MD/OZVoDyNLU6FKdR21d7/b7l9X+kquIjtoCitxEvTG97B11uSI7TNZHJ9Yf
3rUYoRW6MUJXuq5yfsmrvR2ePJ/eGlmiOW9Xvxp8wCvA/mp6pdhDkiwfKuSpe2e0Aom2Uo+aDdbh
ZBqs9BzJLDKwJ+DCDjBJyNbDrNOWzc/mnDvqEWO5cwtuchb1r2/+2noMB91sDqk5xPi79tHFb/MZ
DcQkPIfnmE7eE3a0N6HF7BA2ISom6JpxqRDs6bilxpF8S7ayYg0XIX3cn1DFllh+zgV7mxMjOB8W
YOmOiLmD382MPTuUE5TuItaa/pqBlJpYTeWIcjQ5OdgFREwAJH9Vo3YY+082Q/M4eHHp4sKMToYl
5NTZ97jOBQGeILT0f4n3ykb+ILQ+XtVj3xBxM9fkRPs7c9cs9lgok3zJ3cb1QaLP4U8VXiFyxVvR
akwpSunNLsxaV9s4Iwxrh05J8Su/hB+eI6vwgbMfVh73yTYNRUkmNEu7Ujil0CjGs8jXPiphGIDy
8DCFI1vHTSXMlyMpUR3YYNALWJhzqHFC44oRanYR09iku1xf5zyMpY4QpfY7kMSAP8BhXYF6CsLU
TxDqKHmhHrc77US9zQAMk4hXDYdt3HnRpOLT6fM/GwzmNhrHZEPMtEgDo7+Ow9Cz/+81EWyWgcHd
vVQJsVVDf9J4eGsIZsYVVrjNVlLcnSlKtvFyFBvVMAoV32+YD/XXT0oQc9X3E/NM6rL9+zZjsQiy
AcC/kkyI6B4ZkZS3tlD8KRAxtXz53FkqzrK4cfio7RNrhnw3JYB/4DIrWtnaL/9P2ughF+DBWLD/
yQ39ZkGGS8TcnC1Gn3Hhn2y/ZCFpstlHuqitq91ReuLGBXntb5ASRtpMwR4wNdEfOBC2uR9m4PZB
31/XNPNk3joJnpdASAdxOop4k2VEGXlg+wDxeeOVbMrudiSzZRYF1Nq79u1OCsUB5AqNT5l9O751
Xf/Z5smyTHT4O7C8NDcTwk7keYAvLUpv97Gv32YCJAFbyFoe9243pve1Nu4t5Jo2Zx8Gg6sA1dN7
x7N22SJqpg98AUVJU1CfttsLtrm0kVV1THGIHkonykBpH12WhFww+8Yom8nuAKZYqVEqt/t5AUix
33aUYukWlIEuoF6+3tGwYPNt/FhilwK1iqN/aMwLAOLSvE/7amMn2X44u2nixzZfG9RQ693CH1hx
9PtnYtPLDoI+bMbpVmAWKwzCLsyRJ4XkFDbu7mQDQTFQc/c9zEK07dSZfBYXGTQpL94UC5g9V4fr
HwRDlKjEpQgploGkZyUHyrU9GjXmzAFdStocRaDsxdO1SGzrgpdhTaZaB2kjAWOnWXKtWFh4Dvvs
bnf6/HZYSjKhDnfmkCpJLk/YdbCxsvVg9XqcnrjKNanQE4cz9yAO8CqHiIMPoAkfM6/tBv8qp/ls
5z2IWuE/nRvxfPf5XcFIyzs6PLxGT/NHzW+7dXP6dFilqjs3NOl8mDdoTzJvRoQ2Psfb4mw6sX7u
wdEQrIMxTDdtrZHjuuDHcLVOk+mmZm2MafpK/VNccnv26y4vP0EMYzufppPYDzmZ+NLP6Eq76GaG
0Yx8JSiO1ACnGFX6nZv0nLiWqH8xdX545rU/nWJkhJPOYq7vBVIDzS/JZcjESQfAjC9ZiieqCMOi
4tvgvXz4Dr0jGrmOH7NOT+Chq/WJRMWjfICenrYndJXUPdqPsI9+Oo+BOWwcf8XoElIlQAEdlple
fkT9trm3iE4J7bYwZCRBswg/lNYPGol5taAJ45yXEBmVtgm/8AWffKr2foyx72Jks6FikKPnyaO2
C7U0/7h11MSMJCdupuOA72BbRKk4us935CHrt3D9LGYutZhSF52CpgQ/GLHNXnxg9QsDLkzllCN4
94yHiRxIaa/m7STHkwZ4oTAVCoL/b/txCVkwCugps1Ma/4mxZabO8UqTcBMlIrRid6bsFf8nI+qJ
zDf2U2pYA0lY9Z+CdOhyZCduy/8TuDuB1QV792T2BAdHs2AEI3hBl34CKtEhnfGhI/N46TvBq3QY
XCKY20VFZkbYA8po4fzYL6lFxtb2gWUFAdzaQarG86OPcOSwS2srpB247wHe3kmv4WJuA1qTvPxl
+feT1lkiW7Y/rQ5wsl9E8YqZsFE9m2sfSJPL1F34H+VJVOVYrniz8JkpSSjUdDkTozQUILA7zXzG
IbP37F3rC4mKLiHgT9pfgjf897xa0WBgJqbfKq23uXLZoV6izYSyVRrdQAeU5/s9aLeI50gOf7gt
kYWrWB4a4pRj8Q3HrVWCRuDS8QnDVVqWwbcUV9QRFitLditYoII5iNtWBu2JHQf5MWfOknLsZxdv
leRwi5PV6D0DPpcSlFvfbJy+o2KXanhbZsEENGNNFgdfeBVkx1qdwMawYXGvzfO5piAF9PKqNJux
D3uGPeA/NLPnzusFcQ5FcPq2laEVyIJZ0HVbLZXwxFFEmRx+NB5fXDiFATB+R3ZGVZPMZCPr7aWU
lfra4h6P3dHFm/G542CtrI+b3nE9YTIeNV2v/iHQt4blpyXgkSsRXcwejmwK8fvIvZFTWDpiBP7+
MRj4JCahDYpCXV3v3Zvcf5EZu+QQXOJqQ8klO90ci0KWw49Va0Km3JC4iisJexI1lwx0SLAwPe/R
y4m2tomfkt1uPkh/A/c4Y+w6THE9AKbT46JDT7ieFmufj1k5wYup+OWGFEXaQOLTa379viDbwwB+
N+qJbg2uRts/RBXK/LW1LzVaxHde9ds8ez4TxPvkxJupcCQBrqS3XSmAdxOhrIzNPuZUeqWjY4t+
43hMS6kxEJS09YtLywUnrc1xPgRW/tfooQU1yDSYN4iIBAj2dvvAdPaPijVsf4mDN7qQpIihd4ZH
DcHJIF7optl9fuxt71X0NpJ3rCIj1mHbp2DGSEMYTYh7HRUS/7hr74SLIOtk+d91xtF+OG7/Pqd+
fJbQtkkPY/NoBszJHIxGFJBsjHNQaZyonNek7/nqv3Vi/zCoyiRtV1CHHZ6gzVeamdKaFPVzyhv9
SK8OU25u07AOzbfiH4qonPyQ+fxReafp0egLkdFqMkPPBTuCKiejvwUZEA5YUqr1EJ6cXooWvQCD
77v76x+Ibf5OsZilVMxp/fab4rnZXR27//mu73kRZrvCxYBIfrLbot/zQGboDzip8jjoijm+YLjP
b/XfmZu1b0xe9fDyH1XPhqFIDSgCP8uYVmIjEpWFxLkQZXgxmT0Fdqloa7Yy1p1Ktv/h3OugNjrs
Jev/YdhRhRiFiu6pCZRowZBlwf+5YqV0bWoFSvocOOfE2znhUE6MlpOXDsPgTK0tvVw4p5v+7C+r
ZWRbYxR/g4Rke6E1fxXDTS+xMaojRnampN2fs953wW3b1/ExU/sE17R9aTPcvIfujnLJ+ra7Ugou
L6P+0px3VVbZcTtnDLRqbZ5TLNaAsh9B1OmM215S0pE+Xp1gU7OBSTzl9M2JU2YTPQopw95jnPAt
3o83t4xqyJGYmJ+pZ6uk66b82F5ebfiBUK84TYLaPWic/W5AGaveWIpXdvP1a64MeZQh88RoBbzG
P3yRhHMgyU2CMmJR70mkWqxlDJGcKks9gQbzWgnAtZGyEmmTwlp6XOFLYP2SHU5min/YaS1gApA8
Xn6hWLO/Hj12dvpJjKDo/u6hOs5UDls1GXey+w8b+oQ7p2NtIUZZzAieCQmRJ8ly295OIhdAANP0
Rs8febJr4devsc+JHWFmknWpc0OoHllvy+F+usDbz5Chd7nlGPY3egoxIQrRkHIS9rcwOD4sM8P/
7KuDYQy6QTqa/7vmT6MW45J1NkqXwYIOUlaERf5zIU5AKtltJf6abyYH5l+63zF1B18pUdf4rXvQ
S2M3E/HcEuKtUMsCF/CdWv+48QWDUDbc0vAAL42J8hJvyoxWfwqCOSUJ0HQpLgPGtXiXXLJ+mUeO
Hin62j7G8QrhabxStP2xn6BB4W8uY1FM94q/HSJ3bBkQZVVAmpJauZ0vJBJpsNckkcgfmTPM7wXv
TQQI6pNJ71ZuvyJffR/EO4Pw7ZOwFVLPctvQ0Ddvf7VO9597PLOru9wSD6OAX/LAKm4puPkjLBdK
mRc+VQJa8JqddE+yZCgE2tLOkibiBCA+nUKycc0CUf8tqs1d5+HMLDN2mnwewU64WEFbC6s3UhHY
+TSaQEZcQHzb0+EHqQuNbalZ14qL+fMK6cWY644PRdxxowaDXVHpD52145MZA0WSW2tdYEZH011X
cqE2hRp/QXRtbf0WzQY0ZbSK49OAaAmzUMCdgwuH06Fr3I0bNN431jan+A3qhNJTfw9cr1pPekAj
AJjuvOchnVKiDPBsRC7/DXjcqwhyudvlLfEu7iPTB+n/yAINtWNwoeRQSx1RNacrCtXIswrVl0w9
i/Z0TEm/qEaUi3vjrwMwbWf9WYey9qJBx4Cn+1B6OQNVCHLVe0wfr9WWgDIiXWHabZNWSx0zmml1
6Fyu24ghEfT3rhy+1hoDCPQlDazN0T+Z/Rytk3GOM9rG3jtaFK9rYIAvwg33bntVBQIHAsmEIVgq
RAEDuIibl2pZX4st9e/yUDn26ob9zQK+2WSYEWWs/bBShFa2fVFXBPMXUS+b9lWbX6uoJvOlhYWp
+FPbBwQeismhUn/g+NslowodOgq4dkjKYpauYgA8UCUu3LbOtGN3JA5/ogaquINuzEF7kF99qa2/
QALEK5+qqlrYhsPQvPGCcbdvtJug/9NYuNvBKy1m7Ea+XjxRMojVOFYqghj2TheP5lrcbXKMXo7j
/968klsHiTUsuvOYroT1cSItxZD+Nik6MyDa8qJlrJSe5AEqBxROUXLhyJirm7RO0ajazc89qpbt
jUBFNKXbwSA83OgWx7p6fpYwY2efZT7F1eptxIfI1KxK8YotuBPLVbaAmqkXhEZZbrNWyeO4P2Eu
VQvtC+buuS+e+52J3hGis1doRhjmV+uBG6fMvTUaPQIE/J+EaoFcIvSkPrlEGlW8Vucr8UlnzUPM
ftiXoepSmuTmersah5qozqdxQKhd7FCaP7UMW1LA5o1yH/XgqJwgd3Lxmo3VUFeqst3bOaiw05My
S4CP53YmmZsc//knzT0bufUFrydypMCUVntw11UDJxtU2RBAR5+9z+qRXkGQ2r4n8FHVPU+iUETw
OjEYlIrAFufNdCeEjYF208fvXSrri0Bgi4vkHR6Rt/Vl9ksiumZAu58TiulL8Uf2A1QQmVP2aa8K
jOmBW8wAluGh8Gjb6HBnzLewxHbRcwowoU9afNQ3DC1hAcBXHlFOmkzizcI1r8bhmWG+n7Cw24eP
ZcTcad+CWt6+MA0KJGrfItrOc7kVQ4vzQWc038QvxC4BxwdmwNJlTtBsuAM76lu4nvKgDgXqayC3
JvKtUp4qKwsCEuRtxXC7y7P7QrYTKcOx/qtZd14PZrwfcZ6HOqkELQAMNT0VopGyy4yX7g8hzHHu
05W56YNmCn4lB7j60PdjFVzE2UTOhKXaxsECUyapEoHqIFseIub69a+gLhIQGiVL/RmiGWU5R8GE
01FBeegR5q5trdfG5C2av7x7knPT6KSoVsRqPNjoStc+HQukrYdiCKiIO/Gq81Sp8uB2YHn8MRXM
lTHZOvDUkBkzpXKhTYvPIhbWFBCe4Sya7I0dnKa97jzvzFCfzjCiLFl6vK0y/ded/gGDObgZzHK2
4pAOXAJZGMf+JgdTfdVoKrMS4MNeDoxUNn0xv/QzqtnQHFqIWytTDKQhM//Nk6cuuVtLUV0ciOoz
Dk9mGy8K3zkHdw83WrgUrno4GiTD8gBa1mIDWiPkLqDigIHnegF+GlvFZNqze9Y0/d8BVEiErIFU
XudcDQQ7Zjszwd3fDm5r+fDamKU56LDjHxMC+mSqyf92JugA6gm8/pVv7LSiUaMV0Fb7ce5knW2m
z5qE8rDtnmVYlC8bZ2F17LJGAsKjAMevBqySRzD4+0jyU0sDULPaWmTlmpgPDZ2dnPdYWu10zBTy
g51AGU3M+zRfGatFVObrAW4Z9YG4R1TJCJ1/mmr3RC9IA2LpdcKTQ6zw0TBH2Aa4KlSS/MxqUw2S
xSQaLE+KiLBfzais8TjFkU7/id0id2KCRHgYG3LVv+u6P/s9zO0Wr2PsDbMXPUuC3HMUklt9/FJZ
l5izHaxPLYoU2g/os7MpiGdr3SWtoTjeMRGzULNBCJvqNuqlIy9t6Fogkeszdp4XlBYtgrYuHBXQ
xrTm8Hf412Chs790WCQ3IKi6mHxqhunrhJ/xpF2CRIJcfSDHEdvuYhGmXG3hc7avpUf/4bmAGrCP
8+zlrwEPeeQ65fUMPNwVLEomLSiP23VfbdOJ5L5JORn5EeBX2DYLnxfejXcLWM/VopsJQLb4RJxP
AWheBW9D6QNlK28erOWwxx5a2nFbxrCNFPuFbr1e0Y6svNiqPPvvQt5jqAjjv6N8acYsurOH8jW0
JLUpzgaH4jJV6J8FqlZz09UypHlt1lU40dwqOOO2PDlIWm1+qzUlsl+w7XBdsgOnhRBs77piqrdV
I1xUxSPb8V8KJVcIY3Yf4T0EDtLPSTUeKoPMpp90cqGJuVc6Gnm2ZactIa20fPNM2iD8Jwo+M2VJ
g3/MJ2SYktOUkwoYGcolq82GceSZuoG09FPMG1oCGKv8FPhJa889T4K34OeLmzYk+z94U8OIWYpc
3pjPYGpX+2cEcLkdByLT8MdE7rAsb9DqRDuFmRAstLqGJvwZ2KA0IW0nbpkgtInf+h3DTfgzfAOU
na1oym4N9ylHsgNrLZtmIsbsY34wYy6tjv3rJhdaZtMaVFsaMdAUegi/mhaM0TCOxKcBEzFn1S4o
t1Lm6OKnMG1UtOGgFWx/lgOcHL0/wq2nPIk6vR/qDaaGg2NqhcImlAf4cqywGnPTc9x5XsPCmHkZ
r1N2uTssycbnVU+No7a/Sp7f8qWjays6mAZ2iKFjEqmyw4zsVENK/DKj51ZDe0DDtdwPmEwxeful
bp0YMOL/HbZTKYihv4PUSn4aFQqiNJgxU2NDCg+2gnR8qjXh4mt3S77zoK0zXtUIKaCK4oz2ncSW
dE/Pz++HWmZl2qgkhMjzADiQZkUXNlAeu2WcSZcfvT1pC+m+opGP2AigxRrG3sKq0SmUpsgUP8ZN
uIu1ZjfhZijQQQI4++GQ5IgrLVycjI4/n3e8XCDyZcg/1xAveM5jupJKiO1Km6BAOx4bBPtoJaFJ
z55pDWE1Sj4qyYPgUHKR6yE6y1dDgzduccAemEorwfPK2c5ajfxxhGXXiOf4cyycZL3FHrgQuB2B
sAw0TzkjQxq5PZylQVmjKiXJXG5mnk2IZYBUCK1LtmCce9pbFmIu9WTRftf54fm9OA0YtWVU/nR7
RJ7N55Sg2wInkOoL5OlxJhN6hydEDdlPszKRaexVh2buDRXOtllbknkN2tYMn1F0hu/Vuf5FNwMV
UkS19gjiuNQEz7UTd+tBiN5cb2vSOiQg0VvdRTJjN6APP0J/4waMh6R48aDtrF3p7+JYIOd4Razr
QyxPhNctg99afVJWanmJqu0XB6VkGOZaJlRHFxSchOtZsissXb1VmRyi7tilA78Ag2wM3Jk4X1Ik
M1XRsnI39up+4VjzfKaony5tkqcSi4KoXGYLLUCdbVF6sPa8I7gybKskPTG6uSCbXSNzmdMvaDWl
2vi6DllGLkZeGlm5aqe/fDmaGmn6G1IdcCCsHjZdi97HWiHU/sMuLbJv4nQ+VWwzMhTMIa5OQOFJ
og02ZbxqNjzu4nR5sFXFbKOK7ZLsDGGYbNzBkYwHgHFJDQojznJhe48AJkgHDotIcDrf5jxy1R47
I1KnnQtzjq19Fn1g2Y0G2Uw4qHH0rOPo7Yk/scuxVk/1QhmzQmO2dsWPOSrEazdGfBid0LTIUdv7
BS3czWW9Q1hwgMmz4sGUfWG8XmpsLNLE5JaFkJk3ULZBFg/Fmjc6sRLP/D50i0WQZeWg1eqx0u3K
1tx/u6FZzjAwpf0mnNZCNct0cxLHu7wKkpz7m33dGgXEl1q+9I3M5edTMgLonMCsKQPT920mRseY
OwdZUaQAJLElwGrhloA80q+BA7Q8RCGLrHAQOVeJJtwRPZHLQUz+OMi3B9A7C4wnW6P1dj0kn+WF
bwMkcxWjs14BnGOcv+IdlbghJm5FCLGaW7Pi9ynLW2SGpznrEbax2fU4XQXoSCnBdltajSJCsy9/
NZ158rQGRdD3MKnKpq/SC/CQDn0OxurXTgCohRMspCBABvTDGRk0dNeyjl7/DmqctTygFkvKAiLq
MQxKc89DSkC7K0yt/UrPZ43KaWflaYYSlGECkwJTcE1dz4oNBs1kt0dVnE2ObNPL3jo9Cls6FdA9
uQBKuNXGivWOgh3GxfLe+eHabmZ+C/rku4vso9AfWWq8uOXijt+vu1blk0+jG5jUmSpWJPtDcA6i
d5QVn8WXNFxwAB+AaYeU6Up944xn9CH9ZBBgbCyMfAGv3aVXnjngoxZma37nffNRBOEwpn3CARb5
Y1+BPtlWU+9N6+wrT2uj7ryJJzpN+ST1wFrkQ8AB6pEn/GCGdFhSh7Nr5bW3LsaJSR9aBX32ZBJv
qTS+bvU4HjxqGkBpIwovN1yZyWbK6He9GM3X6m3XuxwgSorifxU3o8VP/fMsCLGvZmXaWvPENHTa
ib1/N2Q3D81IyAdTTiDODmuS3Jex80oICD4lhqxIcXyQdncSLZLQCmxaokMOthomAlrwEV4d2Vnv
bmB4UV4CMJOJ2o/gk2PhxUa3UQNNtOPbDyoQmDB5nTzENSZ2ESzh1st3Hjm/5Mb1wbqSURi7CoWQ
0uyw6sja8IdVjGimhq4Pj8REgAJ1OAU7BoSlp4A9Sm0GKDfNNGP/eHNsz8iQu1h2F7SZaCWUD9u0
WmDrgXtBvlhX6D2oAVR8T+R+3detfhlsShyeRgPSyQnpLSb2tvSDc+24XzM3Ekd6YB2JciFjVzcn
D/mOUq3Gq9SQQIheeYG3NVSZ18sZKaoH6WWStIaCLVOy9mPADsoOKFs/rwrGrYLovbFMAog+Edfq
hpnFoVNidLTT6m9EHNylUOAb8nOOTX+krQ+9KuDckYumnGpImeP+aidZnwkSyNg2AxP6ARogRyGl
X1lB7wnF3/TvOMFLmMw2bPZR0xIp9uKWjw7MaBvUfOTvGsI1hUTxFTxtFvqH/dFMS0jJm5Awl1Cw
rbHaC75MoKcaqXGpbaKiHIm8RhVj+rRlR51BYMiTX21p6FDKH7kRXh0O5WKbjku+HJOrJOobJWdf
HFnlwzcoR2QQtS9XrjS2SBGbFLGxVlpDDqGwCVzfW4q2MCM1cH8Pd9TArcLyyuOdOBnZ6bwManmJ
87aEOJynSq76+pAt/w/S8U/+DJ9S6uzbMbqDSpTQF851vsQxmf2ufh+xGPBw0QiIBJXTHtpupe/7
+BW5CynwuErjcxlz+3lXdRjnWt+SdHciD3o1UxhKJWPNFVOACBNepQr7psAW7VMfptIkggT/awze
TI2m7tn+n7ovuCxRFRUWb5fhO/tfA9iYcq8YG1V+Fh8IhDdOxx2CWBcQID1gN/Xbxj9XT+uhrrFO
K3cL/brlQck5KWOHkzLHiIEJ/gSbM+lRJUWrrD+LrfG52ZEpaNJnqIeQF3g/tc5+UQao3iF899O2
w50bhAJjd2FGzNrqjVEqk3tYIGMXd/54GvIGPR3NbRzK+VCvVZ8Q/fXvY2E7rhUd/Ig8dn6g8JNT
URfhgzuFjhS6Lxp0AYmK0q5hQkFqcCVPo1kOmRoxmK/mAZLBK4cOi6d4bph3LCrmjKRWNHE2bRwf
32aIK+cVTl3uynVaegIutDeQsR8M6Di/iX9/i4WyPuYKI4Zj+/3iz4PR6ida/7crXTJkSnc2nnfD
vo7uO+AwQpCDvJNcughafBCi/jcvTW6vUDNMeXMzXKE/yPHgmEqApY3Vi48+B3r8CVIE+Oyuu/d2
QV9my/ZkOjhzzSoiYDMclZjvTxMe8zBFZVpNwsQAInnjFwq5j/qlwP24edaKVGW26uYT9E2ohEeO
QKLByrAbjQSFZZsdPazxKjLL9z+K5QgEsoNMfXgoHaHNEeItHDCZYu5yjO+LOgHq7O53ugsWTUFJ
08/pYlGCGFgagksZGHyXN7ryEAXPwvZsM+p+lG1tRP8bJI24yzqrhK8EfjWCLNRXv2OAMv5X76Xj
sY18ocJd2sWXFBeiMYNO9p02f9PLSQeE9RD1z+SaG8pmeTxEQXxCLrNFScli4zBRljdmX5Lg6XkF
S+a8z2hLL2a7iqz9U3nVmJVVwDC5tcb2JY9lVIW7Wi++Ea+jTQpFxR0LRzscKmSynfBsqcDUKxoq
XiViRjCHiveKwSwL+Xj+1dSmIqkLd0ZXVzAoGBWGFQegVATNijqTLNa4UuOKLEaUJjOJfRpP4CKj
QPbsegIxbh1cbxsoDfnomFY/HIVkT7XgAy5k4sAyu3pQeyKrN5EKT6fiV302ax5v9wrQWsv4AFgC
tA5O1XRWYNKFlPrxz0eSweFmEaIpsdu3DmjzVp6jAMoQAy/Scer6cXsimVZJkI1d+gIAiK+ZeOVe
0pz9bWzqxPOrMP4MEnhBEBLJ3jtYoibiQ4tQy61xJAkxFL+dVu+yR+/sRtW5cdTg58OapNZFARSS
N1IHfWO8r07v6dRGta91SSZawoxRbQgYhyw4qUN8E2YKRUSKpy8/n9OhUub+XOEAUElaN9GPhcKm
v+eYyGQSVr4w3w9ruvfj1/ZYbGxFKSHVLRKKwTBI3nYuqnX38ERkti30erhc6CITGGE2ZP7wOf55
bI4B3RCzQ0TgSRW48OudwxGKuS7fytk9tN/ByGZt4jO3JDp49x6bR36Zr0v3y8xmu+0vMC2hiMSq
HUUjvZmAMl1d1mbJaAI8Uvs2h6Yr87yztA8InPPNyf22kJAh18seCfCHaJIui7t9mCJTasYNXhYf
MrDjeNZBk0f6ZkkywzSol0wpuD/xZUu8HDjiTy9B3trykYiz6R/M++vhMvV+LG+S2zSnZ8SQvFvL
sTsrD/32QffW433UbbClUoG6d9kULjn3q0OSYjHKphCmjZTSjCxVgqmbpBUgsMPcuOxDxLGrS06m
kuZFMF++yKHJQzWHNYSKp+J+ZXEmfro2ojaxhwL1v9P+/EYvX9HiK0PkXI8K8RpF1rY8mPEv19qk
XCbdco7eevyTc1O4YrdXiwLL2a+jl1/azwIOWCz+YZ0TZ7qpCRGAZcqd05gA3D0Iw6qE/IyYcZxK
G4QPcGm2OVLp7dg7aR/wdTLkcdoRqwI+tl7RmPPKHuMvEjAcLdQ0ASklM6Uu2ENe/7k8FEMjVTp1
dvEdzw1ORbOXycbhYLcXV85MQapFYdJOb4acT87EwVrJ1rWURrux+2Ll75+4Y6wKt+kmmYQosuGO
zdOlk876AIUdbsmfKUCchU9lRqfLd3nZDKCAlcdp3DM4a6pG/mI6K5++vnCe/aAcGQ9S2rjaAW5s
vdIL2O3Lg5fr2VvcLjjFcqSxMwzcw64r+TZkxc7qJZyho/hXHHJ1HDGqlJqNbsJX8QmoLfEx6j/A
UbGNmnV+lWN+65HyWjrDGNg66Za5VawQqR08rv7V9Z0ooSMYqzmaCML41e14G9ZKwRRg0h+J5j38
9c/w7nc/9J+F3lYC5QgbKHgQHp1Ce/YK80Z4LoREDTmxAPWvTnsquLUuU3YKMNZjt0HtgOmIjHei
gdw2TXFlB/S74uNzGMZ4bSbjd8aEZmDUHoZj4a627EU5dN2AL+mZ6IZSzgzKYu/7DoPmRKQFzLWa
ztry9kGRS8MyI5dKudZlcH/OzvZMC8XHPGxJHidWrmsNlNthxfDLNN1vbYV5cP87x+mzNByr4JK6
hUSxxN3EZSvzdCFSY3OJBj16S0qg/Gl2JV3/t1M92yb+QnSapAzozQMQMTQpRNHdkUQvQTmaH8VE
Nt1pToGOykaqqVL6EuqCl08waK7lWaAcpxA8fiihUz7PJVXDkJfe9+mRXLCTx/nxVTmBaa3/VS6t
fb8dBj6uGpMNE5wwgJl/lZ6+0dvm4sWdthzqklu3dVJbAu3uaDcR1pk+GZXVh6Ue17rsaZItkEfG
wxrT+DqmyRN5tE7VToLkV9QFET8B5EAuXTyGGn+JZpqFMVH6Ox68NwEOYYwvaB15YEpL8ZbdUxDO
7bFNv5Nor8aQf2M6si/d1s1n9CUBc3ncE2OccEsWm34aP7PK4Ruk26jvap5B+S5DjTPKLid8BnCn
clw5idgYwo9L+9tRr5Bz/OIKFmNZzHVXko1Z4ua1MK/XwUV6BEC/eEcUVoLnKZ/RSJ+88AU/Zn7X
NpEcm63tEpgjYP8R5Jtp/3qY4+BHKe9Eb5D9oKu4I8fabV+7E/bOS/4NPWv+9v2u7aDEM0gXKw+g
VbSxWe3XB5z2nC3P5xVAYLtHlb2jUPjWhKCKfYm3gWGeXkZ3KGH3BNh6OCPtPZ4xBcTsQsqmAeiB
pV6WMwxRf4Q7jr8/j9UFz+JYyUyeeSuuuHM/+WrddUEgl6TM3ZhlYrTSF2pSr1butr6HexJ0+3U1
4Y6nOCCp16lEh/ubKi2E61bE+0YBcwZKKzK+oYTfaODp9hE9BoLQS0YK1gHNQf820uYbjUSUd3qr
gpVpkoKxMvvSM3gKetW1IJvVAX74SAF14kyKwojzJ/2knxcqRRr+YvSUXpDZ8pHNZ+jGuU16VquH
f3pVH+93Qp8JgkQkVGprC0sKReyTx3Z7w684e+CAkCzhvP05UnW2CUy6AfjKNLTnZ5rXTR6Mm1Tq
ijD6VhW+tOuTgwoiaDNcqNJNL/5DSm4ulnUuW+LgxsUijM3yhVStyMa6U8fG/hw4GqIsP9SMncW1
qg6FbxNupaZZ0VUPUjJvwI358XapnDK87ElYjBbLqDvYmOP2mrzIVWf+Qfg6yg8qOndCHqHtKETA
iNlq6ShWVpV0VGpadmYy2n00fVslaGuItcLwTynqECzLl9+niosIhblJAtJdQiPxmOJMjJ01nHqz
1Qg0uZ3gL7Q9xROdO8U0+70tYJYlUJQXq57Ly6S+sBJMIslehmbcziJXjYw+THHg0QZkbuApP6Zb
AF6lXhC3bfwoO+OJuLtA8ziDclg2kvvLB6UDxmgwZXLEqGVaQ5gs98jC5Qvp8fj+zaDboQgBIaMw
/CUySt2YfwTRqmxDnRSnyHYS66X+M2wxBhYCGyW7OGNyDgdQogmt/UW2dqdi2o6nemkqq7NJ+LNF
rYtcjeW3FQOKxEYTUSiyJO30+fjICV7t33E0pi8HgAqcTwHpHWr2WwplX07Uol5n2XLeEpsvdCaG
SFG2JArU4CdytYEiNJqdiBROMMqRubTca+jjivEi3krAMQow/QvT45CcK7DlSC/dyX2eydW5lPcn
DSkyc32OPfEVx+FPdhWdMw8RoJAUfvXSEh+ik+vnGvdt/eS6CZqj3FkfrI1iY2tV+Nz8oXx2RwYj
yNrSd5hKynpYmLWb/gG9rRhJLzLVdsrS5w+5MpfmAh10MqSceVX0CrbjVNEf1wSI/ybCk0cvruC1
5nd3w3DMy2BtYGeaa834LWvYZ9dRH60iqLCYZ3+jyJEywop39OIDJ3w35zIZDRwt4Bk/qZq73Idc
4Nfv4qvgxrsNwVvCG/tdQV8F/T9UNe150qP6XGj1GFeXjkF2czLoPr07FwKNW7xuArgpyjVagT9b
LU5IlIkU7teTj6hXxrTukTL1dqLj470H7oNhoie0lKBJjkLgDqYVvlA60dQ+mG+DTFIpBUnm441u
mAsWRT4JOwk+T34LzWokiGDuafT54r4BAg4ZyW7Zy8H5+Tpuqgo/n4/NFeygMV7wnK2Kyh5YHTdj
/WaiQ2yhzJ1TKPj9z0jAEWN6pvbGZUH+oIFtoGxPf1oit/Yoi4Lk85R3SjoaCr510RY2qPQKGvza
s6n5YqdgblRxhzQD6iUp820hTJvAa9K6Bv8dWAk8O/kQ5k5PXgeZrLauCMJSDBK8mWwQB37V7eAk
UG5WDJhNT1zReoozFDy0Cuf8YxJn7nRCjAL5YJhefVfiFqL+Y+tVY3Zr6rqZRe997WMeMJlJwJ2y
oEBG6i4p91DNSx0lTl80eYCoLjt34XPXNeIFgVNvqdQG2yovruAptS8Lrz9ZXMxxldrdpfAlt/FW
B0Uoh+QB4hiN4zdQVCHlbjdlCd2eYUziPZy/ZK/tRzIUV1tJOgFhCQOzQPS5EUdkGT9vkLry+yVr
ckkIo62lGtBu8PPoMjdfNbu/G8CXDM3yRTJtFWGxH0tMTK9hL4g/ZNLRSJwNabq7JiB2rqICHiC0
q+kcNOu2goWazGjeJVFdvZAapTAtj5qfXZYA4HC5xDUUVxxBgSw/qh8uxtKv3bS7SDqzPJSW3QvK
LHJy4LNrWte/59alBJa1U6OvKZe5pXoKJWY9AnSnSjZMotgSZNmaCniWHmTdjN7F2alR9VRseaa7
D4zGwLgz92/2JiUa/twYbkdzEzu5/dYt7OAeyTqXo4eOW5m55Bs4ugOaL21ws+y3Z/THP4CY9kwA
2weS7tPT164/xVwviXUY/V/o01Xno81PD2BW1761qXBv8wasrPnOuKudDvLWwfdBI4Pa3Soy+47n
HM1o3rXZ1R4/5kqVj22B0wNQjJUV5MOCIlZO1OtXm/lXUJES+ZGET2JAgBZbF20/38Eydz8CMGSN
xgVrVMVPsA4PJqgTQU/ldS8jCSqVqv9FTCa56eLvLVvpOcosm4CkruCfsMPZmoEzxDuqgr5Xdau5
N2h+kOzTNVP80Bva6e8ZtsOHsmSNbpRnYK6WUQpJF8qomzqVZEhl1oiHrCPZSeDmmPbRBOuzwIJq
fjBZ/nQTd9k4S1k/DVjLscbhN5XFo6rnW7CVM6M8PR4nmINMsHoyGeNbgXkVVC+8zGUrApFASQCZ
Llm+WhL3/SwH+nsDaEXPQ3On22vy4WMtZs7Nn1v65O9YsXchwkrQ5KcFpWKkK+6c/MyXWSB+0dqz
Y6gLU1LfkaP5mIz4VFZks7yUEaDqlluyBn/DYDpKLG2Wa11FLADzancvQa404Vf17HCNTsym0Xa8
z2eklbsGySjSwJI1NsiJP38QlxIHPxcgUToltyauVGZsYdiobrVPc8WJDJz4VofgFACD2FbO7hYe
j3jBdr6o2M+92WMkqLJudoNahqwU1wmFAUdpq5UskfuszitcrKjbsRzscoCDgO81+rZ7xNG1e3s1
frMeCcirouEsOCPAGWCQRkyhDme8PPbcN13GtHraurc3QQcr491fxOyDq/IMY1/V0RnJqrOL13Gb
lLKUowxWE7MAMVioixTfPzJJfZ6G5GGYPQbT903nVmS0VY1hX19hYqxeNusMj2ntqHjbRGsc7BZr
9ZMZK+rd3MldvL0vjDuXUPMwj7ndJ0IKgKoOPra9glQhQ5ZRj5fA10qUWjaabVn1inXfm8S+lSKY
I53hl+0OGZOfQb1QcpO257vul8HLvXVBtAIBkWsQz/s0CuO5jCabWQcarKjI+LC8/tUqwmWmIPrn
ijZEoHZF/pwF5jHfny2q+vivq7xNH9Go8yB2nvY/zcjeRSkIl/HQz83aHXXCe0t1agZ+wijzOJF0
A33VA2bW/n5+tfZxTyYRQ1SezV96Jag2dhmqoZ2A/83b+oUk/lzFzNmIoVc/ti7WdQWvR9UXnlqE
y4dPUQp8V1SEKFJDvoAxhc9JFcTRky+uBciCoZLYkRmW7oP54+/nqQE6RC5HXMesxzak+9yCKZbr
tz1eid37A/KUYAuUO6kU77W5/8XH75uHrpf0AQWY1eYuS4RbWNMK9e642dvLmGUi69FDVRHCHGvQ
FDWiEUlFp2t06fQ3pwyePhF/PJHFZucI+hNmaJeXNdTyfRHuj5leySeH6GzeZLKSOT6kMoASJiV5
LeegL/OXXKzIcYOQZXv7xMqAP/Yl4QTIiue05MVv2BU69fHyWla3LJut+35zKLNzAT/ZsoL9ORiM
bsDZz7FnHOHjVEMaedOJj1NnmFEhgrAIB9tAwAoA7jtNVa9PfBE4/gLkQR+9kJJffqhki+bKl8kY
rWkW5iCSmqRJoplSgaVLtb+NtPCtzD4W+cSFmvOEhd+bm5VguWhb/r3Pg9uDGH9WS7Hh9qRp0G5o
1LoDtQyogB+02sSrz0CxMqdkP1F/WRNYijpBGYdUR5LGw+VZ3Cv0Faa9GYZB5KmGMfk6i7RWO94z
2piUHAZZjgVKRXTkglllbigFpaWd7e/KzbZiHHbeBzfHbC6Olp2C8C0lXe/c+E7AWLs+W0hbuEcx
s9rbyTXa04LRwOvvQaruKhK17L0Ae73gPjPrSg34MfyYL+8mRhnB0/wCG/J2tfChaSI4W5eYNpys
psTlfl5tpvFU3t0pRP442Pwn4gnMg9UcJLWowhoqUxaZ267WYJHKmyVIpJ1geziHYa8CMBVgiX8D
Dw/pz81Ei1nIx9UcgUFmE7rwf98fSnoGx0p4OJmzddtrIRmG6Ufc45aScVq20dhsXIoYupIANr4t
ptk10XP91EFZOTxENkjqZLDac56kLS/+ql961YPi5j5+scJXKjj2HGngRZimJwtqTLTSgHcPfw9E
dB0+fQZ6DnsNF0kED5DLpHTTCfOAfQ9nhxWt8vMM2+Z6mbumzUa4dNpNHxqDSXsUBuk00uiqgneO
0pP/hhizaIG4spyhnL6jRJjP4I+WKfu/zTfbFxFhAuV9FKtcA+PvbSaQxZiRaGGe8h0Xv0Tgkr9f
EGDgd45E4/lsACcTw8misiFbxEz5i5Y4nZc+ea5Hg40iRnfPrDEk6a0CmuVqiyJ2s+DZtL+pyKm9
nPVU5SiZ4ReoFc001/Mo6bsjNzpFDQAkYcuAhObnGryamCE7bppXhisSg60qracN+Sf1IVswX6H/
TA5k+QHUMRmpExWLO29sltDnvFLBdyqhIvQvewZAK+6bTVXKhHBFgJak/Z/vNlooRRZ4ouzJAY3p
TRqdVh5nOhyyDsc83AsAMmCqUmjXv0C+UTmmQ8METhUp0/XNVM/cTk/Rinsj6AIPg+L9JZaAhmEB
vqe8QGlo6+R/DWGYkfBope/Vp+jh5t4Hkbghm/+ZI3GdwHP9HPyeYnZcg1h9pUK2D1vklOhXt7vW
EpyqjvqrBrsfAHGx2dfuPoFKeTeCH8b1Ykqped8Y14HTCbXOs5t7YdV/EinnS2TDlRwTSoiyYkUJ
fDeVLB12oievSCzNfAf6XPxe3yEndyh0SwsBlg9T8EUdgKJXFYzTopIxX5W9bm7kuXQOdGw0YoaW
PrPoPoOpDYdUcvQVz44b3psK0eRZ8Jr2Vdnetkd8w+5Usj6w1Yun8bA3W6lDWHPbM64XF/rAc2EX
IMOfl0TMQBleJIhu0IN1ORWnRwIgSobrf8ivNxQuDofBXhmvCk+DgTftdJHzqDfrm47wKzIEe2nC
nzrDh1J+Cj61Mf4ODcjDM6ZCE8PvABLb61XeAkCvNA5iFswYVX5VXYwY0uyMMQZyErNOLx95pzb4
qevv+LSSCIx//xpQ+xnSPOW46n18u+jJfpURxub6W1CdmJMwzboMVwEXWJ/8UbQyg6B1YkdTGl3l
ZwTmgtB9xqCclm1OvvbMkoD2ai+f64OBuL8SafemCDlqnKyu7fbYLBluWV7wSSh5u7CKZAF8VhvC
O0o7g8IM9CO2VIh9o85OM76MoXFhJU9/AjWPj7/sbNh7+wVGeZpz6jhjjuzwyzP9RP/asUSRsK2M
nRjRH4UsQKnLmuT83LCsXADwvxG9bXmtOh3WKm+7A2O/5ZYIWQ6SZO9j+G8plcHUIBj0stgLGM0l
kx0qKjVN9xO3mbtSQ5fSp6DTsOw0SIwcq6Dy3tGGxxRTScNAylOBDFBj2FDDW6dBkTFpPgxiN8Gi
AfzpdC6nKSWpThqNBC7yHr6QcXATy/WKboEGKPhA3BQzTctmZbufbf/BrOa1Lnedv9bI9UqaBvb6
+Fdx0aKO4yXBBX48ogxPm+V24Eg94f+88SSwOjGf4pmNglq7/6Iu/+TDQ4W7FBSm4WYDrezqgYzv
Q51BWQPXkwQOWJXgmGtiPwMuE4Sxg0ZwdSoeZmbu4y9xawD7XHBtRXMOpP8x6EzuobVD301Kq8ae
ktHJGO3zqxwwvHrQ+96P/D+Uf1GrwXTvKX/CAbqMJfwpDKN8+1DE5kumYYZJzmc4xd1Y1O9FAeCb
tnb9yEaOZaLFwjtjG+T/slKKpw1A9zdXZNANWUdFdhfTCGCwB1YzumPF00HvBTO0ulFQCc6EgyDn
BsWmqO9qwUMOiakVQQfcTRLIoCkp12S6G6JKqHflFrumSiYX6SQuHH1ciwxiA9DBfWJ9xkd5XFzC
PBMPLghE6Emz0Xy4oAwz4Np+Sj8MZls+o9zOMYCkIjX6Mtw7pzcOS8GC52JIfKpXQn1dc0feOV6V
uuz5tzAqJEo0uEAuSiW+KtN0OW0SdBjz4tMy8oNBUmmtWHR0Me/L/mgw2BcWAwJtIPM099E4caju
nWZc5WdRM+m9GHRqKq7GhlpTdvyaS/JJEDE0lflUD5lZUMNMkfMq3YvJv65JmN2UjR97ea8k9H5b
v6jvDbvwifVjzV5ZlNfX9ACf44rh/U9mXX+YUAtarywTmNMShtu4sYaiV3ukbI74FX8Ju+GQVPmn
kxKxg9mVJX7HChq3f02E5ElH7tteRyfSrPou92EGB9Nv0PypYjLPIDPz8Y7L7egdOt6ROpv+6QjT
ri1Yz6qz+ddLKs09xMD7GbUx6o0/+UHN2WZE/aRSHh9VR9kpVDeYyiDjw6z3kPKT6XuB3R0ZwK6W
IfZPNHXBZgGF9CLg3Y71eSZjtrX02b7nm571Fqd2DjJgR2sHykJwDz/VLK3hXp1G7IsdNnJvKbB3
r6cs1ZpzHyOle/sSoVgW94fSVeSFQ8WWUlcuf9tVdPI2gauiUj81KlujMHB0KEFYnWfhmnsS1Fbx
F0wuM/BR9lYUudDXBVQiXlUl1PM+d+VrQWCheEZptBMd1G9UD8z83QryfVmtnKKhSVtMfAQ+Qmjq
tCJfZE2mKBO8TXTojxH56Y5NIr6sVZwW2QIESj9z476W6cSgJD+hEkbYnc30eIJfYPDQzFdtZalS
F0j/4FUFDZywx9Ib3WL+xpOpa93GJVPtXBao3D3zVeywfjh5/2OnNFCGLgZI8k2WZYPfXGe5oGCL
HrDDw18wHwXAM/tx7Hjx59sJI5gM18SvuK+2d2E4FIPvkghLhhVDPHQD7g1Pgi8KUUvkcPYa29Fa
fKy74wm4D4OqA4Gu/GfZ2KUpleIFZi0dTBGgT0BrkeNG2egCQxeFjR+CcKSOnNbuYcje+0b2lTs6
jG6yTeQwGRJrC3Lif9gFrTsI7BJMm4rW0N+oeRH0V8TXOaclzAqO5QNAvTTrzEvhG/hIwhyvdNTt
s1J9e8m1yNERmC8zOw0jBS80oId2jMG0TocJb2l8XIXsWe/H7roOugpSE0/VY2wo8gL43qu6nq58
NAzargbuHlkCh9TozglUIg+cCM4HMN9kxVERTBaf3trHGJmZN6IwuZ2mvz5pvSmpxhE0FXikzg9M
eqlc3YOUGFlnPGz5QlkWHYxMcwr6MBzaz/dLrVFS+IIsZeX6d0+rmD5AjDhANtzaOpPNu41aJVQB
a6lkVeGwfoT2Hm3Zkh05JlA5X1H5OwbLv9N7qvT7Zub43D32sUippxcT7MOHUZjye+CdEphqFm9B
yeZOYM+iLliODyC6fMHou4QT3njnP0V+eDDYW+Wc58IRN9kYAX0edFTTf1zH8Jz1qCnvNr7TMHD2
NbY/DUZTJ90RrM2rbYmTRLq+t/gH+MGekI6Syf3nU+zCcjd7ny5848kc52Z7gmxwXw7uSsS3bfFt
W1TCfQ2G9d+Wm3A9GGAlRcaP5wXJuSpywXL1v7ZmOqNG/N3Lw4IIIdDtqnm0sOZZuZvzupt6zX7N
3VZEUfy49MMsosVcAZw5nQtPsOp+B1LK9qPcAADVqvkjg9DfUkHnsA6P4oWr0u5avdUL+IJKj5rM
9v4Gv2LNFUYhR5D8Yxai5NbWd/r/kGQGXbjgCY8+y6Z81lOBiQqLr/WLqwom4tTF5jq/jYZh1viZ
SB35BoE22qnixSSoKijYAMDGHmVUezv0JtwzeANLX6/8sV/TFASiKqCRbcWRk0ysJBjBvnAS2NJI
19WmSrjGXy6YxvRBWDWQFELFhfVpmoDVQs/2rYchxyvcdRTvx355XUZptn95TREeMuHdEC652AG8
QOSr0WaWEawrAIlu4bTJoSwhGSv5EBsx3WgdpcQOoxMgstMfZ8Uvz5sMhSXxuNYISkDjhEQCO7yD
k2+ZGIlhNWkpvu047KMJ0rFx2MXbe70hjLcA61WRtH0rQaavLxAH0/VkDBYaYOrPss4wUO7OeaYy
kkibGi2VwrzOZbWXeAxJDkCiyacTx9+mzvUmHRPfs271hO/oLjue1S6L7wfcuUCtWvX+tyCu1XRo
98IS76o2u1SfktNORThklcSLNgpm6lijfouMQhEgshXYyPV/npOb1dRWpbqP+j6YBIkuj+Er800o
VVudbYRihBlkunotTlSVaOyWpbS127ykMBY2BYknTOVqnsOJcOI59lmqgwdDTKXniP/p1Jr4pmCQ
XSZnetizulJ5c4WX3rIs5gV84B2t1UIUFbOkhqFqUztVansm8Q5C7GeysrROWj7GKzvYY5krhKV4
RaZMS9HvvPDNSboR7fhOYIPT/QG8Z389xiK2HN/9XyONstvqxWLKvWu+uunD99Z41sl8tRGv6ZmG
Q9UdRu3lxjGWgHc+1yz/cvsy1e07petkKj+HCefUibIi9rYXVb4ulWMOy9FIOPoP3xR6RK4pXjUm
CGM1E38s+aP3/9MbJjmjBwIY2X18qdrPdcG4sRs3e1XUbGa044I+VFBLHDqKiQKFInfw6qPrysx9
L7hB5wD0RO/kGp7pia+PReFiOqjhHW2q6dh0MN1ncv12S/rh+sqT/szcSGTxy0PJF90h1xT28JMu
5hG5QSGG9M6Ep7rWKXbEpbh4grn92IwDArQrPjJaUVCuM6BD3CopKpgP+EhPaE3jEXY/5JZbraE3
9QNSGe9IO5WP9Nxx8sxW71CKP0DuxghaxpSgRwKJ/iqjILMYjo9/vwcmgagD9tzyxmirzHSG+YRx
4QAiKPGFjWLbOv1zfcuOUxRFGl3Lp5ivebGAaUpAmBEvCedqay/r31dQ6WHMLvzHhPaXYLZgJNA0
neMeTQolLwnsANo6RQsSjmDtkoTCZaUOhMBRLdNCHDCtle1gLmfqA8PuDr3gSil8FhERDnwSRjss
kUDV1GxuyOVNiTeCVLreslcIGmo91/2VbN9KghciwNkkaUa4S4odFi+7stzgfXFJtLPzS3xCC3eh
An5Nf2+cj4cvnHM9eCUqPnNDQzDdL7KffuHEhtsh9TpUiKeE88/mry97Z/QQ0kN5WqFBxdBAjfxs
wHCbc3NoUGFOH7r/S3Q26r3L1wNEEtLauhXxl1ulvnqcZOCtSs8Dhi1XnGZ1rxM0ygE7AoE5h4fn
izmJmX6Y4Hoo8cgwv4AD/baeUeAJNSO0MEss1v35Jz9TRiHcCqUHuDCe1o0cXFoouRVhQpARmXTY
CpaxhUEcF1l5rqeUv0z9s1YOymYDXfE7MTdqQoa9hm9kY1s1zA7E4rtWWt95wyudYHOtZLN+2+8P
Kd1ew1GpslwKnbqMmQYlGhWD7TCINPx0lsxuneG/AIfqk5JC/b6qsNTmYVRsOMyRO58cDu0PMuGm
0J4pmqfl/gTdnBR82cH4CP/dotjOv+eYHyS88z6F+KMo7cbAfB1jXUB/qxF1Haa/y5RY5Ecm1LxL
CMUIBCVasmdNlY0W7wAAnUXGlKZsYK3crczbauIu6lim4VZi9YzaiwG/iVV8/rqOTgIuQfAo0EdZ
XZzk/ERWwsAffDRBW9yOajhgrRlEv62B54bka6/dQs+C6t2lD0eadValG3R58P7G7pOVuHvUrLlL
e4Fiez0G9T/BpoKhemFnC0MpmT8E/bInhUDFjQnl9T1GOCINo6xrLIS0dhktJsT3hdLiFdU7VjBR
jYIL60NZOMb3WJUxVnpDl9JLwkx6YsYM17943s9iVHSCnTskqACCJgZf4RyXG7aCz0gCnaspENc4
HxWrzQ+4A32hmhu00dgNXw2mIWtJ4IIkkt03CU2OOIPY7rHe+C7YSwA4h2ceQmTErRF67dux9274
N3t1MJC800CQIrAQeD1dETSqb5mXgFpAu2cALLRRo6du4PakN/z134K1Jz0XZhrtO9YO5CTUw2Ce
CeB6WbFTJSgBRikhc46+jwvndELTWUbQIsN1rnuMeA99vYWr8al5HOeJ2EO1RK/hW58QRm0D7+vJ
d7ICQTpQJu+2aWZyjSI1+iFIEppY8VJ9RpZnBJAsHWW7ojvgjN8h/zjHQkDUvGSl4U5yDDGzPs2P
GrsxYumyqvppQ8qSzJMTJazCzpzpnl6J5K0fRuFrYGSkyZHgQwrITJQlKgM7dQs/s1CUWeC3evB2
/Nh6ScgsVUyv0ior0vtNrp8eG5ivS5OVzNq9Zfu1IUI5ZNWxBDOc6H2v1uTrkZh+As+GwLRTwsfJ
1UQ+F/WH3dkF7SBR8qx98YwsQOMFOumQuPquh49a+notEvgATZGceQKKlvsEN4Wxwf0GhKNhEahv
iIINIMpJaHLhWKvqbt01cxFyANQN/Ymq0fWkgjbH/xzLwRYalH9/Mmy2EPEDH2idVQ4Cwvkfpqnd
WINggDR9dFwxF3VRByoQou4xJB88WdYy4oEg9VX2IftnW4u+5C1cLQyYvUkJjxEMQUp3QX8FEKYY
/JIx5wfLAPCNg5miFaHQqUWW7jB5uUVKic0GWuSkvyTH0X9bqCJUaGHViMhxnuLDcc8iD/hd0x53
dsdamUzgq1XHJsppyUSFa1wTvn7dHJatCsx25vLa6QLYMMJbZfvNaGo4BRP82+gEeoMxvuu4cZl8
eqFf4RoVWYhLnMXiuJV94CQSYeDUcXVv/eE03jsR2cTU2j6MtAsSMB3/wp7B+O1D6o5KApU9K3yC
Coxk9mruzx/d5zHkYLnWnfvT97BqRpd0QfTRsr9PdzTswTzZdIQQSYX5UgkjKIdpB56SAFxDKnHR
V59z5qICelGVsOAb6a9yATmyw5PnTNfJ/i2J5swB6ZLXvARjwywv8S7oZKV0FVs621iIKHglfCdl
XJ5575p9kiEQRRwI02yNEYoPw21pK1F6UMZlAz3SqrwiFbTtgX2Wa/Aub9pVY/6FbP9z8ziLc34W
KElkiBAzE5qmCnUkVtvVBuv6gKVsrWdj1h/rSld6qxI3kLnlPVDfGmhfxz+AEJ4sMDYwA7ZG4yoc
xhWB5HsyGlXavAwKapCpGaOi33IrTn4e5XIeKTOnAsAqmdgAhCbkYWslPeblECPjYshG4KcT96HG
PTezamDDt5PhgmexBeTVZa7+gFLKFLK9SvPNMhl067g2RSkJcGHFMpXWz84iQkcYibQufqp8d/a/
t15JmFXwgX9cUvcFdVI4jnETFgjU5huGDycV0nHXmlNQALEE2EIEWvlwPAOyVarDbMWrESEelqcz
//hjgTv2LiftspZdzb4FRyB0BfH/ZIG5KV/t3+LR5bJomuhueGlGauFiZrPfJzLj+Tp3GgS4Sv0A
Wh4Qdb9sWRMTF9xjMHdy56L5KMM6I+ssBFLD7E31BQfwAskrEj83JUQjK9d/sROhgZI6vYPO3Iaj
7diOthkQJTvUMzHiG6qOLxek8RKV+EX4XEkwxGvSZNeBL/zJrLSv8ERd5e1C9Nv9VTxrUV5T56iw
bVLpZd7KN1ZIyGubX7KYuz2rM/ARwMQTaLXHpfl+muW/VFdcNzmHy//QZ2/Zm+tRUgP5VG1GLzNG
+1qBiTFr3oMpm+DS0h+uuf/7yxfBZvxWcMAnR/FAGdpz2KrJUpPbVCItDXWRLHorS/j42/RlgLqo
lVjinkWWQnD5Wsa4IYwNhpBdDMA35MUYIwiqvwRCyt2+UGYtiqaYSEwCvUIDFAOuM0dwaXqUEzHM
FDCgKCtgULmuomR6k9VdeCuRRVyLiTTb1yH+Mnlr16ljRER9Jm/RrjEdgzscbpFRc0i9BY3j7w0v
SC33IWga06bNmt9PFYp4rBXPDLYXzTyPDJUyViJWsoMG+aHASa7b7VM07/3qNArNJIKfRcCU4ORm
+arvQoDaxFBU5xjP9TasIvlFqSdgs8+T1xT/n/n9Wm2O2QPZVq1iOlswXJGIiEepJNhU2Qhfo91V
SE99xGBaubZqHzrJlmwRkjfnELsA04UkaXX0YGbaRskscnfGXaSEj4Yw+6p1RhdjZJGXOSjLuSx9
3wFZkLtIHhEvncc5zVzr+u73UO9cW5nnYGhc9vnBrlq8ED4w2hJsLUp0YQ/GPCCNpCnt5T7huLRF
HVt51mUJNJH6hELS+5t1y1+soSkYxTF/tuh/evBSYgl8OhSYQ3WASJP2KoDvSoHsmHMx2skqZzMR
KR+xDdSn+xtrlcZN8kAXrPlkAq9gfLG+asrop2yh9PfSEsX3cFASX6/mvmvgtLvNW71DHxWj1Ip5
Xx4+CPKkOISXTnpQqPbr5iPcB463L6oo4nqnYbGlKxTm1D9gGPinzAo0Sr0Uhy9KPi3kFmOkHLnT
eoP/N9LC1lJUGg0F6issMw7sTEfZGELjJYU2p8i04CvkmMPUjyaWvorQwiyzvwn3CDse5B/O9AjB
wCIYqV+w58aWX6eVS3scwIezvR60wK11uAH/1a/s1iOj6tXYlaFQafYO90mhrKyLtB5Op/d2/IVU
hJB6chsxKcgGYitk51DSNxC9n6zDMW60tpS9fWNKBaVwBkM0AKHw2ye5yAiRmYremCbNX6abhE8l
PSjf8HVZiggTAUca0HCURT0zYH6epTISBT/czG2BGbK0pd/kNR/YiKt2DZJyWh8N+XkRWihvYrFj
EqNC2FZ7i0svyDKkQI29N0tY/ifB5HhuRQxIwpI5UtuIYe7f6OQTScTi7FcSJj8QsANJJ5CWwQn2
EEmqUk/W3VK2LPtT0j5oSmLcjQbb9X65eJD8NQjOHSYCQk+u3+BbNT8KtcqGL3s5eIe0WVoa7Sla
07/s36d4bFB5A+3AzgJ9leCzJ8iwDpG5fZ1mN+H1hvHAbHKOtphTL2wqG6tHi15E9/h0xqsdW3qY
4VBgzYX1X1ECd7rDyu/Hloaq2W6paJzKqtWpYdqjIo6Am/cN54inVHpCUK7eTxWz22x9jfUMi33K
LT1hjUHXzGjJSIYhPGuQ8FHFC3saMb5cRUJPkCZ986i3IhjfeWRW0A6jHDqL4McsrPkEiNiFFnr3
zN4GfeePolZn9R/laQwI/6Q8XGzmYuBgL3p6geJC3TNI59HoqSZkLSzP03lFcnhIIvXLhxSUirqk
KNI+BevkRPV5HDdt7M3XQLvIFODceSW/pST9Wsty9OVi4s3KkhDItGwspOfCryPpv3SlS0ihB2v7
OJkom0GRAUgPKKdwLpwsgI54PAB4bK7dtmb4znBTILo0mx1axdvaQeBIWyZHcvPxbaFx60aJbNjd
HmF+Zzl7KkQOj8Wz2zKCrgZI4FJLGTASI4aUsbFsTRCXgoOX+8ElqKIkQaHTrfzakBsM+guAafC/
lEbKE8mNVEliTHffGUoTpUBEKfE6LO+wQSZA46rir0LRwGY6NtRnH2KP+Vv2FLl3Gy7N0GGjdAlt
D1/TEf8O2jQGqKOMiV9hvC8K+0Z0P9FP9OKybfPBirhsrVw0Ql//zB2tHasirmSKhWT7MPdR3Bwl
ftwDeza2EcAX/dkso/vwmm+Cmwd3WjRHwaDp6jbxbTaFHJXLkB+uqDq8LHofqigelMNl2dh5ae6n
lGF3zoy4cXxibb+4vP7KCYGZzj1V5GPh5/gNbymT53F5nvNhsloVlHZ22/F8DlpEHZNFvKcqHU5G
egmNkOJ8G4Q3EsEEAM6E1jBdo7bUdYPzryN66GGcE5uRmG9Lld1t+5fU91mABV6IbaKztasQj+QX
IH4mPFGu64uTP2qiYPLAiEKYD3FZWbiyKo7evownrF+u2Ir4M9C0iKst+QC6hGoHCfvoGXJz3EqP
bU3Yx5yX0mNFasxa1AUemKHlwXepjuBcaIa/wVrqmoYIU+Vyhw/NvCPUd8al03Bwqt0rrMwKnzor
ntQVeVtLfvGai72tPxn2K3aWpDtHj/f6MBKmg6UOEmcT9lCnvqkMm1XHJDoSO40O2+E6wYtmQt4E
d6RowefIV7iI4ymog6Xv510ubZJkAT6xjHlanOEccoCskNwK0/dZIPxriaP3q785+kG0Lw9uu9Ys
PWaOY0CMF+CgiZDzJGsVjUZsvl8XUSju1YOMSN4R1uoHPSNAVwf/JWEAYhlaq088n7vHzdcTXW4l
YaB1H+Uwn8yCZRDzkml1UtcAcTALpECLjepDF/Ky3JQeyuKlJN5YTaxWDd4/QQjePx9iV8IDr15t
o00IOjfZ1Hwb/LKbHjDkdlSJee6qV4kQiZtKDZcgczzj9ziUjYUaTQ7uFvqhqO+KI2BaDolF8bQq
JSknu5Zq2FMTCT4RVdDaaapwiVcebK9R75fdWrbEfUrMiU3eRBzCxcjv2UPEtXdTTMICa/T4l7Gs
GWtCGGj7f2xGTmZs5V0PtrIhXOPGeQiyL7xJEkQQcBNUBEUqLwCCxgBoTiAHrw6b3IxYNq5SVgUT
igj5cgS8WDIB6kzsiMe8pe4E+c2qoLHIxIQbVL/LSpgUlhWx9WsV6hvWC2XqiwQmD5aClqNOccrr
0ce/3al0CUk8d50MoOWDD+B62Inrd33CRtme316FeL7SuOihj1iO6tSVEWt86rkxTtt8VPE4/HeG
yVBxek7yDcSQpUzDzR7kxIm3yz+rUjgyRFExpEFE6Emb+RNsb0ol5D+iYAwprw0al/+qOxxDjeny
NwcgcozyX/ff2sWXCkhC4h8L+SM4/+aCN5G1w2mBfCCn5tfuKqmNL+X8DL4/JTf2Wg4hk+ryhHUY
dUXXSW22J/A//kmEwIrCVFxwDC3xled3EZ2P82cpUUzY85LdNN4kWJT0/8RccSprjvzFcqPrtOo+
tunC3szYTZpP5l7jigZtvAjh3pTwzx8yWs/A1RWdC2gotKyB2j4UrkHvCquLfLeLfIs41LYonQ+v
9YExLcWwq6b8pIiPkmA//vTAk36QoujwKnruxAg8dgWB9Qf21/aaKCjoTtH+t3TMrq7Xt1/2pJ8X
qyIAujFzq2lA+KI8aPA0wqZs7jDc2wXH6x9vqgXzEMeg040FV7pIWAYTGFG5cFzqXXEa9Mi+pKXy
fPXbGnDFGBhHracPdhNVCKRia5k2y7hqhzXQZKsINMYSlkYHdb5vjSC5102MUYmKf0SHesO9N0RC
ufuwWSEvfABvTTElsMzOfxbRF0SSuoT8ckV1LpXI+maJw1uD+x1DMsVEgt5NwA8y6tzkP9/6es6W
42EYONNNiBJK8OsYTZmLgnAJF1P6LEe4OKoiqq6z4R4fJjayWFwyYt+7ZI4VS1KJ81tX4XLXFUsC
yXMndkWSAr5Q+A4tHAOkpWRIuXptSfcd3o0oni8nDIxlzR4/e3NnhON1zjoHwNfdTN7wbYWieJYN
NL+oyQiiJ9v8INnw+cDJSjoP0Csev1YFYy32ko2yCGioDc4yxFZRwIzz8atnxPtjS8G0jgaxH0yT
S23EXXuC1Erx9FfmYAAg4p1WAgs7mk7Mphh97hR0lyYW3YlcBDBUtYXw9X/l3X3jxLHBmUzdKWVG
U+oh2Mivu5/BBpXOKLocZR9i1wFnciVOVSxQ3H4JdyzbZb0OnJ8zQKXaBmkLjhirLdma0Ghc4KeA
UT1RBrI8jrKkw0iRoN7YsuqqNLf1tIQU8L7QaBiwNHBSi3y9S2yD+DuIWh96hoF02RgtDCJ0hxVH
BCI+YVrjzvAdX4JuXvRCODDPnkZ55Q++JrN7vnLbhG4TPdDs74bNKLrLoSSV5ay43SO39D1ovti1
nrlMXRIZEDtWtAwQuYWf9EEj9Mw9HcQKupv0xuSZ85VTGWHwSahDSvAV7chhGGyc/ZRUddXYY/YN
iZ0mgEQs2qSIfY6Y0gxHKU1+w8qHEAG15di7MvLnktlFDDvaryxL/HdA1d1o/NSjsh5TVNNv8bXs
JJGlD/tCi7JP9pedha7Tfb3s18wI2cqbVaxXMC1IvBn+2Dc7SVCv/zdkP4lE1itCNK4ostr7gXK9
ewhiWUjAW/bdPaLrrx95LOsorJVlQ2VYMMqld0ZpzMGedDwzvSK1HC3V6Z5w0LVEWLvuDJUCHz+w
Ls6Rcn9SdeX/4rTGwNiqkma2OESBebN7/irG29l4rQ4VdNrYUbtpUuIf4hVCKDgjxzDTVOqSMr41
9A2yDzylmVMnMTFK37Q7GLmasehQ5JzFRu1Sh5Fm+VxiBZ7+QAwOxfzYxqtCd7v0BjNUPsUygVeN
K3OOgxEkAMzA7N0jVkV0zgsm6KM85U09mOytP44bBytpL1/wxxUZqdgITKXE+FpqSkIO7i5coG0I
q6KyCVrSXGOr87gf7SY1DAwEl/UvUyJmYRkAcfDlHC225LWh1B+4F1w9/6Tg4M75V5M4a2qVuWTc
jIGRxitif1xwTJn3E1KgIVdsUTimRtU6WQnlWs7b8RgPI/t3UU26DfX9ALCtKERdy4UORExaKJEp
tRXiOHwBcBQ22OC/8xU5T2TIlo8KVEmYsPRClgWq1z8W0E5E1qZbyD6vyBX0HFXJNdPT+jZkwk9r
TP/ES5VFlSIQ91Z+eY8VlLsNTHaIXda017H6Euru3h0Z9TBSdq7gvp56MmM7JIoInRafRtbbg1QE
cmbgggJqzfLVARxEpS1NpQlS3NgPXBiM+MCRgU4XSzkookgqjAbnYiLLW8illGoDhVtTkY6JibEa
ZPCddUEPgXU+q2paJK8AIfgLNEAUdBr3PfhX6a+URnshjW+EJomvqX97btvdsnpRWlrqpmt2cJXh
nur4A26pnYXE19VJxsUBp9YSwU5me4yvxgLEDKs4Ft8yktWpDD7uGOWFodWyCBr1EuiEslFkz4uw
/fBrOjudIieLqlJR03Kq/FEaXo4ZaYEtKymv962rIsfAERx/cUFKPqJ9FXj+wvh80Lx2Fkp6k0Fb
Tniw1OpB19HCR519Io5ipLrw6sMbmfuM9VSSVnOnOfALGDs4LGndKFIfLr/M5qzWnt7GMvcoy1UZ
D7qgcSSDq13+iz0k2tv8U5FMc+vxrdI6uCca95j1bY84X5QnDYVhTHuoPcyNh/G3RV/BWcAAhXT3
/DyzE4kiWCYWxa8lmkWGdKYVDvTW51ScQjT/aY8hA5mzXQ2G1CQ4P0vRbDxhwV5Qejk5HC0V2f0f
C8yt1+usZA/v8exyeW/fkSma9HkIiTHTl4xf0ewTPxKY/K7lB83XbLxBI8emX6rUoAOYKfCqTZp4
54nSSl52Kwb+L1ife9YGo8IiCOV4yTytHpUXdypm6NYc1DKEiyu3g66YT7VrWsqdxBSm2ZkfXKUl
nLpRFDZGBCBSYFiGd0nj7e/GTShBWogyxdpCbfMspJ1oX8b1UgJKIG14RtRBM1oAh47+tOSRhyy1
cVQ2YCjsWQCCu/Dnr9ZJm0TKmuTwDBUoJtU97M7a6JYpVhLI4f1Jezgd5Cd4MfPrxrQnaf94ukBu
CdTLLtyTvoOdcLqcvzwyc934ncygl68jOuwaeYGOk1YTCmqjBzmULYzZrgvrV7CkBSgtFQU8pi3L
c1cipQYJYavJLg/VTUJ7js1RkxSc0mDQLX+YJTHsog+jfori2AMYHnB9CNyI0ktZMtxTSPmaSDxs
b7XtzTvl9hIqJ8NvjYGJr3bm/E7Dn7NlD+0Oy5+0/oY0XskAXUMCimKjkhH9K/UXr7tEMpKMPb0k
rzDOUHzze+/m1fwwYqKOlSV71r5XruysFonq2wC7rylf7IsyeWvE6PQkZrlK7iViT4tlp/FOVwFZ
eUlSglg1SsgzG/NDEx4lCDZD3iwKmc5C3zEd9haAUxGJdtGraWSSsM5BgqdAzYmhR3L9dkEXQ6fk
8Y/Pmq+jloPXIizlwhbua2La5Z6PL6rQW9L84MK0eu2astaXi4Q3DQt+FKJ27JjOAIs6YxqhQ70W
/W5kucFPrrPW1jBZK+1QZoRSfKSMS9sxDartth65HdI7ivXWeN2o9FJ/u/C8G7omiuthEjiCwl7Y
Eg84TZzEY6/SYf7xpUzlAmbPhQ6bcTo8No2P/tf0FqaymU7FY9Clyr8JuPALc6Ji4W12EU6iwxFo
dhIXyXE3QK7Agq09dBKF7AWVwxxvnYPyEL3nYIxYfz0GgW/hnYOQUfZBVyKRVBLr+MHvjuvrLb+S
etznu426WT3oyBfLcN/+fbAVQc59SbEbPz+1mHPsqhSfzA9Yixhdi9JQEnFEkbcSlFAXSVLQRgsX
oLcjFQINsgvi+NFYlm9kz0MBlBfxF8Ewe9gEqa6ECqNeWjTNPHTNdn6JWWZxyC4jMijtKYCFTYgP
gsDwFfZVdIwdBSIX9Pcr94dIiSzx6llZzD/XWuoPfD8mTGJ+9shx0KSxv7Gb3pwwZsj0vQKVAhNG
2B0IdLC8gr2NEiIo/G10u2+V9Vcu/p99h4qM0EN4OXiv7wSXgH2jVPYVUM+DSZ/L2qtUbFwiHymx
nUiOYAH5PXkPvPAEbFSa8tZvpFS0oB2XtX8MmeDqprJ9Gk1kVY9H54UoR06v7V2PlJlm/zOw5j+T
fKsYb+nh9KVRJCDEm1PWmsayLstA3236mjyH9pPC4knTwP5ki2fcvqnj90kaQjNvV5YfJCvGgDnv
AMER7hlPO4GKMgtj8xkZKkfQll5ZKXat6FRuez44jfblgAQmmzeasfb8hU8nRwf1ryG212YRgn0P
iwIxGG/Vhox15vNkKkoArQ4A8qmAk4obBPmHQuJgqN8whrzDwRnXDSQr3bVlLwYC8D654IUXYDNn
MeNDwVFgOCxt4W8vXipXYURYLZULKxmCngOa/kiWsyMKl8rPDnOIjGQfKa96GCbHgv20QqLdKfUE
aZ/wzWGYExnQGniey1a+kU6Kr/RWgsqrgOcxeiCUv0ppqbiWZQRs5J5xleiGO8OjuU6Jsjnudpia
fCdYbldDhs7ynxj5ho0WfsnzIP20/6by5AZ0678JEeVBL5KYnBJ+v56dd8gb0JbRp4cQQwc2cjv/
Sa4qi4NH4EyGAq8ctmec9fYv40vNTITJKhHEG5ihzoMkdfDJ8c5ERpTImGy+hped1n/UDjspNMrS
tP4F7Y3+JjK1F8RqycOInSBA6H3XnRX52ExfsNcSx3KTXrabAyrStNSU4J4cDQO9LAVzyngbPE3K
0AziztH1iIjXatPNjXRPsUHh+xHgNANguSNbn5CcqsmnCI/I5rjxGEsYhsmX7Tud88Tgfb1RbiBd
YvytiAhixZM1Kt1pfiSs6Pgs0uVSRYaa0AjpGaFaISccR/tArcZjNLJ9mQwt+lF2uUFin/iThRWk
LdfbbN+OjoAwbjrhE0yHjK1T0s9pZ4vpvf5PqOPNefmp/nKhGBQtlPxOTmFfFPsWoSs124nsqlOi
Lpp2Uf4EUzfLYaAIfXN8I+AcyL8FxH+1KVrPVLXQ9sMr0QNA/EXjGhKMZQAkqN5fqps2AG+seRcL
roGyr3012bY+hu0qTCLlt8/MP6BgpIKEhZ89c2jSYAKYVOuzgZbYQfg09bujetgfWIWnv3arQxyY
yKVb+jG2hZ5rv8nOnEqQMRb8mKB7KQH42tWe0gAM5gEkSTo65nLnbyTI9i/dLsCwg0VySeCDrcjd
JQimwHM8Kec46PunrWTWb0AXi1fq+gC6OlvcdhfDjBd+t9muqFyh8jcf94kiA2Muq73ZWL4H/7kN
08AD9Ct2Ibumyoi3hZvtJuCjjNgCWZed73Tb28v3JZ7TmiIM8kdO0iJjrLHLLT8tuqOQC0sHreXX
NN3e3FGSwCgVcnCWkneYwMPlO+gfQzUnpXno+pnAuIecAXjLAaAK0iOZNGtStuHAfkdh6YvtvIQ0
CAwc506fqoZxGT+3ddC1/Q+SvEUQuCqBHNW772sX2FJxDupK9Nyzw2emzEes1yGn2nk58f/4WFqV
UqTGv8U+htVzTGQItEQX2LjFQKXKRty9Ktpux7wvRax9NIZVgkCZA49vgHSTbWzhF/ao/zW2jSXW
hq3otFfRQqwvbYObQ7+h0DY1ts57z65yGNVb2yCHqE8BYVMLxwAUEfgGYEtM7T/Ha3e6FUnLafza
lZHDYo2kqFUXaiC9FjfnOhskUYI3+qxhua+0QDvWrpz/NJ8/HpS1DrO/beKgQwYdLru6gqHfrU1U
5UhP/EMDwhfAn73Qk2VJO180fYK6/1zr55QIsTdT+dp/xXeK05wL64iO2WKKxAoAymOG8gzr3YLJ
zq5zqejGub3fzXhpnk+yAdYJ0R9Wi2XjMDGvK9gxOOzR9QVvawU9ClxOLWxqgZhy7mG9CxmC8ZJL
tXZm1IuL8duElVBCJFLqgD05BjJmFHwg/BO7pVVAdWap39XZjwccPjRbcaTKWMYlLSAAfA1He1O5
X/xtdLq0DPxstKjf3bvf+cDa5wKyvFF+JR6AG+QnZL6PsGhIiA8E8J1KkhUG8thsBF1p4Tq2XRYX
T8jvNvwkqCkuhXeCcbnV4iGziD9YaOOIja5zYOQuzskp5YGQFpg3r1TXm24nNKIIyLQcPuVQ/Wum
LfHc5EE6kiC9g9qh3YNPoDiHnokRArdegpJRmVV1NIbwUogIQ1kR0RwJxXvMVd+h81DNE14FW78g
DYon3GsXpqv7q2JXOtMS+Pv1qPM4Oq2zAy8uucNjZjXGlzPCC6nJdBs54c87UUknSB8yFvdgDi5s
yhgppRfGB1QT+1e7urJqDAU6KsDNX0dhtY7lI+qMbOOY6sJaTt7Rd/0XjS8m43lNvEcxpDRC8TTD
vuj5yZa1jp/ZnHSVdH1GDS/A1R9ZzcDsUhFQGQ0jmEMJCIU/eJaX1H4sgl3a3ES+UvZ5r94zq1Kc
DYWq8JrLgr8YRBZ1ofTW0xRRh1oI456oVunv5sR9w1VrmvxxZPiuxHMEpxj3Gq0/y2x7AFhAYxg+
jn413cxwHCqowfCdtmu9jxUXyXzsPrQB2wYUTZN3cNQFvAQUNUwyTdR3PwY/1VErm9tA1pgZaPt8
n2+kqCyeWG0lqlpo1yWleD/nNY8uRh4rfEYd+6mZowjGyhf5h9kk+gFI3B6XP2FxsvV2FV3qpJ6e
je5yiniyfif75jRrmKjknJ8Mqx1ou/S+0Reh+kFagBLJYJihkOuL/GJaWgX2B0TxZkX1bj5W8Lfp
/VP36p3rMEcGpimkkRgYMG68Sp6XBKfUWF4k1AZo1h+h59TXOOsBoWINVicIs6mQVo1TX2LoTFbD
hFNA7fBDFo4D0LNXOIikotanWEN7hGwT7NbLh6pFA3pKo4h5JEMJowN3yg84ZIFSI9YEJTNKE09P
hEGUnOHA4ywgFfu26AQFTylkmqYpya/wYEK6FvV/dgeVPoCIJl9WdFGWKUOseMf/7oRUkLJiEHmU
26gN91DZ7bz9yPEwm2Fg/TPAFuGpHVnjcQ0SlMF63KRhiNLjaW75piWSKc2ygn0NtVoC8CXbNtE2
ocMoTq84FGGkF9gpMUFH/6xl11+19cPx5Cz+A2zZIXUrAVlM7V5S9Dg3b5hfOWpkoUoHRY+zPl21
zTsc1DXb+t7HWWNd/mDIxVo2r1JMzx9O8hI0h6ZGkLE2P60i+ZKBHwORviFoq5aUh6b/bRPHLfBT
2w+k0y1USp5i4R/3+GhYwwBGCL1tCoOoVYAC2z+p7IicAX2z9FZSZrHoMvRTgb+DEfNMEp27mg0E
GuCUIPSYgzgxh6rlQ3uq6xvRNsvk24sedsmuWyvIDktoYo3j4mlaWLP0jDCr7zvrnrjuFMv86yyh
Ekfh9kTy6PicJW6ZV1PiF0533pVEX5R3JBSgEv6CcXo5r4sdwM2+HylSoOMOpzaQT0vw5fJqaleX
khJxukXdPjwvHwtyD5KTP4uXHWce/p6Z+9imhr+Vlux3R7TCaYKQ+Maq0JUKJ82K/2cnioIL2P2K
UHODkNFq2BjLZACx3uEUbZcPp8v6F1PNbJoHveUmUWbU29TpziDZh/8B+fZ43dxUUAw56mwuRxmN
NSqm8l2DsNpgBXAInF1B7+AfSSql6KbhHY/pWNJ/VylshXqrQrPt+fvQ6sy0VdWa/Esd5ZUj5LGs
3JD2fEgYT4RNEWNIY8YdFv2zal9/b2zdTGT5DZiCrZ1JHmdDBtdNzz5KAMq3xvAx4bf6eQRyI0he
eQgCJtGnLEUj6rLdyaFQadg/Ug4MBTJXCCS3nRKC960nHO/3pi5ttI0xk5IrXhAzgbhfUuQ8QZ4L
yc8KQ4HMNHp1AgqbJoM3gmImqFjN8xOOgvqDAZ41DGd7YG6DvmtdgVMoQyIc4A4RKoTOx5uFKzgM
rC/8du3UqnWTkNy8kxmdxtCPJSINiunEcnpYKi+Uf+INH8FM9JUKLuJ85Q/hXbqgjKf2okFeG5Fp
Ye3swTKMZr6MbgxwA1Af3c8tMUMpQvIHHQzsu1KyUKc3Yv+eEjqSWPZN01DnLqoXDvnDkMw7sTXM
UdzsCNhkGz+cJgkspizGw7MaiX4cqCENti9ZMgalJIfS1tF2vCo36tBaiX7Nub+1ENoUKomrluzK
SnFm/5KgY0Y+vheXTW4KDLn9B8Dsv9S3kiHK2EiqDoMNaKtGAOuS28OghNbTi+BYvniWIfZprMcE
Rc/z5uvdpk6KLdO2YDjvwPG9lPtA2zycdpiSPHl/KJ/PrgVMi1yl2U9qRy+ncdjvK/XlQ4LxOFj9
jGzVRqFx4hXQ6Mk9qEjQ0Ani3oDCYcDRCoEv4t+ErtKMLF1n3dB1iSubou2TI3x2iCYFRnXHrnUe
wVfCzFB4JiXYKopJ+TQ0WDVD0ZDMYv5dYzIGN/Irpq35651EylB7M3oCmykWKoHTOgdEVczM7NSe
yw4UzcMtl8cFOigdQ7Wwfx15g/UsA01rMJbOBVmB+3nap5hhxIhawc+AMYENIyOX1vvKZe1qsHf/
yJdfm5JaiBTrTP5bPJQmJsLl6LbeXQd07Ld43K3R1mQyS6vvnLMSWzZBkZa9DPmFQ+pxYpPMSlFh
Yokmz3L7rq2AAnr54OyMZvIRD0jBxDIxWrH2oSZdqSELH75Mki5I0qpQhM1mYG7th9uHSjqLQ0Ci
jo0wrqI/ZgOxVHa8DwBqWNZibzkUreMk5MBdmzhPobT91c6hTYfAfaMSzXt/ca0yWtOOF0DlypZo
9BwGwXzYaC+yeosVNJtYLZcSY2bjk/A4H+/i4KbIUDPZ5f/38SbMl+JezQ+R1OQxrluz6lSKR6aN
gYFNRVttouLJyBZrfkpkoo0hSh3lXSinfkbX5J/ha+ql39wsLLWDbICwY7jHDKqlq98KjljDmY06
90b/9pQg04UJ+luU8/9TvRkI5GhuqtxfkzBYte40JS25Y9XbebkRv6EEYtB5F32EDiBVFb7MY2w8
23ZZcexJar9Ah4zL6EszujE3PU5QgkWDwKVxM+I5OXWNMgXxQUxLFgdshvMica3PAEB/451r/dn2
Z+ay7HsFU2QJIGWUlwJIn3tGGUZykLdQDSikuMqas1QihobfqpVUnJwRe5qeFCjZJ0dKk/to5TX2
wYcmU1F3olM1fKZNkEaDRgKS2i5/Hu7eVJLniMDJcpkFgnwwbeXjHHY58IGAHk+I9yjlmvjAwRRd
wC6BP+pOqcZjQUhGX6H8F5/OaujWvushHpoUADjvAd6+9tuZ2yiJR4TlDSC10LSdAqnMvrhhSwN6
FDemyN5iugy0yzZ9x/daLMczd+5JFRos2ZggRMAHdnV5YY1DuHp4HTs+fSLlq0utbA+DW9j2rwh1
BsvIxmP8LW2KnzykHv3KB1rawd/IBkm1YfnfCwUqxoL2VO8uJx/2RI6hxoWjzX2zzX2cqnpwn5UY
Fvi5n+V4GYliJu+u7e0I5D/m/rB8xeHuIwNEt2SfcvDMRf/4wuoVp9WzoQBPdKnFYhEr35NDI8Wm
xGTxBUA3nz5gNNTg5K+LviFM21y3vGxHVou+3qiN/dOtMXGH+GQ3ntAtsQKw7pNt3mFJ3d2yIqr3
PXt3Lgr1esGQaoDkp3g2cEKXIFsW6cn+LBoZiS3hfjGwvwrPtGoFpQMI2/sJ0TiNmFdSS4/hd2Ah
G5P4ExI52zI4KS1ri3kCeXrbW8EWjZOevYl4Pl8UO13nPnQdmlOpNzJAsgZ/am1ZLKfueQ7Vt3N+
8+gPZKC2nOWlpXkoQJepbGaKrK87ogJcBzG81BEntL8pqk8GdJb0LsKRGfQNfaI3GKscpnGDo1a+
wNF6VsMYK6pk31z7JNsA1t+XN1tOEaTaZqtIeALW6iJLniQJ37mmTTrLaHShAnvZXYUQYj5afs5W
U2nqY8saiRB4xpAJTP0mDbSNwCo2ZEsMQT19yR8lC8RI9mZekMV+MmppvG3eBcRENzZ+NCHTt6gH
7SOQymDj2oMQIl5SILsecyim+AKFshArII5dPuxd6rFY8F+D0MAcz1ikQYMBp56Yrlvl60MTQcyB
t5XeiSqVIQMKtoEqLTmCa6mLLw0Clkqve5dKlWa8fNrFRjzmBv16eQrG7ITAWN+9Y2GR0HWc5+42
xDHUK9dXvAQj43aWS+0V6jBOYF3NqZle3II0Z+W6yIPO3iuXXF69b3jNZjW70BHl8CkFAuvvbVC9
egc7MMb61hZfVs5yDXFTAlQh4wUjn/9W1kQwwHYvSOuwb4ZF/eE99/6qHp5oo3ztjkXSnP1GhfQ4
4hU97HNFx986SCYF2gFgv7Jh4DVx20aGvt2lmWPsv2TyVUXSopblm5WXPiMiCp3yCzu8K0gyMWF4
Hqd+CzO5fc5TKyRNdnBlmb+/76BenxIJOwJuhJa9DLrPXHLGnOseFnGU12/+YmgNut6Nm6/yOAaX
RCDblPSi6adTsbv2pDR6gek73GEASs4l24C1OZwiC1mS5PdQO9sJsLQ0SiybsVAK6bvh/NlbYGwo
REk4QMM2ZmQaGx8pAUmx4ggjBcRImkjnvS2rO2qOaZ5uyo7QNVgOf4sC/+ZTcijljMt9xU7Kj5p9
/pMRo0RIP7Le6k5kx1ys0dgEfjLIs0uMiqiFeAlxq0t8a+jZlWAX98/oTvrQ9XqU0vwynfPHzed3
dZ7yYLFSiOVFSjA3unM/L9OWwYQqbv5nXGJxTudhN/5owZYDGB8U/hhHkkW0vDKXNgU9alX8CfsO
/2swRffFkbiV5fzXdHXnLw9KnJ8FUousxYiAn6HkW3jP5WBIyMmOkdGlpANnoaAvIdOProW+W2GW
35+f0qmgdoMTPsxzdahi+xtPP65ChjJT1kFlfuiuMCYAeFbFI+v/DShnUMgwuAR9Hh4uEm3EApA1
vUW9Jw3h7EaajRM6tRK9JpCOKl+iaS2l5fIpSztqOU3JZo18rR/6kONeOXTB5u3VjwtLfkiQJtYt
F+/hH24h9REvONC5jIOTgOWDwnblCKbgZ/9iSHwCBgTQvlyADUNO5KYcnQP1K9zaAKAu/dvW9ZsH
8p3JxHovZVX8nvydrEXIaFOUIykFy27+vdVulkLDwT9S+fgyF3QCnB/wH/pv17SSSp1iu/bvlY4m
f4ypLlnFH9nFuJJSQ7Q9ZyMAi2Vckxe2pr7lz50QiOeMz7oDzu1HdWyUb2uBZKhnQQ70Fe2+VJoL
GiG2HNdCbzoXC6tLx5ZsQ5djlcCdwIOb/CAPNNnSB1K35Rzl+B+bYl/nvZkjorApaq7Fb7FtbnqR
sP76pdImsKRhCFM7hJ73O40/1S9ABjMq4PceC3Kb6TWWizSSZGmW/QilXByEFZ9GHNTrNWZUjPod
F2z0iGE4LeJuNxIlbyFhOfi7xHg1NRqYv9dWqfRFZSwTSDaqhZ6kCYo2OIwAPS6r/u1qviI4vEhq
kfrjuSqPbMiwzRfG2j2JwgsumY25vHaXaf9LbufVNJBBTcQwCwMzyUKlicritHamI9t5Q1qRQkUt
LQPeSOw6d+R4ibAx3nSge1oVltzC8hYpQrO5UmHOwLPpnHDjLCxWXXOkZK1obIx5e/UvSfbAZQUY
58sHccDVcPI9CQPuXu/6TDl3/EdbdtMduQpsAz6mJB6K9tsMVrjpaTGTg0fVrQhOvCX2VtTOs9kC
fxYGz1328ZdNE6f2iyZ70iZo/TZAgY+CDHXSqwgvREO4g5ueUrf969u3RyE3N5rayjgtycsx8Fx8
H6zl3OVBQNj8ZOpSZKO390+g6u+SPrylkhUxArqOQ4QwdMRU2kK7Lu+fO9DLGyY3l9bQ+KP8SpIV
iEmm+9YoWGDYKwptP5aIilbnr1AFwx3RWKSArQy7egb4YCwPG7jEaJR8txbME315qwCwgEgLFUdO
RCH28FMhLIGb4pU+TmDs0AT/7wXMAZL5fMAgTDozIR4v1akeEVpkTk4LprpXJhJr/aj7aqmRRpYo
1JqZjZPW4/lpKG88tomjCiD9X6qfnGWG4OCZ3fgPmnzsQJV1+/tD/0i7n4G2JNe7zJtdd6aVTRUL
KWIox7tMaX4dH18n+ckgJtkoEVSXHLp7/RHeDzciUGAmrh/HiuqR1cxxCgJBbpfTexAdPPKKW/n3
XumU1quI/yjyTunP+OdZn+nhiMvzoeAXmNbutsGLn4/Mb8bl/Fhu9pJePcdOhPjvGmTScHyavRCP
tFpl7S+in1k3X25LF1YmhAqUlOOvoWHHtsV29i5zLCJA/kap12VlPKErcK9FuFe3MsUXX2PhRZvw
CXA9VutI0HAnYz/EBBgBkXJcLuQnYiU+iL9bmgNgI+THN3ZYPIHeMOT/mVDQ5tZept4sLRr2h1Mv
yJ/mHeNQkKok/0tovwhXe5n3bX7FhKMWi8T/i/cfL0ZbOW9R8ctyHIxv6tfb4dOJDpH4sPVWRNuu
i55aG4S1GlvXOWjNzrLIZZE10GgsZzS7ePCZgi61NAH70U6GQiJrGKmvayjFwvqKkr2cyXMF9XVf
ZmHvJZ1LBk9AJ0hf50caAVjkl0De64QQk+eF+cNSkFzOKaPEMNFM/KAnj14QiFZ+AXv12UdP15aT
lKndFXGt+plg6fzg76k6UXAUb88OC01/PfLDgXpRnftSL4yod03qAFqrmvvD5T2L8aPujSIWteWE
2VbBUMN3uA4p9eY78hIQoOc2CMRtC2AgkHTefFcxFxtowRbE5yae1zW6VEwvjYd8/a+3JH3faP24
RLQ824hl/R0+tpMJkwNpOdF54ypSF7hovhmpTNvpeQuNh2r8Z/5G1kiCe3/uzXKktr15Y63E2eY+
1n3qahSO1kUoRvk4SVTPXQxJbKuQpOLJs7lMNZqld+fVG27ltwleV1a5WdEaMZg5GqZii7AzfGm9
swbDvi6Xd3mJH64w6kP68rAcr6JM2z4BH1TpVSZDDyZe5ctc/XxLsFFbziRjI9FOGP3ByZSTpU84
d88zwx85136JmuL0/9cMFPhvnwRS2z2TfrrzYMRYNyyga/kY39BbC1dMYWarpfQ+KtOBXDJ6WguY
j6Vu8XjgC8hLyltQ7TgiCNi6FlYRW1c0XN1QlpQsNDxqBmBkhpthRuJS4ZHsbuA0+4KNbFqsJNiU
XQO070V7/FnogR0kG/Zf9QpqCiZvJOqlNvvTUVjhm8yk+T3i/vTPiCn4ekhUEXGAipjwMoXRPJpK
5vDKvYCB4OVx2oSVeitwRZA+p2niXXyNSOikat0MO6nrlP9NIYCvsHF158j+JnqKIFFZXSn/JTQi
nKbDlTBjwj5VqNTEHz7OxvYY7Ze8wLduWUw3SlLujsxbFBlPwbT886k9xYrG1PTfk0BMWRHK7w4X
fgDWcXKbjWTefsr9969MfVK4hAx1uTizFB3apImkxYs70Rb7sF2Om9rq5w5B+a9e2TKCwY6SAb0g
zaSDUwgB5bnvDBlB6drnMaZcLzGmbLzESuFaZxSFOcaTw7PcHMSMIi8wejamHSQkxKKNspTmnrPL
EOE3wIOC0WlapSvXVfheouYt7DEm3/4ywWk0iH4ThKIYHL86a2MxutQSW+mx7gHbTl5VUrEPSfaU
TA4vkWPkS9nB+9rnjRi6hknCcQIxvcu1hpAdn1XS8Yx5EuPR6Yj9Si7U9pPzBvOjFZIqQo1GvLp6
ymr1An3f7aEgkB6/OSx0S/ZieY+FOtkais+Q8gmdQ7LVRm+4CAz1Dri752NG9gdUBHu5vJQGGVOL
Hqpi1c4xnsullAgaBH6t5asQKT/a89q+ORhhq4JXcDwLqDqnGCTquLRdsU8Bb8KgBh76z9pGJ+/F
P7RByTvZiE76nMJW507aLeU7aLgcr6IRIOBjjRUdEjcsaqwc5QQJvtSK0znGp6hOEbLug4lNGZ8e
3cP+i5x3chKR0sAdEBIQCsG3/6teZomrhpO54x9MOTuLiJEhycAv68ItVz4iBcDhhICTHTmhnPEO
//yJtl7gDkaMuVxSSLcXVCHCLoag1a+jJpzgrVaayyawcIysVqJVeppZS592tfu+//1Zx0q8vj0g
yaFjKTjI1yefD4DbYjqe30LXVz9JZ2MZ4hyeKQ22nJ+kRLQHjvq4ZwOXf4xdhIT98d9i5QdF++Xt
Z6wv+o4dhNgukyHr/dyZWA1RNZeIboq6RINhq1edbVv5KNvTpsD4ixlEPTJtkeLP+9I1dxeKZy2+
D7SyL2jtHpw0lq9mw54WDf85W7xga6tmdM6A5Id5C6pz/WJ2yVFMKgf3ZyK80x4lO0+VSSrAn+SS
sR9lj0HAGluXuh+O1cVND9rixs/iZZyQ1wpzt7Ga1ZS4cT3XuzYn/xl+lGKsVKiQFDerLu3bOebo
p7z7U3X4LVzb+DlZ55Ixlk/juwXV2MZc6UtqYSND4srHVO2LuVFeMeXGYhJLIExQkPtoeiL9Yq+v
EagVeh/2h+NgB4cwkRL3GlBvCBzNfzrASrrUrki3AASyvtub2iFxsC3BQ+PdA132pYexYXPmbkPj
sENZR1Vkp2VlWMwAItGaus0hg6yfTOivYdTtCcoK5D7Qb2QzjmX4UVNXc/Snsrj08FfsjqcZ/L3j
xY/J736Nxp8kwuzOgSooBRdNl0mvDWZlmCQfRgY9+vNgG0eSp33Pw8HYEsSHhOLtJ0RyEAHRjqem
f0zEkdtnWJP9CYFqyiVp4COp5klnVyZwK5c1ftWbyFA1HrKwd5A8jJUQJElwBb7XUZfxkT7KZzrb
LFHtGxtPb7nYZlOF0sLtOipFU2eSTjF/a+e8MU/PDqQGJIscKXirm31HFfj+yeXgN4mriJcu8VFr
IF0dydSQ5asMhIfJuxcE8v0zlpyPIaESGJ05C68trIQg/Adl8J7ET0+EZ8zIpXwiN7naClyHx/5b
FwSiRTkWdpT9ctwSgimU8cAmLKlLiJuZSoiFvILvVXe6q9jx6qvs5ojHsopjaJ+VmKJ+4jvZ3ZHr
sLOeox+RusOR0QO/cceQIpolKoXpek3WT2c7+lhrOu6u/S70itNb1dkAKbtlbq8GxsEDYDggO9E+
/Sx3VCs30pbyNnfS+Mhw2rJIp8NSCEvnlbRAkWD6vvF3BHpOpaJgEwUw8At+qDHnGq3a+gRhutpL
5/YKRrYNGuagNdZDdaTrU5mmqR7byVgaqgOslVHAQeajB+83aXi7/gPsf0gnFa0cmMmi/i+ReuSz
JzJPTzZbd+dJlpHT/EdRRZBmT8IHLrarfsWl3yKvI0gLBVyjST/0r4PITdXtZfqnTOwLtK/B6BTU
FnB+Bo6cEcrAu3rJkZNjsHTk8z0tEFtF5hLCgWIHOvnH7vOnTYKzNes/L8vzTvpBHyn/RuDBship
prIjegvLlvIDG6VImDvrGzhJ3nKyeMvRptyxxM9AfXQ+CKQH6DNygE7q4FC1G5EEi0+B2AM+4log
z9QYvXEtc+XZQpVJzcW+KP/jRfyzutAnyHo/vJcWNpT0jaKDyXvfV76EVg4q183hHPGApMFWr1/H
UrAPrMbtCbwdzujSvYCzTUqc/G2IsZsbSwYMvYaxFNVuzBinDT31MbFBmzQR4LfoGlnN+ZoQ6oCO
Pc4orFEHHjxpH9YqE+Tx2LcDLO06QdVxIce6MwXqpu0cVlcu4NzbZpkCcpFGWuKX0WHSV3lU4pIG
YkksgJfbUxAPiEFE3VlkO5U7kDNftLWxIKavr+CTVQVMLh4HE3E6KhEeeXflDfV5ZyR71PLCC+/R
VNZQTteO3XEwnF+Dxqt21mXH89L1HQR7+keMOFKa91y79V4FIcywom9EYzNsQcXrIvNp7zucuNQ8
ZhONJbo2jizMiI0TPHrUC37UcYO2kewn/9betqW9rEfgH4Llsde9TqQW/tahjowoyqUCfzaNu7dp
tjCtP5ORyAT8wxU8fwOefvBSdkW/C1cdfY9bhh79Pjg6VVLLqR2NY47HliC8mr8I9roZouL51ahG
lnAXZqaYlQ2lwDVrizb/13Y8wEdFzyvYympP9J19LO02x3cl5zxg9tBPrcDx3fl7Ji2gts+hMbGh
SkNJ6fROZa1e0LGCtCqPV1JcJyF+K/bYkCjdo9z6MWG1AourZrG3nKpBCx9E1jYBwQ9b9u9XT8Ns
K7BnzYEAOKQXEWmNRcVXwb/g91QgKNLkLSm9LAJbABo6b/yaNha1gyk8Cke3U1C8QXu9uMqLEmlq
4tNIJe0yFGJg82kyRXIYBaOe526dyiLjxW3/RbvaQnLX+Lb9BsvxNJfLwflhAtFQoEO7pqqFD77m
aEc0u+9XUxjU7Q/H8zIJAR40dwCutGbeY25m+TwANZujsjHJHX0vqZXtzN1vNhd4C/237k+Lv3x6
0p5KSEB1HqH9Wvade0Jxz6WFfFN4A7wXkh30guG4FNsYCkAUOZxhRkGYfeo9gYvRs0F02NpbvQF2
yQBWwOVvDgRM0IVf2w0gKBHNi8LSC6o/bASXI0ltDjkItIAcMhnq8WogqwH+fJCCaL5dx2scjOa1
I28Pk399irwIxVxBzaVZmuER3+sXRQTDxxXbNaHpXFyaJ/t/swtrG+jjRkZrXQC4oPvSYVjsOzko
Ixid1lDc8IpVFVZJnKCtJCJZU7xEvKZQWSmBxT047BTUhc14uaZZJc85sD92bE8T0bXJuHSZfQeW
GnojNoXxFZ1YF9uTrPmYXJR6eKdfz6b9ojW9vLc0yE0PC4e0xadabaE5LzAQQ72QhAaW0BhCDV0M
jFhiS5IGq1JCpHkGBdyHoViuFxYWMSh2tp8+aSkIOJBZ0AqBjQlFt3mX5kYtRibApf1XTUm/h08/
HR9Wvmj/4MGqY0TF8Z5Gd8JyZGxCc2MnqAdJAl6IKuQTqz0i4/yHX21WKWeBDNAHnnSRcX0VD6DH
O079wq37Rx6k/l0pVZsAwNCnI+O7yKggTi6zE9/cXeL2Ew8eg5fOhLaW3L8y7jmjS0bPjc5arkmf
mgiQc/I5/01Tqkv1mP3sJGhkYi0OCjwPR9X/sn3fl6iKxIjS5NEMscec71e3ETeR6Y8na+rOrIRk
T9P1+xKKAzr9EpS6qgDGCXcSY/l21SCyg2P2xRB/5RUPt49FDRujQ27pRLwVhIFpAwqjsSwOJBk3
BIFK5Of2PGlBEFGifaV7RJ/mo/qGkqBw547WigUANSY/ni83ib0z56vdncjhd+vfqr/sW/eGra7J
v4ORukBkz9rrdWmKS4Eb8W73XNno7lUoZdTO1j+PnpgAMzg/8dOUhS2lBy0KvBl2RSMLCKBFJU97
xK6uiQCCBSxdc9ETi9pCAdnrYCW+fPxQCsqZaCGV6QagJuiTWXirx1PUjIteJBhYk3TNKRRTohWm
g1dtQRuUDw2C4hqQx2O3AEwjdkl8X3Vd0bi5YqdV3zLjsjPLzn+fIniFlaXCPV4muHm7yj73XFf1
3t4zyi6xtn1+GPEdOyRaSU6lpzASvhl22wEyEyY8h8MMR7vvGT9n/e27PLlO8Ca3v/u7NTLRYIuQ
DWKf9ATajdQrwrLtBIFVy2hE8SjGOO3Bqg5t0L8V1fMcLAPzK6J/BjnSvygVlj7jD13tu2axpPqf
R8U5C/k2ICzNFppdVgeTR+jfVgA7rGtIErV0V2YOOLk62E/lScPWjygxb658knPPKoTWqJs1dDVJ
LEnfna3/TZmRN/eQQCHT7aZSfFEuKmNHDUXYvoiyLMZd4ddGDADT/T0dTfj7W0NxZhyg4rIqLmGz
onf8H2WgTnDzCrrBmuC73ieQhisOz28tozlH14RUsI7bSEHJgv9Y4aFAjo8hdbDZQlRS9dFY11WV
N3OBoWQhOF4+Uh3yJKEk3KI5/ObG+nXKwXjLmDG/72Mx3IJgyAfMf6xZZdNmcu8NLIslyViLmpNX
eVrI9Cj0vRy4/N1nZbWDEoQeumEB+LVxGKhRo015xlAbCocbtsezYXS0jL+9PzrA2ZVQ/z1TxM2X
eqAX1teOawuQ4uSKXyhSFgntHzHsJJuCzD+YVNqkLbihkKPkqJGIlRhc5qgwmWaoAfEMEhOj75rt
zAR4KTzHJu+cWHn4EQhjN/1wRtYZrPmB69qOZ0bxtWsC1vFuhCDYDXkx/h1eTXcrhA/ciIJLebkR
OOQsDUA9+NShtpnvVTLGyRmAVgW7K9rJst/JGko9hofiD72c0i91JOkITFpTpQTe/+udaSydkPv2
1UOIh52rF9LWL3RB/5A+n50U6kaQFpzQBAwjsEs3lTH3VnfdO+/Yw0fc1MCoBOq4XQqex++Gg82Y
2HhK81MY1w0Tg7hlknHlmUQPBYrOzZ87dqKwJJHxr33NlxKZJTfUhoPb/GpVOJSI2GJnI0VsKE4D
oeY3gehurWkWq3yZVHxpNOvhvNjV54kSfz0BEKrgfyDhcCtPWv9DnfH6duTN4RapN2gNhUnAtnJi
KoIcZhGP0bScyb6gyYS2d81cGNKUdH8HP390KZ6jmVIJIduh2jBLM91btAlaOGkS851JEznRS4nd
BOaw5S1GYtn6v0lGcflGzp+TdqBpFWO1fdYA+5nmR/oNnRIqOGewnq+p/8ZehVd6trDIHw7SshrY
l+1iuioi8XJJJo/KTmPbQVX0hPdWU70V+BDj7Hz2nJDS7Io9NLhtla3BaoHd2h5rAC1qPVXQg/xq
+UgAEeQ6xLIXU/d6qibG9ZNnygjy4qE/064lpe6S2GVEd1o2DkZcAHWfcyHn1s+1pWA3xS8FNcLI
f/el1Rum1kQpuDTrkpfTmIR9RmTLObx7bajV8Adp5GrKXBzk2JnLpB270En4eIlWGMH9S8vPZgJS
Y+wqvaIMp0p2HIxd547PFj1Y7RNS/k3GxNfCOkqbtcCWKZ1k6Esx/OqwJkYKvzANYd6yO7Ds0Ih6
e6yZm6pZV81KT/nUSrmqw8egoQQG5/bmupBOYtcmIAt8TzjVajurLDq5FUqy+YT0mS6yWnScOeP9
rzZtbjG3LZtYzAldte8zNF8hA7tp2VlKONmb7fMa0L8OM4UcGr0tOClkDiAeW3MYn7i0gbjv7Zkk
2UmBxGYgVryVot+uYRkeh6OZixh1vLD+kQFbzdKwJBXZhzuJ8qbvuq+rrcXmYnJp+71mzRsNF1as
RpO7X7dDm0kCbtx9fB4UR/2tDyzfG2rb8kY3szzyszFqQ9BHSVyi9dzt14w1mkudS+3boG+VNV0A
Q9MSSLmivJBb/bXXObKhesS5oyyt8lQgubLfTMnF/D3NaarozsXv+Ic7G3iP6vrjuKOi7hL8Y9+f
2vNtcgFgAbjF4VHi/VKNZ7EFmRYmv7lGFUM9tjh4HaB8D3vu8yQVxJEJ3khj0d2nzoMgJudTfs7j
ug44d18SAcEm5xwlKjOZpAPXVOldsDunzS+0+7+XBwfJwK7kGRjbgMKLs6fwkPym3rIF7y7s+4GG
mrPVyuyM7+bKt7mtkVyyR8095Wo3UzqG5VpogOE4Iz2BZqiMmLCye80Q+4ufnYFUYx1NvdVTAo1n
AvjGSdZN9RGH0FxVNd386A6MG5Nah1eqgif+mS/kWR4B2Agv57U0NbhNXYJ/z6HpbNpuGo5CyAr4
SXRgfQuvTFitlqFIw3lDaldqZb3OtunzRw6AqZKo26iB3xUt8x6t/IP1L9mV16XSB/4RNoiXoCUK
+HuLNQcDYUEUU7AWk/sPYlkBGoqxPUEnQ5qmGrjXF9MCM7Qqd/dRmOMWg7nRA/K4g0bL1t0ObM/m
1sfXOxI6Xnv7xVzTg+ubdyHMiuUada72EEKZJX/E4nMK6ZppKe+7WwJZ70tsaGm/ojcFENKq4lrF
CilwrYxQgNbngvcHsqaJ4iXW26guRKOFHWpD0QLYJ/qzYfEEq5O27CdRTZhEalVbebdYHxb6cd05
+sEL9W/aJHwxvPYw7wo30xygJ/ERNjmAOkSWsdS1NaJGV/oC6xksGDErpbi43me25XCaCejt8MrO
dRbS5KMMK4t4TAceoyTdOfnkCJ4WejdfJ+Te5ldIJ3qu2S58MChaOT1/CYsz8qRF3gmuoTAKXiNF
DGFP/n8hSnEqbHYvM7CT+YSl3TlsrFVkHEbA25U+BBQFDKsnTT8a5zwFsT+alvfvG7XD82NlEfMs
yfRMICGu6oY0ikxuiVovjGxZvNCfedyatEhz5gWn157QcknR56r1lavuqmfEpK+jFq50aXc862Sd
8s4WcKAdBsSOl13QOUKGKwbKZub9Q6YkY5HIZYQjnWHtHUPg6QoHJOxOptPi37g6zntW/Df0Gz2e
cUoj2Y6JR7cdZIswPlII0it/FT641jRkANhMzIvDZ8wVfUmSntUMuEvD17omf0vokYvNNxtJuvbH
1MsHCILQ/vd8T2KBokDHIFEfcuYTUONKfAUAqPeX3jZ2Hhcu9K1wEcejTawBMuyHGTEixwC+8TGX
p6KhDA8Q2q8ro/xGPAGu3S5C2gDckpmHYRYVR1rzPGcHkvZAho7Yw5S5RMsnMQylgVI3+dOs7aqD
vlPjikJtA+MCPsMiqK/ppeMLXhutAofsU4RRRPXB2xKSBa6OrDwC+siH0BnbqMdisWtdm7pXCVdk
tOzfPA1ZzjMmntwPgW4NE3s8W1NaMf2kt03qqzRiul5wx8rJNudgQVozFrXm7ij1ipYnwt4NfpO1
nNy94xT+gpkacIK30xT/CLvQx1vI+6EAxkfwnRYKN1ES8WAjJ7SEYi/bGnbyUTgoa3AHFq42IJrl
jSc7AYgpk9WV9Yz3Y1xPNShXzHdvQRY2lKdPxk8c1I49EY8DrgFLxMGAs4tA1FS2Nke7Txf+DX9p
tYM0IViPe5/FsC3R+UgUC0Aav0pzC9DqKVmNDeSStFoV+rdMOeAa5vUVCuO5knxncCyF3JG636wi
Oa7I8wvFX7OsmMNJsPONTuFP20Kq6O+UbjwVxvS3fIntvMwPFHhRq0xfu0C34Ab2JAd5qDoIj9Tq
iS+oRWvXTiF6XmyUjEsJjzjkzk1VdizXcnuCIrtuWzhZpjvo+E9FMeO2RgifcZODafJbA0A51b7I
0flkJSycaPPH7h/3TrZrIdpi+nQrB6bSjt1ARLcM4J2jWsg0yScWEMLRzXjX9/6LK6OKsjPhY7bn
bGYwHhkBP28AZoUsLgbUA9/RTvcLWsHx7fWBSbKqhsgbBwUK69mw68mpFTdRBd5uPpMG4sl/V+D3
ABqbCtcydtJBtxPUZ4ermaOg4v/qVovukzfPrLhoLd8YLpPiB+Ng2f2PCu3x1jpcRBmakF7rDO6J
SmfLpZnvL+DmZH7V2IXIMl2it26I+6ZcIkSNpvMVJ/uDDYSiqa6zVUfYjcoOGTZYgnyKGjltQ4wX
tTH+rhfSR0HDJjhWPNfQkSkCw7dEtI2iI/Yw5X7zN1a+jHJQIEotbutsueA2sY6iJUXd6D3zLzDP
BDels6ygtsom3RGE3Uhg3Hgg4jgIGr/JI7PzvcskE9HXejxThBZASrxxBDK5w2g9BuPAul+Ooboj
iKmGQ1PS0Rlol8gd/QZyjdGFthUS6hvGJqPQdK9W/lJPXTyivMdvDehFxhptiOJ0a40duaTd8KrY
wc0syOosgfvSlQHgUopFUI8rm3pkZY5xruX3oUo47rxLsOwzEt0jc4NMObDax92RQ1ZX2zAhOVLg
qbPwB4oLyEFFEhMOAKD+TIDjUZ6UfuygUvEkVG/5+yyP3FvJa0nO3XWoAA0WWknzP4q4UnagTQDZ
1gQSbXpoaWo3CWKWTDJDHZ2K3aedJuW3kNg8qgdb/Y3eSt6iUlpUhNKV1kY7L8XvxQ76uV3ggMt4
jVSnmVDig9GCMpRLkLN3tHy/kBwwkoZl39dCYffMo1Rb4xpXEx1IX+z54OCpJbQUJpIZxRCG2wD4
td572Iw5rxkoPdtiOAHxeLlxEDq2Pjis4Fey1x4y71aKIn16bQyCMVFlKGNdQRhO8qHo7KOkPnDj
jSp1TkYSfQn2Of8MqFkz5tm3sSZ9LLvbHfxdRXgXYpNjba6ersqBRnCud0zHgx3tiDP6PTxW6RI4
32kBJKHNPySRltO/lSgWJXsn38E1f1aIrpWDFSk99pJzyK7+rax+GmUlZ3Pc/FYCCep+TysN+K9a
6I3fFeDDpzQz17TTVfJW+8QsFPOHL+SNJtIQgipJDbVpIcbKq9tcQg0LHctiH7GXFCNatIgAdEs7
DpGBS5uDB9RHpKwTdzSK2wPLRNmWrV2ZrIKfBF7gBNYHqs1u3AvD5R2WzczcTNq9IFF3w0MTRpL3
XBQ0VY06ZmUpivECXNk/LocQYK7lDxAnVdjZ270D/7wMBW4ycfhRwDQW5AFnwAPnkZDW0Aw5b/zP
YO1csgjNNsyZ8uLAWRsRv3my2p+uBj398zNKiqHNWKX8zqS8EVrBJY2BU+TpeJtijbQzNXheQP/f
UuT2wQJI5JLgo2EG0J1Eh17Lx7HA7THjsmf0RrwygVC79VknGhHWTz6u72WHenQuQmHHP9uhhmad
P66wAGkAF8OP7NPN7RO8USWXoE4JJZuw4uJwDRs7z6oL2b4UjmionXrIC/7nwPKgI1rJNW0ChIC1
B6GI1Eft5J4LPIDHX0abj/stMhmBAOf0Ygw+27q38T3dZ7pt4Au/GeRHF1dFUTWgsxW3DIXpubS8
DQebvh1xkg4WuZCteJQDNbw9JCtzeLhFDmYjzI+J5thTIVd3EnmA6oTLH1HVNuqRdIH1ULpbVwva
KQXZ2OxK8tte+ZdDG6M7pFtDjV14y6GMctuESPxRu3Ftd5+QeYsGjBeMTvR9idddyLuZy12LMyj8
0kqxQB4d8CzxqQ3F5XUa/xXm9ct93COyW1q2YhixLcAarP2ezslpWqHVy7I8HOuSaxmuDUl4rUfe
tROlFH8E4V81tTU+tHaXBGvkp0KunsC4Oi3xYspRYdnmZfzogr96LXDUlWILNlsvsVxJIXRdRGEX
kHnpUX0IJxLvZaSkkwz2SSocsFBRUzHZVr9Q+Uu/K2EYnueFLf4ROAwbCzL9g0MI7UAY8vJq4pNn
RlvIva1k0LiaL2jbfiInxXAy/xO0l9Tlwvgm9+vMaoeI1T0pVLTUjLhb+QxduX8KmKAA7SyHstWN
xUMY82LKDIj8aV+x//3uXFJSefLSM5g6nZb023Lp6mX0PPkDo+J3DYgdDhRPZZuEpopYfz4+XQPo
3figgS/5waOPRxeDtAWSqRe8fZJLfjSRCXe/eUhkzqpmG4WVbwUKcyv+e9RfyGVRb5cW/aHKMLKa
a+UXWltU7ZpQ94ccIV/olBZgFAAj52xj476nl36hgAVHQJ81NgKqvnLTFq5MqvgqI77kW3+bu2pW
6VO7kXwNKQRlpVSn5FRlwgvtc7Hekku1faHJ0vXTRJUodxMZtZHvtpZhm6TFEZrEA4eM+ox9uhnF
kA0VRpjEIVk8vePwzGB6hvEAfasgfPspzhi/oVjKgmbQSuXHA6u43EuZh7pBPRxz8x4zNZV0aokT
5IuCDx+D16T6vNIAH877vyPDtoyQV8tjAe3lr2ZtlQ/+V3eTdWGK9KGPSLouImH7Qd3y4dxBgFKg
D8BLEcingfNXgMBRYQo+WvNtgcDd64tgSu8jdSYo7Y5dD3sQWmAuN8u8BmIX4buIfRsjnFgyvySF
ZeoRrbXrtVKcm0iAhpGdU8QF90Pii8ikxB4gKo5XZ7lgLw3g5gsD0GXEm6k+VRK1Gpo/HkphGRTi
RdVD0qEWrufKFSiOijvltLfA/rqTruVWDBppKjSSRc9jCtpBQoptkuoboxGeKzKNth46IedjaH2c
ilO+Q36DHHBtfb43jAOS0uAGBQZ6pHIYNFzA6r3x8DNvfG+EmvzR8t6y99STpTQd4U38uny6+R22
J2qcg+6GBBfTLJmPL8V/NPwQuPM/AFanZWIIPgBG02lJ3sUtodEIUKeJaYGDHXQbTE1RQNgWk5yg
tPlxYzvwAt03vkYacTXQY9lEHoncHqSYo+a59T0etTvOKMvOsXyNE/rgamaVhPAoAHL5xbcMUpYM
YfnbjBVM3muoYP8UAlIsrwPjLnOsTqHmj7tKy97O7gW/7bPO8+OsmNUz7C4OvGOiemHSga8DAYjK
HOnYkeqOUniiWF0ILROxfF23OtpEGgfRb71q449SioRzIBeItJybMFYG1D+6JUr5yzBAznHBsSs6
4SrTiJmZzlyzEIxgtE/YQUD0M/J8yDe++HcGOMdunaL6p/HXkXEGVJjr6EaRDMkHss5fqKbA7hUS
IPbxYqT8mEPXLvxsALpaI12ikx1JeTDX/6nTv9Ga3WhqupsWO8wy26UL1fQaxcUcChn4XsuBI6Sf
U32E7vsgtJhNEPcc73N2xUWT2fFEqgbohMsluoleDQhaAXYVbMXf0oyw/jt1XvjU5hB1fHKkPxJq
9nWGvtjj3LgUH45iToiBmzltDpso3sdHDFeZ9Z/D+4e95d6wNYFnzepQ5UDhSeZlgonN0R5KNUck
oTNan/RZZDyb8uBQXITfTzFiB7DQC19/SbXX4eaa5uAxWmCyrgz0XT01RdxqeUvMySL1CC9sOXb7
sLZ5cVBaOGvSO7UJhZ65cKhPSv6Ktrs2kW/1i2sb84Sn8YaQ5zUr4aVyi4TmBUYvQuo11aKYhKJv
NWYojjZLlcPcSpNYVnfkmf0bUrhrsk6zIG1Ou62djjtsnlkBDSo3C8rq/4JE1garLWw0QFlq1Ra6
NOUUHWUZuYdaiAtkgGgSlEaUSJ67ZpbWM5qYq9iww8sNmBQ3vVsSRpPvAQzyF3Jqah1w5qx4EeJc
Z6EB3qg9TByUTXi+dmS7Xp018JzKSZITBHSuVl7SZnLseSWPa8Rt4hqtwS8SiLnZOI7ux5N9yQG5
Lg1rSnqDm+8kd+jscJJLIGf2FQuIdY2JagR4jXs+fhtCxu6BMS5Vn270icT8U+oFLzdyp6L8N1XF
00uTBxbNjyZUEVmA0OJhGITNcYd2Nd/Qk7ZMDa1RoWCdDY/gfsPjtGa/v7nJm/F3V0ZAA/yaJRLx
1r1f0/e/z+o707UA9SlO8D+Oa+Ty+tw1IhM0dpwmh/4AmBd8nDmaLqZL0lmKDBWGQ0Vh2Cpi92In
EWaRPHZZ/ikyhYKEd1phmEZLIuZYeRSSMBhIqVsfNgc/mW2D3u480rjAmncSSZPKwYiKEr50KgQb
WcRYAWsv0lAItJFxaGSE4WyTevPby3j6RPkCL1DXn2r34z2rRNBBJv8bD32EJRjouaeVNjpgZvzI
nJW/dNv4PguRNxwa6Tj4OgcRockNRToEJt54+ny4jFofpz2g0hWh7JK+dghM1Qc2ejl1jCn10ZI2
jMJbzRuOFobAtwL9tA17OHayic26GjLgULv0Yt0UaN6fOMCSucb6h4P9kiW4lPClcOIzfCub6W2F
VdM4f9ISXlhE8XIuKjy562zAu8CFn6jtC+K+EMwNtKG8m/7v9YHPHPRCHhLWyk4OyDq6QN7FV27E
UZ9rSvop02aMOWglYCNneCbhGWsZVl+AACp+/VnVKKXrXxEWqlxr9kRHHkSvOWnTSwL69N2thtrv
cAe+OsVKOqapCJgFAUJt0FllUb9WFyEedNXY3tNxJ39huBSA/CXCyHqlQHcvFoIh0Cge5LL8efnq
r5m9cBrETySRHwtNkJBge5k54atpBn3qn08PjPQ9OTudNGtxEwPSIybjP4JKGWYNQv8oVvfQ6ESh
oXcJcofB08QOU/TS6PKhquGRX4GFnwdn4p6EprrUoVHkswT0OekU/WmuvnTGC30ze9N3Df5AVWDF
BPVXEgZGEqHDTVznVa6P3mxyPwueqCCV9Ekcp4EXMqzxVjmLwU6f3XhK5sBy2Z+4zSO3G/wLET5A
yoyHASF4fEiIui0Bf0WCn/WCncgj+k4gskq+ICfcwAfhciYtkoKPmnO1kILtkLHehuRVHt7JPSRB
8oF4NGXarmJho5vOT/qsvO9uiG0tVG45j6ydO5etRGoQrrmP0kf1huNXiiwl6iN9O/R7fuKZmSPN
Od5g5d9j62mLoZJs+yYBYaF8Y9kCw3FomQ/ayA6eEXhQ55cpEzP7dgg9nTuRslN70izSV+35PV2F
wtlqptXpxnGg8w4mL/6GvCdjZ5Ovobp5Yt049o71Tt61rxLJZEbTywJUkgwuH8fKlKnW2ADYmY3b
o24zIFM5ulFZxSsHVE9Td59kpu6vUYn9iOurbEbSznEq4LVLPN9Xzl/Tvan8kp04PPRzlqUv3EKh
ZdcoaiogeeNCWal63LVKFUhUX08IYDZTdA+Y5np3hHO2l82hp3ANLROh62NSASzZ7brWqNjvkG/l
TfzWaQFcQKjfw+zNd2LrUoULSOcu+t0+Q0JOtdhPXyTcTVq9MiPh/GN8rWpzQYUtIdnHHADnGexN
U0jsJhdipJ5E9F3ZrM6BWOy/3zkYkabCJuuIi7wx1lrsFwgJW+p1sl8iccI0Esmhh4NtTbN7va/d
QE+CmEqU3ubj5LiKzWeaJMgR8KAUfsSoPZ6FK9eHcD3drM2M3FmXpL7bCBWjK6qiAbhL3qPJUA54
/VQNueAkTtDtMmxKROsdcI1yc6jF+fVqC9YiXJifem51aPT96DS4xB1+qSz8TGGmSS/YjrkDg0Kg
XjkYZEEfaSPzdngxlF3yw2FpDewfAgB/nQHleytmA7eRs0eXkUxbOEjGupGhI0ItXkWSEH9dgCGb
YUuZZmG+EWkKmvWop32votKfH3Rs0E822uTpBCpjOYp8ThVUx435+UbcqowkpjxC3uhjkbRQeFI2
CNG3wMRgTDOoX6aRpMV1DNcUt3V3L1VaVSRchf5S+P3Ad+626ZC5HQhR+7LzRG5+gR9+exhM8Gyj
3hmyQp/tmG4FgxeBPS/o0n3Kk6W1duDmMk6rxCFJOsdr+7TNz4swnDZyRmlGfpANTZHTYVnoyZwp
511KLOIutBqAXs2XZNob+OD5FO4+2NEawO4ngWC2IZyd8tgZcPvxtJrPcswcRA1/POxULKqX4WZt
UL2q5GUCC6szrO4yxB7I7WoSbF5ZLzEIbB5kJvcbqXmJriVkPFZfNra1trMM6si02X2gvAlMldPL
M+fGFR7hwfBlPaZqt+fO/ozBshIC8zs7aiWcvNC8mWIhpc4Xm74adNtf0v6er5EHtxBXSPHHYdjA
aO89JbVD3EhSR5m69zR183/jDybuMadwerhCU/+DNdCqv9cNytkakXKw2IIpe1PRhsOyLWHpvmHS
7X6G52q7bqoX0PxDdS/Kz8N9UUDddbC0d7RMVo+HpN/g6yW9BQLm5IjdeV7Z8I+2whAV9h83hF24
qZ7SC5Y14AqGmlSagIjTVPspK3xWpSqn6P4LDfm8JueMVA6xk3M9unQxj/vYshbIyqz4T+K5N/E9
tJDAxJ/1Dsb0V4m8wNB0yW7vDrAtTLORTAOQGADxjLrF+kb+417X3EHi1NP/SNfLBDIA8iHY+KgB
jPITx/a9U2Zmf68r2DbQEis3pMrjeJ6rCJn/BCALnaPf7sm9gEubJrnJpUzP0HoodGD0GGtV1Fw9
qlDZbnNh8aAuHzubd9pIk9wH9ffaz0H3vbGjemd8dBw36DnhPq7fB3Bh5W4PiTqXbQRJ6Dq62dSi
VM9lv7jqniDYlxYeipNpv0piugfr+Hf2L42yrfnMXsa2jOoRDp7b8FNvRio2TtO5C+wFTM9GdpVQ
vgosaLSU9j1NOZDWCaVavTAYK0oWgJDe28as6yie7jsjO4xfqhJFp+/wUqPO4Gdc4oMtktVnQ8ZX
t4iQYSeBUDBN29cjH6hf0MH4W5+fxydIzJWGv5CjTeM6gWyvIwU9aWLUNo8UJgshtTCbqs1nAD6f
FAX+WTzlwHqFddRsLQzV2trbmBxMA/68jEk8VKEIhpsY0ST13M6cHyrxZkJGlVQymqJsU4HI1cG7
lHU4HIPQaX36Q2Ziw5YHoGNy3eavCzsVQICnhQB/iYBmVFFue9xlLKtJ4sPO2FgMFsGA4XFPhxMt
ZgG9bWURve3BJjPMySocQ6HUkrXk66qYkgR6pTaUOU6JcL3+iRkL4JFqxiJ07aOIZ9dgirVLGFZj
4gk0gPSb/DINt4aHrVDgxUABDcE2xpjrxZwCd4o2EKkKAwHsT2CDDoBcqCPrO1A773gK5AMe+MHU
HN/ea8lRcvlCv9KeY96720lV4DEkLBrqSSP11LgxYoIc4JTRYJq5bC32oRcnZtau/JN+Sv+GxA7I
ogL88bps3G5bfWY2WPoVUVU67E/wjQBYyH+2d5YKnaTouYwgdduAQSsGBtpje7uJa87mYtppfGyW
w6/h9G0spu5IKucJjQ2eOkiGTkwJKvjU9/0Le8rDrKnp6510LZl3StOJOJm5hl88nMOkhJ4qj5jL
JYEGDCsaexw+rHhrLEWZRzRnz/dKbE7d6UtnA8Txw12rc9yZ4jf4of/awC5qPxud9SpnIkngGi8m
qXsVfqufNyc7ArWe9raETBhL+YWnZFttICDrHcV8HO4EJAzlu5rHFJwR+3J6xHsw9YKUq0FZrQbn
7JfDsXwOo9Iyx07TiD5hrKoK8JctROnV1CvMKfN7C0elJ5woZ+7yiexIzKwiDjpwmZamUrR1ovb0
x4wk8fgnhNU4OhMNuuqUjZLT1TXizKHDsojxGpaZugyvA0miMzbP2lfeRYIAqMr7+f4YY8Fu51+J
o4/5gRJv7UEHjjyZ2hW3JOuRiYeMSv/It0OyvcH75KgYDQZBJoKNO4w4mFOKPUrax2qoND47Pfox
hTCgULHryIjnidb/g5jJcvuBO9Xbndbj6S/Kv2C5RyHNSmw2nJPccQdUqaMKpmdxBoFpeeEH/4ia
q4doYY0Ou/j3pRyJ8vCrVVrwR1yB44ptRu2qQjbkUVCr2MHlrCiJpiZy/WpXRUKjXUWAsi8UJIeQ
NVfKnajvIeKCkbVfqDkKCC4Qp+5JiuVoo+8r/xbqn39HmK3nDrFogiR803QsSuAN6Ha7NUu3YvCo
LnUq44XitsKSju6luKocgtJxVkzxXKAX6Dvp0GMXEgMPWUhvmM8HcsAGjf0/Qnw/nbRs1fLVrLQd
mwsR028hPM8JmsTkzN/fKTyADZuSQgpbIqBGaMDe2/tVjnLrbL0fl49v7SpUpqN59LObkyjjx0t3
1ra9rtjscBw/RMz/JQH5VkS7VeM7o3EMo0ZxJ9ReST86W5cD2JLYNA60EdVOqoJZ2Sf74narAglX
H9CLwtudWEx0sMNH6nDLW83ZgwBmW7gM5S/W03r2OT/9V8JMakIQ1tsgOfS9T/wRRVbXTViam6mt
iKctgsX3y/9ANItxyYHDS5wHdYWY9Lc3W53BrUisVy3f3MMLa5b0I6J2J19YHrKIE6oAjOXTp7qO
D6PiCEIoHPIdECPEiQMpCFxgtNvU2GPjY4Lqq+65mVJUCJKfqRE3X4sfTi29jzcBvJ5TT5x5319M
8kR71pFWkW1NCRz+Q38fu+Mq9ydNpQpuaKPPWgwolA17XR5XbDd8aptsF9KEFgbyG4t7rFkqPO7R
sm8oy8GLKXaBTvHUs7yQV71h13tsMqzdnPsC94VZFNFIcS05G85HGXsgKlYqI9fWHMxYP2BAWKbB
GdsJ3YzCyFT4ZK8oanGU9HHJjDNvxVnfgp2Gq2RH50tUh9UzkvZcdZ7vSkcjeASvtD2JATTDCbjm
KydKPK1hh+J2IAn0cOgaiT/vnkKVwehjaEQZSh9tZAmJt+RvoluliPwLzqggbMtysnDJVZ7eyJb1
P/pgHbLzV0K1ZD0Ro/YtPXbPUN4Xq/h6pWYNGEbf7UwFlV6vaKcznKiL6+JKgq0Ngo7N8IRXE4Ih
1ZV+j+lV3rXmrCAAaCyqwhvIlpg/nJhBsz+5dJGm9yoUm3zXT1te73exMgF2ljVpLcJZIdcs4pHE
8DRNxRpUHzbpJVaC63mBnBMhUwF780FMHESVTpk3YimZc9cEma8u0+10hjANTMo1xMP7M690qgJt
STZZQsMyJgfhDMC2iv4i9Htjm6cgpG4SttI8UHzqLQar2vfNJZ8kTBe5S3L4x/tQWIO4T8rpYVbY
96/WfaZNwUkae+Z9f5WsUlKvT7fLrZxvlkidhBwkm+jCVkk8uNccj/H9OU9ZfRmgOvY2j7RfLU02
FTYmeK1EpwdQfuURgeR1gm2DTLxukNmAQG4yZdOX5qcGCoMb8VF21ILZv3//ERhX9Ns7pJdLnJl/
rpx9HMJdbdaDBYot7CbSgv3vjABIjmPIkCNkwNNqEUlvmghct4Gb/8ORo1UFKRcPVVO29Jn7IWZc
Zv3R4DgjWhSInhvqAWcUmSSAnU8+X5lR3sFFoFy2ajonN+tERy+fTHmK3hx3nYCbogtR4cASljjW
9jA3Ovcq0NRkahN75cLKFcckoGjW9PWgCXFsbK46Mu2wgQCca9CNovqIHvZdn/MneQgfr/88ZpBg
7sX4lyigJpDkB6QOU+cLmD+WGbmMlCZDPwU9P+XC3IamteSmZ8nuL1oqiodVRBVWhObhJVK4NcwB
129t15+fADv73BbGZyqc3G58NW9mrKUMS0p9TWC/J3XKByq93UeKZAgDnvYwfDdcqeF2MPD1wZ8w
KLiOhAXZNFVchTLFsQv0COiJuvtJ2QrTxmUSIK7ZzNKNwQedBctZRw6iRcuBfwqyIxiU/SRyVJlZ
LKc45N8q9XF8jAFLzJuK+wzxY+7qnVMC/hxnis6tiiRtOiUM0OVRLW5ATayLBWp2D+FFUZhfxpVY
pw3JRH6SM+5kd5S30I5rJ2GdEeUoSSIgw48jIr+h/YP7zEqm7igMxwbTc5MieiSQpY94hgnpnhd4
g0gsBQXUYyPoaiskEbQVbDeDL03yzr3hE3nCfMJ85YzqV3qmZ8fFnKmh8/PqsJfP2LZx5BBQO6VI
buTg5FDv7rY1xgCr9J8d/7G3pC9TRKy6o5hZxLeprhhoRML4DeTzzp8Pa6AHSOlT2ch9KneNxZvR
trYHZDHtGbvKG4B3YCMN2vZcBuFTI4Ku9BunUlN8nAsbogXEO/IlBxbccjiXWNm9oc0luYHdUhoH
UHS8FNr/6FId1YRHPRWLkY7QKoXk3uziLLLMUDFg8zmdJ+h7NDX18w123AZjWoR3gMKLDxDN6uc+
H+aYgUu0EOlrY/veHOtD3Wgfym8erPE1vA7QjKrHcDKK3QCSvg3LiSIYhJve2KBm3crnfTGAsNuN
o+SstshfB/Hi1SO1CUzgrsFozkuEDu4A7Nzl8Au1hklL0ZegY5P+2JIFiErfphRJ3HV6qxux7EXo
4BMz8vaBO5RQ58KH7n9KpEIuPIBQZyFUKk5sU9/uoDSYdsjoqpfZgtsDUjeewpVJLumV5uT+md62
o9Kvn5sIjDnQCGmUTltujxB8Cn4uhGCPgAJpe0IjS4AeX4JQAW3fKn7HSPjBrsmnR6vdDt7ot1fG
71Md5RiKvZoiW+7TfLnYJd90HrIQudleoDQiFlH+oKsOCJJKDV6jxpIRYDXo/8QD7X+8+8tB8zTe
QIxJbV8E9WtgrCyeVsVJAK0KUY8GuWYPmec8AIg1HiJjatL7mA1G1Waqh0WGe6bmPKDjsBzvR0dh
GpeRsE0TmFCbubw8uaYMheunQaCfY0CDFnhWR6qCDIUsVNe2sKo6sPJNLooDrvb+3A2izHaXlA1f
Ijre0Vsx2LwQOmS8+TBhqD6Wlz8GNorDSnIm6+lJfb7FqTZjspt7qlzE611nGMQ5Vn3EyYbEZlW4
68HKi8Efw2ytoDEV5hNbHY05m7ue5ED4SKgxamlQpZu78dmyzXMOJPKRlxKQLVeylNLfBf5BGlWm
Gtjdv/2xpRCtlu8uQMIB7MNudQ27YhZyteKazx98kbOzsbVYR+ZyFY8gnF2jjetzfl6Hh26jU3Gz
JECXdsCZ02T8Ti3xLokgjItaxnjtuLCLaXxC6mb6BBae1+BJLoWQPMXFIAEY6rCHQLJM05/TgkqK
TOfUCABsBEtLxR1zihhUTK2j0vXxBrB5cpVx6vCETNYEEYoks9AwrBif6FcmhGE+kqb0DX5wo1Ir
MBG6v0JrXjG6/KeHtDsaOt/NaEQA9T0JPCsW6ALT4FnCWRvsEkwohjTGwRErWpMb7HyWtFtPne0d
4tb16eQnFi1Vs2E4BUIqgsl0zVKWoMLgHKcdpMg5CugUCKxLm1S7O6WMffeEgwCoE/h+aaSFJDjX
x3gcPdZq/Ze45UmSVTZ9aS0pcRgHH62DGKnrCWYTY1MsHkgkjs4SsHN/75MqPkOhz3chE/+SaJFY
hhezjjeOUehO6ltYnPNnREgpq1Nt6V6D2GAWGIQzoctH6Q806Pl5xHdD7FTT3J6Qp8mBLx61D+R7
CfIjj2YR/9/2+MJoEhqrfxJ2iA6cKr7e4XejMrV9eNSM66nog2NlEp/VOWTjZVnH0GBMvKjaTyth
wZuDFWF6qy9sIqq5JEMmfFqmYVQ5wd7lTU9mak6ZIQcBpFiwN3MbYm70y/sopCTEmnyHRj2U83HD
wGuHxmJxexRceBUQWKCvaItdnCAtO9oQDdRuLeSddl3rU0XxLjcKKco179H3AKrT8QYWslXxssAL
UqhnMpwTHSsg4Lzt6GZOoUZJvXU7Xs5uiohEdqL9RE0ocg7qTB6/F8fNHKN88C4N3hfXFDR8NGyB
8xrV+JQfjNkiJe/FAuMW3BHSD0YAxMxzEMbJMx3DtkCmdMH+czQlqmid4SGXpIhyr5PMxSuORpeo
EsKf0A1oU+D1fntoI7QHUKzZ26n3VqHbuN7ZfOG9z3T1siGUJT3q65x6akLPwlOJYmhXtnba9hWc
vhr5iLjqpmR0l6o1rLu2cy1FtXbiEDbUutC9MZ9KhjUqRfVpToSv0nBmQBFr8bSvBDaFzOPnwOeU
Y9ZLSp41swDe+TlO+B5NQI+h3As91GfnOp8akmnIE+qE7eYSHVOyaA7nUdEdx7pxNX3NAFXcEgp0
0Fd8S0K6N213Djqd6mB8+Ple4mPj3cju7U3tOLgu6ZFZhvJoY/01yiaCrrVwx7Hn/HnUci3p4HWS
F609O2LrZ2UMfXG2g7u6TA/OTvKvDlfX+QCgSz0JXAn/xb+KtGeLOqrQkLx02wNl30/uFCsy3OCK
JuiwKsTi1QpI6BjdcRIvmS6qY11E60uEJ5MgWpW2PoA0DY0flm20/vhQW+0eDeoEjsFbJOKs0r/B
NUC7Cbl8+qXaxkAu6hVAdGffofzxDjx+lWAmuPwELtkz97Q/CnMG6Js9N5mOSsCDLPelqtsvKNyu
EgPVV8IRuOznkyLJd6ohVRC/HMSJqDxOHvJMrCKSDVpSNnWhRD0zasn+l6kkZGrFqT8lpRDzAiKr
mzKuSW1GRoQiO13ek8MrtOS8O/8huqI7wg2c49GgAEe8S8SQ7uMDjYQF6oCTB3NgR8nJaNOK9LSB
+AbsSYN+DfYXUnI0vIVD1qXgbNdgOSbeKnS+UwHQh8vkQ89yJFFB/HaHxhnEJdx0Mnnz7T4gIk7A
/pMn/EM9oQFUgWD56JDiFzzjRt+TuMd33D76UOzXS+6Yh0RnL1K6ouO1/pFCiIql77e9EHfJ3uZP
xQYlJ/PfXDro2fDRNBuVvja3N2hdcqJ1mUJ9e76KhQgMWMn9ceeic47EKWspnOURcW+aGdyXqKi+
FLZshow+EgaI6GGl1kMDF7EdjqPB2dKu5A2yANeY+ZHWyBomasG2rLZf2MN9EeHjgBRK4kFR3ql5
Nu8gWh7CsXK5lgR7YN104QRrtum5ZSL5fQnq6ycWJ8GfTcOdyu10fjyjhOfuCDlUam9jtdKJatLJ
X5lIUiWBaZVQNujCLdX+SN3G+R9/fBMc6UeYYl+a6mB2uMExlgsAIVQs21qtv53hm0/MrSRKg5z2
oGJZ+4HmdG9Ljs0Elxul7u1bRqlhKeU1C+SId1T3FgwPrG8p7Y1ZVX2SaqlAAOUvw/tTkj4HCoRJ
gsEVALf98NuiJZ0aNUDeMJqK3Ka2p/MBvnvQpMhIlCvMjIg1vDX6zxvPxIDAt+19788C8vPnhEsa
+fAEm8LhFR08Kbs0+RJ7nTNdHDUBaKuwM06ggsGvU9Td7dYmJlz/Nl1pKCGR6PHeDjeVCI8jMFqR
IsHNcZkDGTUWg7+stulPyM2wt5P4KsLj5A/shf8iMKVuX4AFsosMgkrmLbrliN5frFWIKbHBw3OC
WkBPeng1PgsaCdH3MptY+yuH8t4ZC0XwubG8/ZQIxVQiVYYi/voDqC27v3/poY8jN3JQHN5ubcnU
vtJsY4HKfIuTyElgwXVCzHym1S6LkHYKCvAGspcXUaWHzM+72DEZ8bP/wx/x10Js115HGkHyCp8u
56k427aYUYINsTNJZMJ20svclJb5eUFY/APzZijcmPChR78eT0NPXQdRoyfoe9I8Zb61O+Bm1yON
jyJjUbjB3M1s9p99eF/4KOIgkmlTcbDSroA81Eg6E2S+L57bgdscbdzcJrQ0XHeJtZtXqHsw4qbt
3cJ8S9ph6It6Zq8ymmva7QQ6bFzgXluWdCunmgL2CjyoiBLqQhbVWpQ9Y78sEiJQgetzWhkCLdkb
hLk4seGpz8FtlJTxaXZk1sejvioGAz9x6oBSBzraL6mZOfG6d0pepMxmMkPlqhAbHZKv5CYadqBt
d2QfxEo447h6hxRCpHG8NoJIM8+ryCprMGn+BTgm3ni+pCsl3hzNxr10DRSoMRZvcEYqDm7uHQ6s
zmW/C/0tJwnm5QCP5dms+DWnvtO0gXyoYhdnZkgXVGTuEueQS5u8zdXfYRFF5aC0yVqlTBiGe6VI
U+2l1PtgnnlYzFOLx9V3dMNZMzP4MJoiGizM/LZUKu5tmTqTZPnffFn5h3pv9zJGclSg5A8e/bxM
UDQSF4H4JmgEMuceQUCWUbgoAcJG2Q6Ha93wLm8c7Eyc/k+AW0XbvWZiQclJlk0nILI9VWBaZdrS
xs3LYOlSpLiTUPyHhc/pAE1iePwoTVEO0yBClDiAkUWHQNgJ/ZAwoVegmPL851HC5HK8b1w7Q0sm
lAHGZiMyjpStSHspQ03GithOMnt3FkK/0a5EXA6sMqSf2VVGPQh0pcB09R2dpt3SIk4ugmCtbI7V
MUKeOE1q2CD7+wzQUlPu9mj5ZOJuCFbYGz9WY1MH/+/o1N4FaP3pTGj3SCyqm0vwuhWqI0CR1moU
iuf3voLwrRPIP5GxQRXW/n52la3sYdxExR/l0fyJhKB7Ak/77CExFY6oxaxZr57STedpdZcTUmoW
K26dJUpwALH7QCqjiwv4jD3v2stXFEWqquhQPIWwla1k47hr4D2qAyqaKMd2Vc6b5sV/KHZ6lLen
EHqK3GxKnQxoiMvD9zVop8psFHVBnwDW6fBDmmvaJSuUzosg04F82/w2iCLtHAXBRQcxna0r0W4f
8uwgKwuz4T4t6FTESZev9uRFrf/Q+WowFMwmQXTD0lr6yneo8WIXJVE2jwJ/Id6TtaMQJR/AR+VY
GiIu5GvX4ev5oiq660MJeSW8GnejzQdphJjCUhWIwM4hdcV8aG2O9hCpm7dnIA6C5PvtsFtqqlZk
Gxc7gR2r/38u/rFFq10uoo/RSyu3Ayk0PuQxnLBH6OYYd53xEFvt+IXl0/1vnOqqeBhmXrH62L6G
8m8oYSXjGymFlQdTKgyrOk1RQCnll+jQ/iG8OjCe+hQV5eanK5eCHuUGv7VKoCMbbbvegDTmfDTM
nZ+Ry8ZvFtgdQJ88QtG4FQ5PKIdXwYflI1yX5JtBFuYsfTHP0+kBUw8GPj9/Z2EEWM6W6ffP26m7
Cdkkc/4sEelxwfXQOPr06HwdFR/hPsN5IipNCY0gVdT8pOgz2Sq19RTzZfibXrCeHL0LsXecl8xK
fWt83mgKx5Q6cDuaZbI8wu9krq9FfliYtpfPseepKdIoWWy76Qi/bPcmG6uqdF4S64XxbM0ekZB4
K0ncPVVTmdtaQENbdz5HLTy9hFBKm6VwFurf2W4sad08p3Qh/hU7jF6w4cW5RsNZcT+q4wgnQe+l
HA8UEM8ooO+EwXABktv4ggGONYbjOi/t/m2Se2JkVTzwZ4pkaNBDbyt3z1c7dpxDPg4dGnOEPU0i
Amm0hCWAV+giofngs0O+Ak+9kJCzL/GLSItTtU9jlD7qB+rQqDka1FPYJd7Vp8ARS3j3CEugne/H
jW/olaZch18Wc4AfQbao+mkgC7E44vlT3iOkBYjy3FPgCni2s8xkOKdWe47uefOLLRIYb3M25K5h
rrcdovkJps4k0f7AXPKPEdXom+nGjoNK+lIcg3y3dx9pQF8Q6qpghEi8j6Vvsej0p7AQ4CGJRpg+
BKjutXg0dWguk8jRZqGPrMa1r2F6ya9UHUTjxkns86BTZA5Zvs3mtjGgGTbGlQfv155S9rsLZxEj
InTer9NsDRMPjse3+xhJVoDsY6CGOzOfHW3Hx8AgEKdHPDsA6fRb/xI6ycu74LTpGBoLE/s1Z6tT
y60tYSQCn5Z3zHh9+k03OkZSF7f1FqwU0tda1pv+QfcgfZEJr7sODIupUzFBs8J6zGicQQX5nAf4
49Cgm+2304KCzF10fFlhUJ6aNYYg0si+NoREMAQkQVs/A9uLaT4Gst78DJm0L3KuvtVyNl51LDZr
WfjQx0cjzMyahu/leZQ79RIwpay530XreRSXSMsR1cTrgEFEPLCjSE3+HM5/u2M0cHxDQdMipkBw
cM71egwWYWp/EZjf2rCZwkcZvGHZ8WF8QH5xGoGcUNi5ox5CsXRF3GlId4a1i9wl4+zFmMfZ2t9y
AZLS7o9GRRXUqoMVx8eqvDpFF/rRf8PbrSjjvHYEw434DqQQbJtjEvsgxeWOU19Thw/Ox6MMuBGm
MA59kMdkDWBXsey55r335k0+HmN7z0QkL8SeaE5h+ooJR0OUcztUsuYPOE3jKrExML24yoj5mLbn
kToSAWZfe/PBkOuxZnZFrJQu8vKp8fB/DWDlSbhp3mSdgRT47sQwc5zlIAf6ZltB6rsTn/DfPShh
ITICq7fJ0gnlY88nbGADZdRZ+IoTPDeXQDTf/uxWt9sMC2K7x3pOeoQiRXBGOdOi5htCdKGW8zEH
I3HdsfjASNY1feVJ+BoVSz0j7n4i35IFwLLEJGUdU35WG+haaF8lE+cvWYkHmkXu+n+dgmj/wR7u
H4x5uS3OzEAYAzClunBx4pfSj/o99d3PPfHzGMDHJBkJIaEelWZep0pvXAWO44uZqihEVYds5W9D
jNC/sKIqtAzCGg6iY9qK8Mdq4hDOZE2NwIXmQkj2Ip+BHbHcXDjMnW8ckbH4E4GJzKmaDRna+L/Q
mXY4SWQbKTTcNpXyoXJZE4mcXY18LJvSnPwYO1tO5ZWKL7PmVuMyhm8ctBJcB0vL7GLIGPzs4m4U
N9LDmwPFXkhyhl2iBuCOSj7AbAqrjYCZGLvK2PseLXECEoVZrkMcUa67hPY7ZoJT55ed/tVapk5C
FsFuMIklNxzzmasw4sVHP3XmbjXRz1VyxDmPRG2NBwNQbvenpEzgGTAn7kFXNAqbA4Yy28VDu8no
D4ek5xyMMhp+EmtiDNYTDPkrhV8KvCrx/UBDjemSFw8GrCbwm0ZfJ4efSvhGS8xs07m5OGiGU6Hg
7Wj6y6Z4QVfrpmcZpARzw2k/yiF4hbSxk1H5ekdFjazAcs9YWK63KKd5UrxmX8HbpqkrDNAvpeNl
CY/44PTqKY6NAnuvRmheqIAXeOHgN+0spODtCgNDnY9w47nBXNM47vI5cpp0/9F1EZHauOkZQWwt
hQ0F11US3S7Sg21kduMpjfPgFtetyL4ldbjJ2ZurvV3WzCpwP6TBpP5xscB+C3TBxBiEmKzBSoLQ
5fr541/aagGwJs3djtgo4/Vup6oM/Bfy8DpoS5hgoxuDRShROJQMGaC1WbHrOao01TjrGYHhKBRZ
PGSfTR8jiTzZ36W/YQeTtFQCB1d5nyG4EOP7klMn7ZG7km5p3UdFSqVX9Go1mHhGtBMPyaiD8utK
gbSoIoIR4sGYbkO/1ZQJdTZPwIyQgIboyv8ULeRhO1XBRJLaR8poF7awTkxL2Ik5NJCdL5PIZSIA
PhOYBZeM1Y4C/EkA6QcTDDG8p2PlSsavUYW85n8pQxVeCW7LeM2MTfhNYMNnk2+Y0/D2gvyYx0jG
qbhEXMsk6WK3cMB19RqOYlqsQB10Fgcho1WSzPYx+Ixkprns/fswspimuf+6zvnY2Q2ajKYrQ0p9
zT5tRnQvc8op1pTpz6OOpVdKFcmS7z6ATtks/p4qj4HreCrOHK/Y3OQghFpdUGg7jcg9C3UXYLgI
Dk+EAc9cO6kT+nroEf9GdQH0VoXTRY+2CQj9ZGF29AsUFLsMroFobB5vH7ba1R3weGE+rBVZNy8d
BJqqYwEOXZjt6Uza4h5j4j0LDxyzj9apEYItD+XzbwtmhGR4Qyqp7nSJLfnl7diClltb7cBKtwBi
zQuaPCbXVEUnVuzcpFJHGkx3Aw1D+qIPOYo6iDDt11OyUlBDY1BzeCLg/7pSPgnxbdqdUmMbeas2
F2Cj0e7hin9C7k/wZKDFzcQdhz0ughSc4XPpDrN+XlMLVun1esq0+U/yfLzn55ZJs5LEVYP+ZfHA
XPsvehb9XbsEk7/FkZ+LSNHxkHZmFtlQ2wK1WMzJibQKeJ+tSxQR914jCGhPps3FVgVnNxf5oAWa
ViaK7HJlk31YSQhqQprHe086/Ve1I1BbruQDL2BHiVyoVyT5rMSGm8ja4Yhg9JW+gPpcd7VTGmM8
mTNv0EqsVQjOWv/IT2xVjS0gkzFcy0KJC/K/GKuVZWK7cjYMjM+GBCQL04B1gpM2YoLVOirxeE1A
77Y4ZTwzxabYZViakJEh8v9BGHEIzw+OwjziknOwzY4RvXBlPDtyQ92+9LBBMq1N3YNVCR9U2qSM
Q2ZBplq5fBsWyLfdf//pl79z4m4oKd/6LgOjoKG85xQ4l/0nDRPGntYLG88VjcbLmn/J1h66SPft
MKB86SBKM4xI1dr954Ce+5H1YnIwcbSr/HC3hqPpovpcUCMeLv6NN8jfiTvmsDCBlihwwv2FCzBX
DxjnNXP2sg7tOo4JYkCgsknIQT7HNtVXwVvZgDd1VOjkvINDwZ1qAwzpY0J0yhKPlbdlxIFmXN1R
npxE/UXhvYESSWThcFhVtKP8MKJTstVY82eNoAz3H7Z4h3ADkPYJGp6HtzGEixowgi162kTTEgY5
+E/eyxQzER05cZXVe0nSQCv4oZivpZYMFyAJf41JitspxIm192+BY0AywQovQjvYCL7RsBxhXbcs
wUYLckZhwcS4Im6v2M2yLDyKUPCGSZy2ajvzmy52A3kC+kpgNvr45aCSupHJxTV3PLIwzZ/GHUI3
hF5FZtpkjkZpHgzluTNS5ynFQMLv6LnKfPnIFbdjWNSbCBqINenC0NoZogz6CVCBw4D8r8i2yKt0
wfZOTnx6oUczCrDbSLFoysVUbFYtYZwd0NRPR+DAhe4jnBouWQJ62oG5rdnHb9YZQEgj2NoiuU1G
kqUYKhPnJtB12v1KZyVMjy4smGkEjddjJRmt8DAwBMvEMt0ePSASD6VqyuwggszrVQjYRdiSgQW5
k0ps57TvLBaaIXd9P/Hh+QI6Tb6A8gSrnOGOcNED36mhLa8Y1DDUdxS/lh7Fz5txJPzMyXfzvY8d
qtwVuyhkpy9LsAJrmSTXtmEKN+GWO2U9GrUZDTt/Y/UPj1OlJxwTKBGuZzGdXZsBc6ibWMXfPxOM
u93yOqmQGz/G5vZIG9ou0aGPPzCOXh/RecGF1b5c/fp6Bf5E0l5cOchLmKZcZpzxLtVI5u+opWV6
2fuRt7fmvt3x0q00FR3MAiS6LuzKpefVTYHA1KuKvzeAMr0Rv6+v2UCGc16zHAuh3oQQxpXvyP4h
d+HcP36TNzqGHlYdzwyXd+ak/ogyt9carJnGcVtrYUe1gfCdftnCoVsxzCUDJpdbcGQjwFL0WXac
/RxE5OZZX4DXavQoSHiq5fdJivWM2y9Spcx2TpqNr05no/71atNzfWeZ/oA1f2hadykl5Zb9ZKKL
PL0Ikr7rIg5I6cWWDe3UzgCpX3Q3z72UICcn6vAyst8U/5ly5rVdgtyo+PXQaAfKDOea1jmSZlDe
VLO8xK9Rgo4YrGkbjikAHaAdY2pez77KKhp5A6KgxEil7GBIhXv5Gnv4/Kt2PwcEjfh4swdMQM7n
cdvRZLKrYU11g1KuCXScVOXWQ4E8PKk6RaS/eH1rpkkbULRq7/hkn5LZJ9+r+ygKhYO5WmUJ50fH
EErGa2KNd1wsmy+H75tcqBBS6U7xq2Clwe+jVzDzNUj1wN0kjXH4szeXyp31iTvzUDDiqAmcbHlj
K7OSGkJnKF5oiolk5fNu6Kn4Wa58+tTQWejqFAO4/2GrOnKkOqJu+exi8IkLMvXRLZoGRAvupCRj
gNAMe7NWQswEd5diGHiPJsIEDkArGn/ZxOyXEh4yBJW3hkqQM1rb+NVVeXBgxsosUB/4WMfH1Btw
w8kqA2mLSNzKkvtRLINVW+OC79g7nELLu7WTSMG1gjIUsA8ilocri8AsKz2WRl3CzROVWegL/Wu7
L3bYr6Pt76GeQOw83YM/eiiFtQwgPHaQhbllnvMvL+8TnlBMpbEoG+hX8tWNRJ5MiykthgFTaY6c
pUfh4oTbjUgNLsBkgq8jbMaGF9vl92HAUZQj5pWjyj3HUBQ2BactSGU620KHGJea9mVOKJ91TqHd
Y6/w4oAiRRLvNAzllMqok2bzol59UfSCjdJhA+cLaU89qm45oJNFueVpILD/OtUXd7USytMr+8IP
DYGMOlsx+pTs7XAtnZOrELAfAAvkU/MfbMF7GG/rJZZL37ZOSHEJW4WzlzrFGwoPmHdOOY259pJL
v3OJo1zV4ugaE3iKvYqbHIXrlsSbRzQnwv6ZDVWGIt90NdjIZFw9BrwL5G1W7riRcPWkOJCCwcLP
EnktPfbt8ero0cY4nKWJ9VpfAh2q0aIgt7eWEUSmGp/qy2OnBzQw76oclaXJpQQpi2yMN792RuQi
6oGAvD2fYSxRQUtp/XOJM7zztrRY8YE/jYBwFyyb1H6jxQQlWVFXsQfPmB6DGJa9dgja6GLbTTP8
ypi2i+S9vHxWXuO3XtsdQsTpgbvDJ6b2E6Pl87zeIoJ1rXUc7zNpDYlhKxdYCDDq/9TBg4IaCvE9
YQboB1oMccebQXi2hwkg0hv0yRyoJXnlnGFbXQa+EEfUkOccRRAZD5IFjVrb8xZvu9Svq5ugFmOm
tHPeGC5ZEdzPEyZQlzEjwcJcwpCQKIlt+5VvHZkZE1xv1gedTduKGqQlX+DoJGg3w/vi+3DaAO3z
Hn4hwws2R5hcae26oHZbCwU3Pufr05xHH/+lGLdGCTAu3p8BGnsF9qldRXG3ucSNxlDupoWiBNJF
Hx5Axkf9/KeemirXHGCYw3tBMHpvlkTySVT86lYdwkNSFP070huit9cE7lCdLhkWCh4+1ReDXkeK
NC+otYWNSs+nRDdeiQH5ktOisw/lDuX78Hje59O3zv71NoTT2zhBFPVHy+NK0I9N/DwQGNgmrkgT
+bp/jvZxDflLIbGVOoVbTc9or7Pi33/RNZmE7JDJeVfhGSyIAoiBHerG1yDOey7NLGSTPagnVpW3
TyZIdBe2oTxEQkiU9dHf9qxOgPg5XKAS6E79CKe9MyM+TaF9+8wI6I05y8z/peL7GFwIjdPqa21I
ZLFkGk5fao9wXPCXP+PyekzQgFsEehbN9u/NANENwaH4BsIMacu8WAiqF8FsQ8AshkFOQBZhT+zm
5h364rAahgR2ytgzpZJwXDTH37i9cov89yi9y7cpzkkUmvHuLSh+lnQysMS16OJ8KXLXxGonyPTu
AK2MNXgk0grrQzBeNNVN5jkfr0Xg+uGKj90lf97HfsVq94aokoZn6HK1QJaMHPYg0Pl+wmXSRILs
HtsrakgZZfFANse79jCeYKkUoyP95DP+Rur/NP7FQvEHcUBlwkyAbcSVyQtEWc2Ik/tH7xn0EFUo
fpxLfH+OTC4rbs9ditWnqFiVB+M1nIBg3Droj5SXPTZNbnn6T6kFM41ANdt9hZAqhkH3H/wHvx4n
TtTqxETw295scJOtJ4V+gxfERcJOIX9EqAzD+ggDq0DKlTxvmJ6L+Wc8eGl2Hzqxqh0EVpYjC0q3
jrij+GwEoxGghvAwKu1qppz271JCF3b3kgasDfURDaXjpuPPokgKqihUICVbCwJ3rz5NeR5ABMke
sdWgFnGPV7MQo9n8ZRYNz7FCQdeSLwuGv6glglRjYg+tqYUueiyXSIQ31OrmdPOT3bZEGnXrxUC6
KVk4AAy4r3lgfOiyiHpoqN07VvijSqLQr6Ylu2NqNJ6A9Z6/iEL2LeCaaznP0ZmDNbDMH7naPpd1
MfLATH6LNErsi7QQUOQ1FgLLA8cswf+KJX1KXdrt4Lpx4hCdLkYo/nCIonA0YBQfX8dKirWfcWBn
C92HNCIw8wpcFcOUxgZ1rpsANQ/4uCWFxloOqILyiRBNyo0ijIely9aA3V0NmRFTJNcfohKMkiiX
7r3zMwFmqtpp7zbpMaEw3eK/wCmBQ0T8BjYLe3cW7C6E7Xe/bvt4kB9YQ5+Ggf0LaDZ4xYWi1eEV
heJuk93zjR2nqX7hUWOpsVPkBsBppJP3t8OfoJe+HHrWbqyBx2+m81hB4wIm0JsWK2wbo/uN8ERF
5XfSPRg6Il0KPoHu6UV84oj5oRAxMQaFwXPjhc02LUtS0RhQ7Su5201hczx+SmhBoRkVNPg9WQX4
VtFsvrTBMGP/w8oTL3ly/uITBmsHWIrzqd23tfre4n/iVnfPPadZDvBCG5TdSdI5O2gdIO3MQyK8
9NF9PNvO+RVB98VTcfoPhzlCqvWTD18GSCZfcOPB2BYo/ZqhY5jAgKOWolIYK0r+pV2O9fCmYbTH
/ai3J2JJyZpNuCaGin8gw5B+e+5xbA5WmozVt14gGAcFTcGsfJSEqo2pwGCZqRz7DOBmcTXm8Ek0
EjW4knTHM+5qVIk51yQK2Zo1IoTnK89PPEXuiDVV+l4DQi/783HFdnFWQ680wbRaWcI5gFr9MOe9
7zvmHpSi8be/1/h0eEuJ0Nas+d4AELjWtF+Xl7YXeVrzitbmLTjD/oq7I5VtiWL/lvmhGiOwzu1J
dif5WfcbcikfbHo6tpAUGKUHNM2VTNiPO+nUOA73se8m+bwdmZwzt2qAX14nSDfqwYbSXcOEMy1r
jF2KXurGyk4SqShetJk1ymOdePctyTJ39L+AD3uZyP9OxQjgXWk3nZsjmLXfESyl1T//97qGA2VX
IgAXo65X7Q5FNwspVIO6m1x2PUa+kIEsWwnrEjETiN7IirKObGjK7KQc4Q3I/bBwNh7K90De7+ma
8KG330d4fE+GZpkMXvYC9Pc1pRkFgBZKNROruhvYktCOr4HuwjDxCkmT3PkWL4d/WuyiM3XYA1mL
m+QSb+g2JVj2OIPDR0geQpwW1eckdNn9Bg2/YjvXLdZyP+JA55+X/jlSPk+9iz4Vl5hlV9849SVE
6RxcKTv9Pht7xYehdJmk2DACZAbiu7wOAR+SxWKJsM8c8AYrGPSfkQlb/LuVDvMQY+TiU+uDNnyL
x/v5TldxLXSivZxrg//uDLoRsyXKknet/YzETMxmHW9pepGUDtYcUVMi6dTEmU08rvpFMnmIJeua
GWqodW1S2EViXOdPIki09vF0DJq4hJzqCVuMN5MCU7Bb6YlTs8J253U5g8uF2C7h0VYc3XiZ5g3H
ntlriJvnS6uH+yY9FwYyV8EnmNe1eMXe6ZnBHZ7zjK3R1V34O68306ynXyklRr3Oyzms7oZOeZFD
w34VUwtNnhaNMI9voo5WA7koguWi2pwlhf4FnHPdLNzc3UjrsLQg6CRGe+1K4hz2fe+YVL4s7LTT
GPjw9CY8suHKaaq8G/kT6DJaoJ3sdbXuJRHNyuaaA38RHeeU57kIBYMc046GUJn12sM071sM6mzZ
j/ySNEZOmNtDO1YaSYmKkHlgebKbJDAIbw/vX4W4CBwueoQLqzQ1Hi6Szvq9/6qsUaziTQN5ap5z
ULmVAy/WwZ5u2hJy8PZRENQx48taEoPqZBockHxhruxW8C0nZorRHYaZ2N0j7wIr1UNkXpYc3aoZ
jF9Byj1E8JwrKB64Rm7YQPT8++YHyq2lF+O2qBYfpF8ETG4Gyvq9SZ1hVkEujulBP0QIUoPfNtgt
gnbE++gCYDBOFNbgMB0MyVMNejdQXGS/FDDBXB4Ky88jysroM87NicykgnU8USJ9c1w65pUn2ZEY
Cqx0RZcyXnJPZ2svRxATjNiosy55j/pxwEZWZPxP2W73uO5mX+IazjkjOGSBobf+fh24z6y6q+B+
WeU5Lk0Vv+drp6DOV78x8fDsihQfn7m3sjCQjErfkZxEkAx06KNW7uEVs9mU1dsqINLlgtMTGQqJ
n2YyKcTUldIjiPoHv3QW+TcWrCfZTtfYitOWzrMYd6X/5KUO1qFnuOOHD+VlAdlq+1yYkuikFtSu
vItOWNUMyjUADBf0AEapezlrx8bqveABJISwtKw8lZ9JQk41xIwmOFNH2/iMljjwmkbbafcpxDOX
OnPv81YW69Bb+Wu3+uG9dk3AYwHbYHsj7ZiZBBZBENWw3NPta833+6fgEBw5s858YkEzyo0MPIIQ
+mf45NLL/4LpFu9K88qgGbJmIANGZE9x+P3MwBxRcQrvDkgqvgou3RDzLIJknbQLjqyQBtP1bMLv
9Xze7h164x8kMiBB4d274MIRE6D0Ttvjl747cJ8xH1z18cSN2gDYaRkM4v7VQMG177k98dK55Alh
lYrbf429jKQjNACaITROU0wkVIX5lNZjLHDCAjvXCh/MmT2Zq8e5+alp82HhBF3eH3wR3+Otlgwh
h8iMaAWIKa/SJbwgpkoSXo6xwE64x815ILV/8BwxdR1SVND3us5Q4iKafOLdKN6A0j+qheZezQ7R
OixyIepURV6aKw9Wv/scDoYz7wPaV8sTokm1zJry8K9/gH5uhOmslhgDJSdACiD0MilBY6sdXf00
/hoWuu+u7o/HFTWDhvScy6rAr0WWO8oH8lesbRdQaRjPEtYsV4lbJ8AF3vhSktzC0zpHR9FySZfO
ISzyN/QMg4SlP4RZOtPgBw/9zRPHOBWUcuHLGI1vTzGF5UwSg7JZdr5i6UbGlwfUYxYgHqNv70SC
Q9sMKFAuwepBs/2P3xk2EJwG31iEG0AFdhMTNgjLrC/e6a/RY55WDx0VKP58Gr9k0Vd57CSLu76q
dasQ3IGVDIgaSbmuqR7WRmbJMIZfgE6nkD0sJY+BSIVYwzwUIN3xpLVeq8KoXQaDTDUCqZzZoIlv
VOOWyRk0OE1kNsinHRe73HXiDZR2nKJt4ik48LuT+n5UoQJgO2IwGTucowzkbtp2seJfxFwU1YcT
HsVY66C/7JMOoCKFHifXMiA+aIp1slgoaPcUi1k2EFYzeS96iVEFlrl7oJPDrVE1Tpy8z0PFdvLL
+aRtsJNs26xpXwjGwQR37llx4EZtMtdPW5t/8g7UIghOP2AORDYcXJFC7h5zCxYbv2eg0fhN4s5Q
lz5OD9SmtNVcj7YBIhb9dPw3ea4tHA5GBcToJI82Lz6Z/zlUf/dqvFmtYG9QlzmqSG6NlZ5YDzXe
WhGVjRrbJwr9Su9LOrmD/lW4sjwRzKeF2HzQiSpgrm+BrJl2aTYgEMxjKO4VhYbi9I/sxgoJVb1W
Tf3yYM+UXQbMP5+KRu9apWpkLb/eKjo2dPaYj0c5mz/D/+cmiRV3xwsN9eGkqpdSvbInhpIO9oBk
VB87jLAZw8vtTUdoRFxQUyU4OF8HEaEzdb6RwPIGbsytsQ2Wd0Th6HOSaeuWdTxHNOEf/9f7Ss8W
JaI6naoMB0B+MXKvTpcwCqY72yrNZ6320mafpyfwiQsi1lhtvwCZYQpAJylZm89YhtlXANyvVW2f
PieU7CjvmSJYk9YGsMafuL8eEtHKWkN3tzvzBqMp7u2ubsMx7qnTiLoEx/zdDhVXIZSmIIskKmqs
52wBCV4ykMXeGjHteSxakn+TesSUBfpwmF+XSU3eaM9Po379dfmDDplDtPm7r6XcTd3AV152K7wH
1pI5O2kT8Sf1GsBmf0x1HsKI57YpUjUzUO8bySmok3UM6M3WeqI1M+8jP8j/5seyn5Tko4iliqzv
cuDzuXHzDi4zgqnagyGeOc7uMQFxlq//VPSHsy4Ga3VRvCraBDSDfK5LxdeIIKXxUVKk/+wBOb3Z
WhvGEJyGnUWMcPwxdtYIKUItENerllZ0WNOrJn7XLjzn3sSN6cWwmWx90e9awAn2UoKz6WWdpRwv
WlJBMuB/i9Ck86Fs//XZ9EGytCJLvUZNYwuD3cBqQchjaiF1luBYBCpzUm4arWObr8KTEcUdWJwm
6UinaXUEaoP0AfhK+xTEJZaf7bXsH7g4YPRe8EW3YyGAIuZcXn/XV41DPerh+PScs/5yKJLNnM7h
as4/Tvw/SJgLPuoGHtr/ofX9U5p4wGztvhRwZJ9YcPvhX0hyj3adJYgR36z9WYelvDz8SllcmfJq
v/4aLqtx5G3ky+LwlIpH5kQVuVh+tvbCW8MCTrPsYxkEmMu1Xj1DmuBLEznSQZ/MRS0NNXnUDLxT
4do/xiQyqW8elvA7laUrWNmKvs/mglNti+DMoF1xqkRhiVu6GyTCPIdwSjWUsY4PdBHLuYj8IA/K
ojD6MiERX7HrGTcg4c1YbOlPb0D5rgjtoOhPWRjLd9AZ440vcAYmYTbqK7aWwo7Y9Ri/9bx0t/mc
oLA23JHpijKavEIl2QttFolpLrpq25tDefzQWCLuZXF33zETNJ5c0hPW9Mpv4kotG6qPgEllqorR
YwOFZBDkWh+X5Tq2NR4xX2K13jXjWe6Nq6LYxIIrX67HLkF0cx6BiaKn9lsyXXC4lgSuXz535DZJ
ofdGwtL9Ln12cK/dsmo6vOjZTsIx/QLMi38NdKyiM4gWtSYHGbxSTM1U8c/neSoENQvMTmF0kP3C
1p1x16nPAAW6GSN1JGDGFaWOEKx/wD9tseu81fa662QkDkkkl5zcjEvS12Norf4k8EyfBfI+ChAY
d32llCZb0GSJJL+C1shT/nqo4hrSYTGDHnbcRoFfl2ripu02UeBLBpS8o/UOsV5SS+Q6r/qoB8wR
ujNXoeoV7/v1gBBnz8a8WqctUywbnjaFFLMXPr3pRBjnc85ShrXmefo5eN58dwMU2GCdxF8RiGRq
HGSxj/zFnRbBI62hNeWMXpnkKnJasfgsuSc/3PzLfQ01qif5mGutiyWhip7AxqCXD2poCwO9kmoH
C0DeDkzbDVjYwzo14jPIWZLoB9kjkdXsJqnyvfIr3Urs7r7xRYj2cm/JZ1hfBL8SFKg41pgoZzne
nlyjfPDlCsxTIrfIco5lIv16WgLjzg1efREOmW+WVWgJA+55ZRxEHNEU/JVFiRscglZ/4BFaIkGj
3F39r48QapfXuph5uRXQq/k4RNdyVoKGXU7vR6zT/3qn7/K/FoePKkAMCRC8wvJcRkHYSZEGGH1B
2AQTYy2ZqkebWNQXXm820+hy2a9UvDD+QrLBObyUX0M7ptfC3nDBprGqNdtW9yiHZnNrrMrdglpc
93S85BTd5Y1spZbuqFUN0xLsCWXrLO9AqsKz9dBgqLzc3D51h50t8RgEIXRXjc/sKxJwyl3LGcEN
LRa67cLSn+QBbSkVwUaYQ8wfccvHLkZeY1X3uMw2MbPcNcs1F/hqw1xb+FT/H+J4DdRqV+jNoptH
Ls3mdPnHddAawuJN1X6jDCSLj9e2urrTk8z4qLynygPNRURbuP0GZIS5BVwvmo48vjieVqntOVtJ
LEMA55IHXDWa/6Bxyym9X5uOs2FMiHO2YK1VCiMJ0ROvQ7X87+eIeGdEcPh4Sup+YfRHt7FT2h3j
qUcrR1sESxVGbAeDqhvDJFv5mO009f5QLzGsJrmqOADq6udtLv/2PWn0pPpHf5Fmto0zyeoYepoS
+FsH0VL0U4TyTX4ys+jAedgNDBRBbu1i30Zo3V0CsaK2hcOt2DJs5cnpPhCK/Lws3P+3+ZaG4FBc
pAFS0pwr5UblZCa3EtGwBBcGTEGz9lLuS/mlMhwIksVkpKd50/9nRZsBMKDq/gmZ4QX9RiOX9aaN
MP9Dw4IpFzw5tnVIC+K6cWBtWJ/5PBx8q5Ye/cqo3R8XOCJbWtkljZz64P/pPmgyn4jSLX3tfJiG
7xIazdt/AlM1BhvMl3uzkwlXWUUS9/Im3j/f4Ood/O54RF4krowfRtDOTEKAECHo7Qlo/rKCrXKR
FAzTYixzrQBLHw9XqWdPPTJNztTI95OJVTVk6lUdyXtB3TA+Gsm6ByIUMtop7ZoEJwGmhBXs9DKG
vzXFhcC1/A+0yELEBJYNn2N9xLOmyfpSmnZyauCtAUI9lSX03ERkY5Zjb1HOG1p6Ch6GbBUfvn7y
OYscChr3pfkVK5dL/Z90SZv7MzKYxuR+7Gn2J6EvOmOS29bQgHWUB9LegtgHeHmirGyI8nZ/9Dmi
w7qwIA7Fepl746XojaarY3IisPxCCvayC876Yy5kg7KW6K0XtMW9LDBo7eHKvMv2GnsUX6+w/Sou
+uOIrGdTt28kSZz/S3VUMZmP9QkvWWV/1RXHmuzObyq9QQDFUwyz/beSPx5VrFz7kr8CbBejSQYt
0XDxS9bpmXZspXQMuYl0DKB3QDY8npvHLTb6sewAJs7QPfj3bmrI0dRnMt7761W/j+7xafr66/Yz
A4598MFbjKVknpiebk4oDT5uv20mUbbl7eYfWucjLvlnRsEY9BWD+BCfbVkBkLfpPAqCpumw66M5
SUGlPNcYVyI3bBrqRCyXqNmJkclyB0ayURkW05QzmyufYoOe0QIOH6vhoVXvqKmmhUrIuiK8KkSO
2bNEbdSyKHzZ31gOuAwW03qRi94HkD8yVURev3Jp4BNgN7yuvvNvHOM/9JIaqnswzkZofkwDwLqc
EVMtOEJuaBagUHHAe/gqDnJhYBQ2gTZpRX04y/o9jLG73h4js0I946TNbxrcVCV3lUOCmmA4XblL
XB/CBOa/EnhWeynqn4yiMkFugBTe+YRkiW9sAPnD08XlwtpPcHad3BZu4fPA99KVYc2QDvXy6m7E
2I/xQk7MiBrhdTtBVUWHExBamx5/DQ5lLZs6Vr27qU1KH37Ta3MdACgvB6RJZ3MAydVFMS/wSGXr
ecdP2QFnN2rwx3IRzghCysKNoldgP4lOoM47Cn7H8B+0BCx8xmGnqTXpUjZgxBluE2SBIDBUZp/5
0DVcxbAZgLD3lpJIuS/TEW7O9oV8nX0b03pg3OdtzuUb9xWeKV6d/+dVQbPivecn9eTpYNe9wT0y
slgAyKzVjfehjPcs4pmpxOq6kEuFbNZknZ/q/P2WMUqYZKlPCNrjw3HR3JSOpNvyHUeMaO8YjLNM
BfBN2EdPxmKPLw2Ldyk+lQYaq66cAZiZhdIpeSPVyd5bgD5PkRSgn/tiFafkSdd72dMAZ9m1NHL5
Fux72cUKGhXgnXGyvQRBe93F8y/oTeRCASw4x+v3oZYj4fN+K55pDo7fTtrCHTkTeugZrnmUmToh
iPgpNnCXQi93eaNubls4Bn53/Fe2A/DBx2RD4k7sXhrE1G4nGeBPQyoSmM2Lv+t4wOOkfaVwU2C4
oCmQ4xKyKdMNXTlH93sb0rLn3V3FHDz13jYE5XSBiVUfNcwKrWsa15OJqUloxpIGfQOyW58/Smyp
UGw7Y3tfc4gLRTaUb85YPD8EI5atzZhomxr3p8Eavd6Tong6QjEAviO5F65z6th993YHtVl+H4Sk
POLjxyoi67Q/CqDBFMpyoRw3tyX/53d7sDbTosKkQKMLdH2G8iqgPn2lcbPDWVxT50KCOgTJf78Y
RXroahDhBzAl+iwu/43LXoe3QY6RIyQ/RxRuiD3gPS4fpGG5TQ8jwkABZbCaPpZYH5XEdxg5581z
fKLrYObsEN8bRYv1xFsZApu3Ij5u1A/fVj+0OvGTNy0mF1LMmo+MeEzg6Ghz6iLNf/WC0MyfNpYS
vq3GItUwBcm0A/LOuNFEpvvzrQUGZ6/nA5pWXL1cB/WxtcsurqWX4EJlUaTYMwfRmj+E2kNdOnKY
5bDeUx++Ibk1/LGRZekJtoVuDLY8kq+caZ0Lubkm1uQ2kkDnEPdbAq/aVkDMj28t7mKrpPU6Frdv
NTPuGsutIVJ8tNoukr5dIISje4UlAH4xgYjqiAaPmlRsuMNXXCJ1J4TbatZzVcFg3ZwyU0j9gxxT
OG9SmgxWFotzPbxGPtRCxzHFFI8lwncOi6gb5Ad8eYH/pTT9bPz4RUqFFI6Mt3HnMAeCjU1KJRPw
V5tlKZCnDpCP8M2DG4DLdfztBiA81SN7J+cedWReDkaC4kKXUh3YUHIt7Rxjcsl83qNsCDgQgsr+
yzhOEc0CZtAVNfX6YfCHINGGt5h/tmcLJHLQd8Lyhne67LagCWDj3xKGFe7Tfy07/Rr0oY5XhwqT
puYULZGTs8p9g+34u2hE3/7buA8FLm+nXkacHwJhQ0PWbABJGGpzpGecw57JkYbJfDKpp9fsVpPK
qDQ7wgctTegeU2MJsvEZ15rTjuikd+a5Ve3q1suf2f1suZYGlkr5mWpKxVt2nZ43RQ/HyICbiHRk
D/y1a8SPkGGAuVm0sqcY4vhmopwFS5lfzKedYCm8GzdbgKQ5hyfqXKhDkPoP4T/GD1FzPnwrvzTh
R3Ps2dPslEZRH1ueUBEuA0rUkboOQcEUqDSlRQTfGJdNq11D907K1K7skxAbTbJ9o5WAZm7V3KFE
1/p+l6HAr6X2aPFXEWrLIfhWz+iVcQ5lqDVeXAKMIdiP4F0LgitN4q1+8eeoLPPcAuBEOV7T3/cv
SY0ru8N47ILMnbQz+hyNlcJyeVRVkdcfopqi7i2vZ/IAwzT0MZnqXJ6moumGAmmq6lrcJHbr9EyC
9FTbAzVpb/SDZ+bT+0L+xV10pKKzpcld1WG1GdxtJ7rgwmpg6ucJ3LCYoEm7eycgXZCLvXzv+QO5
tMZ8OQD4GiQX54zUgI1x9ZDp94+8QY1uWRI2Bshdaa2I+fWMeUbNpak1k7t3SlQU1AAdGKbjjprS
bhfPSlbnvHhLNyHnltWK4IIgeS7wiC4x5gGJ7RSw0+TBDOmlrpx8GVxmuViNSCuO5WTwcFeX+sJ+
oS/KbbN4ozpHKFPR6evxgxZjtIiLS9syW5uWnKiSXs+w7qibdI6FxhZeoz3saMaNeSlO9kocOXlN
GRkZPa8Y68u+jMwJ2Lu5jZrw6A2Heg6/kac3+x+EANPn3+3mDVsIoCzDjvhM+XnmmB3wYepuzx8/
7kkrqiUuKlobhkaiyvu8w1tkRzAkwPZlLpivsogoswgTU7+hQUVGmBhUY3HrEf8UpVnSaP4U+RD0
DLgstkcPJTMkxQByHd3V+7aMeJeYXycaU/Plz52rhjCqMb9hN394MM+RzXby+PAcEjzt2+u3zTPL
JpdFlOMXO+d5WFts9S0IA7+lPSazwsK+xVqtmzDtUC87+vWdVe88MuYweK4J0T97Ib4jU6CTdBP6
HuPiFHCM15bB9m3Ppn964nqTAfgHohdEbkVFOehX3G5ZD/3O0dLqKCozwFTUckAF2udkqoVD2Ua1
+7zUvtN1vHy/cDAA/e7bqLrBaHGrAZ4CLXk/WeXgWTycdlwN/kVevZFutpydiRAp0TAcFbVhge4C
W64VB68UqU6vV8hCBTh2CWGqnkGhL6tT4GGGLf0LSVbjd4VMC77v9JKFgYqCGR+ktkwbFIJ3Mz5E
7BmVtn4DcdGtCKwnAFZalRcIIjDnvCDES4MOs2EXuFSfyZozuaYUFbGfUd11pAQZjM07eio9UUwB
n2puc5PWAPC258dwOCzXRX26nYCOa3pKIFpRUfhZK/ZxGr3Mq8QvzKdFaQvvOaTiV6zi+Fr1yrzD
htFnPxOLO/hcIpCSOJlGfhzXuWMIWWrWP+LN9BoXGhjb0vlDaCRDHw8iP4KOc9fHE2eeYBVIGExR
DuT3a1wtEPiJOg+xwDT/l8/P9ULaxqu68ydoZZt49Y2/HKuRkR7m2jVX2J6ht6SxheL1H0497su1
ZEYiV3t1RtIKvzNB0qdMHEp4u7L2M62Y00s8tf7e1iL7ukBZiaCKYO6p02j+hr3hpeH77bi9TBq9
JLOjLOtGzvsdCY+qKD2jFPfy3JhLVRIHkaK4FNi0kHY+ntxlRqPxahQ8iJISFGF5VsqoLiNrHVCq
SldY7pGB4lo8Y9mjdyTPkrxBKQu0GY4S669sJcXZJ6PKv3BhW3gogDLrCus2PL65AcySHZuB7Scr
RHWCtT8QMzahtpINdnTCtYZrrVl2ev2FhnsJQZqGYTpg1woEE8964BFjmDg8s5TL3OdUj13RKtJj
hy6oe2HP6k/+O4S/FIa2qpDog+qIALDndAsZkHDiMb6GirlIpuz9A8TD4VkFVD/1C95Ekb5ftijK
azP3rYaI65I7KEDK7aZNNTe8Z7qeeCtp1Ar/HtKq9X0oDTZGsdGT42dM6YzciUXpy+HYU3aCN5vn
9vkIPxAPZpqRZdU+SZ0XYH5hYDWY/gA64vokzvIrzwXGvCgMkwc/3jx7+Z5tGjSiRK3gvcHBvDOx
h274NqU1dBrdn66KJfodI0b9XhR5zGKxYZLZqTZXzjZLACJT7kj2Elj9XWx9BxyAZp6NKzGobMG7
jqmIcvh2K/xxnYzgZkg5cc0GNaPHC4Z1+mHozpf0SrIs2yNDcTD4dEyJwDHe3i0ezphkXz3SAtJm
eoeDQRKbtDQ8GFJElkHjWvUNhCrydHip9IjrmycZimPMsbVr7JKF01pXyf71w5o2c3V//qDDHzmP
wYm1maZXBRwGFZZ6qo8tRxsnW6n5D/RTXPkSwqiwFYqtWRCw+EkRCPEAEjMCs86I5XvIaN+7kEEN
ungrgeutxyceSi0N3CdOvkXhACB435OnsYcKe0kUHgB+jFkoCIU9RdRqmsnHv/24tnDjw3rmcDEN
+g4OiiW5lAXJ1nPhRvVrVEzh0pPVC2KPn2hPqRldvq9846jNz5TTo/KylTIUcl7WqFftxsWzgraz
iatIwyXwOvrLlAbg46MggewHGgdA62QG+ezdYIqxgqhpn850iDeF63/hixf3cGyqMrl2ycUfnY0r
+JpmyF3W4GCcy9rAXe6JIrOmNR2+km7jhbgYg/VULLlKDkT+XG1NBMegxd1o81UoQQ0It2YRqBIg
NRVQal0zHxCjWTROwXr+pLvE3vc48Ikb9BZGobipt+fj6QdyzWHgynWtElzH+gFGMeCXjPC7Vndh
SxQMWa1yT+JZT+d0KYvI0B+yLOAUf5GiSiv0JHep6KKFNanmV18HjpRgnrggEMv8UnmJgpRZflpG
PWz24jJULnK3y0eyn4rVhElYKf/CgzAI6wBYJjqrcC4+mBliUZd9ig4copFxTRAiAPrOVEetZzQd
SwBG4Lffk3QkcVgFtA9XX/SbsGh/jp4lH3HrqZejoyzwX8MXbJgAlLJFkYJc7y++zFA7qIezMaKp
D7Bvkb1Wrb4AENBY5QE3AUc2G9mLHdFBt042oRScjxnlkg5ohWObToRDgMHzrGuwsgvv4Sgw3axh
Z7ua4g4PQh6dUdSsxEocx5qzlkFioUyEeR2GE+1+NXN6QU1zH26augNf5YNriPK9EpPt+3AfxkvS
bkOXZUMCI7gwKYvPVaki4cInw+V8wbtjBcbAF+V0RHAse+AzR0rVfx8WKCkN2eJ/x7NxLIOp4CDL
kaUdLFiXvu7eybae4BUGvbHVRWod9/i8dCby0GrEYZYTy/UZNk9/z/ot4ZFSeFnIcdtnpt+ZrLQV
9v6CfivWUUUMWvo+bHGmH2XjuNyufrHgrhBlU7XXkzrZ+yDg0zUUeBrldk0CEsFpBlfbNXqVxKJl
e3BPHWeckXHYVfF81s6zF1gVTdHAJmTU2IHNVwIBLtDJUksZuYAZJcRy5H+UTJHtLT37z3kECUr0
sk48m9kDimcSiAMHqpAV42JVJpx3nyLLHEqho5KO0qwY3vkxxDNlRemGj1JPVAEnxv+jfdO3IRqY
eC0eCtkTCx/kBw7ZO2qvOPIewLOMC5jRPtZY/Q1s3sNLW/HPOiqiio5K2M0xF8wNy5OCcUYaLfn6
G9fHhQd4QwLEirec6kOUdfAMarxO6E93iXh2WnWoNv20apGDcZDJiKiJX1garby0fgleOlKcb8Cn
+acnD/TiNg0VSqKlz2u3TTMWprFKm2dQ1lmLmsk0FQT32w5ftHJynUfK1m+MtYz+3HvorkkYXa1+
uz0NKoPbL4JwEQp5C+e7LgeHJONl50HCU2m8oPzF2obrSwNFlnUrOhI/uo1A5fvOY7l7lAiHql/3
gCNIyDBbrxxtUmtH9IcIvb6Jk/honZe8aWcne1m+gHsGzwmPQOosC/T0cXaRiW1UcY3LiSMob/fE
9IzAp8OBIYVxNN1e4E1pgnG2flu5iejEGHM/iXNs9RZGkT++aSWpUl6M45TvcHM6TBgVtO1/YfaU
O4VvXakByiRIui69QLWB1XsqOJr/HFEXocnc87OKfpV7zSWXOGVmfY2B36l4tB+CdLrzFVkWVo7w
q3evtJg9lg+nT53UBPUk2NS5E1xavpT1t4uYfHSUqQHjgIOrqRThiTjWR2LrmEVo9uxTLu3VFGYz
SJ0pTfuYI29nUK5HKfTtr6eT1ivUPUMpz+jH58y0prVgDR56vUt2ER5QNe63JEIkdB4zuWvLA4GY
Z5KDc8jWuKnxQMN6Nf8tAlLPGgexkZuT+eqtXHyOCW/Tn+ROFcJDhBqUrqGzLKAqXmfEYr2wKJtP
/D1WSXFjwjJMnLY8ONfRFtrx4kQsvF5euHeJxMQGmirp6i4EOHuXbEFDLOcJ2DwGNwUVgOMKpcAX
zrpEdh7Rsj9zGC6aOB8bgC6sdj9BiQKICpT9fR/i0Os9kfjtGaMzUC2QYjYL7+5n0CZhcrHTsnt8
sJ5rXRM2IOeGbHgw98jENDERxTrC9HGSLYslIkUVP5pjqKzb90oxFfxZaQLvG3gafTs3RrBTHJkt
nKEy08ORws2t3cc/Cx4YnPLIrAJ/TZsSKQPczb+R/7jLTlqehmcGDwsA3mEG2m2u/5tZr9KqU8/6
V/dcoLAdLZlpmQSxYXcX7wGE1HRycqXG4Y3LKaBzRfy0RPRQmGKAD585XeO8/b86j5uEwMCM6M+3
Gef0w1LCS7w7RF4zQVSqrJbX7UOjNzfnUhFTVWf/PBYdUl5fQ2PUIgOt/rZaXOc38otamwdxsRlL
vmH0+O7VvEQ+P8HgGO9CnvGgqIcocbv8cqZAxPD2F/Mk2/2UWYhW6u31O0rZWLs90XgIL3WhwgSR
S5K0dRhu2pAivSeXKbRvjSG5VZ3tSu3pqtTtcuT/Ha5YryXWlMwD5jZy5Upn2qsv2Ge6/+4zfuaa
eCbb9UrCs7vu88p/3J62vqsuUESbpGXCReu1fpFdQN8S35wplfqSMh+wbr6mHc4/QIxN5Euyh02f
ppvt85wNBhDw/f8XE1SQmVXQfXK/2eTSJiXwQ6QiTG/S7KvYUWx02xkrwvYeSVs5LL5yyAggFzvX
hX0Droby/rpgYc3O9Dgw3ZhWDcVKEBFpOPmOBnzDAgBJ8GtH38IynWkfLDK0X4clTFCpdk8OLa4E
xlEOdPFyKnAN8JUkJICP0imdKZNguL+4fXdlp0+SeHjdhYzeljd1bbexqP+syhFuqaTfkprviA9W
sVSmOHjmqEkJ9cYiysIigLzxUVeSDxm0jHeHyxTwIUqFr4rrB9vC9qD4lVbtT35DO4jZlxtRMVQ4
JoU+ViwtrJit2zkGpfLFHVcYxGSJggQyWuLW/33SUHxpb+fs4FKYzp4ko4okftkU8WBD++WPLsma
GDr+Vqqr09DXGECYvI4yvqXN/59Chf5LABmJwPGLBAGsaB1updO7fVl+xNKOvQ8zxl0gOkiu1up2
wvziXy/Bj88HhXN5x2dMw6mGE0feSZyUBE6Gj+RqsYwJ4CHE/5dnwE1Aqz4VMkjk76yx0oq4Cnb+
Msfam55pJTB0vka4Myz6gUoX4jl6nXZx1Qm19ZDIjTFyEdtG2Qhisv1mv5M4IH3vni8LH1LbS8xd
qWedBySKvUXwXa/xNswsUjbZP6P+6TMnjjX4QJrw2nf8ptg8jPK0UjZv1442w8xTPJLmILMZlm4S
gFZn06yVypYrzHA307nKK5BMkI+N9cqXCr3ygvZIJWqHsY+0OHxW36QQBisf7zLS4vNOE9W1FR0Y
Cu8Q9s0fHeMxyrOD4qWJliiahkEODuuaq1EGQXAzQK4QyULcJIFMFRtaWbiyMrWGA9c5Ja795lu7
UClp9F1AogXZavNOFMFF2VC677eEffZjeGpM+0ZMwlj1ON3mDmhdeLjpFyhb3g2YrVf3uGoWCXoD
02rIx4sNsIIaMYP6pAEnDT2AUEMOeV4Wj7Xs1/JEQEkFfHkUI3vUD5yfNtKivO71XVsRHGW2kcGn
t5P+L4UFa/w5PIOXUMb51AkjMdsJ/3D2YA0sPcmAstq7s9lM8Lj+ZH5uVMaRkbUSl1hkM4L74E/d
n0i8SngRo2LkA/gnVsil5OHiXg8pQSEKWqtopeFxhLEJN65CJOkGJFQlREemiiaBVD/6+17UkTcs
dXmmdJ/aXHi71oSGR04+qncsGN1CmC9B//oSEApeQ0nbBsQVMe581ew/1vgxbvqfE6CIT5GIYoGR
Xe9Qw9fBpPXybJxObx2blZ4kgRDfPLXMZz5GXp41tt8nVwH+t8Gft8a+jjp6TVEG+iHCO6Qd4dpI
PxkI8mbEcvB+K0gjDl5iCsPwv9KQ//4H8P4qn/TmdPncOdsFspmA+Ic2fDKYASIVcYh391xN4H+E
J6NjxDHM/yB0/fYk4AMdep1sZBoh2feXtGiTieWOcZ94MaOKv4VchTtPUYteyKBpFnP3Hnqtxlkz
UYBQZwcXtRLqKeAcCH/5Tgcvid+rqZI3rPNS56lkZKGxb1vyi8TtuTLQQw/l6kGKnhqhhzRo5vcj
qdbAufBsJBit0wZpJKFiyfBPzakPE9eHHYwb+YvodvhRDydQ9zYIXqoFwKV/oYfDVWGb5KSF3QXG
asX1E3wWc1nvpT3gAZ346RiREG2jQm5uk0mixNP8fT6ARqVEtYKt1GEWK8ghOOu0uNcqfLoWWnQa
P4FeLWCDASYncMNt6uQqyf51boCNjPTaJ7sBy7GgxVluh6EjWzjC2B0kGUeAw8uALkV7zMvaR1xb
qB9hD/yKApJtC531gMEWOJMzzhbcphSqqfhurMdo9IPwFHshgOgO+aPRnQ/TYe4ZdwMxRktqXcBi
wI5upx6J6alU1qEHFW/CLZTr2GUl7Vr+J/o9e0zy461T0yS/Cbw0lPSXUjdmCQZWcmibTg4kcZ3/
hRibXKhe6QgCSsTPXO4zFKnCtD0Zq/csPdJ9e8QzHA3rm5JgecHexbOGjyaKFoWZ7s7yCwOenaAR
F39kza5j8lNWTLlTHBX3z/48xYTeH6I5yr5YqywfQoZg3++ceNv3Goken7BUy21FsDDXgEklec7S
lGUdIO02BpNtQYH0lNx5l4uifAOJEqdhCpe3TALAJYOuZ7lsbpZjkOlAayxEEo30w96AGASJPZYx
fhDimzpV0OKE6JpgBRiPH/BuCHi4OvAZvFpi4a1oeqpv7Y9c18TwewvQR53d/zks1x1RJS+Fuw3y
JjG+bSNfPvPwZBkLd2CrmIqtOPnwCxJmHCHQ6ZrzXKqmv8v0VeMeAZSbpIGBcXBLiYFadkOHa7lA
5M1u9uenBXckimfZaDp0SMPSry/ret/PnEo+y33j5F9g+TnF8XjgaTdZ0HKPg/hln35R0cF+9Ps9
eXdzhmXgYhNUcKJstILEI/zRWrPgb+inwwN4whfTFrBms6ivGrjpkloEJWwr5PqfJKjJiswPEx5z
w83IcHl8oF3l+8svBLKcx2d00Qwe6nzkb/sG+yebuUn3ZbOVD/oImzDEOsRkzjAtA/pXGJN47Gaz
qU2XuqEpI8etpwQ94E4Kawj0MbU2YpbQP2JaUhByK5OVwzTA3bLA7ouTG7dfGVizqu7LmRzXP5nE
HM3zUM16C0nwbv633DPRuKuj6BkEJdj8MtpAQec2ajcQDUkCmPLH0lb+KeZXVsPN+VYSNtyA8/Ey
IFNc+qh1wfJZlambqxY2ndOnNuEVFwQx+GdgwpeXK+fiSg5ssq7zzBeOBEyTM9JOeJckjVH5XRj9
nMPmxYrVic5XJM/I1R7rjNgbRSc9t1WOtm5msKe2W20sr6g+kPL+enRnGeB6t2AuRIQIUUEsmy7D
QUBvKTIYzaR9IL/Gc9LsVfthWiapGyVgVomYaJiBTrqq1ColVKfFcXSj/96XEA/dS/+aKR1DuSH+
XHHOsKt75f/UwqMbhoFerDMQb6eww9B9kr9HYXOJUQNmeNd0aZcAuUFXaWWw1exc5E+KlnbGtQ5q
fQWrWYtzwTaQjK1bizAXNzzb/SdtANQWhYGshpbBf2CAdlnw8+9OhmsDLtxG5Ji0EfMCssSG6Sa5
hB6wWiBX1ewOuo63uHgq5f/PWqZguh9ecxjZGFuR9JpMeozd6arvfX+yjFXutJ9RNvssdMEJLQK/
NzIHQ+8xcKRmKPqHhOdGrDf/1VFMwaBaP3slZ79IgMT3ezVM0Wcl2ew4ZdMK3+lCByAXby2J6l9a
dZoREA0zVhPZTBBzAH+/OuJB5c6V/asPxh5md+c50tUc2+qEzjz1oZyWGaFeyEOvm4DlH87t8lMm
srEgUtfi5v8h4XR4hbZyLeHz7bga2SVtFYi9nrPtneGTRleosrIUdQtq9GagKUSGBJyJ+BfMMDw7
0vTULjQJvc+oj+5jxNd5F5vNy/A70/tyljOHc7Lcg1rV/XACcxhZRvVY9vrfiv59xRob4sTvyubW
GprdEG3tMrQ7D9yOUa1Z0zzaGCRWLZjIJKghpg00r/L4HDcuLwQHeDm52JKQUgcaljflUQ7gEUOO
NKzNJbBquwi4OJyWpOFc8OznWT8WJdjimumplhPmcqiD3RKmgs8P22u4rprxEf39jaAMXeuxhRxB
th1zD46Sx6pVTnkEAwn6ql5yNFwC+VZgCnLi62Y5ZCPc5UjVoVm9WoFWfOwr11vQhNx4te8U/4Cm
yOawylTiyRTd1DCcOYP0f299Hf+bOBleLBfJ3V4ybhAkBMbhaqOMkBFfk2KuBmfwmd5VjsPHVWWs
1KU7JFEjEA8ixW7SmCN2PBNcp3WHRZb63ynPLwA4hCMwl0E8gm0p1CQqpRgKlNGsX3NP+hYmTE28
reT//ETPiXWRpes5Sao+34TieTz64x0pnZCTqxYWYllJIdREN2Ns4F2f9Pk7YFzjdR2zPJyvltR0
H5TM4RwSwHhpXIV+1yStStkdDnUa78gBz2RE7PUVSybnXEgZc5U9fXz6wEpjl4xU4Ogsgm1ZEMZy
TxSGvllsJlC+GSPYuLeK7A3uPdcYBBvhhZ6Y8KyTjxo8+QBmsbgjBjlegyBywJ6FB8rG0KgxDmjg
cL3wOv0wz8UffPGJM0yEtEWnoDbxzOxpOXt1M009BoJSl3soFIgEIz5qvAPsi5yG3mt7vcY/lQVB
sHmuV/qgS125DXr8RxWM773PNVSi3Cmu+Vxa5Femy5Rm8ez+bPyt1j7zkzn1AHbOSxELt97MYRVg
3ouLkYuyuU0floyhWlvT1aMgkGS6EC46mtoEmNq3C3UhRRJgqE2ZVBdWBDb3Ix3dUiVvOKCM+Dhh
n64qkODBOa5kQEhBlIqa/dExn6vT18msIe56Mb/2c9HetHtGVAeduRpfxLr3kRNRyjd5Ke9SxLLW
TbbJ5OfzVjVKLFzum5LEeQXXGNwRTGZ96n20N0n5kMCx97axCEkR5dJcrZ9x1nD7xpaPmxxstti9
0BwsjezwVS7CdRWiU7xBaie/nSUPv7sw8nWVlGSKbxnbLmQ7jN/n1sH+VL9M897aMJCiElESW+LN
HDReFpFsp6jWOSwHoY1mVn1od2WZyy7E/xtynvFoo3zye5EbT4Ba18yjCeGQm5sBw2o2rHUw4nM9
iIjG1wTvHEkxKS7Ay6UT+x4XZCh3LVIJAaOVTgRzctcqouciNN4J3TsCucrSPNBTfMd4pPkXexIy
cItI9x+f+O14oukqUR/DVNx6o6cnZ+b81uMKZmsiQPL1rVWHLgCsaC999V4PQxr2Qf9UZcfv4QSk
UFPi9cXIfeYJts+AK56iZ71/aeYf8kcR4BQXjtVZTcRH3bC53z5KGHmc2m3uNd6bk05Pq63CY+cK
04y7sKHmjYkeG3D8Qq+/LvivSeqqvrx2OZApFFzFZS3j2buLEftSc7Pd4VOkmyZ4vRXctiLB3gPf
wjvK27zyyui2sdp+QnOQJBqIK/xJFab6dT31yAxD+uvWA50i0YuMV6+q0Bwvx6cKhggALLCVV4FJ
60DmuMg/zois0aNema09wAR/g6cvgl6ZBtUNkxlJZtgA1mXVuZcv+7MXoHosUAe2NLk4isM5gNGz
mY5/Q0R2OU34z+U5BcGVpax8Nq+QYWDMy/LpXgCGG6Y8hbERneE3EF+VQmzzbIGrIj6eWIIdjApa
OVrrwJZ997/aP32VZ8TgvhudiXhVxLVw3gafftVQ9FAr5j0bbNovBRkngx6ErkAC8hp9aTfY+lKx
nkl+K5cGZgTvcwrWjb8JYdkdGikgSGczg7Bva9fYT2mBcm+ZIdtQJMrvs28inK8BKWUjvOSAYb1Q
nCQl/9PHutm2hHlCyrHvUVR80sMizDbaWAbRuDUG0ls2QecDmBgyG4+QpL5DVwbWMajtGEdPBAcZ
dZdJ3sQuTNFvuqwVAFRtwxESvHeMUg9lfZfDpaLTwk/QwhjmH7zxFwlppw9vis3WA7IqTGNNe0e8
ReCAEYkD1LWfXa4EE8pqFVAjMgN9jjep9vddRnhQmlCDe1fT5Dl7uVjUb9MjT9XEnsmLAzXlYbtC
sulzL5kIQ11imJ1imQj0IpSGjTXvi+Ymie/DY/am9n9uZuDf4I2M4e0zbX8/7N9KpD9oA8tt3Mec
tKVbYiMJRm61xCOU3PNZjd7zPzHQr7z5+GjHnbxPUbpY4byIxMg5/ro+Bt1VaZoD1QoJ1WLhjJQv
yxypjZy/mikmNU79h3fvCUAZ8khE52YNwGIxxkyM9VJ9CHsIF3pRGDhD2rk0682vzaWVr7jDemYt
mi3d7s8l8iGCKwc/kM4y7Kf8LAGxwNgZX7RqoBVpuufEv7JNXUYBMOYuwSGGrET905G8CcNXB1Xj
SvrN6B9JeEsguizqYEc5zqcrq8aL3Ni6zGyFJgQFaDaqv9gEeWivE7yw+asTnZvZZjNeFDKmrGs7
fOY3JF+QJ+EiYr7fxdbObbLuKY+EOEnzgl21MjgzWV536xy9LQSG/xe+qwCAjiqxEbw/+oBGm1Xm
Epa44Nvrfe/SMeHKoTcExVHVB0JHB/MU2WEu0914xqMDyONRRQslgju+ClDmNkNKii9xvdI+5gZg
r1gSGXOjVkv83mwtP0KnuUHZ4O8bayMFPfZr+vpJjSRbLviuWaniMQC/O5bV6ua9nsadG29UJFvR
RU4CIV80L/GO2zrIlzgEZVa9xWNZ138ITSDCc1BzvjzqChdXwA6s7Aa0H3zPQdZt8CsDThb0/5Yj
fL38Xbdu/Pe3p3N4U4qNQQTprR+Pb3GnjdBP2beZsE0P48o0ES/2fjFenW4r46bSRA0XXaAmAbM1
d4gkExC693OYJwGovk2zNmmSbBAhhJO4eGdAX7EGvT877MQUn0oI1w3fMrJI1S7rZUJ+Pkx+CF2q
6XsJKSEKWuRAzGXNcNQeMifM1T/81aqGCmlNAMFeLMVN8Svw1wXsVNXgeP+tAt71wnjP0+3UEOc8
9UEbUZC2bepijIfqlbXbCIfX+KIRLHozdl17uNGbcv2jh+kxl92zsUttFLtZoHHsD0SOnDuCiYVP
i+R1fwU+n2ZNPu0NS3mBUataoyGKEUtviU/VQnlivwYfg5vP249GdWD5JFGLbML1w6ayTsDsKgOv
zlDXdNY+PPAbVvQbpnVZmaAaiSWDMpNOxoaWvyHDeW7d/awSS7ZgmbqeLjb//WhqvyRr/t1QSRPB
3+M7D8F2pt2TKacfs2fuKaRNZklsFB2VTZBoqcAIeGOemUgeKOfMlrbtMc88eAwkpMjWFrrcfkfk
E1ip5qVQS4XC/Gvm8lavzP7UGhACYW+c7ar57033iO5qswKy77ZtGWvcgYdpRGhB+BZPvPgdpWqF
dSPlhs7mAHr1Lium0DfLzq52jGd/3euRexXauRGZjFtGh/8Pnsj0ZmQs7z4Mmot7LRutiVoAZsOi
dJjwkX/vfQb963x+/tHMzcEE6ABqaspVQlRg3v3XWiE1GayOpSJIJMU6SMk98yQcymNHCR55hzsT
lgTTe1hzJbxiBjKg3fxhoVzRiuRaQiPdGGGZr1M8OF84TfpRL5FcmqBdStz6dJWcrKVoQGpjuIGi
SB6w1OBi6zNCYJGDQ3Cex9m8aDO7df1e1WLlFP9j2LHTrxrvdkpw03oxvbpNlGy78crC4QriFdSn
jK7vzWT12oCWQtrA03Jx/mWgkNMz2N/kU+9CbYSJOQLpkR3uSk4cI0xU86bmZER7iwogad1rE5AW
+qE78ZOcUmTOCBZ5UDtTpFS0dKi4w6Map9cJdkovqk/3S98D92bi4FMFNoF+ryfm1QMp0yXuydsf
LKmCGauvXXmfzFYgBO7gErt8sOYddNoAyxfPMVw+96tSGFdUl1V/zjHMwhGGZlvWpyLL/eNRtHWu
nmwoi+C84O19nWW6xDuwOfusydMgeM4ZBUeodz9chYpmgpE7wA4tLW8bcob6ib7nuttuRA0I47qu
mUR0I2DwoZi8BB1J6eg5R+uI3vWKDkjUqv/1TredBj3iR8PTw64DtDp8jucE1ncQpxq8q8JYI9sQ
qjiGCXa/0ff0WFuxjo7I7y9RTxD9N37OHANMxvynib5DBwZSAeY2fIpEDucfaWL8SsFWuSMGkg2I
ah7zcYVjb7T99LIrRuLLy+e3UnsoOsMZMUf+IuIyiVd4b9EfTAP9j/JoSKb0zz3zUy95To5xcHET
4xtLzLM8F8h6Q0FSONPwWYdpC1Yj9bMcrdTJuLRUUG8MhfCSEdiHL87+LxZuTOf8edulYNXyRKIA
9iSf/52dbxSCK2GK+lwT+n3KE28F4k1jiCDcWV/r40vYeYK7zp6wQF8175I7WbWCY1At/5P14mg+
oXMFYLCyhJmhFutMLW1ZD+qZSlzvAmyAdiCFAgPilVIIWgtKhmJB3noHT27Xe6EsuZEeA/qd0ubb
iwaBqwkVaDiioSqJ7BhhmA62iD3onn239ga2Iqs2ztiZ3dUg9YeiRvoDnvM9yAme9sRFJtoprLZz
annMadg+3n5pNAhdpgMnVKKFTCEF7OUheMYwrI6QECeToHTWY8IXCutCMvMWb803EQ5kfq4OOToo
BAzu5na447Z+V8+YNZqc2q2j+9edsqutvzqgfwbTAZVT+mqtL89QWrQ4kLjNoWI+lYYpKP23Urco
LlXrrPWqNDUtEtapPRWH+hZKklulyEFl8m0MDWvEy+2vQujELVZAOoOFiEuHBhvK7E46m/enPwey
YqjkXJqZwrHuYKYovg4BkmIF4/I8GDyGMGY504SKVwJfdAznAhTLpEBEzp1jX8UCpbUV1aeLloli
bi2hBR2aox0HfU2OVclXdyImfaW6YavMqdEZbI9pRtAs7vS7V4Zv22N3HKD0FWJO636QssizAUEO
IBjRuMzghSfnXWR2F9hrvWE3Et8AC9iKsK8rp6jphyV+UnFyhzjZoq0Q+gbrjbPVV5skLEQR9MH8
3yccUE3M+vBlYS+IZlyRaV+rHGKkYstKPHlrvugNjtjDoi4ujGL5ZNQCwyj/w1l4fdpD0pkcqr6P
J8H7b77d7f9vPhvHb4sRc+Xj+iXegsWcKUyna78r9h5VsZ4Ce+n7O1reugHugDcee0rWD897Xih0
BUGEKrqjSA4vmaVkCX7OD2sBd6/HH8J+AHKCddq+e1O1aE/CRPTYBrq7M1ZXQ6XVoe5mk/oi+krn
CH3tkLXZ+1tuPgjFN0v1kkbzelVgcz2o7w65NQYMivayliijsOrnSE9tW5y+FZPjwhtM8DnK7kwW
9hwomA+pECCYhUO/+BiaiUl/71Rd8cUH5Dsq5dfc/Cyx2Xk/IJV4yyNtbi3oe0bFkFGR6Exoq9TG
A07om55nBT40j+XqJ1FHq4UnkPV3CSxfLWc3kTJGjJYTwIOagwjsQiZjHQOprEcH7pqNCeqMbDP+
7EJBeYLSRaSGXWI5tWAr5h8oim3D4MDWuPr0239GKhrkSIDu5G5CrGytMIHwauU0KSC1qJDcxzYG
Fs516X4wg2scwHMijzvf+m8+LImnmNWoVHgLtJc7R81kz7zJABPXh+nYLE3zZbWu5jeMmUVCJX1k
tTB5U7l2GLeVb7wLsnpecLafgZ+vdKt8PjC056iuMz0y57FxDZjcK//Kg48maIWKab4Ho759j99z
Niuwcp9wuGUhNxy20hBAMtJIEm3ASRJBY+CobVjx2EATJxuyeRou7Xa/DEJ/XgBiaxIESfDuuPQA
4BchbHNdOofjBLfbsjFj13Uv5WKJuESnxdQMR9YWZj0fhKtqVmHSJpGp/SBSuhT6T0VoHolTnq0u
Ay30D4Iyvvy+KEePuQCQxR6W/wTpcK8+JcGb24BPxr2FwnjdpctJUtCP4YvvNSqBTHO05QcuAPSB
SaUK1Sa8BYIZs2byx6Y1gWNtLlqX5BHApVgqyf8W0KbSXciZaLZP249yKsbxUuSdbEGfZPClf4CN
qOBxogoxlAjNuW0oSGt2E2/UdRIjYjZo7uYiPR1IrX/j7VypF9P2MObXpATUD2/FqQfwg10EVNDd
vnAVWz0pBHAqN5XQLCRgrAgqjMk2+BBlDNAkMHNYWWC0dd14tfg6v4bZThjoUJZRqOeXjujqUxWG
GP/JPRAJAk34hRYPXLH4LZk3XwiDEPsrTjYNAWzUKEekIPvlyzyimosZIoY5icKticUgdcDErCjg
t/bTtb+bvGtso4lWhnla0RfP2lxQG+26EAi1zN4EKay7BYsV14ED88DHDx1rXD1uj5QKyLAg4wmo
J4Hyiue0rqKQI9jTsBbbI4NZ7TxVwchlT6PXiitnMjw1MJlsCNpIjM4LI0xRY+Jetdv0cvTbiY3t
eOtDUg3180UsnxEsayjzJTxcpZwa9zgT6casfpkvfiVoqtDL/sOozNbep8VfkTZGoWRz8XHK6cz2
ptNzDGTJpb5ZFq7hjtAIuHp8IW84b6uvovhNQEFT6AjvMNM5kcnf90PBx8EBeQ1vqiNnFs9x/INH
hKwlYhTs5oMzKz7fyeX4dLk2yKeGUIc2ixC8q+62lmrXD0ee4+w9pExFMYvP/J8Z35altWfTa5GS
UmwXcg5o1aJIfJAryadXzM2FLcuTsL2PqyGkWODRXOE4sjHHDAEVViBYurxYza5Ws/SYvKTBKfP8
l9CC+HHF3/fSvOoDwI8F9RrcAxdcdsqflnm4o1+NtQG4R5A/jvoT9yMotZzEh9/fVQEeJr2ByN7Q
Wc9Qui3mYH0Rgv3ia0NgK9DVqhjFV0wqHZiFfgt3mV2Bzdv76je1vZVvrIpPEhEfQdSS8ig1UeMj
4RzWbW+d6vweX6TrYjQJSUuuBEJQ/XgbA0HzYZOelVcIAKE0vTwY0WoTOD1BU46JvrIY1r5Uxr29
aseanfWPwJeTLv0plyHD152V77G9HG1nPfFvgGouhSotaz9Rji29iGUWMIEPj9cABdDZ4Xc7UvY9
lOEbUKj9RK3vc9rffthI5eNaSZne5ROtuq4fR/2NxA6ZagQ4rzz7NM+j0Q3nfhKPVZgoQZxUwcYn
qI2Y0BZJrvS4nLrvfc8IrXL6AM3xNvuDxXXQj3uDWIraD5GD0IelguZwgLgNYunG5SuS5fQ/5xiQ
H4tIRnTO0WJu79oXwQpchbwk97FMu6TiJMaRrt+uz90uN9fc8v5IZwSkUSsIV135mP5eCvVVc2nt
f5tN9xhOySwz+FdRcin3xUK2Cnc8e1wskSltA8lKhgU+yI1ihHD9YyFSgHjQIYGUY5IpNQ1ktKUD
liY+pKLS2CWDgDopeH7q+CvdYMu++lH2z1vvgqZRs+kmoQx8iMT1dtw06TxRIzsPb7ngGzEliO7R
WN9Sv5SqigVF6RqqNID+cFeg+8wdhfH/5QyiMr0HkwLOj/LYYphYtTDl+rwrCkyG0NXIeBvpyqgc
ArdeDhBI0yrKuo13vUP4B7kywCxoNkGTUMl+36aXeDLmk4tPOfadptpHKUEmaZ7x0fLw/StnE0Ft
SjdqTW1Xccm9fkuo4jT0kHyAunmybtd+CDdg/h+wgsnI/JpeehOWDCQ2QbU/vKap/eDgbiGIC6AD
kfS6H4guD0AKip6iM2PvwtGI3q7KjBiGOREFDTqFdD49WfAY4UnXKAkGf1APumr4iMUE9wfDei1v
It0N8famNd0jXMJFwcom9MOOz01MafWV3bAGorjF4b/hAm9UO95FWTKXyoKABmhzIwPw73aVEB8w
KP73Enc7IHAU+j/2Z3GGJa0ay0GJ1EBej8CYbGbq9Qwxkh/CHwdlfJCrQg7Gn0lLiHDjl54SHKHJ
b3zqRF5ydrEu7UWa7GEHnLacJFmBlVrNtvsRCtk7YWYHhOj8Tps7yDYvK7uVOhc9xDuME+AKF82s
UYEVbc2Mw9Xy9iK2oMUwYYPYEHRlXNQam+9BmD9T7NKjAfgHYNzBqkeTu/2ekskRa5rzRWnHqmhq
X3xhjS/VeXXyFq7XnQKypsFUc+TDkFrHPIeu4TUIk9fPs0HbVmp9F/mqkjeo7VqlXG/emFab6gjw
WwyiKPVlukxXY2SsX8hikxhzeozyw3buOzf4IaN6VDJwBuSfSqyLsVAk9j8Cb2tGhLMyaIFyUWGu
z0UgHrjm0TBdqt1GJuAx92rFWkPE5Ng+b7t3aMS9DCjwXY27eQ8dMVq2AnS2ISUA5d4/yPA/mMzb
ludM6N3LFG/sYkAcSEQ7BoC77Qhi+l1ZoOFi5FpOHKjWkzHRKAjhnw9Z8cbt3u4g/jiYHU5++bLj
XbMSACPcymB/cbzfXGrWWDN336jnIw6jtW5aJ4AyVcg0snHWZrtYdJNe58US3A4VHqbul31gyifB
/PqBxwGm6aJ9/te6mYLdCBtqAptrf723mD8JLzKfS9h5yGKAS6DQ42mNX+32+NT5j0jfgHLe9pxa
O0mcUcTvj9zm2ghqPBxclCFdZW2r+GXLjOu8ITbAktGCd+I0uWXe4WP+TWaFN5FqQrXHErjibp0h
rpodwM3fkAMMjnWy+LVPOByjpz1bJS8Yo0oURco565riZ6JneX19HUHs6yS3Z3coVNDOX3QsQ6NQ
eiGZs8V7ojFFXTcANWnpIM11kdVXV7H0iU706QqIP2qx76pjt8D9MfQzycfQ/L6jB6aqcxfcL4zC
aHFGIfCoIfF4JmlGm2uO6P9O8xCSZ63eTxrrIS3s7xkQt3Ew86bvxdEw+IVkmo3Ig+TD6BfTfCnx
OiI8tFeFBSU+CLwFCcseXtH+in8dxvC6VxG32FsHXDIGHCvkCSGymCGFmV+BKF65S7J/R2w1Tnfp
ECay8R1SVgpZxWVpvjhXcFVS4IOonktJzs26Wa9nPNBpt46DmADsyH0yYDF6UXjoY2MBmkEu/e3W
tdyFHf554KEPLUxpwZKtTRrvAnzPc4o+U9aiEjRvA06kbFiQxiOlbV5AVZaKfcIjPDJpt9mizFbo
FxoD3s7hl8hpgyLiE8RefdOuW9AJC8luulZB5vUn8BhVU8PfXLgfwGJeEVHAJTRKiCn2ww1OWnWF
4KqV1PpYV5Me5tlaDwgeigv9XbvNmYTRy2HxBsMnS1UiBkCyInDEmZBV5y3dwZKlXhGro5w0whap
UM2gnAU/9IVp1hIC9HYM1pq1zdfM/rXrAXZYxzjnPV1F1Ur+J4ERqaZkXBcxJMppURwAdpYY+H+4
ABXrwaeM/wIS/cmMIdNevvsx0G6IZmOG7s8f3oYzTDflv6I6OMKfIO2WnVBhe0GVtXrbleZqtWZi
sJC9M7v01z5IwgatEtbWfRnHxagoiIZ5ONcno7mB84bsX5Ev1Xq8ToQkMn47rp3kD0dGLfybFkqE
ldOodRX5REc9/x5jAd+BUklByzUg6iWqpdQDpkj4sJl1T6JEh20lP58s7yrQNKrmjtEdYWUVC4uc
PvmIimwsBMKu/E2geYIpT070qegpyZu9x3+bcOdYHJOFKPqJkCUqepPNwshu/8ewQ1F5/HsvFQOP
wtQyWFI22WjcnGmWj/BR2HYyp68zjWNT9PNWVzrrikI3UDJF7ndlVpzCD0hx01hY09Lbd4JjKaFR
Ckc38W5ud1E7ILIVPgcea9x32IYIqFPmQgiS1gDZD/Ek0qZX4U7c4SNdZm/JQDqiBbqGkOgz/bRE
mENeVyyZHOB08g6UnOVdD7r7ADJXolY9b1zO8p8rP3u55iMk29aQCEI82zrbu3ax2AzjA7QvnXxT
e0VUJN5+DRTGIcBc1XBC7ctKH92uhi2JzxFeqFov6YIZoXXUfc9y1m/WMNILunE475w68PbY1EmH
xOe64Sy7/goAJKWnO036ZdrRNe4S4igBTjlW67N7uNXWVJH6HMpk5hBJjk9csEw5hKFmYZqsSyiv
6HxnJRpMzkAn5gzjtNBPEP9j264FxF16edCP1vZmJQ4X/zEd+6SZh17y6jeBgovroXEFBn1AvmvI
YJgf2MMw4YrT1YxVtduazvlGH0Avj/O3QbH2yMno+eiuSvpJ+2p8cC2KDuPLhdtaFxrFN9mZFRdj
Gc82kHw/Xx115x7MxZyYDdgXmXT5rRLuMnp64PmPW4Fr496Yt82gskhoKBQg7EH3fATTCPrxIJ0d
2hRsdPzlo02yDx2svBBjNGWntuRVf0Z8e1EU+ENW1vTvQm9juQmYY0PXTPC55LFLfUDJ6l9HBxg2
oOQwzrWu/wTFf3chhLy3QYvEU2IeFitbuWsKtplWxs7DNbZFL/STuhIDLLTFULkbLx/+9xfBAFkU
ayj89TltP8lnzz6mJNSIyKaEDvZ+E/HF/lj7NEZZk/mmYFh1xFOGFEMhaQLq6nEnZxQpklsDja1/
VWkLSZ0OXjDBcx8d7GIi6nmfpzpXyZhX0xhE4CN5xrn7EH3liLUrh/gs2TB7U8HGnsg7EYuU58Yu
jmC5bRieCk0ueJpk1LmTBEc9mNWhxIFyRFtLGDgMRp6k0HN89r/j3N3ElDSLH7pL5KTb548yC2cr
GZNE34HyejEnDC1CH5rzuUPLL2jLlcer67E4wHcHsWdqNf/SGt1oERZtPKnY6lGK3voj6PGgVK8m
xJMbZoLGc6SJvKQEPi2hSif1G1FS6/7mtTnKmBmTn4wvxlWg1NfNxh2xNcfLFMVJHodEsN7f3Lp7
HjyBSgM9wN1b00KqylOj78pJW4MfrNxhSOEQ/439sPae+wse+s8/3hPJGMsvYcftPU8QxylW43WY
itWBdZIDE0uJQkZcp5E+sFAqYHVJCkgWyNOTS1BBfU3Kux8MtLG7oORmdgJajOIlQozZh49/y39+
hAsh1Ih+akRd3sK7XOuAOZTVS1qSGE9yKhYDJLKc+t4LaZGC2ko/u3rB/hyQdN5eDfEFvh23l7I3
JhFRT5Snh5eOAPtZysD0213YxkTbD/19w5/TZHo0HGZsRwWM6oHiSWIQdhLyl8I5lVbJ5R0liYxB
gtTUU8peWPYNGOZpWdehOA/cBMJzO77F12+zxDrc6YEiJGbFNMjs1QrEG1q8kGQPiVKfRJ1J3/El
s5JkGWQMTHVysH6lkwaha9AEbzNkuUhPP4LTqW7WW8aXIi/VUQxNMTWkgh0PpbSfPEoRhWjiwQVb
xgC9DtIKWx/OUJ6KrXpBhSqqGqH1tt8TBG6JoKRjjIRoa7xbJQwChVX1VYYAAnCqOYBkG2Inhphi
0kirVNAkBPZs6KGTHGuNTTTAXjrcbbdk0W8AOnji/zQMO3vJUitYqHbCXlfv6B8pu/TjqW7CjPcF
Csk3nTl3+uWEo1F5/66hNHFbVJHQfKF+5bf6GFV0fQhsNLPlkE8x44OmxPcgosAiF2h8ZVjwDLIU
s2FSvHqBt2yJ/EDSh1w0nxY33EtuBABPyYuMLjGogHbi3pTmpzd8fO2Dsi7i5HgcfHlcepdXNILl
M4/kku5PlelVaVZXl2nHJ1n0wqkl3JUC4WP8qiqh+EdAzji+uYpTsYVTEv/ImbRnSTSsO0G5SVhj
TQus1q/TG7E9EdF7BGAsrdf1m4R67aHFgevfZm1ty+As5g6Hmq4UVPo5x6H9kvWIFsXf4HYBLgYl
X4xH66gUPB/SFyZKWiWXac5tRYvbI58TAPEkMlPspH+jyzYJ91Si9PQyBS/eQYOR+V7KthTaLtZc
8HizqFBy7nBj/BjxyfLuyaPc9kp2UxrJxcXPJz7er3PgDhnpY/rq+9KjbPMLtsWcjuLAIH5nR9L5
7mZ16KZnctHm27ZbT76punEqD7QIjX3vVQPgjtCB60rVg3bUXN39pI1OSmcG+I5gtprEDI294Jav
fMzQy/lZ9PfWQyzeA8QuutNo3vcDK41w8Lf4Y5GKvymfYNmRKQ8FuamuNA3de079p1smo2Uhz0gA
/8Q3aG9O7LVP3PRuiw72V8kWqRaBbKo1h8cbwhUc3oRItyGJHqlS+jf0q1YD8wF74Zdr1eYWJy9w
lLXPt8J6NagFWITWDwkGcNWiuhw9skMlrKNAayBcpZSWgLlA/ICg3EMTgvF+UURW1aJCw/Qm+NTL
72X4FoBrSlIQx9vlfxS7dYSOjUFPMIYOMu5U+wQP9gCIXKO7jfwdlhCsTi3OmQCoMtdS6RsEUGQw
/w2skD3gruk/MeiCAThzscsN4O4WSy6N57GMqda54Dk5DgxqwGkxaSjaKSH2jovLIVfNMV1MuB2E
WUWvCtxNjX3C1ScTrs3veTbsZOlwptIlDr0RpIwMtZv0qm7V+u2BeVL9TjU0lJ4sOBjrt8e7NHET
wLHrmBzEIt32QdRvXiL44o3frCFQVZOAruBEC8W7LtnMuE5K3oQzEp46DFFAZBsI4RNWEpTipe97
Jag3MaufLy4lRUOUYy4fkGoE6C2R9iyvQFn9IjcnjfwoHJvcjWlaOt6Dg85JfXBG3FjPCEPfap1I
asD+rti1lEua/N82YhBSrUm9Pw+0NKZfozQedjMl82/8JbTbb0lVZeu5RpCrsVU9O4MegijZtl7O
RpbjrKx4qvYPtZ7wWqZ5z0yah7b7KasjlnxOGZsdQlFfc0To9B3YFKMDUAQ+F5QkLO2Yk/Xw9Yt2
nSBEvlcYu1VkC55OQCWWxZTVvWYaNYp3rVB5KetvfZoTOwvAVtAeIi/9xfyLefSko1mY68D2RFCU
Os1xpS9POe2y4i9BKPcNld0QIchKgjYflCIJIMoFXBYYP2PnQDaZVKtG0KCult1bbSA1mmXZ+oul
oBRSpl/IKjAISFUnd3QvXOfrxd61ewJuJCuRsZHXTjtX7BjphWa57Y9O7BUC/zAYGDkLlwAfEOYE
PRuRF2uCLJ+4070aU32aGqNNXhb27cYyCIwdE1z8hb6FthjH3nmXO2NWaUEHf+XEu/NoIVfOaUYt
RtSgi1Xy/BiU59mX+g3AknWhxn2j7k5wrQMSDgQvkx8JeMBXK1qGYHDYmC/8dL6ZUXNK7ax0VLta
OqvjreF4nM6t4+9WHYFkTK/JVORSP4FTj7uFCb3SQTrCxjMF4CMKpM5wauWho2iSQd81U8twzy2m
NK8Lg5d7Jqjy7xYQokV/ZfBc0LdR/JhM5vBckyxxLPIKCsrJ0NLQnVkRYwOeIv9295EicfnRlo3W
w6rn2Ie8JHs+MZwhmf59Ccm0Sow9+5939hMk9TeclDG4DTG6+JreCTAgOBWAVsWxcRAtuqc+Uknp
EMU8wolfw8IYymUHb84C8DV+1T33ZzaTNolcJZOYvDVthaVeEBlRJ0wvQLbmjfE5C0+iw0aPKy8E
HvLc4KmQBKBeDISgSGgljcmQDAaEuim22mOvRrHf878g2M1TdSrAzyZ6ADVjVFmyed0aSPYFXdcC
YkENERN9rmNedvJCdDGx/wXeG9l66OewZDudTUKnGk7Y89n9PKjwzQtctsGKIBQP69kAk1b9PujD
pfEL/plPxgb+L9m3VGNWu3OMXHI4wWO5JgYE1RIFf1TpK+M8VEA6sRkxth6d3IpsqJNKmK+V1TX1
GBdvqG3Q2tYDY9nTG0ZHVtoFTrUqQnbvnKwZhWr2dwlJYKHns2F74d/5v28wor0jhxu3wYweRMBY
o6wUOD3w9YouNO4sIZQaBsS6taepxWvKL7Vj4f+yQUXQ+BBqN1G404dn55QqQ2UY4coDvecgrCHQ
z5xVC7J/OMMEFv4SY+GKKxmpRk/z+GI4m+HxxE2SEJ0gqZZU4jcH8oM5hMm+EN7EfYLrCiXPWtxh
qSPAnSqtVI++S+PezPuk3+4JXbg9fWnu16Xi7oRvZU2QUKMxLw+PIevUI18iUDnJ8WRQwRvPv/kB
5heonsMQ0UgGlXOrQccScJsLoskuDaZz7U3LBnR3G4K4J6+8HowyUYnLJsL0qDPiQ3I08snNBQy9
2wtYayn1m+XlzXg1JjNAMbmi+2e2gUh8r8Nu1LIYYptO3ltZIHgvCsTWkTTkm5yIeoycKPEjdaA4
dMQQTIxcghj6JUSX6SermjFWHkCsO7WjUPgPdin3xluYClj6aW8oXbctZKHWEvAaEuhYhXChzOTo
ibt56N1fMZHl/PqmYgZNDrg/vP3Jzhg4JTDoAYUfaNN12usF4b0FmKC9sFP4Byd5gcn1OUDh1e32
red82NlIEjwHyV9UqGf1CBLT/325ovOz6O0iRvhqwqsVFRe4kc4XDaV/qXDV9co9Jv9v52ed15gX
oJvN3NQlUOHCK9D3SwM4CSKaPGsYdHF37EXd0LoSpVwGanNMfXzXpuwZT+2PNbGc8lOKwUsalB9C
OUaWYNam5wNQ1/HB5At22Ioe9DFCJxMIf2GhLji+3LdnvcPg+uC9/HH12dQ0p4IcJOj17G6EYzep
EAlUAs3U0Bof+1jLtdQ2LqCe2JeVYpFtvRrY1TLuMeOSnnNemWHvBYeOqFDTLA56xBDznUbNnDOA
eGgu3RHsErMkkeIinyOYxk8gQAguv1um4k8nvOyWapfXg5CJZprRq5c4Zumf8whoEVJwAbp5R01n
oEGVSuJGsCQ2HdRp/giHiYTqScnqWWtpdD82PsLX3FSoqKtYHdDtmH/PXuF3qgfc0B7q8CbsD5+9
kDxSYXY/+0qGaBmcblASWw7uLSigFSfclIKp8t+0l/GrvtWC/N+gI/KLIXcKQJxqloM73BUoO79J
xDoW/tEybb5QCwuRLJdu2dViUl50ztSb1LpWuE7z/8FtyHEXDLZoQRMHDXZy881oxWFT69u8ax1q
eCpxJuXM4QVdryCaokaUosAgWOOaETk5QMuN5hGiNYJNeKKxAsepro7x7STiuqds+PD4pcT0/2WD
njDviApN2DeEOU9sPOxmE9smkAGhU9X+CyBP7WcMS9PZicJZtNmt53/GygrZ22UD3vuHHkQXgYST
g1wbqXNTW87r8B9w+O6lS8ms1/KjS7pOnuXTR7Cn8pMdzZ5xQSPkjSAeXH4MrNncBL/H3LS37e2k
SgHkWJ6RMN0FQ05mMMQovgx+9cm8NufeI5E9SjbmCH3Qz0pVmJHhoxnwOMIJF7I0yd8B8rlu/A2n
ru/v+vmQKNeVMi2BFDCpLK5NSWBKjyN0W8aqWW7Wi7T8z8gNhH2GqW3yI7bhih8fRIlSeHq6IRUU
KbAe/2EeET4jUMoJUL1EhwImnV6tNfUQVrzsuyjzwTimlFe4WfPOizZi3lrsh3GrjNdOug7VhAGI
FhJHIRqidY1q6KhsaqXmCYXK3M38cftw2FxuYHjzo8yCYeUS00u8NY/H53XRmlH7aZ/3t1QbPbcx
c3541TR4MWgl4qtxzU6Pds4E91kWp/4pwFyjEdy9th0JQ6A/7qzlCZGFuT5FW/jG3dqDAOmXOJwk
xLHkk5FOcdxFPMcGdWNhX4qbP3HfgfjWsaxjz6iQAoTt46TxMyvxb5bfO1oHtIfWLtMN/QyxzoD8
KoFwDHPVr2Esaqh3YdZWM/6AZ2O2kyXoE7rRpBnPIC7ZjvsfyR1PLR+WZJrzM/w3Xxuc8oVFgRGG
s8N10pglD2Z/4oIg+lxuFL49iQhgwF0YbU3q766zYTIZHxGKpKtY5MfNaN2el7KUmVleQaJjGx8H
QpKnWTP37BdiPqkMo5k5dsLnZBZb5hVbi9Zwtz1oN0ozD8JsoPBOz8n4/AiFapByrpNSO7IEXc2e
NYqYSUgIyaTnnpGKDLbO5A2cil8moRB2c4xLRA7akTVbU8YJEtDEHM5LX0J8HtIbKX0/6jUhaKF1
s7e/2cxsZNY+ko/mC35REzhw32uRHOVuNrM4rF8iDndvb4raZJzCkoUODsvqCOMdoO5+7Bo7mWkp
AhKzhdyCF3JxF3JvITb1nQtRY6wTIQJ2191aS8rxlOJYw+99XmaPtvveJZCYcR2SkIMmHHd7fvNx
8Y7TTqS2GYrTXMlCaGvTjiqf33D4omGiMyPUDMYpxVfM7lGasMt/FQ7MlW3bdV0C275CHC2Q3pJ2
ZyiL549USbxvoIQHDFEXrBN0gIrDvoA+dD9lBzI8iaF616iGFZfQPs1QWwNKx+W/6W7XDTCPxKx1
e1qNxpvQEbb4uY3jSAnaoymBfkEX8sDxR11obtOFOw18J9UKOStCpQ0rZC7eKbbvGrer2/CIzxYy
oudXtqQD7P8Xy0NR0PBnR7W1/SbhU44S3BS1wgbvg0O+fZf9SEL69csQV4onlhnmTlarGCfWbbsA
RLn+CDid2qMCfW5jH3u6BUOvewed9wGrwPF6neVw0AX1QbRIN9tGdziA1J2jKO2nLqoCgH+cw6PY
0Q1ZdW4tj1VyB0mQ7xskKdnMSwjyrBkm3a0QHRGkgOGLfOY4iiyGIoRA0grMpG+tw1CnxzsWd+55
olo7GWT222PdM4k7aqLeA3AhH4uyb0bUZbbMxz5V9rLrcYRCy30FusLWBh2hOFDeqCfSS8tQ3nNy
9chQ3GZ2p36eM1AsEXYBbc5tk0vBJheaCHL7v+6KpOgevFHqVCZiSu7OAiGW3x3fh22NgMDNDQXb
zvgNC3Lb+5l6Ua6mZYGY3eHl9xQ8NMAEZtLOiY5U1olNLVpuRiUM5qdhDzT/d/2czq1PXCVMd4Ns
oBYXh2Z8NkhX0V+HfTw13fnSX3DcwlbaKg3G311NAjByXIPatI7nTqwbercKQOTrJY5bA4Y3qa59
9C4yAtGAGLOvv2JKzIwGaarhD6XIPqxGg9ttJuQt2mxTv3O2iybt1uVP4I8Qh1FMCorwK/XOKlPM
YaZUGj5DKIwX4iNKlP49rDdj6bSK99IBk1RX3ql0MQK2ObpXyLeVqfYQPRxwMSwc3fC/qKrJuo1r
Y9xMLni2csU43snx9TJEmw4aDlSNY6SIIpaJr7vV/Yaecy4jpUwKRI8irrna8LmnWX+gqWBpuYeP
VbrjvPD3ihYB+cMIuvPfWusAiBYGmm4b+7ubGQ3B1YHYtqEGU7AysFeu3v+SFvSedoXcR1QFTkY+
IeRFzcn9AytzOc4XFxOZsRpVN6lgorrq8Yo8U3jSckSh31CobP557SExwrD+rX344insOSNjxEC1
HAyEM3CC/abdVV2Y1pMSK6eOckLHWuqa758itfSzjfrbq2XDmq1wfASWofGbzwHDoFEUMkBtWJLd
QzyoYdn0XvbdA0NKvJ7rkLKTZqXR4Jt7TwFuUZxzDngu+QCWaek7Eq9+8gBUupWqjho+49lvcdSF
pfUSIA6R2EH7ncE+Emm746LM7/O4MrsXLMAetHNr+kdw9/05LDL5f+HnOrgz5GdxJzWw8x2m09H7
hvXmHJBAPIj65IlfSILs2t4z5O8PbSVZZUxSl/9r7OuytJ6MBQo37Hjmt0jNywbQQCvzjF3VwkBR
eIMsCyiKi5wCnMwgI/YxaGnDn+OJmxrKfgV4w2oR7n7w2q5BcovS7xKGwjan4WXo6OP5TbwhqvML
aheJCrasTV9aYugTRTcsVoH8XlbZRJt2YYl50cwqg7DquxophfhXKHmZq324E0FKr3L9S31C8Pzb
D2NzCKt5NvCArsROZgBvIVaAqqd3ZbU0SSQYGHHML3G2CYjORANFGo2XRUfEim0NIgE2AFU19Du9
4JRTr0+DAc7g/BiBoGgDVnVmGxxxdJuQj1osSc/rC4hepGYq2A+aame0hADxS4FsZPMMw+0Km8dN
eFWvW7LnLwunf+IwsjZc/ZvvZTgFes/hNiVvZaCTNHyvDCeMB7qnrbce1MgdD9IgY3iaIh2w80dx
pFgct5Gob2LXTzzVI6+wjoQEh1PzJbNA+3DyUPMAg3rmkzHC59sq2NQth03tr2v1VGgttWsUhyZA
nXnAU/0uQjrQkdJc4M+ignxOvw7kq4h2it9vUnI5xqWYq3cxMK2tXEEj5ihbM+huH6apcSTNGxxb
nfgKCh5C78B26LzktfrgNENvCCkDlAqS1MrShjnSNjCvNIGKbMcu7EAID8kSvDUGSk55Ltg1W1Xb
e81JKaJpTq8NOw8yqSRAJt5dZnsQGgxvO3n4ZOnR9/JCHjQaF+kma/2uDqUNjp2Mx8hQVEAiZBNT
d8km1Ww0sznZoUdPqCn9LpAmJwcUKg5dIVWExMAt/gxZFefsheHIsjFGMrI96doYilXzU9BOauxH
x3NzYxnfEwcDuAPiaYzbBQYDEnE6WymHlpEYfLuoTKNohc14ds0E09a0kv5oLctpwqwd0RUp1U+B
AlZFoHSE5b1A5VqdWXFo+pOBPYaOdDSjnNxFUzWiMBzsPUYKGFWgjNLzGlSbGJVX3GG3vXtcc75Z
kv0Eh2kPul9I+VSaoL8EwCw8HRkhIhlN/fPW3CEmfLP761GRYAufLysC2YqA57fD635cbWqrvWQ1
NBz9/ETjSXO1qtSIDYzu/Mdu6guHuBea1ItvqyxIPdOLUi0wdJujhSxT3HxhYSruuckopA1xvs2A
3OSGlzXxfcAjACS/h9Tamx4nSJE8/SFRvNNC5nG1pqBJ6u2v0BlfmIlAJj7T0Rn9HeA3lJsCny1h
Cb4w1LHddYSPgN+ZN/LB8d7qVp2RnFznpUfMfTvXp5cz+JpkeNzncd1tofh1SvJo/mmLO/0eX3Ba
DpC86vLS3Z8gz+Iz62NWac2HwoOqwauulOdsQUoqGbYz/OEKyDgfMht/QtFhRIVKX66XvZfBFxAj
E90FWEJ6KB14ikNwAdIWce1mo5hFy0uXokdQIQLVv4yEZ3vbO2mQwUF1/+ipZ6nH+rgbypjUjYSI
79K722ZNl0pU0OPPSr4vMy5Y5raMIIk4nXC6q3fgCdBPtsifIqg1IxxsNrnAzsImriE2EOgnSz6A
xFo/V5CdfRs+0OY7WD1iIxzmdJG9JDysWuvYY2XBXMt6lHsGbhs6Tmb8SpRZR8leAWKSDIrj8AZc
KM6b+pJ/BTXnSBqdIRdeO9360O7+zKSgKxXXU39YNqiIo5wIoTVRHtRR0e4PeMCvIaBOGpfzYAUl
ZgTtC3clTdLIqPHcV7HMcscbUrSNlYqIEU3FW3ch2/HnbUzqOerTjM0CwBAAhTWnBOcQORAqSinI
jcs9t2BfvearGcMY8GSlSrRu9TIHMtKv3eyk1ucvqape+rFl9x8I3fLZ1DG6eSfjEsaorIVUUONd
KEFbZoaG1aDgghcLWWq3BY2N0YkQ9i6sucQJerymP+miR3I/2drWNf2AlsyXTLZ42Qo4BnjxOrFK
OW7mI/SM8cTfg5auF3kBnAEK4uny4aK+7CK7AS7WawRZpju9AO47AeBqluEWuZnmk7G1IHocJXfn
TRMBpYh6uRN6o3W8ea0XHLL8rR7XZM/TRmX5nZaxkxVmWXfZi3zfxueZYHuK/7rhBwHox4IHW51o
jKWNZ1JvgWtbEnUBpdzID3dXvHRfQxdUwveL4Iqz4FE1zjxzc9CZ6WbmgEH+acU0wERSp2eoGKTz
G4rmv5kVD4KOfZPufAp7GILKES6mBZEx1w2Eg/DmO0I1H16yHtVpoy1dITDI525F0IUbXJLdzlVN
lBk6Zrf7rJrhK9+YlO5dpwcJynyIuipebzGUm+AoWpyEKFyG0AHVglqUDuUCbQhEneSwqDCOH0P5
xK9OZwy99bqw5+zIAWydflF5iKHUe0wqjKMRwzzLVVpHKUWoYSiDkg/MsQ0egRPUEF13UjEN89xG
Gf7p0obsBGtADm49DESHHKy1obYQ3MA4dS2VNXX2/4pBwETOwX79zwnYSpyMDYFs5Rzs/UBvTb+s
yxbenU3T2xRXMDdwVsjKlgcLkuXDvRojRd19a6QK3ptRcWpIzIMUqBWERhCwzEAsfv0csZSWf1pZ
3z4ufT+ZCbfWSxuzQil0FacvljUw+99WdNahgjMIcYBav+LCfbnopf1cbnqUhnK15lI395T5LBPb
HRA8TahQaA4TUyWCZHkqTGLdmMbV335wMV73TsRliwSs9VYWNMLZt99W4jAH8VUXr5taKd6gsDZa
Y7H3NTFy+enteDxySD6bmvOKgzTvAqAvxO5Hw5f3LAlfwh+QM8G9kMybx+OjfBQPbOCGf/kFB4og
uuudjDGlrvQu2rq90ALJvnGhuPvFZaMubhVw++At+xIS9RU27/MuUq/CJC+eUz9ZNTYvCFF+Dvng
zAjQKYjrldttXzVl1mc7i7CjykAgBTPFrms3x+q3FivqN2IzfldEVej/uJKN8M0HK7bB6NDksE9d
SMmQM3x2ogM3TVGs01Trp3WoSTxTPhvZobuEDmoxzw0XcZ84npp7Ri2VL+ZLu2JhMsIn+k64fnVP
Wwbwzuks63RFFoW7Bo+olgcNO2AXQ+23NavQ8y2xj2hULzJiHkpD6SJ+QHPBGSWTOuTldtxZDAdt
0LWnFJQND3lssMzIJL1Imn7hVF5F27rxkpAykuMbKVInJhB4MZZpri0MEpGI4Gy42J6CJ5y6P1zj
tlhBkPDFbBzg0KIUC9JktV5CP1ZefsVakpz5RBthwEUee3N5/XrYG3duIPJlbjEPkBIcF3zhgw9F
wpHNfJifSBm1wRRjcBS/HlSYkU466/NQlJnZFnNSZ2m0d38AnAj9CPLH6eqaM4OQwNaa5cFgZ3Ei
Wr+LUAE9FZg03cce7sMbwlYkCmEa7RkyhQ7LFFij6B8/Uhl8ExIPwSpNkvn5Q70z9a/XjLFH812e
XePmap3iR0trjDaHF2MQEy+SurGtHVDFvOo0WXmXjg+pxz6b8VcS1h1REjMl4ARMbIDlFiH97tX5
dTMYYSSIrTvRh7el/40u28+I6ChGzpeAQH5mt7O7n3csNl/wL7UFQMT8wHY86wfrND2zbFPeNhb0
+cekSudzYnhxGo08/gGeAaKkHNOWWCn65uym88IhXDwoMHbhrKqWpM+DSEiCvCMNdun3OAWmbJwm
Y7OAiaeeLM3tawjXpNeaSwI4QkOTdJq6WMI6YuTMqr2fll97HzYMgEOqOGl12NuLrr+eQxb0fe2f
GhtwlSBBS7Py5/DywudRyMIzBbohWcu4irzM5jzww9tiEHUuUMv3rqcvj7Ve9h4SVyeVRgyqyejE
bQtVq1S6iR/R3M4/pHN5dd/NoZdrjm7eIho2MruMjePkOFbABHTYnquh2+s9O+uOqXBdsmo65tmu
yS1qEDA+j1o9KRFKxLB8OukLyxt6KUfVPe/qwWliuR0IPbWQhzWbakL1yiI6+rSH0l+39dNCaRBU
68/mfYWPgEP40gyqKX3oBwgoPvrUCQ50H+cjDostQ4CCDqVR+eUFD0IZK6s7d2iIS5/01/Ryc6+s
M+zM1OAsI2ZSirGumIsWmpQCr75JX5wG35TJts4RQW7zzxRuuNSKN45pRnj2XD0GSPRnnpdwD3A4
kENtfzyJv5Ix43ERRExdbCViP6vSKHww0k7xBizKeUO0Qfml9mQWGTPNkL8F6ByaDoIRz4wbyeii
3IRtb25PkerhibEklHEhAwag6rsY67hUGgh3EOndX1Mj9q4jH+r2NFD0V2GaKSuQRHf8xa71SEZw
1Jq152cmulUnWVMOGpNHv76wV12LNhU7WaBqxG1gmrAnQdT9o/OB7GaIiBci5xSYz3Zj6dTLbKBD
jwN4muT+Y9OjN1qbKqWANnu0WLGd8dYdDq/gaK3Zuy6cZB4Y0+KpHyUtXDMV9ad/6LamrIJlhzSN
lofWMBPdrjhOd3KVG7ThV7J100eKYHEjI9MJI4GiDRGrDhWkKcw2onPYbgtGaClajOitTDYV3lFB
Qb/5LBa2xkO06Mz2hTmp5vFU0C86MMm0/R2odaZ0R5Ex5xyaVPC2G4EVk/x7iSA6GLyzgsTbSFxq
eAdI6ED+d8Uf2M63e5xKCGxC8MVUoQNhD/nyZP6mPofxxcP08PcznmBiHAeA8l0IuL1aTfURFqoG
eOzlF0w/HVJ71cPc4U5RZW5jQJbTpNlfhkwJRHn3kHfrlufVolMih8/2FnTrX7TNwBgxK3l7NSqK
GT+3Stql6BnO1rTDk8NlKj0WwkV1XwBsRFt2ZgHN4VDxQ/bbqYOUI1LxiiYUX97PHMYdRH4bF0vC
ru3dX+kAlGeXaMfBMQ+s2fkUN8U//a4qH5GkGk9WPKc62NYglj5qtYAI4UylxtHJ4Zfo0oCTRRmu
R4u5+669TK0uewcMmng4St2dsWA5zTYqhtYCl8hB83g9go6cHyDvo/+Lxy2yA2tKjoMWx6nxAKda
qKqKXWGy8t0wM/nk6YJIRKuzmYWzAbgO2CQAhhiiT382X7JT3vZllqBwd5J1vS6nOy4vCGYRNjQy
roRS3Tpj8Hk7izV6gTkzu8aP+vUYMqhiAO40qVB2R/vev28tgAiKGj5Zv9M8h0v7AOSiwblzN3+G
g1YHov+ICyPX6R+QOE+dJzGhBElPYBiqk7nRDNWhI6bdwlMPhpLXFsMeCMEAQKjKX0s8YHLVOkj+
F4ZkTM9aN2CWoFgWGa2Idxyc1h3rIZUc0zPrTIu1Q+VMLN3ebcw/QZLDjvRm3vD2EP3/YkttrUpV
4EyhF81k8XrC403hZHTwbgj+AxnQ4XTVNM0Lw+NRpGfeAtGXA85AlldjV0oaEmmrFhVSFEdHwm0u
XpFD5kfdY1IuNslsHP/fuCnpXYu45GPOuXOksUw12BJZqp8DAUoB1QoyZTMULXD/PXZZ3eMfspWz
R2+K4kragRBAwieyx7taBzm4KgXJrf/R1dEvS8g7NEZkh17Vg9jNpmINrtO9FbHam9fBITi4k5/j
fFLNSJmOZTCHZ5YcH0syhExD9UinGNjfNRK/zgX1TtP0YJIgWcXi51xYwckwj9oxtSM84xNi8LF2
zEDFHZGxTAYFJt6635UUMp95h+0hxFUkykixX6R2IwmlExoX8PmSzKm9sIVRi5CqpnPJGl08PcL2
MqjWijLx4D26vqOR08KqnNazNcjRqEwxXeiopOdpdGTA8XyCPkV4K3Kq3e6zE94Jf7kpsAjVFmWM
Gb3oO1iYqJ1PIZlrlkSCewx69zJY2bqqrU2mMx+f2KtFQPj400/M6ITZUGJxZxDbjdUN9/FcGZFH
ixZN77VxofI66XsbjwxyXdcaG+K+TmSdIUg6SF353a+LgtLZIAvBZ/s+lv+c+jh9XkF0gzOIatzI
eb6iugSRh3YSy8teVQAhWLELjY6QYbHeXyoU++GHlqh9MbKuKL0xeYX/coYSlWvaRi850vJY/I6S
PmJQ8YWnveVOD+L1680lWssFnioqF7YXuFSmyd2YokvIo+26A6so9S/FqJQ+bFnkaIsNMNAAh6Bm
U5kHNeNm11y3qnA3ijDImUjBAZWG76X2wko6AKjRU/XAxt1nKAU44T4LGdA+Y6KBiE/55u4WeIJG
NI9DT40jPhkVl+vAWjLhRnjzRsWK+gQ+8gp1Mkj6gUnAuMu2/LQP9hWDpbv1wOYcAsXH1vYyOfwO
ys+uTeUV5NsIhsOtQ8/fapjuHYSfTxqcxTpAX2HWDSDBa5VXqI3dLLPhYFwSExDMsipe2KGpfKh1
njPE8mayz7ATcbOmJeeYYpR7Bbq75kr4/f0SH/I+4uFmUTO7EJ2xvrv77530XNeSseDdmGhArg+2
NnIddLrPa4qUudU0eHII6pzZ9FN2Onj2nTa+2WeVl3ibgmToxrsMklTBXA+pXSHZdHsfvtQagDxK
4GRYRi9AR5flbxPm7OjBGwVN0VVv3s9MzRAc0mRAYdna4oybe7D2U+xU2WBItVg9B5zE/GK5ucn8
6buswJ5GciHZLZ6h3bYmldOP+ns4+wqFi1aD25uH3rk/aN1gO9Bxt6FQqlauORReJxJd9C7fzf5Y
snHReN+iWuedJYiyj7KT5FLtoQTFC8h+jRgWfTH5KRC8lwRnAErmC7E1rvDL8BZbXmorM4OJPXEo
B86N+g8OkjvPn2mDhcZSiFTroCVbKFmdICPP/gfjivVUz9n3SLWgYJQjhMfp9x5suHLAgCA7gpAW
fcBihZF4Q3OV4AckjqLGQp9QZjHTpzDnOizUwp9jU4DKtp6yyDDp6/7HNf0Wi9kGw2+TxuRz9qv+
mDyRFi6SF0Tft9uFWRHoO1qmq55uSH7NhHFfCw+exNo+pNeQ4tSx+OePE8XqFwi2JIQnZAdFRaTS
tH5ERZPT2Avo3gQnx01cy5MHUhu1AeSC7uWRf+kzI2yM/Sm5FW4qzLJZm5J1CU8mfaR8aq4yqyNa
yxpQiqOeT56N27CKHLZlYac3hFCf1BB0bhPeVpLaFVV/mK7Oxt5Xu3jxUpOSzVk2bl6mRRPKkF92
TSzTXufmvtH3AyYsbTSUlnkLSq68AGS8TsnWqruOdM1Y/uFeVDA3Lg36i8LspnQFpMuySDNrmMhk
tePINSTT1nAOOKlCZcKUwJAlUWdFHy1+/EQk0+GrkFqusX4GiTh+Ew+6tvXgTmuTwzUtnZAfDaIr
SqvFADEdo6vaIgbah5lF4bQTFSFXd3va4j9CIVkq4jgDyVDsID9qiN6LwEE2JJJt4uD4efZ0Dv+8
R+cvPX9yb30nuRqMP2mQKo/z1FkS+IpWndHCuoUqXhPF8VK4JeJEHMCI/5WTr9uH5Y7akmHHQCHK
76HKGFk5OBMny0BG+vBM6XS11vHhH0pFTB+374qgm37EMiFcQCHhP7NY9YSKU0MAk7UormUMUMd4
tuT9Vh+MIg0VyRFScpaQ0vHfV5DWACulEvO5ZCJGDKDhG6Ne78ZtrIo4wEsG8RYjE1PkujogG4qt
rpseUdelcax0XfLNChnPFgRYZjl3v9BjT4lCDpUOAzb2xi8XMjJgfRog0paBR1L5S6fJlj4gZekZ
N9Yc+KKBGK/irIvPu5to/Zy06eK+icoJuPW0VyA2A0OSS6tL/7RX0XAJ8IGzrAd+FlrKesk0f6dd
evhxV7gHHLS2uhhAwLEVOh0Ua4zRekiU4vvuOXwlweR44KMb9InlGG62VJTN3EXY+cA1lXsSa4wb
9ykdiQTkmuq4XCu1C1qsU3sYy7f8vNHDf9VRT1KNs+RmJzEbvd4Fd6nOXGJp8/MPN4yysZUiR6Ch
RRBTCdf/6VVTQKMsydAk92iT7KWZnFPlSfJdJdO+crxJe1KFyS4LZa9ZoZvdRRsHBk0GsAYaTJy2
hVAejQMPFko7TXZbbXw/ggMuxXVWyYsv3Tmf9lwfniAyQxNrPf/U1DTGnY3WXoSmINqf49v+jx60
NMWWw8JlkrEWD8LVfbBeZ43B7J+zIbgU6claM8QEP98Qn7kP4NvfN3qLaZm2DjaXAAyoGM0EQ9Dd
YYb1II+j6rtD2btak+01dVXfjFdGGSv9waggiX8cFWoaOIHOPNtUAucO9qUb3a3+Z1Rv/gv36NFp
z8pz9nKSvRy0JEyqzAVv6FxxVs5MlkBLOPbPbKEPLm5dNl4rTYXcVr29rOoOriPJsyrKAaXniFcX
WTP07riIcLxxiXE+nKBf4qay8eBeWLcDprXeKq4Uu3aQkQ/mEbUoy+rfIubTV55xBOMtgoM0c4zU
JYipPHI3kGgJvMNYqAxKxYTel+rU80Qq9nM0WV/SgH6iDwOPe1FQuoLSN/wsfnwtiIMVfGP3o9CR
FU7ERL5p271blA/oGWIIXD1LfGEIGJM8IpeHb+JskxdSBQrSJIWhEOe3VE2YhW71F+RB/ssgUVHU
CRyk7lbItdvZg6imoU2vKae1JNufm8jWeC6QkhiE0xeI1Rhzr9EW4GNXA18FnIoRc2oJ2F3F37Eh
aFIvtEa4Guq96f6IIT//ZvkZTeooiV918pgeeEWKGMZweynTpW5Hah13auLIUCHsjOQANxCDKeW1
2/pToLk2QbDdbNm568U3RSn67+BwJxEAG1+C2AA50cy3h1VNJJscvHHKhE7a0F0I0EYp/4oh0eLf
XBI/WdK/MB+Vomfyv9pHfp2Llj3/xbuxdWNIg1uYRt4QyyTL6cpMJRrdhc3qPtt4DyCElAcK5L6q
45qcmkufVlYTUa2DjeSojoGZeHNlAOLTiTGqnRV0KrNocqAKq799NXg9vjBHOYcSXnFl15101B3U
DP/3UcE8zNnr45oNHekhQs2ldmRy4BXt7I5r2mo4AVza5nX0fqYm5d3676j5Gz2vZhydUBNjUh2H
WhvmrsO2BUWcoWiovfu0Z/KYAAOJOuYLf3dmi7tdm/af5GeIxrOa8uKBWaPhbZ91jc9C2Y3/lLIy
dnjJr9JuASQLQQeFTzqdtBVuoeLwwgABvYmBlcpAC8dDkAW64GAM0Xt0VE/SxmdDNO89Tyfmg1du
cSGphRRVIHVv+Jy+U1TQbQ0O9GoqLh8Tm7xFMYOsNMWe/iFle9USYfzxN9nb65f3DyyeBxutuqH5
G1Y/IhECFzE4lleIy3OtS75NXVfQHGagCII0cUYIOeAJwbCSDxunGkpnrTRuDQ3BsG7zpDj6I5lD
KsjmkpMgxozN+UIb1Ecx4ebN8xqntqZVLxQo2iHSpCONxEMCZTRd3AYoEc6e+Ap3zwSvMEFqx64E
mxBvDYQy4APgmKZVlLoQ9BBjm7bYdtUw7TZRvYRegteQqSBVojRJOh85/JOcvrlwreIJTG8PVK4+
Ft5073arWlR72n6qamD1wDEhfT5o1/5bJRQyKAaQoSZYnAjswHQMx1qb6QzBfzDFTboaI0CIvY5U
IhG9xaEw/1RwbuLziK7YCP5eUWXzMxQXcOz2PL/GEgxZFv6zSvkgXu23CncsUntrbF9tgwcIOo8M
JxJvqQ/r+FhAx2sWfbwYnxCKQx+ZmEb/LVuZE81pfGEyS9us0Z3W7fffho0YRqzh7nB+7WfiftF9
0xZklXuGdHY5amlf5G2JAjsLThxL1+o6JhyfWF7DdtGNRFgDwGlEpYZrN4WJmNgv68NwwTouqtnB
9rCSNZ7s9ih3Ue0U5rsY24rZecDNIPX1XxPvarBL1zurVfh90eulZzmGGhehfbxM65YPjgyjoE4P
KnzTt9ugySMTT9VeRvrNK43/hQGKsIyYtmTtScz3iApGWbwWB5nDBy+TIuCjO2TGVvsv4I5WCltd
e/Oz2eVumL/bHyZA0DnqbZU7B0IfmNgIsDW9Z/79fWIS07knO8h4RTw43Jp55yat0iIs3psU1cxq
SWqrP27zxQ3pu8/Duz33YLEuxEP9jITSBhqEJe1Fx2/Zh4Y+yZUWOAzqkk1Ru6i6tV1Y7Z1XNWPg
qm2OSj9ZD03IjHT9KsMaqjjFx5NGHf3sO+nptNAjVfEuFKFOm60rbuwZkM8Zo5GPGtBq2V2Grzv9
269Vlgkuw4xH0kk+Y2mkeakjwOWbIjk2jus/V3qh6RPLYOp8uQY34VcgdcqWaJb6zJ9bnXHMZLy7
hjZFXRz3kuOcXMARZGsTnwBnWK7a8AoJRJn95FLRrnTREVKciH3Pgq3UTf9A/dCs+EYZI/QwUW49
uCj9Vqc57vVoEEFI39BMJpJSFIjg1j5iwpLh7FkQkv47Vy6BmyjN0vvUEUsISOSizTeYgCRV+EYW
6xyhZ44LwDm+mOuWgXvzeCu1RPJN/HMt04t1GeQuEKaT9T1OTzFQfY21L/A0sCWRItUTHAVouiJX
18jWyEnKUqvv3SnMX2oDKTRgszKCG1RjBJsKRZHM+BKaDRRz1wtM2ochcG0Ch4fP1yGZt3I1qpBf
Gzk0Jvq7zTFhv/77AuhwMcykN/4EWsq7vZPpApUXvTVNC9i+q4FHKxGr9M0Bhh5e5VgmkEU4OirF
Fp1+BQiCEFw3/A8CvV4uz60jtdaW/Das00CZdAEF2sgJPFB8fWLoLq+kz/4GeheSn6QxmKsp78Ox
tvgrlMnDBG5o0G5MtkMZfRfTRVhWkh/CsP41cwmbFi6eeHWup9unTwn+nHeu0RyxvaItBLZkICzX
xcx3LWpAyT3M0PmxzlCxyioXbYFJntdLEy/o/fryEDbcI6z0ZASrHvnw6924X6srvYm47cWjmMxw
QlKzjJMwJUltjgcwpOsNxjYjJMd/fumqMYhvGNiCLxD9UegRNIXjPzfEQocp4CXmCubhuq2dpklz
Cq8EOYwAs2x4KOFptKEPtFQUUmte9GFPTCscGpA42kODYY37kXU5akQY1fpm5m9ROQsaBy9dozRl
MTVVEww1Sz+aHpk55/j08Kln6L0/S5YM5iRdQNCnjjx8+HNzUkn/WjSx+Kk3s0vxf9Pl62RSI2yZ
KeTjChT+FiTvHmmURnk1JNsejgk6aAdt6Q2rlppThr59VP5r+28OpmNtGdJl3QjX2JuGaBjjkC0J
HjkZLax7X+2O3NSK83lAFq+YEnRPwXplRacMeR8p1C/HfLgJCeYVoZXpfktZbpgdlMXE1VCBN1l/
ZsIH/JO6Sg9TEwiHP3ABkNSEdmQFugng443fT9vyrVTIS2/ITKkCU1zvqebj55Rd9pl+gBNHq0WO
lBdYWXV1WpQXsTCYqJEdkYrfZL8nksFFtjaNdS9Q/AE2WVv+t9VVP/TwWynP7Pfw/MyoPkD9q0rs
5REs+PcFrDojFEtZlyb6lmrAyXuueikG/C1O9tigXlvijSrs1nKg7OsramvDIzLtwvy5v6OIy35O
iWVUBrkl+sri/v1Ws7UbJZO2aE0IH4QOhaGy95Lt9q7vFECjjqi9Caxo96S3/NyuObeD1U5N+UdU
zhFrfEq9U5Z9BI/Fz+vlxiD23HBBNqKCiP65KWILluq8Ob57QaaapZwltGVThHEffVBHst3K9iTw
ukz/UDIOTpi4IwALSlOZI6cMxUSqmyIqvphJ4+KcrfGg4MTNoaoNX2e4Ubr4GV9j5I4jET0ojvrI
0BO/TaQzlC9A5BrFPaZWAmBUbgApbMFfWIR0ruAzSmQ76TnsPfXtdONUDAfKx85xQdp6o9Wpbo5T
cDkD4salRjjwY2vSfu6qozy6Vw2ENwHvgVIzg+Vje6s8RvYofEwoCBD9TJQK9OzRGMp2MINMCzA6
Fus3FwQGLWoWHqFu/Y2PO7NPhQB76kk02+bHGtcsTx7bPqxWF3eKVpZTHvkITepAgblPFjnWn7Gj
sNG3u0V+biD3fwKbvyHGnGpp1grpwGdEES5XCjtRfrwQtAf+h1a88UKDuhQX9G9NiN86K1KpS5NP
AMKXImBkI7hQIVG9TdKW9JnyddrtZsPoSTR/VGpxlZMTyi06OvV0d6FTJyU5iol8mwyP6qDRzlVz
t7ERsjoKa/4XDUhZ/c3+vYOqkpjVtMIXLbzUb0+cYPNZ8egnGD6JMFRYQuxeDe0wbRv0ieLOkIlW
R6vqmcquyYgL/WS9IpMGq9+rl7uxz1Xm87G3roHdkFIhrkZ/asohoYb6TcM7IiYpkjN6NubPQowD
OTw8rh0q48Wz4mSXDd88gO0D7clpnkNcPqShZREN6cIXoT3AWMzHt+KzcbujfeipIAoiONyRBqWY
WgdxGRi1NZpcr2VRcxp3mLzZxBiDHSQCi03gzJN0E3fOw41Zj+HYlQJBzHvZtjLusK059vXTAF1T
PrfgG0O0My5OOuaO7gJG3aL2YmHtZdMQkekbI6Mbr+uB4GPWvcew+etRrZrb6ckUbWibI9wVDNoW
I9WTljLF6OiAthj1ehMqvo2Hr2aOOYVZTCf5DvcjRmann57cRo8KgDBCsUPGRUdzDCL/MWJPFXXj
J84NE6OU+qyCRi+J4zpqmt20L8AACzqBH1dFotlxI1F+KczcIp2OS60Y3hScS1J5yhufyqqeyYuq
KlBEQCHpin53Yh90Bhd/rmC89XncpK2Y8YBTVhhfUgQ8vGeMJxpOvsrCEOWOFDOkN9yL/o2hvWRw
FiFP/PuLBynxbdTYBIOFt+0OeVtM94dt4gj8lSikWKWuuvcWAm1EuK+XI9lupQVK8/5ZILeeOBEL
FaQSYLZAPlf7DHFBBGV+sng4MxXlWtu4PBoGSPbIjNNUwBpWt5+vEZ0oq7C1nuhZ9NW6aOsRmPsg
jdjQFlJHwGQfjB9weG+1FG2R6Q8h+1Y/PbbYYigYtVwJHzQmiqozMRKGu7jAK0m9yi/5Eznp7HIT
HNGK3EuuGMan+Q9n9C5mpXMuyzkpAJ7Ubk1WT9SZ9qWcU5Z3bDWOV7EPJtFETuwgkQ6kgu26tFKE
iyKpSRlfy1kDnPhdu5lOtI2JORfATlHKrgaRXkrR/eI9Aurvkxbe28RXC0o4mcGPU4NPzKpa2JAI
QIeIr4ls8i94GJYW2om5hTO2ACkFezZrWAheqFArkUkDA8tSpRec5PWJRGoz8sr8BQFjTjsXu6Ii
Oe0mrZ4Rk0zRZjO66//mj/uLQJJpGDtBJMxZqRQY+7aH3Y5qy8j3pol/cjqETjm5nm9f6QWJRcMU
VQwJKF+diaH1jWE9SNwP+F1N2LbKZ2+W2h1d0/NC6kiOOlXSKOrg+ZSm5ZLVFPbt+klWxC1XSLW0
xmZ5zXdHJsou8GRq4cZVoprdTjNCOKA9YVBBUyUfC4DrjNEJ2mHBZnNY+uXijYAVuhPSY9Cki0fv
SGNsAVGw9aPOemy1OR0e59i0tpcsNHtluqtdDXoyQf5fD+03e4gRso0yVy2yYKLdKsvcPCwDQiXK
W8DkV3ddpvHaoffjTzq9iVvUKsUPxUxI3gi4ZqsHzYj5KXHSYacbytelJkMNoyNDzqwKqRvguZba
45oNWwM9UTj1XWFI0lAQg17wlXNzH6pGNp/Q6+MLG3ujYXdepdy2c39lqagrnvXrPLvcVF67j6lG
uMg69eu3FK9OIiaEa5UIWpohvLfBCslauLkc2OlYg600sBoQy1ARy7uKb7HSV6TBu3YTJK3HZLF7
JV7YpJA4Eqw29pClJl9qV2e7mS0YvplbMZMVMB4Ve+PUnInJOBTD5Qt7n/y7adK1VmsZVCyuIjaV
gdz5/jbb/a4dWydOhWXjWAwR79SkuQus7bBafmNETXmzx/bEM+hIKzYCTsV60fVePzSoGOQ2PA7m
lKoEGIhJv2aYP9Yju44bnNBCLMtKmsDUMai74KYwSu+4t06PzgnlpnvMfCZBVOIr2omC+HOc8/DD
Qx05d+sDM3XUREg6xiPm2ZN6Iy5VkDrXnQa47x5oW3rUvIxZ+d25ZMe+Dgl1AV7vm7JPmqIPAs1Z
RFg+f+jcWeF0MuKeA8aPqoYzPckdiQN/J3D3u5BgWeeU74Wo8TlWpvaT2a1qjB9ICjmL97HedUgo
Kwz4yeLZ8JZN6Rkvp/QWZuNLlVXb2p6pcVTWaFKZKj9e7E2D4WeMGDg1aAYeAMmuUO1KxNi9qEia
VH5S3XiUMR9/AZFLdFXJiKHs0WHe/nUMcL5MhIbs1kfHOcfObUrEvOc7pIZIg4X+PfM6viIP75DZ
2yciBTxGmkvZMnWp0QydrOpQApir0DFMsg18tlwFVjIhPabbu+HHUtQUHU394bGJEi0T2SPupXmC
LSvnP8v/BU3ueNFp5JYnUVxjW7d7PjTm4PCeRPeitOdis0byX4JjUys7o4RlGuMvGhu4Ym8tz57H
8rIgIlsN9+ocHcHA5KxVEX9qrlb9+7m4sp9L8tNHwu1Q1D7bbKFeWir2R7dnhgz5VFw5Lg9Deitc
sWFm++ADyKrjLOxCqnl5tiVwchZkxpnaMVMOMXgPmF/1uOcHWfEpvj8b4FDVP3+n9MTIOa+wNfdO
e/d2MNLwca2lAF6hfT9yKWVZCmDl6ck9BNYmipYvEhNOeX6eOTUQRpICVawmLlqNlUtuvbzJwpNc
7A35JLE4AEGpXDVBf872ax4lbe3sP2+tA+lSmhvkRTZqr35XqXGuK828652LcDpNOedRZnaisw4a
hjmbLBbcCBlsPGGGAgUqt02o7CdfnS3BaUxGldtowfjJLs4jKbKWDdqmboLBlbGRVy9kyUkgFtUW
9oTV126rN4kcDzQ2vNR8PH445pJ7G7X5NH3q2BYUkLsDS49MCzR4P7J3yTZ8t1EXYgTGkEd1Gw3/
lzRrIqRSh6rO5qowtVEjOCmte27L8Rjb3eqpVVPuG9TSA5ItkZDYDtgCy3afNb1EAOkBiH8LbaPP
alwZZx1nw6F/nKLHKPpAn7+Ww7YXjhfzwMJOzETHAC7fHXtuKZ5IWZof/CBwygiJLU6ltmHDT6G0
RV+e1fgcyabbYWW0UkON+akgfTMeCvO5Xmyr93JQIFEg1UhTRLCQMn/YSJ52+hW4nAgJ10B6zslA
CDtQL4zl69vjJFV38SOZSgD0bbDCt3+0rJUPnXwEhH4vweKpC5nT4RiL8tOMPApBB4a2KOJ7d58o
UqY4WtwQ3JHblY1Fs6Ypz0sAQka1msbjAl0kFQT+lrFQTMmOtoN+XbEWzUEG3tBghlMRZ9Zq2cn4
kTGPTnBNzNh6tOXOAQa8aCi9XJoDMvYYUlZxQ/v+3NzRzI00XVUJnzD7sDwXmn9fb64BVN8YBO5Q
I7gLGM28R3Ffk4VjCRfHBe3lS4wcGL7cC8q1nwND+L/Qi8xprtKyGSMeGF3W/dtHwWmNCqI4Iz+O
rXNFQXHUUD/qVmzH8HIROdK0g4L6IcOZ//A/4n/5YsCt2CXFCpe9O8RzwVLIiK0yohcUX4dQzQ2C
zoI1Lx9K9NmC1pjoKVO01sPme+MMJOaYXn9CllyFy/HpkDeJGEcRr2EIdIghX+1iBBrU9D/qQ3yY
kL5RNmBDZhfJP2woc5Trbg3RpXpgkUamX6dRFhZwX6WGWfvRatTZj/oyjm1Ei9QQu44zG7gELofc
wGLkPzN4tjFrRkY4prUp/frAUt5O1fCE860CaG5TrntVG2cxDipRbQ5k4tdqSvbCQZ+yE54PBEgm
tPlP5Ev3wFw5WG3HgWrPvAgIJmh8Hiuk8um6x9egmiz2ToH0aqc5csw1Nq5dhhK40PeSvnnUZM4D
XK9cihQ8iTAn7G3Jyl4SVjXJwJc4xy2RbbEEGTqILjHjhOcCO+KkbbP0xi5UWB5kWHPU6GrvhSve
i/N+9t+MzuGs9fYImO7tGoo75lbo6x3aoqn6UYpKohRtgin47VM7/p1Ms0QYNmACDBz2FxDT29FQ
qNwYkv/4PgGVdQsEEZeSimABj+xNDW2GAwLM/HdYaVsBQjRBW8lP1Mmug4cVezBD62B+Bz/2fGaH
eOdt7SGyqVOTxLwH/zMdKpdymogYXhw99q3VtTRtlURcd91TEeiUNQhZcz52IfZyoKRA9GhpfvLa
ATkb+vowLSirnrpTp6qtb5fqe24qA9lx0arTlbe1Si7lZV5jcVf22MmnOnSG7dKLu3qF4uGMOdz/
zJPF/Cg1eoOLUAMDbW7utW3BbhMTMUXhiM/nF+tDYyweM3mqw36CxGstaq83stZaixXGWj6wKsBP
vadPP8gJIdBmqKlCMDYgtcEtjEJYsCYupRmAm9mZBTZuhNO8OBNVjkFa4qPMSts9e2jKpg5KssZA
jb8P8JhJEUUynVqM1NE1YRu5ozfWKTOj5/xVXjnsjBaPvIue3I4Ohfw+Z0wDIV14sTk8MbGYy27e
tNDFAHzFukUtd0ALZRgmFxLva32QTqrTkhc07dH4LFr3NB/PVcrtlpxp9wEN4WMUImnIFk/++7z7
GeR0N1ho9OiBp7f1eEn9f1iW82GdMg1+oQaykd0gS4g6Ei10Y5dSi5J9kyEoVljFr4y/RtORF2y8
yXRMcYYb841//rfoTCXTbEz8c/F+xQs2F0+iX0zpM3cAo+DmT+/zGEAg5IeAfOJqJmTVm509WcIb
LLsLDasO066ptkc1kZLG6Il7UgMwIhNxwEK045SwHMx+Ls22oiXvoI6qPwPxZ7KzU95MIawxHR3f
daic1IvfF7uDEXINPcurDL64tfrlV8aBByQZNSFon/y8J51zMFQrT0olwrUoh4O9YXlizT0uWHOi
7gt1lYphspLPHjqLNK3htz2jV/zzRY/L5pVMnQB6heHCe1NLYUXLnI/3iMXgCO+VamLP/4zJPeOs
lXleCvEB5vHG2AWn1g5ogGy+NjwsoAKeV8Er00Ih4SuVv4INIQDCh4O6TxGZsgHWGxpc/nVUG3lR
94ZpaBUHF21pdwTbVctzy2l5j+/+eKgGpxxwG2IiqLvp4UvY/h+lAOU1HQF5vhqtYtCqnPmxacud
h9CPWLkscTCmFtddtF1Z58cvjqjUMmJBm33NlKkdR4ELj5vW/2ZIDjyfYiNiOpsyi2EFhzVoUmlB
g/C6Y1w105y9GwRl5+GCLnyJ6CTw7fHQjCkkJaggU5QT/QYPK4Mdn+2QMtDsSkWQS1Shb5m1ztWZ
Howl2o7P8Li+nwqLDxZkZ7I8s+Rpaif9I4CJM5Tk77czUBdgLDWkladM9ow8jhnRIy788g+8n0GL
AZuZBRaerOgVuF4e/B09w8ShLoacHkhJ8mGZ1YqcpFXaIbNIhVZCI18Kv3ZMGMsnk93HlPsf/8pT
1niSvwaTIcGkHuYKYf5xGSn8ZQdGGH5fireAP3vbBAZsNQnwmpPgS2F1oZUgYnU9ejUydaYsLUjK
5mTXLgd4gX0445XhHwGXDXANoXXuw/I0HOcavPb/tNGGIOOWIKyDm1P1T/jyjsgotb6dBmCtSStD
qlhyhwx3G/E8NK+2gBu8AZdxNiFXfzySXxqD9pLICzxL03qMaKBxKzxioqoMPhiPCJCoI/txoZBZ
FkRoWxjdaCluKga7Fa1Fr59jmYK0SYHMunqSYtvCdi9BPM0ADwNXvNZlRLTAdzCIuYUd4P1jjRMQ
q3vKRripx1jk6U3PWYL1rNraLTAyJso+/JhTkARaOSaebrp6h23XPXWnpteOLFNms6KWUE++4ExO
sim0MP8xjQzHI6RX7+VdlakLXSdKs9vbuxRXb9Bgjp/4HYOuFzVH2G/iMUmuFYk4t1tgL2t8Ch1i
a00kyyFg0z6dA6SythIMIoa8S8X+qQv+NMHJSXA+WCwqTSE6VbiXlgrH4g42u2fNYfHX242HA8ZJ
66TjbToT+1QH3AXDFaKyR1OI4/ZCMY545ArDC3ciT8Q9WPAt3sKvEcw/h2vLXV7Y+Vg2rfkYNBmH
4WL5VUzQTlVKQXVe24Qzm0axy4paipPWFTyFkFBUqDPDtfwvftIm0wYYl8LIinAzG/F3grCZCYPD
ANFF733d2LU+K89UI23PcItTUE98NbZr06xt73HrVmBmY57I+2r5NZLW6yf+GlzRbvQMvGIy5rPl
rHMlpxYmk3UdNsq/QvO+Q0QFB+ttHE4d1odvcMCtEv4eyc9qwxrbqn9VySFj3ywI2nTtUZkZEZIk
fyRcwX5J1M5ciLbHSkC/lpeCan6N91ezLkH8Ky3xLjkpOu0wrmgE41uFc2mM187YeEK50BpjCMPr
NTulil4aezFPw2LDAXvdy3AnekOMqgBUD4p5+WqA0InOoMnaHxBLLAX/7EUWZEsCbwa4MVcrJYXl
68TTc4jk0TS+m7k1rNPylIIuP4Be9UH3k8+9EGcXcbHo8xXtLLOdPsJY7c2jCuSLJTT0wIkaoRU8
uejIw/cqzRrTBGhLVFdvSZDGrXUHsgz9e0M5pHD+PDRoKk1k2pNuYt7RtylCe5Os/EJk6AOFTCBT
qDy2nCawzImMykU7+BbnKuDg7qNZXedrk7+MJfxwPsPKDG0FAA0Z8SatAhlccGo0ztBwxWssth8k
d8BGeUuShYQPGkWOPJV4MAxr8/WGAAKu8hJt8zk/T5CbiHHSZ7WNoL1oRQ04aB/WyI1PmX7gGX+a
APY+pMrFCm5efbbME/+9ZHWS1z2lJHeMpUZXc6T+uJPmaRVYjEdnJCzF8gXr0xEpQLMpiy4jZ5PV
4EhXc5XdUUepm7baJfu1mJ76hlZLUkqx157tnc3EnteppbIlEhetloLKVoIGFVylmD+9XKe37cIo
N9MrcL1o57X2/KE+ecil5iTunYK6Gh/n45YuKNpFMMmN12QzoUAighCTEdm8qkXGSdVQQL8smGnq
VJ8YmkEbImxFnQMTQ5ywPlOqPqYYMyMICrwQ049gfCt6CUq8BmJJeZ3YdttLXqM+r/b/jZqyx4wL
Tlq5J8PzYLDim1eXC4ao742yecBGhwAOkQojaomwfltRTOj/GC1k4QejM8uVHiG3s878DCjKrap4
Bmkvq2hWFHsGEYC3vnDjGDRKbSFIFi36nT5dXEwXYMiqtmx24crf1s9a2ye5XSggoVjHJkTZ3kdY
lr4DSUxawhpzLKSVqWnwAraXLoGsOWPWmJyJl8rTDce2h4PlPBNkCLQDk9+K6LunUhMT3eciUgY3
5gKyoVyfYn2ZusFb6BECGBkOi0muGzVeYgUIPK+68qiZEX+B2+hrh+oVCnFNanuW+586smnlu1Rf
W6f/wbv99Sfmgzg6HWPmtaUFOgSKZfsg90squhj3PCAlIGYeTAZYFla/CnQsawfN2rzUcx363pEt
DxoH5y+CotV8GQthjyJs/F5C7HP0ws2wdvPJunYL0E9F8qHDpOmus+MOdtV4UM7VCC4aExOgU132
BRaHwMZQClAL51hmY9/zJTx2a1dKCGf1ArqqM/UUgImoM8R7xoq+KQkVuzI0TVAxAEyfPF2CZFFs
z/+04g2DdF/gFnAHZ2pastulZpA3+oGGsCKA9ePLHn6aa1wuDVou8BdSOvt2w58myE1mxsdLmGkQ
PN7/bf5CDpJzQ1ttSOOXPgkJLEVSft6Ap9ejbwEcgehst2O70kRrFXa6lfEX4MjlH4pmD90wHlXS
0SrgUKcqqszgP1qY1eWOcuA84N9ZTTz0fc2BHlA/HUBNNGnN5zRpsuYyiK/uAhBx8SjA4Sain9bE
JuSuSErWWJpDLTNLep/+W2zCqn3jxPEbxxNMsB+07szioc4cAldwgT1LiBlFHIUKE1QWOKk5VvRv
3cu1lYqugwE8IIT5nnO9koqqm/GtI9Lvp4GVbaGTR1CHagIiPevR2ZxBdypc1NEHmSZGVAZ/1X3L
Tm7Io/0NAeFfgw0Zf3uS62HmTZ8m3OOM8r93UTJqwYe8rMe+6dwQrXulAg2Z8z2h5eGL8R3f7mNC
BIHssMDy95peuRaPFKp2Owq9klClYRln9tbO41FXxS2ZFVPI6hYiLm0YSZDUUY8CiPi9Z7gLhKxP
WbkT1BAOAevDqJQiwyszkS3Sf+MZjvFwEJhWoW86hVVtkeWaKKnBWhReCzOvUifk3jmiolVo2KjP
dM8ja9YHZfnckT661sWCXxNkpNdGNVaIT/zaXDWjbJHzGUn73y2kHHAcKtwrZ6tjlX4TO8aA7F5x
gnyIl9U5ZSUOcqI8TA0CbyUeOwge7ze2h9vJBB5gmzlw5AmQTIQ12QFawOVDPLVSD2RygP5OBrgu
MBLR7/giCLqKzrU//4ChKpnjtvBKKJSU5VwYEdoiczfYzDO3zGGN/QuP+ASgN0xCPPLg9vIKqkEL
GA+4lmarsXUndrBdYOJ9T53CC4ZP+GEMDORhpCJZ/SyGCM3TllObPXVkqVqaZ/1P+sUL24XkJgYt
yBpewlAF0tQYDgPMWjsRs82mrNiLL5jNILonGHJar9Arjcqp4PvsIEv0/Ov7Zl00+oQsBwZPuY6k
gO77SxDSUQpSatNnKWh9c/pOXvikM9PiBSdaS/+AhmgFrvNrPo3WkI0XrQAQKYuDUFDPup2qrU5l
Ig0TBZ/4uuT0UoUCWHc0XHWmGMZlYLbBFay87i2B+B+Eos3gnqf9T+0McweR7+4qcIVUv7dfEd89
j/bgPeBAqJX8lALMjxkP2m042dAB/q/s7kzH7Q5Fwypd20ASRCHqKHYGS85wjVgfnsYV2N1oCq3F
d/QjooSZEhR8e0rvEqCH7fS4PJQhTG/bUZk2b0Qf3IzO681WUcraFEyuq1PrbStWuAIJ/RHumeD6
i6XlVXQ0kAnikqHutwAWQCZtqzFPZLNVhSh5pKrLNSxeTdcpngAe9dnzVxemkShFrkdNcaH6Qp88
drBHwBfoUnpkoXsD7dtDo8BXg9HETzDURju9rv2XbSIWwSkmQT2GNafqeiJ1xR6wxUD7snY6oLca
fMiNVxT4yJmiJ/cxUhwW0myVcsd6u3fENu+2CoKNnrbS6sL00uUohdnweJEMg53oyBnHIuvOCxDU
E7+gujEst6t6pOvfuLmf1e+2ssjPQdngysqQ1BQz1TmBZGHreYJA8253ae6oNGhaoGbSdrmZLfoY
Z/A/ChNjuBQtsl3lAUn2Ee4MpcAHXC5gbbS8s20yJhM3tMgpSQCenAfxxMVTjG+rJA2gHWJmu9l6
Kaa1YSojZEAF59yq3C0AT9LXuqkdbErGUAeFupKnmamCQTufpNHcvjqnlklTEAsl6qn87MzAHerh
tMi8ncBTh9E1JHzRFUXTJk7UtbVaETrzoRXLy7m5P0G119i5jixNu6/F1rLyUbI9vYLKIqXB11RF
XpD5iEyYzTVIXHYLnZV3HeEoQTGTLmp4zK+wI3QGwWDtEH9x8IqoPe0ulMaWT2JbIc2N0D5sdfNL
MszCAO2U6xLzCQfI02zqx3rxRgkxQugCQJktID0I+lxCN0TjLmI876qpM0BCf3Oq4yV+LYQhfdk6
H0Cym4K2Y7pD1Rpuou8A9tCZn3GHPRCFHnNrRKw7dC2zeAbajsvodudNZpxTQ7EDY00LIe8IqcCm
NbHlOMeSW2KgQDRE6CLWTGZnX2qoz/wa5YZFHY8juLfCp46xQJWl5dxa4yt5qm2pYTiCxTteAWAM
FFeIyK5Mc660jjLSc7NtUYXJhHJi0i8dTXc5hV++qOyHxM05653rp61rbG+Ymiwkfs8LuZ5sFD40
HTzhEeHf1CkkR/WE5YgB32VM9PzZkxtyzgPmcJqsAtp6K5ZwEQS7OY9bFekEdv2ZfxL6GvSGISgo
T4Mww8u6bxOnMysWo21xTX4UfV4G2pyj078YM4rgbgT1EKs/1CRHhQaC7Kuk88loj1pIIMKsEwM1
UUBXCd7ylPMGkZ8UXS9HXPEDxW48CBrm0pRGWNtWcYCGU/UnjzaoHrNBJGHl5NXk/5iRkNkYMFHH
Fw/LbXM0GCqVlweX7/5go4lT0y5btK/h8ugHXkR8S5XPrSW36zP5R0K26uySGt0adkJ0gvA4LsFs
KSnyBjZdWkVvSyUWlmTHr15cJ1v8LTAvzsVehnjuuBlSD1RNVdg5ZsYbQSv2fBSRsZsIdWDz9mE4
jfQHSEllXO0A3uWDo3/8D9JjBl3R9kyEeIaD9XYQAXgT88YVBMaBOxfTuP+sGReNO7ZEQgb1/WTs
PMNOhUgXeuELdTg/8oamCLNJr6W/L+cZXW4c9fM3b76DtiinMCrFpSF5Y3ipyljrsi1tZwxZyYJo
Nuh8xOPRex/ItGwxkEPTCUvwvAdBdwcxP1ctK6WYtzUV6KsbaUwyMhT6L4HceLxijm0bhSG8agD7
ClUVqHyV5/UDaOuJJnCWGZutflrGWBJSRciQkqw1LCrbPE1R9rOZMN2hiFSosB4MLpOeVbeLv36L
/1CiYOZCNt4cae12GajX62Eq7pepocsmyn22dJWbNeoCel6rAGPnbuNNFE1XSKu/z5Z3DIf1QC5A
rSNbF0xaycl/WWQswLy6QFQiTpvsqKcncas4GidlMdlPOelbOyDJLZb0QB9sQtZeZdXo3ewGRNJ1
u0IW1516OQ+hGcoDD2rp/yih7cNG3/TK+2j1DerkIKx40NtEv+Gdf9JTlZYyzI7uGuABDlVQqDIk
tB5L6S5CPUkNkV9A3PztHAO4dE+3PJak1cHu3t07X6GnYkOpatxb8/6PCbGt8dRa2au4oXwhHp01
gevATkWPWS+sjPTXSfCY9od8/xpiQhDqerFMFqJTC042DFgMYuIhZuPlq7vFqaqasczzaK7emtYH
FixlLhIpvslRquY7TrXVAMH0EYyVjbCZj7R00aQBLx8cDm+4zbgtBjnxcbKx+R2xOjLwX/YQ7+Ey
rm5FCcZfQa44gnl1lgJ58HjB1YFRvI3zDeCSbd79Hb2vnPZxsgCXuO7SgsoLlklZtsL0+ZzTsLzQ
CH760bsIkZv1OIVuAzjq7nydcdNBq+Y2hJXZ2PZmKlr7XXVnaXPqVtmb//pTN1FV6BiBrf6fqjhW
HzuHClY/1iE+gbB0xQplPOqiBuyFS5hEdBt84WpNxEdQPvNJKH/MRUz6IbHGb4IW0uTvu8a3JtuC
M9a8GpjmVhVPZ8qLv3KYNtCByVis0LKwh3AFwAHOHSCo7sx6C2I/TXf745Rqd5p2KiLNjL69ggQQ
rw1kKqsNXUB+cj7UkPDBGxjTB2zEgFk+qvA4C5HWxs9Foxf35RtuWTDq+aUfVgUPWgLvwAN8CRJx
+30IMKMqG8m/aXqCWo9lVPTHkxxHsUss7Qvx+3hTYiYaYPN28RyAj/1ojzRAyPJfeq5jVN/p8app
mnEJTdQiXk2bnE+unB0vBLM6qMa9C7jkg5+TnuMi4W6+oN9QcwNIQ9BfFEeYl+XxII1HGvXwfTeo
uI+fZzBv8oT8wy00sZpM4bTzGdsxCLa4kGw2/X07W91QZg0CqCHS7/XZ3uZzoQ+exh4xzHBGZG50
57wd9Vif3osI83KbqdDPHtoxg95dY+Z6/jppM2SO4aYlFTqmG7fJimuH/c1roVTOsrmYpO8TWkQ5
woC9lHo5KA4fpZXFhEq+FTIO6f0rMHIszJlh6CmnDdTN9XRrXpuQcIpEvqAK9bRuyXmrabcR9Q/j
Vmyc71YIaQgcYjcQtCJRVlnAXXma1bkhW+IFdjsW07oy4LSUU4kdVPIHBT+VjlAAt4wAB7nSEy/5
xZrWvusQFJGR/XiZ70RvOA5GyY5YOaFyREns6nAXo3cN9FNRtLAkmvPrMXMwscPtnKKu0Sd35GoM
eJCom2n2zjV4q24SA77/AVqdDJs0IfQ16mEnBAd9NqR2YSXAmXzS9Um+xOqvMW4JHNuR0y2uZXMc
y5xg1zrCDdphzgtL9rFxrRX7EQjAbRZ4Z1QxTafmfEjB5IeCwrNn++Km9fhY9PO9Iwzuj8lkjnjo
FCuFrvIiSpdYMCWxsYbMA4rJ/bEK6oCg+3EPXehHa8SFYJY/cRX4YVraW8/Ab99iJYFgg1OZ6Q3f
68RvNzfVjI1Q23mkN4xGVtQzSxRx3tDyrpU2q5YWoYH1dEBPchIoth10xEq1UXbxMjFuFnR1yvlO
dKBLhcgoLlYm6NHh0/dwyisLyaRlFbJHuumeSFIJnLQPgWFzpL6l6CwW7wzCYjIHnggJPtPYBFbv
tjG59BkRYtX4LGPIfPkGd1pjK5wO/OukzZx+vwKUAp1kJbSTToZddOZoZ+wm+uU710V5z3AGd/CC
R4KnLFXC6M1gEfpEgyAvbK9KiChnkJ7snmub16w5ghKVJPyleEJdhVPsfDHakDebXQXaNNWlxa38
tnb5Lsm0lGOMqm0jJ7zggf9MglI/N5NbhFT6ddTbiML71BZJ9C300W4DVv90xey9rvZ9HtQZajDI
TDwiUJZTzkmptxL0g5R63CrxNc1mi4sG3BYjSPIryu3r6Qi4nmStWHfM/zxcskL6IdkeurjWk4oT
DxdhNt/Y+9pbSM1YMVPBF1AN3X6ML4xRTmkz+zIeN5foy8o/c698gpoXbZGDGCO274RjdXNBxnHk
2B3u2zHfzIXOIiK4Zoq25E3SUshgLhBd86vOIit1ywamoq29Rw0uMcVCz2U066GuoZgHVIjD59SJ
pD+/oZpN4vet1hdkZhTdzrjijHLv+vC0XfK+iuGhdefRqZqKwrNceEzn6eLVZPc2yPPs4uEQHAfw
DItZAL8F/YggbNwTGbJ+YmrZDs5KG7DdS1TZhXgtzsE1ynpJ2aA7ok7rVziMBvK0xF/GQpHL9RTc
zbUXbeoQRwL2pZZvQLkukt9wnUAc8AU5CZ6sjb2BUtd08nnAy1uE1hVO6lC8MuJqXevxQvAkCeQv
+Qo4ISZDNJaVLB3yW/J7AsZJe71z+64Ul3m2a+ykxljPgf8Hivh7wMfbNBfaF8LnRvsHi4SDKZmr
bXV+hkCs1o5WeW8dY0/JDCb5sewDO4Dj6KNMAKBU0126sjzZ0HFwmBQrn2K9VE935AgBwFgQiyCG
CuxEiXG/AuQyJdJoB1NC56MHMZgOdT162evAlevC/uDyZX/V2tfJr7e7FYOCun39QK/jfbDvT34c
zjS9iRXwoqu+QRyPmGJUXt6xFP5vHA4B1va+lo7nATPgJyB0DVzKHryPL42KU00hSUTStRBU+3Nl
kxr4w/uZF19XTp1lPJ1T067JPSO958qRLXokCb9cEOhJ28uv/PRhmGFqj3xCeQ7uuhsjTe0KojW+
WUPcOih0CmuBQHA/pW+0WQJmHIaFntK0uh06AqlJS2T/9oJL9dyMLztJxMI9vJb9WfACu+0Ispbu
R9zTp+AZZt2gOvnWrVff/6OmW+u/FE+/NcieBlGoe7BOo36ggT262BO5VSKyB+4/Y2fEdrFXdgdi
9j4egscyVEoeseEn7E+W6nQmXoUEa2x//8NJMUzpQ3HBR7pAJp6s7qiD4rAmp7lpDJ8CylGr5mUk
lCdPtW1QAOHP/E/bANruBBxti7DSkBNvPUlXaEubiUX1qArnYTRDZX+dOF7u5dOWTuDG3mDHEUs1
KpSddQDMLdOsR2/wI4nujFOzJ4GK8Tv18gz3TOBGO/n94eXwmd3O7pVqs1yvOEs3UKZxvXXCoTo9
KsD5dzEwSiAsixOBmm+4zGjJhq4rfXU94di5dspQkZ3CGPwhNPh6w+KF1C36NLCUhjM6EvrMaAxg
PVuC6H9cda9q4k6Vw/wEqi7N76JcKNrdvv+/kCGvP8JabJ0ckazxZuvdwrFisAi6XfSBK9weRS2/
9QobC72WDIYsp0jZ6lcBSbHC3Y9c/GvTG0WMC7144JsmFKu6Z5ITSUeEbab4YxZhGM7uX1M17ZQ3
pu3zEqNAgmy/YzGGIpd1ovH9ZhrsiHHNvB8ZyPjZ86dlyy0trwu7UiajuUK7xAQn+h1215CFph1o
75XHl4ElySvEc+Le/SRoZKGpDRV9idunULGYjU+3JmbbWSp9ANQnQBwf4MMUEn94UMSGoujxMiUI
Znw3gg5iVOLtCuY3wq5r01A+ReE7JOoF9a1bLaNASSEXfpztBQIXqywn8EkvXkezlhdMaD+u9r4h
MbllQrutbGcMe1Df5LcnF4XryJBIlYAVRDCR3+hrDCawCHPkGSqqscf+ffqQA+44ee3G7H1PRRmw
p4nedPAodLzg/YAdocT97PNreocTmw1bIcRJ/3lNTt3GlLWOwoJu2/31oj2NJZL+Dou6FD1mOnv5
Qt137s4AFnjx6NQNQ+s+Mu/VOuqRQZcb9j2rQCCZEwP1V8RGzAdsP7asVITyskriSWWvkztQhbd0
5/YjiInYLXwXy0dd1ksDkPlMSaaZOBfHI+AVfCJGz5thuX+2SNXOUXX8NBh4QFpoeSKmxqG0UVEk
+4poLNfaAqnr3BgMvhsKZ9Pkq189uZbM8SxYeEQ3vfseLA3AiQMnTki4fwksLHuBD+NgIKrSK+X2
G/MigYKyXIdWWRzijEpY6+z7BvB3Akt7x1abVYK9kvGZHBQ537DMNSJMZyLQ9rm7lfYl1ScaYVep
8v8twYmjKL/tGfjRN1Tbg+xo+R3u9BaagSAeEYGFLclaFQqkmm5+3aLQQoCbTe/HWlrcciP5ULx7
LKd/BYIgPivny5fMKMiWIs3luMA2Nvv5Rh4A6wkCMNDyFy6XFYbq6DJ+v1gRrENALVx8s8nzwLb7
BUlx/tPbDq0GV4pg4Q1w6tQR0pRZTWDgEyBGvKBP8hjXN1LwIA1G5Rbdd/537YeVqdZ1Hu4379Jg
13p3cy3BsItPLhJt9P+rxX0wIC9gRNmHjp3ygrAdaThgC4gJEsoVy/IaEMN050v3JNk3K5gwWoxE
6hd0f3k7EdKZRjrUCli90chggQ5gqsloPCHUOvrDE7koxFXN6CxW0O5RlgEcmoDpIRtaIgcAEhkc
1nb8EY/pFnqRpZBGzgOUmTRuNrVcBObQjtJRuRwGM9BXAedctThuDptDx8D/M8dDonguCQfa6HtL
9ATc3GKe/40pMDIow19DO+agEV6TkkUPUieKQwQ3NWPPUoOlum1pW5hGKQio/qM/0HY+0WbqAWci
zHRwR+nupeHEny3rvEl+jCHePF3XquXRcgsu/paEnzXjHlnTwDFCR9z3R+MhUYOxTydo6sOBzcET
jy8WTc4yNIJZ2ZH8jnRoTF61FLvMvKGv9DxtHqaRtRHdJmIstKwQGjb2ZFcch3z1ILJBi9yYszu0
GfLu3AODVF3frUs+rEyBHWT19SFAXTRjCEC6Cndl4r/TT7hmfLrC6b99GkLc/KX0BZy9xnV39NxM
7cbRAy61Hy4QBj3roxyOcS5ujhhLNDPKdN/dcl5vY5vLjyQzrEcChZhVrl4VNn5gMH4QaNzPc/wd
Hdjz1AJ/wx/4Ou5P+KuEb/Od2ehv1ieFvWobyWgks68Jk2KSleI1id0TYucqwdyRQ8h/QTOHr3jb
IJNagTjvKdg0XG9dhd9J+/2RMgO+Oi6jctxKa/uZR/pUBm1CcDSb7xXOAYAupMDxmTWnXbzUA6uV
EBbX+2QqTCiPhYb4naDRDrDFxtDOIbZAFNe5bCR+XgyEXgdcVFdHnJwzO2LqGoVy7L+PZPg15jTF
xWNnt6oVHaBaOzgsNkG7C6Z1Mq9Q6793suztDidXS4m/w5+ym8mf6DPy54mVzPTwSF3zhUeO+xMs
+qBMLKUn2OR0OQIPGTTxqpwHhKi3xthQKR1FEBFqnvSPSxgFZwvrT8mBYKl+Yeak+L+j32cz/rJS
SMSzE9meJWoU1BjZvBYPu2CQqmqOElEvUyVAtsutszN3xBSY4vkdxkVM1+239j1IjrxANc9d3ifj
dqdltqR7zipP5u4WSHQkI/F8kXdUCTsAs11IljCxGM++vgFxgmh3lYH++IaPeowxPoKqodNAuxJk
/9xFZF0ncbbt5kfKlT4WR4KIlBgnGce57WnInUx0L+c6PRbD+2BkoFfAn/n0XlVrZk/J37nmUUMb
md+NHBl6ycemPnjA8o4uA/mqsZ6wq4H5oVOmIr9tmKIF//SqEiIVUichVQp24WrVGnuWvZmH9ROk
yZHe8F2RCFLXRs1VN8OFsmYU4pHh1nMJMIS47ntGQb30A5iLEzZaO4bPfjf8V9JT0ASEeKo3T+It
eZqGzxIVok20f0RL9gNUsNKZsJ3jL45bxX0yigBK0H8Vf0iC6KP+l2en9Voa/01Bp/enfjEDPzRV
VoY0iAEo/JyEqim9LxhNuw1O66F7DORlWwQOIIjVA+3OodmyYOreZzjzd+UaPciDZR3X2C3+IZ0E
WmeSm0XGvxnv0vqHLr7r5MLzdR5Bb1qLYx5jxcO907mll6T4Pn3zDUqHLiWvfDKAhWvxDr5m0WL7
WCpEK+oq6uPAlAv7OWpBNZm/k4Cib9wN4bL26J2gtLzP3uHNlPZq92+Y874G/DW7br4yxRLmLB8v
fi2gcT+tgaEDBlEMTZaQKEmP8luSBXQt8UvwkRb5iM2LtYBt8qZuidplX/tfzYlFLKxSH26umvQu
yJOLuTtDh28QKqpG4oRRIgeTlMNqHolYXuuci8bbt8IGJQ3trxMEf7btJMTMkbbg1iieNpFi6BDH
3bKutVsxs+lPc7/Qb/0spEwgU/LyGbB+kiau1aR9pz4EF2nfHhNZ4xYpszq25ON3sWkTVBGlefF5
83BnT2CTOWfoo4D/g1g1bV8pC1FHVu1wTe1KN4SjqxWbj8Q3L9IxST1sWeqcrYHuaAZfx/YZ3m5z
znI5yXcNpN18C7EvOC+FeuiWs9RQwM3Gf0KJVsBTelilXUjFquHRht1xgFIiyB0C46HzBCeWOlLX
dlSOUJ8FPSiM3AEqvUWkGw6ixHFrZNwtOSSPEmgvvXA8Rp574XckZmlPyTgnejFyNqTa1aaNpmBF
YGFw3K0zUCOHJ+8VsYjMxEGlmJowRtfEniljNhBVBNHntnT4Q4lPEFfsPhyGPkzdad3VRJP1KetY
cjxzgaO9t45+49627Ltm3D7wCBWq5JS2hjv9q9Z0DjPGHeXUNWuEizOQ7GJtl5czApJT6j10gCEb
vtIqtkyv9lFgNOFQdk0u9ZbZAnezPA/hy5IH4FszN+e851HBlGFr20iUrltJeXP28pu8y/bWX5fQ
B5mpM0FFtCURnvO2Bn2OfqDoljBNmttqzWNNRyZ5ljG6JhuH027yD/KNJI/r+scQM9+kIXKk8y+5
/XfqHFnBciSdBToO0EDeVN71QB/oFwLY0QqDDAsD1Aw9FJmTeOECPe7U6JjbQWJsNuT3xkb2YdHQ
6ylSzPwNxrGWVn/pHrpJYCirIFIahjZFaV4Qn8aMN7p1Xil8hEV5zLSGH2Eq5BNu7XlYdse73JMA
TXgYEe1AnVhAw5rSTtHX0MdI/A6wJpnkBg9qTbsOeik17fNoiU1kfuka8WAWhWJb4sPbnz6oPLaK
CCSBCRf8P1hkP0piH+FAtUzlwzXsTuZAo8YFJ89DT4B3Cqhk3aQ8feb4AMoMyXxHDaojb+oMI2H6
C4C3SaXYec+mtMjOiXJSXT38SV8LskB87QMlgVb3S7hd8CDht9pUZsLidjtD+ARNQ1JTNN9i4ALl
rWFJT01QslyjugWoUNIaiQNAEY5WmCgRygj3HL6lhSho25iZ9RZeZ3nbAxSkxFlZAgTGsFL6k7Gi
DKGuCb5oJusmmbu441a8uIRyNu1ga2rjvbhnOhVLuLrvE9rjHRZgDW6DkijKG97Zk2ts4wg+8qM0
/wfKMNV6T+JoDuTkaTOXxYrTkT3tYWSDxYlcdrpJXvKTMH/QlZ7iwzzk9XZfvphtsllAoTdAzHpQ
vGfyIXK8tpRc4pnzQKVZNk+LxOd9pvNzquoPUfj92rBQf60UTe7YMCwTKs8Dzw0JdyGGzMhs6N/0
smf1SakLRapUXtqNKrZptzCwVhdxscdu1O5HeQP5rdZinBgq+vkG/xEZADfUk7uQIQl3Ymycw8yj
dEYU5Kpxw1Se7jXHBgi44dAr3an89Ua9WWpvOvGRQePfgNU7cf6H/qw686juGl5QzOigB6KrGIak
SrcORW2oYmLsuzSaGJLH5SoZQdYMezBPDfpvhqPwBHkd7ueWphTU8XYSsydFtA4WdhJGk4a6Bgz3
szFkg4Ewade89D3fLcmAc/2ywPY8Aun2nlhLh6gMfPnsHGKwnanutC2T2sMqHJiEW3IR5TAjb9TL
VtomLlFl66rciXaXb23sv3t6LT3oJvczXhmsqhbN1rIMePFd8oZOAHDzgPRjvATgV6nmRi3GRQNA
cWpZxyzlUrepsCFBUmO82tm+IjkzsatUpjeQCeaxP/JQEMGk6wyHj8RnuReC4gc98mKy+mTqj2ha
jIA0lTX2EShtjYnOVQJkl8/xgpknx25hR7zl4PeEaHNTWS8IPCvsp0+SLDgkS8ihnyOPfEI0wwfz
mUPxvo2dlc6zhxB7UDSdynQxVutwxFejOJ8JQa4GAyyQSMZ9tN1XU7pYk+1BDL4BoCSHCDIDQ4lK
oLWgsU7Rq7BPrc0LXoDDCMMs33ocPfXpZB1f2QUCARRTtZEco0vv9/1Oy6ZHEAdAt7Tfw1IPi/8t
0NgfY8aLQY0VLUk0ls+P+5lXZOO9h51gq7hKuUeq1mbsvP0hl5Iftol6quV1qNC7+l0qqyHxl4iQ
QeJG1KWJS3h3lzAQ6TQ3n7pViHQN9FFCkfPpq4g5geyBU3b23LMQQD+bZKRkKAoDxA671fMYtvGI
E0p6fROjzgLRv8139N0o9FMueieTA+b6A6YLSHk//6eSl1dWIvwGSt+6a4g+5TiULCKwO4w1gq9z
8oY0u3GTNPv+M+Uj/+0+N2noKDdJHuaSOc+ksT3PT47MuHoIEikDoSwLePWfNWLgB4pGj+nN14cF
VE8+KNVDEwdkLLqW/62M52dP+s5LlqnNF7fDqQ6Jsg8rNF0AdmlCsWugJMcwJP9uLuMS5FOs9FFK
1msQ7nwJGXUogBb8Qj2/pBiKdvaQI1MlNYz/pukxC5C9BPT+fBewtC+fRiaFS5nYV0Ou9sF1M1kU
5mnfn/uudZ7rHUe8HuU1tgoMVuVnkK1DprtjHvFYq3LfdxucGqv3cni5HmG3t8ie/SCdY/QoROFP
BjFivjcyOalTdb6gSzie8gS+/4PbA59du29BJ+lLlh17CtTqAd+vYf2IIy+ZkC67XsisbtlML5EL
3Pe0zKm6J5ubvzJUhgjrqmCr2txblJoghA6gawQhdwuBc/m6F0mXAOO7vzoxHU1g0WfdluV0Jyoy
frE8fMV+solk9csTqEnniy0sanWyGWTsbT2zgw1maOl5YZOjionyFIr5TZB56RpPRabXS4CZ0i+o
TyvYApn3o4PU5g9aabGJ6Sb56dFsnavPx1LC+ZKW/Zp/wT1lqkqp0R/yWCscy1+ZYns1F8NVNZco
CZykgGMkUK4RbPkKOUMWFMSiioNkSdPBCdjTpyEli1mdJj8eVwAKRkvijwgiH/DnH7k+wEMLZ7Er
acG7tLE3hFsCsscguabUXODHawYbq3ijN0mJBeN3YLq3Ow6kj0y9woK8jJ5mRpr/fC+e7vMJJols
T9pqFnY4UY90pHM2oK8pHEXkcOepkkuY6SSd7xKVi9t8yhWvYglTflJh/4sIFCKW44dNi+5o/PJz
7pWVz0RNzgn5vaFW0cmJFB5/ZcYMI0+yOHm7fiSP7VFsdPMG+JH3dOi+PqweF0dG8NGBAWWOnSH9
sKU4MWRQRUGRqDPHuK0v9T1K0Y8QpFOamI5hILjLRXd7LqVF7OS0NmYl2JwtSmqNYQXt+jFvOzvF
0LlcGZFju0wyDpUY6sUFD9JpvsREgaiHrxmfBqr/KM0rt68qE2LBQrUuUnjkK+CCmIhyPnJqBvjR
DoOic+T4CKBZ4N9nY2aaCf0Q4O8HQBAEqE7aED/hQ9cyoW/Rj4uhorv7CyGh/wkrwRSZJ5qQHrQO
7oKaWxzuKnQOL/HXPePfwEPdOQ3sGRD4se6oMQ/VmNd8BtTmodELitRQkaAuRKE4tyFDGIBpw82t
KtNi6SEumflbNBd5KNuJZ/cbTqwsZCNh1XemTL7RVNhfaiNT1PUGozQDL5xm83JgTiPHfgucOfbz
WO9ECnX+KcRkaISSAlGHTHn3wTT2Ll/QsU3vddLyU0wZA10lCzZoy8Bw6JQXcMMoVrFEmy70ys0k
WunwHPAZZbpAqeoF4uzECNK4h4PQSIrFEflI3dYA1lJ/nrNgAQlICHRDri7GTbT4i7JLFVPKIan1
DLhkO5f0zsJB7fWihF34es8PpAN/uQk2D6XHvtsugpkmpBALiNwBEL6TOLAViUrV3DfUTBKtvFh3
Q69+Gei6vyeHSNH7/g6pXxRBOjALoRUpEQUAsuBpuK1+R6BKul+q+kCID/tLeI7jmhrN3DxfKpbv
LA3pzLj7rxiTC/99eUY+zU65vVfxZoRxLsGlQ1ktmo4wS0Iq1t+rCG7joefqLsSy4Q9HtA5SWMjz
aJe3pUgK+QxJJ1/3Am1aY3a4O4AUEO+qtUu1lwmBEDmM46aN9CEwkaYBnVjqxxFXpiokl4o3WXGa
Hd9ILklpWXiP/zI6XvPxBHPTZV5OmPOZssyeaaenglHOCpA6cu7+2JEKoCnJgf0AeRHCuc5/gzV7
N1yUSHkJlGZF6CUZSwyuKHNW9ZPCtn8F0s64tb1O376OT+kd8KPmf2mXTp9wWG+yaqczzalIaJDc
uTI6nQP1yf8wkHGwZpAzj0McRvuyhkk2So7JbLcsxwqLTelAGoo+OwJJN3bIIQ9dJVClweHpgoRD
5JpX5R61YjBJRtpGea4wu0J/FpOzxhBIhlLFuQ7HqHSzwJd3DDhHjspoOLn23tGdFj5eaoY7FRYn
/72M6MioHRFdJNcawmj1z8ovS92PpyZqpWjk1njKph+/ZqddrxrAxEcuyb3d7+t7kaFAqrDcsz5g
HLsfLcCMzuNWXvefKmJAhUDejUSK1nycbN4PmwtN8wWMN45Z/Hz2Pg+DoyRIZfJFH5yWqEV348RA
7csXeATIPjThmydiHum0OFRCe7dE5C8hufRuyzC8tv8OpdQSP0OcyaccXKkHLaG9vg4bBlQ0U1S+
A34mBx6LViaISvW1x5yCGbH7BDxqUJZ6omFaN+W+LFbnPSvB2so0/Im12sVFGxvdPRj51xyqaTi5
/Opi954leLRRY/O9hTeZ5AV1RCo/vvbIxS3l7iLgvwvjUbwhPYoYmWh0GqFQEbaoYsE5ofkvQO7g
aVQ4mUw483zSXgBG5MlEgpjulP4csq3nYW6+s8j9uCF48bgJsIa+S1foptnH0mgKPWaZih9zTnIE
RMiwwwoiaKvmHD7u+m8X31syneGNDhKHE2Jh8S9lK1jAY3/08CsOeTSyi2UrWjbN9Yq3IIUOuukM
PHWEaett797Z+dLouzuCwGvIgIlY5IPfUTQRHlOtY/0KE+mSzg7FsVKVO7b/8yVa5xZhFbCFqxOE
k3vG0Do748IWQets7cJt4XYFpmc6CIZcIg/+sKGHfjAyMaVqTNQsEzC3nNC3ihhRF4cXra86Oc2P
fd9ovyUEbMk+FgrHcAOqnhl6AcPr8/Q1r3HUiK5wPu6k+sbpDDFkQcZ0jVvmLHr/zw8J7Fggu7Su
S9UpdzfJ95RUtdjHL49LBi8hYV/U2IgRavdbmquNJETGRyHIb/+bAOWDMJMPS24JBcbZ77HZmMtx
oy0QcXsGw30xDtWCzsEezs8A7tMgrOecC49qJBns1EMdgS22lz9mQ5w/TdETTw/L+zO4BKcMSLcW
3aqq061OwQMY6wjytdB0quUeX6rWc6dffEJCZ7ZOjroiA7g8gpZHuds7mWOLHI4+uvvgQ4woaUW3
AN9UN5n8SyZ3ox+2wu/UkUlXrIwa+PQl7xpHlR3Hu9Sb7SuyEHfDb21d7lPkiejUad4+gW46RTdY
5EALCZPoqzEuv8NUcJvA7F9el6+Kd9xQNLV6vot9tBL1r+cRfDrZnJh2MO2cFQWlw6FybYEZy4l0
MejlIqkNVSiCtwG+dG/pyAemENNh8d20G1PsSfKOjLjnT5guCKq513c9iUJbv/VEkakFvq1vHdtH
si+h1wMPelABZwXrtikBmSMjaylBR4u9MAzpBjtxXtW87zQgEoHBQpNpgQspW0pzw2uAy/BWreiF
xqktu5hs06GZ7UHKqEKK6EZC7+Uowk+/rT5Y2mPaAtEV6RhHQ3oiglcjiBG0GRz1R9VNmGK2uvoL
tVfFHXOP7ofjIsXVy6t28Ox289rbb2Rdd5SPD9reysX84KPi5KUPOAOroKOHS8FNdaGB+ZhHQaXb
JUvNDMz1wx40rb4j+4axxK67J1RZkIOyztQoIuxWg0wVjaRKIxVndrWhOk4iV4K48bdxDiBVzpUy
EExgr1ERIi0j0RRBLDI+O5Y1q6b2qFqgUV/1Rh98k7YlEAbRwY/txfcUrn2cIEQJUwHyrP7ZrxZI
ld2xuRxOjrTb9aE6Wgm92Ruco86N9SA/NnuewCp9hKnoZsoLW7LS2l2+e3seTTmUQnaHiabyGYoY
ALOMmgp/l/ICFyrSKdiiIMAT7ME7oi3/WysdrXCfF2vEZNSDzGkLrvZTEPluXx5Zj6zB8cgdO6ES
zQVaSBxJS1y92tWFJNmIdVcgMfwqYxwL+pQO5Q/oqHnIZItAwYXCPHadk9rMKstryeVxDysijqaO
0W4yix+mcZbMvgUjWlBcxk9BQ3/RXVqM8MBYoiKqAfj8RIG36SSsTTpZwgvdVUnVXFmQvKNMTQL6
xyYMegx9n1K0Hf1KidezG/uwX8aVQ0jKrbu/YSZIpS3/FHdosOfmJqqV/XG5g05lxE0ZgVInnDXE
oI3UAYy6e2JOtBu4u5c8F1G8+Kh1nXFA11Xm8qOA4XGoO30MmGsvh6TgavA8mdGTb+1+VYLj5IJ6
cZIu1P7FYQPWWbNB4mACpZeUXSPrhSUfOS4jbYE1Pi1lvQol56FvPlJCvipa/Y0N014cB32ofQ2X
XPiHMxe2OC9uscnsUM7IVjreW0zBF7nk1lHyXRYMEu2DofhCf00/Q9D5Jmo8ZzbYe1Sbf/9Er/I1
op0NR1UE/1rTupHo3BbiWI2kaUfnGDRWC89FoEVUPxbDdd6p9viFaMBACXHO2k2v32mVldDWY1n0
6TWwuikv8yNvotv2cey0iWKQy3a4WPpAfdY3Ii55z6tG4cHcceCVNqSKzuN96WEw4zXqhZoV//VB
42w4TgOhHl/U20dtkBZpq7h5eUVkIquOvAMSXXD+vEanCB9pfIsPNsIFelrf3P/Zaspoun88Ph8p
vy2zern2fVIapUIWruNovgx7a/7sqlLOhi5IZXZR9B9d6+E6pkcj3LomKbEC1yAUgZqcE4wWz7PG
Dr2/onLXIFheLQv3LccealALx6FaIvATR9UnVI8m6ucZ0vLb+oNOlHEgEVtWVeXbKq4fFl93366H
A3MbjMNUIIiDNGTkWDy/T6ThGqjm1pFUQRu6J9CEr4IWNmBq33MiKSAvd/U5KnhQvJMjVzFCOcH/
gCXkjsCyC7XKrJizDoiIyg1puFeqcQEUUYf5V2GF9P6slE09UuNp92c/1qeAk4C+EiQkjIjimanT
SmxsQ/QeTZ90mCRNg85ZrE9Fzpee17wrnNsp45+wsEz3z0hxDyd5y8WLG+hB6b4LFxEaTjRgrbtC
J0afl/cFQiOsn6DRttw59WsPud7jo9qmR1KLScxC1c47qA9xbeO6jhFHX+ve9ssM1E1NaD1Wti71
lohpKQ5Q4k/AyP0+blCHkJzEDmpH6UhTD4d6MYd49RcZhyGTxfSnz8PNNbPy3B7q+BD3CCGqgO3j
0LSszNGyi0j8RAxNRts78wbL/diOQWgr/lPNojaO3X4+qypTCd+Y59r8JJU3Aludz0DbwFKwIwM6
aF8+VDHAKJ/rdaQqkjlxP5zj2ssL/NK4WFl65qQFWtmyQCs66+vBK31ruK3Tm6r6mMgtxQJSNmv7
Fw3/JkDENRpMM3FjXFLHaqoA8p0sHqhp3z/5Fz/WIwYCmGA/N8ezku69Yk4PqGVxTvn+AMMr5tII
n45dR1lOS6GkMepMegdgDyJZFIqNo2vrX8SAfbQWTqCiNTpRwGPxYtzbfPRc2E68qTEg6spUPwvW
F7ZAaWFViiY8NmavyRJ3v6XLZUjkObpVBkXmE+CestEqqc7hjLfQxJiWn884IuvDm7KP679hFBU2
TZk+1iv2iWa7JYHd2mRFpbytkSc4vpCaAZMBcGUb7OYzQwEYz77gZ2A5GL8HQcjcvf/Im0fnKfyE
zQMfbHHjxE7qRHHYd+b29aq8AvQiT/rCM4kiWGe8O5WZqaJNm5co50FNxLmJoG4X6NbWU1ZHJB0r
tXrzx1W5zMgnFFYHLSH+ANiNINXr1BtXpAhKboaXQzXjoez7Gg/LhIgAL71XcwNgdoGjMehPDl7B
bHEy7j9owVSS1rJMtiedIvrEOGNtwPYyRWLrXCrOBqBcFWekOw93YYdWQwHYffZ8aXKzzUCThRuq
5YfQUNMYt33NsEn4jyP/+CGFBR5qWbtp3fwnoECgAU1/SUWYUCAIRgTLiKOiHowu4ndmFSetfpsU
wmOGeZb4a7oGUitrwXkp7sXCU7d7sOaODvI/pKqR9a06qRcAK9Cb+YcXWCkDRa7en0/ZWB3KqOv+
sLd5MBzbOJgxOREXxZRCFG9MXdrlbnxUecBudiWer0uABxdgzi0B0XOlAtv0zp5rpD3fvxKc6LJ7
SSKjpyVrWjX6duQ7agpk+ThphrcaMkp2dJPWWjARix2v6Ts462dKSCbX4LpsW9S5gazoHTAaXBIs
1OJm2nXt/7sXE8z4i0D4uXYRqV55RpC6llRNt8QSfkGnRA75y0wkNSdSwEqxFiMgA6CHbmcA37tA
9U0Qfq03GINOYx2dP7LnrcTpRl/0G3uMyi3eG95v2cKB2Lr6Z1MmxSbijE+Kqm6F5NIe3HpRhEY5
xjG/ovwAGmZ2cLllz7QQq9NM6XSPj2t8W6ybBVGl6ivdZmT7PIsOIWJzhC7LfKf4nyh+HDnaC09R
KpdQ6Y8oIIURA81jSp0lbmSNo/MZAwCOkksTBQLUiyvtR7cLYf8NmCYSaL0Qoio/EpIBZwzLKI2+
95CIkKKUV87/quL0l4YZoR33hZQF+Gm1Elw0MOQz+PwG0bIvJ9WPmKSeTXEgWU8+7D9XHq/0JIEc
U/rb26a3RS3GI3G17sFS0frdigX4Nf62qTK64tScq9D8QJfuR7iaWMvAHdwzOmxgEI8Zt1MNDG6f
6Hd+uukjYeYG91w/+NRW2GwEQva90RuIcJaxG7ZBh3nfGdiboEouAIlBRKZ3MJlJpVV54E1l+LPd
KqYOK1BxQIMAbPbgoimoC1JtzhXaKSJQBaVlySSHPNUCjJhQJN70uyGG4Vz9peli2dFk76GZphab
oLg3epZOqj6zv2MFFFBIXgriAHIf71hXCsch498aanHAtwLK4Q8WN/d3rRhmz//SiRTL4uwGNydE
rslPojmneQXHwtiuOjsBGqgO0R7V3PVpVIrVkAofl1qhIK4osSlK3mvTvAH/N8kj7ZFq5umiw7+F
Mzocirns2W7h1U0hCMl1Vu78R+QWz65IHdqkKggKXdd24fkl8QcUPe3TwDxOGs4sMQ5ErGm7CWvj
G8VhAg5Mr3Jeo8p9isrh+wDduxh37jNW+GSXNe8adiVuxlDyDABIICUPfwPJQZR9toGy3IBUzHtt
5+3zMkLWzvZHUYulDaKQWuPiL7nxbzQopTK+oC5XBVKNgByOkJE9uB0qHF1qGF7zcql55uZe/qua
f+DvDtd3GSXML80wgyia5GcUK+0seR/Z29klRchAXLv5TPOgXpdeHTHU5BrjfiSwJgyiUfI5y8lF
iGiB6xbUwLBzWQbjSn6FojMNoISL5ehFDE+12LjNM0V+TrTyWW+iSLdrp9cPYzo8yuXS7jmiTedS
yOaz+8AXwACJnLIvqr5XZnpFpTc5Zf93JWRw1QDKFLT1IZT75r2XqLxQraAQaDVJsRImtHUxAbpI
cTUI5r5BMWbmwhCXev61c2I+2AMM/v5r3p2h6zK1bgy6Eu0GryAjWz/ylSRksETOtQ7NodwCsksx
g6LRJnLnPERcOSaZEEfDkt7E2R0emYgOQhIjAPmL/9z4QdxGY51BAiCqnV2vWeu6Nl3QWhQAqszH
QYl3Y8T+CXW0hVzJzyTSuPo5TlX6frLeplDWnDPgz+N2U+H+4goi0LwZzrjAnHYsp1DJZ1BJvVNO
mrGa9wfdwEG4vHv0gob7mzHB9KUYb0WpKAvp1hZvvAAwLGuQ75yK3OmEYqhi+aNppEVAp6ekje2m
emBN+U8qj01CG+X6k74mELO4kIV8KKzt3RlnN2GY+/QYOD9SqOp0PhHpqaITuVDJmtQICUsJ4GRn
nl55fopFEudPxTpt6OF6WOwApcoIFVY2vSDso3GuA4OmBCp66Y2RUHMFGSFVnCJT+/VammlIS78x
hFmOfjrDyVKwiUPyvDuM0HNivehY4gC0fHnPp5Ci1Bh9R8zMQBN14gPOMKD395j7mPgCdSUkU6PN
gaDWVpjSn/jfOusafG1GYxabxP1FlNJjX4qMOgHDc+EP7ex6SPA4zEmSHRIFGwXcZBjHBJNUVX5i
0BONxiNoJ5RC6Qxc6z+RF1flkXKD4gIqs1ZPYojy6Ai70xS8KaawBuTkG+407ie9+MO4ZXRQ6VXE
Nup3PdImpNuIqymhDdbLKLsghnVyjI4phv0kDie0dgo2a5eWIUS4JTJ17jPelS5pNsGJlaCAHzv4
IW4G/nned7W5u80kSL1qF9SRUbRy4Bw76k19epifATTLoq2+xLWzIk4F+e9oUBC40Mn8wqsfiQ0G
x7bT8txxxfPqAznFtMV7rOafJ3oEWJi8PWCt6/fkelBaQqoXP+1PbvXIgOk1pGE3ptm3uJXyw1bW
0FGEMBn0kLFUhI0+nLS2iEICAu8FCQNlbe3tUEyoCp47Lr59qq6tuHcMITaEDPNUQpjgqr+UAj03
76Y2om0FVCuxiSEsl6DsIGrrKH5OqMGQ5mU7QVYBOqs92bh1P5wHRHNAsEisYpxSRgjRmnmBXj5z
rzYBLz8Mv8PfYZAoimRY80lWSQQHA6oQCvMRPDSVfVssTcYSnDUKOO3MPAyvooO0J/1unLkwAQAX
QKQD3kW4Tni6H4Vi9ON3leBo9CzfTb7Y06vy9CGDWFgZKCkTxSVfvlCnu1HkmNhSC87+EmDY3TAW
4l6VZ5vToHD4U6w+lS2VpLeW5QoYX7ZGI3gDZUMhwS5i5y6a8LEpwBIn3mtxOpDo9++tuOkn0ZGS
Xx2t13+g8CP0/UEDA4ZuMFD0m/vOsUe6NlieslLIRCgxKsiprY+ZgNn+dpKtUHn6V5O6CAlX3QYI
O0a6YBBM0+jpwKhqCxAhgjc48bXPc+x86DA2K8214LmOGdGS+RG4MLhxPuxeZ3ij7xy+5TjGT+EC
n75ISCED52uRyUdrJLwsml0sCTWsLMmouAdS3EsHszdFvnZGXSXt1/v7tGwpmpVdgx8ZV8J1SAWW
D6ed8ffIWB7RTlqOIWjdrzOW+4zUdQMZVvr9Fw+AFZGfCqVAxVutNNRUiOEr3/73nB8TKps7yuT9
SwxN8RKljFVAl3KOMuTnSo8ETVT69ndIUmEohlSchQBNW4wrMyY5gbff4B5dRIi3yD7SmxIaX4gA
V42YUIJNC+SYpylTJ+exBoQMn8IGt1qRjc/xXqGow5DzcKkV9jzQMLH8n7sQGlV+emHiGnL2LmjA
0OocxzgS2Mn5/7Ea18T1oOxrsAvDn1az5wFwpoK6aZ/zuSRK8efGbtf/CiOAIG7WqQDkzaQsoAtT
Fkrvsqg3/f84Xyy8/cbA40G9LBkCL17nCwwnOcRqHz3vX99ONcqYZdeZVCg6PfNmXnKVQB3XBcbP
vKyGMe9HX6J3l/PZVFfLdrXiwq3rwV4uB62de+Oye5e5j8+4kxmzGYxSq+uZ0VvvGyRuVtuNbT23
M6uDMUheO/FjXEkerQsDmK0ZFxQiSmRXSytNlbBOjpj4dUMDGbiPCRXhyTrZvkOVBYtpHIxMMQFX
Et1NXPc14dUI4tP+JCOk4KHa9fuvG/+dAThb/BL3VlOXVFc41HW8RzYdcG4aqx3N6NzFIToxmOly
4xYS297t7Iqm1ISJxp8B39DFyFgqf0Sdl+mb2FRCuOw7RKa3QgXVDTx+fgfdk8P5xVfW6LdR5Lrf
URxhErj1vMiiZ0PADFRrjbYBARExreaZDPQC+QH4AKQ34T86SkPMAPYhhalKIfY+tCdh8vtnQBIS
3iasNRyNjl3IQ8kZB6W8DadzLpDHfRZHJ4aJXAKGa2VZPaqO1CKio7u9IIsjWziRgFLBM6FpMzi+
3gIEmx2zsjcly1ttOaKv/6+b/ISoIC8RvlkZvtl1jLb1Gj1MieK7Ed8CKyp+k7QcBkEOrDNdvoLH
ADuXkm0Iky+x21Ur5rPjasCO4r//mppe0QPfRqMJ0ZiaVkmlxP7OWBippx2ZCdFRgFawcFzJzJ7I
Tob2K5c0ivJwSZYvwa9BWgbyDCX5AneKO5dkxg0IV2FyRUFYbu4czdhaISMP/Hzod6Q96TwVp5qx
C3xbSXKyNG/9wPk9tzjxtbnXLgBGmh/lXgtejwlln5/LJ8VdeE0RhvDxaXVnGIvjKQkQUrAKtiCu
ocOAXUawOkBVtKyb+U6/+VZ/scJ3G414l0DR8sM/v35JiGaIXIW3nhlk/e8OVCbHd4RzxT1Y4u5u
7Syq4fsss5+0ze/tDOaNeAuoWiAC4WTtFRnyl1PT/60sVpWPi/5EkEjrnDo3mX6/JOHC25POsZCS
4ee9BIk7F98SW9BRzK/ROLlihu0TGHIzUZlDX2B/d7yjyo4hHnSG7+9KQsJVgw9rpkacME4GQJ8+
PPnCH9KdCqte+7EoEdlgGLeWC/v5BczzdXtZ/h1OILyIryNVw2ZR7dom5C1tttkR+xvrrItkxFVp
vEY+hMLX2atGx73eSPS76Gu5grDOrhXqUVQl/gIaNKA035WGg3cL0Q+BWYCrXV+Qig/o2Ba47tcL
ljacAl5y4KP/CATxrAgE36neVaOXGX9PFZz75LtvRXB1Dr7uArNP3/Au42serSqgssVvH6x2JmvR
KBWb4XOlH7+L+DCNtlOxyzdgB4PCg/eYV+rzcruovPcLpkcgaSJ1j1GEDXRdq+AV30YFu9KrjbKS
cp9VlIL2iS4+HaekgLNZrnmdUa3LOUjCvnqA+BEtJ3vnWo0LI422XcsLRABtQpxddY/YeCBuKtW4
as3Erg/j+0Montz8M3vrrcvHd+QMGTv6QkBM3l+gR1vPMUtEruybNsWjQ40VFic+cB4AdRMdrtB9
fnpmTuJYbAI+32iNFRmVEaKTtRRSd0c09rGhdriUA/jgYHh2GnNntyAb+tqGgmUNP8EMTujst0wr
fNdKyCwIWT32K3oxcTrA8ge0m+t5fXjn2cl0hs7R4Gp88kmRKxwW848cwczfOZyov2GCKy8EyExH
jDU6J4+hxBuuEFIZkxcRMe3r3e9EybWWKwk7BcGxn2gHxBuuKnsw2L18eRGw44TEUgXmWDpMWZfp
kECP9kbiHcm2/H8P8vIrh8DosVmHpFlCJTJE332GxOgu3qUSTK4qA0zUFcN95A3BRHTzop3qGWOn
uA135lcgod+egigQ64L6VEsj9ZS4scB4D9UO1q6LK7HwXl+IDIcVwb+l1mYNY7D9FzA3Y/51GEfk
MzI6Byih6Ev5JfSFNXzZBkGmSMq6axZj7MtEAhehJAanha+5qnBUA8Vb4kRuJPbxrveOrKccFRce
4qtnnA4aQdPy32jb/6ILlUy/MjpA2+8q57eBj8+6/LqjbAnOdr8uVfs5aSKjSR/DvfZTdi4gKtd7
gUul948SwQj/WykzIk/s0l6UbDQU1F9cZ0j9kkSZYjYvlbTtkiEvDyWeF51+70xh+VoHVRrgAsZY
OO9wB4JKO+zU8/Ld/TlscE/uD7HNtunp5yMDaUoenLO7RWTtoTl+0OXZ0syKuQPEYQRCJLQobjDz
2l1TyslCLGNvk0Zpdg3S/OpU1CYe/V0L4hdi/bMrPCtItSS1+DPXo5zYsds5ik0H+rjMjYhgFZN5
Q/fKH/VESRFMHIlwP5Cch30otlBap2QowZI7SWZ6zc1LgiJ9VAFv5vyXv8bZyYtAE3LwYCB1qlBE
7wwZdgGVDx/AKfHvJsxlFRNLAKNnCa9xJePpyzuUHqyQw6K7tnAJ6lhR6gylyzSA9j4p+C664NPN
Zws8K6TfRjlXjG1PHzFgrMlXQOSTbsgAskPTcCXqzj72fg8sdu5dyZvMnQ/5RRxMXi1vLP1TajJx
eiraJegrd7c/8XRuCiwv1+LOGKHxqUk2BrMnbQmJG/KDkIT+xTCWUObN7c0PwE8efGbTigaRYM53
76LydNm6LLyeX0b2v4vmTvfZRfnbxI3NTNgPRH95DOT6XhyKRIsUgtghvlpSiaEhOhXUPbYJ4mct
eTE6x4hByu6lKyaFgZHbg8k5sRfRZEUoYMZwhRQhExuXXYS8smriPe7e+4SzgshtFi3G6TgZ9nUD
a1hd2MAoNK2UFsJX7TKf/Hbi2Sdi0PUUlzAfRxgGWR5Z4k9eSoRB6m4oGJ6US8SeTQCvc4UGeZb8
Jb7rztlmh6ZXdQazmlHuN9artosrnDmwoRTsZN2c3PUCjlW8tfIgatNMo4WQ4kLV9Day/GCeSwg9
AhmKofRUWxWI6EMnWKh+FXZj8yekSml7Rz70utiXH0jLDMSJ0gEmh8ohGJPG/a+n1QqVsKtOZRll
3gozoF+PpNYAnprnaNLeg/MFtzcHq0gH48SIS4HxPnxPzt7JzL+ESmwtX2Z+i2Y9lcb9Al+G8kB5
XvZzNwBuKoW1+gKa8kfGDGp6LXGafRoR9JqfN7oPiRhH1Lx7/UQyiLyR/uYgmcr1btrWsLaxvt7J
23USlcXN/d2xINIiCO+hK185qCuFwPdz94Xl22UTQ/5T/nBFMikqdEVdZ8QzHFmZ1XVJlVOJJDWX
oax9avIKTIg4pckKlztiOph5yr4RBHtY90y6YN0uqNP1fhwlVd0LUa+1OAl77VrYfIG7iDcGwoPQ
diKdryL7sl+YgHI2/LVzyQBCamUlkHzIXwgJSFbDl7YPbFH9BXwaBZNYfawZZSiFdlEMgw+dwPdf
exz+FG17XbltUVH/SagoZiT1c7I29cS8cFv0Ppzfz3v21SHkGwoUMpdTQCswH13zc3e9629VysPC
Zrj2JlVo9sUNtn4GIi+Zn87qJmwu7dmSQYMgFBIdX19jfhYnqTajKmxabwVrRXPmqd3GbdyF4QFA
gGCCFMrOFtr5Sy64SEjcRe/oRd1r4Yx4QZJ5CqM8KHSQWbkZf5VSM7BMnETfdiL6CFIkkw7bFHGS
gy/1KmOoGL3PbE1wxeytmUOnXtz1r3SCZaD9RX9VxgEAy7odiTNfHgNvFIT2Tt8qiv32JsuYkc74
2ioDrd5DYav+zpwXI/C6PONk+0Y8GeuItTbQ/9of33HYoFZvvDJ41dg2phmT0sAV0I0gUSdCU2aG
Mvz+r9CGObupAtL3WMsUs4IsnfF/KDqCpimbWWqfhxFvmpZDtjwKUbMDaTWOhL+bpbN/VClLG7mP
bH+S7/sacg41tfZEyK9k8mNA3q0IP/O0VhGQYNW/MVB/4xFdCIXp+bJq5yynAsCmLrq/ROsRinhT
utvUYwUwP37245Xnrp5jjzwhID2cgtos1efVXB37/dpOS3Fe17fUywN2A2qMXhuOU5FBlGoCzU+p
qZtBdldkf1ny0d/l/JN/+1Y/6cjfAw3OlAU8k4HWtCIMAPjcdRN7DSFs0krmpUaJCkJG+S+usNln
wbg4JoZd/XkM7jMBpL/7ai7wv2yvPVaGg50sU4EEbBHkNg9tJLsH3UHvgx3F34UF0yRF4sKl7bmp
Voutjyv6mklBSz2zyhYAV3UfjKEeVudjQzIKiZklwP/jsSzU2gsUL2AlL2VzFkHlhRW0vRGC76GO
7smpBX7bw6aIdFT53+LgJ2QzCLK/p/rLFSBWPys5XPjdLoeLs50e3ueCld4ASmbTZC8oq5hvWhfN
u29k3h3xdARZtu0hbnG5r5CxvGNwHIqSJOOjgSRqzaDlaIdvzEokDE8QOwDeFMka/NtbrG2pZn94
0ozPr8z4sZsG2lxTILa0mYe7nL6xkca/nvD8+eicGibxLOswGyN1UXlrDbgpYwkz0oJl5rRvDL3p
2B2AOROBuIMKZRQ/UG+8C77fhatThtoksH+Ru5NSP+Gg0VX1jIPP2teAlkzCKNQHnPW6GdfhdtZd
2KqtctCpmUmmc6Uko8H3UcHXmklDjWsW/J/+1teJ+DwLwrmQAh2sFUz22Tj4w3xWxUF0SWmW/gjD
2R3Pg8/cBx/spsoFBOGQW7YchDpUDIVvO26cEetktPyoIFeyRGGAh8r9Qk+XUDslPt826w/AoM+9
GTASi/dyYmXvwrdb2XGtF9byQanGWP9qOB57YfDxXiT9yaoautp4hNysBn4hlbQMsIUivXsvar9o
2WM08Jrb0Hzac1dk1/x4AtMCR9TI6d3ZUu4Lr09Zqy+G0eTC7PrJBFOelzAOKcT+1FV+FAwSon0d
p74t84NuIPacWRbKZRV+QaJXg8XpciOEZuSTtxtn1UYC4R3F+ucmYXeBtsQMKqEcfb6P0x8PI9Tf
7Zr/hgciJn/aUWV5o/K5VLvqIqr0cVuiDV9ZjqL2nPbhIkY0aCaTeP3OeRtJtBfsmFTBv4uP2pen
fxu39QbZdCSSfxyD5J1rtRP8O70PtJrl5yeFxB9B/59tGOUkutp4wCRyM9JUDLoOzqlz0ozYaPtj
r10NSjC0wEZm/Ru1xg2PI0EyoONI9PTMDvizs9JTuUia+DnCp8iH7yYirwgoYnHf5DHsz4PAQQ/z
sGKO6mdlhO8UqOKKKbJ2bMYvo/YECjljIluUHSBz8k7QcpmMqU1580PmZVUJoDmOBbkWZZeZUyjH
uIyHsGCVwkuw7d+vxSnKgKCICTXpvMKTFHyQ8ttZiDSYiVTX1Elrza7/mUXetsH52+d8QfYY1nzq
F07b8XT5gzdLxq9vpSKXoHHQmVok9o+C/MZu3DseoPb15ruqF3iFuKCJRweaLiTqXaEadROxegST
MJCNnrsvcf58bfFaco9AZ+jju9wtrcSBOmCEc9Z8cFZHRcjvNGr+xkKXGoW2H6J2PaPLI6QnzU9m
nk1k8Gbi5GQB7ZU2p6GHVjk09uy4GasINxmRnt/gX+Fu+ppcHeboz14mzNvOa+MnypeQkM9z4S2q
5iIllfq/bWf9bJF0VeaFLRNPdAtVKGid1gntOpQAetNf851E2+w+/atCY7OVUMi+fYMPbfUkJy0b
sq5PF99ym0VENa+8S0XJfoRboWpltQN1Dslisc0jUSLAT6PsAYygA45V2ak0Y1RqO2vWjG607dMG
liNl6Bffk89guMr3VHHiHgEFhN9s0FjprsXhNpI5ssaJ1WXbi9Kh3xcLBwL/QS4FDvs4w5mhp3c8
3EEpcWEwkIjskhDVZ6lkDCYMJym04Us9gjDpXTbeyub128WVg04SG3C6d1U0glxFoJ8dXC/sjWFb
ntbAmWwIu3RtmEwwokrR524HVn+8OjHA8DKyPwKloPIADRECKtdPjyom3dIgtFinhokbgUqb8MVh
Nr84NdnXc5ylmQB/jvhH5aFDi3H+N8kGtrxcjmOnmtgQqesD2uv4C1beI781JND1GhLqfjaEbZId
zg9QEyvnDR3PfC6x16n6nUlpJK0Ui+gKaDS4n+KTjCLnN4B65IP3vijmK9iykYtZzFynugDsgoSg
2t9HLT+0uDmiFe9UYNH/tNBPTSjDKyjE7V7USx4kONppS09Jer5Vp9MKHhKrK+BBitmY3j1EsASZ
ATFWeiFKeA39aQsM7Fb0sMIgAhZHU4o0hjnGFvD/gECbw6KzgFosL3TG139iRjdN/0w6pM3o4JLg
YVvtILHZhqyEefvsKctWxt99D+1vCB4nBo07K9eltcZ2e/MT3Cd7A6QJd9JwilzvVxPdUDDWm/1U
of6/eNbYF3rjDdszs9oVYi4FAconKuxE3rDvPqVLI0NBKxuU33IDMetACeNY6pj6mb/pJBB3pRO5
5tK+eRgGNCS6i9Lw1giMaIL5iKW4zMjNPKKYOiLfr0aoAU6KUdkKbQSULeYJ7RK2EPvUrEsblhwa
pUF1GaqbvUZ7pu+A31BjbThHj5EaAGboL5CW7o38r2b6D7qnYca+LBonEGOeShFHPeBWuQNCMkHj
sXxj/n11TIVHYRsvpMl8qF8PW9iHrCeZTbEvpsKn01N7U2F6MR5CBH6xHIlvbmYrd+sZnU48wQSO
vtHEg4j+0eFBjLtl2iI2rBDnMQ6NOxWBSL0Kl2EGOpxQXaNRMnIwBQKh5e2krKU2pnh2r67fbOBf
D8C7Hw1VXmEyabMsC/USkueSYWQ/Herq8lDOBOqfBpWdTYvLHM2QLuzm35cg22Hy3jnETMpT3zqB
vmwr45iIRMTkp+4ZQa+QONepCcb4Z52YmMqP9e/cpoJTXnyf5S5Mjv2pU55F8AaQg8gAjoAFZiPs
mOZoU/93wUf4SzvUdiwuvSqc569dLu44pvPiMaqsjxRWM4iLM8GKAadD1yART663+TiwQ4O8PhtR
+5mOnK/FxcJrQhnkpWBDy3eAlTFxf1PBq+8EUrSGAqKMe31HT106hMdvHvzmjT+J6aV7t2qvB8N2
qw1H5OtmzFy5sUmIZdqoR2be22QOjEN5mV31VAgDWS/jxrBWxJqg0EiqH68rEmOWrRopjAEhUYQ6
O5ZmmlKep8pJtT4f5ro/1P5/pgCkeuDpvZpBK6//p7RqKWCOr1ztz8LTyEt0aWBIj6S7E9EtPEKO
q3elVwuVCL273LlT1FHjNpfnMP/6T3gOiM2mYZBC+oP4exYuZg75rz8DYWVYilXNRu9LcNi75Hf+
MCoC6IX2jF/4P8PqnxB1KyGjf8mTqQ6t1RFFsiITQNCrVLOb3dgAmlaKkPDxxw8m7i3oO0hzDn6r
C5gSGocBl1rWgvJI5YVsluXyRa8rnIx3pP6RJRz276nyOo3FPSzPBB8KArTSLLo+/6saRHHbulNM
0Ob/uC7b2uLLQerZhNh2Rz1Gyp80z0EzXtcW2SpR+bB21AEYn7tMgMQgk0DMP6Ol99+ldu8AMAet
AnSbHXN30fopz0HgizzHefHsmsbFjSWvrGbQ6FWpsP0/JebiT4BwKLIzHs7x8S/lGwdOVBatAeDX
ViCGpCTAbJvyKDJbqCCTVYoFNV3x/WFMNT1Cns0dyHjYkHn7KWF0A2YB5+7jrBQSX1IH/7jNiuit
J+YwLucWDDDCwfjIiI8qQDu36LcUoaMABVbESWCs3witqC4MCZZYDnmW+HfOrEC5OAIuXJEYOXiP
2YLGaogf85+xzvBo88EnTyXYYB7BmL7rEFV9iJW5n0xf9n/7umY+q/SafPWOfQm3zR00EThvPNMR
aTWFrK3ufciVWlc/DRVALd0WJ1AgsE+1gWCLqr1aDu3BuvT7jt34OHRJmS62vpSgPMQhR4jK7vqX
yB9gb4Z6j00PAdhwwuc/dyU/BH/Ki8utEP31VzblsVXP/gDG/DSKPOP17bpocrz9hJTrPI/QWgwl
r43Whqh7Idbh5jRA4rv3GfOIdOq1xinDFbbZrR8VZHUV7SB90Re1Tp9NwPfeq2Jiqiue/e9RJSW9
0CDYT8NKIIP2wX1TPTFtKu2osKw0pWwyihVKImbV+93O3Wp92zWXtrqVt3ua4SQVsv5D1DdX0vgf
CxlxATzWu7N5Tqu1XUqlcaZP7MDgMPEXqnoH737cvFw/oOZ1pb1YpyviKih/LbaXRx0C5AWku29C
ZgSF3zeFZjftaMXd5cm7JUK5plf3W6W4nYVRYBssUnwKMcw5k1jTXuqMvS7m4jPQnLVQI0AZ9axS
+j1wGnz68T6aP6Q3Wzb6wX4WQThePjukDKty2k6EHphfmsBIUimzgmm9f03xNxV2Cl1dwE12Mn5L
/QBmGm7qXjLcCreBSSpAwgy8FSnUBmetMqEoLvf6hco8sQtUuYw4mmRmrHp1EKd6yu+UG7iv3MAV
+81dgHaBtSk1o/B/3xVV2W2PlDGuUpr9JrA9AiAtjZErq73UaPUEO8ky4HAMX7dnUOU+nJLNMGf9
SHMHd9/mNd1Uz5p6ufNXJaHIaalr3uXaSPP3NyH4GtKlqO3UWzdscCJY+an6QpC7kuzpV+x6Xt6o
cZ5soCGtiLtKSQhyCNf6QNcsAExh+L3HVGot8PpGpuWDxGJG3oEWyQJK3BFyw1Pv/1jtZgHRfuFT
5d1SYimBfXAhPN1kLwIsqn/Ga3teghUJ1DoG4KL7YuNwnCfM7tDLVDlMuKEr0UhPYaaJDlC2YVOK
GCDhQd0cGj3ysB8pHVifba21JzbMIZxPJn9UVZjFPhSwQj26qs/nHp6b0cE26/T0E03dX88Xhh8H
G6/XT3Al0LFB68UL9jLETeW8FAafjLcYyUJo62m9lyR+w1Ag1Okm8wqaJa+QGX25DXPU+9Qf9bJf
+UVSFOBcPxK3t3ADRUwDjl/z5TnaBINvMniQScUb9JYO8WAmFaLQNQh9RORIwt8Lgt8nJrTP0zuu
kZYzFUUIUBQypoba2cWmXjPmBuR2wcsZHYcsNQeBjB//e0MsSaTfvBFv0GcsNDvDuQEUbwCD/sNw
HOUVQqB7typXpdfjXfNcseJxptKAgaGv751zoiz0Qeefg/YbBv7AM7t6EiSsOYTyoYnaj76LxD+8
jrmk/RLF2gLgsan1QF9nqtYKhtaOua2DcAtLfddznU7+ZobJQ/sHjiU2osk2NGxCUzfzaJjPTyyT
4N+nFUVsWamuR8c/nkNR9k8gSo0MieOP9jSztMRYXdi2gBdoYhkiR3mfSPEw1DMFsQu2U+nLliaO
javh7bJKnLvLr6gJHklE8P1yyS/eapvkuqSbrrShoVZq5uA9FiaN8RolhEWgQ8RgesmY0HV7p+Ct
EK6qrRrPJRgDiCZSO3jT1KQaH7tAe8tSee8uHcgUPjBi1okuDP9ku+v5U8uAfRTCCdzay9SimVix
aKkMskTO8fyKsptx9SCuamwKQ6QUfzTI2tMHipx6x6C8a/TQdF1tcjlBhk1PzQe7uTMquFG8ReJh
1/C+s11REIOL2e2x3ZPo7B5WiDQF9qqhYBkqIAnKE/di9TJ5K3OXbHMTbTC3bS5Vq/XZh4bqwZaX
gIU42xfYt8wlmQqOjfMN2+03Qz89pvwWV/CsZmxJ6lban/RpoC8yhLRiJFj1H5MNgpJniaT3xUT8
zBO4/xg1cEAdzC95clr2PYR+78ZCG63XKg6GLeD6V58IS5yWACq4Ysm7L7hZ0i1OWH3rgo5niLhb
OVFdmlYOx7lXg6i5ugL7p/sAoFA+mOHEG1couJIiXU8mZhoheObJwIabr4u/wZnOUCdzqcTGdAY+
MZTN+wNWYqXyDisXW4b3J6Gw9F1A47e2Ui7zTn9Gc8PiFpeXorniovS0RJ9xdEJqk/UuEdiTl3A6
sox3samN1dbnvsM4lnIlUl0JT6uFWdPdxRLIw1y2jrzZcyKtemyONanu73NSMSkBQmvMt3WLtW4U
2asGLzDOOEexYDwCjjaArr7at3sUqkTaMkHBjqzFtU4ZDSt1YRXBcu5gxkQK8ZTWC3DYgN5si8k1
OhYd09V/xifx5heGpMBYZCdH3DB/tMO8AFf8e5F6LVTqZ7tV1FvLDQklvZ1Fr8oQBqo0QfxIDJCn
5JTtRpUy/GTFwzA0oqGWVsdfHAqn8MeClusYvb62o30rE7bE16a9+FnGaUvMl0BPQDm3CZJxw/Dw
y7ZLxFPMmkZdJhTd2uUI2XU7KnHwGz08YCRMCwX4GiBeNCP3PQI5W2kxabuCm9gHro70apZkbHcP
7eAG8ISCJYoBTgmURanZV7slHC5lLVTCTvjQy+lUojqLddVkrx/JezdA1jfWPryYkmPjj3Fr5ceR
Ga4YkXvY3ofiB/qUtAxOkx7yMIINvACW+uACPcDhy1steYMTWJv4j7Jsfy50ZqStYmbrxsw1OzQY
lFvJseiG/Mfp4HVR2za6PIDVCjaXCZeaTAfLgEuZMeSOVeNov3Hx9HRpgJKbcwkefLlXbPkPRZrm
c8Ks8Gr4XCzqxqDiKzRkhf9wr8PBbzf+UI+ZwO436f45NtM+PIJtfvC5zg3X+3rs/ZVUnu8TaHvN
5e4O9NHnjKw3PeElYE+pIf1PjSCG1CDeikTrLJee4tIg9z+2FzHrlt49FeNaPJMmu1SCLASJmjjD
5LJKSglG7ppJBN+5ElGUVTMkfEWzRFn4EWqKlkhndCF3YP/JNzkLDSxToinpcS6QBWr+00lnZQO7
g+bnr4dinhoi5cuPcb4jGKsvA3DjPn37oJ8SUz73DsF/ycRLbg53CoOWHQzVJu+ROgi5wFpzmIMW
F0+D3p1ZeZNNsOHeBL78q8svgLM7Zp21Px9Ci0kXENLjRoPgHnSpiZxfxj6qM+LvCrbLxF0otz0E
HGpro3wzp/RvkMqx7+8M2wQIg5yKCjMNPZnxFokT6wgohpJXFKH/TgPnarKKb/xKiZQ+i5oNGTqj
l2yvF1bGZKiQIVIxnV6noGLjB9y+KEd/lt1HxsfVsjQR3w62zvxNHoOp+T1m8uNYPg42pGRzuWl2
tPuRCZAwsDfJWm8GuTT5n87izxa2x1dYmf4nY7C1Z9E9J02cvtH8y/BnVrN074A10r/eI32+TRtN
y3KUQomjgNbaJv1GDO4cmcWTyV6KP39GFlDCH9CoGYtBKP/WbHmj/iwdHxZ4rtdG2nCcDSX1zK6G
I8q50Yf2fE5mwqsMKHMk/T+8HlBnUekZro6NuScM8ydCZ4SePKvAZvhZpAqfMjAM2bEVAdYNhKSC
Fj+1NJGV0zR4WqSPY+XG+KLv3JVrkkjjNJ5ewsz6uHJmYA1V3LQA9sQRO42ke9GkNlyImHdYrVSw
X0GYcWi8qthN16+j8/3i2zr/6BgQdLLVu2fzXMV76EGKF/IWhziRmSEuXeJSjQYcYW+6fFcUf3LH
74D1Sl52g4rWnto93wPfBKcrDG+u5pf8INuceZw5FzicXelYRI9HEqmDJBGIWMtce7wJAwBa+qZF
IJHe2LcbEmwaawtBKND0wV0aDmvtu7n1qlmnH5Vri7D/cUlPCZwCk9MIxa6EAr8flrWJ8f7yt1tT
UzLVjkuz2N9eeWHphle08OuPEpxU5nq06bNHrRzu2bR87G2aHUWGB6jpdtkAQFLCVTBI0Ft16xoK
hUZukG7WeBClo4J82M7aew/TAzKWnsC0AWYxcGrDsPSaj5N13lWCfbSYx3n3wlrU+3muBD/OD0PP
qDIgLsZ8dF49vNoBR2szHyKJ+6ifOGNFHIdfR3NtTVtHFohwY2OttDi2Yc3VPZT/3OLKXasmT937
XUnDECOsv7r4t9+e0/tblafqgds6UZf1TYYg6EaKi6i60wVXnGbwLXXaO853Hud66DsuZ3Mk5rfl
p6M3eCqNjVxQMWreQxCl6l01/AFRzlqOGtTIbChnIMyM9UGytr+IsRIhSAZJmckYv4dcG1e3bpkg
5PjdhjzBcuW55ytPkTqvcHzLjtYEmY6Vjd6NR2U9674qL4DLR1SSU3XDvIRs3xNFWrqvsUQk3K9v
gNpWsknUmk8FiG+WrRvSiFKvxmR9LXthJvazJwQWwPj/ZTtc9xuFqcbJ7BayKF6r9V1iBH1QBAYh
j6LzgVTFVXbd7X5BU7SsFTskKHyaiVS7gI656YMadlAAv0rqMRvW7T4fTOpMSCYpUvWi7vbD5yWM
dRNoW9iwSTAoZM92iLgHgXI09m8PlZos2/7DAYTvfj3De4cPpVMys4f/0DRvdGjE1mO7AOiNI5Cv
AHixbcXljqUawUU97z7JiWar75NlNL02xmCjn+n4poFbFBuN66vjLgy5udFAjGkGgh3w1MMmNOoT
6ScCiXwb3bSvXNv9gnxn8eqOOhe1be8Y7wqyVy6bdDgq1BDLLfEX2KzqT+wUpgLS+lhrLwZwqAsN
w7VQpimIP0S9CXSQQ2f0TuQdLccYn0dyshBzjwMDbhS9JOVTRRBJvFDmJZrD7jbvwPVkyTqxzsN1
qSf7IvXs5xqZj39vDpk6EczYmjS6UPjpVvECXnnBc7Bm+r6VIA6XTH2mfKyc7d3ZVIxyjQH5GbMv
fZXzSlH4YOKbAaDUd6jcwp30zhjbxoupopyXWhvohPBicwABKO2iv9eAZkpmwFeDizT/cfdVfme/
oQ4xrc3XlgjDtxxBdZCX3sa5iirujQ9g5lI1IrhLyBiynVvl0eovYGmmRmq01aYMeVGvo6YKsTWS
vIA/sayFU485pKNbdKhebwDTN9ts7WpjYKibNS71JLtTnDDL+COumF3BiFPw2/RvksyDrsgSjHc1
7z5JZvoBAAMsktBTv/qM/+nNJt4Sf4UPliN/yiNHXhknAk8UvvQum6e+/9gNgDRQuuzq1Gj465yn
UKKeqgc7BuNj26jD0w08FtzSwoYiT2INKI2vXdDG7r4WM6JZYqUNdSkioI9meVSzOOSx6eSs5wxx
Gi47lZiyEaJDPs49XLVVfOSrRJKcRfR2j3cTZXAn+caZlIRDUDSLc4V9foKHeEKeb769ryNaA5lC
65com/6FhXkWtqW9q9fs0SeAldurrn5bBV95dMaelEU6+WMJgCdHVW+4Pt1wSvlBL/vJ4OwQQbFr
BIsnyiTWlJ8/6bPHDW2Z2EP4CDGaraWxfjuPmWb3L86s7bao2jvCIzyjTalbPv+Npun+3C5IcKOE
r0wciWtbxknVStGDlZG/R0rEt2HM7IaRpCaB572/k2SqLJZY50hh2x11N/N3nV9gSf/qkuunklHr
+hlCHXAk52vLIvJFFaPZRN5mZwZ2gCgSHV6xx3sT6ksce1RBjPWF/heY21e7oCt5cBvjU178dVYW
KvislfA6dk+Us7LvFSbrdNAntEpKQkazL8W4Q9Wy1YARo/6a1HSJph3o2Pgc2kpy+P/XSvke1twd
RvqYntaO1fAM5lunBT+Axf+saCwVZLHs31sNdR1EGdG6qC6R3PfrHdSL08AkXPB9A4HkfBr403IW
fCuD7RECXMGXwsUTqknj4rg708QuwxmH2cLhpQdHQ/fZ/m/mIY0/0E0fwoPtfZX0VDk39c3/014F
9xs5X0Cm/dU237P40tHfNQ/v9kMWHoiI29qZlqGfUA9odd0YZzEzEMIJlGqcVLDqoeJdjWJfhyR6
lpVL5+Ur1wtbLT17FukEHVgwQbY1q0gV3b4OXv2mQuzcYEmRuKpiuWgl4UVdadTHina0ZNn4aBQw
uoHeULdpCeKDa4cmeqIUgQZza+xX1TPaO1Zb+LUFY+OPHeaypDnCJvQql/LpH/n/njdus1g5Hwv4
t60Z74f1Eov7bgf9BnzLgwU0W93YhQV+4m6HLhZsb8e0/yLtX4UATZnbq3OF58HciaeBz2Ac2jsw
2SfQh6E+AEf4zXyv4m9vimx6HbTQybPA/8n5wW3IDYgy/B283X0ZrhgXLFOgIQ6O1GRDUT91XDnj
htKXFtvqLwyJwFf5MC9x6c2lNDrluUrw+SFAtUAwU2MB8TCBq1hEhUfHWJzYqU/Ti0ckaB1Bflqv
Kyis+EtdI2TtQiipolruxUD36t8m6QPYE//GRSN/A1qAi4enqh/ZwenNI+x/62WntRlVcCv/kzDN
GRapUGeVpeo5LPq2jfT+5+jM3HeN6IHrC9ohF8S29NK/t0dDHknQmMWLdAFk+yESyVeFJmfRnlcW
Y/nt5hM3vu8WL1RbsUlyqC/5adYXmy/mURtrWvNEjuzbtv7PkrbhacmQpHCwcIqy4Lp+hAQQhAZm
HeTSlkrxeLdzEeOl2EQVt7VDbHPzVb8rhMfyR0GoSlqI4tsvsLo//z3DnOi/Ie+g1ygUJ4HjsDof
KF5BeuIOeUDcleeq3jvDCtleeQOTjD6cMX0q3Gxnyk/KSlRpBVAR1oWzJpfUuwydMXPmVdp4wWc/
1sRhX62Y45+Zy9/tiO4ELIR9P9jmhVGpRDWQ4fMkDG5MdgeUQll7fVGwwNRZ8/736aN3Fsn7UiWW
MJ+P/HLGsrESBGBh8NwgaFYtVknr3CFD1oSWrJEJDIgMjcpVzN+eILE01CQ84qOsZhG/yLb/27dE
wIAXnZNsb5dii6QHp6y9/2g9oxlshGoH++UJnyzmyr7tD1wRBhGLoBxNYxRwH8Vj/aRrduT3BiZO
e50CTLDKX4hsCqSnW6VCsOYQwNgR0T7o3tnLhW2icO46TF8VVFktyWN+avPhuSQvA5HVS0N9FE4s
wwc1r92Rk+/7a9LuqquhO4hJ0BW60HsiLKYUGdWuEXm7hbCXj4jKX/za7jnrXExjrzLbGTrQkU1L
bgG0BkvRqhy0doHOQxBm4UAiU1Is3vLB+hOoDY4Q//EwEsIEiOnxCNqnhm67YewWy0QBnJPQ3gUX
ZsiZmDZSCXyG/xgkk7rORWxqd0PnVzEILy7Kggj2XyRKJFyLpq1ZiZwIUjSFk/8dVcNrFsBppz49
KBMdtVfgsYZAJtHGtAjetyStdzFSiA2prWZFAz5Yl6OCDU5PAia0MtgTHV3S8r/FYTQ7nuceFyiv
VXUkfiKnHWYqC3xv41oMGfq9n3ZMnkngrkDYxsXSWEYc6pDLV4UwRuBNLGip44wobf7FIEcYQ/Yq
mWPwzwN8I3AWKamR5NRIsUhPwSvH2s5v+kNXpKKHp2tBKOJYmm8XxOPtCMpdH8tc+2ALalrYEMc1
Mqq+jzEhz78yStKkm3WnBgoKOjz55K1gZp+4utMuyPOwqAQvUYn1A4TvEGtaZgB671FY0wnHc4V/
83aNFD2cOyGTf/fnZRPiWcNdhRF1agNLM3EUe/r4kH+mY2E+0okT5tjH1zDKqFZ50mHpGFwZGEGb
oI7V/GUegaJcIMNioAGURAqEzWUr3PTA6WlI4LYAzb6QKCJ9AqOEY3Kl9Ah2pn1AJclvVDOOeyd0
GKnjQK4QDL+nimoe4FHIjm5LaqFG7GBwIgykqbigQ3mq1nDuEGBxJR8cpzxNdvkQCTOH0R1pjpn+
1OfojOIUQPIgr5gzZYmwXLlbCJqGWpDjvi67fZoHE3T0r/8EIc+eNkZo4OGaybzYch60y5wvJmj3
BiGT0pc5e0pY58RFVzwmMJUsxe/bojKFy5TtlxNPdn6ScFEeANnrPiSBkn9pVDA7O2WRTvGe+ZIZ
S89Uts4wl5fgMU9BsdaH9c3R1Rw7gcIg0EwPJo+gdi4vmuTWvswBs8Rh7eqSXD9yORXRS2a2hc4J
Xj5JkQ1R3l50jVARQEyuDL7Vfufz2e1BdmuyD4oym6psiPjGMOPZT9QXxJdy5gGE3CpcHvAvMUBx
JfBJZoVMFmxASLCkU5ORm0Vs53pmyohBIwxY+FDQF2FePWJLUJfW0TK4z8NxRr/fcNZhnvzo7YBO
nc4ZAgvhUmllYImhiJQMNqGML7F5mfRtZctfm/i34qGRLNdhUDIVsLhiRucIMLlZsDUaNvVTtnEN
4AiFPozMBLoKaO9X9V8wJxtv5XfxrcghA80Z3q+JGcp43BtvC7bD0A3gA8cNH/MLawDz6yWnA4uW
GECRIVSJPOqTRQI9G9GBNEGryLoF3DXSZCJkSz7QWpaEl4kdiPSyIHl+51KlZxA5KsQHKKTRS4sh
RBwTfpOJj6Bo3XCL4+g1ynKX+1Q6fxxcXfRO+Sh+vNcJu7ONjY8a5uK7oveLfb/4bXy910krkdnL
cpax8h2t5C5K2t5vkiDZM1fa4Aaq9jrle0VsR6DgST4KfnUIlYEyJ8gQK+3j/kv2u1WXF/rQbBdU
sbUocFKrWi/qpnfA8/Kx9BYfk0idjc2jfxjZ4ENtMqI3AF3q2MN26KmJOW3tSI+qRSjA8m4qB9t1
ZBYxbp9Q/4QoMzmbmj22erqmcCjfXQlOdHmzH3SaA915N7Ye3MynRWu4Cs+0oUaa8CY834NcK85h
RsjzVHwhboUmJ3LXIJsQMpBNYHBO1YGzProQiB9rJPxypqIXKAaNwMm/tlyVa7YUoLIaFDz8epKq
UUDSgF5XSN1TYViU/H9LPqP2Ws51sRbKXX/Pu7AbYnZtmdZmPfbRrQXVQ4mv1uWuPg2dQtG0Mgiq
oJNzWLm4o2jy8pI+DXoO/72MjmuKbfTs7AmcbyTY+dFr4qggtmVvPt08Y9rMc5DX2uG8J26oorRe
jxVpWd+mKOdbmNbhcrF/H/Vb4bVa82Y7v64w7mWviVvbLJWapkbExTiWfqPJdpBI0MwYso86gQ+0
OtRhcCXOlVH9W5RB8YPKJbFKkQ9mALZIXpidV6HPmdFkWqtF5UQ7GX0qh7IpUSy4WzgSU+pl6Uyu
Rhn2CzI2puMLBg6+Zli9qwWLbRR51wNjHry4JjR7LlwGAELdpAk9GYDfAEH/VmxjZq5OvmOMUAQS
eZHeUhPCq1Y9LjgZy7fvJeuq0QmsFM5BYhNjIUKS9dQeQk7e3tqZ3HOewirdo+a7WMI0k06BHB7d
SXCm8iyt8/Zag3mnD6a5ViVsp3puOxqTiU0vbqXiPVA9qL0PsesCYA2XPjgxhnQKleEeUNM3oxaI
kzIOJLoojnJ/N7MUsJAzGkvOr4Gw1kGMa/upqQlAYkVqNg7N8OpDfgf4bIsXHEbqClw1b0/8m+7Q
0A0R5c8qgomQzGjaJzJW7jV3bUIES40D/Ivqu9QT9EBa/hALjx7MdqgOq+0OnFNnsUhFnQH3xNUD
a0xWbtPbu5963clu0g1D/5hJmWDnMU80gB2rZMXpeF4Nx2DfEUH/uV+RNGAfJulVTDkRX8Hsn9iu
mZuE6fNCL5jefjPBD2YukN5IRD1JqOsqX4/hXPxj1C6S30CBDZSyV5QPEJX8KkXxIwn7iyHaWb1o
PiK8wq4JtlqrS/7QJ67RzUCo9GZ0wnSJ7dPWBsFpe2FK8ss97mvEYJ76jVUDZQV1fArNOJ+Onj/w
RFjdOAb3EqTCggUAAvWFUAcADNz+cxdEbW2mRqFvHqQDtEMGsUq8pIbPhDZbhmiPsJWa2lRuGEST
pBk+yZJsQTHVx3oqVJsViHyBj7cC6RqARPD5n0ZW6l1B8RDB7Rbmhwk/1lxr7TkG0laYoEX74dGM
2m8Fd02rIa+ePlmzbW6ckxurdFWtHaGWTY9gquEBSeTViFjRb6DBEB1dPD61ThpS9N5mwXtBcq+B
ck65Bl0/QQjZAHNJLXx3p5ELOG21QRHaIrJ3zul6x+v3ASFdsCYah+j7VJSVmeHd/JOjKz1TuVXE
RNgAa/E2mqN8Mo5pzISR9dxcrajQrOJnIMmix6w3CKVn1jTNEnBC4++T4rcRxHbUmzKjZUnjcwfk
girlusHbXTSWWW7ZWF798ih7pvLjxxlr/X34LnHsY757hm10Sdq5kfYYSleVUEPD52p8lRmzVVp5
JpcnxQwfwTlQy1jm0u0qhw3xYPYJTo3lmvuc8QA0Nn0zMZ0IDVIg9+9vTwLhQ9jKtzfAT5AyNFFI
D944/LMotu2op7wfOqyCg63sMpIoHgprnGuEi//4e8GDVSIBisuZ+KDPFs9F7T46I4mpmS//TtXw
5L885HuQzXMYxcl/quswmcIB99c9UV/WgBpy5d4DtBCOcQvP9MT3Sx5CVEr/abYwum+E+RrZI5Mg
lggXmqBazjmemIwba1Dr70LdAlexsNm+4ymE6dbbgauAG36CFIchJ30fwsDM8LNEw9RosPrjIsQH
f/xNWtwOB+RXVcbRzAHvf83SzpDNMALoM7Tr/6ocv4yuP1lvbRJOQ1AiyOhwZP3mMgqye7FMD6bt
99dfDjHdWtBF9F5hKDj3KaCxrxSBHnwj6H1QaCisI+csS80chLoarDOnsuu8aqYPq8u4arc3w0WX
akVSsA+QXruP5wtqpnbiWh1wuUv2nNXXIH+QNOEPvSZw/pQkzZngB7Z9Yp7DNA2Qq90hQ5xTUr3r
a+dJ4A51X7IPUly5jozqc8HjXDbuMTHPRV6wTgAbIBk6W8SQny9bHltwbd5MRU3ms1JZ/b39Qjvl
r2quv9+DQhu6AoMYdh7GR14dC+1IW/ryJUQxI7N+kfDI5j1/Ls+i4Tsa/PhGSj8pIuLo6+8Rz4tx
at5IoutpJfOPCn5o1VuXCQSCdtJeGQWONRautWJY7m0rbYaakF+ZzMK8Kc9xMAHkNkWiNtvGs+sM
S3cdJ86vduUY/LNfBoF6nHYZ7yUV8JvU/GEQVtwfNFWcIzw/ZNdVNwM8IvwlHI/Tf6YHahdtJTNV
8jDQrX+Po7GvvSY6lesSaZYpZX2Xzxsj5pPTzZ7ussSKOCRx19hVKVwhiiANT5ypVArEJs8UqteV
dxT73BohFP4lrF5nyXU7hPz+bQNy53VSaw9HU5V/3B8vUe60a3noJf1A2XZ6eOEcEPVO/yV71Cm0
dB6vhmkSyU3lerGtNwU46iGHZF8UIZra9x8JmPTCxSWSr1+Tue1t7PbfDA9t4wZze6hZQDzKjVXB
Kh6gTgvSMOevEwn8IFyRhsD4mSO3QgPWkTXp9zfHgMblUy2YaqVotRNXN5BhIZDwOFkwCq+fciky
bGBZB4KoDc8oYB2qZCh8Uf1Yth2ej5GBqSuU5lK7DvXwsnDUIqA/6zbZQvI1XT+uVZm1fzegDM0s
VyUGZGaKNpB2SUkHgSqQ0GGzkbM3/M3Ueptt0nwNdAO8qHixFoaRtIMqRre/i20UI8Pp0ZsFCZWE
B37QkN+eF5gaEGD/c6NdYUWvsmAmXLGsnVNwhVb3/jFFsEANZyv2cG3TnEtJyW9pTjX/vcBvndgm
fHdqspUcucCDvm9IOsbQ7KMtHtIkn0nmnPLCZGDKxw4CkWIG5B05+qAnOoMXObjjyQC3mwSucYix
jOkCOtbZvWbBeXu7m4cn984ky77yuSpHwN7dW6vrKD7J0MrIHmEtT5rsIBJ6SD9owe2paIZYPHPg
0ZOJ7xhKSGCyaCHmvwZ3Y+eB9z4tv46K7tJ/UT5/MY/2+joB9FyCrZBCD/G0YOXbWgPASeDLKlOx
QKN44D84v3lIOVpnNIhUAy1U4a3IM+FbqgR0he1ike0MfP9QFsT4NFoMivv/7COsqDLVEhXVZz95
ZYcjmbB0TMypQnFV8isyZbk3TBVmwizhBmBgRmEV5OQw15wmSnL1LajjIV5AEu1QYk8uOQUaZ/1b
7wn0dKBQRlt4Tp5PbaMFT/KswKUjU8OTNkF4qRozbZpgDDP7c1zeAnAadfpvTEKJMkfuAp9SkIxJ
aIuL1LWXu+Jg9eUwIYODhTKciJd6x17Rnp9p/JdGTP5hC0ony0qSWqCg77Jpc68HiJiHTknmKd/I
05bJCuPR2YyOAbMtx8/I7GvEzbszH/uACRUbh5Z6zouRhgO4KBNAB04NxweePCnJBNjC20yPcJWe
UTU9Hsh+JpXrKh/hJSRtRmHVV6XAa/f9dhiyi0tK+Fw4m/B3jBp7/yj6zwOJ5z7KI575g4EmZqZy
JIXRNeWkqFEefCjwBQfy1KPN+dDFfadkd7hz5fdRHDfDv0ftRYnEDMn9c2JvJeiyoaNrHbLCKPOg
T01a1jTtDoHXajfG1O233uPF6KHWiKGUOhBK5klO0CTw0H9o2Gx/3vq39zGbKvlyjhmS961fJ6kM
jh71eosIGWsvVPgiN8m1n3dC4ZET+TCfYKEekrTMJly9XEJu+BysGAx6e+AhgS2xKNA36BZCn94m
f7pI3TmSxdSJu7V89ZEUaVBpC+F7axdrbGzjJLcCcptfCU9cWB2mpjbOzSENyEtE3r++oJe7i100
LAJLNZMMBMEYs0xw8S9oIDfdmfSTXGdRMba40cy6CqqaFeeSZ1WpJJhGjb4LFGpmlz1sfBOAn8Ps
RNVPXnLsFddvUQcjlssK0RhKYFSTj5kvtK5kTU7dE6xyZwDqi9G5YgDHqXEyZxBQA0597C+JK/IU
CGLzPpMzhVnYUrF+YQngOnGZBVC0S6bwwqEhp8czE47StEsOjYEWCPPWFvgNDOoaiTJYFVIrjZ9j
+O7rHZvEuuXGCplYqVbEv5ndvD89rxU4fiTiqMiU0ewJ5z65KLFzbvjRop3RVJNukR/4DSM9gSgd
isGNyRgaL2WczYi4+vsG9MQ/LTjHcND8zixmGV2Q23FXC/W17BgNmqzCDu5lUntpDK8YNK4yv0/l
JNP4okZGWb7H8qHTodinAljoYFHAuiq1e53cMgrEyGjbr75lrIwFSmvrOV8ef8c4QypCWC2ktKX1
5gRc87gBaAQUqpoy4MiJtJKQsT5mwOxnSJ2dEcvat8Z/YQn7cKhyo2o3kRpAbbrY/a8Jbpjbe0Mu
sZ9bK9/Hh/SM4+LzldoRbe4iUuQmE+scMxp4umq7P1pEqnsNqq9ekDpl0Yk+nOdj+b2rBujB7NxM
oK/YVyceM4OBHk2nUre5S8pBLIVrDGKx8GDhEwR7UVj7gewFzrw2qJTXwWYYHKhLr70xggoquVsM
BIyx2hh8t0LwUjSXVltqUpIW1Ld5/2lyrlnf7v62PYNqKLy1/OnVidJ+P0SOdxZCbhDkXap3ZBZE
G7+ULia0nTRaW5EuItUA2tCvfy9ghcn+UaKgOzl3fn5uRR+F6lSnl97wVPUP/KDINUkCBlst6LE5
5G5JekHJORzCg8mrtQdX/rv2GGYGrKzvqpz9CFfmeEkjXwexgKYVNukQPnM4tydFK+EgLIf2ZTgF
73doLtQnj0E1ClsIkk3svIjCARzaB72kVJhkji/Pd3xtMK7HJbza6YDnP5lk3pjwonwj3pzfX7yS
KEk8Z0ld9j+jqHKwqxcR3LQ8CkfSaRUgVGM/0cRngMlkxWHU6Y6wNcteR+MDy41bB0MdoZXmjbOt
ay0FzJKz4lqIbuD6ngBdUbvLJov3QVI5+w0qR2tGy0cmKwFeLurjw6oNJMRPG8KoBIKR53aAPN9w
3d7KvNV8LzpnhuXDY1QcClhYFI7nYZmdMo/qFmpnZZEi1Is451S85lNkwr91ecK4+Lx7cB6fUvIy
3Lo0vP0txK8PowqAKWDw2HBD+J7d7epVZ9AVnKiTwQEeYP3cDTgKHp7MiN6sHIu6IdEAnGY8rl7Y
lJvaBsv64t/pf7Hfaxu/uGWTZIOlHwIbs/5y8gTJYUjs/K/w52bwhJtMIL/rR/rHDM85rRfLoCy8
OG480Skt91ek54S9rhTRkU+l6CPSnXNtQN3LRACaVahVA4ETWVm/GWSDeVOgej8KZ5jNjzw7KPWU
XgyE/Mcraa/2gV32guU2R6XCajcULHCFgO8JkYkfOnxGa7o4xEj/67X9OBt1ddcut7Qfr+bnwNWW
EMSemB+Cq65quq+/4tuPnY1ZD5Xh935wT+mAZeLxY5m8H/3urSNHknuZ5rOIDvMqHAat0dfc61ST
na+fh+qjt0SMJePdCor1KqFfpy3H/XHf4kJLCkY9sxksXguRHU28OJxLBo5rvOub4Xn+QvcQovNa
g/lsfm1KjxafDXDkrmMyMOotSP2EN2NSvtNPCAv3kZ4TutNZaQml5IM/Sw2uDtAfbH3nGOe1InRS
eAHcl0GZT02bdUpg90qUb7D4nM++guxz27TJ49hdseEfFPFFQt3TsFsFm0tPVop9EYZx5N9O0v2B
80ibTVhdjOvyegmXtKPPkivFn78Xfs9LiFwfQs26xKUkw4Wt9wXsNOvGCCibx2Yc/2bCHKhMUBR5
NJHy9vOd2D59kPZxkpb9SnOGZXoyu5r40B8SWVXX2AuAVMRybBx8+IDuR9zAjh5ZSt1swZeVeSoL
5PP0kW42/TGKmVGpfeXccIi+6j4iTIQCuf28aWqKNsqceykEXnVjwl9FshAUQ5X4v9BYQk92/jCr
LFXiKVVnDsbbgoUpzUHNdA7mbqUSXk0+31I3Udje+c+vkzt4qkNAag0LE1ls9oQ6vUxYP7Kq9/oK
/uiTgoSYqlMss/z3xNMyhyCxlRzrhiBT6SO/ubdsaWrP+ADhR05XNidARRQVjSWk0X7j+FCWIwC0
Ew0hPYo5kl1o0oiJpqaahVmZxN+vNeo5L8PctPAI3rVuIz93X4MyoYlbXJFCvoyjQrRz3FzGyepI
bn+0yOEmQT3I3JR6p4VLQ1Jj8ZTLEORluwlRTy7x/g5PQwPHEai2Ab8g+DNROZyRTy3EkWlUp/29
x/Zje57uGBtTocqTqhjOJHmIHxPDwspVeysMYDF2AYUpZ0BEkOECpBRGLKCp4cNx7tQ72imw4eUc
gTTA6vCBGyHjkov8UGP9VjK7pIGrJekcs4uWdY8Ld7aCSFqu2t2DKJAZsb8bDKfAxfC9i7ewsFux
WGkqb+qsqvJTlkAY/qZs5SnqGhk52XIUzd7sMTyi0rJ9iUwPgqFHrYvNgMK+zBIntNvjrmpyGfQs
3JMmLHOdWVO8sD2y6JJAgpnS6GzvfaciwYgSuKRJXOxwvrXjkeImDdZVSys448rEcRLSP4ip9CMy
Sw2bw4zCm3x1PHaTiwbaImFMvxfx2m5zWq+D2msjMMwY3vzyC73vDMAULXxIhy/Fkv+RYA6kfK0B
ggrhNXWRgzHuDKaHBkEM4ZkgS7TtF4XOi2jkn1TcS6v1fdPlN5mkEzF+cWFGZYsUXGAT+hKXPT7a
hIbnDHiBGYFAZ0ek0dWAfF5rFso4kkYry8vTuCypDTTfOeksVLvGHzcEg+G4RxKRmChx7bS2MMwv
95ImtBTtK/7l7GDXEbcEYAxuMvzK1UtalA0lmHo8pputyoO9ui5jUn1j064rL0QfxCngMVRDDMi9
jm4a4ebv7wxBBOcuQORQtFmG4k0iJoXiylTCTlSNCVe1dWn6HyCUuiiB550Z3saO9WGlTDfRHgCE
GQetwqRQFeb+Gi42TcEgZEfTRVq+O/VjiU/Z4YPVtGYFnN+60In2oib8HpEOiQWbcbCjMljWuiga
fPokUw+tnbrW95eXffMPUFbI3d9dvQ7wQirdzGg8e4FFe2hSylGzxoLHlT+jkBxwts9L9IN2hfXD
c3xBSfoXXfUsmhUwJUM5UMDOMODKuIiVG9qDRFu29mhzAfKVKRCBEYqCjvVf9B/gpwmtCgOk5aXJ
g2nlGQbgXzdXKYeHgshQtS4UhP1z4ITcotgDBEBNr1MlJU1bLox06biAi4CNVvsx/+ewdMlcl3sM
VUWx1iCGtmg30zqVDLNHLbPUkTV0O3uT6uC+5rG7quzYumya3IJUJygKVgyio75QsLlajMhBOg52
QPj737F+/n0ZVJN9J/hPfH/OjuJCQbHoDuBuefCtsUaCdF2y6amtMembH+9A+0XVDRC/9H71lwW+
gTnHZM6ohazIxAU497dRv2y3zV8nfGjcXgofQZAjX4VaJfJOlnbBaEvaHYlzv/1WwuNwTGUbmPtP
OSc0ZGhWXvS+rSHxpejwaKmeRLj/kS0WxEJyrtQspzjGbSwxtNSCQY7ve5hCBfk8J4R8h4r4jmGE
BIQN9hJTd2GWBlrZAdgvdcwzmT6L/9sNxcDkhVL9HRzj5gEoYPdUx9rmrX8FPa4cZq164V0tEzFJ
5OrZd8cww3lLHv0xCdJpajfuy9cK0sqELEgTdMkkrHwamcP9GWuRFFt7MJ2uPsg81QzKnCTq0mmo
TxDUF2DGD2ZWliObNIF9JinlFt4scXfd7O+0ctgNAVCyenh9tBM0GhnMjxdTZ0Fynh4NkPO7w5Go
4NHen/J29uiqxCvfJvMbx2+xKU7FrC0G577O9Lsn9QJQjV/XOpBDQVaIkDX97eeYvYo11yWS3xOP
8IPpgUqqsPy0/H5G0WKYFH57iQPgqX1DHub8zZrsHUYCxhJK0gVFQ23ybpsNcE2N7AGEAYg1KBf5
+s3Mp6eBusIqwCHlnV9ShXSDQtFv0bFMjAaIfjE/bOKYFDM91eWfEziyXgnsxvvIgwUEYymzxnCd
8qEHefhc4e9XZ7cIixZuE26/iNYkECjzATH5IbL+CGKwagSoORp9tYOxSIn5xIBzQHJoKaGQ+tUs
U9fdU8t0RkmsQI3Yc4PuvDtVQTte68tKldKOodVooY34UQlZ259LKe/1de0yEfjuCSsLlelj8dDC
+Q4qUOlvG0wUI1ONMr3+4eNX5J8mg5uvayfQLtBayWqSfhJAmdWNl/h2trlcBRWwfAfs0Oe7R6fK
+/JFJ4z4LOnqrwoHTm4fguCtdGueuroqAtX74J/h/WFzLo5VSW4RtE/V6hjTHh8aRVTTs0dwglTL
G34ZLpxCkqHhtFiDFNLoIioNB8T8faBrq5rVJ+7KL0K+qoz7knegZ5QnOOcXnO8MScMDqlUTMRz8
sjqmkC3zwo56dEdD8LfBBl6MQQtVEx0KtLrpc5ZPwn86zev2/qIatbDF7xceuhv0TNPy5XpYrivl
mim28t+6wGocpBlemNWS9hr7oSlm80pqpgmSDQG2pHj2yKW8NxaOeMmQBQG8aqxfcafM/89WvGt1
IhZUTvjiKjqgWjkPE1x9DOCwq60QjcyVp8HgPR7qME/F5ZT/JxbdmOPjHichJ4aRDWaO8zpx9zbS
9JI+1gCdpcQ7Pd+a7j0KzV74s9LKu4KSdWer00Z0LwcMyQugqG5sUvTSfJwBwxVlRTdSN06A5170
QzeyT9gzMH49I/h2LGhhKA7INJ41lXUxevfw0X0JHOu/54D+BGxTbOlo328SvcfyWujAuA8JvWLm
NdJIPWVlDSheFvSqpqJXTfHYYOsyRIb4HKFfGvESHfv3dU0KpK/oWDP2nDZEIv7LGDrnHSsw4bNP
0VX/vr5AbO6QTVOhhrRzkhCMcGlmjrjV0dPxyAXY28flIdkX2i65AIVBilWaeKFQybqEn3sf+q20
hbyvJSnKylk40OGSIE+KFOlaNQ8L1FEQZh6SzbmUUvyG8l3gdgE3xdXQTy1hi2Ae4a9AMObFx0ls
u4Hu3k8FqmUIk21ZmJCeJCjx1F/mnwCX9juqrCGTKcrhXBebTi4SxQDtCepXcMrmmvg0wuJY//sG
xmbdxZ5IwG7kI11GTt5NhNNnR+OCH7EN7V0cWVppXJojigYX9bUBf7AoJ9OrMbZ/JILEGOtoixds
2jq9GLAhEN6fmFdw3bbC4DLLJavHP+K8cuR2w2tm+hoyP+Bx66xS0GGGQTaLlJ+FROcEzmKSaE1S
Ul5KW1mwAD8lzlPaBxn1tbfnwvHScUKKbjSFdOjlJe25iaY1wShxp1o8l7CED16M6VGMVXaFfB5U
KKfu+QyWWs1CYB3J0SuDEUKrFfHVb/nD8OMLhTz6kN25ns5CgShgB/aUBJT+vkoLrpmhYG+ca4Hs
/sQ9M+GnahPw7xeLdkD3WLQZdLGc+g1NbSlMYlOH/bIUZJtP+ggywZFc09QXCyt4ayDupAtMEOE7
cmic+Cnt59YzPzc9+SqGA2tyZgj+lTDn6ajJVT+tZvflQTGmmmggSP3HtD57yDeIOI9TL7D9JTT0
dT0t/6gX31Rlo4oJM6HqfxeeeZIh498jv64hgbpa/AoOTFweEEY0IrffZGjAQp+F+Buqar7yeltK
zvbf1D7uOUt0BjNDYmuGhjO4ipUYiXXReHsliTk6ICKhA9kIQKPHReTE2s8e0UCA61bGr22T5q6j
jfwZdADytEH/rf1AVqDBi8WkD3RGyfytJSU7VXJ39rgl3pnSYPxA2mpKAlwoMyklNxSq30Jlr35X
zr7nX455eSWHL2QXA7iK1lvGCX7cBPtFsTj8xFY/Vi05NDo6mgn5/OVE6UDGMzj2aWc5iXbMcIlD
F3g7c5gmU06WUVrzL5tAkV0JV49cSxpoH0nB/1cSobI673qUBD7F8jzI64D1zRTv3OP6qKx0VOFL
/oL2SALXw4OG2ysEsaShMmhG+pissHjIwPq0mk9bshPtIlzWQhTj2F7s7sdmr85q+dgcFkUZG0N9
SqH4aRrhtK72FJeWiLqa8l8O/8RnCgESdX+HduGTgiDgIvHZlqhXvz7pGE+49DEgwxDExO+w4W2i
An0Ez4w6ALO23X+4+EMO+GzKskKjO6j79L1oHaR1bndAwqeAcLLXTI+Jy2WZIUPF0CnvzuRhy0Hs
EnOubjPxqE2osO+QLpjYKK/KX0M+YLuIDwwOY3dqfv6I2THiWmI6q8vJeYghE3yfyPsRcgzi67fK
bgnugpTxlP9klR73VBlFMFNpjJcHwT1S1LTcyWQAa+Ci5Q0t+72T8NtaXBFaaVugiwK1NBBMxKfJ
PMuqeC9IoP60XwZuHqUitXYXE3EmJFml6dUM8RNaj+ODHWEvBcjXUDmZ3UOR9h9C8/715Ccd1XDq
pRYvE8vnbT65UVnRrChJF4Z5A4+MbzroQ3oKOEk2TLj/xpao25XGhNxAa6+d51iTGOyNiIk23+nO
BSxVOKdRXPcXvku/RN8ykMc+5OOVdUdl+hu8PCHNLB38KyQaynLMPe464D2q0KWrU26M0SALjaL5
o/qmbU7oyP/tpZDmhIWr0lDwu6Q82T8lABdzLFm4+ZAN6jQU50fp3frprWVylDIfxz7CN54BShKm
AdJ7yDWkje9yFxo6NHBruRCQSX9EucvIUTgz/4lK+NmdgRLX7DdNycIjpfO8aWHMklXFJeX39lUj
EMzrSD++OZjXN5E5uJv0jHvoDP9j61wsMH2EhTkoEyGJaRYVAu6FTGBn75X9alWD10oHcOcHx83a
cQmJkH73fnXQY1U46Kx0Ox8JB0LyKAFPZMqNUT92sgO2NFmocxKDgJi3781vmOAGNTeJQhsJYQgu
fxwQlzDTgVkfoTuWX8fy6zI+UCbsqNpIL5Sg7txKRW2Fzc1HvkonWij51gQvdnhxEfNzqSTAvKnm
guzsBBeKaxAP+mhq0LDYMDnJFAVNucY9Zb1Hi6UwlLeqMPyFH6LsWX5pZsTUUbHjPhSZ+NI4DPnK
zrg3G+UUesoNMvB1ipaiU+uT0xLH/YReN5CnbXsUJaUmi4l0EAX4/+eLGQg9x9v8PPmLQm7e8jrt
OTjTgMFOEXszsS8FEYWDO5fznaG93t+UEqOZqVIwZA1GRIQ62jFiDbAm9q7JNGVG84sq0qkocgjF
mf7az6bPB1BmOlS/wxmlZcT84S9okXiH6PNq2t3H5vVxUkk8DHUIIvGtIo3Lx6ZXAe0gRl5wTU9O
oPaXhuc3WQx+e23DLLOA2Bqn171c1O2htHM2E0DdCJinieui83YMJ+r3QfKRlC3U7pXxu1SdhTet
gqy5NwyYTvv5VxlLTvZoG7rLOOdNShJsRVyQKqSzleRexgVIy7vmHxR9Zisx1jRDqAl8iWSYgj9M
AbR9HqcMAoAfy5iVSMjiDLXTvo//qSKqvnNcqTxwgSKSeKvv9rgzUBDxS/8gyGoh/lGEeK2d6Hw4
5I3EnS3Sh8hoz1znYmdOkslXrMJKJc15WRpBGbEcMwqwLXwCNTDXCx5Z7xb8LMK/5bMyV4zMZFYi
m9YTzsPHR7alPlqrLsgPlN0834A1apg6VsOZEfc4rsY55OXZ6GQuIWH01cAZKuoSHLXeFz8kEqGR
Yf1YP/efHaBixGy3jewB6ECGU0HYr7zE6Ic4GKWXWWjdTbuIGj/AJHz3tu2AvJIRfPY5XgsEFxzV
Nf4mHc12yc26xb5TQvuDCYU1i9vQDsgiGgFwnyh16wE+XbYl9kSAI0dxRnp9Mmnb0Ne73ddBE6no
Al/SthLgCY73/Toon4oz1+3S/O6zbKg4WhQxx2mY73oVKTH7Xmi8aIZdq2kIQ0W+hadmugXqYagA
c/NkUD/bk02TXKGG+WZoJSvDd/W7bgcV24ww0wkh1V1fchY8Ia6XGyFmTlgkO4fD5eb0pawqn4MV
hOgR1ti34l1ob/9olW10FFsnrGsOSFvL+KPt1ZhkPhW7gNWtynVIVdyDHKAVham6sAUZMYO3ymWG
/HFGD+s4aWzsSdBessaP/Ac85psKDSgZ04Xvexz/BAPlFMOpR2TrlqnV/OjQ1mX3bt0PsdJPPR2j
mT4jmQNKHXG6e1+mHX0yWDpKaapT3SQneTYTN7Dk+bzW/7qX4o1pLcUjhwVgoWxWsEoioz2k6Ujg
PVtHD5L8Z0gF9IsL09BdAEhzFaEwCEnDCe2QqrZ9/l94anvYrJkirCC78BzzL0TOJno+CuO+YISp
MtJ/KIXpHVZbEvEytMTOobWwl/ZfioFgWbqMWQRJxeskR6vZyAYEpA3pMCm7HLbxS1nRS7YFreC4
LkELjfY7Bqb7BIWFXhRNM+Sa9u8x3jM8nco2BBB3dO14BWd01dMJa2qVvGthjTNXy4xmvIKprE0p
Unbux8+6EZfVur8aguF0/1GWMU9dG5fKvl8bQZ511/CnYp903iEB/r8Ku/zl5lP5xqMB8jyHRQto
02D7JILtXzCgTFLXZaJQOVv7V9ULOs5EHQLQoFQzNJ0Ctqjj2diVX9eFHv26SiijlR3Y7tbiVKqW
+N2/KQ1keOTF2sKKq5qKy1xfSUWYXWq5x2JSkPSraRGwplgYsBq0PVQlo5A500GD3ZuTvVh07uGE
0wRUxpIc07Pe9jPF2PmzXgkG6ThKCTGzS+3h/h3pJBnnoKpvCCtwS9MCQowXtfGIBWPY7G5s7ITt
8nCVddydHFUIeplBA4KpChv2grFEVJM6IzdKruaYm5d53BRPgokK+FIu8/+wU6e76pnJlQ8ymNtU
MfCPMtqJjI+p8gC7szitRf1VJMnG8856pYj++eLepVLbODhqL6h9+gndExiKo+dq9mCw60la6ltR
CIzWRrnbZ0GPct+oXovhaJ2dz8qMTehvuYmP3yMPFs2bEetvdAN6xh6lIWrgazNWJSel3YP3tsIs
8Jnzbat0zcYojMwOOSAXBOGn2y9P/faUWqKGoO2UZWYau4Gaxf88hPKdbmkXyFLMYPx+USLDDxbs
fwo8Geeb8n2/Y3WAMZpiUBIg8M1E8ez2wqaLOmkXOfnTOgKBHG0uLuWHcsFgpA0aT8aaRNtX0P4O
e4g67eIwiYfXCUKIZpoQ4d2rBEKViMRinxiH5kR7+nZM25TjCKkUt9Sx8Jncyr/H6vussceJzJI9
z6d22zIjWvnz7bnYAggkqEeqa2mWCUz9GGsMaaW135ZWlyBkBqdfxA2RSd1vfrrPgVN0yKva+HlA
IgiekAq0SbXqS2UjPMKibbjcaGKrXd6d8uhnEAnhwKapDRfQlieFIzFFsfq9yWPNQZtXft7xCRUr
/AbavLb0SL2LjETKRw2uSWRazjOhzraHNcyyNvU1YbW/WJzt+bX+sa7xyQ85DwN7YUsCFBwcGejp
ez/QxBkU7lp3K/PueHL2x8aMT7S2SLS4TYpyKRIS9VerpJBvE1RKosPhn3/ENXHSGTQ7fnOCer0x
IORAzGi4xM5jKDTRANSeOWxO/HdN4aoiyfUABPCwuYKs6746KWbfROcLWLZTAhVB6VlrfXyr4E2t
SyaH01Gba9MpZ61v3j7TMC/9D51W172X5b10MRDwvBKWFzk6D7Cq5CSvHiNb+tjj63ydm3naZPPB
v9pNJaPrHBkGV1YHnOMtYUiH0FbDCs1lPPp2tsCQ5wrLBIqUtIlQsTOo05IW/pbFPknU843lEm95
khuTELUl6RP+FpVVrjqIqdKsWrM2g8BvMzZOuCdVK62dCX1E1PqVJ3RRqpX30XCtJBpUvSLC8sul
RE+FCJ7M/FqyQpeNwJJCTSUFO8JsrkHkO93/dwL0xskzJ/aTagJFTWioM2SYK0uERzqSp1+1OQsW
g9Lgc1016VdPAgHKWd5xD1Z6zqQ2HFLYmE56uXs32NfSZKVbAdYWXowxdcTkeVJI3M/QYsMUAJVM
Vxi6YVBG8hzB1YDZlgoAdvmRpALUkBIFTOI7zKz0bCjy0D6ux4JXiuNPUsU5Q33Qx10D20TF2biq
JnxRhw+Vr9GP7ELV2EpJC/+B40hudk3bjgwpiSf7dlhe/mCRVvedW9yOsZ0lC+qrksnXFI329a7V
P7DWaSJd6UJM/rKTHBFCtEJJI6jBDs+xaOhHXqR3L2v/i8fYruyWklM0p/GoqgMb5ahrzoMfhTIX
XA5A5lBsVDo1EPEE/+HOtRBOypK3ZMlT1PE9G0VFYO35rTiNdk99XPew8ahM+jbv3gJnMhsPbqyR
WWvMj2B1CAAvLBfgvQ8ZcSQvo4ObMZhfNYLOWHhZJtPqF/LyEXIe+EqAvEA86LnHtemtyd6BCcQP
ZkUhnFAnceilg+ZTCwPf3PpqpuNQryiegR9VVTiEV3ky2/2zgPVM3S9SFijRRjleLnBi4LWIUYY1
FYGRgxqR8yFkODxbxoh1md+3TAuAxoUvmKZgTpFQrtPttGCYG6OG1rqYdVVBFV27Hn4gAlNRNokZ
tf+WOLBquHBoO7di77Citc4gYGaSv41KihFtGIrMYhaycwAS9GuWaiEVKTcifoHk8zLGb8Oqoig4
RYnJ8TrRcu4c/KrZXn3PHwNP3uV49rwgrM+50chH3hryTFi4cGylHgESZc72FKMrj08h5iIbYOn/
5/BJg//vldvUiOsdpKi6BSR6UfscmKEZuNAlbknKQLXIVRxmVKHXnEqqfhKdxHME3ugTb5v7KluQ
JlnyF9n+fs8hjj5A3Nev5i2ExDuw91A3r1osdKvOilCJir5kPO+SLjf6wlJc38YH1qezKG+jl3/P
6VYanMwkcS89bfjlMzHP2ytyDv90G2cj6BOeEOqV7A3c1/caurWSOHu5pQEb4RbAZx66S5a2rstr
cWmttFrCFw9WSIXbxJbuanHsxEq9CLwO6ac9mzy9krsBbEws5w5XZm1dt0PdFplCMqBI2mrSoSRA
yePyOxbWRWYloicvUeRztRrY+6ttOwH0Vu3YdYETcSl3sQeYz7332suvZ0xwMfYnT3aj2WCKsIM+
X78Cwe4SnJPL8b9/8zG+PIAp/OqWfDZEOBB4Zoxxaeajaga8jc7fiVIf89oiLIyN0mnOQ2gY42iV
Q6RIQr+jq4ZJvNCnRBKvyVlBEgUspLrl1LL5ZZ2MEYa10TWx5Oigguc3XW9AXe3jsOUzowT8C/I4
kKjGgqHrAyurzlVh+wUiJ/7pGQeCxFeVlaEuMLKLcx3HDjP5S2O0JQDDPZuuc1bGF8635jcXKnXm
98Qmr02a3U6m5bDr/JGgzWRS9H4ot27GMAhOh73mofYThxS0NrhTvjCcavggb2plaBrp05MFFs/F
MebKayKNufstfSRJkzbW3pchJ6DJvY4N5BOe4hcLL7tZKpMqiIbm9twPH+l3HAHbzJ3SncHYFUSG
Vz5Ej3JBJ/aG5OmQojmS30o1AgzijOZyjvXLZNqo3PUcFBHCCWfn9qjoytP2yv7Osapm8L5FB0gc
e4+HWt042Y3BICZ/GftdXGGpxHJ/B1xEqWK5zy+MaRHTl2cPk53s3Jkb1/V8DcG/TYHh2SLJ6XIR
DhlOCUSdmSGvaUeJDAe/kmc5QPXPdq5qj3Fxc2Gc+lK+ZdZIZomfhkJZuRLDGLEYRUByYjaFol+9
THCFFg3yx3JHz9dycD6kwBdWmGJxaAjoyYohFG9WxTmXbQeA3IWkdiwIgrtCaSRZZXV2cnyAYquJ
VSM4PwV1rEWWeFKYUj5tJMs83Dl68NfRUZiOUKOgpSdXR8kXibLagC+CrspcD7cPp6oA8MvxvIgm
G/ljnI8jwpYkWRBUzgSOU+Ac1a19oY4pUJ1xOOg7BUl4V/MmYkNjBroX4fs7K5BSNQ2T+j4bFBUx
4RRbcqv0O2+mjtzvBcgJNvQAGXtyxZ/sX1VTRDmnAPhLCYSpr7NeT71q4328llbKD83Sm7PgxLyD
eWo2misQ9PaO8d9oAi1C22PPrC1Tj2k+bHGueCG1rMzMmdE5IreL084icr4ToIfal4E88VuzVUV/
EaFZVcY/ZvSvTyKJDF3PExxMP3VaRWp8bc8SB//edbYAKZaJbmoDGcwXw+06cfS6gg2xuJCb+Iz5
6QxpH45TqivOAV8M04BHA9D7Hm0neUiZXdNxbT6VXqXTa0A4qEX4tDMbIu3+j6qtKiH8LSOWfsMC
O6T4ztrsVR2NSyBOJVip4545s64TsihhzbYykxP8b0f7EzTDxjJaR7cLAGwymMyNHupm46NgzrrN
HeaFK9cqWL054gDR1QRocTbHQNS/ziXMR1794OkxG6ltdCPJ0FCNDJJ3AyOZMIUxAraaW+RFwuph
jg6e7RlQOEfo5c2YZlZXtB03opna9UhxbLw1cmgq2VkCVzrelj4KhODBRmhnBFREXXrEIxjxk/6E
zeKBFfct+kk0U/AcOfrtYTxUxiaVc+XUJaH8QZzOZqUNV1ye3LJYZhIPRBmnFQgQ+BnFatPmQH1z
pcLVAoR+xnkCfVCoGOeM8FAgc1ecIjCAuuR4NxIgB/xY3dWzesZnOkKaBuPVK/Thjr3T3fVx7OD4
zDq/Q7puW4rVzX3Qs+eqj6xa3IsiGGfhhkz6ZWnu1lqJzGQX4mETS/47TB03IXNEWk2GIEbs5LzF
enxE+/ICnjcsEnFA5RJBKPQc9LP4rQfV/JREm6tOGA0iJqR18njHPsbZsGV/yqv2ojGXIx+vTt1T
XkBOszpLeZhapU0cQQIucbHkIqqRLwe0zZJM13pBu0GARlBXhmPfwbC4MARTa8U8b/arWBIAmoP9
jXrNgzs3oDpltCnMTnj5AjniZGTs9G6V/YSvYsv1FGR3Fn5EiFIKF1XxORmIJRDWkUWqpBJI5bRQ
QnEfbKGKDfSRuwanlGAc+G8zO72FeBOLGiMXkjPd8KxPlFOPDBDPrYNd8yYr3DZ7HWCuTFEyhWt1
BKJ6/vSCAftjRNAUacuoVf7IeeM349nJmDPyeyzbJaHn9VoV1e77HkFUMYTfZxzhhu3pQ6J72fIT
PHKfg8rsIsjtD5tNTZuoaLLZEvxfSuQrLEcJZu7Dq42mFHw89p6BXKrIMNRWrDo70H/i14HoWjvR
mTptqW38yPow1Sa+LwLHL1pDHjRBOjGhBYBoxynsTW3nI0cQ3GU2eI9MT5BmBa1SBKHcjPovj/Oa
kCtaYDhXeSWsClcCm2d/OcZb7ds24HckSUkNfsmO0eAS/jsnPrAjWCdUagO/7Qy8PyGRopEqndzS
XxTL5Z3rmSQJcJp5NoqN28oEFmOtMCZhA65X1sDtRQLVn81Exi4SRIbaQbXhP8qenTtuKER+axbd
Tv3jk45k6YPNcYnSqSIQrWQ8ly5XIpVN1OtCBeFzDBU5/KK6D9yNrCAnWKiFXD7lqcsi6C1YWmZf
fBTxFise9P2n5xy2Ng2G43Do6IluQd1WlEOeRyTQwl9EMNU1kM0UZSEJ/BhqsBvU0aqUcIM3Lcc1
hcmOp9ET+cmShlGrbBuIyltUFJ+u7Rsk5d76TtFH4pRuAwJFpMOYnlhTfUBgpkSAurJue3Pvqvcw
RmSZ75FxhANFU54z1YVhVKV8hgrS9Gl/aJO6ZPeLlybvPCzqvGjVyUvtsKjdHmEnmItjZpuLZm7y
d7bqcOkbMZXjT1STqdYnIdDcJUx3FCy4+qGrj4BbSh9v6er8ac/cARIHpRVqWSQtKRknkJvYbNqr
kc3LVIAtaJcdKhT93e1j+QNnFIfImjP21Cl+KGjpP850hnHghXPtChQj8Ellgevyyml8gNPfKz48
C+oTCQkX0KEgvfWLMXtZhcQ346YrRACKYUtxI4MKKr0VRENck6xZHYC+CNmmctHURayYbG+X0Dpo
j0BdLQI0aYIL3zKgbeHGw5yRkbg6lJgqW0ktBt7YdBXDcaleotEXez+jt0x8KLaKd3oH93CIzG1J
DHnMdQr8cjqEnc9qVoEW1xGPse63e/IIxIft5oVdLvtxJENJbPSgyFYT3SMGpIgOI4AoNJ3QIdPl
IN2RC/hiyNCEIBYhsg/sgDJ7h1L6aBGUUTNoPmiX4kT3u80+f6dbbBsI9TlaC5yB3W/DNI3efj+W
4o8NwBOckBfQALFt2QT7p7p/LDyFoJPgqtLW74P7XX2sFwsZeXKPUnw5mr5YQnN8/68PlQJOYP/F
/aSHh6EWtQICyq1eMk8tOMYlXfbSMHW69riStBiE3lha8fn5t63YEuUEnRGEv+IV2anDWtJMy+r7
FAeyIL7lUMa2thLj01yejSq+Reh3m3egsZiBcIffnbX/2alSyWfSjOggozwMSIzoT/eXDUBXxX7V
qNIAs+vdauL2N06n0/qs2GCAkE7pU0KD7+MGuHydryAERD3cHaVoDwQXYVX271UqhJH1jgu6X7Zx
tQGCeDVS8gcNuTYVztOX8qTfWQUoGWU5DtNQU4z642qVEcIKE4TKoaicXcpw03ZPI0pvQjm0IUWd
WlD1z/Nsco8ygAJAClYs9gU5CyaoEu/VaD7OacukJhQjSIwDW8Kr3M0hzjqKHf1EtTlrPHqy+pEK
aKEnqO+ZH6BMzrc+S/Unecrls6zz9NlV8OKZIEMzqWAGraOJJnTBMLD2OChbZnAPWuY4rBE4tU6H
9CBaHQ2gmpJY1UTCdkaQ/8NRJignmV7mzAqKrhlbrOz9IH2oN4e5MB/FKdbOOrHK2I9vdoXuRw7S
fMkMFj9wicrJP/ZcpDaZ5ftX1Qtm8hkjzn4Aiu2mI7Dv39qWFCbo1FrJLeqmmZFNDztaEjQGIqHP
/tUEWA/PZQTOkW96aL3X1p+C1XiDDI04euhbgyKrj38itRZB64fd9rkbCo4fLkTAUcQFYqTerTnM
ywAdnrMgBy2/3lHbP+NUg4NIkh8PlV/RbGexuNxw71YHJdMTPVxlwb5BKEvyl2JodqNYr1x8wykI
4C7XmX7kH3ydxgso130J5E72gTKVK/ourQY8FJh0MzQ5gHHa7KOuMaIlMGuH6kIbVpYi4XDvDTU/
j1A68nvS3F+Rz2hl8LxDfxqBRVFJDDR9G912xqA39L6Clk8euy4pXx7ZWk10NPBAAn209Ct7pwI8
OCyozA8eOv6GdRWsXxvjYlyt8RDDp6bgh3iPdNw+RR0zQOCiOlEUsDdLdj1yjF+dFroFc26ZXqM8
t0YqzMlXytMAdrulXf+WImrhLtPsjJp6dEB+sMixigNq04m0YIjGDCPdSHpbJXbLVH9A63URTJLO
uqzy8uKp5Y1stfaQxU+GaqGibbTxDEdkoEMp6rFEx7mhPzwWMmVc9sU7q9JnczX2xaCRKgWJiNCS
wNQtqs/SDy73ToXvjZiI16yUGXSKurnQL9CnELKp3WdQx7h62c2yw9Aib8rbT6s6tT2DlLED9PXT
zOvW5gDEsgT+RKo1HO6apiqiCreWHQKbdqosHV8eM12SW4w2kgS1vHXj42mGJBINj7x0Cqf2jw02
uNQZq5hDlGnJwJF0rn/ZCQbHNvilxMWs4DdniAEx3itU5ZklIifHA7GPxBfSuQuDKmUnYhuNS+Xr
oQdP1Upwl21eEDtXhrjIytWatWN385Hq3am1cLjFXilrV8PgwTMvL23k3nwdY5+p5g/+4da7sj0s
jQZq4jvGWAq5tpStrs9xFn5dP4yBhPAxlQ4blsTbLH/+MqRw1l0GqKIDk2Orp0jhOrgEvrFa5IKp
0dT4DRLN4X4uHOTbJ4036L7kFG/IPgdhIEGcHBDRsianPaaxkBLXrlCqrnszSuYuk8jD1XgQk7LF
ly+MY47o0Zafyi/5aiouosERbRLugAWPDMV2tK1h1EYTe39uFXeUvb8KRgeFMajdlogcnhEl5o6a
ncu9FPAYXd4230CyUI85wFPRIP/AoJyBDcVdZuZ8OFmjta96UXGtoX5oxHy7Bb6JcCohSSBg4itz
roPs6aTa5qQqWjMZ5/Pyg+yTz58NnRzdvXNWWBSthmOM0kYeLLxbiBRXo0MQbdMOvYlYPXV5Lde4
476DV41C7uKc839su7bISngNKaNNSIucb/Dp3RR4RxabMdCEYbJEKe0BY+lAy+B5En93dwzeyXbB
nqWpOkNxpg78g9VHUot9SlGo5e8nXixG0Gx3yRpslBGuMs56pa1g6xzIAiC60uVqDZ+9JuniKbUj
ChAYCkxaDMJ1sxKL2l9MhvvSX5dVxK1GS7IxgVaquI8biOpNeNOZpD2MkBx8zCoJC3KwpYta6J1B
ZhuEYB74ke1JxSEZZsbM0VbC9yek+sViOH0m0ZqdebliscNh9erJgXB3XbDDK8YDrNsai2LQPXgO
HM5wUjeQk8fWSVJMua1QpP7B0Y0BGqh6kF146y0bRqLf3kccd4XiJqwzTKRpFOZtKNWl6vYQpDgv
icZAt4Fx3S/xWWi80MbA2sDkpFPfpK9Z+D3k+2YMtJ84kUhb8Jy2k/LA2EkerHdSRRIq/Co1371b
YA/0SmXrT6oshGFojiGSPEyOqlWaeh+mwW+scIURk4o6lmh0XlJo3oe/2m9y0k26hDxgB25cAMLx
7LdkKB27yUE4vodUPIGCSqJySP5rq3SjA7UADez+7jwF69U3GcsSArJvqjjyJu1jtmlFCNYYZ9h9
14UJv5OgJkDu3wB09e7wto9FzKGkBCoyBZqqde4F1pETZaFh+8ndgH7StWFCxyIXVUYTwfe9kQMg
9Z86UcMKaSj2zpDP336KhbaEvrl/uMov8f8HrMrFDmXDcRkTLdu3FNG7idKgEK91r0u6dZd6DZH/
2y1GnNRZnc+YR9Nl48dM3fIoi1Ed3kyyUmQWi9DFr13jZJqmVbejmWD2hXCEz1MnKA8zsuXdyqju
rrh50V/RMeYOU/w3oIXatG+qDUD3/R89fcNHaAloPH66UlhH4O0wh8V+qkAOPT2nTSy8gwa/cYhq
67IVZ5HMYs3o+cy7ld1leFGiJqwCGS0Pnb2c6GOH765iXPvSCsUOttLHPSrIirbaIOTQ/DwH7B0p
XcUIf+w6kGrEI+OeDHbiREwJaRoimd7Pd5BILLyAlXDSkZYbxelVFHKZ4ZXXl65/UrtCmW9EPJlq
vM+2KVmC9DDUJLiVgF65jXVdbIQatgSo5gxENaBWK5fe//qsWXtiEkxmRyW27FAXS0cr69J01PEI
GOlHQT/DGSWDDu6flsmYDVwxCPpwUbuqOu8VMuoy4aPfF/fCRPF0px8jVuVDg0p7BzFsmtQHgsI+
nhXn8roAU6IUcBIwiZDwF2cQYppnf1qHiQ6teclkOct28mrv2yMPVvaGF9Yev2HJTecTjiZ1K4+z
6evPHm96GS+CZTQojyvQBge08irde06E031OKnkMCTEyIBOs167hmvKOFjdsnTJIIwXFqDsPBSrV
CeMlvM8y7LKRyO3Eamj4DoHWwXRMCvMvv4nJzN9GH/T0HiLJy3ygmcmiRJNk6OCph/6aCffvW9X/
K/jX7VyM1uL0tuAaJHKYWZGXeaF/9qIZpQPXbk8MGLaUjDtHaxjOGht+YlZhqzk1NX1W7/oDwaqQ
wAcM9I3qykYz6+CWybrgCrvTNZAGIDthE/VfiLbcx/6XCxpYIMEE0yID1/3P/EXZSHL+9raJCj7a
0wJlStIuTtocPiFRWCbU1XfAfsC8z3YU5+Vi1CXESgzXZvJklruOZBgXHbW9PkBdsu7Oyrx33jjd
rtABUfQKZV9Ku6MyTUPJrWWXrm2QnC2VIydVnveLjKl6EfByfTHWklXHk0+uJ3Ucaw/vYhhjq6tz
go1ZiJ7KSdpW7xn3kZsHFUH8OxIWCwzazo5tafpraNMpQU8jXshjsg/Fw+Grmwtq+VOd66N24GYj
hrp2xPDjQBYRriHICyRRrH1005Yee7gZRlBu0DwRvDodJYmRxOFA0huC/xY5LdDnt4lxQz15mXOP
Y2j7iY09ZTPazipNOEZ9N0VLo7muw16Zw7P4QCfdOLF2r98Sut9PeeMzYTgu/DMbL9dNiUiMc9nc
6GdOof5FBe2UxeLIJMKcYvwguAzvLZCXi15hWAz674liIFKRxKoNz+g/GerBTlkbGiDkLTtqTMW0
6xXCVotDZku42T6Ibc3uB7bXynizoQYOJLshP77vUMjwL2ZUQrxq3xx95+qHEA9ShaPYc5jirFAX
h8JhruYkEBU0TC8E/r02si6KLCmdfdtXHk2fjShRH/2YjzAbiD+cE5UH6Jp+Whl2lKlmCYqmyI/M
c7cXeYVaKrOt4aKxW6IboerdBhGFLVOvzvSdt0LVsqDR36NNT6YqIIYh1rHjAoRZ8+sVVA8YzO5O
caYQTkofz1YiQDTNHm5wwEULGn1b6ct+L7NL5pcFRYVVl3ophidBO7P8pdTsloNFQzsbc/OUHx8h
M5vGZLvX1ITqsg20LxcvfHq8v2aW7n7gmh1dWgu7hGuphc4heTvNROcnw8lkG+ij3y8HcNebdcE0
6LSzzmKxlX2xi0HubuKuSBSDPOMfOZ7klFe91EOTa9DFHLOVtc2by0gFlVFLXC9btApLmYhmtEmb
2udAv338W7ygZjH2kp9EZN7zvJDRv+4bMKCA/vDo/FLZOLw04prN3wCVc2Kk529ttubJwyuJdH8K
QXRsXfBsCP40obI2b+O4HEX3hPc2p/4NJhT0vj5dl3ihxo01Usp5WMtspj4ENg8HMiyYvJA0NGgZ
YiCXU34OJn+FPntoW70St16J4k40rH3eNhXtXZfxqZqAzThXJY8qU9GkwHWkQlAU3pMCQgvELy/e
CQhJSFB09MGVKhRLCnNwVYppjeD6rx9UU81DgRza+uA75YCJkdyc8/M8Z9A/gA/mj6rt4dioNYnU
IdPd28TjFzpxoJhw59fbhDZt4uMAsH1nlnoDdoH7TNUhlbV4IYxtSO53ALAwCXKLeKDjm7HWjyAx
vhWiWht6kGBlNTZ+AactgpXLcHfE4fAEwBFyAOkGKR6RYshaDSBto4vNct4biY488bjZsXLf8O22
XP0Luon63nL2flUBuXPZ5K4Mu6SUdYn4WijbGFM2tSXIWaYV3aT2/Q92iAoqbip2MAeOQby406fx
RF3StWWBS2lnxJfMFC5KTv+IEMv70JYTqaPR/51b46ma0Bf+ubpWPr+LT/TWdU/2Yuonbv3eBfrz
HiZ+5soiY3ZU/+e72E8PhqqWR+t9EPJtIppivNPHD+2WCUyYIJy3ofHgcq/PK+gQpOQ1Fq6BmUen
4JoJ4dKFwPU6T3Ej2lb/WO+UAkOnZo185JCRsD0P34nzxiSDfHyejdJx7j36eI+Kc9KE15+cguEg
iGkAsvfIjXIUCW4u/P6fx/HycpDkSplD8jQOexuPVJs9JH5hR3jD2WLW2VuNv0+34Ek2gXb5urO5
6qHRrYhAYPSLxRryNYP7CAhIw6TRr2ANCXtLN0/itiVkyXpYNUOB96srkehvjA0GtPPW6E5CvZkh
0j87XUmIIbMb70yAQbrlO9T43fhFL4P8Ov50GDrZTBqPvuIC6/Do/pw7ZQRGyW3nfxZzCkBP+kBM
Hqd5tbGytoRXoQc+dCfJjEIXOuke6VGTYr9j4mQc6IkEBRUvpY3WJmMVg09TTgtUqYET23iSW9ri
FCcJdRYS7K4Gu5J2fhXVRW9OUOw2j82Rlb4obMHm81CD1wm7tdmi3gj+imQMXzBxy1w8Kn67DAta
wCMUnXCyLUIM3LqQ/7NwxywlShab0i8Xu40kaXXGdW4PC9Z0FWvm5+65n6rW7Bf5shXK5yKp8eO2
1RwkCC/shmCg7THLx6T4/xKBg2HnZla+yMLMeD21T81e7yUQ/EFcU/kWDZINeSky0av32uSLMLE/
sm/9AtWqoNQtHBxduzsnVVXGLN/BVhWIurz0D1vgwWxDFh2UvUua1P9XxUtZLw6ywIMVlnVE7MDw
MSYeIIV+pMOLqsKMtMvj+j6U7zkC52E7e+pet6x/JyAgq/hjKS4Y69d8tjKhTky+oVhZBXNBUGdw
l0sCzwEgttJTaXRn5sxPzDJKW6mUhSK0Y1K2L30rA2YuMzhYC1/veMs1wPLM+fOCnmhwsCyjJNZt
XStS9RMrEEaw9JVE87WhIyXzmIoXZUAxPV09/yUJXtd0OpZ422fq5tbpft1ADfR3dIC5trfgDqz7
rRZcOpQ91nHo3TKrZ5sHmGETLYH5eBcQQBUs/UPSz5VpqC67jqoz56sOOJOKRR5PnfWalpLs3rIK
zNtoVObsWUXPwgziQ4yWKW4ZWYVVXMdRq09frzZ9mxpGss5qqqVEmbtqm7URpL+Q6C2t8ZteDe7q
Cv8+Ok63Y9aJi52LWDQ31oITWgbMezK2OPKmHGDMLVqkMw4uGb2ldFDKgrFxiMViujf0wfO2rmmM
KICr2Xqmqm4IMERqJOSt9qgen0RLhq2doW/4ABStFnP1EpTLADAGcz+i1RyWTF7TNCdERKdBIV2z
6u2RFqpmncgZFmgDv1+AUAeIl+z5iZjqu4KlDewdX8AqZyeBhhkhV5PoniOtsbFShOk0YUbGmKn/
5i7u3WDjQRzJWDb8+CjTVwJhaZFZsxoo2/PYj554catZSJ/seBP7FIeCAeq7Wf3DWmSg8Yw2bwdz
KUOHHsEIuI2/RcWMFrgslQ+MFATaZYqJr4SDwie8CbOJGlGftumWT6GKlpXBy/YnCA3xvsMC8ytb
CLdRryxmrII/L/GLQFSB1ukvjjYa8M8LViNdJoh+OVzYYALFxEjE21chYAbh37qM7/8HTWeUsKad
u2oS/hj0Kkm08QvmeWgYzmz1SMR5EhZIGUoRal2jaEqtMBYd7SxxT9h0tOI4sUVUto9CGaEjIv6h
rSXkIdRqsoV277eHg67yI4np9hTlsV9RlEnm1S15RUlyw+eBzMMx7xnY+LZ4lNjCztN7Rr5xF+qT
YV0AZFDZLL1yqOlWX0WxG1FkRAyBYUR59dICZAqe2E947PTV2VS+b67ej8vQU8+fHHRHrxzAZHJi
qpVvh94JINcKdZ2BwldCManNoTmfUq9C6wUcZs3BAzppeV4JvgokbEEM2kFv1hWKB/gOLXuxAwoR
DUeoUhnPOI+3sCg9aGaYpvRNGdJ9gK8QhS+SHwaeTE32xkcv6BGcJSHjpnCSmU5j4qEDceMqwwVH
kLlCwsmXhr3KZcsGCPgjmgw3cOel2IbojDTvhlIHghecQzILATJQw3K4x2UfYaJ9bQfnWbxqEDKu
IXjHQIQMsanHPTnFcokojtidMdhV1Xw+8YsRgErG9nM6dsMo1CGWLHPrQrMhDijnYZlbWGPW4vy9
1W4Pn/J+TooSkbo7S8ltk4XiEpyEj22oSeb6R9FTIzyGc1B7LDox+zk/jqUcPytQzGcS7/sn3klg
KRgDLxe0R7PLiTHsJzwfI4gV815EjEdxO4GYOfESqO7WMMiIPcBnolRWFiWnxFiULZrfL6e2paXI
s9nvbI12UyOUAwiYD3ayFj6UjTjX/CfV2OiknqwaKk1P1gub/mdBqmPflU/X/QTP07Nltu3RBtD/
1Eg1Flnug3yOQBI7ZtTjjMfkwXmaHJJL5zf6yM+hkqpx3gy1bWoalZJOu/+p3y9VjaymsVdO9Kw1
67wMudQB7gi0N+/KFH4qMCecEsvTfCVKblfYlIj0gZE4V1qX2MpIjoDmwC34xMkb7AKqlKleoB8w
sgsFckIWRuMSDEwP+gKJ7qTERrjXz+Pl8P9dh/gbFR6iVTTtCLHX+iGTIp/Hz8myBX8h9G2KfzTx
ecEm4ozULdqXYQsudrcjl+qGlcdG1AIbHXJl7+uLniCTEtAsBVqZHn7/hyL8jL7leFHSd3cJVoAV
WvCykuM86OwpUWKtQoXNO2KLfW97RS3MowwU886bM5tSAGSHmX86nQlCi6pZ0+8VXCiQX2pNkhdF
HCn5mNfFsY6cF7rB66FLSyEJ363KrcbkrqvSfq3hUxxoa79F8udr4ty/0gbHvPrOpA9BXVW/hrbD
5bZ5Q4jo3hBURS7NXqTn+HABVWBKBrWS+WYDJgN8sijlbFiRrqqdMmf/sNm8PxLHL97enB/DKRGR
N1i9TEmNmp+TKuUhom/Wd+O4o3a0Wk+DyqESe5oMjyhFAMqVtrmeKMny3uTrURoRVauUY8YL/QCq
JmWKS/w7FXsWLIHfPAQoA+/M0HSJOnmgFQ3aUXRW5GKljAYPrc3f86nDbgwkQnqGAq/bX/UToigZ
Xr8U5ZoMUWuR7ze/tevToUv3wMoWv1EXyDoK2F0ETiY868y+oWi37U7v8fgRqZUbOxWZa/4JOwue
/Ydg8/CDti8Vo9DTPcwfwksXuLXZtx9YokVDQEBdITb8fvvMq/YDuZrGSCO7/iwT8SbyDJzWWOgt
mN46L9HtZ8NqksFWYWD0L20MdQc8iZyqlZ7NQM5Dd95f98WjZmpDzTLmsg2nIdFLBzODmVqJkiDK
ghrSilvH5VZ7Zy0R3lmmkgvDXd9IMBRD3swwBlYKzmP4eiRfO7SNnl7n1zs8s5WPQB4bmiR9kQIE
SbQ+jfljG3QOxwln6EjsYL1gLaVq54PrNREbT+A98T64WCckc0voAvqbDRwsf+1AftWsQVdwg1ZO
bwqa+AYHqQp9NLo1STRaMo22zcsP2x90tlXjkZtK7ZLwaonjgOmUKWm4hrlQzvayu/B9SfMFBw8B
bPemyiVUbkdwqmP3BacAvwwTnSNWXEy/thZhgxJS0szb9kyRu2cbECBesHD3UaCjjsgPjlzUwUUA
+6AI93NGCTwwyz3ETew1sHtOWHOV1rDKIHH4NF4dLM/tRv5bPVaZIdanmQsXnFsz372k4AyyUCXp
QB36OqqCZFg/dBe49aFI/Rq7BOxZff8rnQRoc4+ja0RYvMxX+tKUi6KW2eta5pJDj69SDhoYoNUi
lFyEUwRz66FDwq2LqKIn8ceZQRmAb8y3Kl8OSzfM0yws7hQqCpMv88eSFY8KOPtMMxoaPrPAL+fW
HL2bd2a2HMfPPE9/oUIyyji5Q9hQYOiYnBwLEel0Xq5YV/dC+orJ9NQyp+1qtwHLV/utPRbmyZQX
j/JYnH5OwKOa7G1d7qdY3e7o7UQmJVDkcx/vdigeopSzXVU5U/Xordjn60vLfzsD0wVvM+1Mpbb8
Ts8pBKbCum7zghN5Tz4Te+nUSW8207qD9okem2nei3ip0VHNiTyy/eITQznw420bQctYDStSCSIG
pDzdWHSu6afa8WLa01HECqEx/MibikREW9H9rKiFAVNJDh1Wp92U/+l/JCMP0xF49WKYv9vz0/kq
OsHnoeoPWIMeOir/Hpw2T1gzUxm4wkhCyK3ozggggjJqgLUK5InxzG/6Gz5Bc0or+8O65AcjfURY
IPlF33OUZb2T5Gyqrq93WM2AeeYs98ewwZIZ8NP9ollQUb98XN006U9y9z0HlP4b6vxuR+sZHRfQ
OvO+aEMkchQDKfNFmN58Bn9IyPSdIXutN8ke0XW/+YCd8LkSxJYfOiqtp0qY4DaI0VzcmqTnEJau
g7MrkKlUy0hEqIuOO3xP6OE/Lls0R9fEmbeE0n8dhRlHDR9BSg4Fx2W9xWHkgPajJIIa9/vX1P4n
eDWJfGYPODDaj3kdKy7jNBFtpwuQPYFN4U0ceq9SRS6BrDeFWD5VCh273s09BXZdk0bqf8g2f1cZ
B4n+4ffckbqMcGBz9w0NlaCIx5lZioJPOSPlBQr31OxHQ6LHMwVTSb4jAOj7/3Pn5INirqvi9Glk
4lPR+GBv7NOuWBs7RwZea+jYMgRTDaw5WxdFH62yu4/eyxGmu9p9IuWhmep235ivEEcbdssGif4g
1sPMfg/6EEzyVMgPY+pQhHVJVqaDJjZp9vnXfI0WN+gTa8PUkSnsf0j3EMErP6E6MdAUjfAXhZdC
ca3WEJ19mqeDkGJ8nEOGSJeXrAOeQgq5aQjsU5Jx+anRe/QUntr07LF/nRyAl7P0TtvizUYbgQFl
Mf+geCNEbdG3bAYoFrHM08iETW17zuTxuaOVY5Mdtnmze0cDcPB48guW52JQNsTlGxhFJee7mpwF
AL7lG2NE37fF3kyev01ELdOBMlQYkkl5xR120ztyzuhcAp5e86+n4Hq3eujFAGGbixRcnwAi78/M
ncnkvkJPVX+1j7Y6U0FjI9Xh9R3z9gTRiKHtU8VrAsQ0Ts2kKy0vZwNDEvUtypAL42Bog7Xzd10G
TV4yuH4EDa9RSdXKFyBSfpiMurLhI+UBULwKmQEwNCyD77PxXSK0Z9OZy5SeJncEkez8d9oRASyv
4fs8Rya756OpEhYAdXx65myqE/jaFqtO2NJUOEfrUZwh0plmZjn98Io4ZqiPgfKCLwKaZGsY4/aj
auAGdYtlXMLcU+kFTe1Zycnge1E/bcctzQoV2We6nvlL+j7BiVQQ9UXI5E7RLTUH3qEIDzb2dmXg
MsUpI3Qb0kqtMfnPjg0MeThTavVRCBtBi3vWs2ZqDB2Dmz7HUPDnuFE5eHU+1p8bv4Q1GRmsxHSZ
GKEI33euOw5tnyGl86QTfolLgP2YTtSqXjyq6cbsZ/VMRiXm/p3nHsYbT8E3sbaEmcH1odAAebTi
2wbc5La5ShvZesSGlUiw4GeVvBuXm7AgPzIkgGJNK0Xu228nOBLEqD2EU4yvZqjRNVROGRmJZ+5W
oNoZJZJ8EbPeYOLVm92+vsc+I80VtO1GpmYH7PsrMJP9JjMopfKJXBLa+Nrcic//KGXft+h7Podn
iQcKHqqeCAReRf+oLOJOqT5OsdLVY0guNBSUhFllX57nRgge5/uomTooEpgLwVySEIh0lD3vvLIn
8m3PQM0HAzMNWQRhZgUo7LPNbIpfgUJz++WGtFrjPhgszPcOGB65i/BLZtAr6ZPPNAMFi02y0rG9
GDNOYBwWvek2ZejIv0y5gwWz2GdhwkHvQa2GmXmldi/IATmB5dI9jwgGscWKcojDyebRIxMgeFsA
OgmK786QEbt6u5AAHEVPKlqFxHdaNFWjcJRRDEdo2koZ3HJ9Tz04gVQGlCIATQyhoClr9MIAfYpQ
Vx4g6lifVd4RC69LkYupWwvoOqVAHVoavgLPmWvnxM+Bqq0ftPqiTGp6n1lLpdO/ckZiufn4cWgs
M+xooZUGuDpJXJEm3lJCIgTv0H6Cs7OtOkOKpI6FM95HDOk6LVLKMPqoIpPYJ+TniStjpw156R97
sxGarZbGGpObYOi2g/OzT8xvsX8YgwIQT19L6M3UncR9my7U9vIdMWd7wr6G+5z4qQCSViaA3ntI
QKr7Z/xJy0L1+rydIp4XcsW8PRxJ0ZzreI2gVUqLo0LEWzaOZWhJBgDInnLe9PbqI3WUCRxC3JVh
f+4ieu4EqMPFx9SgQzwAwJPOc3kJ5T0zQLwtQbQtGiQxQFRnEodaINxk/9HDWjXfay5JGAOi6WOo
kUeEnoqdYXfNeJDv6tgu6mCFHTtgLeM1qgPwU7XjYtPoJhg0UFP2ogCbVQWwp313cAUP+yNJxfus
qzKMAFbzvHX03ucbelZ1WXKL5jTMLRxS1TiOESepeYcczDov2uJF83Po9KL9TjIMrCX9nn3MGgXS
dnVyX81H/BMAvUk32S9DDKxTvS4u2ZTsdUG0XmjM4JWftgFcjTFuasyDB1USSeq3G9Ls7OaIePmv
aW5F27JOzohvJ9H285THxAjBbbj4kEmWca/CKIiDPIDUmbkwT7DqxLrR+W3+PST2wo5Qu6gc9K+T
re5BUBSQUiIkgXhZ1x/l0ltmtoexF771sakkmnTUsq1xENbyFd456YjW0DJwfzAjw/cXI1frTu37
DfjOq6pbApPoHemOEvDJSHiBsXFv1BG7pAwSr8naf6R0aeORi/0LAaoVbKOih2c1eBPGQgsboWuS
HV2Nu1FfLGYVCfRadhclhaeyBiK1nxJ5g35WiBxjO0PsbqwTzkgUvla6waj345wJNMg3FzYvU+pC
nTX8AMCyJp6wbv0XwkxesYc2dcvMRKGRw1S3bSQpes8J+PNwSCjzQolTzT+f37ZSM9/R2A1cO7y8
Vf7Nrr3ernffYtPuG8TjkcCibJESZS/Z+A5qKeqFWY7J3Jh5ka+jEPLjy45/qvhgRp9nly1KWrc+
V0VguiYp+m1hIDuD/ZEzb7ebPNVjJyq/BX2TZVKz4ZoQufR4OU+sFfs1ThCoP7mIZys6D//vDvIh
uvQ+VRbujn5XLv2PVPYzsmgBlfu1N2IFukrGkDitt1ZrQb/fAIOL18yQnlEtnx9lCIDvibODIYg3
EvnxjvlODdu+TQT+4FuiOlIgwfLKoAM2jAbifamSgvnRFoXsEXanm1Zf7hArW9rgxtJQUWGCUZoy
BZtqjR1pdJFBKO5Ns5DHpANNTKlhM62tjEOV76UP1u3b1pHg2bBi4FDCMJrbLP7+oBpYItLN2Z+U
dRsqrkvfylOJUZMswS9ubRMADI8+EJkvQI5ijZn/k6c50s//zP30fosEZPhwMpIMNLuJYvayax0f
q3MgrpDqNOb+mSr+rxM1UEO95SmRg9IREMBdQdzGu2yXcOmockxhoauOw1vRgVhIUz/pnuEwC8Iu
0bEQpz6vp36U3KQT5GfuGRoQN+j0yolgNJ7EgtAc7PX4jgsi20kenHWvdB46PHVUTcqqIIbstaW2
KVNJgYm+B+vf8J6TwQP9At8CuGS19zz7IU929i2gm4CtM2spGD9finNgjAi9X+I3IRtyKDBU/sxu
ddY7suyRly8DptLa99gPjcKBdU1aXelBjLg3TqJcssowsWOPF/1PYCJe/mGpovYpTZ+2rk4XwdoF
81EfqKzgOTCWewnQbDWMm8tsMr8ubSms9T1xnqUhOL38PgIiAlrvMgH5uNtBKG0zGYU7zD4ncYRl
t47+iAi52T7JqiEHuK2TnooL+yQeSyWSEXZwoE4PX6TIOUzHGnzJJzMTr9GXfSXrIVd5x9BxED/+
TUKwhVehztHzfOX2ICbtTjixopH1RKmeuYEREjMudQO6n8xloz2yCoixiZXN3Vgw9Ph92175X6F5
DZ+e4CmQ795pQe3wg6eDOmjFNEVnx8F3XrQIMxYQ4r1vhENNvc7yUqb1+KoajReoMQk34jdkwff0
vti/RNLJzls35ECFFTikhv2ZxDosuGun/IN7Pv6rqcpeDe4lDxFGnumqe3BN99VW4SS6BvNwZbgQ
z6FDGzUJQNz7rdUFqo4um3gObJ/QKNVmLUEgdg7Kz/6pLoZmummO/Rl3AsF0pjzvBYTNsBsafADD
yUFtfi1D3SpOK3rSbwWeYEU7z6/Nu8JWu4t/UC9clPgsqbx5YUdx7XyQmr/+Keo9Yx2tw9w8rxy3
/GWgT8EItXBUU4WsyAUbLTmrKQu2kT7pvCfjNOmxwIws7HEbpTQBjzUg/R+jQcgFbknU21RvSA+o
ylmLetISlFP4CCVLAL/1uh6xypwTtk+oERzthavHNHlWH4RNTB+ilDRtj4ZlrWf+IRlOsNKgdp1e
zBuEVFDSoI2qgrizvyGZeqTlByz1P6UpkNa87Us3pao88QTwCgUI80oL7NMfV3ga4nIIzYuZA/A1
flhhn51YBu6yBOur5sKsF+BOpLIXkzAedv98jR0eeT++UEgP9lVDxMNuFe4HZ2ziHWz8aeJ+6MW2
uOk7SnpjeOut0ksLU160FGedYBnC8inZYqbB+F/hUcdAoZtkDPMbcHmp2Xj+KybAcQUEyxJsOrv+
LThawx1em7nyApb6Q8WqU4DKOdHAfwJPiYda0/VZT1EGs7gdEgNx8eMqphK3iMtNY42m4SCib235
A6T+zTV6XumafL5ygf0pi5ZIWqToWl/5I4raXJEqPdFucnKZM7ra5xDleYhq6+JOOiG/jRzw2oVP
FZdOJ8izgdxFUJW8xLsV5r24iO7ARJTMq71yUgheWC4x6/xN+MguCz5z1MCULlQiLwJJ4FvgDOIh
/aMoCnE7M1BnNSZDCW8lO1rlD1YsT/Ki4IeT9EDGXHiej2ubo0YEagXQQr/BABynJ0sDzxNUE5yu
hh6j60qnLi4jHdD7SruEuiBbhplV8Tqccg19ysyUwv9gcy2jobvpWnd9mwGL2WoUQKV/Xin07FOz
+WuOy8S1ulp+CdzRx7i01jB5SvhjIPadRzRCMQgyfn6iBoSNVIUIZ/VfhawUS1FzxheZgfmP9dFZ
sXIEkZcE6gLMl5lt213UgYXOmgwlQv9LH/gzrONR8egdcAksy2C0W40Gb7fYrwlEvxCMUyH4eBFt
3gSlXVgPyrhNXrSYMPAqWYQo48xDX90sYPwLEm5pR0H4w/yXbOqqzbaiPP3DtvOUCNB+RW6dZ0zV
Kxqjx5FJeMvBOzUcQFdreYHlqLdDtPKk7/fHwOKYr5l7h+iJIuX376zbaklyqnBgi7wHAtbaI2qz
O4GnY9yARAE3CeOlZJRb7KfPGxY0kuZIphAOVvaJHa72FstqpMZyFI4qg1nKC5j82x+3RzLkpC7Y
m3S1Old8wD5jhu/HETqCkdOiB24WBjFEh3IURdLgANz9nbhp6637oSGARho9c8x89OHjEIguyHb0
Lsdr7I+2xQAqH5JySyGrZ7yDws/+1k+vc0tYkOebIaUm47zjz9T3M5MQ6gnckOVlOOaOOLq1Ey4a
R5eIEhGYnkQaY/iusmuzNDsujvJLY1ic/BuIaBUQRBZkRqZy3M/IGQoJUQZ+uIf7TtaDc8R/6xpM
+fOu3Gbkmvlo/5kmNbRfxiYaZWw4+YZfklSlersOHZK1eIga9jnsymEuIszA1z3CA4/v5kDrrSWv
3gb4Jn30zvjdBdy2si4gI0qOtzX1dM5vnQYIw4tkPEqAskKSPaxDoiPmIKpnh6AulBDF4+w9JQ9e
Enndj7cyn9x0bh/UB5wJBwuU5jvN61G2NyO7xAFIVN59IVxOa7muH6ynOKCgeZ3K/SdQ0gum13q/
xP/+boXz77o69cqzBAIdkCM3FYTVFlWtIpEOK16y3xhqkSHeQcee+GoOm+BrOR99hghPInQUo3m4
k5OEn8TXFOiaMMdojtTBroV37XynUTYRIoFq4C+Y5BpWoEowbDNSdL3+HauyY2zjR5CehqTeOhSe
s3q6hfOL3Z+vopkTT1UdhUl1B2yD3nxGyBoLdrGq2xXUBzvu+Z5Q0JDAs9Nk5q3DGkfuN4/MJ9HI
/je6VOaWKpguhMx5FREII32OzfYI0Dr903cm3eT+MdsVtP5iSjo3xIrsky50F6HL1Y92UFVAviZ9
2wMaW4wmZ4qom9Clm4wV6Wxm2A7gwyMbrYwecQDxG8OK2oQJcYdLUe8n8EUWId0pHqg12zRWKcd/
Ys5j/lMiePAUWKDXa01o7KJYTR4hgNCEsAbLUiBoVvBr+aWhVfN7d/PqOR9TlI/JOQttU085r5ab
tCxprs7K2JXTAEhL7oyVMpNPkX50XUbfbwGaJO23FShbRzJxkNvXKD8fBWHnsIjIsefntQ3bjO6g
aT1S2g0V3Td1oopQi7fXLhKSuou/6ysAji5OsYTXTUnTXliMpNDzb4syqrrreIdPFlVwEByM4x7s
c6yOMIyTt3vPZSK6GGKfoFT5UZYaIuHqNeC9WTDWEeD+7qIPqrXFp2SNNXbD3n7tqcWdWnW1WsSx
N3AZZsPFgle4Dv+M9uhJgzI9nxgLDBM7G+rWGsMlH20Yhq5ZfDm3xkBxM1Wy1SbLL3caRGf3cLKC
nElZ6M8yM++HhhdHaJeWyNEgbfq5YitR9ruP/hqrKDIP2fOEwq7wk9eFKizU1+Aa7SQo+lMgtT9i
5iK4+TromV7dQJbbmh/UX4Hroo3vhYlquCbGaerfBKu9v9XIJ5DCUOQHt+CcDamNKroGfXy2pBTa
Q2yFa6DizNTOoo5Nf8NOzyQscd0/JuSimXAsl6Q32fw1kY8FnjeOjMRuQkz61o5D7PjrlpFrEv1m
nFaZIM3xDvGh5nq7ckqcyHigYdjPQO9tPigy1GlryS6ChTfJWBrDAvBrNJERsk1EQUkNei/ha5Sw
9VwLRa66rRK2SmewBO9V8LZ6SXm87Y5k1bd/FALmXscz4J0cPg3AtxOkakVMaiuXo6HWwMduZeZH
zReqPU6doz0NtjS2pmy6YkgWdQ888//6n97RmxD7jVYAV54sBy4CULAVFI1fyIxkTrlcLDTlxJOh
Z6oJETQ4KUCropSyDDVD5WGwd/BUWs9Ke8fyjPEBVhegBDoEU7kGlNDtxrS4EXmLR5pZLD4iwzsN
uLHpbg9cQDmk75Kkte2IlzVFJMCNgI9zmmTUw4r3Qgz/dc+y9FxR7URKSzj0GnBoyUq0PWQ9FHcV
J8/WcC6eJaIUxZ+fJhiton1gF8nQtdJHfDnDegap5rJZomuSCx2bxjbdZrk4V00TueyhQIqmaNlJ
eb/Mt4duITqPxVOL5AaGJb7tTitFPxDWxLNY+iqdiZ4sExEV4MbLg6wn+FEtNAFmu65RttVhp0zh
lTuGiZ5DXNr9C71EsgMGvijG1HQJoRAwskbO7mzR30iRQqESnIOovltgLYYHrp6lXJrFPRoXxPh0
/hOhVq9RRvy6/JSiY7kOQMrjCIQZTvBMcwzy9zisGzxWAo/CFGMNXXsIUffjddiBAVm/HcDdvMh+
mBmzpi0wK+K9FwIqdj/HT1T58GS+j6O7N9/V9Hn2a1QQy6i7BnpEodfr0hPyb1cFhXofYyg/rBKr
S0+NaTHbHsySyux08BLsJOCh6oQXZPhArb2xzB+43eW9abQ2mBZEwnQsy19tGPnTb3tSkbLO/QfH
gptPwpa60CTuQjVDgMbZowO8Ayv69Lkg07CYhNdNUZPKJCQ7+VaVFrdNtqqacbY+6bGmP9IlSNYY
ShcK4ku+V4Cr0wTESSkicoOu382aLLh4I8GMWAKszo5BP6gaDPsVLTnmY5y7CPeyLZNIyh8wnwrA
M7HJ15DHcQ1gGWj3rczAUXGwip8/4R4ymBNuYH30DexUkbIEdFG2p6Qb06cglA9Jn83a6kRJKN+h
QTfoWcskofaIXUpehu8Ow5wv68nIkBAA0BaxyUtVWH28qe5jQh7AY8pmCQZsH5Dgnb/xUc8+JXEi
pxjxpRoL2AR+CZ/xYDNf0qvTLc8ysQ8EI47ecPD9Bjv0udDlqFmZaXyGWOBbHK92RRHLOBrwWvqh
JUiQ6GIjarsa8Y2slobxmVeAPg0M2aztjyRtajnSuCV8kMRc9BTD4v92A2ITDLIhXkM8UyTkbIb6
hOev8R6jm4Pa1lcFN3YYgq7Y/QKI+Xg9duaNEzmmtgOpBBzx5CtZPeUg8tZdS0JwwWnvnT7EH2pN
RLIPIQPXHdbWU9QMMRTqEanNSbVSuwqrPGIpD828TIGW4UbaPP7qzA0AbYwip8P2balEcHz2fygl
td5qBJZMljRN6RaQ8Zwa2O9SqvjrbKIpK9kVU+QeFDaxbU/9C8lDwpx2kp/Y9+MtSnPC6JrM2Kvy
6C/iITgLM9e8/z5biEs8GeRAist0cDqBlBsR4hE24aUJ+ERQHAU6dE/frIHx/rRTuNfAFl21iJNF
379zfD7x75oMG3u6ljCzRk/ExESf0VvgiItCh4Vc5InHQVApishzB0PsfGrtlhveKSapBcJ5MOU1
Lx9uG6oeopBEazpC8uB2Fxdw9oNtUGJ9DQcDA/F/wwBnbkQfiW4puzp2FsR7SluA2VxJry3OphDQ
aqnhXMPHxum8hnKZESth7mJy/esTXHTsTpf/1ZV2o851SzLfMzhsdTq/KaeIIgo3zd8oZqIeEmoJ
UQCht9VUs0XAkL7o1ZALsI+I5Flk3dJbRHGFlq+WPuL3mADNPMDMYbDMzFVUXRuDHLJ8U/POL2p7
Q3vwrr1YaTBE9cocQwQFz2c7NHoHJ+5b40m41d3Opb0SOAyzFjzoesYK+d20kW3Qt4r36ZafP4GT
gKQjeJUd0r0nX9WAXjejHsBvlP+k7aCpj6eTAgFYUFU20XNogk4htrDpHoJHPPSo8Lu4h8pzVadR
Owo1L6j+25GvGmbSDV3c62P1unDKuorOvccXy0lJ0mkF/T2nxyM/Hs/xJ3dzdfc3ofjP+LZ8p8DU
lK9bF1h2DhIY6Bx1Q+n+ODNVBCXscki9G16xLu2iGrN8AsK628P2xq7GtgQx9EYZdWWWOBqtLOvz
+P5S4qc17P4EEkjtOA031JAc1B/wS7PfkJ2ya7hX4DUvrzuutLHJsDhFN2zRRIkhsfreLrf5GD00
wtHldgzH+lKY7SeU+7R6oC3uX78M2bsNwpgwfpPXKBV/OlN32DkBNN3DziwXl7WyhKd9YmwheJbf
QGQ3y2QKhfUqb75yvEyNIlblJNkSCKobP9he7lN99fdTawLZGCyDk1vaKv6qhSvqOo7Aj+xqQpGL
z8Uag7BiQgWGJg+2A+T/E6ORwqkO3rhLthAdxkzsFYAIE1By2ddrQSFJds4+qzcHsqYMnVaJ28lx
h1G8ev35Ywqpg+jtSdqjh6C4R1u0pm3WhrLS+PLz0SnzEl4fJ7ZQ13GppjFcCrCpBR3JwoAtnTIA
91ky4t640pJMdx5QenSFk3VFgK7S+y8uWaLNL465tDoHdAGa9ZPiNUO4v5je4AO2brxoPPBQBcWA
4S3Cg0bE8Kej+Nz7rbELud3DR81cb4nBRzjSth0KzlPH04UYKR5JJKFmMxbaPCbcnQtPd203tkI/
SiSieGfrpKTmZKOXuh76CmWbRoTT+p+neQWKJf67dxYDCbm8woMkhwF7zQpu1XV8BCgPFe5AKg/m
hJM1BE5/JNgoONpGsLXxV9Y7eVoOKwQYZxegnqHjd2f8zx17ZvU6pV9Cxjwsd+kB+OTrCljyHGcr
KItY786V9kTlcDYXYFXT47SWrYFaY/D75FiuyaV/OxbtCuIqMDJizwcnN2X4oa9opSxkVrrdZ8g5
1X9soABivxjAAi9wdxPIyCRwMERu4EAKnwSylvkmM6wHs+uPmayrB43M+HV/JPuXGq9yIKrpqNNN
+tvUR34sramWpGoeSsPBjicr23QK7YCLide4s15Uf2e6yZXaBNGHs1nLUmqNV6hFZGJFxLZJ1sO+
lQvEwKVXM/QuVC1T70fZSvnEFrpkeKiB5A2eNeilqqJzI4Y5aQatySvMn+DB/nmaoj6AZRG0mItE
Z+jkOB1FdFv453/T82ebRdkGOMxS8d/xRZRJACc3akAKUmKHo9Uw+QWOFp9rXT3CE0pD+AfbtYfN
beGO1SvoPKvqdymoQsrIUWOSfiXnfAUQ04U6MMYGxwZmMa2LeUPXLGXSOnVIIU06JPLLb+eLujSo
bpMTE82aPsweHWQg0DNRJsVKjiihDGMRbDWP/jMNe4VK+6zLUxXGnUnUpFaa8GK10lkR7nP6N5mX
KSeQjo7pM8qdrU2kulEqqpMOOESWKbzZGIej97AQWYPuvxtG0pElfAiGys3oGYQW/s7ijyGlJbXD
ATnaTOS+nxkHRv5aP884Ady8M+WSieBvDwdEg4qcnILVNywchpQFEghnAlSwSWiD6ajTZhF9bqA4
2Zc8DGl7pk7Xjt9kpMwVp4alEQqdliC5G/xvsAkal7cwjaL2F/059z26iJd4eWgapG3OP+MlqF9Y
2TefUrSm5kEhndfIA82g0lIbHtdZ2fJ9vGoRbbIWWM6nAryjR82iApk//Bu8yp7D0aYswVPWy5aI
hHeag8gUvSve6tdnPymPuxtL6UHGg84mWujwKMumFpEInquc3IM9Mq+Lzj5APV0KA6O5dDl+PLlz
RZvBzRRffah6NZJzt2cx2GIgp9kfFrNl9DaWe9/xKDvyWO8RpdTha7LJYUtW5mgFBZ/ICaeHxr2N
yqQJW1x4pKEvBeJdPogsgh7kzql8WvDAJ8KZRftEcXbGvJ0jSkgaR0uFx4vJaq2zTLv8fsGwx0FJ
ol1I9WrEUADrDyqhkmOKplnoJoGb80mdpOuowWLXzP8Ae95bDraP+epHNouS9UDpnGwDvwTNyiwn
xTFEeN0vnzxTl1ydH/SoIOWGUn0qbD7KeMbk0W++ySsfSeSJpvHd9Wyj5tcdXpjUvS57ei7SsmO5
Z3FDQH7BmBfXBtgQDmzOsPXFuR8Z0Bg9Eh4NlrvlwaDstOzKRbDqKRFMCGTxTs6IPWOPJYw4mk26
UzTdY41nHjmobxGS6AaT+Mi/4WPwFCFpiHOHNB/xRIEKLCuiyyUsrz/C4W7BpstcoLqcrusWSRKl
A/Oc4z7Ejae6T8SudYkl/x/3puaZMTMeRYjAI1/DkX2f+lVx9iVlIox+gvnWCVowzxLy2q6GyYHN
xwWTsgnEjNOmf0Ooxj/IPHt6bKWb3xoBkvn0P6Lnyl5aL76OICKj3dj+Xk2iJeh9llj4DOeLZpKR
myzlM0HjtsLcOMBAA7CXF7s3zqGJpiwLJsU5bZvONqXnIyjoLIBhYhhL1yDpgydk0qJstU4NR4u4
d1Q3B5SL/8BaHOx8ZqLtMXYmw+hdsXgrzXADSPEkh8d+NyVivEmyP4MrLuQRv9LuqEajGVVp5HW4
yJPnUcC6+AFVRAb2KiGSfGnMu0bnbU9DLJm5SkYNptf+whTtlJE+hZsTS6d7Ta4SeJmavane99S1
2GForc1gpe2Qp2BmcuJLnP3yhSyGuItDEhJJrL2j2mrqagqQIEuGbiYpQw+ws1IxPNYd/bj+n/2b
BDTdHTxqrDBY7mS34HVUNizbUo771h3/I6Qq06a5fwW+32JzB6/9gCDnfYuVG4FS/o1rR5BnsEtL
I8qVpC3PmTD8F/Zq3k5XIYvaCWgErhdsGixbNWguLsM3/xj2mALu+7RjuAJSn/q3NecssMpqYWw7
D2PQd4tVbRsA8M+3YLUh/t9LUOrTvkZ2gdBUbQIrhofVCzw0WuJggRODUff+K2BTFjnMhEC0Wt1y
GlVxehXbG5IALzKDlubELLy6EASn7eQ/Sozzf2wY2UkYGDG+HB9qRRnqUx8eLYSh3PCKeXcDCekq
BOq1X5BpD3wWqwYoiNl9gVHIL2FrwhQGTXxDS2A3YLcgi9aIta4C2Ph5a4Zkq4DB9tDn0TQ1I6rT
SvvLEZmZYUa50IFgbIbk+FUGyWPTAD0XZC5NOHey2ays2xn5XGcy/wJYSLlh7E8H4Fe0PvTonRnZ
Eo3JiXqz0qh0RiKDHvDkL3UQra8/2aeQkn9H105ouaFbRA87s83aCmnO0Mg8XK6CVVTDoDaETslA
RrbxB/Hm1Nu6ctL+MIOUA5dHi9Q8KzZKY/B6MtNhAgpbvti/H5/IJGc7SJjyZla6zUv/Tg3FRdhj
WcMU35xJbSQzuvFP/c7Mxp568DyaC1TeTxFCtLgL+cK05emMkllozu+EYHozJW6Dch0endFyVRlF
g6wks3B9adhzCSHQ1PVH//Hk4DzLZU2nzg7fFhXZgtzHxlMhLdNSNom5dAiNrGpj2Swz4lAFQUi8
UEYxyg5sPMiluO6h+OcGnL+TJJ6EcluXj253Le9OjuekOQjiJs1gJ4qJAgbLrqf/qqvCJbyFVcQA
mCitjZcvIYeC7JBNZm1LZABl2LK50VnaaWTHDwfeYHZW2bPcGV5GPhppG/8tzszerfvuNWf9WFio
S4dj2bzb+XqhbEaYz3f/Ha+pvzqM2XjXbF2Xe3xNLeprPK+O8u2SwrtSQK+RpBD8U2iebhPSgNnZ
CY7+I3m87mmCVXemCOYx7zLN310O1KqD//y8TIOzgEiYCfWIRuZU9PW74M2OBEqpVQP1MXh5aS3D
ZZzXTBBCMpb3fsNyZwbWlSbvLywrVmN41hhwU9yR1C84WrycE7z6t4hMNDSFReF1/Jsg48Iwx4rM
7wN5ONALERVQWGgNbouHHkf1MBLPaSR49LpREsMpi7o164BteQGr+gvglmWWPlpOpw/EaomQKtpy
DrM2Akk3wQpDx3vjwiiiw8+m0EJ2yGmM9+gvpxO6lzYSYh7fSC/tyHRe5dsrzpCtAy31A2dwgYql
1CS/aEseuf7/Gn25Z6rQC3sBtPcjzWVmh8Yc7RV4trkw4nT2oQk2kUOAFPmBkJPkSbGUxDtE4YBg
quh4RZdoVpEyAamAGpsTFiMrepG9sHMVwXrFz3nLGH9CsWD7+41qnt/U6n5A6glzrPwvvLeL1FvA
M2JXlPVstSCc1IgBLql1z9Ao2tdlZY5b0XFED/UuI3SqUq3ngxdq1ldBZjmOoTwQfvi8pF53TMxE
Q4SXLDI/suyyIEbiWgDqpyqkB1uHwplyqO5QAdESUz/2J7OGgddkwI+TxvRyXVa1JyjDdkwSxUDX
fDW/88Krs3dzD576t2ehjkkYUoaWtH2Ah0M0GMruV05QFmLNZYSy9cG5qr7Nbmf/yFup5TgHL7E/
1lHvc+mzNlZ5cXpfYEWZXufufLFcSbHuZPX6j/x6/tAuxb+bbRdsHYmDK+cv3SZ0kp5+BuhbhmhB
ZcAik3fdk07rngByZN97nKYc44lmCFifx6GqA+ynrDj9QKtTAkInpCTdh+BkeDgYChf2lGHQtGU0
WsI/fnD9i3dgR4lwFbSD/z+DzvvZTeQ3Shwc6odVwEpcRY9w+LWySJJ6G00uIZei21ucB9+JA8y/
FR5UnxXWlNNCI5W57UBh9EmYYTxmMB5DwAaL0cCIQdXLYoTwY5rcUix1jV9r9H9/DqrKk5Z9IevB
lgI39HwxJLMF7iRZBF9QbvoVClQjZhYL+zMRLrRH1U9hKghr0bxADg+5W09DwAWPSRAtSU03W+2G
M3eYzGghO6iVgrRdrKz3Sx6K8/Dl9NAMaDABd59QXDspNy0e6cV/VNl+WF+voiPKOs6/hIfG4OgW
bRKrCqDsEjBekQoLg1HL/1imzF8IMLw2isdVroBVl7NGUmUcelW90Bg/48ku/HcKYL2yE4+JEEY1
q98obxNmvlPspDZB0Mx3wZBww3jU5QRRHP8GkWYwOlCyQzCuv9ta+w2BBtwdjqZSJp93vfJ31aiK
OQwoPrXRRX1hR6WU70X5ajsVXNdeOaTCH4SsppFOc3pHiLeTKw+XTUBojY5b8v5m5lSrDlh/kRZv
H3EhdOYbxtjpg7KnKPFm5RBbQhgWixr27KtsD8//xhMqfYpt7xShOOhNN8rzDRc/Gh3kW5j4uxVP
VAOTwW4uE5opbNI6e9eYupsj7LvfjJlqUodHbdpDE4ZdN6hBP/mS9waWVMcM+R/LgOUuqHyF5Yky
JpNKcmWVc3SvsFja4cb8K/KtJtqkZhFMvvpMsqhlF6RNmMtSHf9DJaoML+ADiFSxHpIlsjDmij0w
Dt65Lg4IzgmCz8RMFndaG5bkxUx6eoLwWtOJj7KKKRuhDZ+3cCJftQmXPmq1I92RGjRMPEKqMVEr
tKT3N3Tgrn3AavXkAwvuu6td9bAH11JpyEIcsOCiihffOEFAcC5PL36suXg5HLPF+iP4BSlgeVS6
1eGrWo21aFSCJCDMxIPexbgQ39lsYBSYxDaL+rECG/bxdlIQbiakkDRBWhu7vHIX2Eumo+SlzW5/
E2smcLJ6nvshxmhqYgw/fumaI/VsNyVoEpT3h5+II0RFkNU1AEUfu/yvDE+jEr/MKdPUneKI7VVu
WXDzHPW7JkBQ6eP7rF7KM0R4OlWJDOrnVZhTbz42MMJFbd0W0Kn+pmZZbHEfKAZ2MUkgCEGOK3Wg
/BA09YllsNPJq8EmwZ0FnRiO4GFFWgTOGJOdp0PJNUqQ7jQ4mB7HRcYwLlwtl0tK+q2wFuMMGBL1
vHHLyf6EJlV9UI4Wf+OB8LAeAYpapZWhK86ijWW4c5F5aPBH+Jofl7SsLQXqvGxIADUYSnX9OzQe
7P9vMpArAmwdQ+T00GCM1prjPSQRA5C6HCeUGikkvTAXJwSGs7QA63LeqkHVhVt8mETo+MOvawvY
bX83NugvAPn9XOsLS6ICKWALWbhwLglYL1OyjQS0WIzRxi+z0eXpuQom3PvNXVpyTJd7WrHPNEQh
SuxJteSo3VpqBWdu0jtGnJvDazYO+LN4QfYYM+I5lNkIpXB7hyR+jdAnJYUT6J27117Te+50XuWP
0VUjUSQxF5v8R4PSQrgEJWL6tlxgvuwD2du2QQjzXtf2wBKvlvIQ6HO5V3tL6+l+OIlPsQZSjUo2
T33ohdpODn42bqC49MIwl/qbaLx2xD6WfctM1i4T+1kzhpW+egYmY7kL7jpE21eOqF2cuJA+FXad
b5dKY38qFfuDfKCFuJlKmoYQQYHr69VOmUpFDwAqoftMEBhsAXHPwEn3Ljc8JG91ZCifMHZB7G2g
EszbRwIMt2FyqvLdGvn5DByESg2UHhtui/lSvs/T7c4+zPIxgq4anYxm7cYQfnRhpnvNTykPZ9Q/
DLzm5Uw5fIUtxjnj3Enn9NSBTb2BSVkJA61bAJiGEDMvB0+oKOAPVo4JoOXp4QHKpQnN6+v+VUpJ
CXo5St94TRnXgdpTPBRLwBl08GRqZVgi8R5N4U7vM17hp8/9bXop/AejFMDsyy/Rw+146lJaVC5W
zucsdIbJzwNrPs+Imn/XDrQeDdH2Kdgyc8wcaXt+QhdVL5G9dUbhbcpIseKeqH/m1X/z8cGngQ94
716HjZiufHYqQKGSOkbfWrmQBWTnxsR2EYJAIgzLTXniMpKYNi6NTFygvG7nhumG2JR4k2n40Ih+
YIqCyO/SlNDpD/kEPjCxfCKjt0ZOZXdo6YaGoDXN+LARnKkS1qM//vl4kNF94SsGySx1L12fGjKV
yinsBLOb3esJRga0Nm1NIMsq2AKHrJ+lzsOuLn/W+AVWItZ6rfEurVVJ5edp6gxAQDN/vRwyA0+p
fkGuR0E0AyRy19HVdNCZkFCZxjdjXEzfRz2XzixPz55NcGIHPpe9yKu5WiR5CRzvRJLY7ZGyTjHq
vNUyzc5zMqpPW8RuZhgClYMI8oYLgU8GvhMgV8wJUJqYVJf3BfrDRl/lRFPRumVWtFlTt9ebxoqY
jWmEFlA0TyhFhiqByZIoe7/kKlARccr93QWlJ/fKL57YDNvs+v4lpv4uJXD9lK8RJxyAwDdAluZT
0Yua+baOLZ1luOct9UPEo9MvlOQFKA2wnU0+avllJbGrhp6wVJ7PgfqJ01nC/+i8GHoA8jQHewKT
nM0Nnw5vhJ1N1xpC8sO5ioUrfZTYouc09qIpJma534Y7mT6jVpOop+wT4OSE3Kj4tzEXPoPhWYh0
vYDS8UP6XyquPRnWhH+jwcXjpAbJyze4E8eBBTchDDk6Aczn7zBaYYvjGpAyJfV6oSqzb3ZYwdLf
NlunGqBJ1eEKDA9lQPse8cE/ghpwE2MY2FO8ktSmbKAw7R8zuFAE9eyVO9ITWU1UNGXJXaKr5C3J
yKiEqbZH1r9Y+vn3EulUQ4wXG9dNQsugEzobku+qwMREk0EYr6f8xexOUCAdE1G9ndqhXFSYefrd
x6NahcYH0VM/+TORugnS7MROebsGMwqmnoiRow08TPaYULmPTooOc8VZRn7pLt0x7V0VoalCFBjs
pv8v9/j6wnFlhGrHWpnPosCnoFMILJZ8suG86YWHHp02kMWtfwbSLO0VA7+iHmiH+WIcIq9usOdw
FePyT5j8TbdybXt1Keloh0aq2Z7Iu/oBVnJPCYMhUfXXdIhD6T3CSxUd+dgcGvpTpxM7ZIUcq3Ew
RDSC8+4neeJ6bZcqFrRxOrrbGcbcqbiTBawItHr9BxfypbQujK98wMVf9uIZ3utePVXZFlYAZyyc
u8CoRDTfSIhYK4i2LqHvRRO2jIP8KQ7BgyH13zpFVpD3WgqMyK0bKFj+y0qcfudn6cQJI2gpDShl
pocAxQi+yqMYnSKHiUc88xMTYEBPUj7/qZxgiFM/GKXKyPYdSJuLwN8ozzGBmT+A6qyP2hnob290
tetX64BXPEQS0ViHkRPa4+ltWFaEOmbPgSPDmYtO5fJu5fswtzaCsbKadxLPiXLHJULbzV1/u04h
5hWFjlYus6S4wjUwppTviJscutOWEiThu2podztNN6gJFh8FCPIkOzEi9vr8BH4XpJqFk1Ue/w4e
cdx6ggMcGEizvbPde3HLF9uXdBZFNBIQEFtTBR+QdKm6dMK6x5KGLN65yzZgQA90J45Cd4RcjwUj
L9u6bj42GGChv+ndZJNvUvl10mhfU97a78w0jahbk6KtLqhKEpiAa+ilKvHh3RUCyfppBqxqnCnh
bO7Uao0aLLV8usA16TXHdskwaslsV0bb2DrZcaU/WT0k4J1+ys7zA6Wz9IQ21h7xm24WqFIyUg2V
Ltsw4+IF9OWQF7oVErJN9U1NO//BuFSOo5I+GmZVZa5IE3ibxc6IPfioxBuYebIKooKnidnfHVaM
aQe5x1z8uZpJ4I2XbuqJC+hxLgvRnhOEVuiYyNp6C5nrZcMor9WyOjRoqRcGRmGZcInftUBu+SkN
D3DeyP5EutQmRUXnPoarAw/lxCO/KP6Cqc+c9CyzMFRWj9eM8QD+fi7BlNxRwC5Ol+nUBRrkHcFe
ulz8MK0cs7qj+PLS6LPGZ6fM7lZqU8XVu1Da/wY2SCC3YRAI4/fx3EKpU+cjt8MtUubvfAYb55m7
wLH4vMU7TSuaaa4ys0xW2af3z2e9i5FsTZMm66E25Sk5tDcrUtDY3LAkgslQgI4XD4376uk5ZYKb
QvRtHrgia4jUfQgsnK9/7/zSP225NVRIa2EdLMeYM7WlKWlBjBtJsttp6QA3F0Oxv/s4R/gd+ZFN
GGKkT9xSSYtktoXNUNCnd+h9RHlsqFXJRpfLiiGdL1z5AqHmR2TeYteotOIWB75IKTAaII19sqcE
i7wex/9sK8RnZvmB0WVeHQfa26QYlCfH5cHnT5tx5B5Qt1LFPYlbK8jGLZ5DcLPfRQpGmbyKKJkv
tPRtCbHWT0O9KTnYwmMYEo77/tszq7EBjyXquJdf4pQajn088RvnOECWsDkd+vI5b21tSPe837qR
VsP4lrK07QvxZ4b22jERKZVyOrMWMKzO2wl7DG8eZd8X47G3eoyokPEpBhOjpJ29PTqfYdzbu3tQ
nltq/CDCOorYZ8bqIaXoAkoO26aJJGQTlpprkK9lBEj3FF6B9QFR1RYv7w3vmnXiTxoROSBonw9L
RxCwjmInsotVdnGOGjk0ukAwqX4x1KxVxrqveoy8gucL/T83liJYxGvG7R8WtfDxX61balePn5pX
sP1EwZ+KQaB21ISYLBqN2Mq4kvQaiIjjKVPNmL6oSBPch5hvctKyAGQoWfEiJfxPxIXtrTDVsvpP
C/F342/ooNqr533fucCn+sKTC0V8Wq5f0mCQ8tAniQrBQzgii25SVRbsskYu27URFHtXRTxfD4IU
xBLYQcjEdtSJH9xIkwXET3cfu4IMRt+rRklX8FNEs9UNQhurLXEjbiUbIXjpYQ9cIcsfBIaUOVlb
9hA5AF+bULGPDPTvj61NyxwXc8imv2jRibPqOM41DEmkLi/VKyMhNxA2m2J6u0AN1HQpyHtq6/EU
G+IZup4Rb1Ex3o1AFXZZRhjf8o45t35z7lrzXSVw3e8u4fFUpyTPucqM1lc0KyXGxw5/ow2VbgKj
MwI+wMbU5/RvfvGNzmKQpCheQrsntCiorF64IR3UFZr6GaWCa15QaOz24rSonsoEAm9Xb6SkW8T0
WKEdaF5X8VfzckwjefIfTuJCKfZ4XdIuvuWVRo0FsBmGkt3+/6M8zoI+8dJ0iHp3me2gJvG/PNgl
7cgm8/WRycIqYi7w5pstSaQ4RtMfcE8YVQx+Wcwd1akVB7RVCFhT7uGMdehGJ5j45mEcKkpbUgv6
r+AizrsmEdx+mUs7ThnPXE3EFsbdeNlMzAvjaW+V2r5DRyhaN2h8hdYSV3gecYLDGFGCDeT+NI3c
Ie629aA8GupqrAwHn/3e+kbbbLx20xUtzypHJyIZACjOwoS6IQlwCxCNHsUrodvMPqfcXko6/dWn
UnCa8p6odBYzBPtVuXrPpj5cdhvOnXxWy1ecoZ+375BjEMIn7mByZKfulkPFmLkn8nri9nnXREzM
tEKnE8CV06yfd06gpP42F+fwAp3JbfzfzMrG180/TOFmT1LJWBKk2TwSiJep4IWr5///o81oI1bx
lJglZK1FK7ElHST8iyIbuYXs+PGy7/O5WMgisIXP3qrzfLHkmPa8BCh/2P0m/R4VwjKHMuRTBWRM
RDnh4wsxE4a0Xhav71FMQ7IW1cf6l1lFZPAi04eSNNHpyGQneYVbhGtsyS7J+UsymFLwDrF/OXjz
KE1nkfoM2P6wA2KRkehLcMNwoWLg0sOL97e3AhhARoPFlTxzoyOyJx7pX0oLmX5AjymVwLthRJc0
8tAft1p3vqkhahJHqYoV8y31oVUWe4mRMLhdI7VSyHqVSJQ6v385WNiOWAHil6g2OZ3iReVmttkX
pGXuJ61BgqBt90oDUBAWMGzB6mks0fUCf9X7pRC5yXCMc7igr5mzH041N2J6BKe77HU1G11SrY4K
yBVxxpuzUclqb2gA5JBXaWwll61Tcsa5l0pzL/DIlKjT/SXo1jHkk/oub11ZejphQO0E0xjA6QkU
cTLT2SmxkxsQkiMw77RcvpKCsDh9unvHr++5pmu1VlI2X7/l0ysif7efih1eLv0rDCbL4A5dL8pS
WHqdzs14l2ETOfoTeMuMxPd/WLhQW0j3JaSFSaX5s8rtCZfIfQXC19vBWVnu8O/Lhnyry7ebB9Ux
7EiS+eYuuDLoma1erdJqXb0/x25YlLd7MeAyXeREXTLRODBOFi6cS4zr2JFAML+ON85jA7BblSGN
dlPoFf8z4ctgUQ1EgKbBjxAahdQ/PF9Ub9jZ8NJcAmvFEnBk9jQ+UTsvG3UzFmIXJ6Rydux5GVK6
iodenMuWCQ0ssShuKI3LwdOopvsb78v6KIlOfJCCI4qZtQ3bQkTq1LnjQ15Nu61jO3UcTakNv8yu
6BD74rRy0wc/sTbZm/OqdC3JV0LRu//voEnY2Y5jdS7w5zLbEJcZxCcsLyrm4wFpvV8Ipqej6eAu
A8TOS2uQYVgmphVLt/XhdPcjsqbM61eUEterVXv9d1h26LtQ5jwwVo2vDr6NdDusP+IyXNtKcqow
vSKjPtwef1An98CRiqM55qf/8ECpzR1/d+dUcXfbqv4Tqma13ceS7OUp+62H/g0dlaQH8ifwnAFc
g42rNn5a9qCdUUR96xSF0IRee6erCikpJgXLQ+uDpTy9MPUx7GlY7iKaTbW4IJ+v0V0kNV/RlfcV
tikSH6FRV42C+IffP/0nGP9lIyQltFk4dhp8s+MFIYsq1LTp7eDkwSuIYYto24s/0Gn22uWcmQ94
OsKIPUG/jlAVXE2G843JXYTMJYM88wO92QHk+o5aQA2zrHolDBMPQyjA28+KTdcvjeQP1brIniMe
3X6lOfyVjGXzVeZ2AUZcfy7picNh0CveQJ/Kk+EfAkz2gIl2NCuYamUiG9Wf+Gd8YKnckCUc3w3z
8ZYEd4atV/+EbWAaWJrD+0LbCQsavIg4Lsbs+qZnU7PPOUh83Y0p2LS5bGXSGufu+4iEKWK/nMf/
fs0rM3f9DPc2PrCmtOFcB0rVBXrInXkievxCy+5Y1H7Roy6REdCugZgDOqr10qTNkQns5EeNyJMa
JpztMEg/a1j/gg7+n/1h62XVbCXuM98P3mylWhlMu11hbNGxXxFh6DLfJtL64OxP6KUU+6kS61UW
VJYPaTcMIAIhfuI72N0qPdD5ChJnpxZUwN2LEn8c483xi+8AS6l6MDwwLdq2er8yJrEvLt0q+UBu
UmtxRaZeoOVjcA992fCl8qQffISQjHD4uE0erRR3ipf9Cilb0im27AaWU5FglJCe/3/MClHDzvtT
FkXcMd2n7mK6tdVLSOJwxRJDoInhWVYjpQxfUR7E4hBeEqESCyo7TN1y5U5UALqY1fyt8vUr/KEF
n8L/tFbYO8jgPsn97GwGpmhj1cOORNdjIflqrSe7RkgcnYW6/pXtkODRIqBo9adENZXI67ZmHy95
FsWuifxmfMuPiqiXUPMtYp1XuJstWHxZky2r/tRUBAYTZkE0D1U41Wrtpzjesoejfz8AyOmQhOPm
8NRoTTxnuSziwNl+5wgAGr+YffNV5QcJxPNZ0pWQSZOb/LWSEOMl2HH8p/roTC9BnlMMfp27IbIS
d3V5ds2KA4dRoniYMfRWyzm/abC0aI4JF2/2q59QZaeI2pw9rfzZ0XO9u8Lbzyx6A7/w5+IsBjil
vb843WaKLgo0UsdYUaD1WlNcmzzsps46E+JdFUXJkhDEQVv0nMb0Ps2Gug/hW0s1Lf9kldT/vWjJ
LaWkLoiqbXIuqNUcojt0hPexak/9P52yyh72iR6dTfbbZA3elbApHCe/ChZUUsIEwtkExQt/nnfo
IvNkJXoOeLthRwArkAed9nzAkIOtiSDAUOZU0FDDzMT98RFQpaciIA9mbd/i6cTQ8HYcV+zq/QwS
o5c6XJrU04aVKjOWHRwL/CYfoxEV8q1YSocsKfCffMLUpTU4VGh/CISXaa+VBi4IKRVSZeaj/b7d
0imLgCw1lPinFrfTcUDQVbSyMIgiC9pcljPhAYOXChygWq1aRYOlvfMqR/WyDQM+23R08j4RgGf9
/Q9VQ+29sfetnz7y0jvww1w6Z+T0B5q4pudIw03OIlnsU5ZBwZUgDi1Rb3KBpcmXsTBO8YHIXumk
u72yup2i7KKvCyM6jYve7Tfn06dg+dEoyGw0v+GJAXQnmS3agJrRQpFbvt/j1sTkig0JTvZJtyJ5
BIkccC5U2rzLVa7e+d8hVz6gbhK72pRgU89eythQNCI0SAmOMC50gv912NoikH/VU5Rumw6Bi7Ri
1H2MoLfMYc+/U9TkB4lXA5Fu6ckGDaXwmlG1JXk71ATcm2H/0WIO/yUcMVL9+y1F+nkFZJmIayxK
RwH3YPp3X1F+umiLgrVicrfkWCrGZJjkSce2EuGawk11wpNq/Dzq0sgXwx7tFgawK6BHYfwF3SmW
E50RJ3dmKGBoeYsYnv3/bB0Nrkw70qp3mx55F8IZDV2gRTlgjIsBHZaaV/n11ViBctkyw1KoIonS
bWSUbJGuLaUDTa21gD3tFQhbTf2HUM5Zs6KaPM6AheCjjP6JI35wYHTGI/eLZrRFibajq4bxwcy9
LjROwbkmBCL6Am6oKHGqGu8mzRAyaTd1nXuEefxyRKm/o79cz0dX3AzTETFRk+yaN/SZ58NHst+v
CNEABgYAKAL2MhRa/2PAVBkdMZMgKw2KDIklHVvqpU2pVzh4BHX8Yt0EENzqVwdnqCml+8ISTZ1G
zfuKttP4YlVP5YTbzeQgxQwvNBJlaI3IZkT/W2RqvaR6PldqRQ4OdFLXBuKXyDzquFaA825edohk
Llo2jJLhrPhvC23YkQgd1gJovOFi4Dn9ir75Bphzf/Py284M8JIJ6QrksWHLeeJmnxkYSGzrSbx1
l+cUkWWea5YG21f5hIP6oawUrp8x5Wh7B9ewQXhcjteW+xV0DtLKnnpQnu+U8Gyspw7KYwgbjgxx
NTPIh/rKmwptbjBKwSCGepp+utII2P4SLHivYzYK02j+I5AZzJbopioCUizbsezH/vzztozZ+Mk+
eXQnI6VYV/h7PyNE0cG95YqJdrgeCJ2UcnwOKbUnku5h0gAIcipZ8J3+pP/GyAsMZcorDka49nrb
eTQWB0LQazaBGae54886btSE5tAh93xnN8SBK8lxCknL7qukPiEl0T+EcXvq3U9xc5Zo1vy7O8st
USqHNRalZRHhRyKyy2f96q2ye34XADm4PO7wdl6AiDhnsH1HbL7lwRq+7deW0H5Vgipnc7/bFOG1
g74UfJ7bETlrhOWqQOeGxeG69K6VmYX8cHG2BYPgowMK6r1pdqKtMJKQiFQI3ukTitF8Vls1Nq8/
A7t7RS36tt6meqk6N41eGP17hoNytZSzAdXn1HHuHu8czJBofyP2NJK83FNMc4Dfz2+3Qqp1luML
+c7YrWAT0hYfRUqL0nF2ebI4CzMYhMQDywMPwfpEUwD1TGp6brcRBNc0KpSo2L8WhOmluUdnjCIO
WgfuKzG5RBjI8s/MyE7Fk08cDy5q1jVV1uzCNyFbd+/CLjq6UUPxMZoOzMkQyBGNpt0BIyJ5UCT3
eTYEwaLSB+rwtI4bg9WrqqL0RMhRfmNv4xKWuEDggk4j171r2CGwKo73osInbY75hgoJp9xBsZuq
SB0jdPelLx78VEMlHmQ6Qv/MVn2wPVPStHUDZvuDQ8OYHhE20dzJ7f8F5tt0sev3QaUwFZYnSyya
Ja9pfaPqVZtigpAJrxvGGnAYaKiE9MH+V3Qk4INy7uU2f/ZrPFzQmS/3sMuaDDBFJ9xplzEv53e2
wq2kKGEWzpucdDKYvDmSSYwHvc2ITCwfWQwMRJ7ndTZ2kKMqiS1pyUhW5U6VwNLdWZTOhAugqJZd
YX/VqGAsNlRwYFYyU5kyNssi4daMPLIAJyQrWkIIvTbUmn+kARJcSj1p4PIeUMBhKhQ964cAq6dz
6PDH3ShPk3Tt9fmZzZjSxwMGvBVtVehAq0QT3wpa/Pw359fpcxJl4mV5gQPMIdm4BPvkCVP5KPjo
qW9Hk9OkGj61i1oQafGMYsJS23xcI1fGwjPBGAKfqR93LWQlISmq6yDmjQ6YLYhAbnQ4umYezezU
hXP/SrFdlxfFPR9AJBHzliXQHjSrFF0zOlVHnFV6Nhu/RDAHrkn42qBjPGSnuEGJkLxAz4HjFMs4
kjPzAopyk9deN+bxPWQmhh16F+WQjmr/mZe+IK9Ml6jkwHdzvvzgZ599R5MRCPwxrpeFB4UH4Fmv
MGTW9UIbtZ8Vvz7AORPnRrPECPotiaG19HI7JKr8xQua4i6Cniw9cLg/SMku3afjpuwk9B3d0K7l
ijyfpYTa+AbSwmlWGSA2ttCHAJkebnQZmDa1fqQGzIi6eaj5ct3aC8XI9kl0ze1DcPcRnDCwJDUN
gua8rmUbNpUdq3JGqQwaaC+XxmpYmMG+DXAFQX/53wiET1qra4nL7fGil3mXp6eHl2y92w7s+V6E
wO0ZL1Y5iHBkHWcRdAJIUsWSV7ZcDWjTgfFwNZvWCCgoNf3st7BHY4X0ixE/PRwPdo8fBT7jvy4G
3oj3cNntEA0P0o8l1qpDYO00KlGIahuaxnXlKQrUv4ImbT0F7BK1qNa+B6AxPH5ssTlVNG/v5pql
8Z23Nt2oDcAPb2B3bUbhscr41djbdwxM9FAGsp7ZzhDATZSCa7Cft68/ncGj3ArZxaMboNVT5P4q
7mVXbsBSvQZZtnTH4Ag3NPb0vMR8J1OKpiYpW2Btlez4FO77vKMMdb0YtM/y/Bj47pbi9mJREPMn
Pz9okb4HBCseDRRCxHFDtl2LZf7dUR1Bk4ZxqA3xeWVR92+HY5Zk7nhCoyNzoj3m6Mk3puirYztx
/ay1K+/7zCsxGZuWQ0jaRHki3na7RcAGQjAsUnh8KwIfYlJMOb6MlgVdpoUSnwj6N/7VQB6QwF9u
k6jOz/u5iQizn3mqlQDWxfc0evWzJeXRV0bbxwCl3KbUNgBeg87KNQJzkhY0I/1njxCRol9/M794
IwQi/JfXQMxxzIHAfcyFxVbsJbRugjtSuskZKtZIBd/JSA12reFlCBrODba7ytJqt5PnS/56Wjsy
ugWqo27mQCbvLe04bqQ/XHqGl2AYgeVIMh1RG2IaL+FS79EcyzyyyzlxO6uDHROt08DZKq4fY49h
V0luw0UCPcOCbRVWn0Hsbphdr8C8TT1wPQuHQ6TI4RdyOoaKSy38RG5ujrl59P8ENBa79K/QjuIJ
It8oygy6zqEq7yTDzFCinrYkf4Iof/j+1lyy4dvy2gzlud/W6CUJGXF157tenWRp3ezK6UW1TF5F
IHJ7MTLJzQFR9i00+QuY8Z2caYI1zC8/yV8r6i0W8mhsJPN/k4+X+zCRwmu6HlOME6VmQBxmsHeo
WOI4JVUO+Qb6ZE8h5Bn6M5QUZeBy8kk+7foU2SXXJqGFSCElImpAqBVv8l8TOv5JgBf94JMAmaD6
Y1cix9FKQxJ3kWYMW9m24/9s3sHkHrxA3LYDLaAjCAR2MXyDA/fSsqma7RBCtQ6XmT1+/eKVt6V7
FCYprrA7SKJPd0kyR8iwsBCY2vM+qBO57be90o9TrLJIW4aKGZERfbeq6Kz5ZFakvW6HDwdF3iAK
MR7g4TjD9etpjKFXzM/PkR9QmSCcY2zBHyZuJZRGu0CozOaLuopTWb2jhpdcHoQAzqL002rXaH3a
IKnQ1GzqAQ2nK7flnzwY8tfpE2cW/JzFwztgv0d/y3DBalcL1VHelnJh1jbEchRBu7ajX2tUDa+Z
CDIVZB61f+DJSSQ0TaHnUNVVVB80TqtLLRo2MoBnQzBZkObDdMYIfERr+l/deJbHfuz+4c9ibktL
AiatgL9uBXhNNcWGZH+5TZO/Ep5GFFXJ8rsYemKIOvU7jtFppCK5dMzcnvDY2oGn2f+EsY9nlYs7
LaFICjV3VynCTp9MszZZ2qYqdHVinzZoJbU7BQ/Pa8som90FXmoW8+vwMlL7dGO50NmX7sqisKpq
p0X/m+g4qf02Ow/JVX4offtnnBTFmqFjBp5/XbO2h7ABxY+NcV+YELrDMI7j8xp7PiEk7Eky3HKU
H85kKuG0GfgMIeoovvLs5/zVLN/kbcCOgIpekp10WGXVzZ0beS1tXZwMPaCV4SQKDZWQZnn6ZShh
dqOKumjxMzEQ07xuDswwuZt+/i0Ugyz8L9H2FU+6WmQlm9YhVM1hxipreMCnh/oBBaRgFI10j7K6
djl0NwhkBBWcynvdM5Iq23Tzzv5o4MgPwRKuM9giwZ5jexsQhADmWQcyEzFkQFSzYtMP0XRMUHWx
ykoNzank7Dy31sJaQQUpEv4GatJmiMZv6qRnsAM/+m8J/XDrSOeSPB4MKd3MRy0XJyYZwmLPxEwA
fqGfUB/th8N42uxe+Bj9Qn6iZ12beQ1lvX0ad8mi04EBpe/gcqXRpzcO9RkySgn5WIvHHSGXH83l
l3dJCd3WXnuDWLznN8McJwRvSNHPqZLS9lEF2g0Nw6APE+M7VZq2EprL9PN4o2dMyQBAt/2f/Gn4
ONzl1CV7ptnmfip6YRs+SJarIshIxAwXvxpD8GWr9Z1BspYYYbyjfgA0iDlsSbnjGABvqNXZh2Q/
YJmW0IfClZu4KHn8ZjaUJnibnreUDSWYgTiQqCFDC2EZYTJyE6kTHK4tZ4Ec+oqfjzV8WxhwsLGj
nWpjTm4SCj0W6ebF571yk5dgk+ODb51uUPhZSqyJFbk4xd0tDGpc07z7rd0n1rZfzXfo+MJB8y0/
NDBYdB0Z3ng2crDnqc5rXTFG67QalYeM1KDQWx+8LDZwJhrbL5nO5kv73FGbpwvNzF2Akjx7s01T
/OEu+n8Bdkpv3+yYRmsdn/N7zfg8uLIwhL43DivjUoquvye2Bb8ArylfPiPGDsaMvNSEHX7NH8nN
PCpFwn6sJFJkHEW2lEx5zs9JqK63LNVfCBFieHABvjK6CirV+lbUCu383Ocwf0VAJKjX9tfJibpP
duuLEFQhQVPVcYVDyQRvqifKw5kN7IBVR2z3PJTjbMtfFwPNkKj5SzdHu34BfyyRuPkUwOncAE7N
JH8PuKF08woKDBeNqzXMkBWdKE00Bb/z2tc/o52eOgXHcvyo5Tdp99vXVWLMr3ld/zeqBsA7SqWb
LzJnUqseztRDzvDOhZrDRb7mX2lfZS5u0bRsgmmsHU5RHGGwH+G5k4yzglVDDfzCcJwTAaO0o6Ty
JD/b5pWlok2lzBmsjAKP87Wp8R0WLaIUteJGEOB5PnEEEVN0AS4uBiF1PuOVxp3xGaL11fIsNawY
dxj/LnJcnQ859DTvM2s55pwhzRwXIa4i95kptwGD8udjtY/SLVUUWGnT+malEy60OM6YEvMa2hJv
XHs84CPXmkhZ3QSrC+0q3AKwARlPhlib/qByj0IpBIyerDIN0PD5kRCGWoWa3+J+s/cjOHYZElrA
3NWZGmg6q/RJc2kXszOgw2+4Ns+9hdYH7ygWKn/KPTjGHQJN5CBjd0CvTQb+PW4O7YGuxgNPRO5P
S1IPXglv4IRJpIrllQGTkhGjzeizxwwVt0Yt/MoyukHGMoeiVXEE3p6YzUYhOuofk8vYhTwjmak3
JJOpTz9qnT2oHJXLfnKw/ymWoAT60x/TFHqrlTymrGbhkXYlvmHxiZpfGuY+OEy72ZFs3BhlmS0B
L0DHrUWtzRgK+zmkx3blaQ3pakNksnlZ2nhpqYDRrZ/zkCBiFS0mmCOAgUAP88XQg3Jd7RKhaOq/
wKgkozUqS+45rDtqi5HPX/RgejvaaMfsV/KHic3Rl49QNXNxaHY/JfcQl1Ka9Y0zlROcVdVsPxdz
mI4iYP3yRiBHT4d5tuxINrbz1/EMujf3Nc3/RF8ZcJJfbZ1uOriNA5otPoR+YN6+i5UL9MRLtjCp
VHQ4Kai4BWOVSUa/XzNqssw5nKZTDmwc3IKuC3MXTiS1/dZxAQeHdP8AdtnIbZylkdBkd2Xlb25/
TcFkouHODO+/Wy8xyEpDi9XgAdqg3BuosVikqH+v6JD8a9uO69qbkxCOHMv0HQ5nzem90wo8/w+1
iS/anPNMl12E4YuI/VvJ4GlAL7odhc23Dxl3D7aKnZJAPDkRdfDUPXBwtcc6V2bmKq0CgkqDVrMq
8Of59Kg08EysAT8kcgEaN/FP7IBxaVTNqec9Fo+0xUsxdQz9DGBWz1T/yBIqQFXAtaAyotgr5qzX
6od6os9dl2+gp/C01D4/fFVxV19ZXOGwa+//YI+gS2yySvbqjdhl72A8FC77SJksTPdWuqldmvQX
wZXbn9+iqyq6XdBWrYTQqq//OlSaXsaEXR0Aa4uO+5WJQefvOlZ7ieH1sxn1kBytaRB6tRiI4RgM
cBDaEgt0URaV9rZSMMYhONUy4Ru5ryvo50G6O0AdF1F0pRFTV0CgyJf4//RmD9gzhUd/Fs22aOSZ
F22GFBoksQs6wYjWvkQnRbAYaRpdJhXxiYcm9bsTK/XLaQ2RKr6y4vuzkiDf6hCZ/suxdgWMgeYx
EV2iN3t+VNJgwvtLsfYOXopa2Yn6YtKkCAWD9TC/qAqXBI5Cw5arU6rePL8F/7JCsfiEkCkM2p41
GXfnoeQ+K/VHpCQDXDpj0Qn8r8eN1x9NSG7ax3RBW3huxsJt85Sbi38NwmCsBykaaZTJN1uKZOXq
E62T1UET8z1b/dHW0okzNND0hKvvkTz0GXDsEEKtdn36uvqJLUmJy3dDyNJ08+cvUgOq60rh6hjD
yerw4t+ZPui5+TpNkgXuydJtcLIwHOFhprNFtVOuPcdy5G+alHEZpKJgD/D4zoMh+J+baXAnbuVG
NZuB31GGrq+tRlflw75pbJyiTjLrQZfz4/rcHbR6FkXBjSE3fB1OptmCAboHWC+s7Sa7I18heUHQ
csZ9m0A9/FXdY5dZcSNqW1Qu8zTuwjlxZYu7tj5K3oydAMNxWwPbKYJrSVbr+cAPzFo/7vEn1CbE
PvY5j5sdh6cMcnLSUQcS4Qqeoa/J4ozk1bKE/q4ln/3fhySjVjRQqWsZqsMpj0giBkv1cwciwJRT
meRTCK8j30j7h7WIhmRTVqc92ylD9qmGEJPaGssnyh3u5wMafee1xiEh+mOIqF3yPi+w2FaUx3rB
3on0wP0fCn5mGkpH0XvBRj+cV7cGu7Owx7ZkjQnaETp/tCFeloafLjFtDf8wWSf4dv4Bp90pYOgO
TpITX0dyrBtVjkFMxPer6eUV/F/OTeXjR3B787WP8QzqNrIVdgI36MuPKRb8F1dpIpncL+uS3d6Z
3nc/wML1iSh/WsgiGwsP7pK3SaTEECFhKIlzEQ4hED6n9XPKm6QjCUHmNhMC0E472fuVEwmxZjHs
oprtgqKPQl2fygdALn2o8S96foBzYOwhzy2SmS4J6vKkS4Zylx2Tde4qY29Z9MmYE/6oTvD6m0I8
SFiyQTMX2RoPoU4jVV/OCnFDgLcvLxeXDwLcOgxCCW9/d0FipJqBRLxZvvteuLHNd9/a1wY9vPHC
42rCDgIuPujzbfTTL7hOxTw2YUb7v5ehsGMV93doFwrkPNKG3el3fL8nzEd15V/zYYfGa6OsX6tF
AjsdVpfFgDq7PnkLqtzMyLC4SYvQ6lSOYZhu0qjpG5T6xic5T4HNdrXLkpliLF5+4EPpuGNUySxf
SyWvYneevRdNuH/cL9PcaLMZEcZb5V+u2g/5cVfyn81LMhn6Q0TFo6WRG6f3oqf7uoOBFjv+MB9T
TMv1e3jjLVZeI/QTHXwDd3bkI9oE0g0e2QJ/OKRkShtRUUBd8xoR99xjUgklB74yEH0vyA+x6edf
/Gy6xHLjkQDzO95nJsHsVriNNUtTnQ34Kt2C0u5y8kK58qgL21FNTcsGvm/IMZ4FPtFoYYeOOxzC
rLEkKI9gb3XBC7g5PDmViCDsEjoh2QG3+voKWoD3fPRgxcCPJ1nEt0ntMexrdd74OBFjASd0woqQ
t7Uu+cIGVpdy0+BFZCyixREwcEHxlEBbI0FiQcA/X2wqiVjnAY9BM3ACwAAMcizoY6tq6TmgVDET
Kr5MITxVotCk3jsIDwzRMTMU+80C8YnBCWQ6sUxg3CFvwTNJ0vf8XJLOUHNqH1P5CchIqWUSS/3k
H5R2ww6jLkNAjbcvcMi/YTJvohh77lv9qImsf37DgRgczcYWAWcRGqyjPBIDw4LIZ57yEH3F8DHf
xtxQmJbyiVOoXTVNW72W9O0K7gPTyot4ABgNETS+kbsJJY8vBcqtgKdg3WXPO9kpDmSaO0ciVaYW
ui2IrnRTD9U0IdkqBCdVR1V7TMHHqoUx17CHuKQ9oTRg2oSyhHuU9bXHVoO5cttJ+EF5D5yCJAot
aqijnxYYUf2cRO5tUrLZ300We9Lcip84rxBwmMKriqAWUisYnAIa9t+1kZb+3FtJ+bxnmwItu7Qe
Q9mC98qsbXxdj5bGxSQn4wwFCsw8xJYqGBT8WVQka2koNzRAjCiIRGaaAK8l2LQXMRG+xyHJEq3/
R2Ua7CiqI15T/Sg/KJnzvAfxc8rOcipHEpAsA6EgYgQobxnt63TORzvus2ZaHygIesxFePILmiFI
vV9QSVIqEbuXTiUl9OM/J1hi1mW/1u/gxpcCSZQrF8I7dry+ToTOjiFruvSUtx0gMF8YwVUm9LU/
bT4ypjXWvedOdvGB6PUr1uTVX2JRyNh2OkNXHksyIgHAcTj57SMrmbHy6Xhqu6I8bn8y2I6Qu1+p
1970Fm41VjGajzZ6djWws5M0GuxgO21Uglb0JRLixok3nujPs6FQeWZFVOOXMp2gxCwTt0VjCpyN
7HhiP6Up0yNwtFbeuPXcsisdwysljCwlaJW0DhL9utz2TmCHH4oCBVbEJe8uFAfhTlb6+82g7MKY
L+X20EhjOqmYR+kbiTCKpNKzINGVM8l5mzOR/o3FcckAhNJTM+bGjYjU8puhmtdx0F5CVI81e2X4
kGulzg2+jtx1Ei1OWzTsuL3Ydb7B89BxF/OM7CqPlmVOFv9P9vGffbQfLoP+U0p4a0PRpH0r1v6b
smw+6hYLE0iGeNRiFDpXn0k4eGEMjj211O0z0dpK/HxYy8XFq0FFgT+iDYHEmkjaqess+YV5fsVI
HkWwSSEzOHbCAbrp6M2UYnVjuDCo7WJTZ9i/+p7aCxd9P2h37mEVW8mQBLQAluzSSLs7vDkIqPzK
tsMnVTUmuZvr51kB1BAAimGRDOWRp7XwMw59xmxCTcsttu5TS3VCz3Baco70iQzoDJbz+8MmAQr8
EEBnqonFKmJQpgaC+9HZXQ3YIwGuPZc3h5cwIT6jDOx6hMfWNT58ki3xvhZmIagsCtaNhF9JC/c0
Tjeu7if2ojIoCSg3tRoAUBbbHQVnwXGO8bYBRnXMpthU33a0ZW8+MUTMAm190f/tBwvrqc3uzbvf
uTnp0QeI7WO434GJPDMShtAGYmIw1TCD08ujehuCPx5BtT9tzJF4FcuOYq5Vr/Uy9/6YRGJN6pxC
yi3RNG1I0Vl1jdFaAFSolzZD98MvYw7woQf0aCxvoNojv2XprA//t1i0RGW2FKuUm0+6BAMnZj1/
Dp264Rm5rT/KjEM9ErSXrmaLkT2fNy9Hizd/UPY3SyfGmQMx0CUAQm7dXx6qQwSrGoAVvOKOeInS
I6bvjiUWFsGpxR31AznAH2fJEkmH9HCXpSROQ09uHyLLfeA9zPsSFtbmC1BnEnl+0ve+VtkqWEjk
YVNs/MosenjCIIMfFjGxa3m/AD5QNKpP1sLPX2Fm2XaI1Zmu8xc4TVXYtxehdz1yjXUpIM1hH+YD
oE19Q5LJ8933wfmyx4+mq7p2AU+aMWApygZojUycyWyWHoAur+YJfoFzUUioSXKDIK0jrAiBjCYa
dTo3LdlMnB/VjYtqfPObwIoO7Gs1255yAalTJim2sYuK7nIfH5OM0hG0sHo8WFHuNSJ/QDMOwE8G
5QJH0tE2Yx6fSBXJkYT0M2wj78ZO1GFEhrGzVXQHm4+zZByjGIFkgh3CgfBdRsJOu8g0Ku7x8yeB
RbM0eX17c+xgT/0RL+SQZ3MUiGwC1w1l1OaItnOQZ6FHMaF9sPWtUGXerk5/7KGxGi82OyxzCtER
r0GFktvymu57LPOWwqrQziN0x+J5gsNAQOyI2wS1JpRI5m5RZBSNE3BiWmxhoBq0rrzwvXqR3yOo
bRNdI9MoZNM/is6+uEoHNSpRQy893gqBf5nCgSnFUEfPlXS+X9XG6vBuh1n3gtJOTk8G0bIxvlTk
ngojM7pTHGFD97gm1/BMNKDLEO78wpXCLMmsVGzvk4ZkK8TDKnFEkvRISGZxqXQEQP8ZJ0HMsO/v
ExGp8zTkSPln/9ChngP8SoTwBBZBASeNmLwK9IglYmTx3bocFX807JqtT0L7mODt0YcNnkMllnrj
EUfQM8gxykAAvbcZfE5Tm6z0hOhSoyCjx+tOQxwXJlJKe5+V2Myu3SNEYs1q1uoDLK79c6e/t302
1Twx53Gi+ay6uwH+2imjWaAHe4kLL9s5I0J6fxyFSpatl1evM70h98KnuQ6tDt1tm14ttMygbDTH
o+3g7om1aMkeLIezJAyuIqRYlyRlzCURS9BNKlF8Ar5Tpcl0W6fGlCgm0BWb9zfXQ15VZUTh2zDA
QlEQZaH9A7mvTWUuvSKl7YUmDqq4kY9tMpRPddcEEeT+vYNz8X82kqdR2oX5k2qhjbRd/3J+nNro
alykzeeVeS589jfKIvQ/Rj+H3jwgRg9A/XJO0N8Vm02m8VUjOkoUqSDeLX1vmzn6RMdfrQPAp6T8
S1AaWM7YqufwnvqMMD49MxI/TFT+AI6uB8GDpQhCncl2E4ESJTfB+YRPtcHEc8qa5ieNq4yASyIA
nHfAXdWTbhEfKK+98TFV78kbMfdLBJ3GyhsNKKxHZH6DsNjyGVHsqASrn6FN6xZ6ohXE7/Xf5oN6
lYnHXyzuNsNArVxNxXRKu3p3svQ3RPpZL/eCBptUu6AL/+EiN0msXZBXEtuKuEiZKbsrhZJujyFg
XtZs7xEUraulK9+aiHDeml1RRSqVxRTDBciFDMqNDFlwDp0z63UiFKx0O+WrN9jrqrSpbr/op6Gb
tuLt3CSY7elj37WbbhKHL5odIJbxzRDIUGjWdegA8sKVxh630nnBltQTMCKufwtvRHUtPEJtN3jT
32EXIA0MB8iwgIwUIQ7T9qpS1wsG1fVT7GlXnthfvJv/hEC8jvJcDfWhVjb7B9/dJmBZlawi6ijh
XD7B3Tvfs3E3SeUsla95gZ/XSo3gNsMS/g0N1mbaUowO3iczcHt9RJC3JjQcLhiMex/efWPqX6oD
9ueENfDlmnsp78TuGdrq6bsi4k+TGxGyTYydA0GDXUyqUg8o/jye4r0jf/k0QH53jLLbUTrPLGis
QuheDpWeFggB8oJ8LwWCeUoKfvsNnKKDMt2cfvPc6MeJMTEpjZ2DCsJ6kpFwUsXfx5fDRvxp28yn
cWA7bPZhdy5bhI82593X85Roi4l4kGdkU7atS9TKDkwWOHv9G6EXbrr0TfOeE2F31Ifv2tZYRGGf
Lkyo1yU0a61OJfGJgGFsBGYqWxpgOPGJT/U+mu/vfHRCvXH5U15pJyBn90I3sTmlR7Qe5i+tctrS
TmunC0ak5gPV4gBuyBFOwrss3jVXVx9E1u7VNsBnbMSUIYUMBou/Fisi8W8OU3pjMXY1GpsVGdNf
fw4FRCdRpv5OVEXkcNZ99VUdGbhMWDskdia5j92Iv5/69XgeM3Ag4JWjO3ZU+gaI0UFTMlOKQnY+
YQag+5WFoDqRIlrgNV/WphePbviuinlaq3dhqsGGRwTkVSC1lgqgGGr3Auk48SR0Ok0arnSohe0n
9f0Zbu7eKUa08tJNl2GmZ+p777Sk/Ng9DjGbRbJiVbxtN7unPoQMoqIgJ2FSwZ9wR7ZPnfMD03HN
SLenADYVXKQcgvIjkPA5e18fefXaIrQQfy0OSnsL156bKQ2Wd9BrEXv8qyu1Rt0nosAuqBGqmTh0
VILC+LU2O+K6Ot+QCPmdBSQiT9WfBxU7hB/RiKwKMkrx4UbNcYg2JR4XViPz3HEKEp+eLt/CXOol
ox0o8U7OUYZZuenAUM7P0SCZ7LiF2gOR4WV3z8JYvrhBEJtRJY2mLsfk/v4vg2lkIR5UKs1Z4b/a
H4+6uTcWl4nLnrY0AC3QmL7Os99KxEfV1/CBjb9Uy218X0MtehKniNQ0IMNDDuou0skBEsI82jRw
Zf+Fbt6kPM7zejvJdZfizxc8psS12vTZQAAV9Vd7ErwObkcqhOD4clbNDn/htizESD5BJKzbcDJB
dwTjQjctAzqIv2RR4EwFyWaIR7K/Va6aFFCS4cuVC/7fYLrcSJ3NP6y53Gr3gluagxOkpew0lhUk
SiJ9VTX66UYMJTp9PiEju9se/xXnLoMECBEtXNrGCdA6wbfg+O2RyuCL8wG4gkpNaIkPtBUbZJWW
umKk7h7tBr06xBvboKExIqD389b1Tg3YFTXUz/rvRHE35k7GmSdgt0Cu48DqMA3XxZZMcHDM9zkE
Ep+5OK5l0iHoql8etmlh4eUE/IdQD2+/CwVN8RG9YlpKm5UnoAyfckJNrGrKkNbuGNs4keiVFplp
+rscJ+FEyiyVjXsyFmcBUZf1YhshGjq3OJyF5iHAu7Jby8GOg5RUUC+phC4QFuCMHQ6GRKG9fCOz
81vLHyDWX1dS0IH1AOOQAyc2xwDIBYt8oGjsX0NwER68wu86zkeoq0ylITQAwEkL+E2W46mk2zMi
K2dj2lOh/zPth3FiETCpuoFoF/aErHKaEAqg6vEhg7bN33fbr8m+RVxhyUuDdHKLuegvJWn9EaQc
IzNwlOcr2FfGa072bXArllf8JGsvDijhhu8TbqqwCouPDW10Afxmun2sD21sbVXM4MVICPAoplS+
1Djtrkcqj+5G4tL30NTY4xEND7POa951QSNv7VLuA4BP8pMHss706QNlySWZRp5o+EIyYWjyCIcl
R/dYgMPbc1wRkwpUMv5RBXy0335j4auDDDsVdYExP63Keg4rad+b3D3HQljqGsUQoFipq24X6ZUf
NQvG4KofVBahRnjzeAd8qy17Bsw4QPHvqjZxcWFO5OgGdSnSxjVxrHtQF1wQEjdE3TkV6xEESrc6
awcYP/wFG0O3jXZR89rrU/GG1m5QCx8LLrV7KEt4QukiKY/ahcX0h1Qlif1i5wrx8srRrYqG8r+a
bpI1/81PnzEf1MAqwUBa6UOxgP0rDJK+C1I2PR4HnefoFnraQAsW/1DB5s7SNiNR/l7ru6dJyLQ+
QUvkXLYbcBzx9Oe/HQhNVMC/mnSRL8BtBdP4/7TzFD5nB+zYhg4Ikt++POiHR3/wIyYkUrwCRgT5
BoQkmrBUr+G6USNItLc/a1LXJq+2iHt27MpYsNW7QahlJEBIwQoCMihmqiigIImQdiSdPG8MCZ+0
60tPSm2dUEw5dQOykHGJ3AMK44/Csnb0lIsVRavATggNJGTB3Pckvu7MpQsLE33baQdYTqRxAAn0
+95rIqtpoojcV8j1zYmx0moSzf3Ks7Ct0uVScaTAizq17H2HGjmxtp4a4MGFpFdrjCLu6ckKgC74
N/0JiprCuLSYQ2W6W2ifS1sZ8tPnFNf+A08jQWoRkw5rJv2nP+T3vXtJRXEEXIKIk0LuZF03ad44
pgWBdJm71LC+xI4CQTYbncZezDCogkK7T3iefYlecKDIiIcfZI0PJlwViQm5vd6+iNuNbc9eBZw6
0wWeCLuz88OrrUO+DeX3T9Qm5eSL4fL7WIwsvExyRSgE7w0khzF1VlIXzVQH94RTEaumgBmEScYY
tZ25hGw2LvU80EEXuYT2QNSxQMcg4CCkyKDN8FkorDdf1GT0Yxf506FGFjitNnmXmFmzsvctrieB
oDjSC+bLleHmovA7mMIpm5p/fbfqI5B1hp9oexxdGxPk9SvHPDhq4w04jFbtIm+a7SvRwqmRBBO/
I55jS7GIpEh7KYIMBZFKGs9puTexHTdw4QtKGrhV+a5FNTo0s1iCwW+VNjr1n+5ilkNIVHDTW9W/
Mnx/PRuUDcazrYRUYWv8cLNZvASPYZlHpSP5N9m2Ou/Z9zJ76SRhqjEGyQY0YLyMXUtIL6F3W3Hy
2O8P4SiUXC41BFfYXKoL7RsVzf7jr7hZ/02qoCpkzOQsnq5D8bj7mlKa5w/eKq/ARYxjnFAi8pFq
cSJkQGEREB1WpkZiR8kukjKi7JY6IGTNe1/rcvLoip/PPNSFvMxmaf2LLMVVyreznLHirUkEYLtf
uNpPw+KfVPB+fz4C7ehv/UYl/CmzdZXclVJleDCJTH7d9OV+siB7x674Ft9idko0xqzXWcNeAuJn
Vmw059iMo8gp9sXozKNj5MmQOeAyef/xMIQfSXU/TYx5qgCX1qZrKwWw27aA92FcwRtA/ci46/V1
iAHBmyYKi+QFFM+YXRuSU/mXBIAkWwRiNpbFG2mLHs8d3HwkUGUQ9UeP1Y9S+Plj3HYhF97tDgwO
dlBF/7QUZ8FNeQ61DefEWXJxvA8PDWHaQ2tUjhRfmPY+ZDsMjL5PK4pVGsUOFs6XZCmpqNKred2s
zsn9xvC6KL1qB4B+4l4AMvn7418LSgN6Qh2s5i3Kpc6hRlx6m6le/MBaM5Uwq1b8NICQPBa5yZPG
DSH1XFHMbqn6L+CmyUJ5hGBjzHS+47iHNQv+EjejGlN1Ep69IUB/8AaxTtI4MJSIP/rEf4mNKvDW
+L900a8t4oulAVBNuyXq834ER/GA4gysX1FsJkOj412+ds+PTmfn8dRVFoQDZL6j9vMOK/j6TgBW
h7ICpRaxD1yUagqlTA1uc5BIYJJ4lkmwFMelpk6OMb3P4ofbduBxW5EnsrViVAy5LURK3ACjf4Vf
k/TysOl2KeWcRzTLwnnTZZINQkS22igxYpSYJByfvtN4PByoWVkJSgpEVLNhIF7EGY58ImMsI/SP
/ZauV33baSrwIISrHTWfnhwWZ42dhE9JEsh5oEh4mi+R9lsKVjM11yb5TISKtNwpngxn+vqHUcGq
ycQBaRdufAneVWJtwRmeXN7Hyi1OAfciBa9+boLLltGYafrLhPe3AtGQT0Z5WoJHEKwa4gQnC+sL
Slpy2eAnfEzZXwBk3R5KhAF8L+W6ooxiqyu//5CzgdkVt5BWSfwVc1Hjq45v5/Dvb7iB5C3unOJ+
aTFlfP9xr7l5FlsP08cXpGtWSaZ6QmXsY+sf/Y8C130AQsRT0CBbn3C3/qbZqDlFAOLx3JajsW1P
8R8yLnmosVwOwpMmFZvs42RbMVgE5vOtI0aQn20LBGOpteBlvGPjztnfq4ESzoCuZc8LQbv9AOFD
QEf2bj+H+XLrx5DU2UqUYAjQfOPTqE3JDJusC7ZFZmpikati73AU0VDLPOARfX88OaTrJuVpTlUy
JYHYdBaHE1o6DIfeBRc+HPmCdMgDEkN6gh+92+hCeHRbjAld3i+KEX4XRwNbNqPgagRwIoNgTNIM
Cf/2ZF/Xwg3mtfaDLjt4mQuJDOJ6JigrlCsaletxdsgdmRFmeVttC1smhjIucNG5ozt4Bqz6V8Jp
qI+U6wB89DWO+p3Zyc35EdEvoFPFjMQzJIKyWWYH/fQfEDCJ0v3Mc3/kvzPR2yjq050CqWCGSINU
v55Qgvwxv9rnQsdQzuhT552tW6LJhFL7jp2byuwcRYv88PN0/Y6k7DHcm089Od5SUHzuSWcuZhx1
B6YzKoJBYsa4WEcDp+IeUPuDLwnXOmXhAPwhHzyTJABJgsZ0C8Or8VwCdPl1QovG43sK+JMc8BFM
DtDFcq40W7lO30x17rya1vGm4T2TW6Wq7IvR9oPH7v/qfEGRu8QMJEe/i4Qjc2KUThrNh3AYEIHw
jbTdk4luY4OvoExoIPX+3+Q5wBGSHForIrVqVrwYe4+H7mIRjTpIsoOPMqiwQrqqfPMzr969+jjW
JCVJO3/FTcOtbP3pKekQl8mCaKj37ts8Hq7BQ7bQLwADJwzKReHPbD1MJS7NmEgmEi11Evb9Emrg
cOA3Oo2i0eUOotlQgZ+CnPV9mBDzj6ui1JcVVGST/8XqkzgYp0/PXxm1zvm4rehDOG4wJUPkZmAC
SuRzMb8SjhskITcpI8QCUE2ToXE1HjPUWeeEnGI6veEFSX3A4fPLGZj8Czu0eXIMfSAAdIjwQuOj
+XhzCHlYWb3fnD2CL0K8qZAPDGTqZb0Oz1307zusZPybyPH/Sjb9EYQGdIrlJH4jE3ZXpykUkCXA
alRi8BCfvp/BRS11ItUqIbG6IUd4ZX4haEWXMZlRRzQQ8Q0h+f5rVF7QPrWaslZ/VFLBrrYR3lA+
9gXZUfV6t2FFxpqfl5V1tRwTqYbT8FeRlrkCJdx6ZpnRDcjDPq6RXeoNrXA54OSDrjy1bZvLPTEW
ZAi0kcrKHQxw/5cMNnZUIViNitgByRWvRonDO9FZT7veKKaEks6T3Gh9LXRObrzKfBQ/cRgaptkU
sBdW+9eA5xkFp2D9ouPuQlRaVMn+alRj2GvNoHs/5v5xNFYmUU21FKvy9Dd+uvgqbA1rxG+GYJEd
srqan7XoZR4IWzS0d8RJp6SHmevLgKpZPTGBkAqTkcQLz7hOtW3x1oJGepKdC3/TSLBiZG4PQpZ3
eDiJkNKJNKAwhqVKN2ybQL65aDUOVx9p1pRIZLCAq4x1B/Fi8F48otNKD4B3yzc/nAOaDU8AO4ZP
6L01wotcTMWE4KuNdNbRnNmEeH1Kc6rIJjDh9Dkq6uMNV9Ow8GOgA6T0yWHypp3DcBoaJiFLdiYS
9rGorLW/q7AasWH8/cyh5HF7bwJm9CdXI86l9ZGVKkF7PQ1wpm6nysxgfz8oLoy2LKDctpxKlB/F
cr9CEagA4DUFN+AdYutHtfLtW1YJJIQoqYsPrG6atm6VzuPnAu6dpDylpt9iIxw4kvH1FQERd0mD
OGvbwVDdQQ5Jp41b4/3jtzc1moMmYhUx1DaGD76q4ROK097KLR5Gc7bLl9FxTfgz3lr32EMnxPTD
F82a5uPkYWvDYS2KUw7Mw5Wu5i/CJMuOE+lWzdpdL4eoJJXyVUv9HS1VhSxP9IK4CJ3v/GUdzkrN
xzU3ySVKGyYO/kCNffCXIIZM75CQIyUs24peUJ3fHMmNKlSmmjWSQkEqOqgJ8m/3+gzdpM5HnKBM
k09f94Md51v6kFg96rSD+rTJQuPY4VzOidD2lcDVXprIbyjUYq+rvOUA+IktLm5qn0NHKjSWqyic
YCjc0girGlvhYK99ww3Uzfz1naCAWjtA1fJ84Cz8FpUvdiWJU8mfA6Poe9CxH9ibrpL7OjKgERof
v/AYzDzmB6Lrw/V1Daemf4PyLDL4aAFF5cXWrC/ZbMz4tlgOt/88ZefliwzhIK/753aXOxZPeGj5
tDnVTci2Mnc84I1ozOKI3oFXgNDABhq5sb+BfU9DGiHH6eUA6cS35CTStEsqeNXMMht6Uv2ZCLGO
AmGdjqDxOh+5r+o6CuPDmCvwn6m+2tZKVZL4A/njVHwbT7AZZWQ2bMllB+Kr+aOddKyK1uVkpJyO
uJWnTYy4RGFKU2SS4MAd7dYa1I2Uo02yG80Q9IGfig6wqPzQJ4UHO7gUt4/Kemxfa+xTTT4KxRB5
zrc03YJHggxFbJqPUFJ8l3fMfziGuMBSADLR7V0NTcVUdVPRLyRGFvJMWP73XoBrz/9YlIm7siEp
vO1ww9l4itt308yrZB1QyYvRhdQGRXCC5B1L1Fk2WurqUw1CJI99AO3PyxwqUj4dxU7YrQPrcCjC
eil2LmmzG9+j0w+cwlXKbS+CgRDNsOt/PKwPyer0AW+k/r/kplLQpjIusSRNhnw6XaxKnEmI9mCs
BnSIrO0+lHdhOzvpIfWddCkL3H529fkBAQxSIllNYf/BCtHANrtsr8k+FBn37p1C5xQbXjaFRa3q
ThU4HisPUtRNekxDIn+pP2S7yNZOlM1DUfiG6XHWUuF2OY5Pd7RtSPzwba1MHP4v0HcHMfcLDn7x
GiZdAUK85nTfoXXBp3SPBSQoF79PMmWdT0KeFJYfuWY1w+nOZtsr+6K+/9JQBRTvPeoT+8T1n6B1
ZUSb2l/4wrJVFmAgUZGWuSAb56MSdM1gT6a8NaLpsVGKN7MBRFjGLsNsZCuCTPQ5wx9ai6JjD0Ts
6BY0ymWNYAhZaPA3yY4DqJp62Pd2EOe5bdit5PiE6dHudXSZqBduN1nZRfpG935XgWdWTtD73Lfx
8cLxZ5oID/CVWUrGeMum4JbwW6wBB2pqaSJewDCvLWEgVNEy92rJJVzd72Zr6Zvq+4vXTx87LW/0
Dl/xKsa9z6KlUBEGGX0LOYiHQsBbHCyznpd522af5+9MM8MiqnOQhF702yiQscPGLaOC2N7pJdx+
lRddEuwh0wV8AMEz1rgNN2r1v+sjo7BiESSz/STnLwRTZdxCvUdSNJLPYTgGvJB5k/dQBaE+2M5x
Il6K01E6hAGjeDbI2jVAfO/hG6W7EQ0dz2uaEw8Z5DNNJyN9X1RwEoN3/EmpAsumbg3mowKZfkV5
jG6pV6xEJESdSmymfdJmWI4S5qg8o6G7uNvCFJoIj+Nc+ourN+flu7ydmf17ALmj/o/GjerGdESl
d3cutVQxdJK6VKO5aS6PviV7pcNrtgHyorIxtbNJUmzhPWriAh7wJNouzbHpDCyPHXNuxzVinRjx
gvEpW9Nk3YM0rxNOk3aUu2+Gvdfq6fEqRRY5oyYIh1lSDKwCdaX7Ng1Ri+jvyI012VnF4F57rIld
8AWlBaQzhNSF/0LsuoLDdXD/YryWdAcQLbW/0GfMMVVZWXyKBpWtYhgmcd6l986K1qanWWf4c0a7
bXeuVliCyPbyscWfBIrJws99OPS3xdSuB/hoNA4ePK31lz+EJqZEOekS+Q851QyNpKIhEr8EjhfO
JqdoEXHQ9Rv8P9xL+31E9RBjUI4Uvz0g7Q15lTNHCJNxGOM0ni+Bbk9r8L44Mk/LNAsw5LVaNC6r
VLRk2O42BfzrzSCscdyuy/sv0gy/vhCe9YCQnZmjwNOolA8EUjyZCsLRzDGwSjWxiJ0QaT/BUA7m
Yp+q+SRsB0VJLQrondFyYiN39QV4PWcQtZaEoBTqh+erbfuw+bMDeNRypLXbWjyJJZ6SN07d1BP5
LF2MHQZDx7DJxfjzT4yOsAcN7+yj5YizL+E8DfZcqQM7v9W5/D9ifRdNgm6bNuPgrvnJx2SgFpXT
o2PCZf0J2YskRmxAIHx/8xlOLuBxottzpZgSL7yaASxL53Kwlip77nq634ehUoOdOq75UcmuFHKC
vjf2IsA3t+CBjkpK6C+yrCgG7dWFg8Q6AqfMwTHjzfwruimkYAoT0RVGRHPx3tZny+Z4K7LDv4Tk
ynMAEm5OwzUK6nrxZEfsXkP60TXkUhrhSLDE+lkBHP8PeRg6lmg9BOQNfbDxfsmntGT2Z2xFDKby
8pgVzJQvigE+cZvXpn0HorhBo66QJay3F15wBQ6ZOHultkDX/6Y2hc4n5aUkqPRu1df79KU/iZSW
Bm54NabCONU/RqrrInmn3hlwTyKcrLxajLDsxrX8UL/rpFtnwxWgpopJG9jAZeKHBsGHDxfhxeHN
qCPCvCnOciOmXjN3W29m7HPLGVtJLqdncnzPe3rrs8BPteXKwTPaUQaaYsMNQUWHDI8oXOosRule
1Fx1sbdPkud2AvHYGo78u27fGVwUSvNHm/X5eZK1w1fu6RzdhCpcUReTgx0vakA8CDKMPUcCiUcU
+XSCigjrl1gcnO1/t97bY/gFD4RSgezchilInHOg9UiPvCJLMzIs2a+vRFQJpx5yaCDXq9VAO1P8
8LKwBNRNcVhUGuFuinPwUMWzXVAgI0Tm/e0hUfnQRt/dCcGLQoL2D3dOb5jM8+Kk+JvwRoQpDVPN
9fBsNmbu2K49YhjqgzRXg8GzqBrE/nmL5z2HGjt7CF8udLhqyKzAkZ5n5Y8qR3ToRjGo1MWebFw7
ANTLavGNo3u3EFqTg5ulORHJ2n2K9LbNo2AeI25BVSCWjy2NunhtLOOsE83ZziG2KXk07zPJmOfR
FV6yI6M2xvepWVpBo+XVx1nW0wNiafKB2+HhfJdB9qvWLfiqbDAGIhV2mYnEJTjdXAM7tEeGGjjX
PruExzvNnS9s341PWAqs3VvqUjIjb0xKYvoRsbNeAoQpclcV1vJgfzGIJs9vYkRiQhuDtF1X81+5
0rP3AxV6PhrmSIYTn75wpV7gXRWpmUMbL/MTLOg1OCpbWsoJfOTtnpMRmOgdSH6q0c0hVE6G008X
F72kaXhy8I7PjjItBzsyPD+oQ/IrTwKtBB6gdc+aU3Gmik1jmkmczbT4+mtmG+7yG7S0s3VOFUYH
Gyj3kQFp1fcfbIcN0oSUzmH+u2qR/4oDV/1Gh2pfsAiNpPnoXRn9Ay9+7MsAFzr/asx/xGpmZ1dP
IHlNwlsHau0UJgGoawb8/vDTsDhkxmBBgUL66XWK57oS6I6RT3F0vH6mib/QPGt9dz3nOf8VfoNd
3F5Jd3ZyNnozLsvWOi6z9ixsa5fUyrtTZE5CDV14oQIumJS55rzkiRrnV/FRYu3XU6G0Ks/VUzSC
oZT57euS30qo/B+vVuQEuAgoFW7GaMjUm6Zs0dkok8MIaJAQN3VJ7Vg3234EKJxibMk71MEJNWzi
LgtBSxXsGWwtT9sN+4rxiAYmaKkvWShrJv9yx0r9dTcv3wjSVF+a97F1j4ZbMUnDgePoEhB1fY3b
6weCQN7Xsog06CupJ+7ZMW7u9jzIxfbDK0rWtWCkImVSbRAGExKuy3fdfti6QkXXDc5SVEqbl+w5
QaWZonJTO5JQUYij8KEaEMghGVc9oVrPA8qusC/OdE+8xMZ93lvAEaIrOd5QISoxa766wsNVBsU5
0/QpbjANnrutBdKDtMb+AVbrOMyDyx/lZh/YG8D8Ck8UlPFIea2QSA6Q8kFsUeQFzqOOCkqUcpTh
7HS37DCPEYomuCrcpHXXkWw3njs9dIAbwY/7RI6aPyllORUs0RHWRZnMZ4mRvLdrk9ooAE2LqHK3
OiG5OkNiwYv19BkrQCzLruuAR2Qr8w2JtgZl26YGefEaB+hBrAXrRCjtos+5UHltFlOqih83LSqi
S74tHq82DeM0l0oWaCPTzf8hlcmeRkWE6+qhBsGcyd+kGZ1b0UibUXugWcOk/F9sCtfh6qB+OUAo
fPBVHXkC1UGXjyE1D0TTazfNNwG/RtQJ/c+ZnkmLBn64n7pqaCULQGoGtD6rqM74c5MN40Dkj7BF
RyEgi/wwKdtQr1mLCyr4+vlcrVu1b7fVTAJDFqvDcM+osLv6v5QTK7J6e7oViuZiQsi6j6uCLcU9
tdtZwCyWfQUNF3tMCHRfRbNYnZa6PtIEafhlN1H41TxJEncmMkTyK3nQWTxHKAm3HJMOGQPFEjYx
pPLBKy0b1e7BNTMPsmRlvL4canBaVvOs/4muS5BewpJ95owYHczvfr7pO6DzLqaAl8BbTNIU3JUv
TT2Ml2h53XTTVg0LvRmT6rtH4D2HFHcRFiPNUQ5L4a0kfQgNVQ5BYZ2PFbTMX7UGMwRLml9gZ1mJ
y5bXlJv8qrpQdcr4SQV0+uUyiumO9fXArFn9jZXWHW6WjaHAQ5DhGIYMSwrSfIA9syKIpEcEHEM+
62jKdpBQ9vbGQw0yhqQwYiQW7bVD9OjbTrmAJVU76Wgu+3syIqWxHBw7quU2w/YPm1j7A8IUyZjE
yKn98IMLeN0aPMK1uEdikepPginSAqBpebN5WOuBFf1ceY5c5XVGRlISyIPI3O5PYIUH36oVsCqp
xlw696InZ2gZepcCNekyugZm7xKvR0z3/Ub7diGJKaA05w3EoHoL5RP8UCtpujM64niy2abKy2TG
WhviqhXJZZpkDFpe7ecPB8NQLRex3unxp0Huw8I/WX7Tvy28LvwQZP6QSBN4wVIygLOveT8mUeYj
4Wxv/mp/MTDpTq4OZQIs6FxXFA1M/Zp/jFUwngzR6+Vhxc5mx6IWBHdEmo2RbSW3cdohRz0TrJto
kF+Lwya74CYnd/gUPRqD2dCXAYWEFOpQYus9qD0uGwXOgZyd/6hO+bFCNfxdlvfBMAwfDo/ZpOoF
qu1LXsCXM//tCzuad+VbI80eKkxM75bprGLrO3yp9mhpuL6yFzKLSSuIA8p6fmof+zfDg7gNjbIn
ypAJol/6/iercOG/3DcJfLYQh66nAuu1wfJoyWiZGPTGe5KMbw+94cHycxzpYUE9R9ueTwnISQjL
AiM88PJEEFkqR8ruSVcHRCVjh0TmhuuOatv7WP2qo5KldzwZQaYEFhVjCXfMQqcCgvxGuNPXSOEq
NUVSXA8RbZcywtfoNuSAU1lDFV53z/3Ut8IU+nd44fN4eHH76e0qe0dhE5c82dhqVy2Oz6P6UTVv
9xBQb+O9nuoyXBQHslhc8lsTNuX7V3cIonohvKzcGkRyV/L7no9ildMLxT3U719RSAcSwERNrvHN
nMZT/LC1MjrgHpxjOpcK8YOmjOQDxGKj47Ep0MjJjV9VAGdd9t6wribHwbNHWYBBezDwha+LJWVm
hSYfRG8IxLQZFWrw6khoCaR9Sqw7bIc6WMQIq2P4xVSkY0fww/MDbTvnGFEeHL9QVGqvM1MnBZ4u
udHzpAySFJZag4JMjDw27RGzgVXNfVFOEm9ekNlHzydBekMXuuJIzQeaanvU9WCgAAMRrQ9n8wgJ
2CLn2SPkZzEqfKN9ZpxvrqCsnpwXSdWO7CPNH/897KmyfPpLylfRT5P3N1yQ0r++qb0y7BhPmHbw
sZA83bYTIQPiPV3Dmyp4DX4OL6EjR/v+68Yy+dw/Q45mR96RvFe5hjJ/WkRJEKPeH9gX9MWNwS4g
4e1FmyWc8ODiYHckdpCM5Hd60rAYt+dkm+ax1QUvE3GpnnokP+lHxy3gbs4jM53R1rSiImNik8pU
m8mi55jQe43T6OYuYEzOjOZQ2h1cIPea1yhjRvsShoyYId8NHOpOug7BvxncsSrQMpAHp59u5Kqr
EHxaKhNbqqIrctHEqPa1XwQ9zQTIVH61ts56b0rDVghoVWYtOvvUqJ9+1mnnjFeZ7JsEPDjuqhqp
BeaEdZBhn6ljXDGV1T/CdhegdBtOByeqw71SyeUtfc/rP+hPAMcsgvz4yWJ/n8IAjhJhC8YNsqhW
oDoI+z2vxAgyaKmWnqAB8jyR/B9gqvetowaQAKmrslTGRTGO5LPmExT24CVXzuPL4vsdLajwEgHg
itaEj1Ub22dRqEgGqe0UhuFU7ucAB3kelhKn1tMIpX+F4FE2qXdRTI58iCXDjyC5hhoaNJkZUf+D
jM+E4FfgDG2DVxMQ4bRLedneZMKcrvkJcOsqY53pWZEVfrQTnRxtG7fuCqy6aUsqQLKZ/hMpZWO2
j2/bQ5GvTVSfTUaz5gWGsAR6xV2U/99M4vOcy6V22P9EA4iQlp5WEDJghtn8k3vx7A5qiKyLisJB
PaF7uarBog3sZjM4WQu8rMpynKi2N8dYOR89T9aOso11S0W9eYMnpe3Me5nUmqZ8hBFcCwMHls3g
40Q+HYzo4Qw7S/KHo1Jn//ef51zLkefg37lTfHmLXqEkZM+l7h9+GYWCgNY+ErbKdWqmprNWWC5C
CgWL8JkijKiF1NEMX4tETrFA4rqjMNx7RmRIn0V9yJwaSNDoHSJesx9GWS4TtGZEE3yQ7abNacrc
/XjLoXDUnJCGiqKzx5EjmE7o610NIoQ7KADH4kGwUAxSjzlv2rzsTEMPDhOW/l20V210C2hUd6rC
OCccI5FZg64vzMN5X2Cs+Ftwb6O6REwrZhIzx/p4VIpOrTklaNJu+gU8F3RlXV3PEcImJofB4vv/
OXLhd0iq1VnGSZ9EfL5+TbD/lgKhsQNB32GNso6P8sjUFM6eIrZliG3ZvRDzD96jEzuA0EHThoIU
n0opn8IjqmhWMkwKVJcGCPnOfBci7Kag1QwuUfpfPfYOGcF3UJ3DBHDF5d1E+rdZj9eBgyxCnbxB
Gx2caTBWY4Yz3A+vRVGrrUxlG+4vAj+43UybLptbI7+jMsCzdTj8Iz2z72VZiXL+tN3SS3f9uRwP
G2D/kFA1RnTMJwmtDZ9YYZyZOsrPLwfFeLR45aqGJKQQhIPMNa7w+deyQ/4iS/oKf67RGaYPoizN
Bv2Qx3aatuDYRHV/I+J1avfSLgy4cU7EJ4uTUXqr2wIwCdq2wWMyhOvlGRd8dHlq5o+D2C4BXiH7
sy+3jHLMn8JxDAJJt7wZg7+iWnpj3oeNeyO+DcHhO5NzMvF60Dt+M1oQn6Ns0UFiNGhlQzXNBdCK
hFQeFFc2MaRwCCVGz2buNWb4FHfJ17fWZBEyABiqbrkvIKj2dI6wzcyAFEHJX8siliBmP5E/A4gP
xGGDOKrJjgjmhfcFKy/fqXlHRIxOuPRIMuFVUi+XKrlxUgC8Z4mQAGB22TA9jKDqjuRoSa+ZWyjg
xdq4tuY6n/Fxfvk0G1XKDURBDGPobePpAnSB8novkpPM7DMFtsYxdu39ZpL1t7DBKD/iZenv2or5
KoQmivFan/vg6cebyb9OaXxKPfap1HSMLLMaFvv2ug45tXifJKfoYerpaw2dNQqJc4Rg2N8SdluI
hlYdzWRa6/Ki49vdXRjnLiJsd0OvZKcKUtfELwOfmjmIF08QiNUEZzsB7UpC+1584qnEzA4sRK7e
iPzmXGJMYdXbq2KTMNRgYZnaOTHyEnhE5uFMZH1tHn//stYkmjsfg+bb3PiS6xN6+TI2ZDTxDMl2
4reW3wxeREdR3uCsO3P/cw0Z6pkFQhVFtKccpQ59G5TmrvI8A6NUDTDVwA4dP6ms5+L+dxJVSYmX
nCYMHJIc5KWOpDEs42PhWFl9W582Y/XWdgcfWR7wbIRuxXTvkb8MGZkIRB9+JUtKALd21Mm5iDK8
/j5sC0aLkdpX2Na0wOKPuIXqm2uYgh4qbciB+8G62FPKEYHYiBGQSjc+kggeoCXRl6dKYdYhNVJe
0jKPFL3DtAY3k79gAxTLmx0WYkQqY/QeL+HzkM71IxIEjKv838JbFO1o22tUDqURv0gVDZAwmml1
Wi6Ov6epzz+NEb+D9dwMmyhQ7Jom47w9PyoDV698ZRxPC0uR/CIYJr3WLQfHNUVfwSUoTgQyDBLL
bD1/VXHtAy5UqqTJlpAoTbLWiz+JOU1Ltnl1CvDaI12gHOtlUQaASsWEvmtG3n447pS2/wclQ0FB
/B8e80+4qmCpaHO/np1T99dIIgXTI4aU0XvinKv//E6dQPuBaM4HYMtQXS5OdJbw9ZkzL4v6GNiC
jYycF/Y4XNJ7FiU8svfz4LxuttSBMGOgn5O6iD5QEwwBDZordTy9ykzYDiFNCBs/I0501iznX3qQ
IBQaMISXByKXOKrCIlCOqbvAdCOhTYo+0QZMalkLFwCRUQw1ZGegsvSiB7wNTtq8orTVOv1MJtNh
Fq9vyxGH3ctBEdfeVMPB0/86lGcg78EJ6kIR8AqqYmz39k8SaxozO8SGJadHXLUkTB/va54P9OCI
iyUEzRs7Mn7IDD/fDB3iUTHL2j6Ar9hoxc6wkoRxbtJfbdyy3lmqp9K7iJk9Y9m5UUeIUqPZTR4/
doIpmHEFopOAZCLu0wOnt9MUT6wuYEcSiyc/9kyys6ckx8btFnAvj8W//YZQpxcVQkcFRxNmX5lE
pJSdHxUjzTKCqmcZREjB+zjBqpET99qf+8p/k+Q8YthxdCpKk7wZ1RxBaLO3OO8SPa+ukbG5ecJI
yjvleMXMaU7rejzXZqSqTEfdcIMWp3vVW58fPzYL0kobmt+0GOMjWEE0FVN/una3UWMQZKRRqsxA
JKOXFX7o5xnZT+EuRqxc3pi/l57Zs5FjyANwWZiKZtUihlcbrByk8QQuy1qHMCd9XpgigHDQV8lt
mIynX02bJt9Fkho8VasOmG22WpIbDJJkdZq5zuBok+BQtjdcRqilkr1NkarT8OpMYmtZeRjqLtUC
Gu2KQXxN1nHFNX7dROAc0Y852Va+R6WCqvZtonq0Ahek+dp3knQeAQhBTLYiV01hcfE3D0KIc8aT
yzZr4rRMcQv25tO+FtyCnK95RAScC5C7dnFolHrAXh3COy4SlnXXey+Rcdoeykwt9lDf1yvjaJsg
t+/9nSmslIRKmKOgSdPKZqV6YQW9WSXl/OaZmO+5jURLxPmmcgG6Xm1mJhxovNB/Cu85NAXK0FoR
t1+2NfDZXxnvumBFD2LiR3zQ/s7oeG9drr4QfivGWM489qWwmCww5LBL+fvniphVSZl7tS8LFxA5
gLn4G7z+w35Tm8/5w7fqf8sPqzoyZgwUAsowRaaKkQvfQmCXLupWnI8Sg+ixjV6aUQ49V3YGXQLv
o+N7rSHmy0WBfmSsJLLHkRAkml+biOOWLhH+AePTB4ObUv31NRtnMlUzcLd5lA0bhYyk7/rYwADt
fqbBHwnClkOexcEBg1zCLxGv73ROcruI8G/I98FzHSd+zisiSSLMnUy//CtEs0wF970plbgNihWA
yx0O7krIOaE11WTvbw+9Ec9VMXnKdJDTjW0YC8nKyFmHGax0/qF7R8nZVYoMjmMh5Csb1I6TNV35
bRo34PJ7TntS4ZqxypuSdJ1QiKJMlCuFKTX1pGO8etlbk+XxjnupPSIq2XnhZYkuN0x/tvF91B5M
rgkknXD7T8vH3LCtXFZ5fDxAB3AOksPHO+sDVHBSDgSTQqIik0sTFj1kZT4OdhrdUCsXxQxtIo+W
h9fmeGKP+aexlHTXQmAfJOTvB17OhF3Q2H4lbvaJrXc+OOjttJzcXpzuSKvvSFYOxpwFqlThwO7f
Y79m8sk67XNV2ztDoMT8b7wUs24fuyX/Z+/3AtDBkJnP7bOOnsgEywvGhQg5e4ItQSIBm0qOJIIc
T0ij/h9CSDdYWxPelBh+PQwOWOPdk57cJu+iVAhS/uIsZc9EixNkDvmZm3OY0OVWrTmvdVX8xCWX
ATIa69lrQlhsGFf/PGYnCRgyl433VfrDBXMMEEp0pCFBsc8mJrFIzN2HRcMUi2UywUAaI8yrBIwK
qSBGbzwhJ0Y/KWkvKB2gCZAfxnDdhrYWBuPAGmRHRcU6yy3Y2A+d5tagtcPgAojtcOR79XLnzm4w
hreG0s3OjJX3Rs2aQNnCrCMErQ8zE351LhguN7/xJqBbugy+EQsa7z/w1JfYg93ZrnPq/yev0CaM
QXsGjkKriAcQCOuNoiLc1i91ZrL+FVGiQS0iAnoX0OvmMFfPSz8R0uL7bc8GU9fVlglYjF7HYvPa
tke/WGh59nlUdoN1toQ12TP9P99bYBLlogHZ7VEctftRik5fJc6mJNEKOwLdCkDKbu9RSWk8rh7C
anE/J7hTnjeMX/ybTudQ6Vjwc7K57dO3DJXK4W5mvE7c/ljAcjl+yMqub28+TaCXsdbf+jpR7EVh
b6aURWQdlwUIDVcFKi2Nvd+tTrYRwCbkj42884r78UgTyAmh6bhWteclQHyBf4RAovR9jFOuxkch
UNCGUYoDIm0r4K3SqWwDco/hQoCdCPx3KGUOhuDx5yFrA19KOe/IW0WIGfEZzmeRXKwkGWHUs05q
2jbbmwKjSTi/lPM0iG8ecrAMOdOHKQ2KHR2XDcpx2ihoPQ5SkRSZWFHqzpLyfbO9QYhMEeSJJr1d
i1ucdZS+GfeQjFcawKJbOCREuSTXjdbvCRTzbhFWtUwRqZMRuQ0m3OsnUs8oZk4MwIpezUCwkjOc
e3N//g2OI2N87ghJrbYmADPIlZjXa18MvNXeeqgQmMlHrRXbKFQcQBz9Kl6skODrKMK8IS6hzPP8
IR5wyQyS0RFqESe5DLG0SP7TUEBiSdy+hn3GzwkvuwDCHJeKgBExe7R8Brc/rAakOI5Fqm5w85rG
zRUd22m9eme4m6X8y3wMQ1IOMVsxhBcuBK/eUqiWWBEPjVZYluAMQsbhM0MwThHTiOS3oIho2cNq
Wm357wTSnzWbmR0P0m3M0iYYX7o2NC+fIMWFm61p9cVY8RkmVYBEhjrVbuj1HeWbhtU7/Zct47qE
LS2ItpW1huLF7gw9Nb73Wd7sAcAzbz58LksnpguSKH4roEsVjvfOXanqyJtz3Lv7BHnyekQdV7p6
RhSq71e5rHynbBRJuRv22JnQmxbLivZSUPC1m7oPQuiJEl03VNgGY9VdNtBoRbVKV0MFIRx5GxX/
s3RR059wKdkW9jQYvaiYhil9RuFKfWOhLowEM80mb9qmDrNqpJdQGY37dRI0mGf7pLrdl/jLyYJU
vhj2s6RCplsDReMDp7EiDU9ggNYLp6Q68urhVzhz27F5pF2DLZAAiDUWMEDC/FItwDmERSiBCbeU
ozTyc726Z8XzBftygf7ZUmnzG/I6Pr3DGwjkCCxuL/EFamtlf5FH9U+sdKb9gi9NJ8BHdbQzBboc
BMbSqOkxZ2mRNR1lbrnJ6oZmjqlWdZA6uCbxZDZvt8hf5nhGyyzBE3qfqCLwU2WeW+sJIaEeWWD0
NyHUBfzh9G5bR1rSNYc8fkceI8OO48YylEH8xhbva6hCy1u1OStkb344Nm/QLnpdXIhnZTsVSKlu
za0e0DXnh0fKOcVInXgS7pNxcmJr3Vpo3xLMW+GL3KfYAsCP3ldP6UTWoC70qJV2ucPuMyZ/F0Ej
JEcbXzKV+eqyeI9IE2u3zcT2PpOkGSwKTEgg6odvM68RydbcSfawVLkM4w3ou4GbpvSTkN1mwBtb
wjuBRn0NK9eYo7nYA+KKfWiTou1upYUjaxUaSU1i8JkhrVTY+m4Z/6X9mF/YxzX0ruk4nAUDFox8
geWHxhXky5zNdmg2HgLbpbLYOPUcJ38hLRf+JxnqUsDF0B6DYfIIdv63DY89SLrmQxs9+eusN9bg
b0G7+8oLlktbo9S+F/mir4fvZVpKPoq3QMCyBEAomAjQjS3hrq6w59avpGZZ4QyeQzO6t5Y1Ua/h
wSLI2QZnyGzPiaLdPTmAmCt9RTB/jzIz2PLQ5t8AqCfCIWDBSJZKEeCoQkLs8T/EbZoO4uuHaSrl
F+kvi+2QOpLO6MwFiJpW3gxUVkT+T8WGZLIeObu/U8B0V3Db3Npyzd/iHXsehs1mJUeUQwXee141
sYU5oIroNZBXSAaG5WrzPX1BfAKWn3CjkW7XIMQ1TdiSHEODHP8rjRw1HfojWKtZl2i0EtuhSyCY
bNesCLlOLJvfE6qVRiCWqIbLRomqDxhXNxe/5tC2fayO/KAXfxar2WljPk175cPOWPpVrgmN1oir
TTr11OTifBLpooWfT9AXgCIk18EKYmuJobk4ULm5chtUSfhuVpdDvajgj1U2+t8dVBOTWXD4Yo6y
7KSbmVBBmA3vlsvHVe2dRtrP3Y4YPfV0kQ67DzdVIcIat6VgXi3VACrKdzAq0GiORQGvdSYwBy+Q
CVK8TGS0sr3Rg3QmzpmfFXfbkkstJ9MHdRV1LzGFh6GFX4/BSSvKo83ijplOgjcY8w6REGNUvysh
daNheeR9yRIwfP2rE5yGDgVBp5gRsS1vRQ4TQ+d+fpx+DQPEJi+SQpnH95Dx5tShA4FQwsvt30HV
L0GJs74U+pErOdVLptWqr4UCwPlegX6XjWRxfLPyiYqajC89bTzcfgyBjEHrT0HQfRVbFOjX35qa
lvqRD/qYWU4ZjmAHHVmG2P568um+YcdNxYo/m2nVkKahl/LNkRxf1/OEvcg8peaqK45QcSpOvSHN
CgcAVso9EcGJMA2JUPLXWJZuKSkyVZ67aI9GDmM49QpOxRsNV7quf3+79YkjB3PLtSs7hBKVzUcp
B2/p9TGCIQDnubnpzAOaz+B4N5ZeBbhUZKbV8q2Sn05GuuFdYt4Ry+2o8ZpGU/ogO5iK4jH5dcMz
3OwSSKupPjyOkryeqYS+dn83GjjSCP9pWSyDbrrLEyLsaDoRKxh2z5obs/zKncpwqezSE5kGHWMA
zOYWYWQWn4wQ7q3Rg3pHQ7VIodFt5leBbhgTUzPtamOBSxmdce17QOW+rPUHBKdoABAYnYfV6PU+
ckflphfwgs6sLJS60dI7Ql2MwxKHtTqoGLEXHpnRT2ZPDlPkbofckZh4m+w1lETwooyYa4wZkTE2
m5X4rKLI3bjElRBJ34rLC/2tN7UkkinSYBlHJYjzKtxbw5yASu5b2DDQDtjofFGrql/hczqAicfI
1NU9XmAPGmf6hYRX0UQhqNS3ygrMGcxnWT8LoJ0JwGQgG8ln4zORn+YY9WdkTu1eZhvkYBOxsT1w
joJkh2ivptnYu+JOylx92O1O3Sy5dR9scVxuuCWZlTHp/5lt09S4Jv3K3qQqjHG0kmZArL55AUxx
pC1+kZMx9j2riBmEkA5nUqsONgjfdLEhFyzKviWTvZyeNx3MqK20IdVZeS60bN0zzKt7zLfmdTJU
EZhoeh/oeHrKD5R/LTn6A/zLxAPLeeQVcmReNiZut93oUW3yMH2FtJ+w671z0M/lvphdthC1iTVs
eZ5k/vwO0TXSap2tiXgYj3ll6/gJwLTYmofnIXdMnzjGvJG9AWQYaf3/8fy4TgJnejCNxBNN9vf2
RCtiYYj8UEnE+PK9fB/+54tKZBP3CLaHvxN9aXFNPskkJTiXtrAhJsheczqN2kgs4UE1tFnN9jA1
K6lXPhfEcMI8FZpDn8IyPrKBz+NRctBrU194rpQ8wq8lgRwmR0XvzIz7sjrh1w1wwAdeQC8Q+4wU
r9zqBboFzuSwkIugBrDv6WXDnyGfJuS+OEVsZ1eOzSEALjc3IU7f9hPu7B4d2o+RQShlvQt8rcKn
wSJxlSk+/MuUIrk88Xd8KY8m/qtLDRP66Wug3fpPVTY/JXtKnMOZCcxvBVCcQuPnwNZ/GqsOMaUi
VOGYHJ0LE/Ct1oSY33uOjqDYZnc2W5Fl8V3pT/I7eGYzJkMzknDK4CS81mOmZnop2X08p5aEa9OD
Hqs0OxBsLJ5eAxchZ1KnYaKmPA68lAvqh7ia2hCovopNhEnvt64dAd+rgnvPtD7shcoZ5EWj9Fu3
MZL0U3uDnuGPWFwr6NyJyRjveyxNyaJ0k9v3AtHp1NlaHwk6/xtvcKWMLsV8PgOlLnCk8DboNIJA
R0v3PiY3g/6Sh3CLMSKeuFUcLpKLdlFbR5DCvTGgd7gzRqE+oWp8QhGfjEG1ou5wuyS08axoEMQQ
202aDXDdcSbx45McxyP1nHdBWIdMQ4sjEv/OdHZtGuBGbEVHj73AaGDa9jHy6TynfQ3tAzIXCMQj
Vfdsb0XP3HC+KZujp+l3aILQZs564r0MWCBwyeQmamtaV4/NyFqCpiVvYDYIl6QRu3USgRrswRPO
/TzE2WZEO17Z+IDVpMVed+AKVKRqKjIIzGhjMd89q+cKeFzYxd+jJyT6WYMwlyRsaKxn7i17tipw
2drWo3uDDSy0KE5U75+/13aZhck6yaW3wGaVkDxBLuVltgUqXkAaIgNTCvDPtdEUeF0m14yN8omN
z7slA6lsbECG7oXh2HoYzONCuWlo3SMLXfM5JvJdbBPk5l5Ja8pbIX3fZxtxIZcu03R1tYdp/xCl
/UpbA+w7qRH7Wy2YaeJgTCMXJpe6zke6nzkRnkMhws9vMEBaZvngq8pQ2InBriAwpvfTKgpTXih3
iPVr+exu3JclMmc0HrB9ApuVHHopRPXOysHY760SrDRVmwpP2vEgZIyvBD8PAPncqSNjL4WtKttY
Ajwt4RgfW3K6NsZeud8pCmzSqF0mQeryn/PpIaohg5a1WER4/M9ZJW9DEzc9NhaP2u1gwgSWzYsM
en3gbcTez6xqNxXvnoZttJjmjd8ImjMTmfTR05/wW9IDLsPZMoTPCML257ckWRPNCW7Xkpw/W08G
66b3q8AjZVojYyGiSR22JJSMd+rqA8w5Pw2aY7s1aWh31rcRQnncSqrhc+rG1Wv8WRfH93ljjFP3
spPK+0DLGPj5amCp78IWHs36CVzK1uVE3kaAGyqhHiVasqYhbSQfrHZBbJj59o4IupY5soO8gh/r
JciP8+MtyZBrAhVo55gp3c5cUd0qNMQZWZ8ugOu/zql7Jfej9XnCMkwLKKPOC4GZ9vYbomy4b6cB
7afUJo9O8n7yvKAk7XERVktY3GeYXJ54kZnVzljFjT8ivt7FKkmdGQWHQx6IKTqLhdXkh/oJwZv7
nj43Nh8aBQBcOne4An/ZLXGKS/+g8UETfbAp6ZUfw5COJOBNlRo1HAicEspHxil6EC2sSKKVJU/y
0vI6b4/5O1fGRA+8yiHssrghqFNzli/V2R0j0Oi75QrVLLJOHOC4YFpBX8mpLePM89IDuDG2lLA/
EFPfyccOrG7TLpfqeV+5ybZxFue9y0fMPXu4FO1LkzYFoDtwDPuqW4dHohSYRNl2eVn2mHgd7v8K
lmvedBmxb65Z7jzptWV+50+FJb0MWKGUpqTd4iuCVBxNrUagTk7yubMPA0H7S4nOE4Bfe1lc7JIO
w0jWNcvQp6jHpYrY4qvfWPked9MdZ1URjYnbMDUHYAE/0/Z2nFpwm/DyGyXjWW4hCssbyHTX38qt
f0lbiriU5SO7mxtHGttTZ7OOsy0rrZ15u3XmMy3sBqU+0udKgpVUv5NyecLbb24Fjq66sYNAHHzp
AIpGyPo2zwbunW3yl1IS4GWLyTCWjT10Whd36gEDIkw2lbbjglfxgUFac+IUeMzQdcATclbgidJk
TDQRIuL8V/Y7Wt7FQeIZFFbeXnN+S/M1T+osMDhBBfGsK1KALTY8Dbz9eEAg2bWo5ILORWDcmw3+
EosWHkKADacIU721dM9et4OtpDpvc9eECOhCaqawFGXmTMTmmGM0aTa/7TT3Duff7GWv1r/H/97u
/vvo8vTfeLuk8swCbIvyFN5UoHF9pqtF11wJzxUjQPLFY2WZgzS9zf9L+Nh9NhIDgriYX9nudcYC
XXVqp6/KuELFTxCB7Mbb5gq4S82iBIfqjJPeGPGQt1YzPqA9y9iwin8av064hU+xlYHV51o+aYDm
F1xq39BlRef8KzCoocbxUY7RCMr26pgUHzyCNrcfWDLldUmMcmiee7CyeJkV3Sbh3B+ypaD8sSJa
eq8b5/n8GLAh9JSGeuGVZ3I9FmLKUdAFYU47dFNC2h2ez2i9pmCZ57Oy34OUSs8SuteYRybHaT2h
D+Zsp6gkRGEe1WiFdNqfcAQ8VEBzwrY0sWBdkWKjTQkEVC+diOhLr5y+Q+gkGB767ZJA3uAPrESs
OBaEv7SadDTpTQvyzqRHlifGUSEo9NrgZT0a0lH6lmy0n38tJeRPO2njlG5fzBBMTYoK69zX02Ad
ZMuM+xVjTKcZ2dNPtEphXMCV67gXLzp+OSB07QQDert7Ns7/RkOwZiiLpw7tuHLOux6LSVqLPID9
ZW+ZWbfQXowZiNgZDfrXRM5jXrO7N2CAktJb4wXTK++2pQNnpwmaqXqCWpyRbEB42na5ZeOKvGRb
DKFHdXaU+0Nwgd6dgIBC2jWS3LR5vHx0szxRHbYdUhm/H4ekB9qlKojT/4iGwBr/LIHLqjoIHC8/
foR9J0p/347qAVASUvW2+N0iwjhkLWeld73TfbNQLjXczn55JnYDF1PtUrSGgb+aaNcCmn7aW/DT
LP0SUaUH3aeIul+4kPKmWG8VHkHfbMAij+2YDtZrrmYqIaoTlWxUQmPBmFqSTVDdSeo6TDggCOAf
0UMX2v3n4q17VatVB4Et5JRJrHlgnU0ALNdh1SY1JcvdeIMtUCvWdcVzUvrNNnPMmCqXGLPduS84
H+TrtXwOcihouNDk+Uk1u/kCe0iZl+PZ1c5y/kPg/UhqO2CrMzau0ZLDKIsI9eTw2oZWQVPnvFJL
WU28ZulqBwUm+nl/fZQSWY8wvgJO5ZAGiRsaI3Tk+8KecpajvZn5WRE3wWEAcxY6gR29zZctS35L
eW8Gotdhinz0G245qDeIatWtCi6C0Q1oMq4VQeJq98Y18zYA1EsgpHjwYeTq705VgfJGl+GnJYjp
G315YGJB1fIeORG5ABNo71eEYf11JaVM+N6pXqxHhuaVn8DE7seBVzdG/tsRBdWag2NBZhODv1Lp
jvgzYlh+FipePONVGd4hk2U1sGmGE4aAkJSR4/WeTaqcYfPweOELWZWqjqyIp82JpFKdiSc8Vtue
xdQzD56d8NeM3/NK/ZOY671+xrqtMg0yCf3gOzYXi5NJO5cCPmNHhcIruCciGeeHXJvr/6tUwuQn
Bihapq58cXilXXP8kHx/AIqItr4x4ac1yApvFhliCOtH+/Xifxdi7JgCNu3JNqM3iCafioieVU1S
zO522iwI41pmGmUYpNQO+IPPm5O3SbRZJV+6H7yi3UtQESr/U4rCkpQHtJBYFydjuFumqzhS9T0D
kiYUfi8S7xzTQ797t0mrVy+rrRs7d4+zK02I4h0w/CmRMox6Ycm/86X4f3QAhe+DvAaFYUaHb9WE
ScGrzWscA4enQPKYPeUAJq0sj1i+z9PWkXId2OZHkMKq6Ra8Qs55Uu2aS0GBM4FEbzPch79g+g5D
59UwLV9R8cQ6/HzdM9DOffFAOA79XbliUSyOCqpmtsa8lO9BBmwQ7SkDWf+WVkvhQj7Bfw2uMK73
CT3M7sJaeSJzRFLz3SZGr9Zg1aZlMOsj+IcZpdCk40cHRwCuHPDZ17TrzOg9RG8j74aOZh0krSk2
ISq+5SV3OIAI8fXkCk6k1Gz4G3yLa6Y5YNrQaMmcwxiYTbMR3SERdbXJj6mwAtxc69hnCpzAmGYz
8PFo8nEwoiBHpXBIKHKScX3VKkGapJkIpssUzT7BzqId3JK7aHAWBQxOiVmHUlpIX8+RT6WLN4tk
/YJGrESWf0ApgEzHTV13cR8sgln/L5EeZhQLilzwuAjIqMDtMNh/i8UaX45QjpohCvoj5J6JvAMa
pqhrzFBcmBurOnDCSO+LR/O3K+3nthlzNwU2+ZXgNzCGPqeDwy7+ANCr78r2KJ6OUIZInEyzgAQ+
icxxIUy5xSQakjx0MCGv/EvsfetuVO77JTaLBQ/tx9o1rVpeltXYsl9MVmB31F5hNlveSe0Ukfg+
4TMZrtcEgF4nQEtHmP3mq3uXFGkpFEEGRWiVg2uSCpM/wn4hLGXZ+VNWb5X8kNx/Dhu73PhMP6pN
YuNOre6kWEpjKbyy7hsTi/R1diWN/KAcbReVjSyHOgO411SxWaOnmyMm8e83ygx+xvkfR8LZWuPD
7z6lL3uQcJa2Ok4VpXlskr+ui4nXAn6fKJVmHPC9cdr6jSCyYNs6wB+Coxlz6zWXCjR2McnnMJ/w
3kBQ5uTHPkOMa2jSuvbNIqQ5P2ACyRkJl9GDUM//hJTEzQMg37mb6IHFCtAVLvI5HZBpRwdGuH5W
WotHz3kxl1za9UaLtKMtnxz+hNtj8DsosAuDJ1jISOkzlew4m92m7Bd0S1U+BkSKJMA9TRmS2BXs
6icbtdwJu3qVINKZHciY+mlbtler2kBT9b+sOUrK8/GNR6ZeHpDcBcYvnSZMqyyf+c//MYHQ3qi2
X4s3ZelHFmjnkSOIwz85frD7UcsoxgyqRbnzdOo1CuvfbnQydtYYbPudrU7V1C6wLaOZx2NfndOK
h/O6sIDNnfOzqI6EXh76ODq/ksJHUxHlxqSn2ZNlYPFGzrnT7QGHg36O02tXUnxmsabZOcFEhq7D
1PmJQJDrwVTorC2p4elpUsxfj4HvPzimExsXrxNr9wcr2Tj6auc9xBXQUcEXoN5aRvNWGpAARlUf
xbh6/NhU/XSKcZ0RxhOvu/+4KeU6P+MKwmAEZbHiPQjDxK+JNUqq7S5T3RGR9sQpudKYJ+Yeqxgl
uw5NVB0EwKd+rfdbyN4NjLpU2yN1fqm9Sfq8pXLnZ/z5zOLy1iNjkNuwy9uqnZTD2bVX2OzJqs/k
YbH8r5fNntcB+ajeUEpeYr+4k0bSp8YmlU4gUd7Na3oMixMrkUx3tFs9hXovNu4/PR25o/W+9LEa
BO9y4IMBdqnoIreRIVcjbfO8pbh6jCPXuJcrOROJc1MKEVLsq7QK9VCZNrUvc1yM7liTwcR9ZvBj
dtUQmBb7cxXEGCojE0EnljmLDTJhpipW2ojXZoc8GzFOTNxifbRWln+6zfibufBnE2Fslg2HcWP/
0p7fljGM1nap3PYkAG+m0Ie+X5JDVCrnhIHQCKI7JmkMvKW7rufo2RNv23JWi7NYKURGF3zSjJE8
AjUfGO2WdCGhdEH5Tq2yrQ8LDdbc4Nix5ms2OUPNPxjYIyWI3Y7vpWbHhS9Yzs3aM4pOq7uJVAuk
PKbvFlfXso8GGe3eh7d4p1O7ypE3NUKTUSOPkJ04BxNAXPE2neBLv/SX2+MKFXa374wBIq9nIfCn
6s/i+GO5Ay4wDggQtxrYmGEYuzNmpKX+pI6HhaLFo6MUjXg/XaIxzYn3d3NPR+EZ2rWvILjdB2AN
KNAf6k97EKXIK9HXSqKGDNqZymZMgi/VC7Z4Hx6boB+zXYlrGQN9tXC2j5dDvP8zoxZkaxDd9JE3
1vYxeUKnQqpAR3d76R9ber/dUVfCM2xdVDOboTOTrmKbDXwPTieTnTIYAGgVosCUPrW8e+0UfWup
uxmi9XhGWk8B9tK1O4HVhcjCkdl7HEyPP+IhJ+hnuneNlsltfN8N++XsUXYdnGRaLsj48gIqhnBI
RA1GBfDFUibaQ7L+Ns9thviVD0KFMNxZFfkFZcknNYtn11COfYxhBIOuP2T+tkCEKOiIk/eXG5fv
RgaRzO2HgWPV+LFcb0A1i+qYUl/hWtB2or319AA8c1weEUvkKUdzK7NoogFIX0cgnYFCd528nIGi
21N24vM36VtOst71hFcVJ1aEuzeBkFl0+9aBWFkMh/DHjpz8iqr8TnRz501AM85tSr/5dV6C5ZSR
2bamACLHuyBhcQPSiKjnJcY3kFpd71rszAPtxPvE9V7hP001fC91VEaV7m/rqhcOtrwtCrCwtwmj
/djMxf3bTH+uJoaYai77GXB7bhsZydxgMeBjHC6ayBheMs6hU8U2xbQ7vXZgKA17EQvT1I1KW9XD
YNYvi8D0thAflPQ+UjqDfjttFtp0gd040or6RYaE0rZYSLJo/2TrQRAGfMVjbiWukM0RmFT4wJtH
304FRcyUzM5ttPDk5ZeBjHApszdKL+X98AC+gsi2cuDpDja76AjGKlyng+RyY68zt3JSEvvEPsi/
UKoEBRRDaxuZV6wEYIrVk0J7/ghVgWdWXAFEFOvBmJfEnnjXkFYyjxLSEflO3msc2cCKauNzMJ5d
y2sGWut65+pa2jzWKT7N+GuGz8gFLqo/S8vazqf8SVITkFnRDiAgrYQECoYlDCj6HjyjDYe9JbRh
sy73WruMB9ijX81Y1uem1ygsGZ592CtHfDN3wam2STxVXLnggVfxdEWOUoVnnrxRsfKzmhmeklys
H26SPGqNlkwb8BbsB7t2bS26Aor9gMrFUrS91Fjds7LKfK45/TbPx1gI3xnH/DGwXhDnqBSJWycb
yJUOu49oA9VS8cbTnX0pVGtHJAddFS6huUi1PRKwtM3wB49aG9Sj+slsmb1/IYDG1l/Mi/8psqn5
a2z+cW4PxhWTCvym5zQr3db929twJtjFeYAgfkvVO2h30X2GVGY9i43UajsP3RvsH+zA8NHLUWaa
qBuXuEP0OfwLHPv8BobkCiXY7tzxJH7koqpmNYVIfrKghA6bC4VhIXSkStDVcGJxD6Osj4IG3vnl
Wsxs5P3W7xAKGNHZZLRgGwbb6p85IcsDD0yCSntvQjhhvINlGxA/lQCsKkHYIUaXDNvyY3S4MAlS
QrWx/RUlBeznuBg9FV+mqG0OAxg7rxbZuixeF7lM/T7IpC4kg5EuDCGgNMJ1KwpZR6AXr2s118nJ
XUgb009XAAkdbCYDD8PciBOpoy4dmc1MfEUrY9f6gwgo7vd2Etk3JsvbqpS+V0OdnbQlFghx8nrQ
waHASuQ2zAiOLEcgo7D5DShl5vX+4ZJzUwebJpSuHcOkyFsGS4xbTGk04eO6c8esVHsQWYYkJ4Zp
uBu01ribcDsb3obYspyy/wDlGVBXCXVGiugLJMovijw4IuMnjuhoO5ubyA1qtvCbLTpNHPO+dbzm
FgQrCiitoq/9KvSQG6JPnlC1eblfI3W3fC+j0Q3UqZqskJLaRtEZVWTR8KnT8y8fMUvxUX/JZrKY
r/LQ29fbYODkXMSXwak0v7KDaSsUbqMsfxyiint1B371C4iUq4U2Iq/OZHddKt3ajYRKqncU1ulL
givRWl892d8TvpN/PTf2Ui/Hj6Rzw7OIk8BZNGQXNSUyR7x/Ljt4V777s+ydtPu5fwL+sC067HHP
LprIzpRxXKxAjIJTxbEhExGqoXlIdrgdNWMWK/ervdIddg6Hu2VQROmUIfZJLmJMcm9jivwMMBJr
OQrlfSttnVHHasibI1AzXX67hkQxoj+oNmaJQpxTV3nLxtffta5NQILfLHp5iF+qP+APtoIcsUoC
4vyaz7R9S2j4OmnoCv+I0oo5FQS5WfGlxeVksr2J9uDiYsC7/F78ooeARTVmy93WOizNkwJtkNFX
/EJ5/wZ4MpWwbJYK8vSCaJNbEntYj0/p4hja1M+sYYhA8On5fpf63Egb6En+a7UnUH7Do/68/cIt
3ajxgSNnr3H/Evcf51hTNpXjNBaRGkQrRPzizuM+/LvEfR/X55h/Ji1fJdgiElrNz0l906ombalm
uQcuB/bwt6p2GpGZ4qehKr8BU3ivly1B1oIzDjVFPLNR982VtY/lxxO/10qVodCk/+N8lMfs+jjz
Y/6rH8IMvdsQypHdW1SmefBh7P4J9SaspAy2AfDB1KhXJ8ny6Ff4DfhNXeheY5WrHY7ACv5vEr6W
AAd61fTSBBBO1ajXrXNLU9j03xho+J0rau6zvLpHkDlrLnciGBrSQ53AiVFQMqRumQCFA5B/Ehjh
mtomMSID27yk/pp0NtUyaj2t7YG5t7zJ+8qYBYwctYDilwX74vXD2enk/4UyBtHXUy+qtPVt+nB7
GkiWdVmWfFiohXaZ6uUxHEUJGPZT8Q60YmanGZwBmRKmOTZbam0Ib3vx3CBtMLLtjbCITFTmliiU
q+wkGrwjyowqK7twYEM+2L2V2m3MjJBgeRPlqbDtZuUGWzstrIMYIujDX0MbveKS3b6xr4t/FUjU
6D8u8/AlMzBFFPkv2FpOYxEmqTBH6y6If+xhpSh3057QxcjHMfCcmTBZAFQkHTEGaax5+iIsd/rE
W+gnElG4jDZIfA5ttOJD3KKpfUResLQ0lJ4XreSud3yRsdSTqCC0/qDLFj0BWY9PfCGg6tODnN2K
Uoh4GweURRXtN4YZXTrF6Xg9+jiKPkdmK5GBTQWxDAzW73dQNWGFMxgp1P1OiYXvAwT3tMoKnHSi
b+N8CsDlQnCzqaAD88sCaEOzqMb3yVAL0u5DOEBgNaPmCNCu+PdJWRoVrVbLLHMKKl44dLvU1D8d
Vnc/5c1JE7sqJdGoL0+7d2wCcgE2LFDjB0GV6PfkN9BWOMuV/sXGSHMOZvaMyJadv1XMkvzvKlIQ
6Rz/ti3WjMoagnVuOrYmnI2DJ53WrYgxJzPLRWfiQPfp9HC1+1TVmjoymqfSm3Ni7q+zkrKTtZD6
LiIte6ucyYdcKNVveU7sg2rU9kl3a6xUPrvn9A0oawHo3qaV6N7hsBUsUvhn6K2SVHHXgb+f/US5
ub4BAX+OGiumRkFr/zf40nkgqyVNcsssaz0D/9F6Y4m4Ysi9Pti+WKvH4P2+2jOv284EW0yToLlU
uaoZayYUC+XNQs7j8R1YlDaa8MFOu7iFgYalBjGR3Vz3YjDcMOFJkibmBzpdpAWSSNZa15wqgYKL
McH+aSz6/ChLKdIVSivVbPh0KjT642ut/uL2Ep6bZangJhK8o7+QGekWwezUFd0m1QjO4AmEElO5
MWV2mvRzihK6KhoFkqMqp/WjAQWzd91TxuYUB/H08Lz/R/hOQ+uthSsO3KdHYPMZjNx02fWQ2vD9
QYNUD9QOB6F6I+yPY11IwqGn3PCBijrx3PsjQnVfprc1CiFSVu3Ump6uOO+VCjj5IfS/uO0lU4SH
TENnJTxFfqswnmxB7PfwcDIGONdZfaFmvB0GGUMYyyIadZkZBNzNCBGeUPx290Ry2H0tfNrZVo2V
9Jv65OXeiI8r4krqowo7tTX0wmR7Cl2D+BlqlIzJRkGd6J6olf48ydrR6n1BXcqrXOblS5tl5s+5
5b4xj8I/yS62kZKPqIkpxTxjP7VFPCSHG5CEUb6/bCVGn2doBEYaLUtDEDYaVrHiiR8/wcXo1Jtd
uGt1yX/PxIakCEEixzh+v1H+th8wARUGrn+HKI5NIkXUJ7MjMmN+fWmxvh1AbW9seQXm/2gfYY/T
9bJhrq6ueNKV8I3YUpEM1lYkyeCN8fRhD5yGqGEia/jQ0A2TbJ+OK4aqJK6vRGiTW32gG7ziCSMA
ZNoyn/GsGmXlRtHzEBzhDJww7jhAqytL1pDQF/k5sWB4lLdOq9N92Gvy+TD21iWTCgjGahB6Xe8H
bMDoeFim+ndgHPJjOxhlLAKuuGzMEsYM/dINJWss/MVUS3BE4W6jXDofKCuWmrsZDtvI60OIXd5I
JrDHnHVrv861kl/N8n20+CP4Z1pXINejmDd8IUCz1SlfTvPcoVDq5OYFBW+yGJzxigTS7vddAknT
EZ0D4CSyn3hL7BiKcloLNpcYo0LHEVEY7f6Ox097ZKxWSzZOFwzP5ugOiDtuAyBc7kjEXyzlcoUO
ENcQw6J7z2zBSQyUyxWamlD/nZLUwevi3KQL7A6NG/a7g0a33ATMo6kXgnirHy4fAbrjhvkx20hv
1/SbwTu6PrDyP14C/Cww7GDIg3uAA+TNjjoBKghYkLDiWcTIvXjuLT8HTxF0C3lfKZvP9m3SX5cc
u98LJBTLzSLtI7pj5HkwNTcO3OPm9FipY3S+ftwEI1YXj31j4itubowQrs/2B+TDjS3/3hO8IbtR
NCfwFl3FHllLCbuKE70m83BzCKGCu6oafRFerQm8vCR+oa4clKqKK4gbjmU2EIpnu1KJ0Y0fBhuG
bv9F0nvXS1vTiN1jxy+f15gWOjICXNtfz3G27589fAwyUZtbwVrl0KNIg9TUaMAz+HXqtZSk8Fin
VL9n9CiF0YvTfpFA8Cvw6uSFMnPYiIk14yOOP4dDnEsag/7RLT8OaxNiGEOWAYqZm+6XUQMpUXhA
mfpG8DEitOvrlafEzc44ETC7Pn9ZewdXMDrwtH+Z4dDGGrAUaKrombxtrbiLjnwb9xD8i9/y/Oi2
Q3dceiKA2rFoAg7cSONc1TeJukwdNxuYOfWJen7Kt0vZw8L0BJe9GBIFQTGZ3LE7crd81a7PUOyP
f5msO01UtUu3ikqy37H/IHKLbXc16ki+/rODD5x5mik1VF/jwSJ7BRXlxFj9Cv7QIIo1xOZKX2Re
kGD9JGZ12qTVYHYBvw8jI1Bd5oJwoXI2bHDg1w5aBli/0ru1ixQh5Vw2kcw2QZBzQxcZPSa1UWWp
WCiVuC9VTvsiI7Oe53yKFiVcxHMxGPP/zGrTubryFEgBvnO6ntYoNUFDJRVAkB6HKxoRVuAq7kLs
lcggkPfdwKo7ai48Mg3fobR1o24imRUFD0F7KBwnOqYr50phghOSHEQ0XPuNnY0jXkNhXjqtG3Lu
5jbrqV7JPEaznY6ra5VMy1vsItQN6T9Zbpr6t4i/NFz8T53NOM91+yLBB6xnIOvuQBi9O4Ih0W44
3VIB7s6NYY9XpMMDaIFByq29uwE5jCu3NIlAMGSMkWiYATqdVVGFl4NeQzcrG9ez0G03/cG4G/y2
WEbwCjCmKqq59GQY99z/i/lJ8P7qgX96Lhm5+yH2bN13RVr1jBGN4oP/gxy+XpnijC0A1MWEqb6y
7MKDMCHFhQ+Ou6XNx87ENyVVG4OaxL1Hl9YNW/O4jDKZfQDk0+oFc3Eb/UJFAGuz8XHO+JkPB22m
AfS3rWoj6I31hnxyJ7MhoC8giw4p9pds1OOBb0dP3/MW2Gks4X2oQ+nFc4GqO7OPnJrMgFAsOE7n
166150K4hVLe32Fw9G4sWVKN+G6BBGdFBTZrS839K4d7P1gfywZz+C8AC5Ue/CNy+/ihWrESctsa
b1QB7jwqKQnF/6hY2UfVZLHPtPlE36xH5R+OoJh83uBV8FUwNoOfd3D3D6t3MMKk3CKtWE/B3pOm
2Fr1jJ5BpzQUc9Fi8nL77bBI+ryscpF1D1UlTQddqKzwClwKdEZeru7mLak+KumQvUasoqDtfE1L
te9Yl+rzopsu47o+9l/xMpasMGoRvoLxaZIYMtUZfQ7eJ0bTvr85VSK5I2jHgvT1dgVRM1mzW602
LkHVVnkS6LWrDmjD9lP53zrk95o+tuLSgqAqR2qbwc1LsGDqc3VQrD5JxIjkPXqriIqUXsgPwLN4
zigMxkNpWrYXJW1rgXbTC1f3hvrWTtdgdlIrdrtCB83LGMA/Xr09e2702Y9e6es02Ewqr6QKZzwM
1NsD7V1E0YPQRzIGDWO8pLEQQDQ2oXzeI3tJQeH58eXuujKXAQA6j9MKTK5GGINw4/cTSyOqnr80
MAs5GelUYldps3DuPkHxcDIAlMKQKm88ZwvHTPK1KUuFBgvCiZ0QO7MHz1NIb3EjjoQVeaSQMpB9
Wu+rMBwKaUkAol/U0Re78LE0kUWJzBlupui3YUvnwu6EZcN4jJtyamst33zY2S3xpOs1rnM1WWmR
BXnwRvW4HNy2/K+jB1b3Dkpo7qqSRm2YVaMpaxO/ZxjWhRy0xt9BZkgHRt58BgJ4ncLyy8P0upc9
We9nM2+ZyskPBR6VWeQVUpFijhJgzPaSwLJgpNUgE3eGq21e75b2tP7L7Vl5eGojKrJKpG9Y5VSb
OuDcx4EcUkXDNAs5BGK9Wq3JhoCOj2dGwS5M6yviD2tnHw7FBob8k5waXCv8KlVPKsDxCkzaihfj
lCo7aoQM4KtqfdCh8J03tZ7Syo50KHSlRBHnJF8dkfngmILMtOd1ksyoRIJn4WWOEc5uI8uhfK6Y
5NaUOr4jbaK4mLnJiRq5pyuOeB5B4BLSHBn80fHocv0Rx1mtSyeVEqNH8IZSTbXeDLaspH9Ge1wb
hlS7tv9vtEW+2CWCYBhDPUPqCtmyC2eCGpNR7GYqvOqj4lCCuBCPzRvzXk60iLWBHpqObGzf80vL
0Qv871xgpP7EVLxmgZa9dJIlUd67URN36P8+AscRAdPcGkg3ZG4OjUp4r/1NzCdxig7l+dE34UQc
MIWhyqSqICBA1DL4r8Nx3BfsXjHNQ0NyhtPMtgJaox1PItljxPKRS5mgkjGSsnMN+naXhTeYiwEZ
E/Gt26v6Kn7lSdBQHDaF2u8rc8+ie/D9nZHu02Qc8Qr2RJ64gIfGXXj+Id0Np83KaxaM2cP5UvqO
aDw2vY18/8dKNgImKWPQuLDwZTgloeMxC9z5jTWiqA2ZMKxmUypafePd4JR1N/N4wn12eWM4Gtq2
SxSJF1NyDBXkn9WdGBeAxkEeAK8VV/tpoYPma/7AjRGkP0iA+6/EAAJ5RQ2Ii2lm23kut2Kb39oi
1a71oWt8hiEjM2Wd/mSRPBReTTbg1ZSqUTAUIUOduyLJ1NoONFZ2mo4KQe9ax1C1i7Z9nI2HyY3f
Zp3pLvie+DWdj6NY5XjlkMSJn97H7BNv7sLHl7NhKjmZU2W2vQWjjr94MFp79hPu2DxFyX+ilGsq
wPaDHHT0gYr+nSk3vCMynByXe4nqaGY8RzAUwcVw189aKrH1NvWZXoZpiCCsTOEkiab0bDfGJL3C
n52GeKcC1PWFvPkUf0t26JrlCmzoHbCedud6owbbrftvqCfMEnkOBEeokOcAYQT/yDwabRxYau4H
Jq1nppjhdpoxaeXSqTkQSRsKcYZ6amnscJJBwgRtUu1GB3qyJxhY0n1sTV0IlKmjL4RQ4eqyzrdo
6hIywPXXmFeZ4KoTwlk5xywXiReWuKRitgjr0dMuvl2eKPyaSWQ3sYTaqmJGeTzKdQtdBHSjLi3j
76DdI7TQp0yW1gPUmwOHbGzDJVSw7/XBjrLByc/xLW+UOWdUc/Rvm2OjCy4GRsQkCripErZg7U/D
3BeXOTnWxRgFeS9f+bYrCBvUTRiiTk3mpHdEJmhpaG8NsWorVBZlcOnPkvTHFE+EUa9jOcvwlYjw
p5oOP685ok2Vi4pSzuaB2NAXB+jIF3fBENN1OzzCKgg/eRUA9cjVU7kaM1vBxAbs1GV3wKbOgD1b
Jc3zKQ1zffGVS66eq+DBuQHPhl/gD3bzavnLyU//AjkVlJ3Vb+jPcwR3uY7JXrssv4P86Ac8yUNQ
mUo2FBTv0o8c9lmIvFRjcX5Be+B5R8gwBUBehVIC1f+a3e6ffZM1MjuY/FCl3wD4TlOd6fzPudEA
NbISKxhJTssjOd1+m+Qv/4xqXx7tr3D41qidF9kWQJTE5mOkKJZ8PSDIidouYuw680iLpw0sjmyh
i/UNMjIMZm1kYm+HTiQgwaSsy+YgNdCrxRNY80uxI0itg0o7eYK7c8NesolsGmf1lxlbBzcxLsZb
WuZOE5drmN8qJVBtdmX4VobleRWNDpjzYdGYybwXBsXMREnBYie6SOpp6G74MVWS0MdHp/1krSMm
T+fzN/Yq5mXjMyG6UuGYpgbqGANcNCSABWNNXBHMypyCAE/dGl8Iw2YrJ1EnCkAU84ffy4+t0WwZ
T5BJ7NR0WS8KN5j5R5KAU7ua9ATKiBIbHfnkJrahEeUF/7d5/Gt4555ahMdv87eQr0WbFfUhFnRI
9RD/jChxjcnFcXTBEf50FfNLPpjIQAYbJo8g4Pqb+A4YtnmBBh/RxefOZFEf/3+RU1FwoyeQduPM
4khG+xynBzHjwSVARWAWmlIgCwyyHqClRn13npZ3hV3JZfRJzuAREevd3QnpL66pesRQmronzUCP
bNbQouYWZEXotqbLtxMncoRINBLMMc7jxTwtpWP/LZ4e1aIMpOiNItc0Vqt3zM6jDryfHE3bcMBy
25IqG1Dc2XyiwjdQNV2pwFhVKnhRcQ+PNMUnL0qOmDMvBscafFgv0HRFg3q+7QXJxdh4Cqzd1eQs
0SEUKM0sdDwstRokk4Y3QSN0rQrav1n5qxqWHmF1L7qrv71Vp9ukPjvCePTWNx8RXGU7hjN4Fdu2
g/d1nnWHiZGB6xudCYOfoS1uDBH6XXiHRqTt2Qk1BamWpnFiFoJnRxlKm2WRv9APL1w+GDAHc8jo
A5TrSoTyDlMy2TeDr3B2TcsNuI+LrE7NyfgxOQrakOkmjDA8j2ZcT3NaU9nCiaIDdDHBgatVTRAe
X48B5oidojqxdgvg31bCVG1tX7gJ8NH1PelgY3XOv2xvVBXbgEPNARf6118DYrWnt9NSRodgpNDw
9zQCAvaztuTg/gziSXZ4sEcLDeMWIDbDdAu0gnHVi4drK1dBqVoIpwOk5Kj6tofWlsElCkhwDKNd
UzO6AmOzS1ON4XqIYPggVErtmhnmKFDZI/dPIVRrFGNZ+YrDYBKzw8BqcLpjmpZ13HiAnWYct1T7
r/wJS0NySKvi1FjOrPaHxefKFWQBCgSOSX02oWxPkd424SiHBs74AUD8ekTJ7FlbOVr0hKuU2+xN
cifPQyGgUboymz4wDavCjswk9DP6ol9/koozFfj/PMqTGWi8bLU2Wwgnm9j9edKdKsEqLbJXXU/r
BCJlVAvdaRNwI9qakmvKBfjyANJxQvylVeQ53FDBRLcIhPqG/Q0OdVTADRUPHANR8CAiQNzAcWwB
7ZECdjdFL2rdP2Jb+AyDLtsga8KK01vGP3G0sITZNd/BfOh7QtqH9vEEUIsZuC5cZFGUoasm9kVG
XQ1qdz4mn7M5QwiwevQVj/+rDysoz3faG0bzCWsJVgDR/3MZpn0O8AxZ0Cc0GSiHkazcNpVB+8ld
SK6UMk+GLv2kvWux908e6D2td7ScnzTb1GUwoX40w3h02o27LajxSBGui/9hTYDLzfSHaPDMYMn3
wk4t4xxqYCcJ+COC9mfIxifNhlzuaRzm86niPI0ZvwW46MBR+wrcBW0te3KHZC52ERG3wfoCif4N
f6f3e8xufPjwx6fcHjm1uzA/pCwTxbxs0RfGE3I5/5paOerHfCp3RI/6U68IWaPDmAjvbd/mGbYo
TopWT9HTfIAiPesmypiLYD86vX2Dj230N3IcjhHdtZmzhG8nC6xNOJodDWdhu6EaWeRNkjwLXYi6
BFOXqwoFc7War9N1HapE/XjVus3zWjE5wRlPY4vSDofBxeCTE9nCtc6uACRG1XezaM7kvSIttiTh
MHxKu9PaIDGbbfLcB5aJeSoRp9rL6lknZpuCq9vlRL1spNFP7duVFbduuol/OCbbLQ/2+BzaF4IA
h4ZdeVaJxb9tqgfucr9lPV7YqeoDA/WxovQkfIu6gJKiqDEZ8eP2CFfzA+v5bRG8GuC0tAc3Fe7B
fp8JE48wJBF7BWeEFDf/kTpUF7YKJrDwv5PI3JIsmOhuuPCLb/cmPrPSi/jHsWi8548tLcd4Hsaq
1ewKKpxZ1OgczVolCOJgSITSNGmr6Dyg4nDSM66al3UaJtVdrAIqWIS4lxsuDsQ5kBQ2h+LY6ASC
sn/5uqaFHBuHLkFV/EyW7OODo5oDO3nsC6uweI3rAm+BOQoMhKthG95yzbu716uW3fm1Ur0y9Afe
ri12p2e5+vmsoFAwuiG3AbBLuvwoBL6ISTOqReHbrhiUe5yP/BpdHLIhYWRPMkMH8jUnmCtK4eTU
ZYjvCI8vmDYQldvjkXDwRJgjBvBCZvySUhrgyJe63bZ3F3pYxrfhTPFfP6NWff3309C3lwrWGY5S
kdiNxMhck15gPjW2xWm+tN7FodfmOAR1iLiYQ7x2mxs9FhBTzFhD7+Q4Qye3lZttVAWXclHsdc8l
WjzFUR6bJ022fzva3kTR0XGjxL/kZpYwIJ0k4tsEklh1n7der2P/zi9nwBcBBWRKwC2nl0+56BcF
kvjq4VQC54AGBUdp3OBEoyKWU+VTANIkRaMiDl7JkzO4wDzjBC5c/K62toSdeRLD3VQYxMta91EF
OKe92SjeMT7N0WtCIjxdcjGqKu2a0/gtKyVsPUywtxzsErxxS9sygLc9h8ebWdiwIKBXj+spdE3x
Nlu5p9KtLf3TRvNGDFapeRLYmkEd72L7uxYzbAAwTAnmniZ8yjb+EWya/4wjXFmnM5jmnFMVomjU
XKL3lrURlHNvt4T3TMn8w025iuRIn9DGiLGbc+UVJSVcKAMp49MCEMxyCPLjKhRZh4c69Sita8dX
KORsMkuo0gv+w9kX9YWJvGB9t7+a+uoGKsn/87Lbcnw/60kJ7FBmw7ieSCvCZI8XtIwA5LYO/NCZ
Vr7g3359ouZYlUhT7PJdf9osaLuvdenCOL3lA1U6kNVqm8EEQ7UpjCl+NY19lybEKLUhdK1e8ZZD
XHZJW46T9V+rUt8C7m4LRte+PXKVqxHOlZ2kt6+B1wcgIQQMNJioBWizY5tx6E7czAqXT7XjAX3r
ioVmIUr6of9q5BJBWOZPiI7yLvIpnN8fLGeg9jyNUvuFWc6SRnBt5PVTES/DD2MSC7H56MgUn8ow
qZqtPe7JHWDTtSVo3xHZr5LHSKYC6aN5IHYIZiT5S+m4Hr/HgnNHlJLviuctEpbQ4dW4xKk0Bzjk
H3G0S3pyUP2lEEyLNzlk2s1FZzfQw19cyg2njN+zhrSQ5z2QLRHzO1PIbwkQKlEj5UHjTth3x6RE
3BrKXD+dusmc0qs6+CUy8sLoWLEWHC3QzjLlI4LumT7ypUfAyTvZp2U3j+8o6lYwDMHt4KqtNVTR
ZHcQFDaJrsl6KMvoCrBs1LvT9XMsskWYv0ioJlqbvsEfshCGK0GTlsZOLZTZdlYxLizlEKiBmOLG
idqukRAfMxRm9FRLtOBSq/1kw5Wv3xXJVsBkxNS6qn2xIqdPR8JJQcjTEYoYvXo/k8+q+OycefTb
1QRa9HxY9XHY1obHqte6OUtI+GUa5WtACL9AD7q+Z19krgqxzXa9DSr7JdxTI9dqHQdQZRRwq0bY
xOvPu4rV+IcTEjYO3IN+QpLGdlWIWxDSyO3rBF0LIlxBI5cRwA/fAbTuV1uuLiB5aRBalJlOYtCI
bc9JvLrc8B0qdTJ7p+z3Gugt1EDP26OrawaGixCT8+dNy2V8+PsMThqsv3yuNK3FwY+EH7fIP92I
jsNslzb6POuOjSbEC5Cr87urvxGXSbtLimlLBf8uKN2ajurOqOKXxD+pWGkyVoGQRhN6JtjtQ5He
KAtDVANMhmFDEtFl4z5od3VK+9qB9oyWV5ExVZ9K/FGY0fKv6UXx4N7ZNLdLIqpu0RZdM5CU+LCx
HuZxishjrm6lepcUi5mQ63pOOWDljTU0HLxV46jAMIAct33BMLjH10FeSHMpjENlE5D66ZakjSby
PYDTh1flYij7TJcW5rfW3QmBqjIW6JHWFm+HnhYrBqClqWuKRgtuAP4hjU273yN4wiIBD9EcNfRf
RGDm3UbuggL8xiB03sq8O8PouoHfoGxfvnc2prPxXxe94Nm3Y1wTyToiJgtFBwK4p/LhQGvsD7+M
bqpJDz0OMx6P3NvNdAc1bapvOzIMplQTjenLu2WmCfOJeMGmGzuPJibK4GAy2DfdwGAygY+P0jlU
RiUWlYcGOo6kfZ2VS0RNY/pht0xYu7z4tNRaEtkgBDXW0b41NKVsF6EVH0uujkF9wy+x2M+BoNXh
ZezDxqdCA1e0+lq4uMz4bKmkZAARd97PeIYI1xwLWRCiOg6ViiwtNfDJEJHO8G74maff5U8c6G2/
ftRU/hcmVP2zNlua7TrxXGluJgsI3u4owhBE41E7Ka8TjUmesIS38/37ukZERjNYfKCvK1R+U9n9
qr4VZYKLx9KZSOc3wkvkHmuGX2AmUgt9xCp0x8eXjJpuV0t1WC43p/2y5HSUe2JnBedlD9bbUhnw
mnBZOKZQTm51lNV821jz2sr+IhbA0m4kZOcdR3AggqM2r6Q30nA9pfzr9/XCcUwhnqv7w7L9sbKp
8PnFnFOISSUtHUh0kq4LX6grjTGvoHtAFTtJ7+1UG/B9dImw5r0NWYVZkxlp1NM3ugZT9BvuoXke
yXe+SV3rWAT01vf4VSDBpz59BP93p1vaze7u+TTFIfpxJU4RUFSJG1u1MDTSHalYhp7jJrVYWe+Z
YbZYhfmBysfOoq3EJ/KZtq068e/UV5ubqPlwUpo1jxpoFO5HW77nc51lze/thk/yJ1rTcZbAX0Uw
Izjzc3ZSzg5JDCdzIgt4dup/Z1M/If8CpYL3+4UHsI40oYL0ckiJjcYfoXgeTEEH1BTIfraeX7q5
i/aJFo6cOZrzpJSVZt3Pumikqaonh3g6S7rYnPNqapQMLl0MMsQ2SWF91vzAx8jJWj4NGud3KU5S
apYeZLIYEBk6C3L40+7UctU/BohmmhyHRQcoYCFA9pcsopzmfmyuvtwC5s3cbNphdcapWJLvh7jo
dVNB0B2o3iip6kKTnBZT9EC7wyDdS5W2D/aLQihad0nmwRJI2X0NqCMoRNSRge1k0tEmXhAZT9/e
eQPe9zfQ+PfPmAx7rN3bRukneCFWtOOBkXEdKrstaqKXUTpss40b6WEPU2e+u/A8phCBHr6ZsOXT
7x/6SoW01lmN6wQtn7d6AGaTXWPiPtWfF/TnvJERulKunIEGmgEXx2QTDIMEjQ7kNCGsay7rOP2x
auiU9FdTpnmvNb/Rz9wikBqi4nZ36PwhTSFqwj72JlMQEDkzGJsO9STr6cK9CLX03altuTfZUOjS
Rp9HOKxLAcWFeGJVZKykHFGZ3/md7ez+DsNw1U4QQqXYsO7tpLp810/jWfckvwicHHhADd5XRvOE
kcZxVMpZyVj6z9taUw6eomUN5WrgCdEOUauKYWOWEc7l8uXsTMSoH8I7+KgVTJsd9EfapXdUg/vx
FAapb/b8ntYo38pL4r2XbMMPrGz+X3bPDqru4Fli5rdWIXiMzkg5HC/4CZM5Jc/jF/2CbjqhWrQf
ko2vUP9AryYZqy3hSL0JSa2zKL51U9vWyW9abqZUZqRXqbI2ljmP+q0if4lpY+/b+OoFu5sMr7nq
vaP+uCeJMqVB6PxJ2jajLlsLXjXqSiKXV8iKy4yBDfITZGUL8sBTkshk6T/KG9WizO0hN9LpT77W
lXTnkalJZGCr91tR8zCVw3jVAoN+qUWlPN3/JbPNDBvn+DIqjCxrOqTCLebDvbRIlxnSckNk1/Do
Lu3O2lNGyTya9QDnkQKgPD7c8Uu0S5mm3b4jOskXQIX/X5p70VoJLw+PcwiByE48cG0hbcBgowRk
CCPSTGepZ6QilrI5qkAjc2VoFE5rpFR7f3u3P9n/yX2YHNGQ9hsUyAOh4BOMp6t0z87yyG5rvfB1
ISJLP/VT7BrN55baIvMRd4nYb/0GtrbDBUT+jisAC2gu+0MQkZ53xANNyzyQoT5b3awtqHhVkjZo
X3mM9n8J5ZNhPrrg83cu2YgXAe+PQnIA/wy8MT4LsLqnh9ZfSvPQCscr8PA4Na2UKgpYjZD1Lu7T
irEP+Y05sbKdFCOE1Ug6UIoq6tVzm52bFWZXtlCah6nMOG4kcO8YK85yki5/w/RcJ8hAiOrR3IJP
MtdWJZ8hrpjT9CDeUjQ6Xb83mhOmHPdc6+5DLCGQyr9OkRVj03LkmoRoGktIcCcenKVUav1xV945
EUHibrjufWExVgzSypYWKYa9YAPpaighc/7b3lgSB0vOVrMvfKX8QgwiuSTc03MiBW8wv+liolSl
cIPTbhV06vfa6rBRCCJMATP9wmp1aSQRSPExohg2qKEqHA2FaRuzJCIkLqvrgI7Ai9JQ4wiVldkj
WW188iYvyrh1LjaKrCNjybbzoOvhsgKXCsuKHbEOVj2fZUKGP6SrUjfzJ4utyzw3+imb7PKu4NFY
pHcy8IwBLKayybXIiRuZTqTkRpwZYofNByPjFnSuowkBuKy6iysg4K3zFmaYfrhJwDga25YWFH5b
fyvtpEptdWzI7auRMIuUHNC9DkPAhIihWFIi/9ALWOsKx4WxqySx3sy6qYaqum+zEwzTfComLDLl
BXBiROckKakQsOT2DfbDCVnR7iFuJAS3IcSlY/oHuBgnkVpk1qBvbyBoa6NHm5GY6D2cgK62GhC7
kHbQ+1PTO0nV/lwi+tWLxb9+/O8XmOMaRrbTCve5WEnL7iANJ3oIFRPGYVSoRcVT7K0SA5g2AvjN
yOzAASwKHtG03ZWl4hcrTGcDfZx7psKrJ8q4NS5OD7JzhJLepquQ+OlgTf4Mzpqp0orWK3cN/v5X
TgzBOPEHzpNKiG1ymm4Renpeaxg7WGVl1KdGgiQ54fMyenCs6uvweGA1T1iGLeeuQIZpmrEhL48F
r6sgCbDQWRJgq4P76Q8QDKnvpja0OQof86W9YYYr3uo08Q9kdCYU6cc1N1Fr/HepFdPymp5NXUdy
r7dDgHbZRe7mXGYpE2th4EqncczuKfaLo66PceXII9s5MHJNH9kBT//rQ3XwSwNBwRNM3uod85fS
WFYA4yLXVP2+q+bgg/p/LrRNzhXQTJTOzfrmwPFrE+egcntU9p/Af1ZWX23pgOd5ku3WUdDQDMUq
UGforOtjkPiv7Ts9OCy9Q3tkx8D518GbMfqG5FRAtH2ww50Pnyk0CtujrjRZUQNUGD3FT3tHC7p1
a4RbaxWsDPdp8ZZsEyL0cukEOvEt0XxIS3o49MeJ03NSsFIdIRiBxT5arkGvAre+NaPAFYUTuDaW
k9PIvn/0pgMqVjQnNHhXaNgf154vi+sp3tc0TmB7NMIimPTg6W8utTWBhl80lqgRkWvdWlPCN9UM
xvumzQymVQXcLBpodoHVAQwu2asvjhIrDKUgJ7t79sc+lwv9As6Gx/h4Q21l3DEfQEC2Iz1QgZJC
kZ6zgZvtshL2nTFInl27O0ga/qwBRURkMpj7Oo0aRcoCNbmpPuyyJbq5E2V+jkjlKdlfQcT46rOP
K0kFNTEvnUb8V1shgyZLdjthh6SY9vSQ3oSQ7eZQFHRC4t0IeG2CawPJvAujQsC6Anzg+XiyIaCX
VKhHpKVRUQdDDkwVruDZIXQ7i5UqzDv1Xlu52qnaUC5ICB1TP0PNKOsIsTNFlCLL15uj5/UlBaat
K5PFe682IYKsUR60Rc28q3tnFZsivmX0p88NfqeV91novFU4Aff6InNY1/RB6NcMCjEbEsAQptCL
7l8z3Ay4XEalf8XwoPqmOdA1mRX/J5JNxdnG+Kz9ZDQCi45Clv3nIPGM1eWgA8JRpp4/LE2BqNEr
pI7t1vzdJW5fTweVxtaNI2XPA3NKABubeW0DXP+zOJw78fQFOChdS+AIbx024sf226gwDY2ZbXsp
p5EjdD4jE8SzBn8NXO+j3+OT2c87Mm/ipViGT0r6ZQV2Pg/BSlhIloulZGRcBNbY+tQ7iWwFiYXs
rrLbNmZSNuqqBTaSSqIPRDwdUFEc2xFYsCpsoMRsqCKLPQKT+T8Zq2dd1SXp7Iy7KhFfsc/38DM9
kTxaOttY1JkwlX/7SOKa3Xv1z5GIE+2dHgcvsbhRgXvobUE4DHSTASXuKkTGDaI/mKe/BtqKQA8R
Hil9AR5GejZg2WOjdS6YTbWqHJ2c+baW6J+94s6lnzfCuqv6DVpmEJ+uqCoTxkTTfQKq6sWiTpoO
lGEZoN0ScD3GiI6gQdwO1VDmpj1rhkRKc0ogs5gyAeAbfByci+2+cP0E48jQT3dMz1Q5DvulYtIQ
599s2xJTFzkEsA53t9fORaYoy8eIBEX1rSf70tvgV0P36JxY9h2rU9sp5wFmb2I+YWANmJfNEQ/Y
udUObTJ1GzhUuVxai4u8AVrFo7OXYTNHoKmGUmLf3MQbwOGMcuGbxqwCUJSOCRC9Au+yUbot37IV
jW3hg4k6rPFzQjcj4I+OjMTfcd1JzdNUqfKbepUIAT1+RNItoh/UZTEK0u5toyM6JlZEtnvAZ73G
XV/YH3VuVt1LNdLO0869EPazXeUPDrd9FHnWU7EBTgLJK1HQnfbWeNWzY/39WYZo1ReoNoCYve8g
EXA6JtWGfjbTHJyoEca3x6qVUPs/zqI/67uSaTuKR7ckAscn37N8Agxu1vhtw/XEdEbYGDIFKXu2
zAAPDx8PhKcOQ5upBYPe4YcO8GIZXlSqDbRWV8c1GIlrJ3RWXjYi8CMqmPYRsQEjoD1uCf+STmjv
lFDUpi4g8zsYhaF6ZmKYkFuC/6qd4G7OJgUf5fB3eSV5kMK9faufSiLFno2ouIcIJ1Vdu2mt8jff
jPDudptHXD35vsMIVCFpOYWyGHNK4tITu3J8qKcy9wUHH8Eg6Ob4tUepSIGqSPnbFO/hrSN4An0q
WX9dZe9q1h7i5YDT7+NZCiZYCjNSEKcJHKfqU3e4rB2BA105wVhI5SYL5faakax18Nht4IsYuYHm
A4ATiGfjHHW3BRZMzTEfDPxQy/5oD3Jl5Dj3p28sv24cOv7TXL6dJ7ySmZJEAIjK+EtNul5WFF4G
MiyCk33yUAWU7Q79Hi82Da01Y0eDW52a/GguG8drmhbI6gFlQBGlzDNXNY+yNk8UIvmUlUrjXKP1
iiuGWyRFkndsS48Lzo3q259u+UmpcC9V8VMG29jEJhY77GloVNmgdfXgn+GFUp2bGWRYTOMOj9qu
r3yFK2o0xiXUgv86lg7JYQuSwuZ99Fs5DXMEqvNC4NmY71mIJOgSeXbyVVb0YMYtdUjavPRjCOcQ
6M31yyWBddtWsf5rUISdHJnP7L3tb0/yeJ7MM/OoJ2PmIB4sjTEYB1wfkODe6Xaa9QEWdR0CIQ5i
A8MJav4/RdGY/rWfGc70HjdSqpNKS8sjiuF24BnpacQYUZkIZb34Y8Tz0Y7uDImXBd0cgh7p6Mxt
Dd9n5kgUTlX5/jrzR1WWCKZfd5SnIpPxD2OqezTsuIQOMU8zmf23VWIMFPqFamM2TNmWDhcA1yvm
yQ+2/eAenVyiwZstC/mXY9JzEmciPrH2bjyP0Qa9ECAii/ZMsZ5EcTAGGIZN0Ck+/ewdI+oSufue
Wsr0DW0uLFEbsMyWsC8oBs4ttTnsg/038tZDF2LLPTtnb+O/eBo8gAoOq2nopxpNYkCwnwcDylts
kWk+hqqdhYGdqgKpKk/MXwzVHkjxBJHoJ49qTaY1IV7m9xLAs9u6oxEN6zX3T/CXztXr34QPz4Fj
DPn3lYCxh0wbx7Z6AoisGfrS+xkPjS8O5yDSU3coQMPx9uMzq71UL1ZrkDRD0H5FBDElczpTAon4
TkTg9FnMuDEh+2JL5U02KK9RMfAu/KyyFGotAMRNLlF1IfRudSVuQvBNycJBJxBWSn9ntgHNoUnz
RD+hJSGInTVzhiyO99d0lQ4dQMmhqKX+HxkqT64FEGQHUY3y+Q0GOk5XWMxYguqlstQjbI15WqGd
i2186pkBIG3ZSGWQzQKCgkgDHFbFYLPFMT0OoA+3wvIhGF2//PmvAPXHfit1SJDqUSNXXr9NPpXk
mWWxbDuFKogZA5IyUN7foEPgZxC1vL24+XDgMNjKl8JHKCIprLIMRXoxMmzlDdlUQ5GJDAeGu0WP
FtApiCfCxMl+rIgd0NxrtU3A78X5yGzzj1a70crqOdxpWy2q83ENZlsct0+7EZaEI/7MDSS2qUqM
9/LRU4lFuLHpfFrlkD0PtE6kpCT9c1UtVnH1j+2iY1mueWHv6tF6DXAZfcuu/y8WhcxFrG2PoV7/
/OXJIK2Ve4t5F+GpA7/I6e+NeZpvrZ6rhzY9MEgSPHDQPM/U/M3FPV2Ik+jFB03+KuLH2poiGePx
zhQpzloo8Qz8Z/B+xP6tRJhTGyXJCb5xVhGV7OTduDro2vmXnOYzqjfGJsRgau7lPi2ddsxhSP1U
poc96OYv+GztrfxoYjiPxV6FCbjyO+IhFO4jg3fQ5OJK1Fy6XxczmiJWWs5j3gxvwSCrEZLXGZar
s6jKeUe1zCfXoBg2+JYBs/aQjZratWwF2XWi9obE0sxXIkUcS48BVSAL7uf9NxMPkRfx41bEZPzJ
Hz0bLt/c37J47FfpejDx/qEXCJ2rV3w1T2fWgL7fIPNOqe7dOGi7ARz5GdD0RP+05uHVeCUs85qE
zvNNaWt97d0EYoAUcHCBnzCjL/cEI1uOBHNsp8Z7qwX1eJsv93jaYq1cTbL89c6i1D3CV5Fb/kPD
QNdBw25uyTC2X5yN0OD1pk77yd07TR6SDFQ74Znpi3jq407/eEAtsPW3bhANY3rQ6A+gzXss/fhj
3l1aVApnEPLttL0vS0Nc6nAWItdQOSoqw3AvaU2JU5CRHZ/w1Ezhn92AZOmtRg/2TxgLdv8VPjjQ
kzVoFC36hg6D/3KR8T4tUSFPX1+WwMMc39GK04pKbnj/+shUDRARgSJFhPW00V2tvwGREf6nTM2M
RW5KzC+OenxNNND2v6D6qagyG2jz3ViW6POszbfJjqta4+nNX42tQ7UTXFCMMRjihntl1sOhGcQj
KKBxeCIi7vTYpzNBIBYTLoCvxoKfiux10/XSfetpJnoo8n2/PYAaFTKWprAa5kMHJHZFoOnKvXS+
vNZHSO62QJgOCf55Th46nAZQNoNWbkDIQE2lAi/NomWcXUAUVncgpBVhAIr9yOxLguHwUNDklefk
il3c+Doi7XChxtbfz0HRCirgsLcaVK6nPiuVfo72lol0cnZYSgu7uyDl/R0hc4zyYWXrAvWUKdK8
ozzHooZGdo/2Q9yinK3Rav+wIMCsV1lXlcEOFvASIrQbFaACev8nOThGXB3co25hQ9fL8IcEo8MM
tbWFNRZTdlEVaULokCIEt/SwVaV+jojzdKXll/ausyq4lZY0kT/OPCu0hvWHj48+EsXygsyElT7I
OBt+7ZQi6R6a4HKI7+X7sEPzxV4a6hP7diZCWYzHRnGnYInOTtLonAqmUNR+vLlG2imN4G/1gSlj
4hzlMaU70a6Ig8M/ub6xJvnQsVG1sUw1kqjW486iuUdX7afdNiJT+x3cZ0PbmLRF5/sb3CvJUvuT
GonlP1GkRL0joisnDylmyNYrdOQdQG9jIaviJ6o0GTPTS3N1fNjAYqmXBImQ9ooryDDNMmyvGjK5
HEHVW0/dXoHwBYYwRcG1Np+4AYrcxDVanVRKf/r/vC0wnGCT3IzBv4YvLp9Qp9tR/+ZoYLWqIi8V
V2Fn2klFsJK84ObPB71B6kQUtXKFsWpQglSeyteRTgYymFiCuzVsGCyVukvWX9xCgGf3BVJynUUu
Rpl83Neq3slQEDTH1xU4lwNSPhJGp0kevO1taSHPZkifT5zIxh/WgDM+L7uTaxQUOsXU4J7MJk1/
n4lnLICiNjPI9zvpSqF37Un7oghH2TXOuhF490c7DRhRFZbwn9ykDUO+7+h+jRc+dbVTa4b1bVlK
4gE9oV6SBQVWUZ2OKd6F6ESpabHpERxM2N3iipdxqDZOJzzdGLy00JI1jXWKkgKQsVczVU/VN24H
gBaOwkNjBHFuxU9Ku9Qwr2wx5KDo7txqaY/o9MIEpQt/Z9tUpkiD3q9jNG2WMQWLL0XtD3uXPExN
fM9+KaNGfsFxeRe+fyen9tBivmAYBj/X/mZdt7Q9Zt8x4CWd3NpcVbneoZX2oFCYJAzT183xR7T7
oF2awdbc1RVJFR0NPruWEadLZr5OmK2jFLVWTISbMAnzv5MY6gIt1oTWUue8quaTvxsjXaZKejDn
NZ+abkSStX0JnvSYYSdSXs8t1ODrITw/iVUGjPGJ66gpdmBYMmhYfzW/0djeS3wO3JbNJKF1OCIN
5HxPFh289Q1z1gZFvu0AmcAGjshfK8O++kvzXE1Q3LfLjZUu6T61HueOh7sWNp6FJk3gjbNrdaTC
jglwK8Caf+jWBtdgH9/yEWsc+Lc7lvp0eoyXwKjZEW6XC0MqqLfJf4d7FnJA5TphtNAFrqEvCy8G
aXlPKsqdkHTKZwoErGZlBMOYt7j+ispcFEwNG3R25lS2mJnq2lsijCZG4mSK8uu8n9zVDiAKl/Mg
MK4NDqPl0WvTebpYX1li+qE1ApqVUAZgXE9GPRH3b1NlfdkOHuaa93bOx+g+O49HH13uP80c6z9+
fHd8hVT2OIMeDp5hDBF3pTD0jAa+93cF45PlUPEhySMmrIuQo8Xqk3KK9erGKvjP60+8pujczWxo
40CP7Td0bPctdHtBA+HrkR/7+uP6+KrW7y5jS97vQL4dBWpB+hUFxfcO+VQmh+AkhKPogTPtiMnG
R3tUumG5BpjZfkLFNgizWs2Ul/4iaJ38T+QIOQJogMCzyMIFFPJuOeN3/z8fvLJLsdlcqNbBHvbd
qgFDOjUeZ7hfU2HjkYy0cMlQVGhvD3VH1/IUKgGHJ86w8c4RCjDj9FVhYM91lcJBjsHTq/mYUT/3
QhIF2jeLI/DKSx/QLYCosYBf5lC864MK5IG2ONM4KdTWdUW5ovTM2zivkZal+aQSa72gkAJFSbiw
b0Bc6yyggV1y/HmB1K3fkppOpoctmiOjNJ59aeqrGM5w35Q9BX1/tnFshLW7mu+c6biLP+3LjFav
Z6+CjIUCQ+YIo7quHM34EaEegKOvjEbQfg6pUEiZcHVgX1+YYZLT8OTq+eGPTSTQxhGKh31YbuSW
pdizEsd8iK932awNf3f8A4xEIESSjnKkB8BXL8noTwdVtNFOqPQ/uTxWwNGee6NEluPyItIstDPI
wynU9WlJOuZBe31Sc1N3zhIwFYvPQNCFc5yu9gidGwr3tjAd3DmJkEyWm4hI2g4TJyG+I2f9UaBz
DipdNS4XECIgsbMV2zTyfrJmaJyba7d4MhyQwAvsYCJVl3n61sxdd4pTK0buOHAN0hFNXFHrRI3O
xKaWCzCBs7TH5PKXtbNW8X7X67wTrp2YvSH8EFzIu27lvt5k0BjjN+V1EJQ/jzFQLd1+fDNswPfR
GRzkCdBinJBRiZNprU8Sc1ScnBHy/i8dnMIQcMv74A4aj+B6A1EQl18uFEsdN77YzSuepoq4WCju
mDoWU90WVVBIjhHm/vYs9ip7blEW2/Cqu3D/Sze3RrCxkrbch+B7JhU9hlmDWE6QgKK/lTIRq1tL
F4zk3aGgGuvStaz+mdAIuLLcYtTEpr+lLU5mRmKp4t8zhY1/sJeyqX3/C71hj8bPAuVWFTnwx/wM
E4/EMdpU+YMqOFNxtyo2ZFmYBF/Uc6N3rk4//XLB3H6a0YiXos7CqJKIAulC2R7da1J/bQ6xXiRB
7cRIkFuZHcdUr+fqKQfvDH3kVT1vpOTvfhs8a0Ua9oFGJaCHBh7ivIwgUgpB8HblINNUgCVQcFyu
AzSR/korW+z89mTuijABmFTj2AX18BwUdq0Zm7N5LRLqFCiDCCyGH93FPnM4Ii5Bip+QM8u8ifpr
JRdnTQEYhBOxWToMU2aoqw14YNLwnBNfc2RxCpAeiZcv0pxikMInF74ts9sGkUw5IjRjbEgv/oPA
b4V3vmRUmdTQDL/om6n6V2M3gIYMiCwp/anQyQGLtcwVI0LK/zpHpP/gPESQYf1wbcmJ91AZuPHX
TGYXQrOUCPCRqLD8uytr5g3yl8BXckQ1ZCIcGSkbjCb88CJlgekZKaHs0B1gaAwlei5rC9I2e4qZ
2HEZANo1rrR0MEoCsMC0TXI9BO2Z+190bhKc3LOG3DbNkz/V1iASNNIiJHSqQ3A5EzXhHfXZS2Kg
v5TNN6XAQ9/M9i8jxkVyeRSSUA4i+RoChOuuxd6xB+Nry8mAPXuIVQRWV/IJkpihDnWLmWg+HVZL
815RmsUMHkSs6bufia/nkMRbP2aqkkCbdsMTe3wQPoWcEv7y3xpIURLp8N/UV3NeYjygILIC7vlb
cG1mPDc4m2AtWymlnGiqdh52+pARmJJuGvVj+8TZniM4FyH3G2U3gjEeJogdY3NgSfn+saC69WQf
DO4V/ywyJ+kWqsChHw91NHntlip62zG5la8+J0vnZTL9enSFQEDL3qMmSr7zK28sFuRJiAipK28x
e9QMRMpeOviJyufl+z1ezjz/8ehhMfh6elyaIZdkEl/G+s4IDZo6hVSiRSXh0AvLdEbdOS4u+O0S
KyOxJ5uQiNKYZsOIWeRgwo9H3/dDJeoR4dGSgQLN6uLEixtqcfeTKzbEKjQXwywBOznoh3uZeRCn
jqqlRMxbPh7mwtK6uRmXg/smP0zKbt0jDBpyiuXmsft2N0aPDCEnnxONS3oEz53zgoHxUimyA6XY
zg6E+3oBId2msm8yjkl4ZQxHfUQ8DzN2BBfqNAsd5lnwC+M27pwYKUfjAlVP72dEKEHW3ULyi1Yc
nZYfd0rzLi/oAZdNjZMNiFiLURZh9LBdn3twzdmBSRhpjvIcs2pI3s4iXmX9FCH/bdKcYRLZUYM8
7Nrfbpg3kAlcAo4+F3EL9FTTEl2g2xFDIHrM4ySmz6vFu3usz9QqxcmtcvyyT42V8uGFtcarp66h
yCcDtubEKO7a8huY0PVC1cMTvTQRTl00lkpDtcCZyCcFDRJBd/oOEuP/s3wjihvZDzeV1znREai1
YDFaDdnUWv0s5Rv4VlZDU4PRZ0US/GJv+xQ0rQtec1fuie8UmxqLvHSCbEhnhTxjH4kZG6nQB2aG
hsVMTr7zhg48X2uBVk0OacqRmA11L+nLZ1lRQ5jZ3paZZ++iOwiDRNm+FOVixhdCYHxCTV4uHZ1J
CBkC1m3kA1K+ywGujoS0mwuhy7EE7syEePWqEP6fmdm4wnxEXPbA+b0FdHMoH98sBbAXELuaMLes
yfXDu2qyxLp2EI5M0IOX8kBiQPnQ30T2qqxs8omlFtbfNRb+hWvY1WxcHsR2Y1Mtjotx2xsvAK+E
FGh4h7fAo1mdhfjeYjADC65JwiJlgGeY1740QIkkwkrsT/Am0lXKlCQIf9w4W9kDfPO01LI/kDSU
PBhm3ba+rlPFB5jEoQhGrNwExvPW+K4IOyBx11utDf8Qn7eoaNr4JPwsxGmav9dzbKLrrJ30uSph
NNDBDA25oX5wMlPMlFGxZ8e6YZamB8ZXkA36k9/1hu9gl0lWGRwWsi9lR06qg5zJwiWX8KsppKFM
PZjm2fRRAEl0uMfKmEA3rWNSRZ3myF/WMZ4ZPjpEZU8tHbeiZ3pbh7mRocdbHKFnTTitpMmvppj6
969JKgVo76HhQEkXYm8lUNkA0VO6kFmEdPgREdChbvl/ih9CETkW7muJJw8ZQrcjo6XiQCqGTSnN
gXbE7m2WFnZqpYyvDDMjGsRytmladQA/zx4t9kVBBhW/AusdrqEOBifMYx376rp04C+o4923B09f
VaQGatKd7TFotnXDHcIICALsj4Z8c+xgcdKjOjt85xf11r+G9iSO1NAekfyRp5uEaM2UbsFla2tD
KILnJjnFpzyy6uojNiJCy0pGC0Pn8yx3NQzg/a9vkHAhy3cUHDLJmp1bbVS3MZoLXOyDO/3b4DTd
WO+htfmj/iVfqKEthd5ui4XolsBpcm4gOFimBoCWqdmmV/yzK3a3rN52NDgsd890LIl20msOH4X6
rj+bkj8aT2EIYGipk2xPIr6u9f00QkmHQFlo4Jw6awx88unrKblz6DeK+mIVaMjH8JoyW5/awPfI
45a4ABO+M1Ni1Vwy36zpbR0gT1sj9piec2SF+djn8BmX+Tx3Z/mCjkJ8v8VnSv6f80Hw3H4rTaJ4
rFU/CmHk1+ae6vDakcH0vRH83Zb+Vb3Ga9b8a5JvKXeUnxaNTP+ks11/2pLC52fONgGrzFW907Aq
cgKFhQ0zHETOIkDUppRGu2UJfZDLUWKYk5SyxVI/FkEaQPCvpwbPrsu71ohYzTVgQND87UdCN2Aq
DaUTfhEuH0n6jqIarS5txd+eTa1sh4JU8CLRpOUBkKaDLj6JQF29GShSggR9q2L4iyf3SUvR7ZVC
sDBGlmUsCUGYDOLTCVRqKXU6BAGR55V/p4rIiYOs0b2T88kbMoTUQJWe5NtDO4vUUmV0Er2+r66M
/VgP7rHMIekih3lvMuHFXNmK5vidWneeR9I3cEmqOEaumno+4KZR/OTL8x1+3jiqnfTHngN3+OQX
ZZ36G+YVcMtVbRXv596I/KDvzRr8wACrfKhOMijeYKOABJdzzjPe+WH2+Vj8mdRlBnpaV4LKfF1I
iJD2kXOZ+vwNqXOmKs0wbHccDuQI0X6+roMJdEztUhf4MYUa1w+vZk0nlS6hd7nxmLFqqU96K2T8
Qcoa4a3mT+VGvTEL7YFAkltDGQ8lsCYTzUXiS6SLcAP5WBD3l9MdDzMs4Ur2sUM1n3xh1qLmI2MZ
3p8iftCzRNzPTfobv673IeEpHqK8NT8ssIz68i+J1QjixT97ZFCmzrXlkP0Gd/qu3Ld9IdTxebL9
ka/B0X8kLkQUqt52fD60sw9V2F8XKxRw4wryw52rrJsqJhYuvGjKnP/k2tnVrSwSl5ZY+gLkJ+sX
ejxZRITOefDCmDm0pkT0zwctvr4+Ys4f1056SKZH9mfAxoc11MrMIBuIb2/nyBAKX2XGJcXUPGLw
4FPBiclFOCFyM2MMWKsBJpTcjfkyDqOqbpt4xY9s47Gmq+wKVsZCbupXi5zsrHjTSLQR8OMNL5l9
szMFrImxnzOGnGS1ykbl8KdtkDDt6cUZSwNe1OqaWNcA2x2jpWqkN+LL0P8Sd14nlKOogGcdxRqW
uawBxLncnWjO4eVE4JI7MN3a+xgh4EvI5MHNMHej0lD/+feWhODVOAo+S0Y5PELSABCePEggGYMS
WcuVlH1m0eAW0bd22W1F1RUHVgbeDEMPpl3cvUibB1V310PCM6itq9+PxKOKhAs0zCS44Hjx6Xpr
X4JiXlnaK6pXEVIvsx67gekBTpuWeedrmFl+iiXe9iYB7lvq9ehdrZ68l7FK5WyEQMBGSbYvjAhu
TfbQX9jK8ZUOiB43xAwnZF4vrDBR3wxRX8Kgv7+AOC+vtsMmY/pXzlQPphYze5elXmuGifQ+7S/P
7HwPsT/RskfdkmlvrUxryoXXhYqAE/BquBFUpa1m49wwgbu0rQFcyFj/UmNsMVZZN8zQoMJPq17L
hMPjFjw0fKX0fFY673hlgfhEcyJEr8PDJvIZYDYAvdKA16mWCeAqB/NifbypDQpamBMGw5B0PCM1
LZJnTaK8r2rNo78NLWoXqm3aNIIdieW3ZLRp7Ufgjh9x/QAIFxJ8pV5xGUkOH/r1xrtibOBv/TeX
zznoJPVcIELZe/NjqQsI9YiLmn/D06YFWcptAzfI+wUHma5r2bJFEnpaCQErtjdFoKNAsTu+jnQp
dWXC7F7ZWkxrh+83qnLOM4BfUVkf22jYX/+FHLCqimkURiznfDOvyAXLVK+dEHG7w8TLs0ROvPdF
iHlngskRtE4hxd5sew7lx9c5XXiq3tplobubcr77i11jaj5Vp39hLN6n6N9w2fLtUE0mzm0qsaz3
3egBboFvEY+d2FRwpBXIbXJKJAupPaidkiUe9krwwMg+ySOujJ3Wpa7cnfwnSMnpFXagDVIW06DV
SacYKVp3tiRg/RVR72avQk79rlziS/12XjyK9eKjjbq4RVRXfNwE2SeJ3Z1dV1FBQxRe1g/ev8Pg
XeUt9I926hButeKUysBDLfnleU+MtizpR6ttb/kCLo+SDhHleOojgqbf9OLbv41rDCFfVs+Cq2Xk
hznao3OwGzp3VZrOvWThWavIuNobXnoFNZBpZ4zpDLWzUJxatVfgHJMfswPGT++zmzAZaaB8TZsP
k6Wu9v6S9p7SEwd0AgkC+Hu9d5g0s29ZmtSuf2kf/gz5WxO0SySECWeWnD/4BpKGH/88xZSWYgbk
M4M8fYsFzqwuCp9GAqneDInC4Y5EEhvvb55Od/AUk/MWt4gTIlg0E+NHdaTeREm8uTHTn5+B674L
XyvP8hzXqeXHnZnVrs41KR5uguGBQkUGDeo+nKHWQMaeR86Xvo3IGAtuakTfV3RIPfphFCq5ddVr
Dlevdx5gAEpXV9pADPmns8I5JwGaiPDX9XA0tRGUiFTja3W4VvqBYoOw6CdbN04rKSW+dYf8Gg8H
OE2AdmK0QOjvkFoLFP6EFVN833DYsF5+mQxWgI0+4dGrYWfUqNT4GIQJ5UNZHOCm/r993fJZgCjR
SfAoz3x0LcATnPOzYYpB2sl2z+6zu1rCmZJRqOasjZ4AvSRd39sS7m3R3GQfVN776CKqZ9cFQ5do
vQ8+sIsqCo1ShyN4KLBss7oVC5Og8q/GcbSRt7iaKaKPJruf7wtFAePplyIBsIb29H7cKGbeRplA
KrSm6lkAofHSFWSIzyFPKSy/0/3ns26Tx80SLxmJDcxG7F4AVVyIgqK5UiYdpQpDYZR8VxBYsyuJ
xhgiXWBV9GBCbrzzKDFcLZw7ToW3x0xxa451w+xzQIb4MwVhnjnLm5Iw0S/+aF+c0UUsQUNO83EG
Hub9qDYCRQGNaOeUO7k80vHtnnmSSHzbizN7gIvOJ3SuS8iTa1gKjFsIk+iKVmevOoDBRhrETvsQ
XhAUp5pdqQloa9j9Chx4N/V76gObPQGXiDXWHK8DVkiWrVIkhX9XJEuxH0RxCKl4KF0YnYE539JF
HBJXnIxDs4SzSUNFDQ7va3cIg3OLN+OPexAMdXsKEm2DxnggMiDq/9M/8WXqzf2x1F/jim1r1Ooc
YFzNaysAF1pzCcxu/h6/2xHPzqFSLzAB1kDAQrYNnhkBUSwgKmroKi8gsbLmX314VY0782HePCwe
azx062EAZpvZmaVK19fqATIJiGG/SAss8IqvOGI4Lk2+DvwO5Tygeetapk+8FU3VrLJ7PLlDwCTx
VzXF2COz5NE2B/8233fRYtToONEG5Su7Inm93hvc2grycnYEUYBLKd/pvcvkhsAgUm4BsTTn0PdM
USweUO3QLEZF2i9X39S1d13SEDwfMJ496E4sUZsq1+FT3Jbg3lJxWjJDIEzrF056TcIOMiPFLA/x
XxZYJreTgDX5umK4OHc7Y9lknYBH3UzcPZkmoQkkHk6yaaZuOnhrE/QbNtY0cLegoiJ6CbctyQXC
Nfa+6J9C2NWVXzkrzSFxEEs8FdLqqcHILWTMaAafA+9yIRlKdKPuLEbtup2dO1Yirn3dWPZ650yp
uGyuy0Ze+68a4zwczoyYLHkyhXz0p21A8LAaiMhlSZV6GMOF1Iy2E+3DlXT6/lvXac/xzgPVrc/U
EsJBm3Y8NJvdhbN+fH16jpK+dGfpEskez1wjxGrimcIxvncGLYoBlUQKXmfvpZEtvGGiRSUyRctQ
uxRfzisqk3IfQwd6z6t9d/BLr5pBbGgMCk4GKOookCQC8Z6JjNxMfQweByQfVj+zYZIAvCHAb510
EThwRd6Atk850ZZEM8z6I/KnUD0SF6C1yJIa7QVuqcHbBzsHI0+8jYUA32EG5Q98oSgw8/SdbHKw
4CuITE7LMP4fY9zYfaEiDv+/ceO8mt6uYBRtu54OlHtylIXpeHyWILVQuilSujGDvnpQwlt93kKA
GUqlpHkLFZ613zUFDFBiHMaYZVYWolFRhwhEZx4MDutGRp7tUlrwYONiIWveVPrsVyoZDxrAhi6o
fy5RqU96SV/5WdzJxkmgA7Cnr1+OXlJ2ezixhTw5B/oUHnC2wcWKOvDAHsUsRnw7rMtLiIfFvvEe
oriDxAMldFbEhz3FtGB3XZbhwbvFHcoHeeJuklPfqJjZIP2aEm1PrKxorqTARb9mo0Xv3vlRBBxm
wtuWASQGtYiIk9DOcR4jLpFg75ldrNzt1lLsqC5eQ0o//QTvaZ4i+YRaDKQQU6oWLTgL+ruyNLel
xZnfHszKZpznp/6Ci+dDiKpqn/a+g9tVpq7ltluaJrHmddGDp9ivnW9LoTp57aFiRsL+wTGCeJns
yEdEzrvTlen7GI6oNF12AlKPP2hH62uk7HsDVGUvnpIrSAaxbgfTApG9Y7YydNeiR4A5CQSsjfwd
3xhKX15wGwywIDzJvtfI7kShJ+a9VutDHF81MPkBe1HG/cx1WNVCdGQyS3oXrcQ4k6GRd1BhHayl
iR2zsXnjhJuEniL0MRHBQUBTM5yUyZtAvRAcWdPdGDniE5vClYuPcuRN6q7BKYEhVvL6wKVelMS+
AJyfUul+bY8FitILv3NHWAUhqXQ/pzXy826+D0Tfj1MFfecfUJk4RoGitK6WJdmFnWZW0k8VbeAv
6bizx3f81Kh7WNOjm+OzHRuO1/znlRYXIht9Y4wZ5oUtUN6wxet/yd3A6TGBpSoyPq1rFQstnAmJ
RZxTDREzR4xBxSONOizlf7FimXLE3bSHeYRmIrq8bHyYLHXbIzvRwtgA4gOuzLQ8NcIpIR1dELxH
2gVN7k8o169d7P6NJrLquvykIkyzlPRiNdQdIoEItJCgF7+bSsYQot+FhUV7PUpNP2hUrLn8LOJ0
Z7TyBSGopnVcpuYGwWtRFsUSXAsyNVM/N/y0ISoSALmS8rH/E8yIfZc8EgHahfOF5kQ7jBqDB+wE
NmbOOCfSLJ4WxSA7vvzX3OJF4FzodjzAkWd0VtVPT+61oqnbH9pKsPRykbBFc3BG8HlBXzPoJL4+
mF01ljgo9ticZYmqTKG63JX1GJw9jAFQWxDkDOllhPPdF79Zm8ftrO/fLA9WszDaUYylUYKGzGWK
nORFRZKWe49xbD0Q7z3SqF92nw2Jrvip0u2pxz0PM5rXNMsQyVekL5AePsAObE3u7ixDEN93SLhP
1uI0iP8TIgaRBkc/3zIQj2SNeMpGjf/1J3ga5+nT+KL7sxo9XV90vNjgCGqLExXSrYPKwRfBhm9d
qr5RTBXlkcTkfgf51Kd/25W4Yj4l01cta0LL/T3HWp0gKmIb77ucjcj2Z2we0WisyaRFSoXBBN9g
BV3cuqjoketar6U5cl6e7cIf7gxy9osxPIj4mc6NePa5Z9H1dhFmH1IoFTn4Bz6T1eyKpvljaTsR
ueHuzhDgQM/fOj1hXtnHTkw4F+dfSY9pU7Sl6Zxgr5bGU3PXuKm9LZRUR5lq27jG3Og98cJ80/yn
9OKPKEjEGK99LLgwZSfZheMpGtKhkeCnbMuS1kh7abwI24d9SZxITEzy+uJL6eM8PW3NqCsHFVDz
3ClVWSW2cikcy/iOsSK79KaSUK5oQpCtyvQfhjx2OSzShphvj6WYvw2BsuPfDtMy368gRy44HqfI
r4C3RhBrGQuMynBVuwJFMf8gMBi76WTfJn6sAGtj5I7tyCw3Cx0h00kxaFT/2/pje3p4d4NxI8Tl
f/T7+U2x5u1lHSLsKEbkQ9kM1udYdACVKh7eAcRz+zNta9e+sS5Imyc/TfKcG/8t2JmCsi+51lJw
/+b4nfObqfUDzzdnQJtvy+ocRuwXXP/PLu9uZSgTnPA4+M3Hmw4R9ByBL7pMcZofbqvkK9aibkdK
e0kzH9TkLKHNPPPdXafFItm1zn6G4/2p/1n4CjcuVEejqZ+iRnB9zWn7A2M3QzHMlvcs2FpLrRSw
9uHvC9gXUJ5RqpbVFCRsAXkfkwefZ7QAFhBzxoJPe0E24bosx7coDaNo+QOsA78GQNSnYb84+Ixh
bt19k+0BHb4kbcUMonhxgbisoJ4TnvKDmjShfkyTodBcI0lPU6Jds4U931VslnwCP35BLax9ZHm1
W+KIKtQF8N+hVZP/fBUZv2yeZuoBIiIM06W+dkJFDi1uGJirABToXaj+3Axz6IY5fUnCuJmltLFA
iDPQ8l/vgADSvcdbZ6gf+pbJecmyXnxM3sNyvwk7yQl+epQYIeLsk773I1vvVIDrEJUXg+R3EyT8
1GJ5dEeC7LhlbHRn6qX3e+CDIViCH3z1ahcOPTb7DNhB/9S55t89JwDSEBnCv8Ljf8al/BZP17as
BTGnBuuGvlcOHKvbEo1lpev9lpXgWcFQjxajHiQWYz/OBcaxNgDgtVD8yQkDGLH/PWZysJxhqTFn
y7E1ZoBgYMxxo+77ES3YmYOQEy5aA5xgc7bIjJfW0J46GhSIeVoDq1I5ECwi9EY8Nhj3ZPjht5zQ
7aI2CgLVfTDkw5q+StbGzto6hH61OhHNLwp1qgzB8WvirYHhLgpuG0hs256KORGu33f/NWzN1MTc
dx0FQUA1zEoiIMHFUP29NHzhyZ/D4Wa9L5w9e4N/WBFBe0ji4YS3JvEL8NRDCbMjgRwOSanhNxbc
ad8JEnaHlRa657ayHGwK0slleTmRhEM47UBA7vFrokDeRpWtcA/Z8ml8H4zuCUsBAJmndDvFxutu
+EGK/uTh4Rkh7FeQMgGV23idOPlC5CBPG0TS3Mcc5wZr3TafGdGqOkcyVrrRVQ7EIaLeNKeB25nr
IbE2dQIdn38f0n3tB13MBeksYv/sWS+ZJgeef5nkCnzvdoFzW77BMQI3+euZ0kru3kU62mEmmTMn
sAG9gK8qc3fSk6raKAwjG7ytZPo4iOfJoQAo4xAsMtW65EFffJfUyFB6dj1h96Hl42Ht67pr1Mw1
B9Nt2RXZsOlTjNEcKatM7zahcclSn4HrvpVmYCghr6mF37hXTE91LGidTf056qwBBmCFVlH03H8F
G2FnzgO2u+zEp/VkEBIjHJcm0xEw9Hx9I5zTm3eKv0W3IRG0oEUQBzyG6MuoCU0WiR2xoFE7aVC7
iMF5YKBHXpzXr5GZ7fKjsXJTLZsQWh9K2k4LYYGoqZiipjXvraPuQmsLvKznZb4o8K4PkLSPDgCi
UygQl0YrgOg3WP6YO3/E3o3x3A46xWFdw5Zl0yTJ93qB33vDhe4x/ibn3klcKfuVmlTjc27eE1lG
4tpGh4R1ZXVt6VagtI3U/KsH3bRM7ZJOgBANCheIYl+SLI5j/UjU+kaXkAEPhfqU5P1RAWXGM8io
5KDVgKn/JofqIruPFc5d7ec0sgLA3LSJkOdFlF7BD/IvFHf7OzNNlj+twSKdevY/b5GP9Reth2Ny
NZ2UwBd9/FRktOotsAlqN6MoEA2f3GIhD+tPS/gAHDJXKTDI5r7f2SbsAz+nerVzUPpofZiwMKEh
a0CcLGyjlBfdSO6gNi3CZtQ5/CQxDdLvgpprpx8M06DqHZ7QQwmEqLN1tjr0VqkhMlGOi0T2Mfze
3/44TAIUQm0+xMV6hVCH+qlWOgcNftl+NE2Z9sMubTHTIrUWiLKBqfaCizEsjTk+4xeIj235+yvk
FypIAkBIuGTdfdzYlVz2gliOplPmieFpEPgMpjLqL446Vi6sQxSAJB9NtraLvsWJ8oq8NX1JBfsv
zHPbr8kcCTzbBsbN8ijpQ/rhfVIYCkgukibx791p6X9xlKFPT8qh/DCfWtCMfpgbb9rY2bAdLXGX
tcHfuWaLTrf/h10TI4oLb5BVWOl5xdyfRcQaarpy0BKWQb9y2octh0LCjQhTZAAnsOsmTfZXEH55
rsFhjA1Rzt/N6YXV+5XDFgDZUm+38imVGbV8aA/mq2QQMZwrsrdvkhHMYL6/xxM91mTium0t22dS
dTf5NJ+dbDfKB8r8V3NQ3VMw42MFT07nbui9cB0XRWdFt1UGSn52CSsYHKNn195EgmRRDQz3maLL
9IfN519B5dt1TJnlGiG6bNwcUTxMJpc6NUPwL2hY9TkdYyfBfC+kQaRPedyyPoU55ed0NCkVnm+i
cs8EpqYqDCLbHfe+piTaJxz0qvgxihH7M2F5kgj9BE8CFnBmvg/R/92+UwrPBOnf8eDmCPDQgUxW
9YIOjd5xPjsu01VWSchvvvkq0n2tp8148bNC8yvB1uM6pMHCJ4bF7XwCd83wI+sn9W+QOAvwUQIe
GWoHs/7i/2YnOZyH32VsywhJwn/RmO+mS7hitqKOTr2hxbcLV4fQej9BmDszxN3bABNJGHx2JuKW
QhSdafOrOq3QdOWFozcVZymZ6NEvcUpNMX7EANE+D9RToMLh9BzYsYslXHNjN+XruzDF1TmwLH+F
6Xih6bobLaV13perf1qjmRM2fYEuQY1ovHcJ2T09Ou6IhMtvFg+D+t7VvmL0BVxHTFLFZd/ESznj
6flahud54oTV2azIWjT1O7/LAQ59e0xSMXAsvk95JTAzuxOh/vjVrSDEP09rhhZf53ddrP7yN6Dd
sf2X+jD8vu/XOSABVsCZdyxusphgYjo6nHLW/R7MC4ms9RzcyqKNO0QlivxrQPthevUsf4+mnHCQ
As7oBt/mcpNlTmX3SiBm8SDA5lHczmIqPvbX9qiQo8G6+OrmizYxOb0/czO4UhJigkoYHkzvFFA8
L2ETtshcBkOV0B8Jkz2OF7O1AXj9Q6SAdN5sGrVI7O/1/5FeW1M/GYOJWrKYvCUcrz41i73FOeRQ
aej/k2Lqn5gaun+yKsooAq5TwPBBblQcqQEOQGR5SR4LhRLXeDZmFZTSiCVJNUr/Rh0HHvRH4pvA
iOV8G8o6LEcdTgnzrIvFNANGspgZPwMbqcgdzz3iPlnyNjhisNmV95ZMIofN+mrmmWkEdwxymDWz
m3YKvJiGhJjRUYQ1ZGnIFGxS+Bkm+Lryd5YJhOT7k5DYtAdFkLX1c3TrfVm2RaGc7uOALU/Wld8L
sD86OAMW3bwQZBizAwL2krXf5sqyYUT5BE9sF7b8dedGarrKEHRb/dnaKy19wkt20goFsXz/C9iV
K7NqMCdb4rRqKzy7/JX6Em+19xSbf0WROdVOOANRvBUHW6z28J9LFtzZblHtT3BM4dAYzpSc4UDk
2V7T9bN4q2gLb6PjVxEJUFzSijZsxdTntfjfzWFcwIr3k+rZbqL1eLOPQFT8+0cyCM/kZpNH2vY5
T+FSVw6mfxMY0vMrK0DySIMkinFgCTf612BixFpkN+Hbt1t6GU+bKlYRLGJ7NOR0oA26IvBkZArE
5/Pna7t0tdWlB0NCetMK5wDU+KWvvQCCbiwLUr/NuHPXZEmAh+oUl10hlN6MWJXz3SAL1zDu1gTl
bOaQQFWvZprs/uTR8qnpj4WQRUGUp0Phc8B4WUdqfUawBjR9SxG6XJxmoF/IzXs9V417jgVq+i84
uH71iuqGAEj3aLVDSQ8qoZUXSyx3EWuUYrQsD+ymL6HyNQtFhIs3awAWAoWFHR/PYBVpEMomB4X+
rFAQxaMQjPMxliuNgX0oJTAeS8ixuuzxDAz+h4TGHqXfMg8W+8CFLm8Bwqn3CbBZQ9Ubf0cdo7kf
BcfsxWkwxf7lGpSQpvRwRtsv+B5Ifm1Z1Y2ZXQIZ2VMcdsHhfHHqYtkvQIMBVZ3S2hxcIFTl8OCo
Qrl/qLrnNRhmuL72NPSVLHP3Q35ZVKq6GDIWQ4KY/8xy2rYAIi1J6pXDqZtnUWK4oSpsoHLZ++4l
7VPWJMLs4pWAVWovsQ4QUC6YEP0lL1Gvh1OAeI/fRfWBF1AoNT1Qp8GO0K+KgvZvgz4aCteYOCeh
J+IpaKzJ84KXvEhTfyTNh4HBs8oSS1o+IFJuHjDReaQbiQI8bWBnjgG8ljpa37jKj0OwUuCLOrVG
kbyy/Kd6uQ3WuPZdx2xHw8jungeymcA533Cqu0ME84kT+//ONNt6vUt1BTfIUcTF7toZ/4jnfcQj
HZyu8Hf0ViJWLx2xoDovV5iHl1DiCfuT6MquI2A+c5efcZph9wK/ZuIFRANqjsr0MltfsRZpPGdg
Q/Tq1I6MZdLzQ2ouAw7J7CiWvech4XVcZC+JG6UIJDB3luIwriL3agOcl9hkHWs3gdpXi9U2wXtJ
Z+hEOjm8Ki34B6FAhiWdJR96q6jKXDW9ihAty438o/3lTeuqZmTbTIyk3z1v807LJZI+uiKiOxto
hSggmytkFj/XuvmvFQqNQm08Fs2WvdUELNg3tYj59hy3EwYW8UFd5NrNWEXp1IDYgzkXI5zHB+nf
+b4iQuEUa9Z+RJ6+xqVzt+7a97qLJjTdMzo3qmYUZklF54vkOdcY63wJG/ldP7v6+OFrrRqAO73A
3hXHoWts/ejFI+p4BFghq2LG7H6bDe77lRRfAWA5hYq1XudTXyt3An+zG0K4xb+jaG9XriipgwUY
SeTTBTKvJGVjaBB9Ztv9HBB1zLxcgrn5mbnXK7vS7GgARkVlbOnay2/aEQTqAA3TObXWHld8X9cb
4pa81tdAEiyCCMRk4WedRtxNxEIHzpgqpUUxTo09gnW/S88Q/l4wejkDzEiz70mRqVrA3dQSXWKt
jdH3gULbelxGc7wbt+pgmFGwf8eZfv6EkoobmxDJfMKTNjtHe8kJKbNB8hSwJNfjg8+eHRdo+yW1
Fi8M2LCcG1Rq2NwFQMuTBB80Kd09FRolixHvWjQRxMnEPBCkauTZnnhKRxOXw9tYlHneO3vSiVMW
PK2YOe4ef6nTkaCxqtTfXa1f8fIcmESz7mTeBfHiuscbwp3SiIxLpEqkEk97io987wcIDKaXklGd
37TxvClEJ8DcZMNK0Pqd5ZTzOxcT4s6MAJd4OR4K0wVLBsUKet2h+aOmjns8LoCTku4GG6WCyj9Z
hl6Oya+4qkHuPFHHSetIQxRljOIJxt65HGVo4/wvrEyfvOj0H4cTYwy5azccbaVwdYyrhn7CmEwP
gv1MgpFKjP5GAhn2DoRb229sPnbKgeqiY4/F2813Tj5Et0bKYnquvFf40XFiYfwslk/MeALURBhF
293/9K27o+PfFhiZdd738ZNhB2DTKddZ71cf6FY1OeDcBLAUi17JzQK9JDI14n0Yyy31pbUpVn2a
oVR7cluURLIgEjGOCPceccEzqTm6/USZW8rad3V4383gBmHJn0YuYnp/v2FEGfv/PKYwZZJyFRRR
AdMZ6QUeSLcBvsT3adJIDqzm19AOwx7/uQ/5Zeu+qxfqyjJQFO43nfAFVD61UvIi9hbJ3n1vTtN5
6Akl93KB76D9gd75WJS2ZCF0INZqjRnS7SrTMVwv0DNhxlRXDQKBFlnAfxvGr3khQqevSV49Jpdb
g7HuX+aQkLkDaK/6YBZlOH6o5WjzHP1McaMps4XDIpac9rXY/biEEtTsUfy4EKRM7c6w6MqumcUs
h1etZY5Qw7lPmtDj1LCnAbg0BFaPHgPIkybUaYArdJFHn1JCSkbVmEQvHunJBjJqLF36VrFhlqm7
fmAA7T5418zNJ2k3F3GQHHuCyAMneKvkTTD3rToFt1y7sNVVg0Qz5568UGcYBwclh2ugjWJzndjo
2FTD+RMSNPNhKLSzDaYkI2LfeBpkHcWSJGQy9vpw3OwJxWc4zm0d+/VPIGtHYQf2y0Qm1zBMT0bv
lcS8S3x+1B8z9HX3DNLDd7KYy7poeFsxdlF2nmTMllXrO9RL/JlN2+lu2OiBpgbZedA2svT7Kq8H
IXEvzEJZx1vfhskt/3zfG0T+5Fv9kkJaWWJ6LIMvJZMG1aCnIclUe/JV74SJb6hy1wQwTcnGdp/b
hR/87f0BYFKAlb3PplnUWFO01qh0KQrO7m9flBZbzbjYRR9rsTHCZtzrVj4wmCViv6nOQ6ouk3eD
E6RS0PQ66o5IztQhSakmGskW2SWyG6rUmF+xRFeXvzlhpedZ4MBbV2UZcbaD7mu9OYlFg3h3A6uH
J2dy/1k44FHpiInLvCyPrSbdnE0pICqyF1lfqU7oZeI4zC+LDb1WHUMc9bmQkNJ0VjxSwKL0p542
aSqAxQ09QKDJJTEYp0vKKNQrWLqwecP//MacPtwqXwJdfSEQqgDImkMSrUpfRB40+T6gytLpTebK
b9Ey+g0PbgkfJrqeqrxV6ZE0YY61zGbb08VgEImxStXMiyxVUfoAVHytSvAdcZxwwF/f8laO54Sv
Q1K73wgp5UsankTfeGovI7cHEI0oIxic4cx6F8Bninyxggm/j8eoHAPDbSSlU9kDD6Ofr0CLI85H
VwXCPA3n/k7xTskZYbzTMPRkgPoE83B2U8afITPviBQxEkWdJ9uDGrOoo9TTNZtVkuAHPNCORSr8
3L6Pfo5B01TlkOpVc4Kw54fhCVTRodq8eubaUBKHRbzpmR+zyLaXFsxKYzowidPvLmfbOZaadqMp
oXpiP4DDBw0JpQtck66BgW/4iTonYAYDxvKx5hbEwKB1kJcuCQqrb7vWpwm13jQEYh3Y3UTlkoGh
EAqaNyEQvrUpVRivucxrygNoCEr1+X3+GXtVPlZJpa0NotfWZc6jBRBGDNUy4I3rwhR8LJAbVOMl
TCznQBQED4tkzzpyRhMXpAYGNTYTc9G4PgoPGWk7O8oNnnBEl9/kahgiaqFjkxvNpflW4KR6UMXL
F6hdDu+NSF/qEwBEDhi7uv6c1xzndXvsTEwkbmdX0wUgTY/cUHstoF4FuNTDd3UrI4x1PjIkcFW2
AQG4nwub7/fbxqCZy8qfyRk9pQcbyKQW17/jkIQ8nV1qYCT/tpoDfMNq9+hSYL4xMr9jC5xQ3Pm2
jdy2wrCSnDS08grDxUUEc6cccrxovaKZtbEe09Ph8Erb83GtzfU41Q480n5Mo8wrFRhmYFfrfykX
5oHaCnsGyClWLedAV/e8v8kn1bviVt8NsWsSR6oc9P6ikpYyIv1x6jfuCa5+0yu2rehL37FO/LkJ
yuPIl0vbu4cf7xnjnq/Z9cUn7PlNh5xpq30gJoksgn2vjwr7UPBY/wfamNOCZA1zjZaR4tLu1NeU
HEFtGnWhe7AyuFCxgLNegXnbhZpAZezpMZu6zeAL31CfxrJnpd41Eb9qYot0FRMaZVlVqFpJ2S9M
0lTzCaIyuUtLwqB8zJ6LYkXHPGofn3WmYxRjdEsxh4IhNS6cGlcm73EYR7CT20UqiIyjDpF6TvlX
yQkOnUsD77wBr2A8VCqtyNRqkokHPidC0LybCWOu35+CoZIdOWGpUWICZwW3C0xIb7kvkwLYlUcZ
EoV/XEdBfV+Vb+W9pUsUj2EDWdgj7o1YLRYlrUwTBUZIj2amJjqKFuRLZF9irkhxbjwPqOsubHcQ
X4NcMIuSxVmr7b35IvHceRGlhoDS5fr/Lax4IuZfrCuqAViar+vT6WD8NgAIZylbIbZ5XZz9bI/G
KEjjQHmC0ODQ3F40pZgo/A/kQCG30dBdAmY1ZWKVLIQjevPMwA/hVu1iIOB/eolF2K+22zYN+qic
CPWy3GqG/B8xVH8Hns+XQZmrjBdh0d7iuFBJwJY9GSe1woGr8N/azDzumnel9arbx2ez49+8zkbt
q3yMn+btAAXG+WRM5d5lO5b+Rw02QuJTlZUr/8aQbwzFYJbLoZG+F5/P1yrxOvRGyIKIFb8RRe8o
lG19o4ZKNRJdKC1///W7zkQKespLQ06prMVcLXWoI9LxuHjlDdL1hmDqu8Fih9DfkejwxVuBeZSc
+u+cuBMW6qIvUcTb+HPdum77Fc0HxlzIK1/nOVXu9WlvjUbqr65Uws86+SWd+w3urIAbjUVhG3iU
Ngp/tsw+A3vXQoxB+dyvqa3ZwbxtME1574ao/Y/Nzs8APOz011r060u7zB5W0ylH08hhbEIYHN1b
7+lNz/ZcldmPK6WObJE2MW/hL0wpl1gsi9Lbrfv8wv5qUP+UoTrxkSYXdwlIxkB92sTyTOuZfgva
esKXueG4eGJ7UTV7JpCoHQLRxwI0WAUAlewA+/Gpp7w2+pjIrEbIxatu00OCUs1qfRNTEHUV3e3X
atHAUgRe1X1WARAjhgxp6PmL7+X1gqPbPreOLyss15gk1mygX5Wt/5e4r6rAlr/ePKsiRSzarOdF
9b2tuDex1JqP4J2SwM3PxB1e2Vp19Ci2cvSbQab90t4bQj0ZgWgXGJVA19t7kBYsxoKcOekWPZhg
jiPH7O8xIJrzcktQ2qIwbptjeqPABXakmsxJo4q/bMRBEoljgprjAhmmZMfey/Pg7rAf5DbgTxdP
SyQLmDQnk5y/gUr2RIPVIKN3vmhntkei8glC8dxZ0zj5Yic7McCfaA3JqX8pe1UUlgbHa2LEoo34
o5lrHObU+z91QRFa/dTQOZLokwxxIqJ++g9mnSu+pCJDODL1gjAxU73M1yJjRbm8B5+G3kxzpkhQ
mp74wyIu/tXn1P2FnvwK81OlD2sSCsR8CBKdBaxr4XZP+AiKK9Nrzk9fOv5/mgNvc9ed9acsNexZ
uaeewDzKy23A1zgp7MLvziWWHxDkrArUShQvR8qETZwXZyW3olmT/+55nJYiTxFxiCT7SjZ2A+9i
yrs1tr+ajrJo4zRvN6UrBBa9qRFEiz5O5P6e57VnDTJ9r+YOl9TWQFdUB9oVKHlu05E+y4JfVxci
qO+XXxK97TanrXIud9z+IDzwANQNNB0E8CWADBer5LRVJkgtM9XTRpzV9o+3SU2PFRDeMYXYND+J
SP4cuvZWfyVh0tTmu2w94QPr6z2+MSRF2hSj5otbJGsnL3yQwsMi9iIJWdugCFK9vnsTDu2NmLdu
/TPoBhGLyYFj0ZPrCfYPRHA+DW8rja8YtXhqoyfFxigwZqkl7vfNPftuYYMT+qWz9HQvdfePTYzh
Qq5s7pFwiuaUn+GqY2ea78lONbYWJd7PEXNgLcYe5oSalJ7S12FxI4u1z/mkmJcShiw0kEAizeea
eSLxtrodF6Gb6S3XlkohIRtHYB3nfCUxNKyzH+oO3BFLDWR0SxUUfBQldSyUb2yKhYk1wQbqHQ7M
t5Z7TPhxxFrAQbTxpv0RX/wLui7u9J55uPBrBR2Mu1ns+/rs8x4n45khwHvpi8XV4iyGgm1mi23i
VkJMHAyHbkC+3w1XRATDZ+vwiWZd63UCVIkIAdMftaW5yp0mX97A+V05GDejfGTRoSnXLUxz6rmp
DFpq0GB/lYxwpTj3FsMuyBoQd0Q+ad3uOm/1juMEIA5yPbvGwx+iwUsS8IQIxba0NoddWifFT1tG
MWiOceuuWqIuTXTUq3SnLBMhINrRL+eWIZ1SkEQdNaY3j0q9MpPc9j0grdKj7EV7/wsRJvB+5t7f
Xs7rV0v2381PVUPXvr3W1q6MU9LZALBlb8n/4We+3VxSY58tKj5ZD+EgyfcACw/YDB8qKI5lV1ru
tz9JuRSShQqZBfyERoYlN6MG8soLe7imfY27SO9Dx8brPonsRxJjuiGjpxB4e4fAB728vR574fDk
AH0aHHrJp859NLQmetyc4M2rV/eCdqvh9yAdnMl9aj5x8Hi4RWetHipQabrYT4NtEhCexwg5XRIv
/nTV5DMMXTIsPtH3dX+ZPQEClbqYsJkiK7ukdGTUuwjkRR5gx+j0Urd+CAqU6JgKcky46t/p2fmM
Xe2NGNQF8SwLxhw12zM8Gqn57OIVnr6Om9h6VvrtLD3kaGBVmlsv46OEbRqzDJYZFjMfN0KAoqwL
l5Qadfc77UgvoHmtFyboA1FLcApWao200mqQn7WUvCkj5DDGAs+34ad3oQQyz4EfM8c2khxs8r3z
89ouU/cCNRu+BY+hjiqgxjlCpdUP7O753ejI6X3ZiUp3x3RlKAPDStcyRE6S2x9KAft9sWWfHutv
VB8H4vuGpl72mAjjPVW1umlBi4xaXzBva2HH+LaOg6mq/B2NFtlrYSkbx2AjIZP1aHvEBrMX4Ibo
s4hTcBNudyVT658WMEId8U/q98aVM/84jW73DAqycXrlq3DnbrT+GLO+JlgVhNO2SPIjLZDusUdG
/ORn3aITo06169fFmMAE9E3e57fhtULu9rhe6ndIghHnI8lRvmHHMzzmA7fTlBC3IAPlCQBnSUQH
FPukXKhHWO6yRudQOQYmbFJ9r9+oXzTnzk2mhd33Z1+KG6wpfK5nYL4lUH5sFPJJ1lIr4CukceVO
S2MTfdo/eDIrGekbHADu15FdaFi1WexwPo1hTMIjGbGc5lgXv6nphM2eYPXFYaFj4bsOn6dHSkgT
tCvFmxnTzNvcbYVa7MQsPLE9OWcdMDSjDEm3xUkWPjEpMwTDRtv9AUsb+lbZ2jltMQxQGS2jX5Ie
jQ/AyOTkun2ocTGAFm4BJkPlSDYfIpGURCF/pcIiovhjnV0h2U4PO0DP97I8y84mAxZq6fem+fXq
BJKF2g/TFKB9TbAS1jib8/jJpDsVECqXOPjuaBKRUq2ZGQm9l/Ph1DhM6jDCzKVyfHB/GObYwt9E
Jt48OzQ+XsPapEeoaFvhZvmeKSZBQUouCYJkomzrG5kaElu7k7mR7GBl+y1DLNvf5SMlhvR1HIGJ
8uzVVIPhGLD+MDCt92JoAg5JdS8nMHjIlbwuAMIadKf1s58DFNUqa5b7ctWJDOEJ1XWlnItwtTZO
lB10D4GYBs/UGUhXE0n54paN6iExKFD/6jlydcMDJ7+gyYoNsoMpewxti7tUPb6qrj2nrevK1nCs
tuhlzbwrZAsPXtN62rLsbXWPLyCuzweFG6P6L3i6t05OhHlHWTmeWpFe1C12HflrCSG9AUy6g/o5
VLiohz3wBVt8rc8GYVc/JmR8POdoJoECaqYz21GWPhCCg7c2qwK8yw09dW/e2b/WgqG5VM394Zgl
eQEdO7d7eWQNZvrs5dvjy2b+azgeoWKwPZaF87cbpN8/BGczK5fwTLYBJgvKUR6Xv7LmhTfdr3kd
WW1b8lnSRacQvajUIzesQ5Ffs3oU3hUeUP94w06ZS9tlbFqAUW6xLmwHRhvXVxYvXi4ds2k2CPBH
VfGlfx/8EGo6qthBu52C6eQGHEmiE9DJQo0O48urV+8+bhArrjwQlcnZfgnPuh5mLC2runILtUfi
UJWr8zLKZck4n3l/0iDx4NiBTPnI7iBvkZXfnOwonRPvHjebffLr3nXucxUocua8JFjSzoRXxDUb
ePycGak45oTTa03p6KfubpLoCPOB90aTnZmETxyatxJZvCHpf6IOM60qNr8MyWlvFf6xH8Jxi7fq
EBLm+1k1UeOn1iVq8pkIh+XwIuCW/f8ibQMcdckyUMRxw3HleVW2/5QLlzqWIebjpJ60r1LJYVia
GwQrCCwM45WUELFoEXIBpJcaG/UtUeHOoiOf/jKWt/zw32b7a3bNShnFUx84XQsYKLLdWwHx+IRM
EE+5AUL7WL8ZIzaLN1Fx13hs/Dlz4kJl/9rjhdA+FbC9ilHeRk1SoOerJ6UBav4NgjqihTEhcKT6
3R6uVldDrVr8z+8+U08JAaS/lHYk9H56gy2tfXiFYTNF7GLiLqzWwMrFC45/WX/JIA/n9P5M4PHE
RMcdVbqjUbFXdpveJrQFQZl37x3I4Psdw+5vJKxR+4mlNsZLDzEY+Vz7d/NSTLmU892fZUcLNjo2
+FCm3ZBDcaO1qAtr+iMarMdx36SOqZCjLPVY0Zive7ld3+NapHKB/geIkjTHfLn4bgulP0dGeh7u
fml/CCaz+bNS8E8YPPnhK8Er6vw5IF/1nMU+CqfapwtzSU4Bvb+KplgVmaaNk6mami16ucyc1s3f
hhb2ml8Zqtd7b6c4wP03Yl6amdF9OzWpBbzUefESz5WZXm0O7UN/Ku95VT0ngGhe+zbCylmvw2wf
xB4WbU9fHK/AthapcWOCoCgaefYZ3J7QjGXPAoqEP1Lp+IkiH4bfynBHIgrx+TikD544Q2U/JvvO
kmobD9NCcThadAjWHXCH+vWpfUKBd1zpaROMQ5h/QjN9xF4maOZqSdFgw8zvpuOCQtG/si3zLEsk
ShPex617MeyPUPPRCIAxyHD23onkdr3ADBfZqNO/iZnB2JrXyGdKxTuuis+QAzolWyFVZIO0keVN
TmnLmx/AaOa/boBhfyp3J45JNQ9nqRAYy5fkHDpv4f2kpNbuXL2Xc4cApgHy21zWweMmkw2d7cSq
vDHFbaBt2zMp/L5WunEg1s4n1urdSO4wIPDDmJUhsSLOrfYJNvJ7DWszbUm15qUb4L8LuB5OyQbV
Dh305F3sStubV8d51uyLqUEXGKhSVxp6kqnuQmb1r1MnjWZYvmOGksH4Y1FK12klHK9luJH3DV7o
qK0mAkCBN26LqVD6qJuyJI7+ZNcjfT5i/ej4ozWUbJysYiQ8ZnYg6rGDO+Ln16FQli3KP6MFXcUi
PpDKJXt7Zf1Vr+0eWAnzmhnvuahJ2FduyyVWusMwf0qnmhPwF+nUw5sPs0azgzGY8l7hNTruglP1
drg5ITzCs31cL2gUKb25hOakfoSbTn1RM+81dCImTJJlcxdBirwhRGQdkA2XpNPOtjAxLOiiGIH8
czhMzykv9v+xAsMQgKH8L1CSlP4+C58c376+kh5YOSmv1AKAw3ZtTkkFeMCBHsdEI0A76pnSv8Fe
J5S5Jt36/HW7iDePedqFjqTbwroCTNVZZxWw4kPTjB4lAU8phefBpquEWsYaaew38CrvtczFUPFV
2mmNwrMYBG3QtUD5XZKHzHEFeJP6/LfqUrEPupMVlthur6S5K1Mp5fmEju3x7vryv2EO2QpPxv7r
21RAw/cAPTzyx3/3aIe65ukFxmAWusVzOHNDqmw1OrF5Knny3pn59dopgR1vWdRujEbUR5eI2gDn
66ZtpBoOLEjqNTVmKjoyhCxQfEMK16QmaZKY+YNLpCzs7itRpnO4r0AkRg7LWyfMJDKXXwWOWe2Z
ixg7IEdEECx0PiFB+gu70tnjgq9s9biVUW34qD/RepSYRX5rtaJfG49SEvm47lw7fcWZ5Xd5ZbD8
rXZ5IAPNbPCfP0OvcuzI+DFspctZWXcP31VYe3JE7Vn22o2UiPldRRpkx+QHYxvSgrxNn5A7IqE0
KKXcqXzRz34TCmlIw1quIWjHu4L7U0wSvsg0xXy6wdcqOEPZnZXFN6pVSjto0YNhdhxiZ85i5ahk
ETf2iOPdOzk9WuqIVU0E7w+tYOkwyX+dN1hgQJ9qKDP1SJykFClufX2O7jLbSH0lbwA76txZLiKm
m/k6RdLf831EqfW3fkbEzDomIij6dEkHV1xrRdpySDniref9S0hMx2iwP4ySWIo+hsqrGAIsmQnd
JBGcvA1HZ5lRtkG9G6ZJd0N3+vEW3vHCArUFzrMYTAAies1F0xemHKkRu/80GIx4YNF6fL1ZNIXy
jxck2nLkNBvJ3U5GU8F3RYphHeLq6IbniG1w5FmKorhWALvRUYqyOdm5Zu3kNE/LrAUV4hgqt1OW
Ws8nXFt9un7biQkC64DQjg7J3P7JV5N8382G2r91YxylWhb8W1hvc8jK/bgi0617xXoUKb+t73cn
FsHEQrYvfWzf8OpTftjdr7J59xt5pwV8QsbOYl4VfmeL0038zSK3/HBSrLusF7BBI9hiaTYqBFwy
b9pltVpX2K7dyUMfSIbmf/P3fp9tlnfljfucNPfFpOhcmyVk9+0j8izy5zVTtUjvPDc5ZMsLNnES
CVdAVQ8aR4V0cFe2AJ8RzOnhGfvwZg4l76SSKSJh57eQRUkluj4w6ZHR9R6laLC2SWRH2m5jbuGF
djUo7Tf+C1sC9YSS4UNLJMjD1Gm5ldvNZQBjL5axytVujdV5WomAvdx/llW/LjxF1zoFErjDOTzC
HCtWs4drM+DQ8N921OAlPkSx56nxFUXZS8nFX2gqbkVJFmiyoqxL0fO3NA5UrcH5U+eauwM/blXQ
ViUw0j8D+q34IJfGlJeBph38XC09846iOwtpW0SIpQGJ+HYri0mLvvnqSvjfBUoqDkRI4tFY6HeB
pqCEjBEBFKjwhDjfuu/CKgFsMGzwfQ4qndalvJPu7WoxhhMjLNYMF0igRf45OM7oE+KgBrc0tknZ
5wlnUZThYcuCMUaU0jpZXez1PteOvAdEXk8yDdnDuHe1rPHBbrGSVxqsRAOM7oY1d6b8PHGEyloP
DD+GNiCdz7zHL7mFeeqVqCZYsaHHX223azKLqWREeAQbPg/uAQ2+W183lP3xw3WORFwXIl1dxyKE
L6JCm7/eUxJKweiRIFz60fNdUsaQoLMLwcvDrZdSq+34inGpOCpIc/YqKB/HN3Tm1GZEVwrXXYfx
XvBfqV1LE0Wd4tNTT/zTCOLPG/2Rp/96tE9zmAkRqpEm7ukEGqKZ+AYVdHxuOdlwVITaS2gIF7vK
dGTouuNToDSQ24IoI7fALSv4y70B6AfBdcZJNZVkXgb0Qwbx6RuFLXXJv5tGofOrikl/ll+b6GIv
yVv8V+5hxL78USbJ3BSIiJnxnFEVH4YKbFkiCEA8I/JcY3/lBH3yFdXZN07HwMAN5qNrQLdJGDIf
VwqM2p+9dVbJeAl1QJA0gcJXuyNDqwdQ7IA5DXaef33GGbuZpoGL26TFrKOGp2AgK5RMA6BFqe9H
UNBnbxq/zCVf+OARHSpmazeZ60K6fOK//G6Dz0k+ymd5f0J3cChEKKjybG2INNF8N5Wbc4ymBN8Q
rFEurmtbDqv82jrXUtAE094yiSiGlEEdFaS2ie9HE45fe2r89qubuMUgJoFAWm2V6z0Ez8WGi7eg
1M9THky+34NqScZYSP/gNKB/Eo3xTwy27/meVaxBqP0ULNExqxy4DD1WNNhhESkzOSA1taRcgC97
t0aZU7HB6XvXfYDs2HSbaLYQ7eIZzRxBlRW0W4iUbdBjsOIMYE9bBCj26wcDMTVkq3HNSWRC4khw
5uFYQdNmr4vwWFN3NzY4IppIOTkTMt53xndvtblHB6mU7CWzHStWvOqIKQ5xlqyiGR9gWqvRaozm
OziSLbN7THf9RHEHWhd/PLokqTHO1S5jFkteLkBJqH2+mt5gX9NdSVsh2n1BuyuRZIfwO0dB6lGe
aPB2NAIKc10ows+Ho5evq4EykXaEWN87Zptn50gWe6QTua0NK4OEzOdcBcXsA+YiY98K0gkGQK9c
L7m5yBcrG+Upt3KEEvNs2p/i9b5vbvyfO6lR02s4Au9WjYEzhH8diWkDq3tuG8CXoUFTFoov7TZJ
xUxvt6KsSlOdYFVEwjyQbI+iawt/V8kJt7z5RFQUZJrrOBPCc6lr7StPvfmkT5SWulh1xxTN1g91
S3UIVwHdJMB+l/O8DJ3mNpnM17AUDdgCS8aAsQEr1RNS7EV73ydCUJ899RBztH9EKGWJrVcarqR5
iKUCW21Mt3D266erUTeQeYpELG8+D/0s659yivK2ztvLTuafY+G2cvXtKxMy1PfMZn/vCRkrrp39
NpYKr9h5oWszTplqVKtdYE8kVeIMHm5FnBWQ+hnwgVnhTbeimej71ZRBDVmBjtds1iCPFlE6Xi//
1yYS8zoCNu7Ev+CTmqw+jqoJ8Ce7Lc8AwpMsV3JTtaQXpc1hP36gGQjqhNWQlQkcJCsn94qnthB3
0KG/q0kEGadBnozExCjugO1i/gIEVN9FN+Cijlrh/9UjQQoW2mO9WdsLkCVkvvT3asGcAFAiShB6
k2MTGgvDOtZrzQON7rEG/Lml0HbyQFNcRlB+8+EnSHSFxytO62dYAKfvABwJoClSTGXVsQ+wP/j1
w1pbGJ3AW6QDYYarrf7WOESfzJvr93/EuYoYi8HZySxD1eIycFEAWhU5slD20tZ+4AntRxhonypQ
BKUirBCUuUACCz8w310EwB0nZ8r9Hz/YQ+q/i/sZmOWozTyAZbriBMBpYmaGvz8Gd8Du5qOTtv8X
NIsRhlo9tU+hsPJc6wds6KtslSg1F99xh2yzIskt3Ebn5PTFQyC5G3a3e+I1PBKdYR58cRW9RnpJ
EnPGckA8Hjc16dj5nJXutKSVVtS40KbhLpZr0fZ0Ex5McNbpwqOKP7csO0Mk3gAtt8iCF3c/ciZv
ca7gKWkxcx8rxkhiCnOdfNS2uhVt+Hr/0ZSWaGutCzbAXFtAOSx7Wl57WIFbnquVWTbC3nME8cHk
xkX59DnSzdHFVf6u3payay0TqF3+k238YIQGk4xbCMSzyM2ogPJgWhyJWNzZwlBhbcDORlXGutzy
utZv5YgJ0l/v5ACPLiBMd+LcCpallgYd9+sx2ed6xUstk+hl1Qj0qoejeFjmCg0FRxverEf2cdDn
7Tlds4/yZhlS+msRv07Z6XTsQklLrUiXVDMYoEI/SRYyjvJHnH/YRLJQvXTa23JyK4WeZ97SMwn6
xbOXjr8eNaL39CZ6QsAyx5IyP6OSenM+XwiKm9u//R5/aoa/EbM09H250qBBgTvZgR580/SBhgHo
1O1pqpp5FgH2FduybMU6HezSCtjFvuGsP7SuvwRwEf1J97dCO4BxFq2NpADyKxyg564ZoyXRN33Z
6fqvkEI3XGjLQSfAj3FL6b0leavMILcYfVprG9fR5i0Z6Fb0rTB7cGh1vNAfZae5CIF7AFg3VTFF
2b8u++92VNNwxhs80lNOus0jzq6aANwPEIsl0UQDv0ifHBd/3i74ML0xCREGhXoNGM8GvLl1cNR/
5XvRqVKAeTOrQ6xJtbmM5ka4n5lIycEGgtr4LOJwDYDGaVRXozAmQhkgFkCThx6LH8kJQIq93xIf
RBEAz0aphv+CBWinuspWF0XVdi/jMLGvUG2SlwDhJ+YUK7kpR37I0YvXQzeg4hjgW+zJcVS9xtS9
MGHd9FC5VFcO9QHEMliFw8h45yyyaysxwUdrklkKFW2WsaInWpPdc3BkvEu3jiWwtiVk+VhbxzTk
Vm4SLiJp22+fxp3ULBS7KuGF7AYFmQu8/5jPqV9qbhV2DOKOlnRSNVEVa31Yr1WT823Bwyk5wlIo
WRAxvAKsvwYQHGsi26rGnTxK7XREwOqHHd9aL2ebn07Qr5r6/PDTZm/F2CTrihnvKgdk/zgfijI/
c7XiBO9Ljgaw3eYwHRPq3ZF6EsRavSglacawNRLUkK99LEjO/wgSpsAj56dHjFmqCq3BYNOGJtjG
poMVTci95Ce1309zCG12NHP6lQPo3x+R9xcQXFauABdnosFlxMQhs+oqe0CGZAQB6AleCXYAdqh3
74ZyGt9RX4rYnIAysdxlTZRimJGZZtHUaBKo8tdCKT02dADgkhOJOy0ng5OLZy1hRMxnHol7/28m
DTZ41k2rhQJoaywOlj6dow2b0LzWtpLuHFf8dYcy5cT3X7MrmlWm6zhJrSYuAHzWwOIO9YC/vBgv
z3JFBeAJRrCyh9rmoqF55TY8j0kPSMsDyh7nnVOlZgOP9G0V2/ybY6Yghw4xfmhbjNfgBztHvyL0
Y0aa1eeVmDrEb0nhI/TXrj6adaUeWGh2S3b3tnvidPPlj+nFf/DPdPbo8sgg81Rvw2xtBCxRxmVh
SBHfv1Ap4ZN34uCxkLFkq8EuuttfKh4QM6qBTNjXfqYvq8rjM51YYHPWOS4lotabnYBayG8M4kvU
bqvbSKr9ENhVqZawm1MbFfjGcRyuw46EIYNyZHksD3yMEJQY9ltT6Sid/PGricT8YDgiMPrvHoLb
0KfKZagXMwaUzUUWF9ZSjUMUXBInrw8QRgl75apVQPN1R8cerFmOr6ITcxzuPFOioBVIMhTq798x
qMs3K5gFEG/rVuWh2pgLs5n5Kc+mkzjqtiVp/2C39NmTH52n+YxSb77dd14T0BYThKc2AadrHSTT
oUNzvuC0W7aaswQRjmLgPQb1QxaCUJUYtM1bsZimfoZNkdGTgDuNnZ7sTVDDJcGNevWVOZaewLyk
w7Vkmhg1fHGEkHcbnZAqmGFVVh16V5NvgbRE5dOmCcrBvevr7CzmebxRMMe1s1yZXYZEU5J4xKpa
bSmdIssFppFZncYe2dEQ7+iMfsvPON4zVoalv7E62tj3hNSHaeug+65Qd970iPxFFc5vizT/FUbD
9wVyDPg0fxL+N/xfEMEQeRBP+ogeSkaau1HYBNvmdLptW3mtx409T1nTNNzy42orvgCi3B7QeXdz
j7ddc+f2eTWNuYtbVTMY87XkX2+GJKxeBeGD39DH6rCB0pEr3SEupOJIjMCTVFRz/N1CcfISCRs1
kzAkz4ltxklSnYek//M0YcKbia8sE+gHPnu98O27BKiLJlaEnLspW5WTTb3aFQ2tQL7wtGomBrvL
rlQojN8TcuM4OQyA7fEV1gYnnAiEWzBfWxftI1Oh3+3oqrgxlq8qy+wR8L5PcXcgBifDnzEF7Qal
pt4vC9OPLNRupJfIyPvlFbXq7Q65AZi1Blvq5EL2pNghfuK2sd/qnfSuVsCmAtHUUxz8GRA8zXKh
3x9khEPyV1tdq/WrSbouOmfRC2MVMbyPiT3AeVuc5+UqfVa1dCDub+Fz/GeUNw5fmMtKhOMtNZxl
KR6KWj4b4i1vXXsu0RKrSzFLqhbIQ5/gbYpkLtQ3A4mpLllGH+NONx/DnIOkq/0RTBRBndT3X9aj
IqK8il958uxZ2LpzELeTxwk3+E3IyErJf6WyTkPaPEQG30/YRzZ5WrowrAwCp07Zz0s0fYsKpaww
bnA9z6SMVLw9NoQVrrMecCOjywULMc4jCrFouTw0Te9hQ8Pl8xvN9x9tzhqJjrSmYfO8sOXRmX+R
0oAGNcE3gFZh2WxszfWEOXiZVhfAOFPJEIcIgQc2c0beeceibYjnjDOT6hBPwhbEjRloJuZ2JY34
YDVYzePZVdvDQ1RoGjYTXIvCmheZ8OpCZiDDeYA6lWKNOoAXlhoAz/KK+Smar8RruIH/JqECVi8h
I+l+EK+BVC7W4Ed5H9O1LT8lZQK0ggGrfim4cotlvakXpndBw8TpAH/b8jYc73W4Jy4IEhbpyWV/
4nVTmDwrisTaRoIZCODgyaMxu56sYJ/AmwrGVNU2AHJqCTabGInfXEvWQ9866J/xdES+jqdfEnEC
cDZeTIHV1V9dmHEdJyi5ZoBQkR6QBhhfhtUJUqguVfY7RKMUyZt4G5CU4sQ0jAlxYPsThRnnFV/y
x/IICpBsL+F+OAG1DuanUiK3OOrpzqBnk0kL2fllicAutkTbaKWN0PfVAex1Pubry8PUzX9rxlfa
C8ZOE01Rj40HZEegsdKG7mtNm44Vlt6I8ElfzNCl/T+aOiEPvKLZWQDcM/XoDi4Sd/GhaJj2+bg8
Y2QgVlOLt92meuMep8vA90zT4myb6DIenA9PvrddFJZ6/kITmMvBjCkmp2kdfCm+jXoARdtThayS
63ERZns4/kECiKys52fczhegDKPU5z2LRd21RNmFfdGuNj28EctU4jV5hfCpOO8zmaf4jt/3M0HD
5vXCfg8p7EZU4lzom5bUFaVXD5G28dqE7fgirSakqcANW1o2wgnMC3gZFIbt20+YYQeS22NdNwWg
hjl+oHke/HmPu1RZ35YIH/O9lz5o6hPJ6nvo7LhjfhVHkbH7n3ggnYS5TdBmxF/JmNjkWYxK2Ctc
GNRWKkW1goswxnW6KfB7UrkM08jKJNzZ6oRwESqp5APErbuEqGgTBYs+3yiWxj6t9ISQvpyDNkUI
Mi77QSzZWeLNqbsCjgiUcIOqkJQT18K/z+9bfFcsJOJ7uMDz8oP9aMOYedj4LDVqWrDCKh2Nz3aM
jTSr+xJTgwIwvhwYUKaNqcYBTBHKF4/qFblnjmLIq+dO197mdygVbG7ZAOjVEcMyq3edaGnVlydY
CWR/wRlYvmFvj+aLTNtwIfxhGQFfz9SvE9QoPcjuMlGTj+uYRBZ+uIji8dK06mt7GdFqWF0JIR7U
srPl2bOENDmcqbCOHDQkXhXNSIt8gShVw5///S/K6rfZcbTJxrEwtLGhTVC1QqWWBGOqp+Zq73Es
NYBfSW714T2KfKakqVyMdlWUAEMk8pHiKmfEW+aBv+Tkn5v2Ee1IBCgc3P77I6wOe3sDVVcplTeV
0jawdAjwmB+dc8CM8kkHAS4yGoK997SNngalKDWvunxnxjomt9Hhl6R2DSbIibrUR8BqmXESnx/3
HQ8TM5H5KcBGSQE2dxEPug4prI/+fLUEI8ctlJ4Isbib/n1RF1+DVFeW9Tixj55D9HHC8DzhNmT3
KFCCZVcwOlOFjv2JfEF33vCEMrTwRvN+3a1BkDCiSTFMlb9DF8jn0qzCK8R92PqpWE096jYkfGTi
1+aHmHN/WVexWIR22hXmc5JYedLXfbIKliXYjA7Exd82H4P8n4/OqT5Clw54Si5IjhdQSWJGxdv3
E7qk8yxAkVSo4RD2BMHvbTZwn8vNPDtDDVM9wZHMmFYAu0KYVqca2y5lFUS7+6eaL3ROluoP4j9V
YQlaVr6D4wmY3u9st0gSJNJ+OmZTxYjzEBptoRdryeMrYobYL2bzilwILhf02XQVbdxrViD99KHl
jq96DP596onddV/vgjPBvUT5lB+hfNDgaytB1X4u8wAu9Zl9xJcrOAzdEWssK8HK6a/T8WOdwXVL
IH9B5GfAnPYXwpKPh3l8YdKTR1F4XrTf70VfTJtj22eLj1h/7lU3o5fNUYKe5jhPfGtcEm7hAA37
pgeveuHP2cptdkFElncGyYA5hsnnTUCWsySP/ssyKI1toy0bJDXyk35Jlv24sDX0LJTdOlgrr/LV
4CgyYgq0NTLVETBGg1vPej/916OLN7Mdc6c1FRh98RfDD6Qon1ixlrYFPH9/gZW4mmhikmXGoJun
yFQ2+EUxUXGpiRtv5MPdObMjZoHHMKJqpDyRcEqxTX3DYXprkylQkEvozLG/FMzY1OCzksWMnAmi
cZhdlz10Ck9aIQE8XOc+nAIOw1GZvN1/FVYKNblBtcDDxQfuTNyIhCV234mgkZydz1eYqxMV7RCK
Avu47TK4aVsjsoqs5d48CBgtlKtndaiVgLcNePoCTf2cxFX73eVpyRMX3aWDfv7dVcjQ/bVls3dR
kt65XrApRw6Sv+0Ao6r54P7aXJs8rMD4H8naP4f7GLWTKHUvll8/fn6WDvKobdfh+uxXGl2Tmmtw
/+DhwWtJZIqEis22kdms+E4O8BrQEFvniEqthDVljNcUfkp9tGLsSobwrFdd9avf8sNbMPrbnYMw
WiGGJt8enr/6KAnyBRoAYHYjg8GGvBHznZpe5305ssDV018F4YS0zwVEyvL22QQEjvCuTfTWRRIg
sqHjomDCZMLhqGbGEdh130BVwMC//1CVylNlemXEcmDGi2ueTKHOJPZgjQf2A0kY9Qd5yr7IhQcg
PoDNA0f2U//t2EWHZSVUw67jHrD7YkHCpZttfVanIcTgXuAtUBAAceoUMOnNRsbsUdm2TBUAInJN
JVWp4SKxemKjvqFouuLsPC9XePKJ6d7eE9Ksa5BgHNgjznpyaV8WtQ2U4BrFXZRkFTiGg5d9523l
eSaWNrdzIr2BQvApUT/5ZSgo0eM2OZBJb2jP4KnGEU1YGldUYDNhBMGKpg2y+dE+HPkoClNswEUI
yd8Fl4mIz8Bbv6/68ztrp8w0thnGWCnxcyHxIMqJbcRvBLUtAAnnlD/IFomiBBtWsD/jWVgmKwkW
l3v8h28pIm0UmnqK44HfVYv/O5TZkpFyH//vJIVwcGkBq2/hlTfn2hgaHljJyYCtymjAQlaIk1jJ
HGTPavCJIHnDj1ePp2Cu4PvO5ZQWcd5Ya5MIEUeJBUcLyf8mvh7xfyzMfblaSJk8XFzO6IFX/IC5
P+Aw9reVQ2jA98FS+1Fv+lfQt4dXWxUtuxLGVgV2m+CqpW05eJX4S0U70n44LCXmhKjnMV4K2liF
vBRFeql3HiUZylM3r6PmufZQWE5jIw7fNDoZHHsiocfcyffFEiDPMYMUabINFtQuN1RUNr8sxcHH
sjpVp3MYypFIvCQpooaL+bHGwG7YdyD5LlREl5cfpggreHkh0QepENYc+jTHf1VRjRm2i9+OtvHf
pXfKDONSllLW5LxU2vUzoWxdXMSxSzBm3UbR+pbQhXyHS7rta3Q4YdOOVI4HV+u/prPn61ZOw/Av
Drboz3hMMWSDi96Iy6w3A50Lj/HmDWHv6uYod1JwxxFTEqQGUtjCPkbtuT1egBzSBXU177ba7RiO
NA41t9LYlyIu2AGw8Day0D9FqFpcOXa+FtWs1UL1OCJK1otDm0lqRLtI1reDe7AIO9OSb/Fpsbyc
YGJKXUFPSCvQYlcdh4jvPm6/phQoqVwohIgq/hJgUoSyiaecsXB+RnBitMQg4IUQwBvkkIezWN3V
GHAZSVYdTqb7wosD5EEuCW5MEJ1rzo70XTx7hq8vgyfvq5KlIgMzCn6EHSInGeJ7OSgJA4ud2LmV
Qr/UeOBuQrbMYu/gq9TWNS5sLQ/iGI3ERTHhuZ74GjCvI13NHYdxEx98Kr3FHib2obtNjA8cOhVu
ilBbvQMcotvUz1Ulu2pRwZncrVEL6eP2bT2/R14Q0VfS3ndXGUCyA2FZkZDi4DbQc0YmOxd27vWL
tjwlVQ2ZatS1SVZd2cZ7KwzLwe1L4T5c9Rw8cRnaNCg/96L7Dh4FQYHjp3BflZBi3LLAcXL2Tm98
nVuatoMb8IsfaZQP+vJtJ106to+6XJX6bdAiTIqFz7GL8270Y6hzg73YJJlXpIltXGE3iI/WYYSJ
VWUhatPV6+7jsRRldoSsZPQki2nEimMI4AcgLcLh0DEHlsA6D1AQgiWV9aSE7hC6Zn63yOb3zBVS
mfE2QgklPX10EerMX8B9JJCQs34DaRxMS1ywRZfuMhPzN6LT40DKyvzdLyJqVdUZPAIXC8xXXltS
fqoGxW61mnJsSXMf094kZvEQvuGL0FpPLsXjrlw+ThYSCbSbenwQcLmXwjk0zZ55uy6dQ/ttcmio
JBz6V4NAzfFgIbM3V1Gltc+7WShrrOu3LGY7eSFPuTRuBg+Mk7TqLE8B5MeI/xEM7u28E3VrG6gj
cv8UVUKv3O4lmJ1nlgMWVDGoypm3kXRh8pxy02nz20zZBlSahV2HXQ8MAVWsoFnCFa8+DTomfI+k
qo6CaUHBWOGxQCr8yhjAR19bKgfIE3lvlPDdHIV3gxRTVFDbuHg9HtuzhwkTEWdIKAvLb3jusQpa
LsZJmUouyPFzXxxS4tVO/ncZQj+Z7/eMTIQAtqtxQ012PfgfBevwSwDhJkAz75X9YD8Cd46NMwTD
RI2BFV2nJ4n49KzulJD3UenfomIm398Vcv219+VpDul1zb0YhW/af0VUgJcNgufAL1/FBqbUpTqZ
zAbAlv7GSz24CIbaBe1HxkHrWrCCWsMMXVee8JwnFSYXo7y8XGcL7PSatN1Ij6keIApT/xj/LXh/
/5KudwtnKlI6Vl/qDhQesGmoYgs3zfsg2WhUp+4N/LXLXjSPJ110Bsn5fHEKNsb+w9SbHvms4thc
acAp4SYthdzDkZIKmOsyp6X86kPalKB8kFQ+yIRHJ5l9LcthElJc1yR5PygBxmmxD1MO9F1jkOqj
C6Hk3hCus2K3GwZ39FCOCTN+F+QYKeKksr0xq0pOS/9lNdrS5SnKWkwfgxBSjGWbRgor+Cthwl/V
MQem/dbBhH+XbH2ibSGQJzhWQybhzn9jGOsPppJFs2HuMF4XpuqxEHWnFFBrofjmOr9oX2O0KxKJ
8Fig7YKWtcXZ2fzma4rn/G7Z9+htZOIMqbttOVdY7vv7vMxMKtJ5frdIAJK74CY/E4dDiHHjFsew
MgVb0IxjI6BhCi++CIqLifBxUTIxvdoTuD9GkUaaTmBN3T/CCoiPKa6vzrvWmVTvxtXP28loKebK
+qISfJAC4jEITm2vuMp1EDcYMx44jb89/s9vgwH+ZSGvT962RAW7UZd7uAy/sML/WF7i3nPS+PMT
VkktTdJirI3jVOlsHvC5fzRB7wnBYnfqe9HYpwhi8ciDpDzEL2FQWsGHqsbJMPRM+FOspb6bBl/0
mGknwn4FWI9JUSedSsWYx4KJsv3V+bzZpCqwslQxwfT98cJBFsZZvgfH2FKOk00ayq9cF8jUJOWu
vjhv0x2nEAMqHHygbuddR0h1LG9Ch0dk1ggfaJDJiKhw9760jdy0vKqBEPRmg2PwnYlh5UiJbMFW
O1s0TUfGgw7YiR2GvYEI9hBxXge6x0PYgvgfjmNdDYT5PKzekBQrS+GQ6700U8r2VaWAbw+YDl0q
tnKjctAG9nP0KG/u3fW64SnR+XcZ3DTigP7ug5Ri0HX1NXDaOoWED9rTYvXQHnB0Pq7p7st8ec5J
LEANKPfrBTdxIVdZ2jdFHU2MV1xrp39mt1ibQacLxz5B+RVvUayAArGfPL4Lx4zLc2PuYLMb3cWr
4tgklOvM41FTSyIN0wt4S1HXxxAwjbc1qNOHHHD6/w/7uihRCMS2Z57fk52tvNwAZTZVRAi2UiTF
O6dAqhXcHOJ6yZXUrv2xp4HdIG10VSNR6gFqoKE1WVNtNZU5O6Fv9O/Pso25ycGpX3XnvWaHwPqS
6dQL4RPDeN68OgfF7mpKEPl0yZyGCsR+Ii1AYIkqQtaSfSnu0LXkLDqJXpe3x18bCqoH/U6r/qzc
roSum/2XuzRr5Jb63755N47+dz+EiugLcmbPuWbCnjSbcrzFfZACAD9tFlE+P35Fw7fpQUQB7gkO
sTBqmMKkrITLQHOw138ZagGmKJA6WHqRvkPFoRjk0YwDML4FbeWfDPExFRJHcXAlIEuuUT+mx0IC
nEV6/Sue/kC7kzAQ7Xv+PV57AEs6k/o8e4ytPsRmtP/ygSam0blU9pPxicEkesvhiCJYr778LCGS
biMG1HbnKFfXmTv5pwBae09uxmqnTRifESnhiD9UMHoz79eFgv4ogdbA2GJpPa1e0yVXkJknlwTV
1UlVcYyYlNUlUdf1UxKjsF4dytIKCCnnIi9ulegkDG3Gdl31yyDMQk6u4oVz9BQmU1Xj2VCaESmz
qX1fiaTWaxX7W7GVwcGMntJA/rJUvqDUaZSd0TNmo9s+EYxXcuzZNRShII5LR/kTqLFqVKQMOcNl
BWlTr91IaGdJ5L2pK8qYnp807LcJP63aCPLhtpV7LPWAeAk2pXTMctodr+F+AGSQA46gJ/ZKwoVx
qPEbhvhCTkFEDWfjVuhBk6aRCt8mWvXaAA8PVILOqxYUxCcEeWbATP5y7ez790KBShGxKiirR5w7
Qfkt1/aH6MoREzaBoaRcdvmmPZl0lpCg/HVUdEk67GY571W8DdQJsV/7/voEV3n7pmyaRqxD5Woj
T8/NpMDuaMm7RjtTnQFH2Up68l97mIRHoF/iFsUtO1TbFv0kfHfLCVQ+Cg6oOm+rY13iwWDW/Hwx
VVMWvLdq5hG6y4/KRnAOaMBww6LJ0ykVw2C344BLug1VGDEQTnx9ASdiSHRNByJlqwVkEI9cwixQ
EUfYs57hPBkFqvWk1hFyvk79Tkvyh1947arkNTIrPEuXgIZJv4hsP3JcBlnzTy+shUaLfgiCOTuz
Vrhs90AbNQkbrTYlB2jXJ5Lj3COF7ALxq7byJiQuaMwHJTqVf7a2q+Xz9S89VnprX8u6Ng+HN66w
puCr0eCl0bb2xj649a8Y5lHqu9k3vyFAXizVWOR6TURy4h8Ruqda1FQbjXFqsaSTxv+c+itsfFVx
vQ9zbCCEmakndS7gbKmBOsRMysJ1ul5sOke5wSZJqIQhMNcyLWwu7KwAA2X1uQVHwUT5CkLbI7FR
wZhbNqb2fEYIbRQldD3D2d1Ioj9gLUo0v9Vg/f5ya4f0DOMhJH/T9IoCV7Gszo02CWusbV+JZUnE
W7t21lLqvwolZJ8GFnYukIyfKZHhl4PSlskJLI92YdL843x6cIbwR6u5Y4FlyJgo+0J/biSkYvn1
+3b/gwW5moIZ4BXrJGz/uvkOo2hNMXk4RPDs422BFPo5QgSXKmJP1K1o71PVoJxQvy0nsYCtvgw/
umyC6+HfMhjgiXa1xEpH20V3o6ulbuJQz+V+/EEZUvyP7jDTa+cmXVO2YuuXytsr9h41u7cBcbV5
7SCQJUKek2BaeX2+hIdt6RkUuIl8YlcxImh34TV3r34R9I4O+40y5StoPxu3rr8X305cE70nLEyb
vUopsJ1OpTokcFJF1HhdE2Xkuc0A7fOvcbR2dNTFL+J/mQNOAifhLPbl/umCmBtSxfpeN/g7MM/e
mIjsoaI590vmsyA5Fx67pVEOfLi0wSeRlfJE5yZkxBz//bFVJDENGuaewcKUWhPhbrB+jsRMcMqF
1G41WqZ/66BrZTUZLOHHo0fan8GbwWI0G53bfJg3zci89xtUdLO+/+PuKfUNfNO7n5P5DY5EBDjh
t7BdW2AbFR39nznvBuman9croUJMokSag104fsjDes5yLKt2Mgtn/YUoX0nhQySXEBlJk8uwTDg9
q0bQRMK96iMIW/Bb9gxD2k2XNH6QZl5tuvUfN0nhqx6jvoIu9yfR+MgoMgw3DF/8IlDMp3azW9KZ
sL8pnTLc9JQ0vG0UWkjGHIyH4F6Oti8VXia+sda7HoORcAQlezOVX+f7PwtVM9rn2hV3+EdyeKc2
Od08LwHlHg6VYa5Z8Pc3LE9XCrrqNtRTFjSsxhkSKTFw2vxuRLa/CCjmT1DGms5Kn1suFuwEcreM
oStEc+gnCOmDG6uUcJO+fkZsDLSkjC7ePddx9a9ti1NeZQaXOfrHMoYqvB8gC+y2PeUm/LGLFrC0
nQkksMxulBZAZ5rlN3Fx9PhZjXa4RCUZtNJW7+pgi02w2y5W1eaOorImQjS5tGLlIBgTzjMUEY+h
W8zJiTLPRy3zZJ5ibFZjN8lGu5HgQcSAROYUacDz+vWjUp5PcqF/9NYRRWp8FNPT/4/CDeoXcf/m
UlBoE27ah0bGldiZY0M/u81Nqs/4qgM+TCeMzKsQ1fEPqTy5sd+BFHVzrOBl+RX5YKpDNdWJZIop
ZfwOKrggUhT5hkI8NvbRcIJI5eqJuDJMjNEqOfcJmfxbG8W5rVO2cxHWsgJ5DKX3H8m6aOvvHIO0
0gRy/nDVynBSHThg4+FajvPGOwy0b2QoUWHBNMqFcQ/bJcLA3IyO4Qxmtvznatwu/ZahoNeUnh/M
noxRR2TNGkSZVGZKCPCNHI/XBbLlvO3+/6WlbrG2mcJDxqVp8YsqwR0HhT2LhA+5tVa7kivxw84x
sl9OYIkJwJcMV1/uD/MpX2Y86FZDfWz+vmg2rqx2a/UwM9BNG3QZfmrNCuUf+7vBOMP9Bu5gGV4U
WoGsIpvSlhvm0o4feqqzyb6fBwptn+o5IkCmT8qYVKhT0fOkNEQQuiV8zzM02Ch7SDamTkd9T8AG
2ESbVERH/oHo2bMY/623tYD17h7FAYki/XSYOmpaI2IEZNb1dgY+TBu9Bsav2eLeQSfxDiv+GHkC
azo21Y+hC4j54CP43ZhNSZMvHF4fyjyzr2vz2KJPl6Bb4LT4Tt71/s5GwHigOv0A6KFRaL8EsSWa
M9B6TjdNF0LXcRUWyv3rOko+zL1rK3ldZrh/E/NggJS5AWHdoReRuqO1cv0tXriDFQ/TxOhH/toS
KwvT2xL3BUQZph7vKifUvEcwEoIDOjcwF7Q5vbwob0TBR7KMOBMuWy0A3GVBJlOf7oVooukiW9IH
Zr2brWLIAPfOb4TNVRSxXL+9WZQZkMFTdvgAvqcpf2aDCG5EdwjdnC48yKsUvBo+2gYaqbhEU18w
Agw3GvGGee4s2X5/5ukk73toG3hL1xr0KMA15iYmyqLQcnW6lAzFMEIQe4vAc3ktsqrgUeLxIX6j
p5dmcQXn12ZfMfiiNULO+75SUrMo/e0h5PXaM/NlDCtA5F4wNl/kyKODPA8XANwQLc0QJnw77vG/
4OzjQXRVhs+bSQPFpIMiOg2tdU6KDh8GOAg82N+ckQzmpdjw03ZGiDoCuj02A08C7LwP6pgWaAuO
wuOxMQFY3+HBeWL4yV3SShvVdiufotywveX+bx61q0kx8o2E4cq6K/A6u9fPkpHgQ5A7mc3qxNkJ
4vYl1T9qf+64fKX3FUTmaTvO9zOsZU+AKT93kPZkg5ykORbd1n3guciP/lcojGH5rj9xfet6SeyS
hgxc+07BHDATF+IB/1JkPnl7d6gbQCF6K6GDuFirHTmILmsZuYcqih8k6fxNkCMf7AYYkUgk4e8m
nYgfFQlNLgCPSWDQED9EPC61sRoEp9I7isfwqgOioPoNkkcQSlqInqr+ccidqHajoZtTbxuqm0gu
DUM8IUt3OHgTDiqFTcHM30GKakmYML3+WGkZuFZ2/pisC68n1VBq2JMuU9YmLJrXgzWMXbCic+qP
hNgbPwH/zaCCFbn1NjIZvw5sysPRhGt6f8nF5KtmTMjmEjMV0HM/t9CBpdct/T7r4WgzVsU4fFMo
Fx4EJtQxAfVLh9g4TFpN7L1Ovnnar8GppNDQiFFQUYYcFZ4dGC1YETTfhhRMHKOeGyhDnI0F6kVF
Z6QxIbl4HHrhQ4mZe0doRtjbbuwkHDWKdoN10rrYvozUPfU/8ydE2K1Dw5iKdIC53e4Ers+N9Q4x
tr5uQlcWPvQwmIrv3bTy1wzA6f8uO5puY2CtX2U0DeBCefnST9UAgfkDKTV+ylLR7DIy0eEticLh
mk6wkhdd77G6ZHBM4Sk6ZKdDyCEJyvHU+z+HvMth/XLXT9TDrLgR1Di7+Tzxt3yGH+stO+Lg4YfT
z4VHv6cGgbSQbsiAMxB7g5LGR5nmmk0UOvFQnOMo4jOePY1hLcSWTiHvQ0eL59HtuTdQMpmW3WTk
I1BjxDHbmX9VyQjU1DfSmHXo5Nk3uwhu6M3lI5Tz+uFIiSFjbvn4dsJ1U0KtzQbcEgcRvDz87Jm9
r5FbWMfqLdnNezNIS9J3YE8jlbestUtruArVNFVnTa9cza1+5HUU4NbDHveXPjMGDwDGHZWovhZy
XiWrfxXv9jFwNbhoEKfXwpRQedcEFfadxs7ZIgTg93YTegvAYREWIEHGUc0s3MJaA+X7xlYoDbAH
fO6DviN8VdlzH9WYVl8BFgHfpfxj7aMDZCoMhkUXoAiml5QwdajOSsQ3f1mCdr3B7Jj+hzk4seAh
y7TGIvK/BR7tHIU7+yaEL2XGP8Aj1m4sV3r80ucTC4WSwZfmadFloquYUmg7t4c1zLhSLZLLJu+6
u0RwdV9nWH5uzOO27Xx3TEiRrr5//styXxDJmA0dFvTAR3oYddaohvnYvGI9u6kfwliVk/oN3MFU
vW2WGVqaFGVCD+i6CHLh8l7BUC8OFHJnVwCbLUcWRQjcmPHRQEKsv7ui8sXeLnKfwfd50C1B0dnN
lQh0DwmejCxvrWdLBNHnBLHxxuW0PDLRLyI2LZuahOnOltNvke0mi6GRcHihkyJBfufg7qd3cYFb
xNnqa/XNQkGfuIdVvtJ+AGwC0AnSVaz/H1W02AMeOA6EZ4GjoQw9H122PBnI2mg5MHoL9uBxtSr/
09XybwtwjeISWQUEIFwD4prkCvHKbgdIDMP/xbAV06eFdZrwfnVoKVO9FVif+f2p/ES7/Td7nbVp
5RuCOQ+G162EmIZ7JPn3G9wuCNV0KCsxzSbBiFuaT3m/1eGmR/WjtDG+arnGKxzGhPYfCa1fiyp+
5EI4tm9VchpWSlDsASSkvtrZEQddY1qeMJB619iu4NfPksxGWVz3PiR93rkMoSK1wPB5P2YeJISY
xDmsAmllsQTIhILsaGrRTJWOvDsFBLrY/5GOLvFO0OcGcijLByuP29pEkTF2WBMWAg54uMyfnDAT
1led1t/dUUvYU3OBcLTAJBE88wTfcx4NU4naeShkd2fbxP/e4CdrUIPHtiOeOBJu2qIZdedLxnyB
87x7TivhbQFPXMEFlR57CCUQG8SrhjdQNvwsnIHxqYNwCFj5b/4lMms1OgX/kwyl8vhE7hTjTOij
U5z5KawU7VjDtuk2BeyThTSe+BOpmN861BjF7gYy6qr1jLajB41kuQBmAbGI3sXXklDqafFVAI/P
65QIPylfQW5vNLoc+Y1FfLJNZmaryeTWAy2Nw2kjnat/ESG0er8TmjjAYTAg8CVMh98lDR//F4YU
lCYbseThaBLKv6+R8NxK9I+SB2KQ+5X5VP1dcAqHrmcLbU5kWhR9ClUMaCdAb7cQQtcvdKESQBGo
gXK42YQjkz5g/EbbU4NXsi+Q1xch7NlL2HQ7V3HWE+pQSxC2oS+p0lRqiIB5E5HtPPsHK6kYPIQQ
easpnd6o1CpCS5nPoH50Hs8BDafMGV5DEBF4vgo3EqeYMQSPjGEbD9O+NRG7QAanO6DhPIVAo7gJ
G+uMOXBReRqWBds5xVtdrq834gt+WYgfOGWQmW+yAn6OPZ+uSDHmCHVcwglNz3U5g1KcC/McY+qn
bpSkq0hAH5hQGA7wP9u0SkrpMcEnlLVSYieq9SgVLXx5AZuBGl26tNrycNGJO2m4knjmqCzu+pQA
Q/pNIhBgLwNLpH262uEE7mgkXg8EE+QOOnm7okAvn3tdyAx7QiDRCINPK4Ghc9pzQV9+6o+xizAs
4LZIVCKa76IpsHuXs+Khib7SkvYlH/+ShpTlI8D1v2mXOjHNwTB2aEoe0iHTPB1LOrUekgdMFmJV
Rp2egeEI5MSPIZqd30fmuIJqZQNPm8bjeCUskISJQqyGbmVfGQfrgavNkt/c4/g5v9N7K/r1KwsQ
vO5YNTqMowlT5bQnyGBTvoglRtuBrkJbEcX746u/9jdx2anNk/3mCZLb9QPCRj9JC6R9CGTy6+dG
gyzFdAgf9U46nSRfOK2Tzon6lix0b0sqS3FWq0fvqMdqqzPrIfhvp2sRbEv4W5yw7uMHfhcTYYfC
K4lFyMeU2v9W6bx4tSnllqNV+eVJ2XklJCphicmhEvpVtmAGSlwCi8z8KhMTdNoWcZLnqysBvGxF
1owppm6D/l30k827Fln77r6pj7wZVk7ZcOAgbwYrd4l264FWEQRvdyi3idX8JEYCPxWlda6C488h
ic/vE984Aovuemz6A1EHWE6qi/PPxmOCuB67o2mEs7YqCp2B1ceNgVj0c5n8WSgbeSqj+pU7xWHX
i0cHueQbtoBw5L/CC9+vjMR7g+EX8Em7RH5LUbZ/N3yW9NtTlR1MpW6cY3MCM7xGH4/Ymhy7C3yr
9ociJJ1l6+ttHUsdh4Gl44VBwOyIGI1o11fIfN0pTS1jweqOAKa3wr9iG2PIuMAr31EKFwX1MowV
jGr31KEMqJ3KPlY3ipNbvhSohtbtz74fZ8UGzWfUld/I1cAGbavI4EANw04XFEMGAaKLjoGNSWtw
yTAO1CA4qkhwzXoDjNbbuKxtu3herFW5+sWV0QZm4Z7F+WSQZ2QYAss3X96MDNEvHeb3fXGz3vRW
SyydhVrzbAEYhqjW1f1Xw9bkxH0oNdIjb8r05ijLqLvUuIi8o9oKXkWTEMFURjXcq+BAosJftpTv
LGDgKg1ZjwMCArrl6AaGwkBbZjw75HFdKUJw1aVKJQRBPx81TmcfTH7GJ5tgABTpReRTuAJijeYf
kSsjZ3lXqI4UdIj5GtD3A/Q3gGt3QMAkVpGiyqN1Lm6F7/XmkYzPrJi5hzXTFjvJfTVSNY5Rsplx
sFyV2Yrp5SbVIfJZZ2uCl5rQG149iJzOHYr2cSRRo5ZwBOm8JOf0YVfyYpvM99gXa04pEu70p5wK
c35KhCiRxP2POuO6cEI13Rdf8ciCkzevkbBIJGo3+4kKegj+ax20VicZM+h+oFZTeQF6PamQvPML
FhVNtp2u8AFE6Xf9qo4c233M6rC4pqQvv4GdwD4wJEfHxqylbEk/SDJXsQ3QOYrWqmkIt/MgHpa/
Fosd9TZriGenz+Ki6Q+6N1PAES88QTBP/8VEHhQ7d4tPWfi6fPfQPrEJg368/o4rRH3S17rSvdRI
/eAFgge1vZNnSB5rTajJrllKixc6JjcAxJmhWeGqWLqqcsCd4WlDkmx+veA0PufRFxhwor0WIm4y
zwoh59g+hpEKxzbSiiAA8wLnLXJ+4AZW9ysEuF1besbahSBCIuIoq7U4R7iZoX9sV2cFKBaORiEk
gBfn8aip7j8NQd5Lbs5Dhz/6QK4QsFX81rBIPYXRpuAloHtVauReANbr+Vsb0b5/ATgIzkva+2oD
p2Hxajpze79UXa3IIhjheM9Q3+BLW1FycX5H+3ppBGvPdEr9vdqrn4JaJqxDjjszIywdK17CtrR+
xV7zqYWF8udco7Wmf5H9hI2o95d0906K+9yy5xA6CNFGgrwBAJvkOAqSgLHdF+IYdxw/VJanu+IH
UWML59Cg7kMkxTjSb5bt80I+wAynyOJ1FID/JNjYlufKdKnBiZynlqAHKmybdJbnhuIEt0LPiVWa
5V8Jjre9kMz/5dlc3rqnTwgPzGJWx4OP1GaDcmh4QClZNr9SIPhHmTlrreOX1AOQsoXyRI+nISl/
WJbIWHEToy3ZoxsrRMiUwX7zfAo5rK+ZdtcVwlQMct8bhi0Pt4v4ZGp9vqrp9zfNPWg7HnhwoaYn
uvks56OfWx1j677nFZSCJHwapFo8fQrqc0ejFdhO3S9Ab1rM2u85f+oGI57w6hoAYHZy1uXC7RGE
5gB4Tgy+TWZo04++upXjUdqLBmOsJ0uaPhUEDZSM/gxxkHHwV+8+1TH7cPIeWuB1OHH/F5aMKbvT
cdaUMbbJZmY6qzmEWbHtQFDfwDaXc8fV0/9bcoTJ/lr1nEN9d1/qcCBDJEaOQsqmB/wVq70q4K+0
DTjhLtE5VecXrtrtaVkOMXs+UbACyNXvk+2t131mH4+VYPBtVPjPOL4ALLS6jYgf1vCFLaJohgZF
8WlGcNn3vNsH1WXNjfM/ba4f0RzV0+q6DtcevtLSNK63F+jQu3iMQkN6IDkp91H6EATfzELUgTju
l3Uc5h1o6y0jv1uTra9mvYngwYKQaI+1iwt+BSNlg+6P4kogA+ozLkG1/fvP2brDgCnxOKkOx3CX
X4cQYC/jMEuwkdTlYAuvM4EQJk9aHFvyWSMOwOir7FGd+p1AaIjNZiTOm05O4VbGwGRj6sDyrwPk
V0j6eMYGO3lmS4qLF2s1r8rnYwQihYzO9+4kuTMkSej+5Mq0P1dUOTMc/1OH1I5kps9XlZRsHTgL
9QUMf6yft+Gkz01Vz3JR89gtSHa2LutFvVmevq5uRmDBMapIr2p2P6OgtwMl8LFrIDCtfaKnxZNb
CiqARc4gLOStsXsYsY1UEcTDYXxH/B3Cbd49EfLSWxMT8V3LWbYppgta3H1RsLSJDdFY5hQ4ni2v
C+3NrfdTGhA+GRwcrtaLimW/8gV9fHMA4FXXHY4yZqIFaci3gQQargSiQftN/N7W1DHn6J2s4E3q
jqwjRngqmRoPjeaoveyXmQELBeJ1ZtTUVEacFCcFpKhl3FYQoj0iVMXAR5BxqHAf7RK5mF+GFipI
4jzxJ0nm9nunBrzppy+5hjT2VZvrf/yDzrQdyH5hNEd2zzitFZrzV1M9vbXBu24sCHgRa0gG226M
BPjskvOLwFRxwk10ej4vMZRVn3OAsrDL8CqVkN61ApDM0L6xdVbD8+QmMIcqA3ssEcaNwnOMICPo
OYktJZbG1WQpW1M6FhFruxi8cH4WAkNHtNlzy+O47H/5buR6vbMF8YaqklVoeYXtMomlTkZ8QNGW
EaQtsXnBRLF6jPefujn3GC7fZu6wwPvRRUxd5BEgYIaH6LqtfArIrjWjDOGzsrH2HyNfRI5rd2Rs
iYhmGzcSwqyO5qWWimnAo9Hgg/XYLr58mT2+UHFozrOKjiqOTETzRtAVQDSb2d0GmWqrIAMMtryb
YXWz/I3RnE6DTvqlU7uF6WG/qitJlghr0iUg1equSPybOQ8uYfH9wmRO/J705OcdvHnW2VXIUSUM
8urzz2vDQLll7aBEH7JIKQWfEfsf5usyhh3yxGYVCMrwAkpil11gKiVn8OTeoeoWgpq5jeiShO0F
5nXE8ghfHBUbyh4fYfLuD93OUPhGqvGCZG+ro66iLHErIMtyVJPslw7cRADsww3bILAtsbLVy6c2
7u51Z9OoPPeyLKj9r+5uzZpsIpNcp0hNyn0kSQ4TYh5mAcrea+mBboEp/TvYZMbb3urpu7ov89JD
KynSfeypZ/SnycCRRf1ulgs9RLzVSNzJfPC8Toh9mhgPEH1dKhYYv4n5kMn6Ic0CyIyf/2V0lRNg
GPNfe85iYrLT9B/ZUCcruKLe4PUoDuZ3vXALSI1U1jJ1ib/71OBigc8TTLf7VAtlXnAQwM7lk9kS
Y0YqUTFNoK1E6bUVy11ZmpGuXWA6FzsZl4BKEXr5yKhtUccEopQ0IdTWLntyDk9knv+EmzinbJp9
9y5lUNHMCwsfaMad40pzVw4cakaLYbj6Cyidrox8lpJe/q6VnqfRWvlIJqvQJ+pzUC6H2/FhnCz6
Cc6C84fkKuVwq3kzgFNNZgqx61NyqrseT+h1E5/RXtJLjr8iB4MUSfG2GR3LkQlcE6LVlx14djpC
lXihx+eP7c3wUCTiOztMFmVIB8BjvfckB4xeSUlSlQo9fNQH4d3pd90D4sJGkLchy13dvdkywifm
Gt3Y49rSWmISJ/cRZRh3Cn1zdx4ph2B6Z7ebgs0Jv/bdqShtkOy/aZrvYsaO796OVy7oDtylKBRg
QUizY/rRgk5JRVYWdLErW0u36YwqYg6jdzR9OJbn14KWhPNXgnUI+JvKxVGtKSgnIziC190n+uZp
EHjMVbz8jx1wtrVEiyNo6PUYPkvqbRv5K+3ZCx325cCTrBnu/+2RXHxXn4rFqZ8qWfd7+JV46ndp
N7JFsmFj+J0PkB5+kCEGO7R6sZZWsx29tpmYKele5w0efYz+hdvIvN4ZJ1vWMlU+SJsc1ZZgkyU4
QTpnCMJQ0Zerg02xKV7HQADjSeEx5jarxeNiEvwBEF9t2HA+LUcErZOe9+00Vz0kvKTQPCEIbxzM
KmVnM/kfZ4XZi7GEYwHZ5qfbUjaeJZpS5R9KELN5BOxtQ6Kia9V3RHOiNNaVxe0olBTGa5tJ5gSn
KhyNGJqYaN9QLtp38HCgU16/jER5c8tnW007LQGqf4V6oddLZ1QfrELkVD9CNg94UttgGUPUeWjx
0RdWXGX9yFkxSEIMtynHbjSAJG1qAP4vc6lRXMVw2x2itqXGYvRNPxItg/tsMfVZ/eZjicapyjHe
FAKU/txIgBYhQOOHsQQTFPv+zOJOAvak36SgR5SHokJrZu7DsK0NL+POWYT8xFTQhTKaWR/YeELn
hZxEi3d0I36aqHqmJRDi39cqwekLUdnZBLjlzk+isgQCBnTEyhRvUMMMH5Qbg/bEtpnNP7EOot0o
gj2SGJsxiPJp0rxUltF/K6TxRm4kIAijfkzfGxLf4StI5gaZLtLMaKjZrjG8hckAm5hTWLUWYD0W
HDoG6rFQrJevW/fRbKHefESvBv/B/rV9UKjjlasHI8knyQGJ88IQF6AT3EaUTIHl+eXoF8S2VyUh
zpRv7xd0+YEHx/ixqSPLo5s3+xOIHcqSnin86XNIop/4Y0HE8CtJqzfNgqTHpNKawRBJBXNgiyI5
14l53yOVtypXVKMpQm/SH787a1LaogxndnqmhxTOtbBjUMJDoiLvVJoOF4uuFEpALg8aOBT6f+Jp
c11XNGh2NthyQsDkCQ657eI31JS4cboS0fv3rjpVj7QxigvGNczPpwBMF4C77WsxfT2yATvVT6BI
QXP3v5b4UNvqFTz/AiR1ijQDJ4Oqn1c/MkDm977jdF11uXJxrAuiZvVO3eX7CwI4oK5iHsQIs8xg
VjNoQ2Pwl/ScBWCHCoKbPo7PKaO8SX4f5wpbFdf/xrX5HAvOm529cc4uXXq4572fw1qkqWrjt5dr
6T1H0pgY0gWQC2+A4vra0ZNF8gckp0jvc5tGIjuWMMUGlprJUNsUXgCPT9r92rq/5/NcGCthGAns
qah8vIHLgzZILzbqhrHD1/9WErR4qX87A+8RZfEtvf1Bh6aUEgmuENKZ3VuzT30WyHj7MsJtX9ZY
hKN+w7ik5L+i3df4GRP/VkV9irCLaOYXpb8ywgJR9jd+BjSFLJT6kSxP6YCryBNNn00kN7txYzP4
EhKua79sYv3AJz1Mp+2vSPNMmDGDN9FQZ6u3sXwY+LASUgr/Stxt9kISfEPqqLC9HANxbBHmF1tI
ptdKou9CzORwxoEqbBDWNdRT4pDrdAITATneLQs1DK6x1M9LmiKpQshRzWp8GkX7bU/JPdHyiIrJ
ANcxzq1D03/34GlLxDs3MsnXr0hX4t4spHs4ox/Hq+Iktn9tzQf4d7lbp0Ewaw/TRfV1zf6AYeju
LYQBqVW80zV2gHGIIZ6hO8uac00HhxQfOblVXhZ5/9bPmZ09SvEKNplzHUBWGULFg1US+6ivRrg/
NRw0PtHafWgH2D2cSzjW7Mt4A41Y4FUwxTKt6KcgYmcClAcHDdf1t/A25BUu0uyp7jkZsIqw6jfN
dg5+XdHUTZlqOgr15+/VI9gIJ3ORHQW0dhJBIQDQRYmIn+pQTyambUro6kF0wwPOG2VsOvmbPzse
br/E7r7gkMwSeyIxDgUaRHdSwvkFWK6YwTWN4t06ou4hILJnq5tZRYCkVMao8DdP9CBSjQdrhgmk
orJ5rfh/qyww8NdZHwZtrzwD1X21yPIdyaUSbuRRgqcAEiTsHKsxJIRGrOoFp/9UgGLgB/EI9GpJ
o5XxdkW2mfB9dh42SsZicgB8blyhF/pJQQ68PNi0WZBaajn6S34PUA2S77th0G+CARGnDn/NjK9c
oJBjxbZ8mfUszMYCLNUS00DgKYiE7PSN8py3uXTQjir+dNV0fewq0+G1bRs2vV+/eV3kf3w4m+q/
BIWK3wwTs2qylTlIc73Ge5BrpKuiX1+6fFYYqoisN6TlwEA5rsDdDftjOP1Nv9NzAnSHKRfYG8Ps
QtF+XsnMGu4LFTjyfOENdIle94CxL4qMAgY1WJ7cThSfsTSq36iLs+lX11tVREsjy9udVU6TdgV7
gVp30pnNmra5RbbFcmZpYZlQaNjxrpJgS2b1Bb2aUBqnM73qEV8fk+6eejBBpaT2pYfmIjgFyO0e
8Ak1wkb22FUhlDVoItOq9pDxa4kT/BVwkb5jsfLHwHjb5HmblJDxQhrXWDJD/IsuJbtp9jY/o86p
NAOGhexSbTBseTsMWcK0/A2JVk6gHu13DLzivsqjRJaG6bsN4TQDlDBSxG2N2VLLtyP5z3rYa8Tj
K9M68Muaw31TVqcl/aS8pYCJFX1dueAf42u/NpBvBlUKNYYJ1/laEpeigfigLEVfKmHhvzh0jZqy
xGAWkWhnKzmDWpWriK2r3OYZiqvouLodmr9M+rNgsuv7wCMJuQgq2YdW76x8kN+bSBX3A9JofMzG
NUcKcIE2M+whnV5h9xEAdk8o16zGGSDZObIEja4Bvd2YrutvuY1u56AryMLP0ghDFl9A8tKDNal7
pgC1xQiYI3MEg1eTWXEb7A9ef53HDkDE2xmysDOOMI3ybm+xVsBe6zQf93o6l2VDXPqX8ugbO8+p
HGQjdq+t066R7fprwteQppACHNY0+4EyHTEjRKD/cFWgoDRoMln23v8mn/znC5zEmzu+bOd4F5iR
t9tjyW8L006Aqml62abTeVhffWsOVp2AExPkU7pmZrw+fDLsTRMY63aZCzzDevGnhKPM9hs+jZzi
8PzSxsbhH59PWdBadFCnQ5NJ5UY15CirZZyCbjxuT2qS0Xd0+V5MX4F4dHG4Okwb11t8HyxuPgcC
7xWfVwFo6z2aEYQ7AlVskt8qc/iYYBmR34VdSXvTblgmuqLlFjo9PXLs3hCNcmUYVXVAEEDAOKE6
AOZMlv1XaOQi+8Pn/e7VPtbfCMGc9+idMntA7BLQ3CAjoWiQjWEEvFWsqo7+Kpcsh8u9WBfKGdpD
AwTNITH7P3MexuaIukL9/Bq2wPMY0f8j469E2Hq12q3IBgNBsUHO2wQ85x2HgIMWSKpRaKTZvsGT
qwOqvujdFikJqGxlnSEutGy83FJcvfuP6y4biKrAHkv9GkvugqE2wPZHc2qucgVH4EB7n8MPbfdo
gZ6pUWISlYFuIVWhqIY40hfGInaDFEOLiKt1kYZ08PTwCZ76HzPmklkT2WhRhqOBaePWOv3Z0W38
jJMTjA1atqGLGOhfKxoU5A0iqIWJtc0bqBovNSgMKA63RHzQNaY5ktLcGDkGW9i38721gCBhqS0T
enVPSkQG1AVpi1VYR99tSB8TIe61c9yDeG/Nz5ofE35yZ4DW7kwaeY5YWrqAOWczrjWUExFC1pVb
86/Putd5VRcwb4JmWc+h4N7urFsotA8amSDfaEmDooRiDaVRmwj4rE05otNHve4am3whC5Tb+jVC
mV9nL764YbKvm6g1fuh16NP8cCyc5dn/s5Xe6rm6kcyHYyj72KlbUrF425fiC0Bh5V5oJFxJFNAY
UbgRmdYaHRDHezZvLlxAeTvy+i9uCiHRTBXdVrkAcPT4TVUqPBJCO59ndIZmwruHAPNjHaxIyxZ7
P/vIJeiNfb7CKpVjn5K4lOtv7W+CTXrMhiJ2AD4qzzmtw256VBsJNAmJPL9csrWESNLegVu2/PFO
l+dySy9Eq0UIm+VRIjB2IpLng/GOJMlKmB7iZqqIVmaYCl83Gbx1gP9CW5/EQCVuhmuwGUkQtRyt
lnIyIgSF4aG+xXyksy/h8UrT+6Rw1kdEbLODm30won/ezaqnq17a9y1f46mktml2y895UqPaEMR3
hM9o4iBX/uxy2PCSkSYlVC3auIh2pOoyJ+EVHcyMWSZA1dzRziqXy2LY4YhlYY/E142Gutxjatr8
Da4dxEX3eRO+E9y0SJmsVqe0SFBk5bqu5Ep72OHKOxm5AS27v7tqRjwuxKvuq41oJHr+qu97bARr
WFj3FQ0AyWFbCol24RxFOx3pyqprYvl281LTEMg9F7Pqt+zzhPG6FTt5zAKrbiWqV1vpAc4vHB6F
rR9HzMs+FaseFC7xdVNeTA8I4k0xmXvexfnu2zYWQ64P7lWkvSHnDR29qHrlMCfpvVqxQpHew8eg
dMdDkebfMLaNRVx3lyHuDfvgULmmwfw7MXYKU28pXJ20kDu57bHckNcjjA+RmKymqxhhCoiRb5O7
tWUFjc7NLfU1kWqg/1EjT0cugReMnW/eltv2f+z1i5Ig5OeJnZClfsc0G+A02gOfGZy6vs1S7aMv
RBw83xP9HutFk+9Af1jEzYmAVvwsNWPcX73w7LHPX0dB5CqkWDMNa8J0cqHkaViOsifXvdrcZ1dI
uNFRtwNqI+62uLmNg0kCw4fi8Od+L8sj+c/PTQ9bK6aPrGSitwebXj9/kSSiDt3KzoFXpOoLKZjf
uCdfiUAEtUBG0ypv8EJwD+6wQnOJXu9netTPQ9pCpIpjJ5bi3n/WsYjllOsY6Js4ix7r5+YVhMaI
Zdsx+odEttet91mq7AKvQ5UnRlNkhEwxGq8ORmfNRi3mZpuGDmbxMD29CdmmHeVaigqojRiaaGRV
mF1zfbRbak1cVU5Vr0Qg4xJeRvqqsDxWTnXwmCm8CgIAd8z6fL2BP9rvSaGL/HmtefhTPomyvmV6
VdX/8oarcwrBgUs7WXvIWEgqeHJANaxIZLXv1ZrK9QDTiXG1CU4WZsRRnPdOh+YrtFCtc8dNc2X+
36uKdZCdCvg+QoXAJ97Nz3E0/KzXEglae2njjxBnB7QLQI9EKKuPyhaINSfKJ0X6zdonUAf5qv6M
64wFKxWR1QNjR1ov7F0nBXxZTCmJH8WBSwcqCzm+NqPMWvDylZ5MHLTEF1yQau8W+upojrdhiuEG
v7IQdAYACGtZPo2J5aXb88Pc7ms2zJJDce+5Dd9s0vSqFUVwZT3nVFXflLXWQTW1vXUBXOyyLHrz
U9IHsE1d7XYi986U+IPwxUvx/jp1VbqaJ/HM2iYcYlzoJBUoN/tuam1S0xm6BGOVaapVCAY4W60M
5UVU1KqoFMYIuRvpf1HxeDqigILxSp3nzkFc6+07jPK7PIrkQFOi7KMVPu/aF6g3hDM14TCnlL8J
3VOJiBKBxWoicevC6f/Vbc2SNVQPi/mPWw9dzAenN66vRy1QJwPsTv282xXe4xRw8ILeKDcfhICd
LYMpryEGR9Q6Sgrj8+dbHzrb8TjuvzO9AfTxQji1nFpVrFZHwRadYoIa1N+F6Kf/bBWJ1yC5ZwLp
1pPIU82W6HPrvHkbr0WWuGDwXDo7fYyd30VxL2OHCsD3s3BJ1jCVZeSVPtnjZwSoCmZD0gHwZYsP
wvLWf1cEw8iipCWIiwaHVK+evdW6IIzvoNR7C/hDdDtNN8JLsGjB1VD4LOgIqw8j/IJcQf7P1zeH
h1gEppZwe2nZB3/qoCRwhB/gDgbvwt3NdidF/JEypS3iSuAM+TyADUkRtP5DDjZinWX3/I2LNnLX
lPiUORxqi4MxQFWou5jBrXXkyzg3PAAQGle0f8dOv5FngKZ+9KCo+PQNdMfgzpUIq+Hxivc4F3Gb
A8QNHYsnwo0kTv0X9yS+ahH8rDUW8WVYSceN3/F/91l+3IJnln+dciKSEEIB2wumHyKJ4H1jzxkI
H+MLl9WxK5vvVmeCQGN4XD3qcJHPRIFNMx7H9SL6KlXCP9dS0JZ2KKoDCSyr+rLI6YPPp99MHPZH
Dm5DLLCO2nxiNgAmbe4eDzXXZlvwNp9xPA78T4XXBkie1l90/V8ZN9KzT10DZuwKv8G5IcSxnS9S
2bnc/a6gy7OjR0LSa3WbV/IaV3D+AKoc9bfJqOTU6qRXgKRI8WpqzKkOTTjmC7N5MFjeshVfEz0f
fTu/vhV54Z1jPqYJQUw5DTKV4eyrr7G/bjIXQJnmNU6AM2LfbcXhNeq4FOWMlg4SYB/t1aQEJWhQ
SlERdhUwgZNEpOLngfHUy+gNnSlv6shjjFe96F6oqen/rOWvRkh/6Axuzu3QixyQPspNXmX+8hxN
Hl/M3dlzfmpe/SJLhBpJucjxTTSLrRzQ/mSz0YMY7tRtXkur1384d9b9xcx0OQI/m34IyKf8IcjB
Itux80gJWMYknpuVZOBJxh9miZpn2E5dNR0vRi8E30aGMrQ2One8PNW660uoAHA7nCvnevWtP8cS
xnsAyaUtV5GcAOZes72rQkGYS5bouqfv+i+UPiXdL8PK9cD/Ue7NKAlq04gft0U2SYlTIVPtMCk6
UCVZjrnDvp3Kb0j7DlIEtfwFPwfNpUWxPM8uGwdiax4fJutM0l58DPp2cZGh0vfiP7UMjF/KvYV/
QN03Sp1qva6M8f+/lLLGdbBrayiJC4mnpm2xhdl5DncljPWEGAWdQafloekP2gdzFuUfej4IpaeN
w/MuJpFCrkQne6SRLHMCZ+HLDC33MgeOmPo9Z94vJyz+bbkIpiqc+k9y32XDq6Rwse//CTo0lGra
VjX+G9UvsugLIcsr2kCktBOSGeGTW6S6viV7ppX/ldoa1BM+TYlqzVTav/BGqOnp9cSdiqeeqYyw
q5oSTFZOaLsItkF+vryLvkx41tVxtyZ9yJ573kIdG3GCsQAw9mrI4kEIFgQE1LkS7atLfnEAWWwC
M/22z0MR6ZSxYrMDYz8Vut0Cn1nGosDHEXncRARK8uB6nrogXpdiFrbJ+vYjcswcX6uceCY1aXoY
dqJWKnwQgpip1fXpy9xWo2ZgyfydziWh3+oeJDyxcRrdp98sjvGdUuHdMaJ0lijmDHaukmrLsT2u
y2cpKK1iBkgmrUEB2GS4Z2JgA1l1ITjxmSXPUaakqrMKtWVR6Ae4cuHG/f03FfEl/BmcFwKeS9ZK
wC9Dd+0Vd1T9iSufo30iKFplQYR0gp3i6Ei8YzxcHBdaLd9BnSdimUOio8YP+wR2bih6ovfEzpBw
hm1aBEDI7HaL4JryDsi9rlXpCSRYfgVCAFAbSQ2QTNjp20KGkJqrO+o3c9D44+cdN0Os7oAuVkJS
pL5QCVP9lyXT1OERuzzFkc2qf9iHMKcWUEbKtlsUI5uXJ8Swi+EwLqL0RGzJaR/D4+w3Vl0viJA6
SN3Z2Fj23jy/pQbL7n1qdXrzEBNqihEo4pY48UpxG1Nz3XtibhNQsbXqj60rFYnUnps9LVpz+7nS
Ejd0fxVnUF2SaAgyT3lXaeBrBE1A6N4e6zTqsJw5JRsiOvrhyuHY/5KMq4kA+P6P2ALPlAXGgzCp
vBVHCnYqyBQ6oDgMeCAK1W/zNaJbz2RG68Pqx4my4HQXfx2YSsskhnxhdzlCAY28TrFNNlhapsJc
CKKJFdPHSyF7K7b7AllShe5zQVURCJbXel0XXKLBI/NjyUivPNOd3gp59Rii6aEip2AEuWI2gUys
S7ipKnigh7y2sJzQEkGmffY2QwZE4uMsyONiaLNxabyDaAZp7Z3jx1skoZfy59JI3lIK6poMlE+E
mgjzND0MBF0tk3GUTAzD6reDDXvJHdsFNGP1pkcD6jNqgtO/9YR27mhK5yhnG/lIB2xaI+tBgG7J
jvWHzNtI4lJWDHYWtC4PzwgmPKftQwtb7kt84IVTPs73NLZnUZv0agHOe0FM579IoFQ9sBvuFK+/
TmE3xwwzqbkCu9NCM69I7nNXyQqt+h4Jnkv9m01etIYuxUxdo+4tQyoBgsOgbEyGa0uYLGpm5BAJ
uRnwZJj18ayDLB47/jfiaVLlC9nTH7xw50dM3DUDbcU9wJFdLP5SJswygMkA6rGi/u5mKC2TTyri
Qij5uwR8WyVUIb70yBCYLdDdwLJIcCF20edlFjXHkEB9VoA7s0RtfTHMmNKHdJijUX9oA3rLF2ks
XQJLRr81BNNTPbE6z4R6cgz+X8VCm8GGFiTNQ+Gd7ik2Ky2sUjPRKnJpuW1K8K5yPHVPidKmgZZx
BOCP1OuosTvFPP6gQ6Ov48oSPucQlKR/6vp3nZ0wSGYAd3/1/rsEgCRl0w76upgv2t3IlPu+9uyz
GeA/yQeL7XWeTFo9ll02xJ8+rl6G+NyiGHDaJAK9ItyuAMctWY6szvc4QNe2jKggnVjYoVC5tKN4
Y1ITnZfBN/zCkRHfnUp9q3qNCGEJo+yXgthfgQT+wm+fhQ4C1eZXotka2v/A1ZvA5bLUbnJbjGcJ
+ENJOBjxdVkDgrjfnlHZFjDC8Z4qOQ9lth5dTqFvSnwlZCTmVCtcRbObmKuhCZpUZafG3lny7jwb
4f5aN3LR9EGmSx1Ka/JfPxAHEABzqu/I+R2wgle/dnjC6URzhb21p842s/r+sA/HR6L1tJAPOV8L
MeXqrBO2U40Nl1l5gQKXTm6NbeJYVmUMIUf/5bmOTa1M0bEAq+Dbza4jdaaOtTC7nk2N+0dtCBz5
YS6S4cgXwu8NdJjbeq5MR7qhYdBpIIvToDnH58KJzKHDpwKkn9aeQi7bg8PP/sg2vJPixNWOsVqT
OzwDQbTJD9jKzowvWwUXBtBi65cGbDRmFhkjSi2XXO2cp6crPQ9F/3M+bF6c+Smdyue+dgq/hhLK
GjbeNvOxYICoFhqzcBJv5Stwxg5bb5oGsvE/+BMxohuCkNqy0rGDEA5tUSfJ+FyWxSGUvHxOoN6g
yyBCL1e3D/dNZL9NWvy3HQs8RVBQDpvh4BwpBUaDerW86EXYN7Dd8/NebKUeIma3nfrdzuFZwWF4
fMePSAkD+1kZOZB+br1IeObAFYZZ3eY1kX1bgcM+g42Q3LYGSEYuh5uS19qk/ScoDi/zaLcT9kx6
xgYfL026lTmlkjEGJY1cLfSAxgTb/1KiEtPLNK26yNglcLBSODtJWVxTYE9TzJnY+5M7naGzpp0u
CGB0WVAKe2mqKSKqgytFEM/O3jnQ6nxNXqDV1Us/BvNbOpZ971xtXasPsXQjD1p9MjFMovelHMU/
wAxBu/VncjoUSZluAAK2prJuTlLEXDEbChW8ccRLyTiXmIndSUjrlo1xZKGITwy6JyHlNgN1nvdW
Bgn9eRGp2lJzf0IMfGiPjuIaAYQETCgyC2yTa3d+RoeSoSXK6l6tFITHZRUYUg5ETMmNDm/D8jMo
YQc5YCOu2YUOqmzO8o1GvodG/xvCPqnh0LGs496vBmXcfv78R4OLNXtD/YgedP6lRTKDZeXNoa4v
fgRtCiAx1UpNkHYpyvZ1ND7H+W1h6vzb5fsF4ojW+YaD7f0tFyTFI1KCjpCDsEtMktTbeG1I8VEK
mTu1LWZSAFlwgzHP2bYw23JWd7KCPPvN419/ec956gHXpS2SZhpNKsFPJBww9bSCiwMf1FrE0Jje
OhSiGo/g91yGL8FOL9XkX7n/nXY3jXpzUygzKF1Srhzbn4WHTCcSnwINXCDV43e0E0KC7CfwARP+
kS7DdNwllbx5SvAuz5tYuPQAnkUcr7wsgJuwpkkif9VRpYKpKaj62hiSQauzFIKdnb8tup9V6vXl
AFtXFBCYVlHeDTE3ODL3NFCtvLUYmvRVFDNcYPe7EuX9efMVnK5mdyEERf2X0vxgyKP37pee/inA
bzNAGOzhLvqI0+D4FwqketR1Tl1bE4iUuWudq/sf7a5xc8ambrqLdN6AlCGa3PyBahk3AVL0g9lj
GxCGVQOZT07cZtIZsaVrc/QoTmt5w5oYJQrE4yoJO4mN3IMabehSs/uIb7yNLHwPw+NXZts+2pkA
v0kYEkKIAOkw0rSXQlxg96IrP+PTLS/CcXso5Mt+BVnBR+Z/xr40I1P8bMv3C3g/xCy7MACjwGFM
RK4PN1U1Fa+6O2ZwnxzTinMGq+oE1d+8M8I1NW0oiMh6oiJ+M783+17IjvffXJjivo61rVOGq5l0
5gj/2L5arcHxU3XLdd/68KhaNBn1Ea4q00JyAUeujCqcMLwXTxIFpmrJiGiKkGzYMlBhgjAckSFe
3Qw0SuwoCLX4jyFp1PijvXEO1vQxA2/j4dysJN0cBKSES3x852uHJnBLLR2OoAh9vIDJCIkvyQRn
Y1bI7sARSrgZsp+2l4LxXAlWYo1LDoKEECOKJO5AeZAElw8MtBWcrBKmN6UNs6Fmx+IEhLQa5OAv
/i9s6nGOtzjKks23nt2QdLGvPcs8gUYr6NYfqn1f6HptFx1ZNGoQOqwPeQgI3QfrA3G+TlNAfJ9x
CFxh0AB10hUuO8edhypFYiryZkSDNLFq631ENWodq8q9y2BoM4CMUzKVp0d+F3pWSbNOJTymRgqS
y2slIF2SoFPylPO6DntXcdKksrKnkPv18pNLEZqkV60kcp1/A/yxQ25KzCKyWIWRuZ7cYsxuoEJZ
hV8JrocUgljNgYP7Q4uwt6NeGKBEWoCBbavkolMuKt+wv7oCJqx79E7LKGQxzPulBiqHJqDSlq7b
yxnWrWYFK1Pt+9eFblmudZ8m2+xNqoPy6duBNZIrJzdNF8gHLpqt3byEGWQQQNOMUm96xN66Ksti
t30GWr8A4g3sPFDEZwevcjjdH2Rhof7K5WlV95ZGG2YwRxHLWdcFN++BVM2nP7SG6aj0+6VxIF9m
sDRnZD70wJQEMrZkeZdmWpuyIY+6Dh1PlBWd3Chww8xFpx7IeHIvkiTHQX539mA6y1ydVu3xjeGE
bKdlNSggcuLi7r35i5fLeNngkQL+7JLNJaX/Z9SNbUjUq3Bozmh5GMi5jMCPZZSZ9CP7dt4zj6By
NpC/UsTSdROCOMJhz+8TJemqLThqa5fu81CIam1b/wAQc3dfxhj90Xik4C1A8GXJ13f7THPYYEIi
FSu2ckVP4XaYT/dvs58IFcR1LQ1HLeoMGid+PNJy4mrk8NsPsxMv6RY0FyxY6CF67eCSXvJDCZAZ
TWystL9Vldt+wdUbdDj4WOVr2d38M9yDHj4ucxuSsfeaQKbBCVkkcwWfa3vsnhlpsKNTk1KDuNwR
p6wPXBIJSKG51vXdu64A+7IiEd509dEMG1u00xlpXlSevnVMW+mQQDOzOJ59ZHFDhu/khvWStGo8
Qp5UFuXs+nHs0PV5qO+71E08jtpUgdbL+2/jev4eWylf2/BtffgYGbJak0oliHSautI8hsG1BJU/
64cKdCS0bDEYebdE/Rl7SEtdZpHq3ykeU6n336t7lz5rt5D3C3Tf9pkQvrXqtv2leHh2wmlQD1L4
jPKLx63iYg44FCPknzRy6oKB7VrRfDRbJnEAi6MDdsi3Czgu9W5wNrsTJ6Gjl8gPxKlGbfGJdKzM
MakgeQCLywzwUzTXrrVCcO29v68vZq4TrcVIuG6c85k+njXgj9yjQ3KhZ0COHtuUfs2ogyC1Nf40
JhtP3U85tifu0QF+IJE6U2BKi4QQmKos34vKGd5ODV+yQcqlY31Ojk0sAzpEPMUpz/3XYgkcVNbg
gR3QfSFN3nwfsSMDqH5ANJ6fMAVunHPT5S2AemO9IoMb7RJKhHUMIC8viKnrD9cyS6xrNw1owhTd
WFelNT2fwfpPzUzCO6xnjYa8V02wV0qqtUm0diTE5suKKsoEUFCVYVXPnjOE4QPGWAQ23n/ozkn7
X7Cf95S3CDbGG5uQfQZLjGCdx7AUVHlwy5wKRPv/An4vadcfLS9BLrSDLw6agu1N8bYcCshgHvt0
0J2SDruG1Qbq2kDqxJFb8aadIzS9OtXqtedL8hIL8x9iGgwYSm2pNfAxZDbnTvv+wqe5qxnB3dX7
DjygVcFvY1RJOb8PDO0Xd4SANbcbbh7Qswz8JhnOV5BRVdHDFp71yJR0Rjt0iAbaj1VVuuPvRGC1
xLf351ybtwNMN91PDv1gBJTKNo04mmQqJyDOFCZCeLdkS19wR7XHgo4Yu6WesvIbfFs7eGK/tEFq
VFr0A8cB+kiLaUshsoKB1YD8i8/xgS27WA5bIxTnhijNBHydF+VIceIASiD5bWS7UjQajUuXi7lF
Xg/YkG8Fen/AKnaJt4Luwysw5T15GI5BJo64ZjbgS1M1i1vMrPpLECB1JKoK33EjZ9bXAP5FK2QG
6dZ2DvR4Kv6Cm4X/qVNs2w/tTag+GDZf09Mqn50S0lYwQ3QYMksDSrN+9RdJ2QGl82Z6+Tv69MFF
0zcAvWqEjlLEiAscsHf9pHn0bmMyiHu/B/LN70pXNPBH/19FG8bj17uUU0gPgmiINItrZy3Qq0HI
wSj/qIjqjouiAhucCRjGMRDdzppCeZu7a8WGS/10LCxiVKk4vU6kcZcTT8lLJsoVFkaERePC8wYr
KYt0wb7esWIDQxxGksovpAXRDLQqdpVlU1fmKFI52Jj4yX3WuUNquVBpxDvN1yqZAJyaF2ZR8+gM
A2//KCMAtBaKd8wPLWtUkXYpuNduthRngjj0/InZZaqpyZh7J05pweDtoXlQG8wNtsYDO5MsAAOl
AwPrfIH+8Wz6L8XnpSYnMTQF25AfXcbp2ukKkagZcoAWyBGzCKggZT0FV3QwwwMh36wlj512Styd
kB4t7kY95kFbMoqVY5MaqsEERLD1G70rCICYFZ0gyApjSpKX8Fgjc5FAzq0tJA9dEEOfkT6+8XvJ
amMRXjtNhlv+B1MWzp8+GDwLwvNLuvDgdfDB4Ei+5jQdtUa3nmeWEDFxMM7kYtu92aa1AX+cM9wb
GrNcAOjkJ3RZABaQ6F6DKofJl2tjdZcVqJeBeennzgK3ubxILRPMb+0InGb0LvjwQO66Xk835M/Q
Hr9YkdAp+yzlULGvCTYskApXk5DAIZok+vlvRKC14Fo4iwWPGk8hzFuW7oH38IGMJdMBvz0b9f5p
SaUYhKTbhIcOeGkwfzIuC9PuGIIPoqfjpLD9V11AoLbFfiAYxmEsGmaRhGPbo5eydbwh3rNDmKn/
EhtOgmC1ZWtJwdkNa93xsWWIAXqlJfnKV8OsQIecmJt4L9l0S8plJeg666tYtduejNEnyzhkx2m0
T5tzu13w4E/7FFLXBdMUsEXIfPc36CaJ1mk0rhtE6CL1/To3HdLgwHPkEHCeI0a+EnbKZC8yx0Vw
KSROLRhSYXwh97MnJBneXmQ+XViZnEYMb9BBNUKIpwdt8r7yaw/XEHy7aIXcwAIM5ifrhRC+KuLt
j/sWm86hKY5rbE6EQlbeN+F5wi/RD6CE86dqyFPS+mHGM+Fjydp0Z9Aah7GwnYjEngEj75xTJ9/W
rdzHQJfCkVol2MO9xF5uOBBoYEol1I3bvEuPY9HTTC2xpgfoL15ZgP6EKYizU2W4wE4YyMUtwT8z
4xO3epWdc8HUvjbla9Rr4OQSLoIdo9dfGwdjkm5eFk0KKydwU2KK3780rxjpcDyyNsRIzVMxKpml
w4LHkJnLe/y0DBUHdHF+ffwnZwpZIdtMOJlT1XhbqAbCWjqgMG2dca/TLXJxxpvfJIjzO9RS3w97
F50nAPzKgv2N/9+vF2K4NDU+ou21J0/UHRqoD38a3rtdwMEFLQEtGLgi4uuOXhVAK2yo84AMc+HU
gRZZUXTmV3d7lrXn1qdLOv5ibwWMCLhfpKCwnzOEhxHqKzZZx2dVBbVXp9grq7BbIpDWCYyFGaW+
DdQkaQxW3ANYicGpAJ2B3BIIxDluRcIKrbrNVWSOQVKiAubfmcE5sskqsmTXWYQGVI8NTU2+hD3y
ozhmb1iUdhSw5CrvWiALpZGY0szTY0YRdKDOPzYp/4sC0989SFVYT40xgmrExxM1IJhsUUlyN9VQ
jPML4HPn92oZEN274BPBv5BwijCR0kNGIG3xgMA2FqU7jo7bQc8JgvrJTqhSix4pnCN3OwkcVNWI
YoIMaYmu/w7sR+OEdA/zyxDYlaQSOuqukzOLdGaCoDQ8N01mVpezSxyduAa4rRohHoH4uAYyMHMs
qdInHupF7mDrQP01yL9BGEJkyMXw5IxHFYCpZmH82cMURSE6JKGAD3JAiCqXlNn6UolodkWDzLbX
rr1kg7dJcHnzF6ewKzdIAAPv3L+6ai/WrzpfO3hvB1jV+UP7WMO0ngfyLFusGrsMxZt9lpdTVmtu
qHPZOpW/Yja6F7F+4kkMk2S7H089VYdggM0ln5d0x3YAzHfNWwN7lUflcZ3i9nAT1AGdWAThtwtu
GqtSpMTIUGiQo7y8Y+RC+mScocEMEw/prKbbMnp9G45nxgHZs8Hv9GpRQ+L07K5/LadVZU1xKe61
zCUivSu3+1/PJ7lsdtV/ugSgC74BlkS05AcGOUzXESYSdtob2/jW4C2co5+cWfTjldIhjSJrZ2hu
Ooo+plVIKAHfBLfL98ZL6z78qhcw0gXp7TRqQvCb8kBUvk/HSj1+8WmqVU4HbRMKqHAXf3u/cJC8
3TYx1uQ8q2KVs9OgoyvPy5fhdKQ0XtYn1dHDqe/An5e/1H7Ob6NBwFO9KDMGtZN/PFOUZdzq39vP
lvZgt1gFEdeIZOc9ZizLt5powsuKFna+Q6R/rlACdL/068WwI15eIv5Uy4ZaAvw9xSSfEWnOBio2
lU4Ahc9iwtg1ivHV6g7QBKdnKxPzh6zw+lBzcz7nEvNYh2Io8nRTgmzcLXJq9FkFYqHpkaW9NQsn
Q0fJMGmjQnFYqaJV/ruD8jj0RpzNWL6wLz1buh5HMbuUrhnqGqxDOe9dOE764i5m9lgT3rc0oBZP
KVcCFzUeKtx0piebSIWJGfASpuR4yLeEtnpNn/e5Z4En5ltqRS2sHZzZxmmE5uQvIE1yxaHXYCLY
1e/cPeCIMskq2/pk9rm2dQ8klIrbJp+gmN8tDap2vl9F4HXWYmhJ74fG5fZZK4cMe8vtYdPiPmsB
yXj7DkxOPMXpyqqm9mD3/yuZ19AoWagGg/UMoAPpiZyQDOg+H6n3NKL+fg657IMrQG6F0eTE9VBs
klRu+MbdlB06uF5+/LiVdWsyQ6SO6uBZZJ/fp9VJC6NHVFW0u35Rg7IcchWTKFu8RMz6FabxnXEa
B8HYyh9fBnb6Pchyxp69YKVJ+PGd0dZDK0LNbe05SDHDuj2MYG5e6RoJSTJRit1djoJI1tSsGPvp
FQOQSzO9GRii86sfCMXdR7lApuhdAPV45BfQa+8cR3ClbfocdcbMHEfb8BlslGIAMsQDjoKXxP7Z
u755Ro6GMLRJ0eC42YWVHm8AhhyDXtzwRaFffflDqB4nI5YooU/bQJC1RnEAirufKI8/kkToFCdI
IN1AEerFwqK+upTC+S8C4MSWRwMaknyi4TYgxNcipoY/hyUxlaqvr8ghFhbETG7y6Y+st9IQfEp0
JXqGCppYl7eppnvONDXPXfR81uUiTQqrbrHO/72RN5TYM4Gi3nO5fme+xpXgcM/8u6dsIM1748lZ
ZFjh4wiLrGDnZ9vqenZzfRAHNtjFJ5RRd5FsfBnC2wC/Va/7UwdI7RtmpdgMXMNkK2iaM+YD+Jef
H21sQPCNOSCh4am5uTZK+lorIDWkG7YUZWvXHVSmuljjE3eNhvlIKsGDfrnEKilORNeu4YYEBgPl
c8yeTlPVRS4dNzbfYEBmLLKFXO7pfJs7np747Ge6rFMsatiO/xPN/ZIIT6Rn+IH/RF8HRVCyrnKs
mo44vJATp/XwdAawiL8zwbILUi2Spe0QrO+y+pDlNBLaZ+IHTAZSxJ2/qBRo6EuMwFEz8srQ0ZPq
lcrqNA3p9f2og5ygvzHnDr51weISnlJA6xzg74Ds9Z5YivkBZDDETJripSFHLXROtwwaVvAwnt+s
wzwmp7ldm79qijxR3yhTj16W31r3e0CE/R3Xn+g86g7fyNm1b8H8gwLtg4N0AvqCkZiKg3aSeyjA
IQPPBz/fCij9Q+1SoNXAX76AwMRAt2WReljcvDXSyVgblKRWwzoP2y6G2twnNAEiA9rd7sI86x3g
ta0YOHNX0mA2Vw8xJcgXYbiK1vcH1kb3GBPi6HNMjWQ+AHiSAYtbn99mbSPQEqzpJKRvTrUitaaf
ExfQnjdfPS2etG+XvUsntmJVLHzRlFJH9rf+zMIQXIvdAbOAL4wkoA7w2/mUV800/TaXS2V+r4ZA
3/GUQM6ac7B5jcNU3KTXxfUrdrgelEZ4fnI5pwJE6bt7jIjYPK7TTSplcHXje4A+miZ9B2BlUndG
0Tk0kn7D1sGeCcRf3gFoUzI14i/TuPu/7+KXW3UhZzoEgG/PTl8mu+Y9HvyjYigfcE/BZaopGWtL
lo6DX/RSFfp+2cbmcNo+rxcx00beaBXd4+Wvnx0QbdTDGIPcg5knVvZZ+oxbgRp9wvvzCgQgYdH1
GiDJIJcpjZ97+XvdesVwFoRdzquqazG9q9HvR/FnJy3LL5eTZQ6kegDTXv1fMWG+saQbOVP9FFZ0
yu6kNG+Fu8sE1MmxRAJKh83YaHDKOMsAOkkqhRn0n2kQkB0IgQXhzBA+obl8ximSXvLxhVHPkYkg
cwQYp9zeCAwBZZuYAL16eh2bwf05kqGRc51tp2bg0MMSl1GFrJ+g++FHChjKZJqoFHr8eOUtuAuH
brhYsyRC9fN4kL+oNjAOR7AoY33sgMEHt49AmCYD/3GE9BAMrEz1o838taNTyx0fMKEy9e+a/lF7
dpaIi86q2t85HEjRfGSbeNBpEQeT70RnkNoUVfwFIVXOtVUTaFiUVQU1on2TwwgFO1YvNcj5v4Vo
azuLM+sCRaCkI4o78+thd7kfmL8/sfrXIMGakJcdy8TefwG1RhD5fl1PDODPurIRva7oBC1v2Grb
XsdZbJsVNEZnP4WbCAq8YpkJcN464AXdTDU2Pslut3SyzY27k8rE3y8cRL6/zwvxl6BqjYGyJxwG
EcPSZIs4LtPc+G2hDEUAru2MIq3W6HED/aucLwWl0yb39EMl/DUVFI89zC+6gfTv+UbVKuKufKRR
LPw37//dxEeVz3/kaqhI9qE0owegUIqmDOeiqLBUYDYyfcY4Gs2B6DTawxQfa0qF4Loc9igoFWQn
slI2Mg4/2KffSeor6b8FOCp/dFuMqwDAAOyIjYl5Z/CIkQdgiTvu3DuFZFI2FLPUxiG5Y7OgDqqw
qbMlRpn6s+S4wfa2qMKu2cx7ZKB03TQOQMFxM+LNi8aTFqwmgEDoddgvKQ7cerzRySquc8+udYRs
ACQnECatcTXAkY1J6LEHl1ngaoxNzizAdurgtUt3CBgbOkL3LDbofXL3gx7+9zbipezBJQ17tPi7
P8w5A2shdVcIIb7Cy9PW+NSnLXADlwJjWGRmgKk3HC9KowTnHSJMjHCeOLt+xHu56tiWguOpo9oN
yfQqvftxsRMjKH9qc2j1Btd8dDvN5RbMR1OhqwnQ2G0RZ6RU3HxXfHUB2zZtIbY/Dwxt/szdtgWK
hUW8PNzW27kQyMpO1tvvkSLIJAQmWGq86koX+bFAluUu2lJ994ybOl3rq2IGFmH6BI68sgWOT/r7
EfdALsduxYBlnAN+Dnm+O/3vfZgZMVKMXO76wrH8sTZSxcJXyiOhNViTGDwqxZ9PLQJJHqpv249d
/jMggGvPAwxQIFloO+Gg1Jh46O3teY2/YGAX6rqRsXtScVJ7dfzZPAOOyjxN1wCjW4bN8zJMl+FN
oR//JjwHB/Zx0Z0pImMt88dUJ8O61OsFEs9AvG8x8rVVKnRU8HVvErB0fXhidGtvjmIDxZoY4Gla
ZBVMhcWCZI/mCb28yve2WrYdOd0UC4Pqoqz1Rsl+fWwA9pJyoXMuiOg6gP6b9vQiYBAqPLzJjxWy
rSKO9vYnQFzQehkQpeQwtVOWXmwvoDL0EGPfplyShFfGQyPHzyn5keLP4AJPEyrc3i8tSTKopz/V
/eiHBiGgGtgJu/fHdn5d9rxqAP4daT05WOs/X+w4TmIvPF0RWBQJNNfyp0vYnfS7romylKo7wp4t
GJQPIkMBSeDqBE4Rq2Whx9NvWZG44CvuT+haAeLeyhi6LJgZZD5dp+QT18jf5kbldBz+5LqWimBa
HBaij3qOxqi128+7mn3UKqCwBQtowK1CB/OEykDx82mmATOYL1OmU+/xPMdmTAGnimuzOgLKWipU
PrX6oKJwgAY7dI46xjkGgH3n3TsiCbJIKP1c0Fs0DDVTYn83M5eJAbmO/58Om4skLpw/emsXMsuw
Q5QBivJlXHSEW5rZjJLtPYTGQGkUHB7wCYq671cVD3lulJZrvzekjEwXWdmqEbe4HrBJle4PalAr
PjXQIgXlv9wY61kAM8HoWrj1ZlV6ywxFJoF2cDpWTBSiDKaZ2Xip1RWaVPINmAoG8FdR6yzb1Z8J
pkwvIQqAf2u521wVuH0D6cK8gQwEYntfAl8eh7jbTopP9KIh2ieNOvzUfpt7BYVngShSCJo3lzXt
P6mmWn7pKUIA/UOV6u0nM4pTD26G/isCvev+ICC/8rR+CV2OSFVz0BRqlAM21IEzHEhlXjPmf+7c
BlO98L33km0VfYdQT38ebF8idELN3JtRQPR3iwkqLyCvVxiNKzVY+QLb8L0ZS8MaKzsuZIshO1zo
JjZfuNncJm5NC+AYmHm6LAY97cMnQ26/9fsRsdt5sGHDu+2f+rFE/c+XlicH4ne1pyAwRCkOXvv+
bcMkDCzKW/aWJG8XL56UB3RNkoi/FrbdljQlmkjOdt475RAv+4AN+U2GNopBOo7U8epiQb35J9Ey
LwAVJqy+F/ETuKo5rMq58pwqKvHzBD/oiKmUPl0xW3Uk8MEXLmDMKMdH9u3SAk1PqMZhOAs6ipWY
uGLcc5dFYO1KpZ85BZ4IX5HCN+GCbUIeTryRPlyd505yoSicxms74F8NNJ0S4G+Xt/H5os5ECafo
wdzB1V1wGlvDAu9dwJN6liGgJXPsNKaKVYizr5ku94aPYx4xUPE1W9eTJRGjMXb08x+msebEMwwC
5YaSf8R0rtYnBIgMYyvNhnf66m7B9PX0QBpI5Inl4pKfJOAVH8Z1XWuSvEbnVqStYRl+ApTJWro6
m0Xt7BwBhiTI1iHaUsJUg5PoxnAnbtCuIvombjzU2WG9IrTda4Pc7DLwOAUQVXHz7avAbFc4ro4C
5pjnZ1kJAiEQspSda+WT92k0nKceqRrpR0WPO+xbRKGZhpH5QLJrdhS+OTurZ0lcITRzLYCoSJ+7
FtT0mE2kT1QjaPgI+VOL4F2QE33Pib4u+avcBTgrOU12qlOD4msBTWBBnTH6f+aWcXndu6Tn41CO
Fio55i3Sgve/Meerz/gizkgQhg33PQqtc7Au51XGmAg5FyoMuKmwOHgn5/Pdo3E2WPKqB5WHn1kY
01qUXMFoJwwGQtL5JVD1hd/0aTs8Ae1nbCGZoWN1BJmcBFIqeBIfhSXC0B5FH9NfzisjyOFNvTsR
dLie0o6NQIoE/UfT9Blxinte4w1ilNm7x8V39c4ncFJ3xrbChExlzx1WP6z81anSnPKRxck3dIv0
awEjvzOaRy7+glY2FX64Yqdfeiiid4grfySzsmLC3mqK6/nAH8qrAzza4LYtwVnaxrMKeRGajRj0
Na+yDfQ0mZ7ElH1fy9uuEhLNa/uMzDi/NFXlcPqig6eBgEmOLunfSvKiIbc0Qul3XnCP+9YFC7W/
yor8P1HGt7EO+trmh4lXpP3nMgbgi3RxxvGFwXVjXcs5UvQpOmHqt70Gmy2zcA69Fmtl6cwXk/J7
pp0Y2CAK2sjpbFQ1Y0JfhVUojiEpLdlpsDZIfp0KwlNwanWs3rPr7HeirWjTAv/EB+oRcnvuy5WH
fgrljV//InWsDjpr9vAPG5819CDc4fr0dyTriTtVoE94TKO8oYhamlsrBiTTlCGl3aaR+2ZzFO/m
cnrujOb/6aK6c3d7/N4eJk6qYLJO0sgWDNTumw016HFThqfwZQ94NTGQ0op9+n14s50wWHBU9AB8
XO0ggAmnKQbEVcIScPelU01m/KB8g6L+Kho9pKy61/2ANGH4f44xyqjP0OOAzWcoTedaZXrOBMpn
zGF0n5KAXnEi3GsqlMse4UF844XHwmZMnqCYP4kMlhD9vccSpf2t5eal2elKgs2L+bMfUbAPjI99
uY2iJJ3rd2S6St2Uwu2U3Rcmi4PT3QnoZC1RvAUA/uA9wOd2gvL+yhMpew/Lh0BZ+HOQXDAOpnFm
bkVX5b4fVRiVt8Lxnjql/zCVyK51dA2B4v66rRoYQd/5OFemZtWEoHbkWR99gz+7aFNUgz7jl+ci
hdK/VMT+BAnqcM1DN3EyimoWw5TKLnvvm1boY0g4soIjP3LhngsriwOsuRhujoIUkN4QKV857bSa
38u3uAbNYmOHV6uLIDnAPtK1ECFTJFPn+FEFhGyFY9ynfOrackcfmJ5eShBRABo6x3cyq/N8I9Bm
UCQnX9iRM5+/5znCWSW+XJ8oX27m5oR6FGZfpQxmPNa0SAtHjnwa/sSPHNnCD/B19vHKyZl+pl8t
J38+4ikYzIXFn7TUPPDtm+SDzJvXdEFX5TRk1tDbUXbyOzMUoOTqphJL2JtkPGMRPvp+gLAwKcFz
DS37oqNikRXRF1cPqV++3M+CzriQVieiaqI1MM7A2Dxv5LWihYHUbgkBm0dOsajMgtsWpEJvjy/L
VEsbHPDD1RSotvJhJjFMUukAkcVwgMffOCsX388Wo/Wxt5RrC9Ws4uy2U9XUeBplodr5jNOBNk0Z
rfPfqN/u1HSlGnKQOGHTrvmTvGtR8dHbFctAwNMMephDUNlaIr8ImEh9Zz1Hvex/oEcd/5AhUqxT
etk5ewLBVnnGLjK9goOq7NbobSnDTCqxYGMkYeCQKDM+rMEYDswKhG6NOn8fDVpGmqfTFjolEiT3
MCrJ8KM+uP1s739qoI7jA1SNX7ZoknWo60GT4Pwga3yM7vMzT5Q55yipIIbkjjEUUxGrz25BReI2
RDlotKf1lVi2jwIdocX3ud1idrx7NQq6hLruc60dNriYedSuFSPtpCXN7u7FJhxtDEiEXPx6I74G
YpdR8Er68kGx4ChJgwhXDLwW+epgiF2j3R6QEUd5b8YAOLGWfYV4+V522Sii0DViplueKy/AmALY
Cz7QfctWqhyC7tmVyviUv/by8Aw1qIJOCJjVeKEww/dPHyayBqauY7akxdyQ5wLStnwLCLSnUoyQ
NM7fnk/jmFkAjH8vWI51DvC3As5/P2nZGuSGRVgzvr2plnihvTMexKpt9EgQCdJY1x/G1PMO1lzr
tyr/dvKpom+EnnYDGTfyiyzGnfORDULRQp35CFzttrirKS3Z4WbUj9kmweJzefLD56aZbyqWwLmt
Yyky673b7NX3dlF238cxgxCOdxNaee0g4jYgbMxnw7DsYhdDnCBzmOh1xfHc9k8LbRwKcWhQgKnR
gROOJOxpHLQminEVEoZWq9Dhqucg3E5F3T/BqmmrEnkJVVr3G6uSbjGRfKbGxuhFs+1u3CoONRH5
44GYyHnj4USxRQpFI8BDyAfxqRsIIeMzWE4KSZgJu64BcyK0e30HgNmNZ1C6Bb9UVjXKdRDrD+y9
QWFvxG13tX6zO5x5Svdm1Jeq78CdeXHMfYWU35ErtRQKWdW//wQtUKuBDdyNyW8sEg4UCP/ZCjwu
nuHCEE488PPIY4amID0Yfv6SNFzdcGJ26p1XK3gTyqCPb+ljiqgpdZ7Qw/LTG496DYCFrC+hQ4kd
S6NwhsO8Lg8TjNFWJd7WziX4l7MkVJsRB8oyorQCWQVnDYDPfTpNe+yUO2mByudiM1DaUEaH0kBV
OL67pI/mtXTY17B3cpxrKEoN0a8wa1hPGSoVhMYhhYzU5ZxOpfRgaWUqqmM6thwVy4ji3sWOLFar
eBR/6fyh4OPjibB8AmtE4IMFOwl41hPewX6TJc1xk1QU6MXFy5aiJcKmZn9prO2DLMmSEI5gSJCB
SyerlFNAhJiFbR1G2/NH/hhVvwKMYQNs8f73xU9GdjBCmqF6YKBnyf2o5wX4XowXDaRIDcdFS96o
7S0uouPaCTK43Jcdy6K9L5Q9SMz+bi7dDv9nadJx8Q0dMcOuV/dhlwOT1WrLFNv4xqUb067lUQfm
AjaIXmZP3+M+A9gFuWT516Kiky7lXj2onLZviAuzSJL9yXbVpQKu3uYx149zy7Be/uTX6/3+/pTf
GIVYXCbSDyFOjrOf4ajiNbcVtF20V5SN2vZX+6+BABXWa2NyJmNr73vW0N9LdH9AvWS5BlBe/rnf
PgS49XvvHfWHZBwjgVrYvHXnul57w3nJ4fHCnVLDmHn1kC+eHRNfMaKJQyqw2r8ZOU0yEfP2XJ+S
wAeND1gaW04KTQfEKG31EHvB3o4pthQmMITLNJuKV6DFJG0JYNDe+bPUu1grZ/542Hmhh6MnyGFL
U9yF9RJmayD8WFYFdeDo7LhMIEz2KHv7PSoCk7iqzOyMktjpVV3raKnLi4C3CKaRJxAVHBXuV343
grOL7VGG7n4XhkR8Q9YUqzf5LOlhyV4sEIQvf0iRQ3Ripyu7591acCH+RtSd5NXPI95V0KncPu3i
c4MxZ4CDekJhKPMeLaxFJ2YYdVPun0KNWbXvCpNXeo7T71IPyqoj68bAj+sm9RrVjscjQ4rAbdz7
IMcgtq76AWT0t6FQJUyJWU8CquoOT9ehP7pXPpb6CPwTnA3WKoxRmk7ocBTe6ZcTNsmcjNMHtaGw
QofsSzRQcAT1LRVddFza135ly1uiUmwU7yfd7Nz3/u/mDN9NkeOteK4YxcXl5V8Ui8HRMdSc2GLP
Yb2S7Uaf3opMvSj46j1OwqihRtKUs3T0zgN91zVlZcAZYe3sKrp9NrZNCs5hoOLDY7/RcrPxtFTm
PCzpWnZZ64JwSeASimKRFGAJZ6phTEK06QBST2I+A5ttOpVKU/dZ9p5o6uL0E8UlhuXaCmyhT8Mt
gNDIYzgX/IGE3px49bXcMLM7jcVPf7mGdbYe3cp2+VGVWjdJeXszeRcqlY16rjK9mHMY2mULoyeU
UWKQya5RsHL3EMqyFoydOf4Yg7eyoga4kPWLGf6UWumzoWN/flpiNyEXetkXN7lFNrzKLh6fXdqt
q0yIEPsuX9wriQkImngFZ7Bs1coGeU7lm78cZW526Rn7QJDNMOGhFxrnn+Jfhnn/o4To3j6cRwjM
Mk8cBT1MVHEZRrtBARR8ERlVmjsd6079LvrpWtZnjqyIPyXZAuilNRb7DA4Ddv9x6MJrcBEBKr20
yz9QdWjpx8gvQGEFHLiHf3Z6gnMgkCMjAVxWffVY+M1FD1/51XHCevsgcfnJRZ4YOM031s3Q4Bwb
nN3xQ7qX8ut1IzJfabLbLqkUGF0Eq4rLUVFCMLlYJDvAiTsCupg9FfRYPc40cTK+DJmFJRfTcsEf
uUfoTtbzNofV3CL1Zm34Lb0H7ev6+suEwtuJPhsDT1hUi9zPhJmOohqoE6D41CfQTiKia6q/R8bH
8QY8Ok0qnfrSWH6P1NDs/1yFRx0NjqMdGPbzn2etXG6DT87hzlqYMglEP7uLIBJjlAvc3U9OyEfy
eZKUBzioyMgDhgSGtK/cCfhOCYfeXvUR0uYl+u0SIGqCCdNTsxOxuurDaVwfdQdOecSuIHXxgUOB
B95LFhysiuEG6xd1MxLgKCUuBaTugsSlmnjp7W0+F871Shyta6Vbf1lc4+DPXwchEkOAGBzil92N
CmNAEjccRSZPOR7SFnKbAj8gnMKvGKci1VltRfAD2ijbWBGbj5fMODsCXqIwlHu3A4KYz1PAx57H
wBsnUengeKR0EizNHCYbaKiVXWXL4BZf2pnlBObcmTl60A4fmyIGowbqtZa2rlUlDn5hxD5EgybT
4x6mooLICJuCOszmZ/94Q0QO65Tu8na/QeCL+X9NM2fkWROTRQjxHYyq65tDGF8hv5VzCtfQ/+Hj
zwAHdxwJ7fvkwaZyGwuHfVFyyJVOedqEcojyO3+cK55A/aFVJ2mEnNGUpvZCIiTKi6i5WeuiGkYr
B1qSprbA6GcKe2BRGpmk/2hHL3CW4VP5aBdYmCdXi7Dp3sUkFtBLpTRGYHWv4X24ZFAHP9YmS5Kd
vLQKhJKtMGbJFxc4VgOnH8AX5Woqe0SxSIIv0DG71zkyC+S2GqXqoM7EqD2/lYDI3lDCGQDfu07O
vEk++dGw8fG6j8SbGeQrjgq4DfFJIhz8Fgj90b3AIDP/A4B7TmOkrcK0j4RW+mq0vzrEq0sMIAA0
1QBb+UxAvJb4xPMJQUzh09F4w2lZsiK+jZnUQxteDzBqEcLF9cFxpzEmrE3LF7ahFoa9tPEXLpeN
gw7Wv1MvPhsTB8iFZlX4qp+RRsmWxi/7ezXlNS9pt4to/TSCmJ9+H6i1lfvuNg5Fukr/Os4YrPHT
UNVdSpuL12NqMYp5D+sK8oFCwmS3TEb4EWr4eQs3QBJZVts4aBjcXQhWq8v/A1XwJ4SakIkc3sFk
ge3nEGRpZT3dx0lvUGufYUzH/Q1+sDoSS+fQIVuSQhVTGSfyRHGPsREpLYmsCUDRBlN4Ur+jvVj4
7BD+hYfTr3xvWNC9hSPO0HlejLVgCf9nQsqUwxyUchxAPIWcfSACT0zHI5Q3JSvUG9bglHQBCim8
ZjqPqUb14TEbqgSaVj8Lvy5u3dwgJKfRm79kTBzvkmD2XM5+2sKxjt3yy5nQez9XDQLoN4Q3KL+O
C2GYfNtn2GgonBQk+KRERiq5qv9B1EhvE3DECqRIAAcfYJ1de5A+l3q+kCvtU52azNoeieiLrlBI
yMppB+iFBUPoQm8ZO7sXI6M2pHFHNmbEI2h9PAjdbIxrUQ3fRhfbFVhEzznZMNPTJ+Z1v+tO3LNh
aglQQw/G58v6oBrLOKBK2ujqy9R6VOqa35N0z0W3aDVND4m0CN3DUBYX9mTZL0AvyhOdtClyGlzY
cNJyurBAnNQFqU8TLRSa8YcAnbTrgWTfJcl0un133MR2JcIVoPMuQwbQ0rsvExh7dY6tiD19l1UF
rNHefgZLGK6hD/7RxfbliTcDMhYT4WM5AIBrzMQmGV99/C+phSao+VijjVgPlPJWFDERHbUxtjys
foDmNRek6yeWfqNWgOYXHj4FLPVYCfoJpWi+rigKIv0UrDiDhvo+RyVDR0ZP9paxfsjzApgzhT6T
dc2y6vmLVyjBLAioXVLZDZF9Pgv+psyq63wA3aQqXD4KQBBeNzKOd7eOubS5XgRZab3GJufVYDng
qfF3tc42gyBmnPWSBEMviu38wpv9nOn1SF1t1G0YKv1Vej9vj8QiY4PbrWGIEWYvupj37wAsKsb2
4xgK7imY6a2Twu63G2trl7wBZGZyqGTfMvw/o+cu1UNxpL0uPZhCXK+5V3qQJ2FGApHW/Q+Gb/lj
WmUKJFcII2xxtqtZ+SvBJRnd26QK0sfymZKmDdRh7+g9xQ08uWGbkShdOhOtYNZhUbINPaK9XRJa
QIRbNieYf43xS/4Wh+sq2B8X7KaqE/zsuaqZF3TFs4xZeSwMe/Qm6TLh5uFgH4SzW/jcnmbcyVvM
TkEBdWiCydzHHKlKakIrvXMYHmVJ+iycOb2P+YXfcHYeq/Z8hzSMF48yz7LdbyiG1rvSF6W3o6na
keXc51oVzu9aptXw8hFZSZhMhDlXJizOjSJSR8eOiHVEObeEcJddIfrMm5sRHfwPCI6ZC18Fim8P
OvNKANdUngRq4Rt/aal579dQh6hqOX/UkTTgZtpD3fs1TfjCcGwHhPlVXSjwZVXvHWJXzXKu61zB
oIpyVrxijYXiFSh1zhi3tD7XJHObeO3IrOV8sP4IFJbTcrPK11l4+vtY4BjGiZTHfaosNAPV62me
EoZobSJVOXmLELzDoHYoo0fGNYYYBbeNnTxEcLJrzuBpFjMJkZkdBvhgvpLs4m5It97hN1Zzs4oH
YPyMNxsW3WdWasD20FZd7Lhwz5cZFHw0EUhjgdf34yaPBijveziOBdfez80gevIqDfGKqGb7eX5g
0fSE3Cz37dK/Xv3QcVVzie2Uhw52bfrwZARxEUiCn11cNv862SqZLsdOfoi5MIsp+g677Kb1FMV6
dMQA5GU+CTEXCkdvgfjHwoEyImXpYDDFH9Bzn+V2cGQJcdf0RySKeI1nvDargYCMuiwM3nfINbbq
CHTfQGK3zEeepGTUnlyJlnSIS01Xh48bLsthd4XypU5aRhKrOI4HL4mfnAn/yza4JniaxjpuLcK0
ZT6gzGqNNkzI1BqgoVFjljdO9r5fT2N0ByxorJ+j2rqq2tLwy097Ovkn/VpFJalPygWlnSjAHAFx
r0vNixWt01ewvOoIP4uW1lUYKx9grxChLDNDPjhEz/7mzAeOJVVZ06BLwUtg7b4iQBGAIdKh5TYq
pd+GqHl+5KEzh3xc71zD7QGvUx19K54vZrm3i+Fda0jcqd91FNNtMkaEVCXIWUXSAxaYZ9BgjQEn
xhmH0SLoPk0WvNrCxSLCVrybLjPJ+BiiQQaM8dYEdS/LLmE3L8/DKMxBcq5ygLxWPRMYU9KEjJLI
wb9JBQh3UKeNg6osTIRSQvmafI0kjZQ/ZCQIzUhsx/C0SwK31N3g8WneCr8BahWHcn7WBWQj1q42
90iT4eCEY38lgmIsOfjArkbRosjE7PkitLyHftOvU22UjLLi7LUwIFEwEnjhWPgiQ9jqa+cYkMr+
DKbqzlr61Alb2arpYaT6fYq1yMX1u+VD8S2ZI8FnSdkHM8i7Eq93YjRtmfcwHrAFw15ns/0QsrLp
MgHyvy6M1RvmWoMXy9n4FdgThkgXY4wenauNOmbv0bPZvS95gIYOoc+CgYsK149cf5Spu8oxtL/d
3pZyO72/F3u0Ej3egtc9Y65GiJAbBm5jAaSDl2d6l8AXiD8kPut4cNTG4TE5uFt+/P8ZWMTV6IOn
3yByHrrV35spUUdMG24YKyKvBEqcIpwjxdBT4YX8oUE2wPTQ2YmO8FtfN+zg3smpOqOiJF+ggsWl
VHApyOzl/8sltR9WlFUbfqNWJKp2nMBHrnY1CrhAyWB9rqCLod7nTHffv1WSwGhxeF4Z5TOqqok0
cuZFi4gd9AiksCBHmJ3uWq43c08Ybhu9c+TmKP33reJceR9Mle27vn6EjqOfPb0sjil+7sYD47E+
2bYKt2vM4+m8XacjtLvDbJj/R6rzY6DPaxhuwEgDXP8MNoA5GRRPsZLG2rAtOq1g/PNr1W/u4obF
Z/NFaUqx3sxQPl1dDKx+i4x0Kx4N/w//W8oOQRGxDSt/Ydn7zeWGU2d4zSyTrjSSNsUfqhErPYmK
t2scsBpvvOG5TRQn457kxBy4F5gyzzwDWZ6VVzGXmzSdU7XkNzTke6iZx2cTQEpb097aEAad70Ch
spxz2isYeqJzwA3zJy5vDSA4UYxoMBbVXrYc5UuOkEDGFKp6HDRW1x2IYMJtl3vniNrklGTzJ5Ol
6OMSsvIDvbNDjPaQh9cTYWXy6pXVrmPwzi49wQ5unMFEJKZ47UekJwTrT1fzmsy8TOilm9RgxTC+
WMaoTL6WdobpFitWDW4T2S2xTPrQ7oGtQOSATN2gRXyOGDd6vq4sZ3VR6E5ngU3M577otPO6Rth5
7WRCwyraV2JzV3v4FGdC2yUkDAuo6hTs3kHHI7KIEhgkHV8uDo+eH+EtqDvQTSvBgfv01s9fCgNE
423HWNbqNQqytcYEXjRSLo+AJYdAIjTaX3gxU/qhXanSNQW/EmX5/+biF2WkgODjqesl96Wj+mk+
4jC9nRNGsRrrlo99nKefXrx39AZqbHZ60Bpa3JIvSYLS1Ispm42xSRKOUkQIbkL06LRoI0iJFDWa
1lzGF4pSq2+ApzX50NpyR5T+c3Givxv1pwuxM55jYMMlbB/653U6QwI+OxtQ5eLK6TcAHf6m98y8
CDyj6O/e/DgShvg5ceB7O8CQFUEFtGsbjxZ6fZRHySWeLjNCc9wNiddrveOOQL78KSKLFFYTKf6m
vubDktQ9TqpXcF3Xxlsj1yvb576BU1cqWKgwft3ByEcCctdzAoiwy8OA4BZA4xgBrsdWsec45K0E
dRTwxsWfr0tKRO7gtJ69dJWy9TMw1Qf1KK2rB1rCP4Z4ojNTAqmuWFUm7aUum+8d72QDz6g0xsOj
iwxO+smqOSbGWFACdjrBgf3xuMim6loUfxWoVY5eX+6SBJSJAYBH3VLbLBbpseIvH61HpJ/4s/tq
xN580G4muM2TjdIH40YKuVca0ciLyVu2uwNua5lHM/MRxPGXKT06QnMI+cMNN5YEsS/zKPRFKYpx
AFKLXwfRHolAqxe9KM8M9oqJ/lHJ/+QDpY0xIQ/vsBjB3mT7v0sIC/n7lHvnwopuU5hSIJCSvuKU
+1y8Es/1DVAhLPFDTvSPPehxycr9UaXr8LGOidmzDW5gB6mSZQ7R2ngCBN+DK0lUVtkaDrkItPze
eUAZPey2/vRG/HlFm2v+VBRY0UUQcuvd9mFriMJvzVh2f3yXiz3e2Yk13j7uFOzNFcRuXcGhQugj
eerWcaeKoW5/Lbe5X5ARQ2LhsCl3LQbcQeuX815TzLqB3Z4wTOD4bHTPhCTVXIiMhMYswz7Es2CG
3veyOY5fQ+PTGzC+dtzYzYwVgFMMPunRCIcFkjIydpvzgsuLa2b5cnyBuY1ad7PRrjrGyCUb8ZCw
SisxzDmh7hW443Moz3bjUfnG9c2AlYCwKn7keFEjy5RJkzNkIU/jl6i6fge1yKMA34+uhQ0K5Bpb
BDVuJwKZIVRHlS+DrH2eiAZWwmncwlKCsEjdGz04NuNz2HBIayULGOK7r3ML+cKXoG4kNlMNGRaD
pHm1m14+FHQVOExcfi4vUGhBmvbzWHbC0CO9YUAoQUB9jlGRAZDalS5QqzCbUh35gw223sxPthbI
UU1i/UU2P9fluEe+nSGCfX+pVt8MPQPj5qlpmn5/YGUhfrmdi/dv7WANm0FRItZvtTgMTyUZCYHY
+BKBECP+DyBgealdAnueGEQGr1ZxQXw4swEaA+H481/uaksrvDUL78xQUB0u7rFD+GY8iEQiYH2F
tOqhYOsFKsSPGMPVTDpo49Ny/KFD9DBpsRZPtHdOH2/XXM4rzTwDBHWvZ+Cnr02BI/XIhU3bD0dC
Sz5JSesefLdovBJzM53fiGqRGu4ejIfpaQMcC0nb3gvOK8X1zz6gZpm4blTNHeDyyZ+Pvzzbu4b5
R/Zkjy79dEdLEcgTSUbC2zmdKtzUp1829UXT8inMSj0Quonuge61Kpi2q4vobJn1+KCYzf1K1xBS
P9OgtMOyzt/heTPpDtMrox7gjYFF4v1I8vMrJIqLGcR3wughT+mibjy7/C1OEpkK2NVUtnXCZUPx
h0zpa2D9nyoJ8wIJ3AW0h8Q/oVQxD/zsMl8yz2XZ0eQR0qKCs8P/CASJTeASIhy86cbfeXNtKyFT
ami5CvrpqJgVIz8O3AaPiqGO45S4F75uTHJIJtr/0O2y81ysW2fCK69cuhhC4QP8bnY3HIruZuWV
UencRV63s6jxOpYyUNqrr+FfK+i2E2fWi+xopOfxlzVx+d0gnsg+tubGR19IDSD9UoE+o75WjL88
Yc7uysqnij6tgHwGpdpCq1Yp+StJg8WrNSTmXhTlJlfTv7MLyk4+DfkNc3rtXW3yuumHmGRPmK4A
x0mCnw/xde0sB2K2SGKJzOj5Ce1ci+BzAGnRJ+DKSQciQIbXLUOtg74wVf0kYgoWeRNcufrbq6Fc
/gBXOXoEgyRpi6nimC2v3MUuJ1e6Kj7RyR5dCl4RYLNFSV+6cgmTkJdX5bX0ns1XOJaqSb/A9DxI
UzWjFrt/M/dYjxIsBlWW2fuqLwEiLPep7VbLH4g4R/qEsjMn6wM3R35YiNeOr7ZEn7fbhUPwhPT3
k45LPGfTygSiEW6ZFFeqSpjmyMKN4ZaB56wXXqR6/WPZmg1+4Tz0SBuZPjVD8HnkdQA0vG2H7BfM
Txje7GBt2LlR8/hxifcxFCXeDQtK31wfn+BBO+r+IIxZPk/ZEkkMUgPc7c87dlXhBQjWhhLkSn/8
eeiVklkytbqWAmLfNnaudpEJ8NADGMBcUA4pCbtB1Tm7dSkth9d2ePR23ujxO96y7JSMoV43O0bh
bi+IvcRyfdsRg0ue0sygyvp+8cUUFhGAxawFB3A8wmqaP5moP0qvrdxazoSq1+3cdt/BQCzlvleT
wVaASEIa9ZCTIbvibyeMABXbqQoS2uO6ePzwChsfN8/gBtF7POVfI/vd/AgHMaUlVoBt+Gta+R4M
iVFY7Scc3teXJWrkABCW/SrHJQpq9EWAgGoEi7YuhnyczaAi+c73znZdQbSkVHspgp1MD6+9y/Vp
i9re7YDlu2xjhuNWCB3MgRwJ7FvfiKtgV6EI1x9D/OFJ/DZWaOYEMquDWbQ40ZI5lGeqYC5BHV3N
wVgj2WdIZP1VZKLi/EYDwhw92xgECgk1dn+zdjXp76uZFtANsiKaUle3RAmEr+uGfp+dPH8ouZsU
xoEK54UV8y3V7vVNmZEid7rgyM7tpnsDLfNVHR8fdiqflIRtfTyzpLpazUfkJbbKtl3a8NBk8Gci
2/yxUD55Mzrns97DN4uL6dI7+qPA+UzMxxH3UZYz+olRclh5GriQhF9LbeVqTGz/wXr6fMRzhJXP
Fkx0YTTc2xC8+U2q+5fRNmR/veVN+gKf1lUkVUE4A7ppvWhx/I93rvARhL/EbiUi7/iqjhd6kyTf
WZyfZ4kv8OVxPGbXhFjoAw5AM10OIPRueMa/V/TnFOgG+9VEyfCFirVU9RvfJgxm0sEvfnyvtDqs
oEJgIdaymR2fX+qqAa5IX4coZo/gWrB313yDezT2RxSrgOKh6O2X4s3EfSPH1CWOR9chRLNQzM/c
ufClA56hrWofo9pCAxxMAXx7Jp9pZn+c4KsBXQpejm5H0kK5+rkq/k2i25gjGySd0fVXJSiqa7v8
s0RfncBgFXJrxEZcuc/7fCvgDkAelML76MQVXkK+d+Lxl2Fg+WMJxBGvZHjxe+sXNcTAzR3/XC9M
T4F8tG0Uyotv7LcNep1qdnxILEm2UADjT04QZU7253OQYEKU1Yi8XGgyXpikF5e00z3sn71ih5ow
5YQejd7X771nYxrCX85DfIcyQbFSPZ9+234ePywoNV3bUFCpZIuItOLF/Vg5u/5EfbkQYxzs4EB+
p3dotl9OFyXtX0mvQltSmyl1K6WG8ZelCeEUDR8DxWjCg67b5dSrmRqF/yGJnOUYqufPtN+NCoDg
W1Btqih3cYhumqJL42vJEPnjc1m7e6bDgA+RN7zkHPLxzBchnzUNYxaBfsdG9tTZRaqe8Go9G/qa
bojKaLN2FpKOcFUPb+abK7th0tTDzindVIPBZ2dMBm0amwXvlm6fVoy+pgByZ3sDAD8TJQa6uXWA
thYDkxv8uPbvkwwD+D7sQqleuNRXpdNdkzLMPrXmk94Hid3gm/iJHuCYiB/4oTuiC/Cu2yIfKBZr
95I8xrrxCFc5Vnq8kFMYtMH9YNzmxjnRmQSQbL7F8eP3B7F4nmp6969Jd7GC2X5d65xAXHcwzyET
pGiHdLhCh0Msq2ado+yEz9wXWMjIt4cz7cQ8pqLUIOv0Sr8HBwk8d+Aluz61STNopRJQ0JNH7slO
iUOIMYC5pwSWQSts7mrJkdGBb4EbXyp0bF5Jlhsn3qL0d7LxO996V8YFqV+Pp8MAObUqcoD53gJ4
MSyGcQ0fDQF3r/PjMf6/j3SPBhuZxc8AAY0l36Z5upO940SZfTLsl48vBi7UYxljRNIcXzF/iHdu
Hhrp/eCg+tRuMq4or6nvt1ql/f+zt1jaUaf+7e515GxB3iAj6EQOnFm4nTWztrODjVt4hbW9SNe4
UD4QKzUd7q44APqp3b+GYASWp96GzbkF96VrpBAI0qfGwIesyVNtHpQiY7K3wCLDzuxpHJSWyMCH
Tcvi/R6X02eivS5qbxTJ7zKemINTCit5G+kP0Xlb5L7vKRZpNJZRkr8o5uazTSsGmMxeM/M3y+0m
BYbXZrxijfNoioXQpjLnIaFeTO/flnH/vnwWChWjwPxJk3+dDi1wQY0yVY8tJgOmRR4qL/znMrYr
goPAsgwfyhw0RMAjk/TUe1uU8O1l68gGHPLEFpsHPrHl1dG6Gvwy+e+ll5usEn6v0NDv2ZVWh+ws
o8e0wBQHT72ltpc2wXqV32DRn8MTDXLDln0RLkIwD0H5HeOSxHotXAeId0/YNasnEL9sV5tTQsOe
opAwgzJ4sN7R+rxLteYcZgZ5hbqo7z4/iD7jR1rOFwPL0hEznvYvDmEThcCNQyMKcL66xZibRmuL
L8GzfMkXjsiXPMhogGTmJehqvCJuJPebQG+2rXMeYd0Q9TQnvofuuBmYtYQ5O7t7NgemZKT18bSX
F38X2h/t7HNTHOlImFUGbHsej7CAH6Eh7QgHcrbacanqo8TaV2G12YuUiZsm/YqtZize4skX+PJ6
kJVioD5h7FICVdkJoTvLZh5WoIBVCrmEwLD0TT49EeFlgW7ZqmkObP/VuYtzH1WPtwlKhqcc0WVQ
9APHdkNHS2dx8LyKpdyVEE9D5bh4tmrDFcM7683j4lPXZW0gi2abphtTe2kzUrWKrY+mkGO1Sj1a
DilQjmYhN7hSUz8JLiClzg6uB3xY4W+JBjszfpa/4IiA5IuVORml5fNCJ4x7YQkBfw1ZqFaqZ1HB
TEDxnHKBNuv9mVn0ADXZzXzqNghZWHK2f2IeUtMe9/QuMxmbNho/F+N7YOxfaZl1tlum/YTbT86Q
fGu5/3K/HkIXHAbLptGwnWc/TKEh5VMU8/gnZczpE/1a1sSHHBujaK/x6B5D8+nrmK9SPsNCjC46
nGvWdfzXVJT9703MyeTGLi1ZhvCiPrMdYAU43Up9TgFe4NCJaqxSi6uT94vua4ZZctMpY9gL1LU4
4AGTWCYFwpwSKpwgjmABY+7rxXhnWeevm+OQFdlRFdqHltCkYbcGHl+GfaEJg8IxxirC0U3D90ev
OXL6xOUGq0ZyUxZWvUPLSEthRk2frNswgJHIZStOIKrLBpphNHyc9Uj4+XDP+Rb9w3TcuH4zQuVK
xit2cfFZVZaxiaMvlBnAuhDG4UqdkGuxPRhd+bD5xedH941gmMJLauh8uBe86Sb85uVF1cv1Olhp
ZkytN4yrt9NN7vvkziM8hDtUCAhVCvA8yz2au+mOa7V+J0QE/1Hd/h3nqRsVp2NlPNALbjjeSft6
bleO2WuYMkv2cv6hb0RT8vqZiOkUPSP6NhEXMkdFFP+KMy57KRkbTY89NePyNVw0wJcj4AqVcxk7
yEsrEbpnbVU9FSeZ5mtHshwglaAOd9Uxct/yBGivgt/LNsMgVg3TeaTNCi1ZicRZK1GWQA9ErMpZ
wc2dz7K3ST5Iy42vV6eXW1v4Zz21bGnsvFjPfOjAuWE1JaioRIT2ZYOBOV0gfRFAFrlhccD08Hwr
EYTOqGy/21VhXuUPrBp4U4eWBbnnozmbYeoSm3NZ9nlMFgX1YY3mEsG7tOmdJ0T1Pu/HvVRyUEWV
MI65x63fz5Ps8+GFxxXPqi8UKpB7j0o+ynlfnFqbj/L6H3cSMMfjUjGfVEZk4towE7ANk/BrS/bP
A9yXaYlmsd5C7UD9B+yrmnlMxIQNy1i7OP/O3IIn+tFX7gQGy8GHCQPtT+Z/Di5CQw54VS9nf9TQ
PQnwVY9ObYS9RDW+PcVQUg7bWSFvaL8OgNqgTzQv8h8rWjIYpnUUZ6J+gCuAkl0qP2jPdSPc3/Vp
zKHKTPMI8n5rPH7mc8v+Vk36W64DNepVr2/A0qS7FqmF7MpBR8V/YNBq3wRiim7by3+TV1bybRoo
9VeNz7wKF1UfW31DG/Btm5FeSW7id9gD3XusLYtacVs53IkLJ127KGgR1SmPCkx8/3gfnkv6yS8T
b/oQBIgOBY/ph3CQYzFNN+WsExw5chR9HuTVyprEKvPq0E5VwUCTmpfpNza1ngdHGBDuwKbH5+Xc
aRrWL4+Ft1dNjgsrQrp6ZrUv8tA7loDZoAKCqKjxw4OfVhzCUrGZIOPdn8OOSZyi6hTsBm19gCbd
z8zTC60xniryi58dzKlAEi2I9HpN9p1EwPvNA1MsNbZTYg644iVk4YctGTNdYfXZEViM9FNUbPxx
7YoFwG1Fxb9EuJ+jFEKo8/9IaKKa6Nr9U3Ch9naMoQe3F40RyG8keEmyTxjPR9HZA6daetBXo+IE
KobGh0S86XBqL/HLxKpZC5+yXo983zcpybkPSR4LtUSmrdrJXjfAmDIkwlstWoyUXK2gFFP+KplO
S3U027/zweJ/bo00Td+8PeetJZLvBg1rbd1lWtOP5pcjXWcI9zMoWe+NTvdV2hZfSCgeI0asstx8
/l1RzH/dvQ7MJHtkKcooF+k8X494vp1l48xiCfNcQ39VgGReDzYXGkOH1sLnofDw+EUSLWpgiEQg
4IPqY1bVMc9+jF/1ZNtG0dBe1bld15tO068kQs6+ZZMX7daLAy7i6o32WAOruWAN/K/j0A3Fq7+c
YB1qnZfjUFaQq/4S6HzL0L7E5M3/egzdusHvZKAEBJVosnl/VuzksU7r84JImr3RlwVQTKVP0bi1
l8ogpAJ4LPSH/8edW6Zb3j9bpXEMOAVKjxv7odeP+jqOkfBAv1Cr9qW1hkqxWiFxhjbrKxpCeYVM
PLFi7GZ33rQlLyFNN+UDr82uTpFp85xX/1wqnaGRSybEg13ABM3DC7TWONAMPksIYmno8zZj8vDJ
6c4J5rfmTtbsnxCRK/HSSS4gOsK5G2YSUXiBk3eZtLK0xp2va0LKldN5ErU9ZBMG45bBQV6GaCwV
iS/dsanSLPssh23Y+pec3Qo4lY6LDoPAmgbKPph0bfV5WXrXLzadzOa0tTAoOnnvHPGxsFZ0DLkz
FUP6LEeju05OhEWhvAXKofaomX+Xr/dDeUZE/3AvUNte/cbKHYcGS0zQbEIGgyjLT1OwWV8/NjUG
Pf7PIaWiOB8SBhuuFH18OgS6vpeMxjGTnNMOMh5ESAioCCgXgILwULoxlYNYyLke9wjSH66Ix8sr
yfhu1wyKdZMWwSyOKvEomydl/yYQq0T3StHGOcpyNJjvr+/Q1x6CqiY0obXCHdVazCPWPIOUwgzV
WbHgqK3KxCRS6gOEbRvy1cdJjKKfm6zmPbO1ijOSDfhKeCyySKESDwZ5xUZcXz7WuIa6fSc23vjC
SjJK88gH/E5ebZCtgHOhbcrfX+wMz9sTj+6T33GV5huqYTbZMCAY8TTddlDuW7xnU8VTnvOVwUtQ
DjE1V9th2KClpiM9tPqp/do48qBOrXGlFz8NEVm94vUavzR1TftFQXEgz5iwymrLcnIo41v0X1qx
TJErmaZquywm/bFEHLCRAJj/g+Ee+3920Ka2q4U8D06A9ZgjJImQdARmnqLdXgJf8fwlrdMyaX4U
vP2i45skMBu2ph3N6m1zZd5x+bSdMJSr3XTduG1RP7WiuR/eheoajzM9lR3NhTOAX1Ctqrwe9nmP
DUbOkEDEgKVnaoarGmywQFhNEfW8a8SlxwFgXM47ym5HdHGB4uTY4yldz1kkg4XorJDw/ojactTj
5lODvs/kX57kkagfffo8UClbOpvU1U/VFxUTOe2qzhxqblCntEr+WtV69x9XReAb/YtL4OBRVEex
A4eAvyZdqY317yWc90B523IwtN6l31pTmCA/pDKOcOJVbKRBulu0KYqHLZnRUtO9tqj+0udfOPpy
F3iDvTGk21N+HHevw0ZUsBRnyKsfAaVPcHU646RKH9i/Y2R1t4bTpF88YMq0Rn1SA6rn7gaFT6Ta
HJJh+47yuYjg9kDFeD6iAXEBjDkr5dtGKTGle7YzgQUyzZiMtLM4iCiVvlrRwiOQvBu+DcQPvGaN
RkgXvvYRBic7ysxW4XQ3M12X7u82v5iEr5gnpvu6o67ABS7VH7NEPamBxTido6CeqtP8FhYAfOSl
pvKC5H1C+lBfD/CVPoNeq2BtKq0yrgi5dLpU9VDZt1LNWvMyJ1eQcqW5UKWbv13QUjSSbgZL6sTZ
JPGO/wyC1CAwCqI/Lt5u20qDltNraVJGY77Qi3dexMrLDNvxTY4l+3V4pVprIksCOFtMQH0gJIDU
vztf/4sVwv0IL5zKDlrgXRBeUfbgWU80zTqMUcthAcMY4aFiBeW6Vutuju4xkz/TTT/pivfGwPpf
rQgs8SM6xzyIjnyx8VPfBHlvUThKAjlDlOBpGb/vEPsxxAEIiVR0iADhMwbczDh0mMNz4cWQ2bIc
MaTkrAic8BzwLAnJ++gGdxNybRBGt/VoH4EpVw9LNKp963pGJmKi5GlYwTzYbU/lb2c+Iqty0bCz
PawOm+jmkVsrzJamerjhNsnArXDtnpu/6ZZBqFnkbq1NglaYVpoM7ly7KrFX3j/1AHVUlQKuPLpB
yoyG5xutebIEruzBOXJKLwCbkMtkS51ukqcMn1ykx5UFDoFVgPECMFl8NacO3UTGL8MQhhwR8Ghp
GZdGTD55bXGNXLln0SD5vnboPsqztz1vEI8EwORPwHc0SXt/C8b3HUdCCC+we4SUkqMAyJSQu8FB
MGSks7PRUcUTUv5kApF03dNGGkDC8O9hPHqb1b4QhWWsLnjch5gYooGgSGGgWpBBO2EEl/XF3I0+
qNSjkQQyYftC7qk9kF0WTY2MahMksKlDGhIBxeXZsyLSFbXoK1a4ODxQ/hnpth1W6m2vCMSGX5oq
AKR3eZ/gNO22brxWJURjH32AimXnoRs/2xji2VNtDDQGNWz8cI6nUWxf1PKKNBMg/f/Lz0IEmhT9
uEl0BNUKB3S/ussDoTAgZswk8KkemtYQHRDQ0Hezz2uU4SFCBZrTtcF19p2ZoAXLLL3b1s+fcJTZ
qlrzaBpnkf0E0uoowatkaU1Y6yjdQe6IAjUyGuvumMwBY6cS0JZTSFdbj/yiGnyFnYrmMV4eCfFt
IEHKREpEbtdAcuQK4Jq6EWOk/Qu+TT+P3zGQll9kESRBnvEWJdnge839b3seOURaaqtMyAGmlnyn
DQ7GE6EvaQemhkTRu0lFcRBn34vw+U9jGrN8o/6cqYRNttw2bTCyFlK2kaBzDZ31W2CEdJal+58t
3LqhHxZWPp+uY+5T09Orv2Fvo0RKk7LNiOtbWTGJKvn8/0xJDFU0nsQYF5mNHkyf4KDBVy7fvAdZ
VLsBODH8wMDJiYrz5IU3/UDBxJfV17gTZJatoQfJJkXFd1+AQ1kuCxEYCnxgP6SZNr2KWRjlBKkl
N6GjzZoMu7Bf1Q2l3i9ITLmOdfGNzFpVYSIKoyPgTyDjh1RfRikftIqUWHcYCOz6TR4WD2Zslg4B
dS69pYu3VSDVNN+X8SLhLpGm4WDO+Erq8Xu32Nh7VZO018mwWmpdsbKn7fftwPBKfD5lZK+Nc0n7
d7Um/k+idrWp3X+G9yj4ZjyZ0xfw2AT4oJ4HGKFA1I/4QJS39ax4ghUr1hOLkOX9xmf1m3T6Q/vw
4OMqTlsADgPl/+i1pxrLE9+weZInGahX0djqF6qpkTHb6XLuWgUrQxAUa74Hv3kjgYl/2y7exr8w
3nzNagEpoB5XpcJr6IJjTAk9+2ox9Id3OflaLRnwDg3Y0ypxujP+2+MODjh25w0bk0JHEo+1V6aB
vtzHBlXrTxehsh8s9hRc7/wz3OyTpUusv6smsEcSjMl8mAgdulRU3q2tW5cLjv4Dzggm4gEXOYFC
s/+1psevySSIQgSSFy6NjOJdlcMhIXWTY4EqWiJv4TYsvVJCPBjFr5SxDk7LRXbHZH4kEMzqBh1C
nFuRfQKDFB0Lefrvdv5RP/in/5W1f/dBGBi4UETTpPimUycp+efrbVWrmN5dvJVTM1zFNyd16d4T
dn/OWkRFGEVAnJcNBVudTBJUWXTqoilABFe/bHfC2ZBW1ZAFz8MN3XbuHW7CzEvErVnUskLWNwuO
z3XY14hUFFuJUnIG9kO5pewgcRlr+D79xw2gNTT7/VIfT+xI3hdbAez2VVU9i9vwryhRj0Z8t1qq
dIYlo5KlMVyGHi7L6GMacUKGtzl/aSLqFFdlWneoxYjEeqMLwKYgvfZ9yFlq1I9ZXu1R7nZFC7VT
r31xUMcnmf3Anxxteh/lVolziemK7HgddlqHT4qXI3QiWqkpR+U01y3v06oC6YrujDz3K6zuX2Nv
+HHiYnGIaTIhadExqAdhA7E7CxeIlz220aGLWdpiaIk3Y+fyRnImXcFV3BjTq54JrDIt3J8Ew/ay
qc+9b7d6Q1WDqJsPN0IYykd26MF0PdqX9vvn5nz/H+H687urxQRltyC9yhGazjIqWFtVn89K4zZj
j3A515ZnQFWp6Mo6osajq8O0/UKWPtFzciMiV2Blg6hhg6UNwNnJ+469NWQHKv+RkcmJ4ZIU933n
wIKd3tKeGMDctCEAY7POedrqtwVomFGppdTbV1tfv/LQ3M2j9QdDcV+MP4tbpi5Qaw31yB7tMSLH
HOeieVSGFf5tjZvAdyqNTxzaDLjDm01NMyAIAazZsf1VaO3+4LGciRhrwU1xbh4DC7dErfZLlsOn
hqS10566LEAazZAxwErYcnHTfR2Gh4zwV7m4Ol11QzFZb/DhiT00iJaRYpcL+j++C9dv/gSkJtsv
L48IkRfF55c9TQPzzyHFBNKe9Kr3dx0gASbOKlSdaxrnwLJyY//jD3TYdl1jH+uAVpMK8ReDm89P
eovUhabTF/yw+lRK+/Tm5sARg06cbfCKcEZbhPMQHSabCbJ06lrSwwGmQswFkF66UO8P/Il0Jh2x
2Gjje6dnk/X2FC01BXIqxT1lJ4ykHdXwsMdC+AD0BNxXgT+zozRprrJvvHf8fyfasfSQGlXQp22F
ajwy1UivKnFBpajTgX4lyFNOv8yxldr/4lAN6AdcFYXWW1ikQz28VfT6JIJL1zvHeZw5rFIMLTV1
dGumq6ApKTZkYJ9YZWatj8E4HhBi2M7acoLr2VVYtH2KzYdcgpzUhJOiliaw+T/JYQDuAB9jdRXx
yfMhf2rWxJYy+8EVis/4c3c2NcduhaYcQUhvvezyMke/8Pw3hPPXP6Rv2p32IS6w9LcbkHcPN3ss
22aT8Mo+YGkBjtYfao9eNO9pat5u51QNkzv+P1dLaTLmTwrlStewrPNZxjd+yq6c7mEfTtn+HfAf
GGVwt1KwFDnUzUhufxQtl50Lsk7p7F2V30HGYvot4AoLrzJNxjTyippN4CjO3bxyAp5Y8sT6p/kf
iSdX6X03EZk7YXjMOjl5+AXegQTiRl8mpXlDThKrK2NWOwk4SY5o55mP4Z8VsMebtFg7vYfr3yTH
c1kK5u5917WUWfy7uFah//06fjE3jA6rlEG+p/B99KrhrVztlubPEQ+v209l0SNUfs2auZygKlQq
O5BFw0zDzmNzpVy8IKLoRXlbYscQAhvqCCjVqw4vRq0Y8YiYLFrCIZ8Hu/WAmbZ20S4rGuses/40
Smk8JRwDsxSIJ6ATsmbLZ0VtgeOwqgbOV6lqPb77/BuEc58Xo1HJ+7glOzltyljlRYvM4rnTk83p
ucQFRSQ/ru1p4VMaS+sV4HkuvpEKxdHOB1yF9rvWgBz4FhDiJGvTlDjliIVrfFqawo/OV8VF4pG7
uEeAjneiu34FYWn4GbrO8uawCMfUxUifrtB38l8eeXWVE6WPQA0LF/LEdA97N5H3tBsPghlAvzRM
BgRZk3l2mcTEAk8wDvpCRIjj3gWbmCCOw7YcFGRBzEYAFMhQG7QbIk+DLJ5xWZnursA5zRi10MYM
da+2jQnMyceMB42/wIHxSKPkIyG2ENjLnD+X7K7tWWr1zrL06jch23b8BudF/DAPcTCw1dNOIzXx
3IZBGyAvHCIQu0wcaimKqYffB5t0jvnYfl8DumKRPTVuN5Q0uDHhCwwLhlAcshxajisHXnznx71d
DDM+QpqTC3xR6yChycCcvWQedQ2BUCf29fqDdDwfrGZntJBiIVghHu2jsm1nklg3NcIPLg5K2grQ
Mh7gNlMWBzAJ5RZ2c3bGoN/chsm2jf9FipEf0WPCz6ljXeuDJoAuXLYMO2D03xnpu61LdHCAZIY/
08jK7QbSYaf02M9N79CU/fGan4dAaXqzNsQ3peLY1iKJ1eR3orLobqWqkOpsXzWZapZXtHQgye1L
pBRTUKX9LPpnxENq2KZNDOyoLnj0Z+vnCHpVi9yM15VDU+Uj+J3j8nPb1XqXonA93ue/O1cpgy4h
XTj6huwyGKRKhDVdsiO1WkIKUVnwpUow2mU2DODTy1EEu4fyeLdPIbaYDp3x+RIEKscWGcRTxsHS
Abd6lNztUr+rEQpOSFhANOqRN2GVtQSPr7PNGgSpkuvl5/Ft3xAwiB4Whd3g3sYLhV9UqGGPUcuy
Xdkbw0n1S8gCEk+PPV3ZpVrc7jbhxELKF5njMtXUuEPanWMIR4CocCkn4PbEAugiUQyhFcPuM9Eq
fH7wZDp6e6pTjXfyzMZehwNjoQHHUBVPxpcg/vYJX1ax4mhf31qm3OYnymcmO3Eh6voOpnjfB47A
r/8GJ3QncxeOH6u/eaAjyUo3ZeMe7xjFhvRTFG4VhTOHi8NJojK2wvDJs8cVRhioXcQ1CEo0MmNN
IGprIRjuCvDeXH4xA/ociT1AvMmd1lTmOeYPUQb2B/yIK05kEoezuYScDhqbhtO0iuoUO7KGbTS6
xLj7Uu8DWlYSK5MDvDfP6poizD78Frx7bI/Ok7s4ju9/B7lWW0ubnZRAvivadoAJCRmhSkcAsIgw
/ySW/Pcb7DMwVHW7xymL9s+8HRj5hjGS+ZgU+3L+28FdBFqzJOEkzwpy7czRv5kxP9XCRXdcKWyX
KqQfMl9gHqvEDclp5ygZf0gkWDxhNGWSLmruSuoaH56qGzqm7uCBj3nWsV1JuMTAX8llnp2I2CMP
YV2wdP/9IiSjJ3WtHaflYZsRdogWsoxLFGbGCd6xQadrHBWXXsF8zgRdshoLIRBKcZwHZLPqIV3M
Q7tdlTArh6z1uAF9CqHWMRutkFKZKWxy0SB95wj1dq3uyU6bNtnHn1WHJgyyNYYv5d4e75BEaonI
dTvhP4NN5u54h4yPvpeZykSeBtYjfqp6KqoxN2fGPlz3pAPnrOv5rgjwMZoj0lnfvv+ZIWnKAvXT
YPJKMAXWxyUxaX9sOdOZxAxevKHiYuO/RHWJX5HrWqZff/CHW+tfNzlwMw0/YUZcAD0oB72daPL3
1VDuT7dAARG80T6UtyOwk5gdSN1bsBHBXdpEnmAzi89Pzm8FFjolPf0l0MKWaE5ZHfco5ej5HxLp
siyS/uhJF9KYTf3XEpYNnphWtefPNngsX8Kw28Y4UtV6ndiuFEQYRRo7r/K/y2c9XmX2cU/hwnig
D57MvzAc/a1e9+1XHGYffj7wqttMVuV/yh3rMfFl5C2L2rSmPFTZ6TCwS9oeI1QbHTzP6+MyIUZW
B3CmUJEkfehvkESPI57M3mvcB27ZsJOcHz4WFh88SxCHqi5GD9jEr1pnEyC68wl8+0D4mSD60WEd
xWBZonrHlT5mNl8hQC2Q40yYDZDw7DqcqtTU4kdKDRkfsemE987HKkFY1xiYy+er60pdDwy6nctf
rxoOYq0jcPVldaWxvTHX4Uv0ySV+Myvs9sgmNzmXLJjvd7kj6ZxD8OpJWBojrd4lfHuulQHEyRkk
Fmno6nSuyIR0Bczw1vVIw8sMMY/EPg06EywgWsWhUryER5eP/pXTpWmbZzPRBS5L3MbcMjeFwp//
7d2rXOQSe92rdka14JYdSTCrhiI8jowbiU9ftCtbTOPwHsRd9wAvORDOEpUaFXJCgxw0fpxUXwgR
8N/XujTZewGr/Wd2pYqoUmZsrmCqLFMG2aYOjlIo2zajLNBLX6pbLRlCRvpRQtRxAU3w7iMwSU8G
kZf3jUnLOGRC2CmvgP5Bv8itp+AqjXUlBC5rSJNCU3EZsrMcVR4QJrgS/+dYstYTiZQwNrb9SWFL
xinpY3bmy0Zxincne8s19lf1pTNt49VSUZJC8lb3ljf0GgMnIg+CNkhutoLVYO28gCuc1wFbLNvT
336uDm0Kerx44ej4qXNtm/kxvUtnPsNqkr8cevxuKxuskODEKuNzdruAR+jwexf9I9GB/HjLOKlJ
WEjJAEAIf3/MzqZAzkt99mP3/cq70AwJ0YQuLC0Ivb9n9lR2g1ubr1e4D7QX06CNN5fo7HYSogaI
T0K6rTZLHLLieGm9b/tDG+OWAcGp+XaQQbdU2X3OekRzX4yVeFveM3sdhfYbfxE/f4cKSd0ye7FD
Y0d8GJPZ8u9NL7PnYlp5bTjeqIEk1TnlqR8dKfYtCNMYPKzB8gAXtHGRfeFWzvjv0o52SQ1F1Bat
Ul/yflIsWVj8wI2TLxRu/PHlbInNq5ugJVgyKqWUfkTglGgW1IXhDjxPUaZucbBKG7JrNq+c4xg3
/MH6txiJXMYKkisfIIJjyRcgJgDZTeqrzxL0eKKyjGrBSosU9++CzrVSgFK1IzjF4Y5rPAzV2DJ1
PpjLulE+mRQcPUgfXXpmkpWlLVH05o8P8Kg4LtAL92RUK3WQdUOXDgrtbQ2t9oefOLLZ9aTWr0EK
kyDYZ3MDh3Q2wcz61XlVE/Y7LjxXS7YDDG1ckzJx4qiFwwn6XRcbtCT/j4Fub0HtwmVmxb84W4H/
Q4bJn9fKop37WkSkRdRkCOzABGRS2jwmeXj/HPlQ1ZVjWjcPPXFp6vHVFC7Kk1l8eRzarpzMP4ID
sLB+z0zSpF1ZPWIbfgiFK/wHvF1SJFrVyT1sj+ycm41hpLTsMLhQv4G1gFd0XCLda4HC2BmCg4rZ
mmNaHgmAs4IVwqNEut++GDwBQjeujw7hj6xPegBYjX97d2T/CHhgd47d3bQXE8hs4Wx/ExVao26z
AoiqIs9mAlUbIqAa/ZigVhezJy3kgumUu9JQBrMB/gj0idpEvO0B1OL++DuUjKdrUjbKkqysOMO5
FJjC3brr8ZTJdat1uBR3REZNXkM05FHMO9aXAK1zPoytrN0liEQeuWV5AMxuG97c8cbU1o8VBvTm
2iABCwAoqQCNUFYRHZpBvP2qTtmlV5aEeAf12gjv6ArXlWJgezFtcwwyArxyJ2AEm+deevm/bHjz
HfyD02JGhaPI36ym7j+yY4dZvVPyk+3AD38w+YLdTkwc5lHGsHHHbhreTq1jfQy/twA7bWSRTuhd
DM5QWW2S4YUTPMEkirDuvxIJkZywu17x0yS/6nToUflqCKRdUbtPdnAEpxoH6Yt+M2/JslJ1FMAB
sfVT6g2P0Bqv8FZqAxfZxVjZG/5bSLCkCGdCf+2b/PmSBUNB0srKLxwL8f+uRXoq0kQnVXvv1kmn
IK6sjw4djDDR+gsY2HXPQlBmFr7QeWl5AKd7N3MKOohZgO4egGSAa//XCgnYXocDDJK6VgQ6e2o9
mTLXjSjyTJzpls9DGhjgk0poiBRzKLtiUnEBkBXaWnQOu5dfWB4M/yheUyq5mKtJBqH+7AWu9nHA
FnBm1/PROKb+g8P3PYIzkLU0xMgT93nL62k+aIl/Qyszoif8GcvbKpljZMynRPIJEQxtDHoo9G44
U4OVLwL62WS14HmIUrZqomBcEZr3xwNMEG9TgWqYclyhIv2OOWAlKFC4GGrdrnYrrqK00iOBkfnz
DZMaT2LRyBMKF7CD6zqVeMEMNXMRvWuyr8g5qwLMAGAD9xJOljPl1N/0z6wVPC1OluDEEhg1rtsc
/GrjtoAv08F2L7Ss3uOXUk3ndJN4ZEa92xpmJBncyIt6CbE7yAQDUavsVosTk0EDlyV/ZIkF/ycO
i3hSGUJmgQQRm57JhNgYujs6gMZ7lo5c+YUu/277Kbp+pGk+OE3VPQBqCiaFhAGgfnO1KvVftI6J
48tnmQ5Wf3xn9tptfngCpP3kmcGgRUBXMf/w34oCjj5wLhSES/NHMMlwtg9rdc6DMrjzqIsqS0Xz
BWdXAhk+imftM7Uo4/SkAA2xTgDPcEFXKa/ZtjqjXlaBS6osKP98lNbsiYf9osQ8P2EgdmMqIZFh
drAUgZu2Cgd8BdVm4a87AxcpWRVwpRCyFRjWnKT9fGDNn4bqMtc9dylOvqXLxCmHl5hra4FC3u1R
xlee1iTtneYq34ixPYdkIcZEDk52srFTyXokYAqJe+a63CW1YxewWvHLHtm3bVB3E51RjLtcadeI
LUNdNZzy2sBt/gqmG3AMDo6y2Fy0WupEvjkuynipYQ+lD6ypAj3KhG4xVzafFlSjnYjqvw4KjZAm
h+ON5QLmOFmMkkIvS8MTzcAMlC9ZKETVrdRxGNvgIctqT27g+bsW+tamivZlT/098pOmn4UF585H
90vXgAE/FUziCTgVgyH/XanyICSCfC+sb4s/4obAvnkfNj9XISp4+c+L9nSeei2EraW61i2QDZQl
HoSFkzs83IwogCHuGKOoZWM7QhNBco5VuhdMtXlTGyWFzqVRXWDNvBL5ko8G2e1xdWB+YgKNrDpA
E6cJ0ZnSVMhcDVS+m5VLmSuXURZW2E1DCqBWK//Ztf/uG11kfjLwP5pTLTknRwXy+p08NsAEplyP
XYj3l9W+bjOKOrjC7nAvsnS7PVvJW+j2p3j5K/IpIAykSOLZwW7yAd16OATD2b+NktDSN8dKlmz0
GShWLaW6pbMEnlTZf/g+t9s5366pW2nMyRzog/GYf2GzH8HVkstXxmsN0LKDK94fn/5pcFwjRR7l
hCpsXd1fHMnpIrzeXNswMMO3O4twrFyH9owj9FiFT+Syf6F5jBAB3xV5ZrRN45wFBlCynArHZ0PW
hoJAViQFVPUE89AF2VtxtJ4cR5p05TJUtU7ob7aXzSMfrhIIsQmy/OvtNpmqzQ+dZF/H+JvWKeSu
ttnyMjPTtj1O8CqgPaglkqdvHpWs2tNc+ZpjrAJE8amWDR9606s8lLj3VDIixFxXZKUgLjqOWjCe
3gHDLx7GSvKW7iFYlHmYjIfAquUKUWdvITMZbeQV3bHu0sbu/fRpIiwc3RWb/71H1WKUH4Khn6wP
IfEBdmN6n/U/FeVCpn45WRXjIMbQLqnWOeCF6K/Q7IZepnj3FDO2vUd+ReAOEVM3oWSbTFmFWYQa
u4br4PkoeM72DUMRuvZvinQf2jRE49CfyBJP80U+O/NIWJhy4IvseUqqFHni3XQwP91R69RZcGnN
NCWxTPKxMCREng3oC335zZqnNguGbheOW33/Rsr0jKDwcXxnWwcikiGzweifXaVaLyECv1E6jhVN
Vo9b/ai7TVG8yqMSVL2hYLVVB2SAnj8v4y2bsJB36spxvYvfaXtTpbgScjRDLW5gZITHBWT9uW7i
zKrC/5+x9flceO5RQ/DxLs32WfaW8AnKjPFGD21K+3wKA0CZW4wJPNpunA/FWhw4oxPHS733LtK1
uEO+dMBySyn9a7HPq3OfwLNHe59UFC7Cfod6HZQ4UN8IvFoBKObOfbSIw2kEgaCSfFJ7YK4V2dbq
Goy3UXPaHzPQk3Cpj7G+SYhsfUfbSwDe81Mtc5TyrV2Zv4301V73m4Ku8UTc9f9uEC9ZZGxzE5Uu
XmuNnGWpoDIGKMGTVwgjDYCURLrjciNyW/9ql7MQvajoy/bbusrmnVrCscOkcxWnWWqLP7ttdIkM
+UbYV7CAs7Sr3De7AaAiJZkIuRl2SF7h9qdLx5XtkRU2rQQvgnmNMQnJsE7Wj7lE85VShaMd3Ok4
1ZhR7HJ90XTW+0WUKxzGZfUGQWfIrIXH4b31wmIAW+ddWDXGEmVB4LhP+ZMsnlCo2e+tRYD4d23M
0nkZe2Nt6QaEyh1U4t9kAkEIjk1QcfMVnGzmjw+Kfg4em+I3GhHwsV9vVtVxut/qZLVyo2xzVTrx
/TwP3DkSozw0EvdkeQ0zjszcPhS+8ZfXzkRlWIgDcEYamJFatcYEPSAWNZ2yeZZSyIvR0OCVeJif
rz/CKM+9eOZ5JTiR68hdKQIWBEUTBbcekjOuDVziHrZZaA8ardrh9wF9GICt6NZByfMwDeSpLkjk
Wz12VAMYR4+eIqCiH1LweufeMC7tqfXohA5JsHS6V8km8AH3VzqE3DafRK8IZjc5rjp4V2lArRAB
Z1HhKSIRo65Ms2441eDRBipF0EQzz6UFpjs+BRJnZYEveO8AsPmr/YF6TKQxDR5BZbhT/JMtT6W8
6lPCIbCzWCTVwXftDRxSeDl3n9912Fq2HWYssTAQAN8hN6sNcw2tUWjxu47NrUCF6K9SCs2cT5zj
trfykqBgdbnMKQvQ2ZMCctFJM6iCJSs7JzmmBj8xxR+Q8BobLv27BeMeuCm2XhV95PYoccw7OvB0
MIJbQaOVjwXo9gnbbcfEGmhzsmGneYfb7dr4dod3iRncaP/IdlpbnA94v8UqbqOyZQHVfI89Y6ye
7FqoO9YW4WiFypMjm0sKn29BWJOjkvyDQcoIjD8ibWvDY8sFLujy+StwTqB/vRpmpI0deVRU/uQs
qKHIzjh/0VL1LT6/k2gdinXWPO4w1oc4uYnUxJy+5YXmYwidPDwQlejZNVlqHPXfn0DLVTbcumFJ
7owmfzAnblUMMNBN492gLTZsnV1yEl6c5xyxC3RVRlOH4cAxFbTGY27m6xft4qcYPvd6Hx5RdvRq
5PI+7CdvRR6Kth6toQVhOV3qb3v2PWZt4hleDjuLoMHRDRLSltvXwp4uE5VRJ9xLp4FwaDVPlDdW
Hz7mCBWNEotpyZp/bsb3gLWQlXv/7AWm6CmVsItUpLUbt+Pt/zfcK1T/J6ApGsJXU0G49Dlsu8oH
Goj8F/6ZeYJWdgFdyv0wcbMjZDM+MuMxgn0yI3K+XGeefAbRVc7eFuIaSfV4IxOMywPt0ijO0za+
IRP0su5tYGnHiMaE7uDfRrW9ImayO9/04iNhuHdzfglVjbWKlhLtsE9/c5HssmguE3Zm8SXI1l4z
iWJolkNzpmMTIACEsHQQExD+kDJ8Tbb/WJJeyfzJrckchHH57jORyC1YG5eu4EVzHwzavBK1BOin
v0fmiiCmHz8dC947t8UN0XBdCq8ktofExm7KjsX+1m+g/jSacvzLuS2zPektBpqB02hjEJM8U82Z
KAU+NNDj+XJkUJiYCeNolsJE6wHxI05NhhCnf/Al/sM4f20ShyORA2l6QMN5RdAUSLAEBD5m5XJ5
ZWXncYFfU8IBm05GFhO8cqrxTiVlwFuhHuc8un2E5ijMeI9ayaTxznh7xJ7HyP02UiLgi0cNfwWS
mTAAZDoblUo7DcbpJ2Lr9ygvOyb/R3O8JkVjnxIoyNaQp8idV3YtdsrVsPvXjtEfv5/d0RGJejSt
jepOBtn5x/ViPM2uVI+Cj2a43cdhaeVE2hLkony/5z6h/uHfdngupQ5XOX+F17aEpvPgQ4ve0Gv7
fZ9dniLABJfeUDqA8EC+3mlbuqJ+g+LCZlj9U3wfych0xLlZpMoZA/A9e/hv6hgBTEO+5MuPdH4q
IqPuF9wXYMmZRkii8qPr4tBaB0CuUB1l1PN2BFFyAReO8Tq9Wi0W0nErwClICcbQqK1AMHJJ2voH
+eIUp7kBa1ThpBSJsKBXrCM6Le6llpZM9ueOhRPqAT9KP2m16LTEOL7/yMAPfU8dMtQOU2p3epZF
07yaCAKzk46up6x1OnqZsLlDg8ImbF3tvyqLb50T6pb6QISS61eZ3l/W0Q8BTbMYbEGtPykNGrTc
gzqkE/xETn78QU9ICkl4OF2BYl6zzepuPv/m442KqC98CUwSZ3NsmUJz/k1SfPloF2igQqxgytHK
Ir5GwlHPPoGLNqdAEFDDn9miv3NuF4K3kio9TtnYGurlphz1OgSU6xmvBCOGYZpzg0x8teHSrH2P
p8km62qfg2A/3hEw+Ps8eBr/yzS2iK2HbCyQQcm+xztRHB4WtR168AFN8f46xwO7QGXnC9IXEo1l
utHz3Ev2oObukZ+NgObtHPINmhrKIJ+kUW7t/0fWOD+sXh7u4NE7H74ENzp+qFM1W4spZVdzys1a
Fu2OvGG3rZH79Zx8hKrqx8adPBHaNN6M0ZTmfqiBVHRjx+mztQM7mr/gRZIY0WOv3rvsbXj7t1w9
Eo0ztrLVHxYm86nazPMDgTDvhd9RlS87361/Cs4VQ3I8evQnwgj0agy9a9E/jAa5dklS25Xh/Joz
Tw18kW3ofuK4bf02S61jZT9UVZ8dW0v3AWZsLOKfdLOhoy5nwDUkq+w0SXT6WP8f0Prr2WwYA8zh
zX8uJecwbvcwxY48o/n1FkHTXYMGF0R6xceGVdmUcVoGqys6wern8oJDf+yRYLG1qTTHy2aj8FPr
d5ZKQJOX4/AYj0mygXCnaAW6cLuKxMz487sd9G7R2bgfytkeIS3N73DxfJGZSI40gFcLKfhRHZ8j
5HJKGgNM71ov98HDQ4A8ZilB2vjFDd+lm7wwensiSMsJtDdfe4+jQPu1/HMhpryIPnEhBBIriAEe
pTOnJPwVJ0LZj1PmY+Gihf1M3TDr5VOEEjsgmGkFOMGaYdBuOKUG3PgPmbAp6NNXzio6mpYK+Bvw
+hVUEZy0tzGeS0UHd6vLYDBn27wSlPsK9z6QZAtHGmPo+GAZ4WjHLsSkeEpjbA/uIyXd/UriGJvp
JgayP8dQebsxMS9TiH7tD/983a+PCmi34dhZfxhxdmNflSnDqMKu2QdRs+iD90muU8sRXJz3jHJy
N6LGkdItu11tD1IpLXQNyD0Wgpzlo+AM8m05jcVzl0XtRPCzWQSXiJ3vui52d5k0ZG3NZYOOsBst
A+Skq4rmN8qgb/Po64AQnd8zDldyJFVD4QxM1bqWqwXgI8KxaD+OfZEFCjd2YB25O0H8zg/5jlJg
ikuFvyuqMKZFv47y8QlinCbdo2D5XZ7qiNc/sW2RLqWai20p/l93WvMDAvx5Cgca0q1t49xRpds8
8daRafAOswZBJdckdr4OOZGICZjViuG8vtYzVxC82OSkTzkEQ2GtxRKjtVn0l+GwMEqEtFG/JaML
REEm5n3tBeQ2Tz5U+VgvJYxvnoFT2M1NfLCGi9LIG8N0IoiuEo+XJ4MxUGu5WHLQUSeO3aLmRaqq
obMz5CdZntCqyIc487zfw48C6+/gv+TKZUJ7UD6+EyrGN2Uiqz70lUeFA+GR4vPkTXVjyJeXOGPL
xSoLYbZyHLEykdD/42yrM363vYj3jW/cJU0YeE7jrKbtRKe/JT7pMWEZIQjdBuC4OHDep00bG9Zh
8HU83/SwSxKGjOvvuyPHKEytuOihN0TP+qDSQoR6yOpalkP/iQgW/M49uTWFUB3ZXps1AVlKvFyO
WOPTzhSP1hmKSV0Oahz2FV8h4NxXsB7b5+YFp0VYuOVA9nOQeQ63kXPUhWfJGNPT1l+FhpwOsTlQ
i0uIZgiRCiccxlE0vG9knDtm8k2MRaCMWLwctGgH6UBu4jSLnLxGy7jbbh0zGKCYoKJUCA0soYsY
ulF9egqLtGHvaoonp6uO9hs7H60zT2pNIfNoU0BT/l9SDK/1UK2k6xXeIJvvUcrmssHw43rtDWg7
7QTwn/3HWSXVqOk4zBeZhpz1qP5yh2rAJgOzxvG96n74h4QKzEG9/N6ASh8r/lrcJWKHHMC3cO7A
UYomgMukIQ/nbYtaS97h7/fqd/dfL/cuTf03t3YTDCd0wan+ynk/zsfQ1e8bdXOgYQbmC9qG8VEC
HdeQp8YVvzrq1SYVNtv7UOhwdseGw9v3a7xXvwVIPzdDJkmh5tYjK5thhE/7D1mXD/yEweLfLoVS
LZEBfR+yZ4SVKojQy5rf1+pdFndlrdOztiGx6y8a9RZ3XMjN+ZbRHwwWjvqiWdSXY+PGCS0h1s2K
Xml2on0C0AsUcIX/pi0SyjcnODKbhkhcytzBTlkQZQkDUSnvvwZiCnZfFNPawJaIsL1VZeL869lL
mHHsDdcP7CRgQp6sqEOuq4Jf6YiLW1yn8kKVdfJYS0FZTIQDqJTCimtK/bbTtPWPmjnM+rhBed2c
LsVhjPS3Y5Qgqk+cvtskPYhzseoxRNhUa2VhbEuYZPjQDUvVsi3gdNqUTxyWJ958OycuXZxIaq0F
xT0aq7ptArLotV6fG1V0HCj4N50ScMUkA3UGlEvM36SiQSCNhUQN+ObJFVdnQNSuxgI5cBPkvu1Q
GRvxwfLIhTEAHapJYHRIhBH7OGNM652Zt+SNj+x2QA8i/g/qn5SPJh6n4IM4k/ql/qy+h0NN0Lxm
EPqiISFi0t5hf9R72BXE6xWcM9LhFLTq6HD+MAl6PNBcfzlm4SKdgn3tNrxPeVGnRw/IBJFdDq/X
D8/q4057YuB6KzNTZFAGrEhldQJy3EJYG+IZ4pTnIzCgqmTgnqPCxR07c8daV12IiR2WdqEGw286
vf4ycugY9/6uWDyl4KAr5LXFXv/VfnaPvqPtbpYQQVqHggdxWOpaFGR7EI7NpGG76+QZKf7sFZfs
QCVfFnv6x8vNhMtWuvMQI+wK7aLnLlZyza483Bi/iKOXERhUWkHn5NpHOzxEnGM6Gn9P+d+8PUUg
aa2Tty83yY6PRMlim+5fJLFLac5jx9WV6oA2MRa1fOvQZKjHwEcqtCrFLiZeugcPGuVRnS7rfECg
4ecetqC/Nqy9t1wpgZqeOiCd1vhnhVmfuO9cM6DeA5Oe4sNuSC3qXzj38bklPJOspqlXoPOne3Ba
FEUfeNKHVw8ALs682b6Depgb/tpGUufKbl/2Pw3ljNT4c/r9Z8v61JU2qY1GfzM+khNJRq/TrOYS
7hoX92KBizmUGaW6SHuCnOyybpawzwsqYjhX36RJpS5HvoThyqmyAWQdZGh/gfd8IUlTgImPNluy
N81lYw+zjH+7DbkJ3h6LnF+i0s5/tVw3buQopNL+NyjFcUeXAG788El09UVd6YV0vAWJwSFzoN22
rSHLxUYUD5mePumAbeme/tCn3qTcjXE7/fKBQ67Pzt8GGR/kf7kF35/gaHaReEFkek1aiwcKzLSz
gY/e167qz523rvWr/FNE+OlVzpIvP1loNXln/Zjfe1/uiipvM33qZOvc0D+LfdP5u0tSaZAtKcZW
cz2iL8kfaW7djyifs43yy5uqQgntg3NMCkU9s+RL2xeM1GNK/ZRfzP8paCuKW/wlFRBAQSuqVkz1
FNPpBcoFQfZh3CgoAehB9nYTKGYFGwkvAeFawWTZPdJGVK+nGjkHp13rqscPPjk88j2sAcJ5AzVq
g9RnGL5TBGY86k4bwW7en+fAx6mi+H+mOrhihd+dkS2lTq/z52hCzH5VeF6cXn/6htgmddVgDtaH
Y4UAUvhhgzhXrBXIMESZBmMhb3S7aO9dC0Cs2AKL88/bIC0x1D3MiDNn9eimkiRSOfRFPYRPPM5U
DNaFKT9NyCXFQ+b9uOJ4w9q45Zhr4r9Zoe2g2py/ToRFhZ8spPgxyhxbehpdyC/gIPooZ/a8zksJ
0z/ZJJ5fsfsaNqQrINwvbBGwkmf3oa8PPU9t2oEHzK/sUzdzxz+WXTPD3vfSQaez4Tt/6QRtusVY
nrmPb2MXo3XRPciSR3PY27hU+THN7kW1LdZbXsPOL+581JmcY/HiSxZQyVuJGYxYMe5JKm+bsmMD
htPc8Ms0GjLj5yPQ/y5ezkpFEEQk89aXV3j1qTwVxiAZnHztBsCeTuUhEu+RmdfGOFBIYxs2SC+r
IFPN8aPsoCWWjK3rAuxPWXX/FgBGIG4NX3oKvSkGz6vytity3aJ7IC4fsXMlzHBtsu2hH2s240m0
NOPO6hV9DSFkSg4L+iIDwOq2bjWvUqJrNR+VWNzydZWLV1gRd9oBZPP/ICWR4e9mfPEQ0r4bTIiY
ab7mvyFX8mf1IdxYeq4lg08wQQ5LeQJMeSsCNKGgq7NeGnfuKKGumfaofzTD7LPGBGP1PNc6QPHX
ZIX7gu5GSiko4NnFykFA+cdg2T9OsIWaV7D90QmRMJ6D6dDtDwuPHhkbSHatheuYPGgI2yqktLIi
8Qf9Ad4zSKcY68Jts3+nAEo07ozalWWCNO0iGFDea2iX0C7dUkFxwOuAe2B4MdVeS0otpBMRBNej
31bwjZJBzqZbXq/DRD82gyM98B4/Gj6ngO/GjqwXzDPmmDJ6GbgieACxE337yg3IIe4GLwP1hM25
Bg2tyvSyiKp/Ik+s0dd6InpNWOxvqTu9HBGNF20g6GNf7g4hFZ85PVUHhhfzXstcG+uk3vgFv/g5
h7Qy34Bh6dZF2kNciS9Mwv4hNZp6QBhxN9yPX3PqKZC0pRvVI1vH+oy/p1+2F3g0zzFIZaESU3FJ
FpuM0Ec8psHIbR4vUX61P9K+ilFPdLNHHGh2lfKaWKm5bwtw8wzA6dtuO1XhO1ErGRUik93uYuYF
JDObxbbhlfY5s+H+WcfPTtkoPPCZaoyWqhYjuitq4td2Eb6Ug0omWXxL64/TJ1fX9xfaMReVBuZ1
nqmBXVrNtO/5HR2a51aRKZDXCiDSCtuBPMQ01zBgx1a1dUHqxmnUF1y1d8rqON+yV8vu7vWa4mfw
bEQED7T1NyMSZyrjTWr31VmRmEVmHMxLWGyRGb3S9t/k6phDwKz6fXU7KH0bunYmhZn4PZps9eVu
hrN7QZn3CgDpSjXPTBJqakMND2zANWK4ZAaDLfhdRYsCrFk35v1bNVAMtlfOG0cwx8e2cOUe9lM8
4PTc4rw7CWpDimxUSO8x8zZzBbjeRnD8RGh2542T/wIdi3anpuq5iJvzr9c5KpHAnejm+9KQOH4o
3YTxv2l9Wy9/4nZdh3gYv64T9Ob7cjomNPnHszGr5D7WuIw35ZL8oSjtCwJ/7EcFi67vmowppt2K
Pnz2moh/ds8+r7rGQa+aMt5Pia/FujQFFbdYuIpHMhkqZYitsSCH4v4Sjhr6da/a6MGm0fSZ7AuZ
YSIDAnBIiLTbV29a5w3WyU6aD3vHgqLRGZguocPWGLmz94/tGbNEOGss5MeehaQAB2GLhWzLTHjg
owaJYSEJuyql/jICBAutb5oWNa+61qWssa0PgSV+ugQmPUqQ5zxMIMVP6FhWRpN7j2T3tN22Q3YY
rVjh9uzcVi5cn3UOJXY/lo4hAHz/4wpmPTjPHxQfnAU8vtiwEbePdvwa9F+82jetZ2V+F3TALe+O
/9ptND4dAOI1vfSaylGanUr+TqeHZtoJuiI+Gn69EZMiOPeqpw7J3eiEg0TRKseD4pw9inMP0/SF
fr+PI+cKP2lSEGDqntdIiM3nwTehgobyyqOyBpFe09sF1na9vOj+aGqv2fdtvi2k7xK4YawOZmY/
l1aEpd4MxN45uN+vdKLxrFyInm/lXF1E5Ja/B+wG08WDfEJffwhPcK24xjaBXAHotIVlyJB5SGWg
7coMfh0nwP2C0u8Ceqmd00Nwa/l/O9kZzNtIrDsDJozZA+ZhIQSUHSgTMjji5BTwXT3Ixstghfv3
JMcNDeqtO7BYgFDFdTP5TPml9ryxl1oeCHGs59i6X+/pM/AUOHf8lU6ioBVgFPgVev2fLhgXa/DM
y6NGOlN2+iRqc+gLZkP5N//s7773ikF21aSAz88JCPLvkZjTAnxFyegGRg9arLXgbavQju7USmQn
8R/9wwl/zFlw3ezFgehaiiE1FRiHFFAkUsI7o+i4CE2hXOPMfXBmoadFugxVRpRW+PRBcaoOO3St
+MJGJCtONXi4PnOwJSMeC/bqbCf6+LmSUAP4Hq+vCaVVbl4mknGk7qOEdNCR2cV+B12zfKRpk/IQ
MNBVfSoVd1u1yqVp8pdnavbesIdWPdk04FLjZohIfKx2lyQtD3HZtyRTwnYms2NnRCwfezjKXdqC
47xg8qvuB9HPjXIwNKnpiwmw1768JxhCj41axVmigCzl26Iih9G3AkH3zGvLeoblIVtq5VYxukJU
ZWgPax2XLZqrJPwh0Vn9y07fVMhPIptI3kfaVDTpMnkivF/bQnXshCQqotj/RSfOlzbpla45pTRQ
veI+AsANrRviBWbq6zuPJv7K66jFgOYhcBk1odzI+bxT/NN570lfbO9ikktyBo0rn+WjRXSkTZcq
cxaYRpFUhTns6j3dOO0yE+HSmCnqegcG0GMJFZ4tIyeR0qlr9W5OcQIh3/aqzpGnR5eLWgz7wwRS
sHVR8i9RuezwIOP+XwA2DPkZXwxrxHc/jU7J90NWkmv0BsVeMYo4vAUk4zI5DO4TSIT2zBVZa8bX
o017/OUvBatgl/08lTQfWCcTLUKbx/f8lm/w+7wJ2FYsaKDOEWp1kRtO7Q2ccXaxEcgNRMmKN8La
QF41ho1m1dw5rxqzwQ2tDVZaNauUWZpFONb5wEkrq0e9ncsCy1xzVw3It5LUBnMQRI54UjGhoGFD
lR+fEztMIKUVcmd7nF2nQ+DADMV7PKrU2E3WRemG2+cd9wJ+4jPLhOD+LLk/n2n2lnicLq2yZI1m
/r1AujcAZ/X5sfuA8MxV+HaTGNQG7OiqIcQVSJftFVsUxDbE6gXNHVZVNnmFepf/UwRjr27gv+Fu
rZFAtThFEKx66r4dhO1/5M6NQ8yCUs4qMTmOfDPqpCdT//DkcBHtXeRyQn/pciZaSroSqh8qQMzr
uynIzcL3XmiGNLcM32f3fAU4aNG/H/fXOOgq3eIFvkORPXM47Dr4QsiP58tngMnXM4BL+uPjYqRz
75F797edeg2nQytPB6A2tSbVoc2wFHnOE0AuxoSxS+QMNsRhhDXLpLCoOo9RQG039U1DqbR4ys5u
EVMo3z0FCSVjivmdYv34BU/m10utaLMu01lpc0Q5Kht8t++sWIvKipNTdgu/GsN4+KJgXRUzlZb3
UccLo5lGWfABRfxLlaZ2iCIuGIShYlSORHmxb8YvrZsv5DJkWbx+PIBMofonOcn9xN9eZbcUjGL2
Em822GFTGaTJQFTjpVEF0K3HHcuHmYQl/LTKLt+r4pYVjQgxf/rp5KRalPU8q57R4Le44rrnBANI
8u9LzO9Njv62ciJWF49Nubp8u9bXj9pCsB5Fpo8J4AA5auOVNNQK3sUb+wf0L/bB+tJxA+FPoxBq
6GZ+SDWambMg898+rW08AxPK5kUb/CUt8zT3sqc0RS021vp09vJlKrLr5NAUQH5RN26wewqtk0+F
euPzR/+ac0XVhtNuzK0YraUzVfCMvcmkQA80pY6n8ckf9hUgBeXTUWjhUAoGHPzJL++o17oqIAd8
mOpLKLqMh2yNpNQ6ozkgRxjstDfFpIr9GI6CUBbfbPjtSFxrPkiAroCXKmKDTzk4NdU16cjbmtFL
xXnwz9jMJBm0yxj7p7VNSYR5qZd9MUbbEFfRaIzqdzwQXt/lAZopV25TOOfUBUuzi7Q8Iy/dWCab
qEyR8qLbBJZnKv4VYLUp2pUplpK76u2JlkzEeZ8e71yAL39GcP0mrh8nbzVUzoTpI48bMo2QPn25
tCS22fPIPXWI4apCiwv1e8NfRn6AMCQiMTVtBl+4NvoTywMsX3nJd14kBA4NJi+77dL8yXkZCPSb
cNMXX97egph1D0wj78FUyHEAEA5Jr49r+ciEhLQVxesPCclb9DaZAdEhM+1Fa4SJOPGzdmdu2DDl
k8sSVjUCCKStDYnDYKMsBQ6P7jzaOI9xXKEqHE91MPS79OAEVyzaZJa6Gd1/KSms8HpksfJV3tRZ
ghMZSm9+pXOpczShaScB/eGDZ0EiUOl5dG6TSqGNknfVsst49TO56UNCNn6vgfMBFxoktjcmEmff
SJhhDP6l2vs94g406GzuXshaBwzQCgHyoem1FoOfcsQQxTyNncjf3OYnYsIkNTGCfRZKmDEAZndO
X9RVpYpFZ6zQIBxbZmWBulgk8BzdKGpQsqIZXfhlAtMqf2oWvvo3oiHw1VqOrkvepS66Hc8VLqmt
frB4oG0JznaQxyj/jvJZjzD0ihyaPidJ8E0LUjLsl0wKXEj/b21tv2i2Y1UCcfQWWHVRCN3Im8rj
9/xdeIHpYfk8CxXoFidjLgzu6uQXZR5Uz4AbWay6PWs8NlJZ37/aVs6MSAD9Jh/GBye2XrzxYAPt
KXVu9wrZx3qRGP5WXvLAPHeS+0HYxxMo+9YchKovhqqwCqe94CuUdm4RtWHNhDeptjzQ1aeIjFRJ
97F6UimB/0S/YHbanxluWG87Gf3AzQbG70QwUYlVNZ3r7k5drWXrWB7HM728BwdDneddCU8NVB+7
yTiqArb7ro2xIZxo479OajFTJ3Fj4He6VzGxzAbjYURbVW0tx+kuFfOUFgHpl2mOth0e9lSQzWtw
y/bYA3dOkcfgORU7UgbW/Hj5xSsxtQA6QUNX+2pY4Roasc1X0EadEe90Mby0rickLImVfddFrh5T
TVXPfjyCSNA152Z25/olk8/XHv315koIzcQi5nb6NNOAnuGm8GGai7NrYXDCdOuSu1cHbxITNeAf
zQ6/537/e2WoWtjQFTnc70eTn2CwBGqswjuBFzK9y0EkI9jwe7tDyPjVlTT3me0grkHfRh0TDBf2
68StUlUHUV364/ZEZALV0QgT88kGS9/m/Ahe0xPKidQNfs/ZIXgOFXcJACICljPyuDFhJWVRNm5U
nHT+7Rk+CguDL/ftddqhFg2L+/VNo4MjQhY/T3ZWWP25N/VFh9t1W3Ve6QQMPi/AksDQ7SCylT0E
XV8eZj6QbDDyJj1PQHhzaQjv0ix59fFlh7+gc0bMTRrPmjviflJnUtGbln5QXhabMQUnT6NZpwVE
YmNEjtc/ArkD9TGqh9goqteGrotTZY66XRd7NjBC2uHgEzojooPsDm3NCDWQDPQDXab6c2MnzCTy
Dq718qDRYFsFnFdT6ypimYICqgpdpLhLbuKK3DaQWcpdw3jX9MoP72wyrLeRZ+ipG9dZLoCkUQN/
Ksiz82JPHVXAHghblF8UlM+4yLFUBq/Xs7w+t6XIxvGZ/CNhWqhMeD8PWGozZVDCB169a5NfrKD/
DUb7gj1eXQBvY/G/P0nmDCvnu05h2WIMQIcHg0L2SODJSYTtgJyoJ/RMVuHfR/zUC87ZrLBuC9/T
4dyvWfj7y9s/IbBh2r2GKF3Oy53Y4vLpBDQiB5HVBEI7VIoTPFW+6W2hPaIPfq9kOxd6j5q/4vN1
jSHtSkohsO0ekygpAZJOGIlcArQXBaNrl9zd0nzzXwfejZRWsdiDsEETM6KryHK4fGEduDPClivh
OUyJbTWwOHoN+QCiqSIUzFEg6bQWw/yoCHjPnUTDYrUc3cT7QOoZo9NPb37R/PK22oA3wpcchq8I
LPzGbnUOeXE98BGgT03PpyGi9WlvTyhRIA/MBSLriSU03plAmerUjqBQlrb/jmFkQrsgJB1AELsQ
xDnZl6TSURK02lw5/vZINMDZS5QQBIDNcrTaJv5n+X/dZTNmLXZfMKwQOw3mGchCUHaoHbSqvuaN
oPmPq9kLSaljoQwl+6EX4Zz9IMP5Ov7NF0+OGxGOpMnvkKGZIq/DPj8YpSH5DDp4Mx+p9no19OVn
ZXgth3If5sUP0RqvKS3WYN+E7DCPaPR+Oz8LIoyC6s2ztj7nOfAzYJ3XwMsI0iE/FBtVfqaDUk6V
TAxfRMFk1Ct1NjucHtPjNR29PYPpQjCkNDwmP7C2HNyIVf/EGltBsKFzysvYyoqmNSLm9tVwdapk
ciqLPtzlylEEwV2t8zVvTa6BYc0tcCZoP5u/QnZNrVO4BPIkqusWlvI75qK5HR3upHyjP8twwgwS
JW6NxFo3g0HSJnT25I0AT5re+ClJxI0WBSDEmiP7pAGU33j9DFGnBdMGqS5tJpRskjjffnX+Y4YW
Fxp6GwF8zcOeButMWi17GUlD+tozHWK57QE9pjaiBbslwFPugeU9jNsUyqa5PEBkp+grxhIUXiOa
AnCTQTRlCSMbOB1HSyD0sPefOziTvMkTy5hwcx+voKv4uJxv23z6+6QBY66FzvQYFIpsZW6Ch8iY
jjmQSih4eXCEb/sDHTQOxBDaKB7nxzYVgh4mqucUMC7u1AjChow+TpHm2unFUZFbwzLQCIqJouag
tpTRgaJzioDLI8yuApVcTBnUnohJzth6p26LO7prLlC68uyWzZT0/hhUcmopVGKmIquqGXQ54KN2
jvazjy8qUoK19AljujG7zNr0o6oQxM878l/MAKbyGTynBWJriW03WQostkgrzooMIVxtD9gNan40
V4Gy+2CU+/jJXKNLYgkvYumgLHaTr1hhsQj57TqDp542s7gIQI9tQXYXpUQ0UMFjh/rHms1hTm50
B8WtV/jtD7d6/1qfz5eOrvm4ILWi/+RU+/I/uzq3zEEOI5lQrbGLjFuKJqMLKwJtmPIOzydVb2xM
oYlPqmsiT0p/mg6+0lDEr9Ju/0kqx7F4GlQ8D11kx3TgPwga/qLxWk1DApLeG258GNIzkxvpMnWF
eOhZjNVFsQacjsKCFZGhrSrfFmMNj/ONaaMjr3ilC4bVGiQBM/ISixAY+mQShOljFUwTsWJH1hXG
cMAmk0OCYfWCM7SFkp07dZCv3XTruF9M1t7mNYJPCDQ6PUTdZuczOVnkS6I44Oq1C8ZAWXHxHxvh
l9IHnT5RXXYT0Y0c9A4y9MwJU2E4eT8eR+srxFx+bM7kBYofagsVpcPa5fcXVQqxMe4HtOCRa93n
y8gDKhaW4t4+6DaiH3JNhq4N3a3ZGvVNo6wyHgwoAMpOl8OhVDNqsWq9DruAPYLIOXLxNMBkQguc
kTBqenc70YMNotHIf6u/mYElDDM+BF+ZWqZ8r6yZyDm64I1EQzHXzZiNSI+i88h/uuiFmVpiYCrm
e29MhVqbitudl43jQnhkNKvq4KSDKOBGcW4Ve/goCyUbFkBJaAOZaGMU3S/9pEZjZ7uZSHQWNFAa
n60llRRle5eGOAbUrXxVBW/YFspdcf2W8e31IIQhXXJ0fB52iBhU2h2optvGifj+azfD4Z8d+RTg
/yiQ0l6W3RfJuuoTguJ5qVUPMbu4E83FdzLJDQQR73junasOBegGaBfl2+UuKekp+bPKtN/IU3s+
QliDm5RuBAFcCej0xLPN5nnOoI7lSdYGBc10aQf6CnDe8CvMQTmgOFC824qvpqj4+HaZKpC36Q9T
fadU7rix32XQaGrGaT98WMbSXw+lWbUloSvJuZ65Lp402DBZeMRAtGbqMIqB1iKQB3TQfCeHxN9U
USPcVrEXnb+/yF1HLqmCcX16IuXNs8FpYYcYl1rxr8xCLlNtO9+YtMDaPkQJ+3yuX1IIQDGhJD/X
7t/pbEvI8WC5OuwEHnSfceI+Ip5pIcvYq+fJ8izL4UWiGsUZCz250THQu3RmfZXynYMGTWXKgIxQ
5eHwZZFQ11U1OpTK295oRNoyNtrq5uRWFz07wrCOKPT+s0eT8zEtZbqIu6qlRpRIee2xxlww2Ajh
ZKQYYRm1hORsyqXv7utPNSwCQs7XPEQgIP1TdiwGfTSHoXt+g40vLx7qWf4yEd6MH+zxzueV5YAL
dXVo/wADVEQk2PpCuKjMta6NMRK6S0aAhpNWHaxfJ67j4tzrtoaLt1yj5n2XguRafqdjqoe4jqJ2
kRgJerC3T1jZwFQlro2Zb4ULssczyC+/ofx4syzfYltXb36mqkineynmzClR00ZUn2wdoGBhg92b
GaTYbj6x9bKycHujgdzxMJOf4T3jzxTNXx1IZr61cOKX2pX7ZAnWrc4P+212PghawQOQZzNDvCHF
XNK0ochySTztkWxAzgfAkpkmwKMR5vEFvjckfYRrjgZX1rXzokJMf/3nrSpbDyysWgVhydxB9hzW
yp3FyORXog6UlOt7mw0iXpM+eAMopx7kw3JRY86OuI+hxT+zwmndL8ahqll1kCLsdbT94HckmONm
vP8n232AHiFEdmz9HBjv/p6bO4Z08j6K+UFNRibe57pCvJR7Bh6JBzofDLYQpExk50hw82YxYwd5
LEa2p4j8ykGLHboiCPJ7UGGnKsm4ZAmdg7UpLp2nWmqg67b9mMuGcu8e2FcMzviflOoggbIB9VDd
4cRakFWNcdkJSC9po+jmb+MqmcIFqHxvjLPlhnHQz9bV9n98RLbNx9sLHM/QCtwaJ91iAf6EbfnJ
E+95ZmLMD9QPQEP7lmH8jJ/G5/PxU9Uh2ZXM/TMs16nftyAQIF+rdt9Qd8/XCPXhz/NwARFmsdnv
vMbRmycRZrEC8oT127240l7YjxuTUjMqctv8tBhlazhBX3UHxMbo4pk2GJ6Q19Zt5sqIzXR5Lo3c
YnPw8m5ygSILHvFFF9XuHVI3ZGCgXL6acCMNvw/D+k+4yJWjtO5OejH9UWU2o1xm9ErVHWRkBggJ
yjavWpOPGjshaU6wD2A14W5bJ0670vuZGUaHDOioSXXmrIiE6oxHH6fDFTpAxcUNVPx3gCKrwsH5
6i/aKsNTqf8bm+GIUB3cMNWKHto/u7/ATqhFmTM5IAU3itCfKZuPl2ThGyr1Y8POUj6uHDO/zesh
E9fo2rn0VNftdBmX/SfDaYqR27m1NdDn1dwfSwqOZcR7jVtDPgbLbczSRJorXD94X3EPoAO2F/wr
Y2x8mjgeRA58K9fp/fA7K2F6XcMdlbI5PzorZcWmIRJNDt+NlHt0U2Y3zpcAX6N5jCf4sqL9U5nn
FtRgapgePGIoyy1Q6XE3izm/VZyOQte3Fm2ygMtpejztzgHztDKTRbbJ0/+VZaOFViRAz5zaohI5
5509D+vE3+fW1NewstLxX5OtCqcNMBNtt6l2yOGwjWv17gwWXGIBXgqiB0hmdXR0KpjZrPK2s2gR
Vdbj+ykutjgowof2g1fzc46u4U9NcGSvbneqgMaBCNJVYvBPTOiZ8KQ33z5NVYUuiT4oIk8lBlCn
UH5kIgULv+YgVznBiFlxuZaH0Tmvi3P3ysOpb9C3A+w4is//nGbJe5Bp9Mwcvu6jovuCKcFD8Vp4
tseqVPbClK17JUGkH4LWW2tK2yf35jB2XSgfFDi5fN9ON/SNamtFwbvryTUm+qxRogZIsBxoLb3f
FuVUyIoNgtLvAYVbSjVCQV11zVu+YJ7YuTRXRMVvlgxdw3agNdWNp+RBOXf3xVOvQ9R6lSZs1HUw
DKqm122Wi2PVuvZ7ROskGDy93KDJo22D/SriMMYhvuV5OWf7Ts3m8eWVgZD1EbwDez4/RxrG6U98
2UL2w12lCFwJ1yGK1dot801g1J7lbYDcAK4ITuyLcgDBmZLvZuva0kcqmeIwbFwNxXb88hKgZd7P
iVcuhQTPDkbrc/z9gnha9KLQEJr8OswlBh6WTEf3M33byXliYgZlbm3cne6N0LCSiB1SAjB5hQ6K
GQ5fbAr0f0EIblxLcdA6k1z9Ym6KIPZ4pYnSXpTiZ/MM6dLs+461MQo3/oBsiFLxuKaco2RUMbcY
FiHAmncv04p4/G7XbNlrI/h936AQXvf3oW5n7YwsvHLCXCGoK1Hn1v4OmptDpZJyWPm0dx5icz0W
yEetfIshu0wtEvG/1oIHuJLKcRjG7cXdW78YeZGEYZfpnyGxelytJMsoa+Hskemenuq5wMR6YPIo
XjIYi8T6ld9spozEk3MHnmcJaxnM0ybhGCXZ+39n9cr38tUyWfRkhcp2DfVxuuS7FmdiJJ+JigiD
cQCxb08Nsf8IBNMY2zqAbT4f6dbMwMiQoIF7YjtPtE2KIEW25DAXc7VBQI7nH6j4m3ePCklBUs7H
3kdA3xti5miaTIJXN5K7SBFs5CSuFPVl7X8kQjXerOmuViSNBf/3wNzUV69sURBSEqdGB2Li0of4
Xwg2aA1nNX5VOcb19/pv0PLXZHk1SIo7EG2k5qqfRbs1f9XvQfIW9oF+J6z/rUNYfQBBHb9LZCTC
Kr0LlwVT4XWmrkvnK3ayMIt/Hyh0LXd9v+bbEpTS7bK+nXHxlP4l8RAbQ2A8cqhPTKph78Spz9kY
ECzoItUuvW5SeLEoVWeCzwsMSSgzvOql6OKFqho1bpAyWu97ZcaydfXOjQfpJdLMEbMETb65e75o
SkjliMwy1okTRrGyHQlgNrbPC/NT5YKRFEPM5YJRwrq2pv9X0KnbexiD7y7fUb8eRO20bl4w03UI
vKQHUIRt9EJNA00XYqrn6KErV1q3bgz8vvTbc3OeG3qfNMHa7jMfKeC2LeHAlx3/3Tvo1+asCJUU
bOI2j1wqVVRzBbFTaEiT7wH6YRLyxkh3f/4tz0kaSbo21gsNZzq2GPHBKD1tnW/Z7Io+6YemR0yc
o+NkszpWjUTSGh+GmxpDqd8NAi9uNZMJmaOzmtUS69uUN/1r992myDI/4pIwLTaJaezZP7c314XJ
nbN8l4vBmU7H3zl2mo3qHRQ9bLEXHHPLe3DiXGuuLlcFeqpdX78d8s28oDBWxWgIR2ntJ4Km5wK0
nKVajl9Ama970H090vdPGzZdV1jZT8V5r6SPSgHVbDHRfeMJQqWD+ZhYJ1CROY1/Z7yTUqJLi7dX
2DnSPHCeUloBCeINPz8PM+qTrrrgTAvNJT8OTP1ZqfQ+rroUW0kaKiANbywqEcS9gOUnqiNzbkNN
PYSkpmydKgYFSBSP3wr1KrL+MaBrXhyH04eLDjGU6V/8skFsIlkjEBf0dGK7lHj5t8OybEcJ17OU
BpGMWnovdHPiPix0qo+uAQ1EHnajE5ioxHO5c+m7QlJ9RpJ0sF1fJ8GVuxoB5QWgsW/uxDNPdVQE
SOUZ+19nq8lRlwh49XFTO0aqpBL40OLVLLK/J5XGPyHfRpAzTb+llax+joL6m6nGlS9ni3D459s4
0p/wz8IWytI3pl0mhDB8upCQOwcjLRGeWodNjlMdvE1rXQ1WpsbSkj9233zBdnBAjjh9OGkH/4E/
dkNhal/Qs/y1BZc2bCWOBxvP87UEj4QYJwdna34Xv8ysQOKIB5s1DbkrT6OR89yA294VRIwwVlym
yv0aWZU307qVJXbsiq+vmfWOZJdEEt1bTiQR4ByONapNgtqmzTojcZOBV2tSCnXTWyh5hJHngl9c
D2oKlB1draeHDFEAwhj4y7i/698A4nzF4uR0RBDF55jHVolgpAFKT+cNGWd7qN8XQ0MEP7/WYOQo
bQGVojts6K8fquvQqaZEuCcx6xjl1aeZDZpkeas8QxrnlWLdlwpjZ2FouqafLlBmYFiZEhSfMC5M
CxEqDzXpH9XvJT6NdWXiQDdVkFQvbyEBgLCA0tTQfSzx/cOYTGa/5gGbxyAj9+GWGbHDxq9D+tQ3
Er73g27IYz1KISQX4W2CigUpqJc03tpCO43wwZw4AQ1M/75kk8PvoBCT5tp7aC/CeGeEWFlXBLjM
kG6d364GCh2szCZ3qOG1bs+X9a3PDgApjYKWxv2Ksu2avmSCTRb4svBB6RxALr2cEthJBQr1Pz5y
+AjJaZisc1VRcgyfCehixloH/QIPsUd3vpzZv9KAAvNJok2cjzqPb5bF0omWHsysACjB8rMrZAIP
rM66zPgfronfke9zEN6mQhRx0z8RbcdM96BD0r6BGIu8HWv0hrcQR+OwdcU/WQtHDd0dc1Zle4aV
KBPXMUNw0RnhVbwAatgJBzGkef/s9nt0+Xt4zlGwlQWVqG3lAFv0Pheeles3kPLsOC59/nhJZn7M
rsZwts4zZXj31lr67mxSZbmmawFE+FFD4UxNffp05KuO17erO5taYZkQ5fwVcYHXLpgKy4gIWFoG
jcngQJWaFFIJRZsY+Rr2eHjlhbsEOP6ywCAIQQ+peSbtelZls0szJpGOpzoAXRu9IK2nwkDVAWrL
eBa1GO3XeP88v8Icuv3LmWNLnHpeLDzM6WV5YnAtadWP3ne8g2UI8/39l9smPt2zsvqV0/cAYaFK
MUTNxvxWt3CIm0kY+6jfBkaDTYAOYLJ5BQ0EPTK0AhTKfsLgun5u5DYPcfBZJ+Vl6D6dORo8vmck
v1Pq/UrySpjQL6lBzxyRz0/2lsjUAj7CqONiTZElXWjrQKuzk7Aondh1o0DLDnclkivDwCfbhH+z
J+TV/1ZvQZR3ifbLD1vmFZKwGDxvDjG70tR++qNlm4VMTjDt0UoT9x7kMqc/bXnKKkQrpqH1Avth
/CwTned3jZr+MKEB3Od70W3N5QDRdTnplIdWZ1TPW0qvmkLEj2cEvc0Ly4+lML/vcc7RHFd6/DXk
RVQOUc9XMniudVyYDGdOM2+SR8Upu/tLDK8iSCGoWPlxLLnpST4inNoBB07xKT5T1EG1MpSfibhd
MErCBCgbznVJafe4YQvVJyODrZjX3AzSTTimmYGStlU4a5glWZabZDBnq97h/skDSDuM3UcnNM48
z7vjwFmP5/dsb0+Ohk+Yf8TyuSxF6UYEnRMOy5er15IY1azOyG55HK23PPS1d6nd7Q88OxXotrRN
lvmqTP7K9zFtXTx8wQNJvuMyIp2/vQJ+wfQaeU/0Y5hb530SGI0VKrRlQokrnAKL/rXs1jn+bes5
vXCczfcsCk3xXCwx2aIXV8kP8ZRXyPFthrLUlPadNnwN9vngRZf++UB2pQXBeRvl+jn8D6i2HSLf
pN3794ESucX08FSOqNP1oxQfLQIM1p/Iml529h6QWMDy+rN4LskW6YBSX4E1xCowtG3DMpGHDfjs
uyRRTJuj+ftxw0jZBHRGW0YCf0Cp09dlsq+Ys6T9BDXq4KrObhazbmconH+Y/xgQ5pmKSj16tASe
/22EMmAplcepTZdssoycGuhD0BZ6l1pl7kzDhyk2AY9/P7aqZQ/TtBduMfKKy6/yccbyeSEGZgTm
9xVh3PLdsMi1nRCUFTxCuokfzKilw8CB3x+YITz85vZS8V0INYn0
`protect end_protected

