

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Z1qTni396T8iV2R8fY9HyG8eslMc+IRW3v+hG8xZdQngNe97GclFhsyPupWq+OKGifq0gIWSbSAq
GKczz5JUQw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ngr2Ns4J4TLYxu5Rb9qxmsaC8oZ5i3v7hFzsbUIWxuc/aGCvN+Ig/e3uzREfWM8l0yT5FJX+JwGa
/joX07r8LM+k1WExdIkIwR9Y8LNxnjKgDveQQRBJUr1FrgWZ3kJ1Nku2y/eaPhxKCkHdbspLfiK2
nLMtx19dp/OxU/pUkUk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mEajCWc2cVvt5aBBTN9qxYj8nmXGU+b5aY/Z+76lvXGCoafJOiBEPfYD3+/UzJKCAYd5FMV82u+5
N3yfi/qdQI2t9r7HHmAMuzMDltJntkmky7IfphJQelHxjIq4B0pjCmio+KZQIBxCV2L1LA7hRa29
P4ikRuu1b/eDcDvNSkwkq5fdFSGckN5mgz43nZhFhfDRRi+v8o6cqHF079JovOvt650pyJG66qqM
a856O4k0HRRWDzmx8T193c5BjoB4U1z8H2NEXTAeWKX+NtJ2bDE4v9N5ib4fPXCNpwF5Kn1VegR/
h2eSUe2DQ61M/5edHexnZIr/lH4YNJMogqf/dg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LfEe0E/llANgtXATlcZvjMcXUNf+JJY+bvJJrPEoE34UzOFvrxs8XP5WPZSL9vNSuh2Qg6+dogs5
y1CIIXPnBhLvQ9b8uwHUoKrachLXExKd/D5qFxOjEylTsCK7ISyXq73hba2Nh21EeK87oUnERcUp
mEWPrFdonIVran5dCLM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LvkSLaIkI75VgfPL+LOvkb1M22AiFuawpUO8wCZL9l532TC84ZzoNgZO+q0zTkNQIRrl+7yw3FRI
c4NtSBUPkKSfKGLxYkg0ccBK5Zav6jgGKll6nl9OOPf8j/cPnHDmRp6Y4dOMOdA+5FvZW0UFAn5y
T3v9dq4JHzmLj9JlxEGY+tMETWuXJrNlexAhelXM85DfExSN5xMPGWmgiO0AEPOg4F37LiuVeSDd
V3OTTxiCje5lsh9lR0QLRrLntnqiyJKQKRoh0faT0lMkQYWb/637Khxp0XKjIoWVxB3PFA50OJi5
19t5V2hahLXTaMBOr4n4ehdVX2WKCSqwQfVmnA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5680)
`protect data_block
MBzfJJd4GdF1KIeiPJ2xYM1c6KIOWNnc+Mnth3gyBP0E422LM2+vAKMVRQUwu1dF0T+Xa9UmChO1
7I6m+zH7bZtFHp0ssrqOEE7wSDJO2bEczkCma0cO99Dwf3z8acxJ7IE+WfKVX5PJb0Fq4K4UJjpP
mSSuaOxyOkD/bttyw9rF10e86IhgF5GFGFJTYzu+dR7HCXEv2xvHcRynt0sNq5YiIC2h8Vtk4Ubs
wbYo2X4T1eOsPkylxxBZ9ejkTPtYXo5NmHMvbGgmXGxzl7/E44kcSg7EcsqRTfMCAcenqxXxs5+n
R3gtytDIU/10IL2anBFOKaPkzyd+snCycdp5c7+gBGuf7tuON0BdNI+H5CgWaW07KoEubxN505aY
7lBeH8I9Hg4NjxKs0qAC3FFKxkiYmsauSetKmysX7qgJomz7StHDBEbh9VGXDPaoQI1S7Boxin7c
JWkWLl+hyp2b1fluoncKsqm8EXHYJk47gZIunkG1gqFQQw4NgL/Io9O22qJX2EEkqVTY+P0us6sj
kB1Kh4pwpwqM1c+z0vlJcarsdqTNfjr19wg27yoYKlpNj1PMUwuly2Fii7ag4zxfmwRTdP2Brft2
toZ5v7Inipw6+qfPJ8qnYw/+p8bl/QaNpM2qBKH3Vc2UdAIRr7gpRE4eVgL6w3BzHjjJfWp/CV//
nMZQpL2yXxJrOyP7qwMsaTmCVaD62A+Krhyit3k7TfjtIsijKpsAhiaWGXoUZU37X3/w6I/QXm1C
wKnjmTuaAHQxgxjP/mz1OEIIu0QsxYg0JOWisk30yzg9MHG2xF3jalCqpekasUkLpH011sB8KniM
NDEYxLaEyxKl5DyV4p8OKEnbXoRryMoLQQ5d3dF1xcm+p4kNzwNTod8EGCZyugtvGXIvK7jCVGGo
2Qjb2P+42GQTuYQe3KnSWbaDTTF1KRJZay/vJcOY60ZbT/MfqHldupKcJQZfE8Ou56LUqqc6K7/E
yBOI3p5hbT8kKaGbKhVmqrPS9w9CU4HR/nUnkDvT/2RqfR8/IiijbPAngGEkbqgE1vXu76XbptdE
6lvmlQAB8FBj2ISH3qnavjXBHrAgfi4RYEf63S6df8WjoKj2coph7oQ52nhjwMReTfwWdFxPmReb
AQ3xzCce+OGopOdZmGfKtgyCrTPt8X0HAVHnuk/xyM/4BtDeV9N3yQJgQ4EOxDkMRSmwCS2VClri
IA00rer0Br99oE5NySiu+MNuIpBb+7WbUCL0V2FcbeQ10laWFImhKOY8ytmXdySt9pDGkdz42TkC
IgUaDiC7f2b6ouWzTdPE1jENQ/frlXO5NAw2rkRsXSivIKsyknOgV4TBzYlqWKUMbf2Huq37UEaZ
2ieiaZa4Y348rhFAQKMXc7O0JipDJalB1RwHLCuWwHCgs9V8DkFW/pKLSIyzpYavm4Mzzxv0Gose
ZxDnEQMVOjuQRvBSiUkXWgB+j5W3DZJXT4nfRFCj/rnLk8rimacj41YrE8RoDa2MX7Mw66H8SKWg
Y/Gt8OuFSxOxjlSunqmsICqL0TRy9zH2ytrj2A+UhmTodPoiwGMnEdlZnrdzFQtTYGlZIuh4h88P
+pbB0+POUCmG48ugI0QNmOfvz/9t8vx5WGhsLhRWVStDGZSAtLOzp0wqQvYvK9zcRsvwtF2FJVzh
0K0W2LmuBjy8BlFmY8EIf1az46MA16HA/bZErZ9xeXFGLU3FU4dDUGo2m+o4ZLzpsAfCQkjNQDQj
4gKfqxxD91KF6SdAEX21MFQXNX2bOAfRx9EF3v9ZHG/gKUwO+cWO+jGhPiKEf/L2Zr93A6+yxwsg
pD2PyRxQJgzpJZrKt5p99lomJZzkjQzs3s1UNBUNzzmVrerY07WT1rLnMNAf01s4+XoQe13ch5G/
wPF+p0gL/gGR77TNJtARKYHULhekv4jnSnkp/NjHg3QrDhO8F7Hy+pM2AgdSkWs20jAnBMUgYOXV
tlBH29c1wXCtmTh0p1eEz7BxdhkL5iKpH46QZiPoBLrI58SGjZoVEx2kqFEy0FFW1SxNdvCB7QzA
BsPIXPCiMXgpCRMMt1evJYeAJ4z74oPkflTfLL2VY7dX7MW+6fhwGCOPJzpRLAASD52XvirY0dVB
f9ikOPdKpQNHdFG2gajN5c14JI6acnsYYHBdYjuko7LkPUx69XLXomD4PncqMilb5WRsceyeZ4b7
FG1AVTpHi6+PoPktf6bcuQn1fgXlx0AMhDFgrW/pl31s2wbN13rgYYsIBvkIdizfr2wE5x8MWydW
TkHqcaYpcuyZqq8BIEE9NtFOS2gC9LdPUEoWb07AvSYqGSmr4ImEBxFuxV8+bIBiosVlvMQqnya4
XerEJzj/+7Jsl2Gf/E3mxcL2kgc16GzWU2/Cn07sV2Ak6tM9QAZHQudhfWKJSWyvxd/oWh/HU5as
r6S5hmldrN366mDtn3W7/H+tYMdw/vA65ibpQRdvfCsMQSYS6/GE5ZrvFYpf7Qn2IKSnEolctki1
ZKgMVh08ytx8xO2UBybrNs8hhonJUe0cW1WTdiu8q5LYeZUcX5QSeMC9jdlNKOyuQQyhjJVDbY9j
e3fJrRA2fisZYKvLJHcr7hrwJg4XwZdW/lvToiKifR8XSh8zvACzCeMtbknhw8Shbb7748I631Vj
9pzzAwVird43aTzqiiKiz1ufCgclTFhkj93ZQMoOEoBYZpblUbJex3n34vPVy6gUwAB19zjQmKTi
mW/Nv+B/w4SpjcBbNPiOxMrJTr7wQS2X344KoERDx7lsXW58novVajQMFTuqI0kcZWFJ+K8dalC0
2X84DDFEBYeni5eERI9Hseh6lnjZMJCCG+b9FzfB6n4l9xsh0zqaHnGM3PytBPRcAOeiLGtTNm5i
usfETkxaYTYErifCVGVeWJw2bIzUZQ6Tf7dmMIX/kLCTVVue+5wwf/lt75C3TNJVI1vCgT3rpl4m
1Hf4Bpxqwv6YO9xglZBxgrNEiNV5GDNQTnsFP2DTKtGiPTgsbXED5ghKniJ2Y+wjN3G05/S1dySr
zlpgji+ENMCWxarD3R29dbrDDPWG8twHe38ZKlPqF11gt5yrtdekpmpHVwP4GQuFYruCxHEnDANl
ay5LgIcoIShXlqMgVCMm4+RaA8tk9+SS/Ix7Q/GePIkDV4OQUo4YF54MmLG9T1fK307DVIGah/Et
70NZYdRavt49uKwLU7P9ZLJSJDJTRJERkebzoEYEjvWaZJq+sAq4Dlqan3hG62q1QwGq0DGmPOff
M3yc2CUd1i1IBi6Hi6dfTpYcbF+LTv0bUZKnPUdSPAlrxJv4th5qsc3CK0dWVBW98uwcV2zI0GvI
2F9ORC9QVTT/rADxbTe4aHbBfOiPSvrN0kA35cJV1OL21XzFWpdvK3/G2QKHPQNDErsDgbnu78mm
/ep8MjbeRe0vaSxuYfIgDwGkFTR1omintuWfva4ggYgT02kE9f7m1oZvt2ohcFd5MP4kfd+KxbqI
cDpp1oiRCOH0tTx+TNfXkFDBgOvvrHLftfDrg84rlDOgyWtDjtTNYif+CnaXJEM9vA1CgeTVrLPI
hS+Wz9vB6a8H8qIXM2iGD5+kLRqEbe5UtyRL9gfYSn0YsHHDM2xLqdmcApoLw0ylsjsvry+C+kjX
0hrHhPFCOEaCqU8Qltix1H2iZ2PPIA2nGsoSF9PgCawdt8HSoERrtUz8/T9qq0wP3bNXDQpflrrC
+poSqtSQFc6UlCFXcQPB0wLf1bGI2gc9hfgubJ0MlPePdyYCN1w3lDXJqIj36Du9MUSw8C6HRKup
+nbInl6lLMTOkwjlln9Fwm13Nf5G+GBOIKEDD8inaoWQMouBy3a3wBL/nJaNYzrKDx13nva8cn+6
547GvLJGPf3E6N4220yctepRx8wiEfL4URWD67LZrtZE1H8sbE/VZaXq27p2lLsqBiway96WBe7y
JA7UVAKr75FFMNe1WRWDEvBr56BPAysP4Iqw6gSkBj4mR3M7TkQLSVqYwJhCUihg44GCz8T02izC
MVx+PNndKc3IMmAdiKVXHXow9rHiA5XPxKvL52cQbGdsHmG7paSWoysuMup3VZTKTuJNbBjRw0Be
BIp2L/koo1upnnoP+OHkHl5iiONQiHMzmiAcQgm4cEeoG3V7q8eBRq8ZU7AJLycEMx0vVfa6Uq6L
Ti6/8fTd9pytVGWlkxL0Rw7SDI6pNDsfgSqX+iwgd66MzJDx4FYno1c9q5FtOFVy4lR7d+ZX/eNS
97KDLxJgEBmB0oVE+WsC3fxLAAjPeGtMaVvKww1bJVb5CkVZq9NJ3KCUlyFEWKwiV6CmsLsdhupy
ZTr2ffczZy7pOj/NKoH9QocYczEthuT1DlbQC3sCJQi2TyzozxKr3jnM+jsp7AhicGZlYg4kJlqy
0VYrCiA7rMg7VAyjpOiq/JIMCH/950UcM+M9Ymy0cmzkj7a0GYraXzadT2f0zWdKwD59EV4n+Ik5
8hDr96T4hi4B4/pYDi1tw0mcEzLZ6aK3Rj0x2egxSL5aWXxknshx4qtajySPshzTqt0/EPk5bVMx
cGUTWuL5XV2X7l73t6SeDaAi+cmXfCtTUAEWY+pCUD+0gWFkU/jGz3h55YDBhxhLSAdUCnqQEEVL
M1wYMnT7JBk2QpiJSVangAIi3cZBZmxc1V+bWTWN7kEYRG+MkX1afUN6bQ6A+/rBRtMRkDI1yvbk
Besy9EMLIPEZFHJgYU7xN9W32DbQ9hhJXC+g1ZiCThyY+zl1B0jbl8nR0WY6LiHeNi9Jwg8Nr/vt
s9r6DX7Ji90qMv9NiAdSuM0We1674y07Y5mKDTKgDTZkWzaCjzEGiUXeBwba+FvV5DnshW11altB
UFEEWTYbeFKswzT1gUHCuvT3Smslc+djgKay/9MuVqXf4CrnfKuqT7cUS+mxN3DhIFcfpy8xg3mH
yo1DkhxXqtvoAnaGYu39GlouChzx3jSgbMrDsXJkao8E5r/HcS6xw3kHDBFP2UpFuCfV0YyG6pSZ
W7zUQT++AtaZ5Z8pZmZteZ0tZOXXt3jrCZAFcZPisGjwKJ6/XB5nT2o/DtUVBibwDTPV4LWRTrRv
SQUGs28+8O57z08SoQ+/52Yl+1W/+QlEWb2XyrjHZ5roarnvY0jtsUf715W3/SaFdk9jKdGtWj3e
XynrGITgKS5BmQrer/NdMMAOxclZJJnD5RHLgeWhtf0UgzeHIH44YgXa33AFUbLjR9A3AdqRUcwN
I53fQSvveoqsRVBFSUKz/wD1gfzHZn+4hS9YDWdd6pOobMSjEAmoRxJUFn0I5gAnk0uNAn1QwxA/
tpIacQJKQwsYQvIK/RV6080lr/FKwof5LnSxGVhfvpbvzhdibo1XFV0TyEw4Zp56fWQH+Wv8qwJj
3+i970F8Ie7nnntKXWqdpkSYKFAv9JFvaAhDScjxXIH5OWDRwSYSVLMJ+jf6/adnBanB+ARkHq81
UaSTUn9Cvx+V9BMYvWwz2LdvDNStoe9hLVV94NUX4EZ318D+5fQzdv0WkYnL2XanJ7YMOtUsY4Vz
QXOXqmL3HpCLWr8Jb2LscdrC3/DU1O6MOqeh4fK/qACliB+PscW9YwZuuAA011+RJH8aWL/5whwP
41ayBppv/Ii9fpoqQWQl4HbAegIk5Iz9REaeJY2YUi1gkjAFl1K/XPp9F4KjYOvkcItl12g5QMyf
J6r5mltD+tMl+TdE/yhNNHRd/t2x1vntsn47wiXPJc+E6arEW4VJuFpsSC0FveBx3GAfaYiK7A6j
Uyou6ohTtGlMmLDCaTehheVBnx/SIQn6j4Tg5WYsPWtN55f70sIwIImarVfa4fhTCt6ORg26oQFW
4tk0Ky5Hk8G7PjXZDgh+08g3eHLCAs1cgXY9sGwRl/hhpKDPQMRVFIaW57Pq+fnaB5kiJYSB4O3+
CXDJhrnIwq7Bd2FXFe9V0AppNi1L27TUlSXo93LQviepn7UCvHWTBIJqXMqWFmTkAfcYQxNporD5
Tyd5AO70xIRAvCZri+cwmxW5XZOxkeRsB9F8/Ki521SE0UDdlv6kN9D3GJcpMMZT5V7NrJ356eyz
7abvY7BY+KyafHCJOrt7NUgwqEJJN9EzcHOrT9PbyCNwYp1WQelCiPvYeKyXvO+nAcPB+Faua5sS
EDEwonfQ9f9XuyI2CSMeXrWz2Njc+ufxQucquy6l9ZPNDFPqVS48Y4uqu4s7PdiCd/aJ+b07KfYM
6YmfKvtvey6mK69/XwEc0t1dGhZd5jvH+oFhn3lDclca2zjW88gtXIk40jd9vgLCvBMTh61gLBO+
GHxEY61xBrjllesrYRnTQ1K/1K0wzRpRcv3hzyX/F20qU8KlyhCDoa/usJBJcu62HsCj09CGdmJx
FYUiVyRvrJxJTm/WUAyeRZb5l8f1SMVDGTLxs7jyxXdCZ1Vs+WZqn1lBsb/M6xndESNUuzBwBZHB
XukIDswE/o+t4WSqVtOONn3+gQlRmTmNdI6MuX0XmKN4K5Ag/wYvKo0Hy3TJ1N7oGOIdoto/dbML
QyyCS+ix3ji3O2yXDOi7oIMJLqMyhTbDA31ztnbrWMFifVEU2Hpt5KRly9depU0cO17kimc5MJ68
m7k13E7WpaNR4UrEd2G9OXRVCa8zCBjM+/LGi5gmfKZXpmV6HInEYpvH/DwP6ZC4YiiMkbXh+a3a
xMXy3FQ0XMGoP1vvZNV3WfMBHrE6BVRFj9p1bDNvkLT4Z+sKM04Ay2PotEtzKpw3M4w3H1UIkl6C
uSttD1PRDlGupIKqBFIm7oFle6q1mkuqNzhgNdg3RewEWHhDezcHGJC1HD7R/Q2chXKJHwSd7H/4
VWt1svmam8lNWh3rJGiVOkk3vcwNGmg8lJ4867BGzkXvrsALeYq7bEE1/nqEhX3wY0GRcCnOO97a
RALqhVplPRwk0T1sHU9UY6xgZMSD3kzFDTYTDgx/4hW9ZHcEiPfVq10LWyzSze0uwN2jxWytvqg7
kjeVv9H0NkVJu0TfIwON/u96uFWCjLtpk3RNEtgmNYUjeCAa+cMFOlwUNLHqAV5B+Au06yk+W1m7
7XVv8CnLmRBTUxPOezDLeORcb5LjmEPs1Gebn8M8Pf4gtbrEyJBnN7B83spaGu5KYcma6uedADRD
aksLfs/plHsuJ3wUeHVKaOjYZZyurnNsMsfXM8mGlh1mZWE4ZBPo8AS3jCOWbBLOc+yfHzbguA5u
RPSFKVHoFyjSWfQybxkYH0D0RVN2eOUslyRWHaXead7VP+zBNfw9/rozo3HCM4b0Zps5iUgvkq9Q
2Ia5OysD2KvtfdxVfJQeeh3ZLLghWYGfYL+3DMTiU+nNwB0A9X6s1N2Tal9g5hX1rvtnhaLAEMBt
YBTu4B6BgdQvKHVHQw5N5T6Vm4R+1Ccso0MkUq2SVlvC3tXjJOqISZtVQNUCbJxIt3A4ZbqG0F13
l1hPg5I+paJCB+NmXw/9YXeVwZDf2GgN57IKt3F75v2VF8OAgCG+nUvR+3rXjxGahUKlWJiE28AK
Gg3DiYbYXZvZSD6TWJJP5uVzx1Qeubdxt075xXue/vYJRyA3fg==
`protect end_protected

