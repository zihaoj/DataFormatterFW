

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
W8f/qc2qrdavIx2U7Mhf3ZSFqORNFIP5j8w/AHOpvXDOUEHtEkxRIZCo9fi2oSi7xMRTI2kXsIbh
aFj8siJGnw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HkyDRyLCEu6STzQL4sJSASr34nv9eU9yqQ2V6W1dCGzZcG1+J/umLTz59veK9/MRw4g7sf0NyuB5
W0D188aR3UTqFQ7qrfBtR4ILaoiI2GYfTD8ZGeOhZPNv3xcKpT+5+GW1egVKTx7y3PbZU317NsOt
ZEGbZavff2ZnuQKhqlQ=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gRUr7OvnT6/ETrGLEWwcf5wmsEf2Hi4Qsi8ViX+WIOih1N3byHevDD+l54lIquIxFvymZjqPZ4ex
RhJ3q8MIh6derf+RDcebP9t9+xTBCh5rJNV/zOnRx1P9HIBrKubnv27FFodu167e09Xq+2BO5J+n
qu5SguWy+TRFTGD9L68P1PyFVRTuDaEed0fFBH7iChokNJUAXjZrtWI+rJv+CRd172EIzqTjGGji
aJzDpmEspVIBzU3gF1hYBdOTOpJFzR8u00CaK49gFeCJMAggxl21tE//ag8lLD5VHefOYnj1G6Do
0E1TiHzu/dAVyVkDQqngoWbnP1J+kkugH/k7IA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MxTBRI1frfMrKbgZLNsMzglLMo3Ubdq+IiX/2EM9v325LeeqJwxr32xeS3wgmRx+RgTVWWZ+SoT1
Cyc5oRPSt57ODiIlmJb2I97Qoo0d7stWC/JZHFqmwjvhOmbx6VYbXxRZl5KpiSgfsyyQ1WsNM+EH
7WcSrwHI0AdSAFUzIpI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HdJS5G91Q5B0eQs+h7uQyUlVxMqclStqMea8nYyQeWpamRkqC2eurlPAQyNWxj2PQk2sUV7HaMr/
POCdGYsWGXUvf5tnGeaydaiQp3ylhCKanOHW8kA8sj5n/n9vhFy7BdbWbFqlGTsNs9ZxWWQzZdDv
ljKSPaxFWtihDHRbA0Q+XeuWSlgXGzyEOLtL4L+PJWRYYRScpMiGSET9PzewaztTDsjlJfMbCDth
LeOWlOwLC+7f3gCeJExbobuYPzSdAjdeZINszxPHPoa7FcLgQ2TUwTvDDRqrx1o8XpAnX/TaKD+a
5i3mF/BDg5iCfywPaW7/PgqN5mDptLpuGf7qUQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4256)
`protect data_block
SW77mkOHY1/dqMmyVJpYRshK8DC1z7tjiKD3vga1ANT2mLl6ncwHQp+0cKbo7wNdH9PyO/YRBeuq
7wrps2ybYIFEp+wZKZrK8xQcfxKHIxyITbq8BoyWwf4Ra8Pgg1jgoR87GbhBFxXVWKodYRWcmOe1
Fil4nnKu3uZFOwFHccEsFULewni0c+QEtcpeXI6Dm0IR1WK/1iGjkq9VsVDyVxBsElELvTrrB9xX
LTm+WRD5oFaVzK8dBGoYUGf8jPaNUOg4KhI2zpqnA6N8FDl3SP6cv5crdjSmWHk4tL6aNPvvBL6C
PTQOUiJgSUv4QNIgDoVKeqNV1WDcclZrOlET8/tAxbYau+Svh3jmeFIXkadP77A1GDYD3UXXO97V
g9gOTig8W9PUa2Mr8rKMlUlH4PkDorMgw2hVarn0UyqOy8EB0Myu/FIWnBoO99hXWGbKrAw2teEr
dKEI9yMFJiTyZuNHj+fukVObwtJreePn1e+vvKs67U7aiGlaQ5qg5xw6YR3LYKQVLWQxzAgxX9bn
6uk3uH1TFjhd5I4Z43SKvIFOdkF+GtlkantaEBR9zMCUvbT3xPcYv1i3TD0gqrh0rNWHWyYHH+YG
a/9Ze9SjVvXKIGv6/s20R7m4+BQm12c7bZxt0rOXLvrcXKzkKvANZl/SDC2znfFC+KhPt+FxZhdL
9s7HmRae1+6ycX/mL/gjOX2FKB+aASVIKc93k1tIan7uZ4Q9nPIc1VoypSu52Wzye+HA6QkCZbcO
ij0/BQhw3yQKtaUbdBNiBmw37oxNndmuV3VZSDeULfXMq2fpHql92lmDlw9vZgfMhS4zBKfn7euK
jbxpykMobt2qaDk4aNYelpf/52aUHHZB1sw50ZCAiulAtBxOuh1d85JG19taBbWbFN1gdLW4Ymei
3e+m48/8pDxzSfDKJCklffpQO6AaNhFZDQGC841sHZuIhxnyxLbnxXa4Pj3EWyF3GhGf6lCZQlHL
Nv/Bp9UOsq6dNNzF/pTya6ibiCH2ZoztWdQa8YXSw4ErJjabLV2oIYK377UtDoB2ltEDYcAUdcPz
uwlirTXGPVAGy0OmoTpVxYhljuCkM216dO9jGtMg0pi9si/GJBTz8aC9ghkl0cWeB4cQxg3Lr9CX
KogfXmHrQD8M3tEyViW3GU6lCTb1SEQLfSkVFQNwMZDtvxcmm5kfbau+ojEgGBv822msz/NV+Aco
lxLM75W0ujgUCrkY/c5ebralYHXd7kd9dcSleWevHELZrlw93HWygLusT5H5Wm+FvCcflOtQbhi8
zrtzEkbx54MGatPFP8fPjmIQK3Ec9VN5qQ/l6WvSjYbP6EbpeV11m5/NBHwWDq3zvk+EOxAOCKOB
RY3BZVoZvdpdlTNTJRFSs+VLshx80enpBJnnRr7vABjVZihR9MrOPsJF0DicZTkMOmNJlUNZcjGD
mW6TsttpxAUVIxEs64/Uye3x5YuZFPe159V6IBoh/u8W2c6d/XKr51ly82DeuIccFnTKMy65dRDW
2Njg98CU40XXpbKqcnVB6A6lWc0TsPqaNJX//SpIyIltMqdlOUwO1V1pq9uP16tMmpy7aNYvovBm
gD7wD26NVV943xMOTCSf/7Zdx7dqXnjfaYourQWuPXA9qRWF9rGBOF48U453XQPkNeb1BDm05K6w
47ZUypgKT9Gi//zU+cRqq50lDfh4FswRRJ2fbSkOsDvmBfW1rU0U6PtIGXBKjFzVEiazcFbzdpBp
if1QstwXVFhVhXVnWcBEAM+uc2n65mdBfOLFeHm3ZRl4JiydZPtRuPuq/vYzgGRDkc1b6z035Wok
TMrCFn2hlnJYkyn39ghm+RycC5JhxN9qvCrJioBjb8aCMWdVvIuiZrOf/TyPN6UU3Y8dh2K4Rh/I
xnbfb7TlqxzpAeUDLvkoeR6udEyPQ+sfTM5Jq42AYBUkSBxBKZpLyazbS6SELjH7wybKi3SYz8ys
DpTkj9DhLmfG4mWr+PPeRd03kX4bxoEA6J+3JzqmjRIT9np4vFmYvgiN+e7PPLsgqAL8KU7esOa9
ZLx8Ud0jD2n0NCoWCT4N+xk6VKYVq2OYy4k3wqnxM8DAlo9qQUU4oh2ARJwvArx/ktQTV4RtNf7v
LCtOvPzO5wU/rCKhlcGpBKV6dwO7mNcPKpfrrqsWgIMGGoQ+yKL3HxgZg+/N8GjDXzj/xAsy41z2
krugtbySaM/3X0Mc+wyv0VeAyYfFm7JSLmRUHOrZ2G70A+JwXup7OjQAZ61q3KL+J/QtdGbCyzeK
DKov/9dTlseKLNurOeDMNnXNEJq8W4arf0cZL3DNbjgu8sjxI1Zj68w7V/6PP5Y3QZEApS8m/q3c
jeyzsG9U8F83RSkwsl4/ieY1buoEZY/r9ESGszI9aCG+K1rB5UeaBIWCWooKX2ZAV4N3CqX7RL32
oQ7rbir0smqDt1vc6xIfU6EIP5N0M0xQzlwd5/l2Mh5mix4GxWw6/U6YMXk9ZX08Zoi2V0VMG30d
jtvfP4MJO0cj9dp0G8o8H//myO/q0MvbqGMaXOeUNbgtcfUKD8TbwwW1WYFyApI2OaAvnturufWM
xOrKQswnitMmZvQQqJpXfPulKpzTuGObnjGOtsqOMxFdARtmpRh3u0ibv2eBXYAnbRcuUD08DCYO
FM6F3MB9T8K937Yfig1OxLLLlhYbpTKjPzQzjMC79GiKBQj3d6zfrDyQ9Yu4Kboh7U8MoqjptxLL
w6rxfx21WnWNcooIbJ4BqWGKFK5K4laG++GO0N3pUMar7MHzg5F1cn0c3fT7F9rdqeZUq+p2ef3N
Y5uQVtzQQMdjUHl6AN1L9V/v7xiLGnl+DvypICgeRUar7NC/TL+xHkqlNHN0KLNnTJzsHyNJbLo3
aCON93+Mc2aBBk7qlnDw3LTCuicAlFx7C4Ha+qaCinGT70zZiLCokZGR2a+wrqPXqnRzDa0Ml1T3
xWswTJS+L6kGYVnbhkUvDbT+uRJjCbaK3oxJ/3QAWdduF4O4kqGPtgggJhXca2wIr3VsOULjyEQz
7amUluLdxSZ1DYmjCnRTzpfYY0BGKlwJTlAlYZchI3UBgb2EvuyAzYEcNlETzhHGSw/3c9AsVj/h
nt9ybestaZZyNzvRwW3YkJDKHVi4bVVdC3wTs8Cx9Uijby9F8fzqzPdxHM5w0btvVspPIihfUbQT
SX2WM8NdHDtmZ+8yO0pRgSV/EulaMnh1VB5+KgXRvY+TgqFpcW40viEcqzxfRqrzN/tP1YnJau6v
1JfiRMpxbq24OmnMkM58bHnQO7qBD2pxhDOKN0dfS+nNtUcmfX7ESjj66kZp72e5OHNjBwoPoj+0
jR6iXIianXNvh078LBM8LplwpyWxj3JLWpw+QphD7AzXMqjlB7g6pZ/INU/eVVEUCH3D4YGvGoYx
emdl2ZSCVzQJU29tzuBKIzW+p35rwyASOpOxGUXyJTKdi08DPLYnpzSgo035ejIz1+0ThQzrAZ7r
7jtJ6HFAlWs7JXQtnRbNw/obRcQFUSdtrecXW0N6i+dzcZmoI6AN5hW21EIN3NtIwwhKDjB9NFnu
szLUuJOirpQxhnmPOmosqqJLt/DRtwFdGOW3fn7w53BAS+Rc6V7op5UgzwmD52MkWhsPMNJUKlrV
UbVXvHoIIV6Se7OCbfbFn7gUMW7VDp2SSRRkpuyPS+9BXAJdBSkzjJQ82QLBR/XVYYWBDGXPFE0S
Oo0ITN5ANC0IPFSQv5xK8uPmDFRJ5KXQvPDPfaM1z8hq5ERdIFeCcZLZEHs8JtIknVfhaOPIV6dI
feQsNPgpka9iqd6gt5pI4gXcRwgnIkrWmnfrenL989pOlsJ/dweTQUvYBgK/rEw/9KedK+gqq+Ha
FQv/5WQDlZEVuQhnwfMpn6xm8X5YPun59DJU2yTIs0ilcKer9n4KnN946qSKDq+GaHlpE6JAEmC/
LOj/4kVOAXxVaQJCQOHPrKu7LwgcN36vt8fopFE/PcLbN+kgAMxMoMdWdi27UWNMFRAglTJB8U46
ib0QjZf42c+hXq0Pb6d1Lc/b6Fzw/h2cN92Fzpagh3ZgxkY6NFC5T66/Rz+Jca6E5H3n2hE9d+SA
whTVaNg8zA6tEGHAa/+Vz3cq+7izzgAjwwzbI7b3h1n7HiGJKF05LXYmj7JpvElUPgYMfzlf0cH8
tIwY3Nw4FyPw1hJ3bHRIYyX7BgpxftB+Y5QeeRVqdwhZ6EqrcNGZlKk3Am5/BA4lAVmF8YIzIWfx
fSGysvcet4DH+AYfCAcDae/c/yoyxL91rOoIK8cNK/J7Lp4QZ4sGk6+Z88YSeoDaBbO5+4YaQMNN
kD1qWIUWVaWxfb1fmELS/Ni+gl4+xQcUs1feJXgoGjArFFJQ/W+4LbY+8dyCiWrY01vDoddbzVA7
uMwRIqLjvn6Bs0Xw1YH8N72rmbBzqUiZgRiLWZJTiaZ9P5TYldqHsPtVr08GKwjZ6aBu4ks4Hxo9
g9S+3Ej+7ialFrKcsD1DEom8ytMUmsW9m9Y1K2vFeVcBv889mmkMhB4WaDZCyA2rJ5fkhzbg/hUs
0HNHgu41xwtDDGXXOwAfn7/2O38lCXC+kp72nSoiEpO0dz0Ec6kyyDkBIJ3uvQ32jMYmrxu3i9jU
3OJzPxgEY+6qd8pq7yfJdpB7T1VJ/VqvVrLCj8uHS1QBQcj9BgoUPR9/DOXKhCHGTMCEFEzh19IF
r373mtLdGEN4rD9uf96OsJa2tBgdaChwWjIEBPKeFfsDFn8aGkK5aOCcJDMXJL8XAmwVAVIul59I
ZnrnI+yA4iWCQUSS1WGu61jht6yi7GBHbRFs8Hc9509iX8Mik/D+doQUlDNY9kA4Gdpmax010ceb
ljAA/EQltEbFzhXQfyu6xgoifqvBPAVnlCX4DrVn8NCndURl6Le2Hz7YMOCw+nne7DZ5bHuto6x8
Zcwg/tjmVqnC0RKv119Q05AdOGye+NmjhZEQJUFenaXzGyS/lVJXJBVjnvXZSgZUwC6d8Qb0t4RR
wTOhM9vDk70A2p1+mM6vZEDso9xqOXu6zO0OoJvylVK/M1xych+l5ZNWFdgMeLvCxQY4ev9hRtEX
Bn3q0j8rpXMoPUGjo6a+SVlFDYD/k5kHgnmc2EwMtozHZjJdn9gUMH6Q29YdrY75WCZkAmSzma3S
fh12bH1bwSNfPJ6V1NXSFh0S+U1NjHuuXFhDGS6Ik4OTW3slF+7knnBB252PRXcI7Iqt+xBipsyW
fnj6u/+K/AxExaLx1XEms8VRXX5+lQHvqxqoKLu3P128+LUtr/26pcw3Gs4DU4/upqDUINnmBNTS
VNoWv5H52X1yntXm3ILqnNDBMhGC3NXMNO7TVrXY1ost3Wg7i/cU/uMwQJFEBnW26RFjkPh69EQB
bRdf+uytuSjsTr+2+lUNbAoRu9500cTrwTDpltjk2ywWO2vL1wM78VF3jynWtfF1av12NPcdohUx
0Z0C4R0bdZnd6IlwK2qONrHJ8X28YdqmcpkYUkNd5d47+ISNdEtnel0QJYDGclzF8Ucpn/NFesKP
Yw+QJyaJQ3/t0qIMcBkK79nmUcSCL4PhlHm8YhnW8pck6uS5uFPm0WYG0GO+uBvx2ang2X8YYFKM
9GhhKp62+jY6NwDCKMZO74pHHdmkJoEsXwLcXuuVs5nn7qXrWmU=
`protect end_protected

