

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PHhkNkpzHyCJ02b/zcKKV4H67KRxpe36QtGSXZ4oANg/Tq5UCNDHZf3jnecctZQreioRQ/cc6TC1
6ycytB0hyQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bWdkQD7iXQyADDoBhEMorxDwaorw5ZE+71aQZ7Jppo6RMyIponN+UMss01BI1N2b3FJS4Zu3aLYO
px6cO+Vs57h+OQYvM5Rj4nWKlm9nBZ41CnWAwleG5eX8bZY42EI0UWD2fk3svZhWuYfYksxWdUez
7k4lE0NIPu9XIkcIeyo=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o0D8irmB4btVuZMHr7825UqIRFmxWPRwnlzuAQTRAkVGag0/uZxMccyUEuNVjWpjJLtX9sBqvYWy
icHrTQtTi0KfJrS8ikJrBTfSeheDRWxGwQbktHiSZlVIs9ZXDCQSHR9RLWTw+n7qd5CPOqFF2ZBz
CDIGHs3Y2Z49vgia3VU0kO3DEW2bnOB7tyT+k0mbUU9gtzpb2sMIdNXoECla96Il3oPqhOn6wnqG
fxyvNEDXX+9ggv/b3AJ8f7vQxhTiWZRghRRZKvz/tDenZJMI9gW1b+QTVFaCpXETDE3gVUMo+pDT
gkeaydaT0UUCdzbodNgTDg5EzKNdDk7z2pWJpQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bZ9fmUhBpgsyORCOIb7xGyx21bVvbIGX22TkOkC4OYVBlblOkFTGwpEfpvP1tBLXeWHsaAsYDaky
+MMNQXyXlzUHdky+SJLxX8DromtiDW0Twg97DXw9QoHET/lH0ZfTOCzNqJMGsxq4/5CuYlwtSt63
Ens5BOQgrG5RRH4Xbgw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fgb81NiSq62dSzr2ywLopRavTEU3BAdPPDhwK9GAYtd64X7TbKUCX2vkWpAUxqNGlnbwV5x+UovV
u/ZXmGRsX+eBE1EPykp4L/3bM3DF2RydBDoHDxeMmK2h+VrqiSaJktj/VTY2xfqO+bNMcU39RNml
fvwPsqHTJOMpNsEG2KsbtSnC9aPwzo5OxbfrsYwLtETkRL+nMXUlixjY6elVH0lotf5n9KrLTEVj
WB4Jxad1k9nwwYOxN3dJ6njufJIBiBpOT8n8lJTiWbAdxhlaZDH8rzWrGbPsBS/2MHuGWVgaznBU
bEpdCIot1kexUpnYXmm6yrI2OYokdfrieezi0A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20960)
`protect data_block
McnLczamM4B+bHS1ZVX9i7jQw1VdXH4BQ+tY0uyRm0Mo1Pxjc6Mrmx9GkpqI/G+mCOa3daMTD55Q
69SsDxiHqJXVErQCEX85h8Iz5B/gGBYJgf3na5+wJC8sXZ0CfolgWkwAAl8+FMwKdPrGHu2DDYyl
sm8Z6tJCAnRE0MijpFxa4ER2yDgrKgmby+XhLK2tzK2m4aTvl9asATSQnwW6aKdt2gklAjdGlyoP
N0oSsIiTVAHK6ntkWB5Xxct6DbSUeR6IOB2YvMshKoKGjK1NztASWyRxIK70YZyScofdnmZ6xug4
QMcdHwFC5yMzZ9kCWgPJOOfrd15wHAy1bPiylPrvuUmME+3ev8qIKWgeuyBy7fMp1aKrbUYvspdq
dCAQUwobvOR+bejt3J8dIwYw1Nkit/TCsNY/Uw9p6tMwG9wjKg4GcU73K17LbnYJkhVSyzbtXI9N
YRA3qNCF32FaOUvvuQKS9fPJnL56e4+q0fB71S8kUv2cr9tsmxFISEZrcP8aWjvxmVjalYhSeuka
zWf8ejYm0+fWB3tTreLyhhV2S9wu/p3VkwjSgU7cE4l3G6+hv3I6bceWNIcOPO01LQ4gJAwCynob
oJP8jSzY1oTwsWJO51Yrg/z+FoWMo9SMtZra/hLD9Z/F0D//BC2zO7zp4Z4tCmzS9HadNFUmEb5g
VloUoV4i1ts2xcHTKxR+CK+2kAg5Z82nZ1kh5BsXRpCPcZU95U43v4NhSAFVzPVLSDDZo/K0TkVy
JE+FQ15iOhufMFJQ5F71LTu1gqM1rW9u33QYqWyzqiLk29iGDspergNLcBmTK5FiGs2dmzS7/EbZ
dmu4JHUHT91RS6qLBbMaR0mn4BoUsv0bjGwb8SU2l98wj63msNx6Co7zrwhZFKY8SoBhEtW0qUG+
I+1aJ2L7fdOiR6Zf4gotNQ6DC4Q188BfPshQF+gAzXFBm39HcbkndK6wW8npYy4B1nw0xbXLSB9w
HXpNpYMANycaVMjBRWiBZtrctUjBAutUOfRihrIJ//5G6XX8Fh41zHRyCfAoaYhAGlGDOIRak/cm
5MN5joEOnt6Vd/AuGh5tlPBPfrRhDHeU9zvgRd8x6N0mUGUOzJs04bI1BhdvKPxm1TA0WZrGxn1U
5p0i9Vs2+W265kKH4rJHYrbSIVwX6AvnJWL42KZfyG2CWEIYmZJpwkj+ySUv+R13mmBt+Lyox/HZ
3Difo6cqNDD+8Ia/0q7bPIGQsXxsAZhF+TfnXT56+TTvln1UscKG+sruX1n6lFG1wICvXq+7K4fy
/KA+kP5XqAXnslq5vbbSDPYOpE43vB3NUmUgDgOSeVcPCd+vxuE2/nNXfijCa5LvxJmovSeB0OCg
uwEq8dcg4P7L/79aiQD50hF9rbpZi4+bbF/aVTjazv30xnrgQigSTbrcBED4knhTb/aUI500uMLT
4iboeo/lnh6DMXNKBYPQjE7C09gwPUjdrQnHdNfZfA5Bi6hskQcxI06ozw54Pbu88aZS56Ma2NWi
atV6vt9QNUNTv6PE3hu1DReeyDismQRJ2+j1Zbl74WUnlpuPhywQK1nFsgkQpCL1Mnw3lKMxy5fA
/+HcsLhVfl5lH4UTOxxzhVNkil2T8nulzcNIL+6F8475eWCYi9J5OHDpd9XI817SGBTPIsEXX56h
O8ht/a7uwW//5uAJhcd6Y8TpULPheP3QF3gvakC34Y7X3SDuvoaoIJGE6rxQjWDZ5DYKcR/CZSj6
dE1nPZB2ipo1IZjfu8c9VTnQhEa2u7TisKPckV9VD4ee00qXGCKoEKTBcYVSbmEYkxX64yja/oOS
BiPsKeSzmEg/Pw8keDu4JaoHFEPNBEUkHsZNAxpTSPR3NKqBT4NQZhctIPivKneC5WmvREAgqxOm
E9x3DSBqfGV8sw0yUFTMTdflSWxDp1lp3I/OYdsSSbss/5wSeugZn1L5l/DgUpH7ZpdNYffMGCmj
/agcqhsZBIFo75qnKhr7JVXH2dm6Fj/n8LKiShg9HmcGfMGwuaOuKMRkcTfYYIZH4Z+rqiqSSzFg
ZXIoNMo0jIsj4PH5pOPhwOgp1R3XGlsrUXOHdQdM5smU+MObCEoVRLY7glxqrrZAF9KJXqL0rd+3
HXC3nicYrpob1k0zR6dbBx6tBM05RlKqWIEzJxei8FJO77ajiIJ8vxoqALPuEAei07pKGswo0Cb5
yiXutLfZRHiTBsgO9OgOncu2Rma/Co8AOYVWGbh40ze8A107H+YnWky+wIJtO5x0oSTLiiIiL4+c
qBLFc+layeo+WQRDWMF1obEa/NrycWMq2markNGHtgjBIJdxRfwbSYgd1Wtr52k+696UL9seo//D
VChloj3+Rk9ZtoMQOkDbxY7hGFlu/9aYP9JfMBOW9H8VMu7ql80SJhMcycAxvJ0/B0JPVLSjVUs3
WyJCNSWrkRspfWAG6N9JZlreHCeRmV1U9hgtUJG/rmSerLWJIrqn+g/dI9PUUKogH3zcfVdmHIRd
uCBRX5yIQgA8pZ3DR779N19akauPZLRRq6Y/O4/kMJZBhbtooHmqDmtuFhgQeiegasgpqj35Kc4E
X4Zhb8xOkTKlzXaTbdkP0yzc/QVvjh+V6LGef+eQaRvWeOn8jpgox5MKriEpOa5Gnf4ArwnmVR9C
kmhMSIjYR4g1SKt+/Zs+GWkYssDV26VYcTg9qUb3+gcZ1FzTlZEt5OLaAv6bS6aROoUrJixZisbn
fmDkjoYgULJ2e+Ngefsq9DZc2ijcmTADNQsuIJEKh+IaVrC6qaIuFdHpz4SXN78+zwnuiGUqVHV2
46bnrTTa27f22e7hBShCFuKMDGWFloG0IZCcB1sgNWUKtm3K73/d4r9/CwUZWzVIOBvD/Rdsvbxy
dQc+ca4ef/4Apyy/EardyD0/A2V83aCV72YiZZDBKZyiruo0BZE6qrWIkNqxULypMkxqoA58JCXu
x98sk/xxh1ivu9/EdKjRGsZzeayHztvvNGv/kWktFWwmjKpQYPV7ul6pUgZ9JezWF7wGRzb8pmN3
DJrOm6/y0SGYR3mh6CNICUBAxv2WlCZkoQNm1rt6KICQOblnw2uQtmm7bQbHpETKTcUuX6NGqtxw
pocFZ2cVCpdTt9mt6KWzeHum2xfKQTeDXmD+iliydNYRFVO7VDbc3d+e+mM5Pj/0K+g377/t4duc
H54SYIygUvKyeZf50f0BWbcqe4NnAPsZ3WQXbHCbYvS/AbckKOQCIp2yLFEmjI9I+R635buMZR+z
CNic6aCU7ey51ACCC3jROmi8tW1GFBvL4pjBlFbM037k4q3e+hH2HGMI0PQtQ4x1Ifi4ZnW1Lpjn
+0Xh8ujTQle3YESnK/SPHtufBalnvOtVcWczMRjXwn6B+F5KEF5Txxm4ZRJwUEjvP3VKdfPMZF6N
EHUhywhb1819U6CnQJdTcdt2f4xp4ycs6O8AQnAT0dyjlBpT6P2N5wHqTkk0/gPnm1jxpNKCSHbn
NtZ93xrOSjW51s4aQzAOSxHVdMiTCpIlht6U9CFKv3fUFYCFmuPhRGwhBGJ+MHMesI2QnQg6IY3S
MeBe8+z3kJq6u0nZdtMFi5urEWR6ZdB/toMs5RoGomdpwtcLGzgGmGaOtCuamkwTMDIM67Ebglhx
/ATT0A2jUgOrS9hLXdVs5rIjpII+LZROmzu/BlNmYq6AdrC05/MiFwcf8RSfuy1ELDla7TfTDAVK
i7WxgIIjLqXCzfFNRj2VpGnTOR0tsKLLdmNj/tjhlyL+xsC33o5JJTvACE0niWLpUpjsPXOwVMZC
Li8718eJMSj7XfBVeVNBsShb/41QYMVFulQ4bkRr0Itt/QvvlZjlt4/Bq+Ww30n1xOPcMIkZv5VD
lReubu/iR9QTK7/nGr8bqqvYygITBQwdTnhzdsxmYuMr3Os04/MYQE6uSEruxSqsb6SdsP2AmNuj
jg4kqrmsigXtizm0ylkdJqgoVPbxQTm911FcOhtRmya9Cbz3TmuzMVJZClDtHQRKCIH0YBf8A9NP
9ngnfAFOUu2wCewGUUvdcecfcXY1hP523Jvi5GtI6D4rdWRxfBGKSaTMf8/7zprULBAvVqPt4l1N
4vmzOv4RpUkfk0jlBeI/9blXSBwgv1Y6yo3CeTKH0RrD86EeaKZI1QqNnaxAibDXDOX8KvJEyZsK
+MRAKsyosoQ41bFhvM+kBYQknwlefCJ2OYzWdrCXYvyxBQEokmFSdMbaaV6R/0zcd7QSUUAaZGGu
uJgEMtJkIzyLdTmF6/xbSC0/MY8l3083Jfxct4tWU3zV2unGCPva9lXORNWaU/vdxINs6BZsz2/Y
sK+GAFXu27zwPeO0wJrobusblKPbfVzjpRy4govzFqT0WNE6ktu/JQkCPNj9cF1JYjt+v8ZyORI4
MRIypTYHLbaX24dbUtW8F0X31ZJYHX7uSkscuHU4+9j7+6JctoncKvvFJoiw3mCeHc7H7dFinSxB
kqr+277zEVEf7ytXBJiWfZHx6z8c/dm9bVl5AxQCnzVFgP+YZHd8kZOmldnf7eVS4vEEeejJiCYh
5A8hC3O3JqJCUW+QWHC8GD7wPUMSIGn+poJDuhbTVaEeURq6GeHMlcXXvKtVSwP0lW3nXhW0iaxS
vEwF6RQFfEsWH2n01fKlK2x9UpkoJzCcTX2Qbc1NIj1Qp1ANEYMgl/wd94wyEAqHaC+DYBJcXERA
EdascCOJ25u8eWf7rHO/YRnKVzj0TKslr33whaq4CnuTmRaqWO/mJlpXP4yimeTRiomefTcMJYXy
0vWRAuB5gWW98COLvXimuI45+6g/mzJqC6MxmNXWxFqMLdCJ9L4Bqk2kcj6WJlqlwpgi8lJaHVgU
cfwQjWNXlGjfMsp2hnoYABZ2VFY5lzawPHFrGddzV3EmPVGgC/j7ZOxqQwiI0t2tnbNvBD4JyIzZ
OpK55uhCgM+YddDQULI0m4Zzq1ViiQVbaTMIfgf2+yskivbuSQsdgqCKS3XMTeneKrW3VJ1z0np4
vbMsXQiuZ6uxMmjlRuzeyQjG/0hGBlZHuaHbE6KD1RDp++QUmJcHKWQXgLuQDxFMQXE3VrYCNEVg
f9O9tW3QiwD64KKGDBOsfDzPIyNyYtBGQYRABeenPft0A0bEwlGlV4biIR679fm7G4MgFYd7WCLl
eXEkvD9KiBLvnQzYG+w+GAfIdEIp6K4O09vX2ncmhpbfX/01D26F1JSxbuaxA5JTQi9JgV4aZMhc
1vIzFAK28kFDaAsRp4UBSVgiq5roY9PgGCbY36e1uzoWy9WGn/CBMt/vJh4rKJ719fvZDecco3HQ
5pRLJOZAkqzgOHHEHTzqkeE1L0qC6O37EWeMj+B6drbbWX3aRiIXH/U3B0QYwuxuEoLqF/UhoRCL
lG/vPmH1eCV57kkbBCEO4Ncn3HbLrE4/5asE69wK1nNk4ztbCDp0l9fnv5vNp3uYFb45zi47/A4E
xVLvux7B1L0VMLmbdbfLvavnMWrEMoZQS5XWHBAOULpBplkfEQU5Ctswx/e1gcIj9Jrr2nwpxKUA
nMeRkfOkGjfs/lX2Yy2D/PUiCJmpSEQRTx0cwcCklN2c3VBMpEi9Jp7hJJrYHI7XT7rnCXqGAKfu
pqERvOy65MSVhspd00bvhtwC3nd7HQ7iCx5Iwh/CXg45903YA/oH15GFBdbrKAh49Uzq1YcEh+Wa
WpjJBnuIrXjgG1I6dyAJGYRMZ5KbQGNr8EsQCG0AlRYUZLTrAiUHkC6CEE/pU6n80GQz2NKqsyAK
ZpZupoWvaq+2qM0PAml53H44ZJqJ/ChmOJnkoYP8XtVsxZlf5S2+q8/LT3Ki0EGVaYQOR66Aa51d
6QUl3JYCf+csbTFAJsCQeHZ8i20i1ZrayFILEDueewPMD+M3IxvUvRO3vmWoBmCL8082JBK1zE6i
N5u86N4NQveS+tkk33aIkzRpxQA7UOCKv09YTYdvWm8dLw2uJM+r2RnJtrsJbCQLWGBKBKqGCkjV
cfvD1qXJHKV3vvyTS+PJu/sbZqFIfImv+mToJHRe5lFOx3QC8qTRfuqCXGiZwobxfe0X092bBoCW
XJWBxewmTEsPgC8fQQiP4CgcKXekjlaVG7NB6VVMINMrtdf94i+PT56h5RKGskn0PYpqulHH4wZq
xSCFSoWvxVz61Lybb3xw1SDtF8bh2T3SkUPPB9FbJdUCj+vlAlDgp4olJLgNZrnEzILc4MbjBymT
0dGdJjypC72wBAutb536jN28MLMVHlSa6xkzV6K6IsT+78HOBFIDz2I+uAPxVBh42CjO6GgSnUj9
dCNN2HfIDQOwc8YYg8kjMR/fP0KiP8lv+0oRT4JHdzcvFGNubHVPU7J2S3GQmzZKkEstf6TVf8uw
px+w4iU17jJ/exMccmomrx0EmLeqWfwYwQ6GitTvD1pS54/22OMdMlu/NR+yFVxjRxup4hnq+FEu
NPon/lA4glxkS4q6WE7wqi3+1SeH68tkC4atv2dr9pBAeXVkRZ9TWuR86EqxH0zmUh5UaNnSvivK
J7EDlHN/I5OyhDr7IbQ+zq4hFvHTMIrJl/hDFtshoSuVSJzi6Vxland2/X+N0pdOEPecp/NxOTvk
gqDse55JGnrfPQv+snbGmGF5BOVYsRhbg0/OTqRJpxIpD7J/N5VN45Efw6+YxyPKMU3yZpCT6/MB
nYIU3zU7izo9q3D2b5JWCwU/36228bM0CWJ6wzYX/SBko1TY5e1G6s5vnwh7c0eSkxmBVpNblhpv
CQYvb/RbviSYWiQEG135XnzXVenHetsTiLYDuLED0iHbf2lf7ZS1NvMdWzexav6m3uOkYfr3zi2W
rENUMz7x88EU89gf5GSfJJlcrOjRTlTNHiYrLZqnn5yAm64wqZw7rqH7het9TXKwef3wQQzy/WBX
bHTcd+346LJ4vVmRkFbn8z7e+7fHqDYR30EiuOQeq+NK6HWL9xLGtthCMwJ3qFcQtCXPTh4CwKpp
BkAAlKqMRxI7c6K2V9T8DTZmb5BemhZsYiqc5yVE16MW+YnpKigYR6agl0O4gb8iJ60JD4l/gcsB
PSAan93lRQOvnQ9R30kAIN3BP0fE+pceURZGl3ROATJkdzerS4zNDSVzjvwVN83CMVnBvo+mdBoM
xiAPZyoQMVVjkyekEJslBXpS0LvZ3Ou3C0SO777qecce5ZhDxiiivNz4n0nJqzqmy5rv25NlaGf9
w6LPBD8nf5Hfrj5RfMkiSgsHbQhqYrKS0n7+UNYazt8H+JjF3qTqCZDZAQLOekm7bDkFwgBjSjri
6v2cJ+yrG1Sd46pFhuk4X0ue5+IA1kalDTSJxEcLKlcELWM+5ir2oYFGdr2qWaHY1QSPnBfXHfYT
yNz5Qw+nIy1mBK7tT8u83uZhsgsGI7WqSwkmz+QFwWIZbxtjfxRSEWOZjYKKdUWmHbgPOYl9YGwm
6jVJbZTrfcchEfzf78hh/T5HMA2BBMomT2R2AyoBU8zNOaknMfb92+Y8VPzqQFnf/LkvbGKzCaOG
xvq22dORy42TEEQWG3xwlFp4SRIi1FNdvLAhhvyZQkt4ClW9vaeB+TkOB7S71vhDI0f2OXHhRCm7
ylAKSj21cmbYux2+dkRgxovx7U5YGs1yMnexHlFzFKeJIUEuElVBhcZAh316ANEnlUjqFDOXXCEs
QPR72W8hwE4s9hXEwHxP0mtKEIeNCpHg94FORDajKYBQ3eWIAkYV0ioDFfeNtfJlJcIiCHFBkA3m
CQERLcpkEjAtarGZ5m77nBW5+7/ycXZ8oqBB3q2CnxNXIgyVPRZ0MKUIhiRqUBijDCC2VRkV1KJb
69S0TpKDPcOYcAdLk28UKwqS4U7DDgDPeuwiMfbzhY3EgUnJV9p5FKnRvK9AWgUOoosRnJI2OQFC
XniQJqRNY10UimknNwDHNstMd9ICToCBCfUXJ7/kZIJnes1cVMJcVo3IsBzgKeW+Z31mB4UQqrKe
+PpHWlmiRXskfU+ZOydDLtjfskp0oNopLRHXiLMk6mW4hjbgHWhmY2TDO7WX9P6fU8EonjppdJ5J
IYVbpRHB4jFiA4JuO0SOaio7tcWWImvQ/OqnvzbZ94g1wwLAueX6P23j54nXD/BgocTzGmvo/+Bm
+x1482cmT1JdsnTZISQL5qY3HMzYQHwy3OqBLqxeb2COy2PCDa45c6qFLfm9+y0khdSCoHdU9Cyt
9K2Pz3kOcT80P4+ETd5FFg4VymJv34WcnrE5Cxd9KOZhB/0d9B4txHWoZHrrkCih5UYLWoXHmvuh
k2xVUf5ZD3K75raq1evuJNClyd38u1xIVNiJs5UYNxC5WOwIhQrQLw/xN37GUgaoX2dJ4BRVEBkQ
c6cwZz5n3sgeMaRjCq4+CepvQ+fDfQw+YKutGuKCtkgh8PPs6Xb5zdAoO2GIGUg+p2VCD11ie17b
ebT0I90k8oyYB3wOWJJCUWt+Bs3Y320F5kuxcQOByePzdRkLzVLu+1tE+c/I8F0uIm3j8BwW/cXQ
efvpn/lw2CP62jbx2218bPHtbswDH/NczXXFxbW+IicaKK9ejXxg4bAxYNBAPa6vDZHMX3qNN78W
qKn3snCfPkE0Zh9q+PasrOor0qhxUMcy/2OE7qWRupzW0Msc+DZafuCfxCMHV3mbKCotlXK9PJjd
kVmrRE7X0Ke7jSmzNzNaPR47RP5MH9QcOpBp6y/P+n3VUVNekAJ75dApxio9JSAudTcRRTlVFp+2
EpRD/PWMthAdYqJ0P1opw0ANMa55s6vR3yZQKohCnIhi5cvzSNAAqIJ4M3j8EWz5xaUR03tGO+RM
Pp+5eWr9GLAyvUAykXr+nXpqvueUh8JtveqHSTBuWsAXLc+OOeVCU/QGAawR1BrV9XfpyKh7Sely
Hm6KXJUtrb+q2G8209STeAdmdMlyFQaynSA+Oi9Iy8ys4U3zTY4ZlCMpT5Nh1vdzbutjepeAqJ/C
DrdoAspoqFA/iq8aeI5RdOlpF6nTYaEUnmMwIU7X2i2e3FkNsFml5r4oOrXBhJoSHi3DcM4aoQwD
vh3OeL7CIvFHoJ5KGCi+RHPDxitzvSaKZXi7blL9Y3Fv6c4WGwCkDJtnsZ8byFDIBBDbwICL8/e+
WMPSJnWutYKP82qOYzsqPYqdYVwcxGPGlYdp69L3PnNStvMsUg39N0HjjmSAKwf+l5fTEpXj9cCY
jnIrVFDDrDDQzTokFfkf3L3koP3BJubyeFaBgwqDcOGhFaNvxFL4MbSjpavajGwwEer0XVnzI/Fd
po04UA6+c5EhFQqJ8j6x4qmJYljWp5zKf9MRH7Qap/FMPVSMA3vjrjl2AboQlyEjcheuIiJCSYfc
C0Jf/wB1vXiIS/n/AygOY4An0Z3XJykRzka6Qrk9LwBYNUtXYbf7h2JUHO3O6FyxZx3Qde8WUuWn
dsAgwLd7Gsxwbnjp2FdVpb7u1pNPuYQrCziHaSBb3DjBHyeaIA7JXoFGt79iWRhYndBWT28nz09W
1aqrotC1norj1yNH+tlt9cWxbHLc8LJj3Z4EJIHPDQ8jmJ/bAGstk76Az4364Ak6NsmzWxnWKjYf
SolmQWNkKYUbsWqmirplO4C7wCNPfH+tA/R9hu870GhtWU3QhKbm2kDoINgD3sNZya2I/c1ZI3N+
4Hskz6Segp1dtsaBbw3sQ7CF0C37RtL+/sGfRcOb5k8tCuNIOgzZDxtjeiu2ou0J8uJouj/M3bRU
ToAr2GaFijm7+s6tJHJcot+qZQP8hlHJfv7vzqIdWcn/YGq9wmMXQvSz9ISjbqqQJfNeS9AxcLN1
19fmOHGFdDZWpF0K96vLKCPg3M/ldDWjGxtCB1EIoE9COo6NlvTqq6dMgqmFcf9P7BGvGNmKKlK9
/4JvdsLBoeEBgz5R/lYwqciUPzUylFE8AiiQutK+TbhMLV8gpbpXoYxMht07o7OsOUO2QVn7qGwq
VUdz/8kLHKBiU/BveNhONTOmoKb8EVEAUgcjUzTGqtEw9W51HoSQFdh5ZhvGGyXYuaVRyDFIASSs
RsDPx732bHmQQFFxMBYZfVLmDiiUAYIsQXUjJmvGlhPlZuhsjJyZOv1ds8RoyGSkoWIEpLpj4kJc
KcTFMvtEXklsmRfwJtN3X6nhPFOS0m9DDo3T9rhCmkaMmMvRnrEWD31jEUrRD8L+JnAyXLHzmlds
tlaNxwZCa09LrdofZoqriSkaUHGLiuLlKilRo4tnp74uupL4XukbTBjuKMeYGtKNYFLoU0mwnq01
PHwseO8xUKLYcReQW0PfjyFflL0NgIr3g8uy/KX9Jmy0AAYaJR3rQdeqpCxlvsExPZcTMGUbqXDP
Niyt+XFdQkIDi4XbINZWgsOc/+QPXjbgoJ5+ORi3Z7K8/uu/SEh2wPUgFMjqOOQLcG3mQZHiseoL
mMUictJQX8xp8wxPo8mYHfJ/Rgh7gTfxz2ECrH2bv//LB4M8eohWmVB19oiuXk5A2c9jSKQwxpwX
ADHkmfaGxkjkDHvCsXA0j3ccn5UFR2MogcFcGO2B9p/+RMMbObAIQiqSQWtgOFbTbtO0AEHt8fI9
pNcuf0SaL0H/0G/7L7/f/7tPpYUnZcT3AwXOtm3D5Fh3SYz9rPzH9zZL+5ABGClJo/LsAEqJBxyB
5ZpX66YdM1V67mcPVZ/dfGWpMXOzVhYRTaVtpuGedvu4MukjCOsKXYHLFQB6UszgVUXfl2aJy5Yp
H2qQNBOwScHXEi9PFk4mxss6eYKsnqZH2Gq9JNcLc3TFPm7R5LuDzYcyPNDvBGtCCAKHRnjcK9ar
qn2sAoyHA361V/7WqRqsfWu8/NryR0hz5RIwGVHVEv6bmFgl1xRyF6qpkjP3zPy6cDmJKnmfb7aC
mDD6f41squ7aos8Kx/nC+Q5UEdt3EewS4mvZYMEKmLpD8rsrAX2M8rFMXIL6nV7hkjuhr3inMwOH
KT0oesjf8mUjkOnoi8kOjfvFQFEzNehMQNu/xU0U2FFAA78rkWRq/1gxPKq1IuBKaREGk4Znra0o
alZSN4q5a410LrxsxqAFKS5tL/+V0a0i6KkSxH6Ka+BZII5F3t1tQZupS3my4pqrrcSn80+LvhHY
g0dPhWxSrKHGZK9YZTJAbZuiMJy33u3GERNX1ff9JpsmXBkVLi6gOyQb+gUrrL/By7JQIw9G2M+f
Y4MFjVwNw4UZl8Dy6dNmOhIQ956qsgQuVGSfWyEwM2FPZ6N/4KaYcnCA4IY4FYrsui9z2DqaWww7
T1Wpe/ondCqma8plPAcPtObTLncYxoJaIyqKWnhqyIj56hbSzYaLJo07lYEOW3cvHdOQDT1fBMPh
nYb9NvQf8qNvoL3/nGA8NHTcEjtEqbRbRBeGTTGPGPegEtSpqQ45PPULciFSY34C0k340JpZnMaU
Y/eDNbHKat07COYt0z+SfBOn1c2zfS5zdujXAf9MnlkSMSwS1CcDyI6+Xit5NQmYaaYd4mv1efKH
ihZHnlXT9/VQl4a5A7Xk7vtqsyKwriKKrKlM7Ws/YuJ8tpxmfVf85A1SuwyizFwY/tDJPyKDtZ0X
pUYFKCk0wnhrmZxXFhcz7M8vdMXXlWtLCrgaIlTlFU2UlEQPcFbYghM0cSC1Y7YDMnUwjVp6xpMc
LGf82mfQcI6RmXwmMfzMOlKQUkeJd/E9ghrvegGj+E9zEpbDRIUyAEXXGLO3hRz3HarmwfmGUspJ
fQq9awjtJPZbl0Oj9DywLG2/AXtRTRqZH3JKLOzTBV1mCUNOpTMvpihHVGHNvcDIJpJXwQ/dObRJ
7yysmvG6s7u1YBnBENEvdPtoiVUSjxEpX3N/rysxBZ56/ktDwryP4WDes/REOG227QnCAAHEhIoq
AFMhiiFYKJ41vAieiRDzYiNZe2d49xLA89K3aPF8l4RwQXutFp3MS7OtgeL0tNApVhttTfwuhhqi
whQ/oKcf3yxy0sQWOVI/Cniua0TCjxRjz+/UyYyIJievbrd3RCKn4iETMT3z/T2mr9eXcqbtIUUY
JjfbbAScPRouxku+OAwcy3s/a+O6mTMEKSAy/DjN1gcGnUkIqXJw8QqAHHZaQBYVmB1Bhgx0k1MG
gzdyaO0wLG0qEiRP375/8orjalxtkYKN5jAMglxQPicGmUwT5N6pF1ZXKLtWpPPkWHzr6aFLJBGM
+h//9HXIOVM+r7nw/FLnibCXV3Q6roAWmDDu6kmsKkO/WxlBazewqXGO0mOxmLNzqkfUem/mb+GE
klGrOYpQ8X+6l/IxpMAJyUczdEpvuTovx+0nusYbUxhWekITJKiTNPQKO1IJvUQIXoMPo09fJUbr
EcTOXNrTfdWxO8OexsodCMV1S9tMKNOdHfBEXl8rAee+cmwqrJt7TCoOQQcqC9oKGlKbTIg5sQ+W
1Hp6Hwc6lnipy/VjwTCBuNGEKALKowRgNSUh1QRZJVzI1nPvGW7Q8jI7ARkFm8q1ZuJqp44HGBjw
3ToBoUSbnZO3mZL6Rcw62etMLATmVH+bhsyoEni6dqPI45AcNqLpodFrrnxcL5+99hbKkajuogmw
oAYM6Ji4uymP5iZ/MZKHfDTm+svk9bnW35w+YJma6HIdmweNq9LqIp/pyWIFaaVFHz3aewFVvtIj
T4128camFQEEPbs+0Wkp6570fqNjhlsLtd1vi1PIv0H+eoenynkRe3wItUX02zmurZWyM5vrBPOy
TAY36fTnEYX4al48Fr7gLg45fchl3oJciX82WDuBkda4QJvSE5d3WRtAhRbkjxzk7W1SDTvFyo/W
RC6SfDnazFeH4+nUl3TPuSciS/WkDr/ZdPcl1Nf21RD7KKZUaFGBklPdAmckDQGCdW0YVhIWyAwV
RuZhbJ11Sr7p/J9qy2DG+g67m8yUZmyg8ir2lLsxSY4RB2Wa3nKG6yvdlS2UWNRLhhI44nVoBWPh
9PpR1FvoXG15BPN2vOpz42WwyYiANiXP2oIs34roG5ybNb0UXl9aG5GX1ITT6UGnnHFL98GPZWVw
ITiX+irtUuMRE8+/SFfxW9foGeKG1s/kuRTe/tSYUzVsrLNtEi/HEs9NaC+1nX+jfFKoZcBPjZUj
t2DSc+6cQpsTQS9yYVRMNn8SMRjE89T3MBL0xmV4Bv9ILgyc1N1CsxOi8TV2hO3YdDTJUN3lNdZC
nfxhVf8Pz3z34JXzYUFYvY7ShKsHqR83imY342viqSwgC13m9tQL0Pe5uxdJkfxQ9vnYI1eKpv15
JoURbNDzrbqP7RsveyMSPgTQoquLyLAFh5dqd4kVt+0e8aWV7bsWn9pdmR79mCVzRz12IsK75j/Q
ODXNUMOdaUkIo4hd0rbN85t4e/Djyrgm/sAvfmFadh/Lzxa14SjXbTUy0cp6L6Y55/YEDRFZ7QBs
+VYsNNp+pXfC+RFI5U1M+USB4ovPTkQXmdIQ1ydn7+ISJhVGvOG9sD8r1C2r0BfnZGmZ7BwhltjF
8yFQvpKyJeJcSYrkNkWUgd0ZqTM2w3Liwrqctj1JxIM8LyH/Z0TidEmleNpAtApj8/Zlmq6f7C3J
bENQapcdJZa6XYFdzcLnC37E89qZ05T62/YJjCeJcE6NtWXcpcIU4PBgL8i3s+Pv6vO7EHOrJDcc
F4TleIr7UV4rb6uuJog0fwHi5Qj6aG/bplmhgeFALIppbztzZmllChYoF+lGN2OcHiugLwpaa7Hg
4HvBUsh5xblELRUJvsoQFnTtBwlqQioGvePRW+G2tPHwJofKGM4bySSLFsPoD3GEtUDramqA0on+
dFkKkaHapcNa0tGS56b54RXPQvb+N93AJKAktdS3zUqXgIJv+KGtcVrAScBO5NwV/KUl3KpPp0Ye
sXaiXHI++vBAiuU6GVNBUPJ1AjNSl5XaBXbqvXvp9P3w44a48OU4T3Rd8146deb4fvQeb0CA8UEE
GRHC2jVUdOQRRiyH0SxCB5a62OL3u0XqmaDCrp+ENqiMZ8numb389e6vh+JPwb2vczFekdqL1sr3
ItGhaa6F6Q8S+LdTeTwFIt9Mbkn0b8rjd7ZUX263GSnMUFqsDOg2+bap5FrEV9g5D0qVU57vqzIj
gh4kDEb+XEINj5l+ngrDjtsVfhTFghGn0hKQ22qKe6+VE2I0S0HK5YYrCBaKJA8TSPHyZ1EUHG+D
dt4ZCtcwepAd6iQj/ls3HUkzLj3ulARuGD9zSWcM0qbF/7Xf3tAwx2Jv9TO2pMGeUboDT1ks2Rk/
xGcUdHgWkiqcgmFbCLTF9oun8sPc13f006Z5mpixd3NQuuECEGpw1Ep0fFdOaqfz8gEjvxzWVhnP
VvLYPWjKUwI4rmdVwX5bfS6dN11mDRo82H6HNEX1e6+7hL3j8w7DVtsRIDC9vA6/mrmFzWVQw9Sp
MGNiJOyX6tUaGb6RRBizRR/755cov6y7EVm+e/+c5G0jyciiGnHvhKWt1x2RbXZmhFyL8V6eTlht
yTu47rEubV414EHwfXX/P8v20GQYacl/Bi/+E7utaxh0teeCC5BRVjmtnmBETvqOhrriksgL/9TT
1ZDRDvMX9vlbIhpEcmaJYIPPGj9Po1c8QF9Mqa6ixxkd3KvKuyH+HEHjMPM3dL8Ubiv70cj3yoTr
TB5IeJ3RvwlAfpyi95t+2Rcc4DEa/WItfTrRHk/BA1JOxme8XED/bRpQLvWbTk79rZ5NSiB55xXO
pob8i5Yf+bgsresZtyHxOeYvQXq7XpIn1aypUdYGz6xk6IbubnZmnqxbFH0ONgJfxXQlttGTbcRH
dEy1hUI8evBQR760ZCu1n71TEgX4keQVDRzln+wK0g61yMmnjAX5MCekMRtEfgUwH+TLQHV9gI4a
AxWV+3tylcXJnax1pAW1JSW61c/80tpY0x76Pxv/GYq8Kb89TtyZcHN5PqyHvq04wNVonh9hQoRk
YVQAFmyl/PqNacAxen4o/VqN0a7IOWgM1Msq7gJ2sct9FEH6PYqwxaJNPLlynu43sVOydmlX8etI
7WhowhDfg5RWsUBPCB4zFc78uashIKxXcXk8mgrU37COGDL3brSywxVDyFqopxNQ6/9zHbwQVpfY
vi8OscFnYCeRVR+5d77E/aEVwbkQZCEG/qaCOkLf8KWA5M8l2FkLQieLak8g2WLsfZuXDN15S7nS
HTNNkClUg5u3GXUUFnGRQoCFtpMrpTrPdX8Ld7ufVoDRKxtKfuivNy3tugrkKgVu4wgDA4E0W/Q8
1Qjqn4tcWGJjLaQqrr717kZcrTJONblABsEk5dVB3SMOKkZBmqAygTFHeIAgUCAX9fnpV+9AY4uM
fYSmMa8XCy3mEJsbSgMu69QdezXpp1GKz5Kd31y0McJ8tIDegJEUWfe10rxZwaqeoVRjuHm7xrtw
1YlEuCit6jo5vSEujA0j1U5V1eFUnaDHYuEWpqZoLS1Xzfp+RkqMxOZF0AOMECkqaPgmXC6iQEqY
Adj6WGWd8q873SG18T7aq+48SjyQPKNjToaNXHrBV2jaqud3XlERJ+5DhbfOXZHgguapa3STrRed
v2Yk6ynlNfOuPyngb0czDOEKkmXKX77tyb/2VAxK4c2zve/Errq1G4sJFE4eBuY4l9lzQgivz3bB
h2gEkFHstz/VLVM+/S8CC11fHuR6UeHo7r+RlEzLZSz7UDG+oov8idPJxsNIqeq8D+Cs1A1P6/3h
K+FmjqEVYUZQuA1zG1bijMTHjj093N4JZlBdwf1XU7J30kFOOvPc8Q6a/+WwSa2hWJc49936atO0
De1PeE52xsrGIDC/EGvWNF6bcIFwGtfBefPuKzAEiCmwN5FPw5ylVlnn4Ecmf+twYHBM+UC3n1dM
8iMDtPpxnqXMvugzpWjeP7pTzN9WoCY2toKdEaVKp+CqgSXAlLsudcoCHa08cU79BwWs74LEJA4I
q49WHJ58Lj1GKHyWXEwmvAzNIbrSNN/fuUqowfJuWPu2c5vcQNbZB28OTDlwhCQkk+jW8KbHH4Qf
6uvNURZWMNkqYerWnC9y4cDlP8hYn6R+qwriTCDPTPm6jf3ROB163H/ZpwOkN7sUAHDRLM0ReWi7
jy0UtaOz07YaftT2I2SmOG196vi7AZH9iiCzwDTaV9kf+qt9Ny1RtA6tEiszKusjTlzZj5hQoM1O
ATuiM5NAPzQ8g2LAWPl6pn1RW3j5Z9VhZT4JQiIFgDWhDkr07HLrOAXB81nZnAk4ZZJB/g2VWnHb
wI7rTRHBJS5/ltEvg3+jKkxmIWh6ZmG5tt+WhWvVI4qYUZQTDoElTjdDL6HBKF8esPh1pLtXXGyp
oyI/qa9ThrYroSPpPZu7L+aiaJUJMO7l4wmkoSrfGgz8uHViEqI5TnuNm8Nd8mRS1oMjN04pzm98
ixVHSDWwKuUEBHvNF/Lf8dG8E+N31oYOwh4UtTczUkI9xxhOH0N/EfDeELdE6lEBwkwhGF9kHYsu
XVRvu/SDtp+l/jgcEJYc3+XeUVQ7qDQM6HK5n8L09FFx3kte1++a0zpKu+LGFPZ7vlN8IjXm6fnr
7Ds5i36hdeDqk9o82WxArnRufqZrH7aKjjPXnmqkwNJoX/3ItE7JDXCFyBedsxS9Q4SOG+HDWcZE
mDOFg/IeV21dwDvLnJvP9mPSTBDdCduEUBno9ppGUrb9/IpXr7sdhEVR0cHMP9PVNUkux/HrWtfq
h6pa4zJ6383qrojmYj1HZeB7PQL7+hbNcTuYR+n46uxhY0+1WlRidDdCLRxenD/JHE8HhS3y7CnG
5G1fzuSidUTow0dExuBg0wsb86GxgCByVoQm9TzXVUk4KThplFZuucffJ56uVa7boTSOXjSaiAaE
uzOzCXDck4gJRoCj2Jf5/yO0LwFd+BwxpdETgap01O7AX2co9oKonrMmOahh0QSmkOEEEsQdROmV
R1Gc9r7ZObeRfBGJsH76OTOZUEuim3q0gOXcp227SQ5EidXgOsl+J5u9GqAiWyh22eVEECSJuDjz
lD3Nzpje5IENzpIm7kN4YeSuuiI6KlTMTQLzBJkGKJK3THbpVrMz3+Yuuw5ef243lJhUOzeUlHNy
kUZTC2ICRMMGBoZ/Gf6BDDLo+wNsZlr0F3wNg6FXgfOJocdCQe6q9iV8yfURLwSXALH1bR1E6HoN
Axpm50t2GYByGboun4u6groDUom/41Ox2/nl/o0y49Cqlbt9v9Ie8u9fmcwqZhVTa28yAeeozUXr
2v5wNUKz7dYWTmuicEeO82JRVGzgen/TqdiMaRv9KHy/cbBeYx7xOOWaiOklyqPpN7wP3mCjUPQR
TT3hK+dv/yOgrM4DtbqmRdha1LEvwEFsWHl4O01tAj5862h6SlcZZt3MQ2keeyGSALR0Q2ML/Z7j
fIXa15D/GIiuSS8qkkcrd+Zv28OjxHF+WxxLOy7TemrLuvXEGhNv8nQeCi3iRJh1b4xKRGpz5GTE
47rbyZDjIeWO1PYSEZBdBNzBK1ly5wc94z1y4kdm2W+7TOkDWprya1XyIUv3AX1D+aaI/r5r1PPA
/bCRc2+obPdMcGcY0zTnLN2RXK/M8zkOsYzh5opV47XsIXVT18iv50MXzEujZKkZ8MJyB5H/qPJj
mSgAbMZgnEDDgtELXSNrqNfJ+Dt/4whbpkH33Nk2y8baw9VNY3A2TQSxd2QgDZ15NwGD+91LNwe8
8OtX2pCzRRHkNceFr1GqfzcQ4DIuC7ax2Yulg+Zf1mkeR1KeqfaBDEAVIafwkZl5Nm2UOd0O4YXM
Zb2an/t+Y+9V4NpPZlflGlI6xk+df1RyDytAtdQCZ65KbO3wTi+UnjD00inOYjdOq6JiUZkQxOKX
yHczl7g1EpZB5hAYggfu+6CLgHbff045FMYIBGF2akiLS9NE7M/XTNbWgE3JmTJgau11hvAdlP8D
9+znUWVduYbZrM2d/OSw5db5t4jHGo9IVBqQAIkfM4uLTKSqB3y6ArZqR4ZidIr/BWlP4x/Mi+49
GSl2DvxiuTf7DcRMcGOlCxTDddPBMPI8JCJVGuQGbnLgWBovjQxh1py62p73uRmg3LQfWOgoqBd0
FmL5Ma04eSLof9QwQxqnigdlbaSfwB3JywFGaa1ndnKHbG5Xq/ZHY34mYEnu7G22qdGFnEGUIjQI
jxWKk4Ngc+JYPfvbDyy0llPt0hYGXaaeVJcHCiPzUVoJW5YUrOLOBLQgFv2tOwxE/I088KoMxG1M
38gWpTljjsLIS6uPsmJwetfO0rH0Ii/DqPfFlxwL1t6WaR0Cd7Fe2beQvI9ZG5+K7xOXVpjCSbK8
qan0IBcO1WFLMh9z2+Ce2Y7u1d8gZoQdw02zy/ZZsK9JwmapHlfqAbmnZRsT4zzpJyt6keRzA+y1
fcv4QjADI8R/GhLwBL1MxQypL+2E8p9R2PhouPpVw88HBqGx/9hKolH/BCjytO0iPooI/kEz6cL1
Yd+/OxF41EAhNLnyKlQsh9trgKT/IuMuwJTO2viVIiOvK9PrnzvTtPIBqq+vlnR6Nnsh9br0OY6R
ijWZd3ym+Gz78BeduVH0r7B1KGZLlgVle/Qd+hp93o07xQMRl+owS3gNKcxyEHet2Pip/dNfZhbX
LHRTx5TmCbKygnvL+u9HZPVKAd2ImiF/WZ6lChOSf71Kf7xJ1SJlEe9Q4w4CbMjfEgzivGHHj5y3
xkQNIYcqMO5mFFQSjDiSpeHMSnxkS4RI17UkvVGTduOaBk9T9BrhlHz4SEm7jzC8/ujcrKqRwgWY
0+fCJJbKFGnTZesfGZvm/ANFad11WUqEfSXqcr5JqCKeUbCTOMf5WwRoy4fHbUJqGgASOn/uONHZ
X36O2FUm+luWXgu/JJlecFDwgK++WrfYj+dDfzjpFGxh/AplLLbSUDpi5cCfRCb72CtMFfVioUxe
R/mJDQBAWBhpu/5U0PsgGFdBIePuOO5bAuKvziaXPqQsq8LLuv59LqfDsNvYw5zJd02I6daw1JGH
22mvlWclNfkRRpmzrKr1DmilYDqn4VoQbmsnKKZSAFGjANgrPUSlQqInf7P2Nks6Gna/xD5M8Fc4
Kup0QYzxNUs+xF/GF5XkRwGCaRlKIuvO8lhF6AHO/s/gShY+D2B74dn97h5t6+GQamFCvjCMzkRz
26QcI7K7KRR9pJONQch5NF1NbnayIV+VJ2Ix474mhNq7YrUvsdO+rn7TvZgkrTBJjEbE0+83/9HW
CUHRYI5x2qqxML+F8woYaFDwMJQUTjMIQKq6udP9dfdTGH6XwoIP3SBoJ925fziN8IrVdP5cxs4s
AX+DIjAYYzyGYEfJAZ01am+OoliCj9ihKxZpKN92/OOdXlp9qjGqpZX5fa4SQIuDM0tcuVze9Ld8
nDSN1yQCu0oWD7uY8KOxVrpv5GFr1qRHlx2lTtGHawuOuzH0soSnsr5xhnXFqkg5X5xP+TZNBi4H
zFZPmMEjN06hit/9cuk2AOYmaCENeU87UYDTeSK4MxMWGLeLX2Dth5kHUEZ0pzVaBOETfUZovdUj
W7Hdhpvwncd3EwsOiD2wNfIeNS59pKYMF+RQgOASwvAtZCdf5rhK/RTuYkLx89n+NX4Qwm1h+2VZ
A/UilNdKOTm50pkyF60vgk03e21jOtW9uycMr1osyqORZC0cVC71qiJDnJfCKM/pYPiXV7oHeMI+
/3yp0OfYbaLBlc3buLNJkpYwPTYoBekXkZemkyyhC93j1JMUXLz9xUIntd9yz+FVxt833uF1HHJp
/BfPDaNhhM0x8jeSRvJXGvRt53dJhALnLw42We4g4BPSlhQKDeyKcLziewtTNwpFTguYtgjRn8/Z
+bh5S9+rGMulsizGZo5ma+xZWfVNXlb3gyMvy2M6kn+rjiUlhJACKXVu2YW+0acOLnqGU4demae9
eEpzYkwZ3TzxZgJBBGBgAr7kr38A8qGVwW1Iin/kZHDZ3yWEvvpF53yADxuMXGbrt7vI3A3w9lWf
Vi8BWTg7zO7moYE6LtH0SoO+Xwvv/24OxfUN93t7/5KAaIZ6hkyUIrUSb8QuXfUnzHuc+2WtOr+1
fXNl1mxmKyl7ZtT++jMq2wxKJ5luR36CP3RX8qKII7+5LW0KjLMMd32tggn7Lht6tHMhsY70XE7h
eQwzeaMW2bb+rx358ps+jZRIQOLxFuQoK66842bATF4smoes02PBGaMnkZuuH4kVDhU8GevnO/93
QddrqCGA95LM6OLzV3IykO/muH5HdjG9b3TmgJD5Lf2iccNaASjgetc0NuL4qrpKBCT2CujuVG0s
JP9t3np9RGLXQE5RJsFrxYpsmbNpCwGy/Y1CwsDqo+ND6o+qFrSIMD9T/iSJHFSbgMRoMJwk2xiq
D5s0wylbEYZIpkuJnP2sWeoe6YiYh6O6mfzmv4q4bsZyEC/jC1Ff3GdQUpW8FYeAG/ZD9rricpPH
ukMgtSTdLbmxemY+1Cd0wnKyQ4uzJNBVoUywyZx3uML27H2asj4xyN7Y/GayRmIg7ozWv1wmKYIw
hOddb9cCtQqahSUI59Bvy8zNWF/XMgiNhZb+qHgLBiHoMSPCR8DV0qaFFHAqAwmeDxcwKahkaBEv
hwkS/lK6IGtiV7wyXn/caRv7XZqco/lS6BTe7IJrrIRY9B6FXMPiAUcT6Qofc/bjq9KAm4w+LeYI
V1J+qm0bYllgU9/W5eoGEYjpq7Ola4pUg9VVDz+A/ogdU4YHKX7tCz96nGWgI/C2llsYsSWLeIU3
BsGNZo/BEXP0OcHGOUhljst8KySQdsrxy2gZbV26fQqMwqeJntV+WGRlm3bKSJvM9jMusSUF816a
ZceqY4cQBI3gr+52cpeRAaQjsmZTILtdbB/fRVkECbGmutSTk+dbvE4/JDWHDmQ9ACB5WBog3u2x
PDkJD/o+XqXa7ORWKoW2k7UZzMMGXn8HQfZqIVcon9xhKHqDUNPrvL4DTGb2YfhmMLn7E8rI1Wk8
ZjpYtmCuEZkq0noJ/A2ja6Wdh/uIpMoqUZq/qPGpmh9CiCKxaCSa4eilDbjmGKv6YduCbeVqK5tR
11TsUufMuucuDpqvEnaDv9hPpm8V5In9zd0SCWgKVfjg33DMa7j7ujiZFgdni/Xmat36iH2pzzKC
AUgk2GDI235cZEwvyhDRtYgojMhO4vgDEjpDjfd5Eh33uRAmukyLZ2UTbZwp+tNvwD+z6R9pzh6N
UYWeBSUMo4YfEDfYEQW7fJMi1P2fr0VubwRz4/hDPotyfb+T02fz7uhblT0dExRghHO6D03BpLb5
SeufpyTToeRAazFftWagn+buRSf6A5n/RqNwaC1BBkp0wr9tqV1IOlJ0GI5lqJt/+VCEMQoR6Pkd
luJbtpuafn4WCXn8DppTaH788NGHOeLykoL7K9kffMVbX8rPGnaRfJ4rCmo5pby/g4jyWPvptO+i
1WMrUTjH6mrX8mq6e7AERI4e0U/8xNfkFPPqvM+1N5Dl4Sa299qsO9VXAB+HdaXP/XS6Kgr9UusM
gfTwnoQGz1Bd4m+8fKnekiTjF9TLdJ4cnhSs5xpUYB8pSFrDmyS4imwkpf0j+hJWUB33pApEm842
RdeMYHA9jCqPKgNI7I4evF6l0BrlCxqbJcn5DGEFLVBzyLSyKEg/3By1jm1gyryUsRS8pI1q/8jL
jUPpgAnpPx1TeSLh8NXIh+Ab2emtvjaNCCU+fHyc3JYZk0N32ioH9e3ukL22cDmiXnYqY2/PVQV9
iFo68fvnr5tSa26Pl/69K0Fxb4pWy/VE4Vw1TF/VYbfpcoxDhFFOjikmNjeaw9UvOwcG0/c7j8NK
Z3MMyOfkFrE6x2XWaEIxH97vI1L0d4JCHv+SeBk6OaGB4FdMvyyyGqGtxWB+QjlwiTqytLYVzJkM
SbU3dsDLA/L/4kcS5BCX7u69VBSL8fa9wqAEf8sbgbSioyxG2s+0pAmScW6zKUzIcGuzwhm+2bWa
kzGh+LD4Oyk6TsBXavBQEjRILcYJwZ/+jNeFp8+l2OJXo659kGRzkkNocTvB93XEnTC5g6MiYoWo
96QklihpQIzwF1/Ao2ugrs89EFMY3gutqQUn1m6Pcm9BlAuwEVpyVZKdScY5N2TivXIzGyF9a0lf
wRgbmiy5PGS+Tr2X0PmivRyz0RYDJDrlOXSWkyHZ2iru4h8oNPpNThoNH1xbdgybslTkhjLIdOg4
P0awvtAg3H00ADjwNty+tJKTPcs+5mXQ5Ki1vV7/BoARJzhb/dAVQz2LAdtHcxHcIO+RW4OHQ21h
Zjzl+Os/Mb5NkOmYgCRHG6QfSIdxcx+aFPRq7phNpL32zCGHLmKUteKSe44sSX1bcW7GRWuDufB6
+0fWD/d/wxKebZmszMCxMjA55/Bw55+oSTH2eEgOqcT9MyMvzZTNXJ5zK0NnoUPPbCzqpCOkF7Kt
9h41OxJK8pAlo9y8h/FW+puP4FjCWC5YcrijdTGA9YIyCkH0WoX4pLjO1psGN33ybS7+j4cJBKyK
aOwObztubgvDnU70oGBohjapWaqdQ96swgQs0nP1yJQvezxjGVbyvrolXC7Nn5kUFjYGsCK0n0K9
cSifbjnepWMXMp09TxA+evMAQ0IzE5XSXKwbeceIRn1D7aEUKAYeHP0z/etjfm3FGhvoq4WvRSpC
vWUl/x32+ZaGD+eHqjmazaQS152Q3yPYs/Gqqy7rBYhGJY75MO5TehH3gY5ehkhF58ga7//j+YdC
/OPIcvPez2nJHa71f59aOnj7Qte05Iy7IpNL/kA4FgtDW9f0sM6gRTsJG4ZAStt7iTyDQr5oqTxI
aIJV0KuqfKsWQx+baFAefWRQ1RBtpG3e334Y2DIqYt7H8hz4Ar/Y02RoPIshBCHpFbMetstkeIXH
NgW2VWOchKkcVMp0zn6OxgDHkEUTrKDrG6jTa8G7GOnk0XARGgZ2OgrIu6APTcN5tL2SYrAlAMpf
Qk5QuQTmqAfkdTXlqN+FAVMv2GhE6V6E8H5qQeE2M5jH4dcDqYeosuo5kcbWdz1YKXlwaLCFS7V5
3GbfzXxc4Rwe+tM1ZI3DOOW0ehxITSfac1Y5gZWyKF9u1pzlhAANRZhkwsf/dZZn3PTftLtJ7zz7
sLyuQdCHDDupJIw4Jq8xU+szyW/7bZKYjGxa/NxvP89sGVZmOrD4eeTXnvlvuu5UXTGxQrX/gKlQ
ttvd/lBNKxPLgBiMsojoSzL83dtDFS354D39CUv7M1ZY2YgRfW/L8mgzLJO4lzZ3crd9dn2i0p/3
YVoEZ7h8lKfnLJtYcQQaS49Mzhb0wh4prnMp/H95NgcBm4QQ4mrGI07Iv7FE1Nc3+oIg6jZc+kUr
pvVSy1xQFa58ZJ/HPs4tN+z4WWg7ily2S/pQTY+LSZjdkrmRC7WHCXik1o2qxDPc7/2MEQzbtrMn
Fvr+nVw2aXGBtWScSu/t9YEUxy7SW2YdpeidkILEZ43V0DzZdC3IQf7Etww+T8fHOf4q5QBrenI6
gQb6PcTBOo5P+iGCZyvpVr4H7gb/1I2Ee7z/hKudYK9I07RrOAnX75F3oihTXyPLuxBvYulEhebM
cC6QdZFGlOyh+7RkcYt+m3A0jBPJHqTPYuoNWd2Cv8GkYuJ4gPHGQeh18ya3CMb7xVzH93MCJt/B
aXULsARgQ5I+DIWfQFs2/WPo1i2aNx1/+vh5xAE6eqQRWhAEA63Q/PKAWzQFedaugY92Y8RlvOE5
PVgQaHRzEqOmRkxWRgiQB+hTjS4WCqcW6F/1ZZWClAMLoAnNDaQNl0gHUPskfTgL5C14Vd7X+s/4
PKOzlYkjHn0J0H5f1sZhJOHYFJyyWB0F9/sVyZtwOWldURBWC5giwvU5zdy21Ny5QWdbNUtAcXEt
ARQVohAWWIn+ZJAOKIJ1ohBtp0Vx9auKxxIzBv6V81NSOcOM1VmufLM437k5e4ODHARggAWHlJBe
TP9tSYbGgU8zj+nXplfzat/Pu9DsR9DXcfk6VahgsU9A4W62mhbrIHKVTP9gU+ixCkXlnW6UqGfy
yUelaPGq6vVPIZs3yJmi+dF62IlP1x2Oq43TCu1WFGw+2EIBJBFVjKiOBniCJc8EB7lfmoRXVH8V
7ssK91u4VjEnZquKkqKcKFC774uVutLLbWzzJ5SjSyKQKo6SQVudkDDh3KPQyiiAIxeVxdyvuUnH
SCAUH8qaGmFO+SKHHJ+6gUk66VBgyuO2aKQ9rhtpsz3TJw9g2WZxcTNM0x9KCwuqVR8VvLCQDfGe
E2uP9z4lRfaYrbAlJirlQIcwZMDfBKspt9GGuUfTWd+1z8Kh3fC/Zj7nKTzBCAdS1UGC9x7DmLEG
pHznKzhcF8KgXYAxQm7D25Eqy+2ZN1ZeKu/Ml7dyN9kYQvFT3IAFr/B9jHiCrnhUlldhkCXY6+rz
w8eTZCDjdd9+GPPRSQVEROwmZrrpCVh1B3GzaIfJqlFLeby5iN0npnOV4TCd+jDfUa6AyYLY3vpm
Swb4z5A+yK7MbqwoSTLK5rCkDq9Dj3FSg+83BTF1rg6bVk3RiA+s3G0ESFvVLy8doD5WRc/zFEe5
d6EudgkKu1X61G1xZ418r5LRttSuNSWywbDUwPAqPt11I31y3IRQ9TpJcIoJ339vUgoKdoQOWjAa
4T6k4P1MyguAUXbRtP+MkW83ogiCM+SNsse5daBX7zo/axkWeLpirKFak/jr0ZAVieVsZMjPT+5v
m8tkJFdWf3mGCkjv6mZZmsMY/pa2SNrdy1LZHfbFKYrjUXe8H5P7BvW23ow4zLz9VZJ1tEbyDqFe
Vx6WBFQ/hsDjZ58GR5fD730xPQQo7kwRzs9yN5tNrDLusduHY5VyDN/HaEIv0PRZjvzobgoDreyJ
xqnn5aICtdaQM3ehrihZ1B+cI/X2vlIptiDmHwl+ec7KybuxdILBojf52hcS52ioW5Eb8q1GcRLT
k8kuAtZLsZCU91dBO6I+d0oxIeJ+4c/CICGkmE2SHrYxJyRxs/GTfFzYC9MlVx25TkaPMXuzERNJ
sEERASg8IRhY8CkyBKGyqnF0sIvijPfQPh15X+yrsxN9cep1ZlYiZf1ZaCyciNQE7rlK95fAAOV8
j/fmwKDrpLsFuh+XQn6t9cXXc2DUSTTWnSbsKSFcA72KVOGOrgzmSafiWgqmsy/FaDiGMiqeNf4A
yF7TqzJKquDr1Bio63G2yPZY3BgBvZX7v518iiCiHNsN8wW5aWSLeTK9pvKgVq14Vck9k9WRcxwB
ZpRf8E2yUQqd5IZExgUUwXGokOXAJI1U+oT1BCMOk7DrmzZ5JJMJ5VS8WJvjfzpRtt4/st+8VfZQ
AuqEErnv+J7kq78fLlXn+/2IgL/qniC3Fz8LKLxm2cLI3b7zx3SLtoZ3KE/Xi38kazK1r9txY7k1
zV3E+7HWHRHexG8OLmu9bcyQlxSvk44MU5svIp2+cnRm+cm92hgfG64pD46pogd1hYMqJdUH38E8
0ckqwvcqhMxgccoLcVHTNC4sPuPg2kG0PeGGohE4+TNZxN3GrJQTl9TT7MILxHxMWlCiWTyNYZG8
xzvBQcGq1keLV/SPX7qg7Wjf//UfFD8lZXRHCtsXI6AcuY7/Fr8V6c3Dt7CuWEcZtQl3MaPZgde1
4unHkeDDXEZetwhk0/uoPx306DS+C211NjDSlSlLNYzr+r4FElZKMWUv0H1tcUumr7idDv+QcM0i
e52YDdDXbfwng8Zofqito3jqUT/jr6Y8FezOSrMtkweui4EhViRmtEU9DcvwqfV4oyzyjz9SDpBg
n0WsjI0/aeD2hj+Jm+WmHjMU/UYR15rWO6iw47VoSrLXF1T4pK3TrpJaT/62mS+SJ8sU0CdJwx+6
jH3TM5mdm6gK7f4+3WPn6EL9RNLUkIzbtAXvERSu8GAOt6pTvO15fUi/pRspJDBjHRcnIK9r07Uh
4BeffIKmrc6gRXy2kmYi93p+X+2LV5vVtg/Z7sne1agDz9C6F1W6CuJlM6kdTT7qoR8SFKfCJPfw
fTYyS8YtlbsnECVE7gkLEgoY60K6sNAf3cBmoVUe4zM7L1JbJfn549vnG5WIcA87jbsq5cKmyOIO
ku4a3qqDAXryevRdXak2WHZKOSTZhoI1eXEGE6jxegQ4ixkMesVzPJUXXPn7z+GJ79Gjo/TgvThE
hX3CpTAmbyq1R1PXQyhppHiN3OzPcwpx5u90CBOMOHkFRSwdj8Tg36Oo3OCUG6cY7eIVn4+Tkv8T
If0kpOKrVTgm09gdUvudJGVvDpW4UJUb9alySyGbU7RpYJMus7D1pJA7DCpfPvsKGurUmXTkvuFK
4+6ESpsmwhONKLXMowUG9BkASdK6vJMCxfXOXJO3f/vkB49gBRmQXuie/j4H9mqKm0QVXKSMooJW
vHUBo1G8j92AjUJ0tSrJgcZ9E/YE/0VfyevFkK8kaMK+Jx/ObMTg4/8FvfAUqs37hbhMpXvJTkJl
yI47uPPUDgru3Dg1bG6WjT6ACJ7CmsmutrCI7gY78LVZvfnYbs3LMIgIddNvBQE75IaHLv8Occmv
rR9JLG0ZwOImNcb1UF4u9Mn9PJxrRgXEdFj3h76qnvJKp1FgB+fUTHiPNZ4sgQBK6YwTB66Bb2k9
D4ecaBhfMxUMIAIPCtApEAfJIpqZ0ELSht2uHugV9YBo/+Z105yJlRzx9xG0rniW0vhaQoBHoYr/
mdez4U6jizrviRkFAoO2+palBGe3yJsvgmAhOMvWNF8jBP5Tqpc12uXtfcLpwH7ptcpEnJxZD/Ie
FQ3mAv42c5DOrfDiv58wPMtNPdWXAcz4idIRe3CxrN9Pqv1kXurvH28TChdkmYA11gbI9nv+zja+
ZneFCD5mH7Evr5+7oWEez0oXr6WtzJFy4xJra1hkvXVmzPoCAgtOSrRyqeTU7f+TL4+QowrJsFWc
e3/VXB+xRZR4wljhRH1mST0e6DHAD8sYAaYQyZlWoF3RTsXwczsrxSXC11/0QhY9hf462LFh3SEC
dNGMNpZF970gFhLRdI4q/FG0lQOEQqiMHcmS1xw82MYW0l9bhKLcbxyLw8zmEnI0xL20Xm7oBtvY
QBLbMpAOk92uKIDEox9ZhpAtdprwpDw/UsAO3VsfGpYK651+osDoP5fsN/zhwoZ2dsvN90iCiLi5
0RVdO2Spmn4mgD1l3bium6lTIWAQ3LpgQ/OzXeU+r69fYhipTSsPaxnwRbfRcK2hEeWUEGL2cuB1
/Tpu5fo37j4nPqRBPSM07CaCbyLK3ZqQIRoVv2taxoULHc/3SOXFZlAxIflcJnwdgKpPZUI+9Jk3
GfbVwC5QChGCq38vZCOlODPTgL4AUeOEPiKQL5e3ZAtr9hEo/YjoVa2ICUTgpIZPi4T18iS0KEtE
/gVCEAYpDQszYGVJEZ341Edxe9RA5QOU3R7RUSLf0KtKwMuAThrzWpy3Zlmxi3KBat0nTfOx1E/8
e2xuajLy3yiaMY9ULOYOGP9JSRiMigNHP9zcaWKDb81EXWPqMMDlF3reUHuvv3riapFYMAgFMbSn
2UTmppWslYdcVJSpCV7OnM7M0ccdGy+NkU3EJA1F1hGN902EqyGjziWb2vgEsD4w+dhIcBXpGBDc
o8YZY7gLXeZR1hzkVpzOTlrPrGLfiRhn3mrqsv0/Sk8WvCJzrjw1VC7Yxx90KXWN6EUxK93rfQ5o
SC9Mc8cgDxDWp1Bu5ZIGykQNB/cCH+2ZUVnDXqdojaCKydcr2l4J2fXYBjuTEmxHkUqgDKU0/48C
4GrbSWygssiRSoGaGbKKHx6Imu+hLUxJO4wCtvvT6DcFaOLCyJrqmbex4ZUZuRxDoOJ7mwhrcJXt
Yer8WRGZ0Zv0AAsgoPTa4JoNea5njjL+oyPIPQqs2blwaGgrsmDKz3jGZqmbYEnNxOLqdJIjk0QI
1aBHCD1QWxgUGvwfLXC/DO0bVAR5pcwulXM87NpAlSY/NX6hawQ4pFBoRtwPGwmnLomPYp1ADCj+
FvrE+2YVfljjHrr5nyFBDEuok42wZMuw8VWZKDbOpEvSV6S2/lMJ8XQ=
`protect end_protected

