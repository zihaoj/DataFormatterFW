

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
b22tRkeiupS35dek/Hkr+WHJ8ZMw5n66iwDYOxpZOA4pMaDh4QW4WUyNRCbyS1nf2GOGjUGEz8Eh
9CM9L/D1PQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QmlHIUCUQnQnCGdP5KuuogznuOT5piwQJTGETTKer4fvWEesY8KTtUUhXXsXG0EQfnSwZEEd+PXI
nv1bGiHabL8eH4t+tzoO/eQJKfcer1rfuXtef+SODtC+2WKEJrEExu1dnhSbmobF2Q/1pqkxNKJf
pVnNjqDDKVdVrkd4rZs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HOH3uQt0bFlggIjU0Lw70GBBUXIJmuvp3qf/6qEU3B+SnULGx3XUPgSqTmIT/Tq/VtZizj64jEo2
EYCYh6wt393WkhXVvM/cAIt17OIfwsCoTQ5XsM8q9bNU3L6oJdmr+4ZMPLZliVlCWAsth8o4J6ht
BEqlNap4dyIZtGO2iCeAT9DK4QDQIi9DayarWjGJtS2oZpFWTc08Nc3gbZ8E6LHDyxbXBrb3NdiB
UeA/aqLM5ohBTbBNyLEZSDnnBm0e3xDa+Df7YgRFa2enWfKdr4IxfqP06RSHdDeCxKfy9qIvFwyj
pAEKImirk0HZZZbDqULePCLm+rbCzdDlE5JnRg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b30Vn2xdhhzDO3Ryt6KVG7VoNpzw8KYKUvhTeEArFERmRnGS3mcRpfuO9G8UOU4lJlmcmjnGxswR
VKN186Illndl1jl3rSr8RXVOVRZviKJ7A8d+LKG3We6R7NndLmdOyNWMcB21NnAnc9YDBgJF18mA
QY/fS6fWhxo7wMkVGXc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gCCdkronRD8oFjhdaX9depvt/0rVX9g246RNh619xQxXLQrkEtypLcbwpRwe6/0AwuEgsBGvAWON
DQSRgbagmijf+5YLz+j2UeFr630i3tUg95eRW6RJBg3Th3K195e7zqo55QzTXzkST9tx17ch4NGW
eqDKAesoNI1JJA4KzgFtkimvHCbw364nHqR3bNe/jyysj8uWdlppb4NS1ORCfBEbEQxiHMdueRI9
LIwt5m8VtnwY7kHA2ieY0x/mYWvNY/cwQm0HyldrMxcfI5363pVRH8rAp/upI2lem+EbbhQw8Ywt
MDdGzoUDUVgsnrHb0ZZlcyMGD8iBWQuxGwDgiw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4192)
`protect data_block
+l1k83IR1XP15sUAC5W2SMo8R9k1H/sq6vdUWvQMyEvQrJhFRCnvn0b+QkY5XYHS1IxI1m4ggSGa
UsJZWogy6pPBxxgJHuDHgZJvnOirkfT5bDGJUXRQFXqBfqyAj6DZABDQm7Hsiuru4ty2nLZ/XgFp
rtTGeZdaTaw+GaLdG++DmipQ50yQdYLPr2L/23VKu4KXjTn0Pnze6Vg1M27sRO4QthGtGl83A95z
YORM8Lclt/C+MAtwdb3P6t63ooAIns7ri6OtuYyXxlBrjyJ33WB9PK9dpkzy4z0DNg++IYVJM/pn
M/G52XM5qYKA2c3YOCvYIJhEP5FB7dStfr2hCsClyzu0ZsQiGz/Rcf0QbqywqgEdERcZEP6IrXqm
3CXnKF5W3hfR8RHSZY04WIYj0QUVQ/FjYwZl6qv5XFvngipHkhGFz4CfIe30KrhxtJ29WSSpNtUm
lKGt8lOz7hs47xbK9pV3G8bSd/nRFgs44oFLbHRR1gOpZm+v/zONeKQgs0fPc0U5RYyytqJ96YCA
32CRijRN/ev5l2o9dKCw8V0BXVoyjPFjK8u4w+Zf+ya1ldKgbVNKOPor7vZAlXuLI5/4BdlAjUzX
3sgPNRrxPaaiyx9uTqunMSd25F4sH8ibGcdKp7A9apzGI7WABVbAc7dVlfEJOukGmyBPIOuu3tN6
9O/PuGVM5BGehpNW3IVgM75zMmv24EO7Qm8QDhwXuqu/7HGn8uNGScEo/+7rHJReBzwlz6qgU/VB
AA88XfI+o6nB1XuPxT6e9jnjXz1aYhdA0tQHqytmI/6Ulrr/7xQtywcPB0nvEHTXlPBnBd0eAMUo
lQUOGlBT7BmGff7kxStPRXI5h4AqdpSMoEFSsRcrv2/TZ4qiZFVV/TKChApNWqj5bytzkCRJ/jS4
xVF2J02Byios91lF2aLj6uDFGHr/kWl4QRJj1BGnO6Lr7N8FIvyxQMGnUJ+9CItpxiaVWdRKyDFx
X2nfUGYQjyRTSDrbl5AMKXGMKPs1Y3hnO8cTiU99X1RhtqEyk75gZ5z2RKAwIoRqETtoGL+5R4ka
hgRXAiPmNhGgZqgbeXEMyDkS/lqURjphDx09wNKWVxZiXkr0wSl4CXDxQrxmIZA6Z74dHoRExhH3
1SBglrDZ69HdPL/UE6OJ2NIzkOJH0JMWGVl/0K77k84F/z2+ha0ASMgyHpd4o2MDw43FlJiqrdj9
RBvpZusmlg3N0tzn6QFUWd9T4uHBFBguwGVQGrQCggbw8/XyY0pbUlbMkQ5p7XPRLEVD6RQOKeTI
RT/D+UWdudKT5PcbChiF3OUYX8ZZ+HqS9JoXVduQj79Un+mHYFB9wgoeb8EKXSoPaSaTOgj5xycv
JwH+o/Gtk7Ox+Z+ErrqGBMC+I+VM6RRg34ISmQoV0esb1gYlVO+0d3t2CUZsbDoeq+NZ254gqYJo
xp0r1YMW/0PATnTVYv4JIGMtv+6lBnvZzP+KLnguZJsK7OGaNDJIhP9p2k0unFJMcwZRAINVQJgO
Ackq9wb+Eze9yrkq0ArbvmwsZxBfTnbG/eR67/6qH7Nq25llKT8LFlgEE1apG/YYj5G60DgFvbqk
hBpHOaQPAvgabkMXxiyKjuHtej1yD5s47YBDDyIqdlV37VCnPpiL4YgU099XEdLvWcgp8z/msTL8
pB9N0MV4JAz/S+zVh8JJ3h/gB+ofZbCHwflzKtTrMJFhSBaHB2xtwDo/YxzIjO3c/Ky/cVUuUNsQ
+OpREu5DxCN0CMFg1Ptl2D2XKHYEUadGrBwTKdieU1ZO14rPErEC5KLbBQTlnfKzUC/cWkvwMwuH
BA8zJsQjwlYOJ9sS+S5ImKjJGYFW15LtFc0mnbBLdt59HrCKggNk6W+0vlwPGJSjVjkjx1OLkM7E
6wkzuHyKX+Pa6hIQMX2bdoeoYmAQbgw11y7GwIlKMFLRsn0zqu/NDKWnK7vwFxYJOr0v+mx45ND4
+naR77Yi1mI2a28+0MIMIab8jc8byXhoaJaQcOHtFux+fUusFt8kKkfeyjOj7Zvmmq9TZdbBoZtM
PkP4VEfB2JjjFvh4UP6xqk6GHLl4agf8WW3LbFDvQZjT+Zi/PrBpp6/yy/jHRyeoz2EQ4sw0nmFi
hsiL7uHC2OY9TvbvYa63WZ7AUsBeEUHkASi3Nc59iSdnQvrJHB1r6cKuJ71UlQU+J3oOCIg1Y2Hw
7bI4EOyyUZmWYqZq7BcnIlaUedXp63cos8gIgB1R02rUt0NerrXY0AesIXKs3ZtQgoI6PeZVQb7O
RhSs0Lg/tOUltD1i3cvTjpWRYpxzi7o9+VNx9xJrad1ci/JxR71UIrsdVy+rn8JJaGQcHmEYSFcI
eg166bAUAEPYz7N3atWEJcuMCSTOSZfViRsGCDdkS3zLsHrMd2asVp2qpcxCQwgVQAPUSMH1LlYe
8STjZ7z7bbATMEeYLUtXOnvZQYXOtIuaWzqLInlh1MEYbhhRr6aR3fEUnv+AlKq229+yGMvKtJ9v
RIPvtnMMHUEL8/v/8uFEWrJ5uOl6ivBljiN+S59NwPBvIt41LuPbn39rHkMwpDJhaPJ/INYYQdEE
aVoOcwQIle7vB3EnGJ/3FN1Ij4WC032z3q/u+SRatcXjT0HX59Hs0NycZ8TTxKDIxVGKogP4AF0q
Yy+6X/yfOtgqXPG3DQ7fqtRqx9LlG81geNL62vm+7ACRxU3iKfU/yLJ33URAvvipEsnHkJhgBqqc
bMnyAr2MQuLo6pcLGyE0hUpjpJNuTcJlmLZya9grsuBLUhrMG0IjfhaVUS2/3apdiwqTnpKDqAUX
0xuL7pw/sH5B9KrLPnJE5yyXi3Yr1rXNRlg4VU+cdO5yLaAsmJgKvoMmeDXQ87eIMxKwnBfEAbY7
4sW2cwSb9mUvpTCkGnyoLUKBlXiTFilwEy/gCvn/LAtmVS1+osuLfJrKchAopZM1cNe/FfOLPvSx
wRpYTQ15eCJU2VIAnOfRtqBn5Ia1NruDSm1X7PTfGbc6Z3s/IoyThAc9A83hihSzGXxKCqNzyAjg
M2QVZv2VqMPuFIuhPKZb5cPhmRjHsiggRH3J5cjPY7JhU3JDUpA6NoW7L2Oj2WoowL1AZohtTSFF
c2k5lNznoJCPV5d248yafzXFtxeS/TY4l76cr1WHGYVCeJ2xc6sXpwzkw3rk8fNJ3RWeh27NCoOL
kSXUEr8de+53kKCgPLtRXuvGuqSN7Vh6m6UM/UQUoKy91KzxzucPjA9BFtGoBy0UQQZpsk1BGXVy
zrp/jGhpbKXOfEnuZ49Q/hyQeRJlYJuEbY3ekwnja97d3rttF8wRmXWoR7UxAkniq49LHMRScTON
YOteXNMjREiOXGKgcWLs3XKyf7EsrpNzKD+M4GIpw9r2LrHgk1zK1fYKzZggx3g1cPRzpx/R8MPG
vmvsKMzROnoJBqKu5sFTCIXbvjHvj3vHfu1HcuhBYCo9iaZKY+8ixMABtKz26cV0D3yOsfDXqxje
454en9wGE8akSGHEjk1rg2nF6iD5aB7xGPBo3OWpKUCCo+fvQI3KUQcXxcNWWUjduHUGxPVjrA02
XYK7tTdwq0W3sunRisJnkB/87eTOvZqmcn/U0iafps58mvreCaujM0a2VcQ1gkCWTPOyViHQG5Mz
nMZQ9YyxuwCbiylzTEIdLxfvcvTrP4aHZuxqB41TXk2gZHyutsdr62k4JJ6skNpuWkdPu49qWa2R
OZUVHrklD5R/XAA606senNiEJxzk635wVgFUWv8Ln6M3jq2PUXsSQuJx4ppklTfdqCDMrqrFu1ui
73YdUuKVs4xd5TghrP3qxxufekkfQH0MEfu8WKQHuqaQ4cWf+5+TmgdSD61wBUShyPZabt3EucoQ
e1HeY5ocecvQYaifTErSIYmcEizPYofgPR7luR8Qi68QTy63vzr+V0TR2uEF0/qP9+to1MUW4ftm
vEM0i2wiFjXkQYNDfMP8+51MRQqzKUc7xD6SBjilrhjgeBfEQFvjTQLlC7AMBMuVmU1wowg5LFmx
pp77uAGRHb4KoXE+gJlyk/2hHBgcHZw4E9fkN0X0QUdH17veV2eP3Wr+ozDdHiegvCVM7KueNFMS
dPlE6arQ8XInwzdK1syp33Oj9bHZC6wf1xVS4KHG25tA/Bm4p2vb/mqLR5TMZqWIF7s4f49sCUWv
70xEqHhOsBWYcdn2Ml+oMNqDgdK+CtebvmWRxpbRdTHZTA9YXE5tQcPrWXZnPG7JE2KiGLNjNh5t
CGnnj5Q41cTTWShp3vEFPTPzGn4PvdIks8JMeQBj+dwmW4V2ExjiiPTXSkZ1zSx5Ha8bELaVHX2F
UQfKRLne+O/azvJ1jjLCVK1AvNrmZ47cC1ddvRDqSzQ0b46kkIlJUfQem17XHu5T4001KTMpSaDv
FCtUzrjMhM2gCZUP2G8m4VPv3Kulp1vb1teS8A/eKdAWJyKk7C/PE20hNr0w4xfXOg0z/WdrcwWU
rH7q9JZfoWXZr1bsvH8SKiBT8wB2gdXeTrACdfB9VBpJgeG3lZbdg0cXyOiDxPKtxwDpwnZEP91q
p/06r2sD/W4ew4+SEiRhscLREl9pmVeYfjT8ZYi/ya7pyTze88QMPmDsFJvNH5BYYEFkwLu/4R3f
LAPZyBzRTQxtg2tGwSUtR/98o/7QJH/hU1Z3wyQXTm76xnHGAxKC2LCa3pWb0AbvXhvLFoGwZbV3
9ZoJqjr2QW6y7I5NP/RnbyHrkR8xFHLsW6D8m1C/7rIyxYaT4LI9bgOa50dLG2LsqYlclsmOFt+B
QzrpnzdlZQbv4WMbfMg16GRZ5iEVH3iV3JXXFKyx7fiYH0ypBWaEVNssfGwgLFexBTRN3j3ncrNP
6VsAQnmQDNZirGsxytabWteVHWlWq75DWCc9Amkdfi549FkaC1MQ4uAhF93y6uEauMHAvOyPk1bn
Z1jL7nQ2PsRTyulbsEu3yF++uaOapuujnl5iHShJajZBk4EdTFTy4/8JxyPJETCHBZXwLQ2a7tdX
w/yU29Z4KN6jaqpVM98KgdySsxEijxxx/j+hME/MivN69BoYongQWFiO5WMYh5Zvp1vyhx1Jcbs+
yf6jofy0ObcINYAadU+L7gK8JlJGvFmK5MX5kAdnnSOmbP+Sl87pXeXLwuDZDYBD+5f0eW1kH2B+
sBV+mMF3fQLj3otAyUaRJMkY7rGFTrMC9LP5MtJ/rHCTJex5hRI4iThubKcx7/X++WOt1/Yk9rH5
tLSoZrXzdaTYODVMwHGs3sjwVcu67wsWwRYoxdLsvdYlXEiVW0SehaFt9JS/i5F8dTKALfbzpyG7
/fPZsrYyfVux4I7++1FimbymGZ13z4OB9728kfow0iYGjVCXfFL5I6KEr5O4InoQCdJkbfjzaHyG
m2cO/CU5crZwAlD8wgNPVd00U9Z0hAgp2lZBiPrfJ3AI0Yz02VnaWq6yJpo7sei0wh7CYmPfK0X6
eHkECAxSXtYRbgSrCRoY+pdx2Zu1qEXFSvDWsO7IDbjIQQ0UG8FDoz/BetGHNaqZhPHqXsRx2SxH
9hMDHpisZL+bAWhHK5IBnWaEAgaeMO7oxPpfrMsEnw==
`protect end_protected

