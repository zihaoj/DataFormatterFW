

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g8r/7sde1iyR0STftzcYOcdH/3R+q3JXUCZQpPRz/VObMWWqrxZsHW7lLAXgWiq4LPjiaWHF+vPi
AECUpOzjEg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WO7DgZGyzsVW5LpO/Eo3jPkPwTvvisAARwFpj2ThVqKHqWqYz+cfigwxmDVkJRua0WFfWGJfALzZ
wH9inJ1f2CNVtaotQX0lZ5c362qhx1ui46ZI+45doxR7KHnJYjtJt0bjBJRxWiG1ibF5Ibq1Vypq
pWOz4nlaE+qETERLz8k=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l/QRLOPuCKHCQg9QTQMR7jaNBVIni483AUdnDJbuUz9G/TnesoE+ckhte/F0j4T0BnQXltD2Tnpx
iVDzBTduCY+rrKSf4BDtqZQWJixR7872ZqBGdzwwbc3lZRFia4ykuBaMAKWhpB3egOY8nll78wm0
IlvLFfiXsSWw6JaF5MsY2IumW7cs9XxYvVrO4NCsL96xF17E8iSUPKLB2HRiNN0435RV6oaVGuFP
6dDpS/axWCBwmIlrR1/AJYmARBBTb/HJMKmuWtKGLARg5e4GekIKL5niXM5CaBOaK1N2RkA9p8cv
1ZaBmtz4Yz5BlqinZppN0hM7m21yUJeY3vk0LA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SIPc+Pr9P1+9JsBFlLDSyhr56wAGsokSTHVRjBnYtNQRv2Cm5GaMw9a4/GZLBPH4gUodqp7zeOyV
CWSlDOlDpo/32Shb9Z69I9aAKcLsfexMWcoMotgY/7e+Q0QLV7cYrd/z/ObLMAAUU5jChSdYnzlS
+7VMeKlMLT2qVS51Zgk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Pasliv+gc6ueSrwDi8CYMLQuGH7X/hw+ACS+RP+c7r6sIaXZM3oFjtvI/1vDkQwJt1DRpzLcGPpf
nX1SRapBAYpWFD/ImY3wBJ8C2f4pksIHaMrjA1wpWFNCX9VFKYl/zBBBB3CLfQ/oAH+HyUHSfuky
Q11Q+PE56TbXHxVkPRT3n1MMU6Dz1GmFhKhauQh4dtuk68rUVbIj1iVkOAV/24pJz11QsRqZTsaY
omz9cQKbLN2TrFSoAkUJgbRAynTACbr8zvFgBQybG7Ha8oZ9TmwUMCoCzJ51TocJML5Wa3hez2Gv
PJVH7QQFGyJyKD2iA/1Cm51lM15588DZ6VeZ5w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fitjjbF+Uadig+MOn0ROwIXMOGmAsKF+ai2aPPzK1LuoHEybEUjV3Ow+S4tCN3XQ0vXQwlJ9qrkh
XjAxKmcndINrHSnUQUnxaTr0eUO3vd2WqvZ7Ju0XJDR4+PjdZ4oM1DsnXl/hmdtnOjsCyplOs60m
9W9MbYlqrIN0NheOVo+Zaea/RQAZCCYgUcu9j2btQONsOmorBJXqpSvBA2MTjrhGQONrMBGpIptc
e9X97HPIpJ+DVROxngOntMcwYa41rY0znA1gjAtxPvzggRWl9qqUkQqmAlth9BjTr5K+UBTT1aTi
YdQaO4qgUwRsHEtK35jViPEl7DIlbfQ25Evt2A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4032)
`protect data_block
Gn3q1/b6Uzor+Ot9pFP8ZeQ1c8jJsbmmDWH63tY2WsTdbvhStKOG0k3TZCYT/eQscHrs721KphDH
AQCPS8WOXatoW7i9qlqt0/zGKJkK5rUacEFDYlUK47lNAt5d5bSffqHhYdbb/cOFB6z5VRy+zqAT
zYjSA0akdc27aABAPP5byGTF66vBsOR4lnD7Yh22MFFCCjMTPh2BAqX3jnmsWE8yLWVzlyiWTmb/
rDOVk4bChqGT6Qx+s3EySvLEY0q39VAO2757bNzlWAgQqd4xGUENd/60YVhCbM0PVCujhM+Jy6fU
1nL9sbxafWGJy9ignToowfiiOUUQxpdsLO1wouMdx1doFBJHVOo7Wtt2ps52YHSnsfXxpoPeOVP+
n13/bbCzeTJBm3bV75LaE9ZdRK1w4cnEkpFysFDlbXwWix9929kjdBaCALfLkVLRLe3VpAOVH3AN
Q9grHItOjx8hJSfpPKBFVwqv3Ou4jD4XxQJSEUcu6xSdZxUCnHRuyMCAtFhSsz78Spli1V8mVkQd
X1TPKtKEgGDkJtRLFW+5r6ae95nDOF1sd8o0jSkUR/FaaA7xkMbB/eO7aby1dlZ2t70vGUaC06sT
ep6gv+IRKqGoouAhINau0WICMzbopMvjbuVl4GtwkiJr0Sc5DYxogm9mfeniCaSCnCNnfuZQ0mKf
jhJp+M5oz+iM4gN/pMFqgF9QF0DY4SFA/U6cuLEq08b7N43rTbSgoNO52AuE63LECcy6xBYF1vsM
hISCKJIeB7u5NA9BbXE02HngSGnTAKOd9dLRMkttalp6n5IHK3cuDafWDuHTQoGlbMG9ZcdmTaGt
5Ma0/c4BCCVZdgMlaFWkJR2VqroQTk0TkQOUNq8dsSmN6TRxdegGbjp2QofRvwnRWmn6OhjHBnxh
Ba0ocq+WukrztYmIWa5VmCYhg2YmjtO1KxI0ZTFmM/74Kn7xE83YaOoxgsihdx89IsKddCjulYLM
d6rA2kq19mceKjd/4PI4q/qc0Pdcb69OTWpp245kASfzqmc78ag20flZNuRP3iBGyp0ui9xHRm7R
HFRObbCfb4pz4UWffe+8I1xXVIKiD8LjHrUATJcB0NYetFm4vu+mAwTNjPENfhKc0zVeBIqy8f/P
67JZ2XImvmrfG2fl67MONe2an7aUXx2tOebUVANLuv5xsyn9KMxF6oq3BQqgF2Co4fb32QrOW7AL
YeY1xm3pk43DqtcPyKqs1edDiFZnk5oSn/FlEtHKEF1y63g3iAd3PPdV6fOLNHYDS0DtNWI7ZtVv
QAOZjgsjZkdy5cJIkmQTkHqplEBwxCm/UHD1Htunj4lkPFAi6l+1P0tVljGs5ujiBkGUwsUpCUh8
nqYmpDzq+xh6WmXUAgY2At8pnlTmONv33gmrJqam3WRKvSyej3EoYpgeoH3WCBlC0jzANS65Y5u2
qxvz1GE/Fv4WofQ8DraS2Ja6cdlhKCugeIJ27FFGYZBhe397MhUPbiaYVi8g/6e19eE+Vx559J1T
+IVXSNJEbLbde0CP9n2frPXXGGQUvuhesj/vUmfwd0q8uMkzeTUwg2Jtouo2ymFWxlthcxwavuSp
6ba1q1ZPL3W7bOmyEV1GaP8Xb14NlLKDsTuup5ibtxPhJgdkcWpfQ+3Be4IPnz0X9/rNwZdzmRIo
2qrNMEV/Zut8rieMbgtNoD324Qob9Ttb/6KFAgfw9JjTgawcqu0w97IBh9QAA+6OOETyC1Ibf1CP
2Gsf4qOjsjU7uiIazednoOLl0MyzQN+Y/+MkFiiovfQoTvS0ywvDM8ttvNKZYY0ycGISzZ+TC+e+
TywO92fr+tksZkTb059ZbIMf1rjSKc74PdsD62WI1jGwOwZGOYkFKn6U5W2/KSyIv79+eSJKjyfx
3/ta7XkWEWVFQ5TN/H3o95xkTUMwetgW3Rvt7Ty9+QTgnwR65DSpvq5lKSLiOe026l9uz1wBf71n
JPj/Uj5W3nRHmJI53TDlUJNjoKrh/83bNVVWsJ0PQdgLQz7PurB+ZjhtS0IqhJOc38wm0zTY4/4m
dd+m3J5+tGSKolXOMmMCqMxdF2ry3lZdoLjuRVpVylm8azX9aJMIDE+8hTMhCBbiTN+5oRtaCmYs
fAaOc+6ccpL/JtaciVGl5mfAs6JkMCyU3C8n9C5GBP703vDr6mW363MY/gRK1QX1vNSB4Nj6lbWo
r1BoZMGeEz5Jy+XIIIyg61i0OFgTgde1DHbDMc5vagV2UhbVy3ruOfpfnhZdveiLchVVh3Hrzab+
hCG76TqxNdZbw5F2a0a+I1Ipmb4ZR/4P1fYAyMiX5nknqPSB4t4eaDWcOUIiwJVFdjlTPQY4VEVX
7N470X0mU15h+uogsRB5r9I/+URc2CAgIxVI70SybjEiApd/D1lUcvlt/r0R3TLXqfJkMkE+grmf
Bd9CgT/gO73cPAB0cN69EY5kpq6pIHPA+tPqfWYMR0yNbhLkJ0O2dXYJ1uLEijvUZm/M8+GWM/a/
78YLIApPXp+fHCQdEM9LoPqhMAEYU3vGLOou8JBm3gJitBEp5ikt46JAPvvSwpBnrB6JwEsB8O9P
8YZGakudC7/ruHPFPF9cKtJEMUPH9TvPm59btrnXNlTZ9Ev7TMQIDqZZL4hEG6jpgrd1eSgNywEC
PTS2rjzjXEOMiMNI/RjliWG5fpgjEG9KgB0BwiSnFCfjOvHXpvUpA0Kh70YLTFh1mLG0/xtmXIJ9
FL7Qj+SqlJzuqiwG78jNPIXNFvlVAPVfA5i3e8FgQ8Pj+EsOHz6JEGXgyFbWM8MUsI3tPov+VAmN
2S9DJTIghVfD+gRvsyAYhDC/dPhLvL/1aMYn+YwkNA1n+Q6X6RoQ8lUvp108rDrNtYdF1Nl/DAk9
r145wOsqfBZUIh738XpE/TiXrFihbqTFpOKhAZChrF28QJ9p3UGZSJMQB1mZz/jBs6bRn8w8bbGY
2V3664AN4J5rY7RnJBtZp7X3Gt47y4HHDUfJdMkYuZxQ2UVqTxn4x2+sDAdodW7QXyzeiCZcCo5Z
1hnG8MYf+TukH8ad+eDX/YtUUPVjaW4tk5HGHS6cfqYBcGecwoOORxqaLOh6n6znJ6rRDyhltZ54
25qnR5pnNG5tH1SH52y23WNLqsyt2BAaPrSDiRULBZwaKMOgrysFgso8L6MCw6/fj8wl0ktDYomX
3+FE5wUWxaZO8r1DyP5qsH8jaedx0ICH9iF4VMyrPQKB7q2lI9QkdBLX5Fv3XNFJ6AFzzWIP4wKP
EsKGn2MkIjoX8Qj4QbMNeYw1O3LOwypFWv/fhhlH83rhhVkh+sEde9lgGWrphUUmx9UMyQj4VGuf
Cq+EL6Lo3GNCvQo/So771P8I15ErEOmJ/w2V1MoIDPMJPcfoa0pHjxxR9uGmKEk6mbHzoJlLjSDw
8HKrHZbwSGtclDBkwTwaGG3q2fmeqU6O7NukVtq8jp7TqmMvJ9rgOpjucqzZLT+56msSkNRDOapL
/QmULvsiXKulfoBQCQ+yR7UU2dz3SiUHWlUlY147K3GLli0mkLl5z5Q7RIV1ObAfNaZtbh6mG+pl
x1WxYShGeDlM203+QHLMeVJoE2d/yudTrZD1To/HFzeXqaqaRzmY6po38cikSJ5TF6KRZwEKBOzC
x7Y/N1u6BCIpAN2dZEBUe5EGJ+BPmv/HPEtclNnvcim36rcJCj82Xp6sGnyOxjTHqpExHbu3w0uY
Wb6QjF+cejHVanKXfGZCTE4r+MI1AnCL/TTC64K8DceJNArLfc8j6nALsHo1TX0Gz6PZU8H93d1z
m/TD2EUhLNgwAZQm1f+4VI4P8f3rvF4/FAhTprnX/Gjx57HyW2ADqEj5ZeVQ0LWgXJD757BjIxBz
N+zQT4VekxgnlpVjmZCvTTam1x+g6FJAVg7rDeGhfkeUA6Nm521rR/a9KVnlCQcCNSdpk/iYjNe6
vdBVTgixi6e5ScC+MJ5TSxRWiCody5lmoSZgfU2F1b136pRFnppPwpa6iIEZ6NJsELmvS4vViJQk
qHHDKzkEMKv/dnBZRSntZpH3DyU3mB9HP3Blsbsp38TdITokPd55aCikqnC6RTLSQrGf5ZHMWhjI
/3d+z4AkOotKIJN3k93nEVb/o4iukzb00Oiyj134XnECAS8AIBk5lre7KgY29ua8I4REyGv8miQk
Ljkw0OLTLFKUSS2H11Tqvx1iit7PCIrU+fCPypY3dZhhakYHCSRdMR1VEGpYsyh0cow06X5vENaS
JlMD28D2bxoCnY0geEZWyvAz60NVPD2lIN/vYgmNA3qnjkwv2bRepc3GRYIn7UCvXQw1erHv/Cxv
YVJWUHRpP5ZPro/y/sqAvE4nJODYWk2LZM2G/Jq3qoqG+HAspUA9AfAvBKmPNacylbgzB4PAQ2yE
kDcIuOnhtemco4Qnkop2FEcVUuRxDSc1W56rbCXv6XZpU2finP8CX0iWmBSDgh7QeDjWNRLcnKCP
akAc1KV8o6iN80OLyNkVN3KNbEVpAidD7Xc0U1BBAppLwawbfL6xZC4ZFVZ0Lm4yIwP2PyswA+t/
lEJ8qcvsSfGG46euYjWpJZva0xtx+UtXE4/ZJRBhkzveZjlSoVVA1AkDiQLEsDwkZWJ6bDXB7175
mfxhphIy1iqGqNPh7sfh5v1Wrmryfh+228ydZywDvhGKMvtbI7FVbPaEBeqn7yasv+oX3EbjJqQW
EuHumTYzqHp1QaG88z3Fx9kQpju0in6vT8CkY/PAEwzWEOyTeFCWPrMsGegRbbQu8UnDMfDEPmwW
IfAHuN0r0LLb8jEJAIulxSNKNIeGzmpq0Knbjd/o89td7CaiI1UIyt9pG0IOJBAER1vaQJglVbP0
w736djwFBU5JA/jHz2ZGtaXueGqNcZTOAsVozEqFr1KTkQjBRFq9RB9pU2KU6L/ZXCbaJfzE4/3e
7LNQoMdXjtQLhtVZGlsWcxd4Vdp3U1CgVCwX5T2EVDdmqFOIHPABxqJlz2fJ4j3YeQjl+snjTB4Z
BDiT2v3PwRNZ+DrBnpwJDSoU5NNtEWwpC+tUC0UaHPJ+NfW2RBdj/9GmU2WwA0TMfZkN7BSwL7Jh
76CTM9Tygme4ey41+TBq0dn9Vvu6sFYemIhZwS+P1m/RUCUrjzhoID6iFwNqtt7zcLYyiKsUG2VT
kutaJpP6fwEBKZ1qNa5cFrNeI5ovdDKhsptzOPZtOBLoEnlq/U0rdRcMn+FdPYtdXagQEUc3c8cV
TSDfzuGHlFEhkw0WWnQuNXngatCXzLr1ebaa7skiWOv/6kUf5towP7UW52rFSgYo+YOPAQQwSIWu
h4tYbKjRyVCnk9oe8itd8oE0pY+7QBsj+IBDIb8quYVQhYACpwBdtDU6
`protect end_protected

