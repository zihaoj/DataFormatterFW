------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.3
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : gt625_fab20_init.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--  Description : This module instantiates the modules required for
--                reset and initialisation of the Transceiver
--
-- Module gt625_fab20_init
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;

--***********************************Entity Declaration************************

entity gt625_fab20_init is
generic
(
    EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "TRUE";     -- simulation setting for GT SecureIP model
    EXAMPLE_SIMULATION                      : integer   := 0;          -- Set to 1 for simulation
 
    STABLE_CLOCK_PERIOD                     : integer   := 20;  
        -- Set to 1 for simulation
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 0           -- Set to 1 to use Chipscope to drive resets

);
port
(
    SYSCLK_IN                               : in   std_logic;
    SOFT_RESET_IN                           : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT1_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT1_DATA_VALID_IN                       : in   std_logic;
    GT2_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT2_DATA_VALID_IN                       : in   std_logic;
    GT3_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT3_DATA_VALID_IN                       : in   std_logic;
    GT4_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT4_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT4_DATA_VALID_IN                       : in   std_logic;
    GT5_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT5_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT5_DATA_VALID_IN                       : in   std_logic;
    GT6_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT6_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT6_DATA_VALID_IN                       : in   std_logic;
    GT7_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT7_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT7_DATA_VALID_IN                       : in   std_logic;
    GT8_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT8_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT8_DATA_VALID_IN                       : in   std_logic;
    GT9_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT9_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT9_DATA_VALID_IN                       : in   std_logic;
    GT10_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT10_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT10_DATA_VALID_IN                      : in   std_logic;
    GT11_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT11_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT11_DATA_VALID_IN                      : in   std_logic;
    GT12_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT12_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT12_DATA_VALID_IN                      : in   std_logic;
    GT13_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT13_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT13_DATA_VALID_IN                      : in   std_logic;
    GT14_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT14_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT14_DATA_VALID_IN                      : in   std_logic;
    GT15_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT15_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT15_DATA_VALID_IN                      : in   std_logic;
    GT16_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT16_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT16_DATA_VALID_IN                      : in   std_logic;
    GT17_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT17_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT17_DATA_VALID_IN                      : in   std_logic;
    GT18_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT18_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT18_DATA_VALID_IN                      : in   std_logic;
    GT19_TX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT19_RX_FSM_RESET_DONE_OUT              : out  std_logic;
    GT19_DATA_VALID_IN                      : in   std_logic;

    --_________________________________________________________________________
    --GT0  (X1Y8)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt0_cpllfbclklost_out                   : out  std_logic;
    gt0_cplllock_out                        : out  std_logic;
    gt0_cplllockdetclk_in                   : in   std_logic;
    gt0_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt0_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxbyteisaligned_out                 : out  std_logic;
    gt0_rxmcommaalignen_in                  : in   std_logic;
    gt0_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt0_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt0_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt0_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT1  (X1Y9)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt1_cpllfbclklost_out                   : out  std_logic;
    gt1_cplllock_out                        : out  std_logic;
    gt1_cplllockdetclk_in                   : in   std_logic;
    gt1_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt1_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpclk_in                           : in   std_logic;
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxbyteisaligned_out                 : out  std_logic;
    gt1_rxmcommaalignen_in                  : in   std_logic;
    gt1_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt1_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt1_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt1_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT2  (X1Y10)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt2_cpllfbclklost_out                   : out  std_logic;
    gt2_cplllock_out                        : out  std_logic;
    gt2_cplllockdetclk_in                   : in   std_logic;
    gt2_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt2_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpclk_in                           : in   std_logic;
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxbyteisaligned_out                 : out  std_logic;
    gt2_rxmcommaalignen_in                  : in   std_logic;
    gt2_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt2_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt2_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt2_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT3  (X1Y11)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt3_cpllfbclklost_out                   : out  std_logic;
    gt3_cplllock_out                        : out  std_logic;
    gt3_cplllockdetclk_in                   : in   std_logic;
    gt3_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt3_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpclk_in                           : in   std_logic;
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxbyteisaligned_out                 : out  std_logic;
    gt3_rxmcommaalignen_in                  : in   std_logic;
    gt3_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt3_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt3_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt3_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT4  (X1Y12)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt4_cpllfbclklost_out                   : out  std_logic;
    gt4_cplllock_out                        : out  std_logic;
    gt4_cplllockdetclk_in                   : in   std_logic;
    gt4_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt4_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt4_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt4_drpclk_in                           : in   std_logic;
    gt4_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt4_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt4_drpen_in                            : in   std_logic;
    gt4_drprdy_out                          : out  std_logic;
    gt4_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt4_eyescanreset_in                     : in   std_logic;
    gt4_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt4_eyescandataerror_out                : out  std_logic;
    gt4_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt4_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt4_rxusrclk_in                         : in   std_logic;
    gt4_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt4_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt4_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt4_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt4_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt4_rxbyteisaligned_out                 : out  std_logic;
    gt4_rxmcommaalignen_in                  : in   std_logic;
    gt4_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt4_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt4_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt4_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt4_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt4_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt4_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt4_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt4_gttxreset_in                        : in   std_logic;
    gt4_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt4_txusrclk_in                         : in   std_logic;
    gt4_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt4_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt4_gthtxn_out                          : out  std_logic;
    gt4_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt4_txoutclk_out                        : out  std_logic;
    gt4_txoutclkfabric_out                  : out  std_logic;
    gt4_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt4_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt4_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt4_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT5  (X1Y13)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt5_cpllfbclklost_out                   : out  std_logic;
    gt5_cplllock_out                        : out  std_logic;
    gt5_cplllockdetclk_in                   : in   std_logic;
    gt5_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt5_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt5_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt5_drpclk_in                           : in   std_logic;
    gt5_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt5_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt5_drpen_in                            : in   std_logic;
    gt5_drprdy_out                          : out  std_logic;
    gt5_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt5_eyescanreset_in                     : in   std_logic;
    gt5_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt5_eyescandataerror_out                : out  std_logic;
    gt5_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt5_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt5_rxusrclk_in                         : in   std_logic;
    gt5_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt5_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt5_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt5_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt5_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt5_rxbyteisaligned_out                 : out  std_logic;
    gt5_rxmcommaalignen_in                  : in   std_logic;
    gt5_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt5_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt5_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt5_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt5_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt5_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt5_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt5_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt5_gttxreset_in                        : in   std_logic;
    gt5_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt5_txusrclk_in                         : in   std_logic;
    gt5_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt5_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt5_gthtxn_out                          : out  std_logic;
    gt5_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt5_txoutclk_out                        : out  std_logic;
    gt5_txoutclkfabric_out                  : out  std_logic;
    gt5_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt5_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt5_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt5_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT6  (X1Y14)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt6_cpllfbclklost_out                   : out  std_logic;
    gt6_cplllock_out                        : out  std_logic;
    gt6_cplllockdetclk_in                   : in   std_logic;
    gt6_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt6_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt6_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt6_drpclk_in                           : in   std_logic;
    gt6_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt6_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt6_drpen_in                            : in   std_logic;
    gt6_drprdy_out                          : out  std_logic;
    gt6_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt6_eyescanreset_in                     : in   std_logic;
    gt6_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt6_eyescandataerror_out                : out  std_logic;
    gt6_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt6_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt6_rxusrclk_in                         : in   std_logic;
    gt6_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt6_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt6_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt6_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt6_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt6_rxbyteisaligned_out                 : out  std_logic;
    gt6_rxmcommaalignen_in                  : in   std_logic;
    gt6_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt6_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt6_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt6_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt6_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt6_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt6_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt6_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt6_gttxreset_in                        : in   std_logic;
    gt6_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt6_txusrclk_in                         : in   std_logic;
    gt6_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt6_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt6_gthtxn_out                          : out  std_logic;
    gt6_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt6_txoutclk_out                        : out  std_logic;
    gt6_txoutclkfabric_out                  : out  std_logic;
    gt6_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt6_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt6_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt6_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT7  (X1Y15)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt7_cpllfbclklost_out                   : out  std_logic;
    gt7_cplllock_out                        : out  std_logic;
    gt7_cplllockdetclk_in                   : in   std_logic;
    gt7_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt7_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt7_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt7_drpclk_in                           : in   std_logic;
    gt7_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt7_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt7_drpen_in                            : in   std_logic;
    gt7_drprdy_out                          : out  std_logic;
    gt7_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt7_eyescanreset_in                     : in   std_logic;
    gt7_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt7_eyescandataerror_out                : out  std_logic;
    gt7_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt7_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt7_rxusrclk_in                         : in   std_logic;
    gt7_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt7_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt7_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt7_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt7_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt7_rxbyteisaligned_out                 : out  std_logic;
    gt7_rxmcommaalignen_in                  : in   std_logic;
    gt7_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt7_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt7_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt7_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt7_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt7_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt7_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt7_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt7_gttxreset_in                        : in   std_logic;
    gt7_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt7_txusrclk_in                         : in   std_logic;
    gt7_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt7_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt7_gthtxn_out                          : out  std_logic;
    gt7_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt7_txoutclk_out                        : out  std_logic;
    gt7_txoutclkfabric_out                  : out  std_logic;
    gt7_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt7_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt7_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt7_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT8  (X1Y16)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt8_cpllfbclklost_out                   : out  std_logic;
    gt8_cplllock_out                        : out  std_logic;
    gt8_cplllockdetclk_in                   : in   std_logic;
    gt8_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt8_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt8_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt8_drpclk_in                           : in   std_logic;
    gt8_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt8_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt8_drpen_in                            : in   std_logic;
    gt8_drprdy_out                          : out  std_logic;
    gt8_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt8_eyescanreset_in                     : in   std_logic;
    gt8_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt8_eyescandataerror_out                : out  std_logic;
    gt8_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt8_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt8_rxusrclk_in                         : in   std_logic;
    gt8_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt8_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt8_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt8_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt8_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt8_rxbyteisaligned_out                 : out  std_logic;
    gt8_rxmcommaalignen_in                  : in   std_logic;
    gt8_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt8_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt8_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt8_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt8_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt8_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt8_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt8_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt8_gttxreset_in                        : in   std_logic;
    gt8_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt8_txusrclk_in                         : in   std_logic;
    gt8_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt8_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt8_gthtxn_out                          : out  std_logic;
    gt8_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt8_txoutclk_out                        : out  std_logic;
    gt8_txoutclkfabric_out                  : out  std_logic;
    gt8_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt8_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt8_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt8_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT9  (X1Y17)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt9_cpllfbclklost_out                   : out  std_logic;
    gt9_cplllock_out                        : out  std_logic;
    gt9_cplllockdetclk_in                   : in   std_logic;
    gt9_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt9_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt9_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt9_drpclk_in                           : in   std_logic;
    gt9_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt9_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt9_drpen_in                            : in   std_logic;
    gt9_drprdy_out                          : out  std_logic;
    gt9_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt9_eyescanreset_in                     : in   std_logic;
    gt9_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt9_eyescandataerror_out                : out  std_logic;
    gt9_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt9_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt9_rxusrclk_in                         : in   std_logic;
    gt9_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt9_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt9_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt9_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt9_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt9_rxbyteisaligned_out                 : out  std_logic;
    gt9_rxmcommaalignen_in                  : in   std_logic;
    gt9_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt9_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt9_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt9_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt9_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt9_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt9_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt9_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt9_gttxreset_in                        : in   std_logic;
    gt9_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt9_txusrclk_in                         : in   std_logic;
    gt9_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt9_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt9_gthtxn_out                          : out  std_logic;
    gt9_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt9_txoutclk_out                        : out  std_logic;
    gt9_txoutclkfabric_out                  : out  std_logic;
    gt9_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt9_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt9_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt9_txcharisk_in                        : in   std_logic_vector(3 downto 0);

    --GT10  (X1Y18)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt10_cpllfbclklost_out                  : out  std_logic;
    gt10_cplllock_out                       : out  std_logic;
    gt10_cplllockdetclk_in                  : in   std_logic;
    gt10_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt10_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt10_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt10_drpclk_in                          : in   std_logic;
    gt10_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt10_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt10_drpen_in                           : in   std_logic;
    gt10_drprdy_out                         : out  std_logic;
    gt10_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt10_eyescanreset_in                    : in   std_logic;
    gt10_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt10_eyescandataerror_out               : out  std_logic;
    gt10_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt10_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt10_rxusrclk_in                        : in   std_logic;
    gt10_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt10_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt10_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt10_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt10_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt10_rxbyteisaligned_out                : out  std_logic;
    gt10_rxmcommaalignen_in                 : in   std_logic;
    gt10_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt10_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt10_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt10_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt10_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt10_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt10_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt10_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt10_gttxreset_in                       : in   std_logic;
    gt10_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt10_txusrclk_in                        : in   std_logic;
    gt10_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt10_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt10_gthtxn_out                         : out  std_logic;
    gt10_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt10_txoutclk_out                       : out  std_logic;
    gt10_txoutclkfabric_out                 : out  std_logic;
    gt10_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt10_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt10_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt10_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT11  (X1Y19)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt11_cpllfbclklost_out                  : out  std_logic;
    gt11_cplllock_out                       : out  std_logic;
    gt11_cplllockdetclk_in                  : in   std_logic;
    gt11_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt11_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt11_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt11_drpclk_in                          : in   std_logic;
    gt11_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt11_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt11_drpen_in                           : in   std_logic;
    gt11_drprdy_out                         : out  std_logic;
    gt11_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt11_eyescanreset_in                    : in   std_logic;
    gt11_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt11_eyescandataerror_out               : out  std_logic;
    gt11_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt11_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt11_rxusrclk_in                        : in   std_logic;
    gt11_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt11_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt11_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt11_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt11_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt11_rxbyteisaligned_out                : out  std_logic;
    gt11_rxmcommaalignen_in                 : in   std_logic;
    gt11_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt11_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt11_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt11_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt11_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt11_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt11_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt11_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt11_gttxreset_in                       : in   std_logic;
    gt11_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt11_txusrclk_in                        : in   std_logic;
    gt11_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt11_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt11_gthtxn_out                         : out  std_logic;
    gt11_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt11_txoutclk_out                       : out  std_logic;
    gt11_txoutclkfabric_out                 : out  std_logic;
    gt11_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt11_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt11_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt11_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT12  (X1Y20)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt12_cpllfbclklost_out                  : out  std_logic;
    gt12_cplllock_out                       : out  std_logic;
    gt12_cplllockdetclk_in                  : in   std_logic;
    gt12_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt12_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt12_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt12_drpclk_in                          : in   std_logic;
    gt12_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt12_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt12_drpen_in                           : in   std_logic;
    gt12_drprdy_out                         : out  std_logic;
    gt12_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt12_eyescanreset_in                    : in   std_logic;
    gt12_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt12_eyescandataerror_out               : out  std_logic;
    gt12_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt12_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt12_rxusrclk_in                        : in   std_logic;
    gt12_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt12_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt12_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt12_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt12_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt12_rxbyteisaligned_out                : out  std_logic;
    gt12_rxmcommaalignen_in                 : in   std_logic;
    gt12_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt12_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt12_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt12_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt12_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt12_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt12_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt12_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt12_gttxreset_in                       : in   std_logic;
    gt12_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt12_txusrclk_in                        : in   std_logic;
    gt12_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt12_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt12_gthtxn_out                         : out  std_logic;
    gt12_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt12_txoutclk_out                       : out  std_logic;
    gt12_txoutclkfabric_out                 : out  std_logic;
    gt12_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt12_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt12_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt12_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT13  (X1Y21)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt13_cpllfbclklost_out                  : out  std_logic;
    gt13_cplllock_out                       : out  std_logic;
    gt13_cplllockdetclk_in                  : in   std_logic;
    gt13_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt13_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt13_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt13_drpclk_in                          : in   std_logic;
    gt13_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt13_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt13_drpen_in                           : in   std_logic;
    gt13_drprdy_out                         : out  std_logic;
    gt13_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt13_eyescanreset_in                    : in   std_logic;
    gt13_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt13_eyescandataerror_out               : out  std_logic;
    gt13_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt13_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt13_rxusrclk_in                        : in   std_logic;
    gt13_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt13_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt13_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt13_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt13_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt13_rxbyteisaligned_out                : out  std_logic;
    gt13_rxmcommaalignen_in                 : in   std_logic;
    gt13_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt13_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt13_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt13_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt13_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt13_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt13_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt13_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt13_gttxreset_in                       : in   std_logic;
    gt13_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt13_txusrclk_in                        : in   std_logic;
    gt13_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt13_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt13_gthtxn_out                         : out  std_logic;
    gt13_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt13_txoutclk_out                       : out  std_logic;
    gt13_txoutclkfabric_out                 : out  std_logic;
    gt13_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt13_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt13_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt13_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT14  (X1Y22)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt14_cpllfbclklost_out                  : out  std_logic;
    gt14_cplllock_out                       : out  std_logic;
    gt14_cplllockdetclk_in                  : in   std_logic;
    gt14_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt14_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt14_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt14_drpclk_in                          : in   std_logic;
    gt14_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt14_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt14_drpen_in                           : in   std_logic;
    gt14_drprdy_out                         : out  std_logic;
    gt14_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt14_eyescanreset_in                    : in   std_logic;
    gt14_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt14_eyescandataerror_out               : out  std_logic;
    gt14_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt14_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt14_rxusrclk_in                        : in   std_logic;
    gt14_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt14_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt14_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt14_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt14_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt14_rxbyteisaligned_out                : out  std_logic;
    gt14_rxmcommaalignen_in                 : in   std_logic;
    gt14_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt14_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt14_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt14_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt14_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt14_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt14_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt14_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt14_gttxreset_in                       : in   std_logic;
    gt14_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt14_txusrclk_in                        : in   std_logic;
    gt14_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt14_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt14_gthtxn_out                         : out  std_logic;
    gt14_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt14_txoutclk_out                       : out  std_logic;
    gt14_txoutclkfabric_out                 : out  std_logic;
    gt14_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt14_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt14_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt14_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT15  (X1Y23)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt15_cpllfbclklost_out                  : out  std_logic;
    gt15_cplllock_out                       : out  std_logic;
    gt15_cplllockdetclk_in                  : in   std_logic;
    gt15_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt15_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt15_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt15_drpclk_in                          : in   std_logic;
    gt15_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt15_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt15_drpen_in                           : in   std_logic;
    gt15_drprdy_out                         : out  std_logic;
    gt15_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt15_eyescanreset_in                    : in   std_logic;
    gt15_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt15_eyescandataerror_out               : out  std_logic;
    gt15_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt15_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt15_rxusrclk_in                        : in   std_logic;
    gt15_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt15_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt15_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt15_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt15_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt15_rxbyteisaligned_out                : out  std_logic;
    gt15_rxmcommaalignen_in                 : in   std_logic;
    gt15_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt15_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt15_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt15_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt15_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt15_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt15_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt15_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt15_gttxreset_in                       : in   std_logic;
    gt15_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt15_txusrclk_in                        : in   std_logic;
    gt15_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt15_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt15_gthtxn_out                         : out  std_logic;
    gt15_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt15_txoutclk_out                       : out  std_logic;
    gt15_txoutclkfabric_out                 : out  std_logic;
    gt15_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt15_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt15_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt15_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT16  (X1Y24)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt16_cpllfbclklost_out                  : out  std_logic;
    gt16_cplllock_out                       : out  std_logic;
    gt16_cplllockdetclk_in                  : in   std_logic;
    gt16_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt16_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt16_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt16_drpclk_in                          : in   std_logic;
    gt16_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt16_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt16_drpen_in                           : in   std_logic;
    gt16_drprdy_out                         : out  std_logic;
    gt16_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt16_eyescanreset_in                    : in   std_logic;
    gt16_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt16_eyescandataerror_out               : out  std_logic;
    gt16_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt16_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt16_rxusrclk_in                        : in   std_logic;
    gt16_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt16_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt16_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt16_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt16_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt16_rxbyteisaligned_out                : out  std_logic;
    gt16_rxmcommaalignen_in                 : in   std_logic;
    gt16_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt16_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt16_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt16_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt16_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt16_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt16_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt16_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt16_gttxreset_in                       : in   std_logic;
    gt16_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt16_txusrclk_in                        : in   std_logic;
    gt16_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt16_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt16_gthtxn_out                         : out  std_logic;
    gt16_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt16_txoutclk_out                       : out  std_logic;
    gt16_txoutclkfabric_out                 : out  std_logic;
    gt16_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt16_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt16_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt16_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT17  (X1Y25)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt17_cpllfbclklost_out                  : out  std_logic;
    gt17_cplllock_out                       : out  std_logic;
    gt17_cplllockdetclk_in                  : in   std_logic;
    gt17_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt17_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt17_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt17_drpclk_in                          : in   std_logic;
    gt17_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt17_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt17_drpen_in                           : in   std_logic;
    gt17_drprdy_out                         : out  std_logic;
    gt17_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt17_eyescanreset_in                    : in   std_logic;
    gt17_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt17_eyescandataerror_out               : out  std_logic;
    gt17_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt17_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt17_rxusrclk_in                        : in   std_logic;
    gt17_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt17_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt17_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt17_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt17_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt17_rxbyteisaligned_out                : out  std_logic;
    gt17_rxmcommaalignen_in                 : in   std_logic;
    gt17_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt17_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt17_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt17_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt17_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt17_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt17_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt17_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt17_gttxreset_in                       : in   std_logic;
    gt17_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt17_txusrclk_in                        : in   std_logic;
    gt17_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt17_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt17_gthtxn_out                         : out  std_logic;
    gt17_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt17_txoutclk_out                       : out  std_logic;
    gt17_txoutclkfabric_out                 : out  std_logic;
    gt17_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt17_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt17_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt17_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT18  (X1Y26)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt18_cpllfbclklost_out                  : out  std_logic;
    gt18_cplllock_out                       : out  std_logic;
    gt18_cplllockdetclk_in                  : in   std_logic;
    gt18_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt18_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt18_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt18_drpclk_in                          : in   std_logic;
    gt18_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt18_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt18_drpen_in                           : in   std_logic;
    gt18_drprdy_out                         : out  std_logic;
    gt18_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt18_eyescanreset_in                    : in   std_logic;
    gt18_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt18_eyescandataerror_out               : out  std_logic;
    gt18_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt18_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt18_rxusrclk_in                        : in   std_logic;
    gt18_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt18_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt18_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt18_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt18_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt18_rxbyteisaligned_out                : out  std_logic;
    gt18_rxmcommaalignen_in                 : in   std_logic;
    gt18_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt18_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt18_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt18_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt18_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt18_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt18_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt18_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt18_gttxreset_in                       : in   std_logic;
    gt18_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt18_txusrclk_in                        : in   std_logic;
    gt18_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt18_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt18_gthtxn_out                         : out  std_logic;
    gt18_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt18_txoutclk_out                       : out  std_logic;
    gt18_txoutclkfabric_out                 : out  std_logic;
    gt18_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt18_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt18_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt18_txcharisk_in                       : in   std_logic_vector(3 downto 0);

    --GT19  (X1Y27)
    --____________________________CHANNEL PORTS________________________________
    --------------------------------- CPLL Ports -------------------------------
    gt19_cpllfbclklost_out                  : out  std_logic;
    gt19_cplllock_out                       : out  std_logic;
    gt19_cplllockdetclk_in                  : in   std_logic;
    gt19_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt19_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt19_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt19_drpclk_in                          : in   std_logic;
    gt19_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt19_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt19_drpen_in                           : in   std_logic;
    gt19_drprdy_out                         : out  std_logic;
    gt19_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt19_eyescanreset_in                    : in   std_logic;
    gt19_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt19_eyescandataerror_out               : out  std_logic;
    gt19_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt19_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt19_rxusrclk_in                        : in   std_logic;
    gt19_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt19_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt19_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt19_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt19_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt19_rxbyteisaligned_out                : out  std_logic;
    gt19_rxmcommaalignen_in                 : in   std_logic;
    gt19_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt19_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt19_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt19_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt19_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt19_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt19_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt19_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt19_gttxreset_in                       : in   std_logic;
    gt19_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt19_txusrclk_in                        : in   std_logic;
    gt19_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt19_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt19_gthtxn_out                         : out  std_logic;
    gt19_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt19_txoutclk_out                       : out  std_logic;
    gt19_txoutclkfabric_out                 : out  std_logic;
    gt19_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt19_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt19_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt19_txcharisk_in                       : in   std_logic_vector(3 downto 0);


    --____________________________COMMON PORTS________________________________
     GT0_QPLLOUTCLK_IN  : in std_logic;
     GT0_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT1_QPLLOUTCLK_IN  : in std_logic;
     GT1_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT2_QPLLOUTCLK_IN  : in std_logic;
     GT2_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT3_QPLLOUTCLK_IN  : in std_logic;
     GT3_QPLLOUTREFCLK_IN : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT4_QPLLOUTCLK_IN  : in std_logic;
     GT4_QPLLOUTREFCLK_IN : in std_logic

);

end gt625_fab20_init;
    
architecture RTL of gt625_fab20_init is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

--**************************Component Declarations*****************************


component gt625_fab20_multi_gt 
generic
(
    -- Simulation attributes
    EXAMPLE_SIMULATION             : integer   := 0;      -- Set to 1 for simulation
    WRAPPER_SIM_GTRESET_SPEEDUP    : string    := "FALSE" -- Set to "TRUE" to speed up sim reset

);
port
(

    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT0  (X1Y8)
    --____________________________CHANNEL PORTS________________________________
    GT0_RXPMARESETDONE_OUT                        : out  std_logic;
    GT0_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt0_cpllfbclklost_out                   : out  std_logic;
    gt0_cplllock_out                        : out  std_logic;
    gt0_cplllockdetclk_in                   : in   std_logic;
    gt0_cpllrefclklost_out                  : out  std_logic;
    gt0_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt0_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxbyteisaligned_out                 : out  std_logic;
    gt0_rxmcommaalignen_in                  : in   std_logic;
    gt0_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt0_rxdfeagchold_in                     : in   std_logic;
    gt0_rxdfelfhold_in                      : in   std_logic;
    gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt0_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt0_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt0_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt0_gthtxn_out                          : out  std_logic;
    gt0_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt0_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt0_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT1  (X1Y9)
    --____________________________CHANNEL PORTS________________________________
    GT1_RXPMARESETDONE_OUT                        : out  std_logic;
    GT1_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt1_cpllfbclklost_out                   : out  std_logic;
    gt1_cplllock_out                        : out  std_logic;
    gt1_cplllockdetclk_in                   : in   std_logic;
    gt1_cpllrefclklost_out                  : out  std_logic;
    gt1_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt1_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt1_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt1_drpclk_in                           : in   std_logic;
    gt1_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt1_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt1_drpen_in                            : in   std_logic;
    gt1_drprdy_out                          : out  std_logic;
    gt1_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt1_eyescanreset_in                     : in   std_logic;
    gt1_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt1_eyescandataerror_out                : out  std_logic;
    gt1_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt1_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt1_rxusrclk_in                         : in   std_logic;
    gt1_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt1_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt1_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt1_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt1_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt1_rxbyteisaligned_out                 : out  std_logic;
    gt1_rxmcommaalignen_in                  : in   std_logic;
    gt1_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt1_rxdfeagchold_in                     : in   std_logic;
    gt1_rxdfelfhold_in                      : in   std_logic;
    gt1_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt1_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt1_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt1_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt1_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt1_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt1_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt1_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt1_gttxreset_in                        : in   std_logic;
    gt1_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt1_txusrclk_in                         : in   std_logic;
    gt1_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt1_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt1_gthtxn_out                          : out  std_logic;
    gt1_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt1_txoutclk_out                        : out  std_logic;
    gt1_txoutclkfabric_out                  : out  std_logic;
    gt1_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt1_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt1_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt1_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT2  (X1Y10)
    --____________________________CHANNEL PORTS________________________________
    GT2_RXPMARESETDONE_OUT                        : out  std_logic;
    GT2_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt2_cpllfbclklost_out                   : out  std_logic;
    gt2_cplllock_out                        : out  std_logic;
    gt2_cplllockdetclk_in                   : in   std_logic;
    gt2_cpllrefclklost_out                  : out  std_logic;
    gt2_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt2_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt2_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt2_drpclk_in                           : in   std_logic;
    gt2_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt2_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt2_drpen_in                            : in   std_logic;
    gt2_drprdy_out                          : out  std_logic;
    gt2_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt2_eyescanreset_in                     : in   std_logic;
    gt2_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt2_eyescandataerror_out                : out  std_logic;
    gt2_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt2_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt2_rxusrclk_in                         : in   std_logic;
    gt2_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt2_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt2_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt2_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt2_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt2_rxbyteisaligned_out                 : out  std_logic;
    gt2_rxmcommaalignen_in                  : in   std_logic;
    gt2_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt2_rxdfeagchold_in                     : in   std_logic;
    gt2_rxdfelfhold_in                      : in   std_logic;
    gt2_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt2_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt2_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt2_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt2_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt2_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt2_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt2_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt2_gttxreset_in                        : in   std_logic;
    gt2_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt2_txusrclk_in                         : in   std_logic;
    gt2_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt2_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt2_gthtxn_out                          : out  std_logic;
    gt2_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt2_txoutclk_out                        : out  std_logic;
    gt2_txoutclkfabric_out                  : out  std_logic;
    gt2_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt2_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt2_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt2_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT3  (X1Y11)
    --____________________________CHANNEL PORTS________________________________
    GT3_RXPMARESETDONE_OUT                        : out  std_logic;
    GT3_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt3_cpllfbclklost_out                   : out  std_logic;
    gt3_cplllock_out                        : out  std_logic;
    gt3_cplllockdetclk_in                   : in   std_logic;
    gt3_cpllrefclklost_out                  : out  std_logic;
    gt3_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt3_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt3_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt3_drpclk_in                           : in   std_logic;
    gt3_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt3_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt3_drpen_in                            : in   std_logic;
    gt3_drprdy_out                          : out  std_logic;
    gt3_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt3_eyescanreset_in                     : in   std_logic;
    gt3_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt3_eyescandataerror_out                : out  std_logic;
    gt3_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt3_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt3_rxusrclk_in                         : in   std_logic;
    gt3_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt3_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt3_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt3_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt3_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt3_rxbyteisaligned_out                 : out  std_logic;
    gt3_rxmcommaalignen_in                  : in   std_logic;
    gt3_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt3_rxdfeagchold_in                     : in   std_logic;
    gt3_rxdfelfhold_in                      : in   std_logic;
    gt3_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt3_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt3_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt3_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt3_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt3_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt3_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt3_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt3_gttxreset_in                        : in   std_logic;
    gt3_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt3_txusrclk_in                         : in   std_logic;
    gt3_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt3_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt3_gthtxn_out                          : out  std_logic;
    gt3_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt3_txoutclk_out                        : out  std_logic;
    gt3_txoutclkfabric_out                  : out  std_logic;
    gt3_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt3_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt3_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt3_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT4  (X1Y12)
    --____________________________CHANNEL PORTS________________________________
    GT4_RXPMARESETDONE_OUT                        : out  std_logic;
    GT4_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt4_cpllfbclklost_out                   : out  std_logic;
    gt4_cplllock_out                        : out  std_logic;
    gt4_cplllockdetclk_in                   : in   std_logic;
    gt4_cpllrefclklost_out                  : out  std_logic;
    gt4_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt4_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt4_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt4_drpclk_in                           : in   std_logic;
    gt4_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt4_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt4_drpen_in                            : in   std_logic;
    gt4_drprdy_out                          : out  std_logic;
    gt4_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt4_eyescanreset_in                     : in   std_logic;
    gt4_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt4_eyescandataerror_out                : out  std_logic;
    gt4_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt4_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt4_rxusrclk_in                         : in   std_logic;
    gt4_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt4_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt4_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt4_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt4_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt4_rxbyteisaligned_out                 : out  std_logic;
    gt4_rxmcommaalignen_in                  : in   std_logic;
    gt4_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt4_rxdfeagchold_in                     : in   std_logic;
    gt4_rxdfelfhold_in                      : in   std_logic;
    gt4_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt4_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt4_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt4_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt4_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt4_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt4_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt4_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt4_gttxreset_in                        : in   std_logic;
    gt4_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt4_txusrclk_in                         : in   std_logic;
    gt4_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt4_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt4_gthtxn_out                          : out  std_logic;
    gt4_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt4_txoutclk_out                        : out  std_logic;
    gt4_txoutclkfabric_out                  : out  std_logic;
    gt4_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt4_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt4_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt4_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT5  (X1Y13)
    --____________________________CHANNEL PORTS________________________________
    GT5_RXPMARESETDONE_OUT                        : out  std_logic;
    GT5_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt5_cpllfbclklost_out                   : out  std_logic;
    gt5_cplllock_out                        : out  std_logic;
    gt5_cplllockdetclk_in                   : in   std_logic;
    gt5_cpllrefclklost_out                  : out  std_logic;
    gt5_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt5_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt5_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt5_drpclk_in                           : in   std_logic;
    gt5_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt5_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt5_drpen_in                            : in   std_logic;
    gt5_drprdy_out                          : out  std_logic;
    gt5_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt5_eyescanreset_in                     : in   std_logic;
    gt5_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt5_eyescandataerror_out                : out  std_logic;
    gt5_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt5_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt5_rxusrclk_in                         : in   std_logic;
    gt5_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt5_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt5_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt5_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt5_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt5_rxbyteisaligned_out                 : out  std_logic;
    gt5_rxmcommaalignen_in                  : in   std_logic;
    gt5_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt5_rxdfeagchold_in                     : in   std_logic;
    gt5_rxdfelfhold_in                      : in   std_logic;
    gt5_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt5_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt5_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt5_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt5_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt5_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt5_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt5_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt5_gttxreset_in                        : in   std_logic;
    gt5_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt5_txusrclk_in                         : in   std_logic;
    gt5_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt5_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt5_gthtxn_out                          : out  std_logic;
    gt5_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt5_txoutclk_out                        : out  std_logic;
    gt5_txoutclkfabric_out                  : out  std_logic;
    gt5_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt5_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt5_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt5_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT6  (X1Y14)
    --____________________________CHANNEL PORTS________________________________
    GT6_RXPMARESETDONE_OUT                        : out  std_logic;
    GT6_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt6_cpllfbclklost_out                   : out  std_logic;
    gt6_cplllock_out                        : out  std_logic;
    gt6_cplllockdetclk_in                   : in   std_logic;
    gt6_cpllrefclklost_out                  : out  std_logic;
    gt6_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt6_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt6_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt6_drpclk_in                           : in   std_logic;
    gt6_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt6_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt6_drpen_in                            : in   std_logic;
    gt6_drprdy_out                          : out  std_logic;
    gt6_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt6_eyescanreset_in                     : in   std_logic;
    gt6_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt6_eyescandataerror_out                : out  std_logic;
    gt6_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt6_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt6_rxusrclk_in                         : in   std_logic;
    gt6_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt6_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt6_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt6_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt6_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt6_rxbyteisaligned_out                 : out  std_logic;
    gt6_rxmcommaalignen_in                  : in   std_logic;
    gt6_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt6_rxdfeagchold_in                     : in   std_logic;
    gt6_rxdfelfhold_in                      : in   std_logic;
    gt6_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt6_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt6_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt6_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt6_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt6_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt6_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt6_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt6_gttxreset_in                        : in   std_logic;
    gt6_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt6_txusrclk_in                         : in   std_logic;
    gt6_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt6_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt6_gthtxn_out                          : out  std_logic;
    gt6_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt6_txoutclk_out                        : out  std_logic;
    gt6_txoutclkfabric_out                  : out  std_logic;
    gt6_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt6_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt6_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt6_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT7  (X1Y15)
    --____________________________CHANNEL PORTS________________________________
    GT7_RXPMARESETDONE_OUT                        : out  std_logic;
    GT7_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt7_cpllfbclklost_out                   : out  std_logic;
    gt7_cplllock_out                        : out  std_logic;
    gt7_cplllockdetclk_in                   : in   std_logic;
    gt7_cpllrefclklost_out                  : out  std_logic;
    gt7_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt7_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt7_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt7_drpclk_in                           : in   std_logic;
    gt7_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt7_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt7_drpen_in                            : in   std_logic;
    gt7_drprdy_out                          : out  std_logic;
    gt7_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt7_eyescanreset_in                     : in   std_logic;
    gt7_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt7_eyescandataerror_out                : out  std_logic;
    gt7_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt7_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt7_rxusrclk_in                         : in   std_logic;
    gt7_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt7_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt7_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt7_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt7_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt7_rxbyteisaligned_out                 : out  std_logic;
    gt7_rxmcommaalignen_in                  : in   std_logic;
    gt7_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt7_rxdfeagchold_in                     : in   std_logic;
    gt7_rxdfelfhold_in                      : in   std_logic;
    gt7_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt7_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt7_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt7_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt7_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt7_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt7_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt7_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt7_gttxreset_in                        : in   std_logic;
    gt7_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt7_txusrclk_in                         : in   std_logic;
    gt7_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt7_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt7_gthtxn_out                          : out  std_logic;
    gt7_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt7_txoutclk_out                        : out  std_logic;
    gt7_txoutclkfabric_out                  : out  std_logic;
    gt7_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt7_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt7_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt7_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT8  (X1Y16)
    --____________________________CHANNEL PORTS________________________________
    GT8_RXPMARESETDONE_OUT                        : out  std_logic;
    GT8_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt8_cpllfbclklost_out                   : out  std_logic;
    gt8_cplllock_out                        : out  std_logic;
    gt8_cplllockdetclk_in                   : in   std_logic;
    gt8_cpllrefclklost_out                  : out  std_logic;
    gt8_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt8_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt8_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt8_drpclk_in                           : in   std_logic;
    gt8_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt8_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt8_drpen_in                            : in   std_logic;
    gt8_drprdy_out                          : out  std_logic;
    gt8_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt8_eyescanreset_in                     : in   std_logic;
    gt8_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt8_eyescandataerror_out                : out  std_logic;
    gt8_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt8_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt8_rxusrclk_in                         : in   std_logic;
    gt8_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt8_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt8_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt8_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt8_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt8_rxbyteisaligned_out                 : out  std_logic;
    gt8_rxmcommaalignen_in                  : in   std_logic;
    gt8_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt8_rxdfeagchold_in                     : in   std_logic;
    gt8_rxdfelfhold_in                      : in   std_logic;
    gt8_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt8_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt8_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt8_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt8_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt8_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt8_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt8_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt8_gttxreset_in                        : in   std_logic;
    gt8_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt8_txusrclk_in                         : in   std_logic;
    gt8_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt8_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt8_gthtxn_out                          : out  std_logic;
    gt8_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt8_txoutclk_out                        : out  std_logic;
    gt8_txoutclkfabric_out                  : out  std_logic;
    gt8_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt8_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt8_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt8_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT9  (X1Y17)
    --____________________________CHANNEL PORTS________________________________
    GT9_RXPMARESETDONE_OUT                        : out  std_logic;
    GT9_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt9_cpllfbclklost_out                   : out  std_logic;
    gt9_cplllock_out                        : out  std_logic;
    gt9_cplllockdetclk_in                   : in   std_logic;
    gt9_cpllrefclklost_out                  : out  std_logic;
    gt9_cpllreset_in                        : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt9_gtrefclk0_in                        : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt9_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt9_drpclk_in                           : in   std_logic;
    gt9_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt9_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt9_drpen_in                            : in   std_logic;
    gt9_drprdy_out                          : out  std_logic;
    gt9_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt9_eyescanreset_in                     : in   std_logic;
    gt9_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt9_eyescandataerror_out                : out  std_logic;
    gt9_eyescantrigger_in                   : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt9_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt9_rxusrclk_in                         : in   std_logic;
    gt9_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt9_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt9_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt9_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt9_gthrxn_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt9_rxbyteisaligned_out                 : out  std_logic;
    gt9_rxmcommaalignen_in                  : in   std_logic;
    gt9_rxpcommaalignen_in                  : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt9_rxdfeagchold_in                     : in   std_logic;
    gt9_rxdfelfhold_in                      : in   std_logic;
    gt9_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
    gt9_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt9_rxoutclk_out                        : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt9_gtrxreset_in                        : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt9_rxpolarity_in                       : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt9_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt9_gthrxp_in                           : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt9_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt9_gttxreset_in                        : in   std_logic;
    gt9_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt9_txusrclk_in                         : in   std_logic;
    gt9_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt9_txdata_in                           : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt9_gthtxn_out                          : out  std_logic;
    gt9_gthtxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt9_txoutclk_out                        : out  std_logic;
    gt9_txoutclkfabric_out                  : out  std_logic;
    gt9_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt9_txresetdone_out                     : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt9_txpolarity_in                       : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt9_txcharisk_in                        : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT10  (X1Y18)
    --____________________________CHANNEL PORTS________________________________
    GT10_RXPMARESETDONE_OUT                        : out  std_logic;
    GT10_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt10_cpllfbclklost_out                  : out  std_logic;
    gt10_cplllock_out                       : out  std_logic;
    gt10_cplllockdetclk_in                  : in   std_logic;
    gt10_cpllrefclklost_out                 : out  std_logic;
    gt10_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt10_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt10_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt10_drpclk_in                          : in   std_logic;
    gt10_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt10_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt10_drpen_in                           : in   std_logic;
    gt10_drprdy_out                         : out  std_logic;
    gt10_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt10_eyescanreset_in                    : in   std_logic;
    gt10_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt10_eyescandataerror_out               : out  std_logic;
    gt10_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt10_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt10_rxusrclk_in                        : in   std_logic;
    gt10_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt10_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt10_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt10_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt10_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt10_rxbyteisaligned_out                : out  std_logic;
    gt10_rxmcommaalignen_in                 : in   std_logic;
    gt10_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt10_rxdfeagchold_in                    : in   std_logic;
    gt10_rxdfelfhold_in                     : in   std_logic;
    gt10_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt10_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt10_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt10_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt10_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt10_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt10_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt10_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt10_gttxreset_in                       : in   std_logic;
    gt10_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt10_txusrclk_in                        : in   std_logic;
    gt10_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt10_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt10_gthtxn_out                         : out  std_logic;
    gt10_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt10_txoutclk_out                       : out  std_logic;
    gt10_txoutclkfabric_out                 : out  std_logic;
    gt10_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt10_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt10_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt10_txcharisk_in                       : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT11  (X1Y19)
    --____________________________CHANNEL PORTS________________________________
    GT11_RXPMARESETDONE_OUT                        : out  std_logic;
    GT11_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt11_cpllfbclklost_out                  : out  std_logic;
    gt11_cplllock_out                       : out  std_logic;
    gt11_cplllockdetclk_in                  : in   std_logic;
    gt11_cpllrefclklost_out                 : out  std_logic;
    gt11_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt11_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt11_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt11_drpclk_in                          : in   std_logic;
    gt11_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt11_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt11_drpen_in                           : in   std_logic;
    gt11_drprdy_out                         : out  std_logic;
    gt11_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt11_eyescanreset_in                    : in   std_logic;
    gt11_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt11_eyescandataerror_out               : out  std_logic;
    gt11_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt11_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt11_rxusrclk_in                        : in   std_logic;
    gt11_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt11_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt11_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt11_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt11_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt11_rxbyteisaligned_out                : out  std_logic;
    gt11_rxmcommaalignen_in                 : in   std_logic;
    gt11_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt11_rxdfeagchold_in                    : in   std_logic;
    gt11_rxdfelfhold_in                     : in   std_logic;
    gt11_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt11_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt11_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt11_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt11_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt11_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt11_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt11_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt11_gttxreset_in                       : in   std_logic;
    gt11_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt11_txusrclk_in                        : in   std_logic;
    gt11_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt11_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt11_gthtxn_out                         : out  std_logic;
    gt11_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt11_txoutclk_out                       : out  std_logic;
    gt11_txoutclkfabric_out                 : out  std_logic;
    gt11_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt11_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt11_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt11_txcharisk_in                       : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT12  (X1Y20)
    --____________________________CHANNEL PORTS________________________________
    GT12_RXPMARESETDONE_OUT                        : out  std_logic;
    GT12_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt12_cpllfbclklost_out                  : out  std_logic;
    gt12_cplllock_out                       : out  std_logic;
    gt12_cplllockdetclk_in                  : in   std_logic;
    gt12_cpllrefclklost_out                 : out  std_logic;
    gt12_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt12_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt12_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt12_drpclk_in                          : in   std_logic;
    gt12_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt12_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt12_drpen_in                           : in   std_logic;
    gt12_drprdy_out                         : out  std_logic;
    gt12_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt12_eyescanreset_in                    : in   std_logic;
    gt12_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt12_eyescandataerror_out               : out  std_logic;
    gt12_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt12_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt12_rxusrclk_in                        : in   std_logic;
    gt12_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt12_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt12_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt12_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt12_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt12_rxbyteisaligned_out                : out  std_logic;
    gt12_rxmcommaalignen_in                 : in   std_logic;
    gt12_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt12_rxdfeagchold_in                    : in   std_logic;
    gt12_rxdfelfhold_in                     : in   std_logic;
    gt12_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt12_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt12_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt12_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt12_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt12_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt12_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt12_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt12_gttxreset_in                       : in   std_logic;
    gt12_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt12_txusrclk_in                        : in   std_logic;
    gt12_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt12_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt12_gthtxn_out                         : out  std_logic;
    gt12_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt12_txoutclk_out                       : out  std_logic;
    gt12_txoutclkfabric_out                 : out  std_logic;
    gt12_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt12_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt12_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt12_txcharisk_in                       : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT13  (X1Y21)
    --____________________________CHANNEL PORTS________________________________
    GT13_RXPMARESETDONE_OUT                        : out  std_logic;
    GT13_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt13_cpllfbclklost_out                  : out  std_logic;
    gt13_cplllock_out                       : out  std_logic;
    gt13_cplllockdetclk_in                  : in   std_logic;
    gt13_cpllrefclklost_out                 : out  std_logic;
    gt13_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt13_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt13_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt13_drpclk_in                          : in   std_logic;
    gt13_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt13_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt13_drpen_in                           : in   std_logic;
    gt13_drprdy_out                         : out  std_logic;
    gt13_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt13_eyescanreset_in                    : in   std_logic;
    gt13_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt13_eyescandataerror_out               : out  std_logic;
    gt13_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt13_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt13_rxusrclk_in                        : in   std_logic;
    gt13_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt13_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt13_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt13_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt13_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt13_rxbyteisaligned_out                : out  std_logic;
    gt13_rxmcommaalignen_in                 : in   std_logic;
    gt13_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt13_rxdfeagchold_in                    : in   std_logic;
    gt13_rxdfelfhold_in                     : in   std_logic;
    gt13_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt13_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt13_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt13_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt13_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt13_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt13_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt13_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt13_gttxreset_in                       : in   std_logic;
    gt13_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt13_txusrclk_in                        : in   std_logic;
    gt13_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt13_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt13_gthtxn_out                         : out  std_logic;
    gt13_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt13_txoutclk_out                       : out  std_logic;
    gt13_txoutclkfabric_out                 : out  std_logic;
    gt13_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt13_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt13_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt13_txcharisk_in                       : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT14  (X1Y22)
    --____________________________CHANNEL PORTS________________________________
    GT14_RXPMARESETDONE_OUT                        : out  std_logic;
    GT14_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt14_cpllfbclklost_out                  : out  std_logic;
    gt14_cplllock_out                       : out  std_logic;
    gt14_cplllockdetclk_in                  : in   std_logic;
    gt14_cpllrefclklost_out                 : out  std_logic;
    gt14_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt14_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt14_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt14_drpclk_in                          : in   std_logic;
    gt14_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt14_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt14_drpen_in                           : in   std_logic;
    gt14_drprdy_out                         : out  std_logic;
    gt14_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt14_eyescanreset_in                    : in   std_logic;
    gt14_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt14_eyescandataerror_out               : out  std_logic;
    gt14_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt14_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt14_rxusrclk_in                        : in   std_logic;
    gt14_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt14_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt14_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt14_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt14_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt14_rxbyteisaligned_out                : out  std_logic;
    gt14_rxmcommaalignen_in                 : in   std_logic;
    gt14_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt14_rxdfeagchold_in                    : in   std_logic;
    gt14_rxdfelfhold_in                     : in   std_logic;
    gt14_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt14_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt14_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt14_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt14_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt14_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt14_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt14_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt14_gttxreset_in                       : in   std_logic;
    gt14_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt14_txusrclk_in                        : in   std_logic;
    gt14_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt14_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt14_gthtxn_out                         : out  std_logic;
    gt14_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt14_txoutclk_out                       : out  std_logic;
    gt14_txoutclkfabric_out                 : out  std_logic;
    gt14_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt14_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt14_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt14_txcharisk_in                       : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT15  (X1Y23)
    --____________________________CHANNEL PORTS________________________________
    GT15_RXPMARESETDONE_OUT                        : out  std_logic;
    GT15_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt15_cpllfbclklost_out                  : out  std_logic;
    gt15_cplllock_out                       : out  std_logic;
    gt15_cplllockdetclk_in                  : in   std_logic;
    gt15_cpllrefclklost_out                 : out  std_logic;
    gt15_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt15_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt15_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt15_drpclk_in                          : in   std_logic;
    gt15_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt15_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt15_drpen_in                           : in   std_logic;
    gt15_drprdy_out                         : out  std_logic;
    gt15_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt15_eyescanreset_in                    : in   std_logic;
    gt15_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt15_eyescandataerror_out               : out  std_logic;
    gt15_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt15_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt15_rxusrclk_in                        : in   std_logic;
    gt15_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt15_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt15_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt15_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt15_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt15_rxbyteisaligned_out                : out  std_logic;
    gt15_rxmcommaalignen_in                 : in   std_logic;
    gt15_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt15_rxdfeagchold_in                    : in   std_logic;
    gt15_rxdfelfhold_in                     : in   std_logic;
    gt15_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt15_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt15_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt15_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt15_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt15_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt15_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt15_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt15_gttxreset_in                       : in   std_logic;
    gt15_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt15_txusrclk_in                        : in   std_logic;
    gt15_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt15_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt15_gthtxn_out                         : out  std_logic;
    gt15_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt15_txoutclk_out                       : out  std_logic;
    gt15_txoutclkfabric_out                 : out  std_logic;
    gt15_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt15_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt15_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt15_txcharisk_in                       : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT16  (X1Y24)
    --____________________________CHANNEL PORTS________________________________
    GT16_RXPMARESETDONE_OUT                        : out  std_logic;
    GT16_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt16_cpllfbclklost_out                  : out  std_logic;
    gt16_cplllock_out                       : out  std_logic;
    gt16_cplllockdetclk_in                  : in   std_logic;
    gt16_cpllrefclklost_out                 : out  std_logic;
    gt16_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt16_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt16_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt16_drpclk_in                          : in   std_logic;
    gt16_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt16_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt16_drpen_in                           : in   std_logic;
    gt16_drprdy_out                         : out  std_logic;
    gt16_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt16_eyescanreset_in                    : in   std_logic;
    gt16_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt16_eyescandataerror_out               : out  std_logic;
    gt16_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt16_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt16_rxusrclk_in                        : in   std_logic;
    gt16_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt16_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt16_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt16_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt16_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt16_rxbyteisaligned_out                : out  std_logic;
    gt16_rxmcommaalignen_in                 : in   std_logic;
    gt16_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt16_rxdfeagchold_in                    : in   std_logic;
    gt16_rxdfelfhold_in                     : in   std_logic;
    gt16_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt16_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt16_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt16_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt16_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt16_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt16_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt16_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt16_gttxreset_in                       : in   std_logic;
    gt16_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt16_txusrclk_in                        : in   std_logic;
    gt16_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt16_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt16_gthtxn_out                         : out  std_logic;
    gt16_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt16_txoutclk_out                       : out  std_logic;
    gt16_txoutclkfabric_out                 : out  std_logic;
    gt16_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt16_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt16_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt16_txcharisk_in                       : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT17  (X1Y25)
    --____________________________CHANNEL PORTS________________________________
    GT17_RXPMARESETDONE_OUT                        : out  std_logic;
    GT17_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt17_cpllfbclklost_out                  : out  std_logic;
    gt17_cplllock_out                       : out  std_logic;
    gt17_cplllockdetclk_in                  : in   std_logic;
    gt17_cpllrefclklost_out                 : out  std_logic;
    gt17_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt17_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt17_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt17_drpclk_in                          : in   std_logic;
    gt17_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt17_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt17_drpen_in                           : in   std_logic;
    gt17_drprdy_out                         : out  std_logic;
    gt17_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt17_eyescanreset_in                    : in   std_logic;
    gt17_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt17_eyescandataerror_out               : out  std_logic;
    gt17_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt17_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt17_rxusrclk_in                        : in   std_logic;
    gt17_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt17_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt17_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt17_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt17_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt17_rxbyteisaligned_out                : out  std_logic;
    gt17_rxmcommaalignen_in                 : in   std_logic;
    gt17_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt17_rxdfeagchold_in                    : in   std_logic;
    gt17_rxdfelfhold_in                     : in   std_logic;
    gt17_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt17_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt17_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt17_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt17_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt17_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt17_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt17_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt17_gttxreset_in                       : in   std_logic;
    gt17_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt17_txusrclk_in                        : in   std_logic;
    gt17_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt17_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt17_gthtxn_out                         : out  std_logic;
    gt17_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt17_txoutclk_out                       : out  std_logic;
    gt17_txoutclkfabric_out                 : out  std_logic;
    gt17_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt17_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt17_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt17_txcharisk_in                       : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT18  (X1Y26)
    --____________________________CHANNEL PORTS________________________________
    GT18_RXPMARESETDONE_OUT                        : out  std_logic;
    GT18_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt18_cpllfbclklost_out                  : out  std_logic;
    gt18_cplllock_out                       : out  std_logic;
    gt18_cplllockdetclk_in                  : in   std_logic;
    gt18_cpllrefclklost_out                 : out  std_logic;
    gt18_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt18_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt18_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt18_drpclk_in                          : in   std_logic;
    gt18_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt18_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt18_drpen_in                           : in   std_logic;
    gt18_drprdy_out                         : out  std_logic;
    gt18_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt18_eyescanreset_in                    : in   std_logic;
    gt18_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt18_eyescandataerror_out               : out  std_logic;
    gt18_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt18_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt18_rxusrclk_in                        : in   std_logic;
    gt18_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt18_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt18_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt18_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt18_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt18_rxbyteisaligned_out                : out  std_logic;
    gt18_rxmcommaalignen_in                 : in   std_logic;
    gt18_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt18_rxdfeagchold_in                    : in   std_logic;
    gt18_rxdfelfhold_in                     : in   std_logic;
    gt18_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt18_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt18_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt18_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt18_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt18_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt18_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt18_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt18_gttxreset_in                       : in   std_logic;
    gt18_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt18_txusrclk_in                        : in   std_logic;
    gt18_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt18_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt18_gthtxn_out                         : out  std_logic;
    gt18_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt18_txoutclk_out                       : out  std_logic;
    gt18_txoutclkfabric_out                 : out  std_logic;
    gt18_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt18_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt18_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt18_txcharisk_in                       : in   std_logic_vector(3 downto 0);
   
    --_________________________________________________________________________
    --_________________________________________________________________________
    --GT19  (X1Y27)
    --____________________________CHANNEL PORTS________________________________
    GT19_RXPMARESETDONE_OUT                        : out  std_logic;
    GT19_TXPMARESETDONE_OUT                        : out  std_logic;

    --------------------------------- CPLL Ports -------------------------------
    gt19_cpllfbclklost_out                  : out  std_logic;
    gt19_cplllock_out                       : out  std_logic;
    gt19_cplllockdetclk_in                  : in   std_logic;
    gt19_cpllrefclklost_out                 : out  std_logic;
    gt19_cpllreset_in                       : in   std_logic;
    -------------------------- Channel - Clocking Ports ------------------------
    gt19_gtrefclk0_in                       : in   std_logic;
    ---------------------------- Channel - DRP Ports  --------------------------
    gt19_drpaddr_in                         : in   std_logic_vector(8 downto 0);
    gt19_drpclk_in                          : in   std_logic;
    gt19_drpdi_in                           : in   std_logic_vector(15 downto 0);
    gt19_drpdo_out                          : out  std_logic_vector(15 downto 0);
    gt19_drpen_in                           : in   std_logic;
    gt19_drprdy_out                         : out  std_logic;
    gt19_drpwe_in                           : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt19_eyescanreset_in                    : in   std_logic;
    gt19_rxuserrdy_in                       : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt19_eyescandataerror_out               : out  std_logic;
    gt19_eyescantrigger_in                  : in   std_logic;
    ------------------- Receive Ports - Digital Monitor Ports ------------------
    gt19_dmonitorout_out                    : out  std_logic_vector(14 downto 0);
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt19_rxusrclk_in                        : in   std_logic;
    gt19_rxusrclk2_in                       : in   std_logic;
    ------------------ Receive Ports - FPGA RX interface Ports -----------------
    gt19_rxdata_out                         : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt19_rxdisperr_out                      : out  std_logic_vector(3 downto 0);
    gt19_rxnotintable_out                   : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt19_gthrxn_in                          : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt19_rxbyteisaligned_out                : out  std_logic;
    gt19_rxmcommaalignen_in                 : in   std_logic;
    gt19_rxpcommaalignen_in                 : in   std_logic;
    --------------------- Receive Ports - RX Equalizer Ports -------------------
    gt19_rxdfeagchold_in                    : in   std_logic;
    gt19_rxdfelfhold_in                     : in   std_logic;
    gt19_rxmonitorout_out                   : out  std_logic_vector(6 downto 0);
    gt19_rxmonitorsel_in                    : in   std_logic_vector(1 downto 0);
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt19_rxoutclk_out                       : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt19_gtrxreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt19_rxpolarity_in                      : in   std_logic;
    ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    gt19_rxcharisk_out                      : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports -RX AFE Ports -----------------------
    gt19_gthrxp_in                          : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt19_rxresetdone_out                    : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt19_gttxreset_in                       : in   std_logic;
    gt19_txuserrdy_in                       : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt19_txusrclk_in                        : in   std_logic;
    gt19_txusrclk2_in                       : in   std_logic;
    ------------------ Transmit Ports - TX Data Path interface -----------------
    gt19_txdata_in                          : in   std_logic_vector(31 downto 0);
    ---------------- Transmit Ports - TX Driver and OOB signaling --------------
    gt19_gthtxn_out                         : out  std_logic;
    gt19_gthtxp_out                         : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt19_txoutclk_out                       : out  std_logic;
    gt19_txoutclkfabric_out                 : out  std_logic;
    gt19_txoutclkpcs_out                    : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt19_txresetdone_out                    : out  std_logic;
    ----------------- Transmit Ports - TX Polarity Control Ports ---------------
    gt19_txpolarity_in                      : in   std_logic;
    ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
    gt19_txcharisk_in                       : in   std_logic_vector(3 downto 0);
   

    --____________________________COMMON PORTS________________________________
     GT0_QPLLOUTCLK_IN   : in std_logic;
     GT0_QPLLOUTREFCLK_IN   : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT1_QPLLOUTCLK_IN   : in std_logic;
     GT1_QPLLOUTREFCLK_IN   : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT2_QPLLOUTCLK_IN   : in std_logic;
     GT2_QPLLOUTREFCLK_IN   : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT3_QPLLOUTCLK_IN   : in std_logic;
     GT3_QPLLOUTREFCLK_IN   : in std_logic;
    --____________________________COMMON PORTS________________________________
     GT4_QPLLOUTCLK_IN   : in std_logic;
     GT4_QPLLOUTREFCLK_IN   : in std_logic

);
end component;

component gt625_fab20_TX_STARTUP_FSM
  Generic(
           EXAMPLE_SIMULATION       : integer := 0;
           STABLE_CLOCK_PERIOD      : integer range 4 to 250 := 8; --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   : integer range 2 to 8  := 8; 
           TX_QPLL_USED             : boolean := False;           -- the TX and RX Reset FSMs must
           RX_QPLL_USED             : boolean := False;           -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   : boolean := True             -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                  -- is enough. For single-lane applications the automatic alignment is 
                                                                  -- sufficient              
         );     
    Port ( STABLE_CLOCK             : in  STD_LOGIC;              --Stable Clock, either a stable clock from the PCB
                                                                  --or reference-clock present at startup.
           TXUSERCLK                : in  STD_LOGIC;              --TXUSERCLK as used in the design
           SOFT_RESET               : in  STD_LOGIC;              --User Reset, can be pulled any time
           QPLLREFCLKLOST           : in  STD_LOGIC;              --QPLL Reference-clock for the GT is lost
           CPLLREFCLKLOST           : in  STD_LOGIC;              --CPLL Reference-clock for the GT is lost
           QPLLLOCK                 : in  STD_LOGIC;              --Lock Detect from the QPLL of the GT
           CPLLLOCK                 : in  STD_LOGIC;              --Lock Detect from the CPLL of the GT
           TXRESETDONE              : in  STD_LOGIC;      
           MMCM_LOCK                : in  STD_LOGIC;      
           GTTXRESET                : out STD_LOGIC:='0';      
           MMCM_RESET               : out STD_LOGIC:='0';      
           QPLL_RESET               : out STD_LOGIC:='0';        --Reset QPLL
           CPLL_RESET               : out STD_LOGIC:='0';        --Reset CPLL
           TX_FSM_RESET_DONE        : out STD_LOGIC:='0';        --Reset-sequence has sucessfully been finished.
           TXUSERRDY                : out STD_LOGIC:='0';
           RUN_PHALIGNMENT          : out STD_LOGIC:='0';
           RESET_PHALIGNMENT        : out STD_LOGIC:='0';
           PHALIGNMENT_DONE         : in  STD_LOGIC;
           
           RETRY_COUNTER            : out  STD_LOGIC_VECTOR (RETRY_COUNTER_BITWIDTH-1 downto 0):=(others=>'0')-- Number of 
                                                            -- Retries it took to get the transceiver up and running
           );
end component;

component gt625_fab20_RX_STARTUP_FSM
  Generic(
           EXAMPLE_SIMULATION       : integer := 0;
           EQ_MODE                  : string := "DFE";
           STABLE_CLOCK_PERIOD      : integer range 4 to 250 := 8; --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   : integer range 2 to 8  := 8; 
           TX_QPLL_USED             : boolean := False;           -- the TX and RX Reset FSMs must
           RX_QPLL_USED             : boolean := False;           -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   : boolean := True             -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                  -- is enough. For single-lane applications the automatic alignment is 
                                                                  -- sufficient                         
         );     
    Port ( STABLE_CLOCK             : in  STD_LOGIC;        --Stable Clock, either a stable clock from the PCB
                                                            --or reference-clock present at startup.
           RXUSERCLK                : in  STD_LOGIC;        --RXUSERCLK as used in the design
           SOFT_RESET               : in  STD_LOGIC;        --User Reset, can be pulled any time
           RXPMARESETDONE               : in  STD_LOGIC;              
           RXOUTCLK               : in  STD_LOGIC; 
           TXPMARESETDONE               : in  STD_LOGIC;              
           TXOUTCLK               : in  STD_LOGIC; 
             
           QPLLREFCLKLOST           : in  STD_LOGIC;        --QPLL Reference-clock for the GT is lost
           CPLLREFCLKLOST           : in  STD_LOGIC;        --CPLL Reference-clock for the GT is lost
           QPLLLOCK                 : in  STD_LOGIC;        --Lock Detect from the QPLL of the GT
           CPLLLOCK                 : in  STD_LOGIC;        --Lock Detect from the CPLL of the GT
           RXRESETDONE              : in  STD_LOGIC;
           MMCM_LOCK                : in  STD_LOGIC;
           RECCLK_STABLE            : in  STD_LOGIC;
           RECCLK_MONITOR_RESTART   : in  STD_LOGIC;
           DATA_VALID               : in  STD_LOGIC;
           TXUSERRDY                : in  STD_LOGIC;       --TXUSERRDY from GT 
           DONT_RESET_ON_DATA_ERROR : in  STD_LOGIC;
           GTRXRESET                : out STD_LOGIC:='0';
           MMCM_RESET               : out STD_LOGIC:='0';
           QPLL_RESET               : out STD_LOGIC:='0';  --Reset QPLL (only if RX uses QPLL)
           CPLL_RESET               : out STD_LOGIC:='0';  --Reset CPLL (only if RX uses CPLL)
           RX_FSM_RESET_DONE        : out STD_LOGIC:='0';  --Reset-sequence has sucessfully been finished.
           RXUSERRDY                : out STD_LOGIC:='0';
           RUN_PHALIGNMENT          : out STD_LOGIC;
           PHALIGNMENT_DONE         : in  STD_LOGIC; 
           RESET_PHALIGNMENT        : out STD_LOGIC:='0';           
           RXDFEAGCHOLD             : out STD_LOGIC;
           RXDFELFHOLD              : out STD_LOGIC;
           RXLPMLFHOLD              : out STD_LOGIC;
           RXLPMHFHOLD              : out STD_LOGIC;
           RETRY_COUNTER            : out STD_LOGIC_VECTOR (RETRY_COUNTER_BITWIDTH-1 downto 0):=(others=>'0')-- Number of 
                                                            -- Retries it took to get the transceiver up and running
           );
end component;






  function get_cdrlock_time(is_sim : in integer) return integer is
    variable lock_time: integer;
  begin
    if (is_sim = 1) then
      lock_time := 1000;
    else
      lock_time := 50000 / integer(6.25); --Typical CDR lock time is 50,000UI as per DS183
    end if;
    return lock_time;
  end function;


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;
    constant RX_CDRLOCK_TIME      : integer := get_cdrlock_time(EXAMPLE_SIMULATION);       -- 200us
    constant WAIT_TIME_CDRLOCK    : integer := RX_CDRLOCK_TIME / STABLE_CLOCK_PERIOD;      -- 200 us time-out

    -------------------------- GT Wrapper Wires ------------------------------
    signal   gt0_txpmaresetdone_i            : std_logic;
    signal   gt0_rxpmaresetdone_i            : std_logic;
    signal   gt0_cpllreset_i                 : std_logic;
    signal   gt0_cpllreset_t                 : std_logic;
    signal   gt0_cpllrefclklost_i            : std_logic;
    signal   gt0_cplllock_i                  : std_logic;
    signal   gt0_txresetdone_i               : std_logic;
    signal   gt0_rxresetdone_i               : std_logic;
    signal   gt0_gttxreset_i                 : std_logic;
    signal   gt0_gttxreset_t                 : std_logic;
    signal   gt0_gtrxreset_i                 : std_logic;
    signal   gt0_gtrxreset_t                 : std_logic;
    signal   gt0_txuserrdy_i                 : std_logic;
    signal   gt0_txuserrdy_t                 : std_logic;
    signal   gt0_rxuserrdy_i                 : std_logic;
    signal   gt0_rxuserrdy_t                 : std_logic;

    signal   gt0_rxdfeagchold_i              : std_logic;
    signal   gt0_rxdfelfhold_i               : std_logic;
    signal   gt0_rxlpmlfhold_i               : std_logic;
    signal   gt0_rxlpmhfhold_i               : std_logic;


    signal   gt1_txpmaresetdone_i            : std_logic;
    signal   gt1_rxpmaresetdone_i            : std_logic;
    signal   gt1_cpllreset_i                 : std_logic;
    signal   gt1_cpllreset_t                 : std_logic;
    signal   gt1_cpllrefclklost_i            : std_logic;
    signal   gt1_cplllock_i                  : std_logic;
    signal   gt1_txresetdone_i               : std_logic;
    signal   gt1_rxresetdone_i               : std_logic;
    signal   gt1_gttxreset_i                 : std_logic;
    signal   gt1_gttxreset_t                 : std_logic;
    signal   gt1_gtrxreset_i                 : std_logic;
    signal   gt1_gtrxreset_t                 : std_logic;
    signal   gt1_txuserrdy_i                 : std_logic;
    signal   gt1_txuserrdy_t                 : std_logic;
    signal   gt1_rxuserrdy_i                 : std_logic;
    signal   gt1_rxuserrdy_t                 : std_logic;

    signal   gt1_rxdfeagchold_i              : std_logic;
    signal   gt1_rxdfelfhold_i               : std_logic;
    signal   gt1_rxlpmlfhold_i               : std_logic;
    signal   gt1_rxlpmhfhold_i               : std_logic;


    signal   gt2_txpmaresetdone_i            : std_logic;
    signal   gt2_rxpmaresetdone_i            : std_logic;
    signal   gt2_cpllreset_i                 : std_logic;
    signal   gt2_cpllreset_t                 : std_logic;
    signal   gt2_cpllrefclklost_i            : std_logic;
    signal   gt2_cplllock_i                  : std_logic;
    signal   gt2_txresetdone_i               : std_logic;
    signal   gt2_rxresetdone_i               : std_logic;
    signal   gt2_gttxreset_i                 : std_logic;
    signal   gt2_gttxreset_t                 : std_logic;
    signal   gt2_gtrxreset_i                 : std_logic;
    signal   gt2_gtrxreset_t                 : std_logic;
    signal   gt2_txuserrdy_i                 : std_logic;
    signal   gt2_txuserrdy_t                 : std_logic;
    signal   gt2_rxuserrdy_i                 : std_logic;
    signal   gt2_rxuserrdy_t                 : std_logic;

    signal   gt2_rxdfeagchold_i              : std_logic;
    signal   gt2_rxdfelfhold_i               : std_logic;
    signal   gt2_rxlpmlfhold_i               : std_logic;
    signal   gt2_rxlpmhfhold_i               : std_logic;


    signal   gt3_txpmaresetdone_i            : std_logic;
    signal   gt3_rxpmaresetdone_i            : std_logic;
    signal   gt3_cpllreset_i                 : std_logic;
    signal   gt3_cpllreset_t                 : std_logic;
    signal   gt3_cpllrefclklost_i            : std_logic;
    signal   gt3_cplllock_i                  : std_logic;
    signal   gt3_txresetdone_i               : std_logic;
    signal   gt3_rxresetdone_i               : std_logic;
    signal   gt3_gttxreset_i                 : std_logic;
    signal   gt3_gttxreset_t                 : std_logic;
    signal   gt3_gtrxreset_i                 : std_logic;
    signal   gt3_gtrxreset_t                 : std_logic;
    signal   gt3_txuserrdy_i                 : std_logic;
    signal   gt3_txuserrdy_t                 : std_logic;
    signal   gt3_rxuserrdy_i                 : std_logic;
    signal   gt3_rxuserrdy_t                 : std_logic;

    signal   gt3_rxdfeagchold_i              : std_logic;
    signal   gt3_rxdfelfhold_i               : std_logic;
    signal   gt3_rxlpmlfhold_i               : std_logic;
    signal   gt3_rxlpmhfhold_i               : std_logic;


    signal   gt4_txpmaresetdone_i            : std_logic;
    signal   gt4_rxpmaresetdone_i            : std_logic;
    signal   gt4_cpllreset_i                 : std_logic;
    signal   gt4_cpllreset_t                 : std_logic;
    signal   gt4_cpllrefclklost_i            : std_logic;
    signal   gt4_cplllock_i                  : std_logic;
    signal   gt4_txresetdone_i               : std_logic;
    signal   gt4_rxresetdone_i               : std_logic;
    signal   gt4_gttxreset_i                 : std_logic;
    signal   gt4_gttxreset_t                 : std_logic;
    signal   gt4_gtrxreset_i                 : std_logic;
    signal   gt4_gtrxreset_t                 : std_logic;
    signal   gt4_txuserrdy_i                 : std_logic;
    signal   gt4_txuserrdy_t                 : std_logic;
    signal   gt4_rxuserrdy_i                 : std_logic;
    signal   gt4_rxuserrdy_t                 : std_logic;

    signal   gt4_rxdfeagchold_i              : std_logic;
    signal   gt4_rxdfelfhold_i               : std_logic;
    signal   gt4_rxlpmlfhold_i               : std_logic;
    signal   gt4_rxlpmhfhold_i               : std_logic;


    signal   gt5_txpmaresetdone_i            : std_logic;
    signal   gt5_rxpmaresetdone_i            : std_logic;
    signal   gt5_cpllreset_i                 : std_logic;
    signal   gt5_cpllreset_t                 : std_logic;
    signal   gt5_cpllrefclklost_i            : std_logic;
    signal   gt5_cplllock_i                  : std_logic;
    signal   gt5_txresetdone_i               : std_logic;
    signal   gt5_rxresetdone_i               : std_logic;
    signal   gt5_gttxreset_i                 : std_logic;
    signal   gt5_gttxreset_t                 : std_logic;
    signal   gt5_gtrxreset_i                 : std_logic;
    signal   gt5_gtrxreset_t                 : std_logic;
    signal   gt5_txuserrdy_i                 : std_logic;
    signal   gt5_txuserrdy_t                 : std_logic;
    signal   gt5_rxuserrdy_i                 : std_logic;
    signal   gt5_rxuserrdy_t                 : std_logic;

    signal   gt5_rxdfeagchold_i              : std_logic;
    signal   gt5_rxdfelfhold_i               : std_logic;
    signal   gt5_rxlpmlfhold_i               : std_logic;
    signal   gt5_rxlpmhfhold_i               : std_logic;


    signal   gt6_txpmaresetdone_i            : std_logic;
    signal   gt6_rxpmaresetdone_i            : std_logic;
    signal   gt6_cpllreset_i                 : std_logic;
    signal   gt6_cpllreset_t                 : std_logic;
    signal   gt6_cpllrefclklost_i            : std_logic;
    signal   gt6_cplllock_i                  : std_logic;
    signal   gt6_txresetdone_i               : std_logic;
    signal   gt6_rxresetdone_i               : std_logic;
    signal   gt6_gttxreset_i                 : std_logic;
    signal   gt6_gttxreset_t                 : std_logic;
    signal   gt6_gtrxreset_i                 : std_logic;
    signal   gt6_gtrxreset_t                 : std_logic;
    signal   gt6_txuserrdy_i                 : std_logic;
    signal   gt6_txuserrdy_t                 : std_logic;
    signal   gt6_rxuserrdy_i                 : std_logic;
    signal   gt6_rxuserrdy_t                 : std_logic;

    signal   gt6_rxdfeagchold_i              : std_logic;
    signal   gt6_rxdfelfhold_i               : std_logic;
    signal   gt6_rxlpmlfhold_i               : std_logic;
    signal   gt6_rxlpmhfhold_i               : std_logic;


    signal   gt7_txpmaresetdone_i            : std_logic;
    signal   gt7_rxpmaresetdone_i            : std_logic;
    signal   gt7_cpllreset_i                 : std_logic;
    signal   gt7_cpllreset_t                 : std_logic;
    signal   gt7_cpllrefclklost_i            : std_logic;
    signal   gt7_cplllock_i                  : std_logic;
    signal   gt7_txresetdone_i               : std_logic;
    signal   gt7_rxresetdone_i               : std_logic;
    signal   gt7_gttxreset_i                 : std_logic;
    signal   gt7_gttxreset_t                 : std_logic;
    signal   gt7_gtrxreset_i                 : std_logic;
    signal   gt7_gtrxreset_t                 : std_logic;
    signal   gt7_txuserrdy_i                 : std_logic;
    signal   gt7_txuserrdy_t                 : std_logic;
    signal   gt7_rxuserrdy_i                 : std_logic;
    signal   gt7_rxuserrdy_t                 : std_logic;

    signal   gt7_rxdfeagchold_i              : std_logic;
    signal   gt7_rxdfelfhold_i               : std_logic;
    signal   gt7_rxlpmlfhold_i               : std_logic;
    signal   gt7_rxlpmhfhold_i               : std_logic;


    signal   gt8_txpmaresetdone_i            : std_logic;
    signal   gt8_rxpmaresetdone_i            : std_logic;
    signal   gt8_cpllreset_i                 : std_logic;
    signal   gt8_cpllreset_t                 : std_logic;
    signal   gt8_cpllrefclklost_i            : std_logic;
    signal   gt8_cplllock_i                  : std_logic;
    signal   gt8_txresetdone_i               : std_logic;
    signal   gt8_rxresetdone_i               : std_logic;
    signal   gt8_gttxreset_i                 : std_logic;
    signal   gt8_gttxreset_t                 : std_logic;
    signal   gt8_gtrxreset_i                 : std_logic;
    signal   gt8_gtrxreset_t                 : std_logic;
    signal   gt8_txuserrdy_i                 : std_logic;
    signal   gt8_txuserrdy_t                 : std_logic;
    signal   gt8_rxuserrdy_i                 : std_logic;
    signal   gt8_rxuserrdy_t                 : std_logic;

    signal   gt8_rxdfeagchold_i              : std_logic;
    signal   gt8_rxdfelfhold_i               : std_logic;
    signal   gt8_rxlpmlfhold_i               : std_logic;
    signal   gt8_rxlpmhfhold_i               : std_logic;


    signal   gt9_txpmaresetdone_i            : std_logic;
    signal   gt9_rxpmaresetdone_i            : std_logic;
    signal   gt9_cpllreset_i                 : std_logic;
    signal   gt9_cpllreset_t                 : std_logic;
    signal   gt9_cpllrefclklost_i            : std_logic;
    signal   gt9_cplllock_i                  : std_logic;
    signal   gt9_txresetdone_i               : std_logic;
    signal   gt9_rxresetdone_i               : std_logic;
    signal   gt9_gttxreset_i                 : std_logic;
    signal   gt9_gttxreset_t                 : std_logic;
    signal   gt9_gtrxreset_i                 : std_logic;
    signal   gt9_gtrxreset_t                 : std_logic;
    signal   gt9_txuserrdy_i                 : std_logic;
    signal   gt9_txuserrdy_t                 : std_logic;
    signal   gt9_rxuserrdy_i                 : std_logic;
    signal   gt9_rxuserrdy_t                 : std_logic;

    signal   gt9_rxdfeagchold_i              : std_logic;
    signal   gt9_rxdfelfhold_i               : std_logic;
    signal   gt9_rxlpmlfhold_i               : std_logic;
    signal   gt9_rxlpmhfhold_i               : std_logic;


    signal   gt10_txpmaresetdone_i           : std_logic;
    signal   gt10_rxpmaresetdone_i           : std_logic;
    signal   gt10_cpllreset_i                : std_logic;
    signal   gt10_cpllreset_t                : std_logic;
    signal   gt10_cpllrefclklost_i           : std_logic;
    signal   gt10_cplllock_i                 : std_logic;
    signal   gt10_txresetdone_i              : std_logic;
    signal   gt10_rxresetdone_i              : std_logic;
    signal   gt10_gttxreset_i                : std_logic;
    signal   gt10_gttxreset_t                : std_logic;
    signal   gt10_gtrxreset_i                : std_logic;
    signal   gt10_gtrxreset_t                : std_logic;
    signal   gt10_txuserrdy_i                : std_logic;
    signal   gt10_txuserrdy_t                : std_logic;
    signal   gt10_rxuserrdy_i                : std_logic;
    signal   gt10_rxuserrdy_t                : std_logic;

    signal   gt10_rxdfeagchold_i             : std_logic;
    signal   gt10_rxdfelfhold_i              : std_logic;
    signal   gt10_rxlpmlfhold_i              : std_logic;
    signal   gt10_rxlpmhfhold_i              : std_logic;


    signal   gt11_txpmaresetdone_i           : std_logic;
    signal   gt11_rxpmaresetdone_i           : std_logic;
    signal   gt11_cpllreset_i                : std_logic;
    signal   gt11_cpllreset_t                : std_logic;
    signal   gt11_cpllrefclklost_i           : std_logic;
    signal   gt11_cplllock_i                 : std_logic;
    signal   gt11_txresetdone_i              : std_logic;
    signal   gt11_rxresetdone_i              : std_logic;
    signal   gt11_gttxreset_i                : std_logic;
    signal   gt11_gttxreset_t                : std_logic;
    signal   gt11_gtrxreset_i                : std_logic;
    signal   gt11_gtrxreset_t                : std_logic;
    signal   gt11_txuserrdy_i                : std_logic;
    signal   gt11_txuserrdy_t                : std_logic;
    signal   gt11_rxuserrdy_i                : std_logic;
    signal   gt11_rxuserrdy_t                : std_logic;

    signal   gt11_rxdfeagchold_i             : std_logic;
    signal   gt11_rxdfelfhold_i              : std_logic;
    signal   gt11_rxlpmlfhold_i              : std_logic;
    signal   gt11_rxlpmhfhold_i              : std_logic;


    signal   gt12_txpmaresetdone_i           : std_logic;
    signal   gt12_rxpmaresetdone_i           : std_logic;
    signal   gt12_cpllreset_i                : std_logic;
    signal   gt12_cpllreset_t                : std_logic;
    signal   gt12_cpllrefclklost_i           : std_logic;
    signal   gt12_cplllock_i                 : std_logic;
    signal   gt12_txresetdone_i              : std_logic;
    signal   gt12_rxresetdone_i              : std_logic;
    signal   gt12_gttxreset_i                : std_logic;
    signal   gt12_gttxreset_t                : std_logic;
    signal   gt12_gtrxreset_i                : std_logic;
    signal   gt12_gtrxreset_t                : std_logic;
    signal   gt12_txuserrdy_i                : std_logic;
    signal   gt12_txuserrdy_t                : std_logic;
    signal   gt12_rxuserrdy_i                : std_logic;
    signal   gt12_rxuserrdy_t                : std_logic;

    signal   gt12_rxdfeagchold_i             : std_logic;
    signal   gt12_rxdfelfhold_i              : std_logic;
    signal   gt12_rxlpmlfhold_i              : std_logic;
    signal   gt12_rxlpmhfhold_i              : std_logic;


    signal   gt13_txpmaresetdone_i           : std_logic;
    signal   gt13_rxpmaresetdone_i           : std_logic;
    signal   gt13_cpllreset_i                : std_logic;
    signal   gt13_cpllreset_t                : std_logic;
    signal   gt13_cpllrefclklost_i           : std_logic;
    signal   gt13_cplllock_i                 : std_logic;
    signal   gt13_txresetdone_i              : std_logic;
    signal   gt13_rxresetdone_i              : std_logic;
    signal   gt13_gttxreset_i                : std_logic;
    signal   gt13_gttxreset_t                : std_logic;
    signal   gt13_gtrxreset_i                : std_logic;
    signal   gt13_gtrxreset_t                : std_logic;
    signal   gt13_txuserrdy_i                : std_logic;
    signal   gt13_txuserrdy_t                : std_logic;
    signal   gt13_rxuserrdy_i                : std_logic;
    signal   gt13_rxuserrdy_t                : std_logic;

    signal   gt13_rxdfeagchold_i             : std_logic;
    signal   gt13_rxdfelfhold_i              : std_logic;
    signal   gt13_rxlpmlfhold_i              : std_logic;
    signal   gt13_rxlpmhfhold_i              : std_logic;


    signal   gt14_txpmaresetdone_i           : std_logic;
    signal   gt14_rxpmaresetdone_i           : std_logic;
    signal   gt14_cpllreset_i                : std_logic;
    signal   gt14_cpllreset_t                : std_logic;
    signal   gt14_cpllrefclklost_i           : std_logic;
    signal   gt14_cplllock_i                 : std_logic;
    signal   gt14_txresetdone_i              : std_logic;
    signal   gt14_rxresetdone_i              : std_logic;
    signal   gt14_gttxreset_i                : std_logic;
    signal   gt14_gttxreset_t                : std_logic;
    signal   gt14_gtrxreset_i                : std_logic;
    signal   gt14_gtrxreset_t                : std_logic;
    signal   gt14_txuserrdy_i                : std_logic;
    signal   gt14_txuserrdy_t                : std_logic;
    signal   gt14_rxuserrdy_i                : std_logic;
    signal   gt14_rxuserrdy_t                : std_logic;

    signal   gt14_rxdfeagchold_i             : std_logic;
    signal   gt14_rxdfelfhold_i              : std_logic;
    signal   gt14_rxlpmlfhold_i              : std_logic;
    signal   gt14_rxlpmhfhold_i              : std_logic;


    signal   gt15_txpmaresetdone_i           : std_logic;
    signal   gt15_rxpmaresetdone_i           : std_logic;
    signal   gt15_cpllreset_i                : std_logic;
    signal   gt15_cpllreset_t                : std_logic;
    signal   gt15_cpllrefclklost_i           : std_logic;
    signal   gt15_cplllock_i                 : std_logic;
    signal   gt15_txresetdone_i              : std_logic;
    signal   gt15_rxresetdone_i              : std_logic;
    signal   gt15_gttxreset_i                : std_logic;
    signal   gt15_gttxreset_t                : std_logic;
    signal   gt15_gtrxreset_i                : std_logic;
    signal   gt15_gtrxreset_t                : std_logic;
    signal   gt15_txuserrdy_i                : std_logic;
    signal   gt15_txuserrdy_t                : std_logic;
    signal   gt15_rxuserrdy_i                : std_logic;
    signal   gt15_rxuserrdy_t                : std_logic;

    signal   gt15_rxdfeagchold_i             : std_logic;
    signal   gt15_rxdfelfhold_i              : std_logic;
    signal   gt15_rxlpmlfhold_i              : std_logic;
    signal   gt15_rxlpmhfhold_i              : std_logic;


    signal   gt16_txpmaresetdone_i           : std_logic;
    signal   gt16_rxpmaresetdone_i           : std_logic;
    signal   gt16_cpllreset_i                : std_logic;
    signal   gt16_cpllreset_t                : std_logic;
    signal   gt16_cpllrefclklost_i           : std_logic;
    signal   gt16_cplllock_i                 : std_logic;
    signal   gt16_txresetdone_i              : std_logic;
    signal   gt16_rxresetdone_i              : std_logic;
    signal   gt16_gttxreset_i                : std_logic;
    signal   gt16_gttxreset_t                : std_logic;
    signal   gt16_gtrxreset_i                : std_logic;
    signal   gt16_gtrxreset_t                : std_logic;
    signal   gt16_txuserrdy_i                : std_logic;
    signal   gt16_txuserrdy_t                : std_logic;
    signal   gt16_rxuserrdy_i                : std_logic;
    signal   gt16_rxuserrdy_t                : std_logic;

    signal   gt16_rxdfeagchold_i             : std_logic;
    signal   gt16_rxdfelfhold_i              : std_logic;
    signal   gt16_rxlpmlfhold_i              : std_logic;
    signal   gt16_rxlpmhfhold_i              : std_logic;


    signal   gt17_txpmaresetdone_i           : std_logic;
    signal   gt17_rxpmaresetdone_i           : std_logic;
    signal   gt17_cpllreset_i                : std_logic;
    signal   gt17_cpllreset_t                : std_logic;
    signal   gt17_cpllrefclklost_i           : std_logic;
    signal   gt17_cplllock_i                 : std_logic;
    signal   gt17_txresetdone_i              : std_logic;
    signal   gt17_rxresetdone_i              : std_logic;
    signal   gt17_gttxreset_i                : std_logic;
    signal   gt17_gttxreset_t                : std_logic;
    signal   gt17_gtrxreset_i                : std_logic;
    signal   gt17_gtrxreset_t                : std_logic;
    signal   gt17_txuserrdy_i                : std_logic;
    signal   gt17_txuserrdy_t                : std_logic;
    signal   gt17_rxuserrdy_i                : std_logic;
    signal   gt17_rxuserrdy_t                : std_logic;

    signal   gt17_rxdfeagchold_i             : std_logic;
    signal   gt17_rxdfelfhold_i              : std_logic;
    signal   gt17_rxlpmlfhold_i              : std_logic;
    signal   gt17_rxlpmhfhold_i              : std_logic;


    signal   gt18_txpmaresetdone_i           : std_logic;
    signal   gt18_rxpmaresetdone_i           : std_logic;
    signal   gt18_cpllreset_i                : std_logic;
    signal   gt18_cpllreset_t                : std_logic;
    signal   gt18_cpllrefclklost_i           : std_logic;
    signal   gt18_cplllock_i                 : std_logic;
    signal   gt18_txresetdone_i              : std_logic;
    signal   gt18_rxresetdone_i              : std_logic;
    signal   gt18_gttxreset_i                : std_logic;
    signal   gt18_gttxreset_t                : std_logic;
    signal   gt18_gtrxreset_i                : std_logic;
    signal   gt18_gtrxreset_t                : std_logic;
    signal   gt18_txuserrdy_i                : std_logic;
    signal   gt18_txuserrdy_t                : std_logic;
    signal   gt18_rxuserrdy_i                : std_logic;
    signal   gt18_rxuserrdy_t                : std_logic;

    signal   gt18_rxdfeagchold_i             : std_logic;
    signal   gt18_rxdfelfhold_i              : std_logic;
    signal   gt18_rxlpmlfhold_i              : std_logic;
    signal   gt18_rxlpmhfhold_i              : std_logic;


    signal   gt19_txpmaresetdone_i           : std_logic;
    signal   gt19_rxpmaresetdone_i           : std_logic;
    signal   gt19_cpllreset_i                : std_logic;
    signal   gt19_cpllreset_t                : std_logic;
    signal   gt19_cpllrefclklost_i           : std_logic;
    signal   gt19_cplllock_i                 : std_logic;
    signal   gt19_txresetdone_i              : std_logic;
    signal   gt19_rxresetdone_i              : std_logic;
    signal   gt19_gttxreset_i                : std_logic;
    signal   gt19_gttxreset_t                : std_logic;
    signal   gt19_gtrxreset_i                : std_logic;
    signal   gt19_gtrxreset_t                : std_logic;
    signal   gt19_txuserrdy_i                : std_logic;
    signal   gt19_txuserrdy_t                : std_logic;
    signal   gt19_rxuserrdy_i                : std_logic;
    signal   gt19_rxuserrdy_t                : std_logic;

    signal   gt19_rxdfeagchold_i             : std_logic;
    signal   gt19_rxdfelfhold_i              : std_logic;
    signal   gt19_rxlpmlfhold_i              : std_logic;
    signal   gt19_rxlpmhfhold_i              : std_logic;



    signal   gt0_qpllreset_i                 : std_logic;
    signal   gt0_qpllreset_t                 : std_logic;
    signal   gt0_qpllrefclklost_i            : std_logic;
    signal   gt0_qplllock_i                  : std_logic;
    signal   gt1_qpllreset_i                 : std_logic;
    signal   gt1_qpllreset_t                 : std_logic;
    signal   gt1_qpllrefclklost_i            : std_logic;
    signal   gt1_qplllock_i                  : std_logic;
    signal   gt2_qpllreset_i                 : std_logic;
    signal   gt2_qpllreset_t                 : std_logic;
    signal   gt2_qpllrefclklost_i            : std_logic;
    signal   gt2_qplllock_i                  : std_logic;
    signal   gt3_qpllreset_i                 : std_logic;
    signal   gt3_qpllreset_t                 : std_logic;
    signal   gt3_qpllrefclklost_i            : std_logic;
    signal   gt3_qplllock_i                  : std_logic;
    signal   gt4_qpllreset_i                 : std_logic;
    signal   gt4_qpllreset_t                 : std_logic;
    signal   gt4_qpllrefclklost_i            : std_logic;
    signal   gt4_qplllock_i                  : std_logic;


    ------------------------------- Global Signals -----------------------------
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_vcc_i                   : std_logic;

    signal   gt0_txoutclk_i                  : std_logic;
    signal   gt0_rxoutclk_i                  : std_logic;
    signal   gt0_rxoutclk_i2                 : std_logic;
    signal   gt0_txoutclk_i2                 : std_logic;
    signal   gt0_recclk_stable_i             : std_logic;
    signal   gt0_rx_cdrlocked                : std_logic;
    signal   gt0_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt1_txoutclk_i                  : std_logic;
    signal   gt1_rxoutclk_i                  : std_logic;
    signal   gt1_rxoutclk_i2                 : std_logic;
    signal   gt1_txoutclk_i2                 : std_logic;
    signal   gt1_recclk_stable_i             : std_logic;
    signal   gt1_rx_cdrlocked                : std_logic;
    signal   gt1_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt2_txoutclk_i                  : std_logic;
    signal   gt2_rxoutclk_i                  : std_logic;
    signal   gt2_rxoutclk_i2                 : std_logic;
    signal   gt2_txoutclk_i2                 : std_logic;
    signal   gt2_recclk_stable_i             : std_logic;
    signal   gt2_rx_cdrlocked                : std_logic;
    signal   gt2_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt3_txoutclk_i                  : std_logic;
    signal   gt3_rxoutclk_i                  : std_logic;
    signal   gt3_rxoutclk_i2                 : std_logic;
    signal   gt3_txoutclk_i2                 : std_logic;
    signal   gt3_recclk_stable_i             : std_logic;
    signal   gt3_rx_cdrlocked                : std_logic;
    signal   gt3_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt4_txoutclk_i                  : std_logic;
    signal   gt4_rxoutclk_i                  : std_logic;
    signal   gt4_rxoutclk_i2                 : std_logic;
    signal   gt4_txoutclk_i2                 : std_logic;
    signal   gt4_recclk_stable_i             : std_logic;
    signal   gt4_rx_cdrlocked                : std_logic;
    signal   gt4_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt5_txoutclk_i                  : std_logic;
    signal   gt5_rxoutclk_i                  : std_logic;
    signal   gt5_rxoutclk_i2                 : std_logic;
    signal   gt5_txoutclk_i2                 : std_logic;
    signal   gt5_recclk_stable_i             : std_logic;
    signal   gt5_rx_cdrlocked                : std_logic;
    signal   gt5_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt6_txoutclk_i                  : std_logic;
    signal   gt6_rxoutclk_i                  : std_logic;
    signal   gt6_rxoutclk_i2                 : std_logic;
    signal   gt6_txoutclk_i2                 : std_logic;
    signal   gt6_recclk_stable_i             : std_logic;
    signal   gt6_rx_cdrlocked                : std_logic;
    signal   gt6_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt7_txoutclk_i                  : std_logic;
    signal   gt7_rxoutclk_i                  : std_logic;
    signal   gt7_rxoutclk_i2                 : std_logic;
    signal   gt7_txoutclk_i2                 : std_logic;
    signal   gt7_recclk_stable_i             : std_logic;
    signal   gt7_rx_cdrlocked                : std_logic;
    signal   gt7_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt8_txoutclk_i                  : std_logic;
    signal   gt8_rxoutclk_i                  : std_logic;
    signal   gt8_rxoutclk_i2                 : std_logic;
    signal   gt8_txoutclk_i2                 : std_logic;
    signal   gt8_recclk_stable_i             : std_logic;
    signal   gt8_rx_cdrlocked                : std_logic;
    signal   gt8_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt9_txoutclk_i                  : std_logic;
    signal   gt9_rxoutclk_i                  : std_logic;
    signal   gt9_rxoutclk_i2                 : std_logic;
    signal   gt9_txoutclk_i2                 : std_logic;
    signal   gt9_recclk_stable_i             : std_logic;
    signal   gt9_rx_cdrlocked                : std_logic;
    signal   gt9_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt10_txoutclk_i                 : std_logic;
    signal   gt10_rxoutclk_i                 : std_logic;
    signal   gt10_rxoutclk_i2                : std_logic;
    signal   gt10_txoutclk_i2                : std_logic;
    signal   gt10_recclk_stable_i            : std_logic;
    signal   gt10_rx_cdrlocked               : std_logic;
    signal   gt10_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt11_txoutclk_i                 : std_logic;
    signal   gt11_rxoutclk_i                 : std_logic;
    signal   gt11_rxoutclk_i2                : std_logic;
    signal   gt11_txoutclk_i2                : std_logic;
    signal   gt11_recclk_stable_i            : std_logic;
    signal   gt11_rx_cdrlocked               : std_logic;
    signal   gt11_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt12_txoutclk_i                 : std_logic;
    signal   gt12_rxoutclk_i                 : std_logic;
    signal   gt12_rxoutclk_i2                : std_logic;
    signal   gt12_txoutclk_i2                : std_logic;
    signal   gt12_recclk_stable_i            : std_logic;
    signal   gt12_rx_cdrlocked               : std_logic;
    signal   gt12_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt13_txoutclk_i                 : std_logic;
    signal   gt13_rxoutclk_i                 : std_logic;
    signal   gt13_rxoutclk_i2                : std_logic;
    signal   gt13_txoutclk_i2                : std_logic;
    signal   gt13_recclk_stable_i            : std_logic;
    signal   gt13_rx_cdrlocked               : std_logic;
    signal   gt13_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt14_txoutclk_i                 : std_logic;
    signal   gt14_rxoutclk_i                 : std_logic;
    signal   gt14_rxoutclk_i2                : std_logic;
    signal   gt14_txoutclk_i2                : std_logic;
    signal   gt14_recclk_stable_i            : std_logic;
    signal   gt14_rx_cdrlocked               : std_logic;
    signal   gt14_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt15_txoutclk_i                 : std_logic;
    signal   gt15_rxoutclk_i                 : std_logic;
    signal   gt15_rxoutclk_i2                : std_logic;
    signal   gt15_txoutclk_i2                : std_logic;
    signal   gt15_recclk_stable_i            : std_logic;
    signal   gt15_rx_cdrlocked               : std_logic;
    signal   gt15_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt16_txoutclk_i                 : std_logic;
    signal   gt16_rxoutclk_i                 : std_logic;
    signal   gt16_rxoutclk_i2                : std_logic;
    signal   gt16_txoutclk_i2                : std_logic;
    signal   gt16_recclk_stable_i            : std_logic;
    signal   gt16_rx_cdrlocked               : std_logic;
    signal   gt16_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt17_txoutclk_i                 : std_logic;
    signal   gt17_rxoutclk_i                 : std_logic;
    signal   gt17_rxoutclk_i2                : std_logic;
    signal   gt17_txoutclk_i2                : std_logic;
    signal   gt17_recclk_stable_i            : std_logic;
    signal   gt17_rx_cdrlocked               : std_logic;
    signal   gt17_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt18_txoutclk_i                 : std_logic;
    signal   gt18_rxoutclk_i                 : std_logic;
    signal   gt18_rxoutclk_i2                : std_logic;
    signal   gt18_txoutclk_i2                : std_logic;
    signal   gt18_recclk_stable_i            : std_logic;
    signal   gt18_rx_cdrlocked               : std_logic;
    signal   gt18_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;

    signal   gt19_txoutclk_i                 : std_logic;
    signal   gt19_rxoutclk_i                 : std_logic;
    signal   gt19_rxoutclk_i2                : std_logic;
    signal   gt19_txoutclk_i2                : std_logic;
    signal   gt19_recclk_stable_i            : std_logic;
    signal   gt19_rx_cdrlocked               : std_logic;
    signal   gt19_rx_cdrlock_counter  :   integer range 0 to WAIT_TIME_CDRLOCK:= 0 ;






    signal      rx_cdrlocked                    : std_logic;


 


--**************************** Main Body of Code *******************************
begin
    --  Static signal Assigments
    tied_to_ground_i                             <= '0';
    tied_to_vcc_i                                <= '1';

    ----------------------------- The GT Wrapper -----------------------------
    
    -- Use the instantiation template in the example directory to add the GT wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.


    gt625_fab20_i : gt625_fab20_multi_gt
    generic map
    (
        EXAMPLE_SIMULATION              =>      EXAMPLE_SIMULATION,
        WRAPPER_SIM_GTRESET_SPEEDUP     =>      EXAMPLE_SIM_GTRESET_SPEEDUP
    )
    port map
    (
        GT0_RXPMARESETDONE_OUT          =>      gt0_rxpmaresetdone_i,
        GT0_TXPMARESETDONE_OUT          =>      gt0_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT0  (X1Y8)

        --------------------------------- CPLL Ports -------------------------------
        gt0_cpllfbclklost_out           =>      gt0_cpllfbclklost_out,
        gt0_cplllock_out                =>      gt0_cplllock_i,
        gt0_cplllockdetclk_in           =>      gt0_cplllockdetclk_in,
        gt0_cpllrefclklost_out          =>      gt0_cpllrefclklost_i,
        gt0_cpllreset_in                =>      gt0_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt0_gtrefclk0_in                =>      gt0_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt0_drpaddr_in                  =>      gt0_drpaddr_in,
        gt0_drpclk_in                   =>      gt0_drpclk_in,
        gt0_drpdi_in                    =>      gt0_drpdi_in,
        gt0_drpdo_out                   =>      gt0_drpdo_out,
        gt0_drpen_in                    =>      gt0_drpen_in,
        gt0_drprdy_out                  =>      gt0_drprdy_out,
        gt0_drpwe_in                    =>      gt0_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt0_eyescanreset_in             =>      gt0_eyescanreset_in,
        gt0_rxuserrdy_in                =>      gt0_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt0_eyescandataerror_out        =>      gt0_eyescandataerror_out,
        gt0_eyescantrigger_in           =>      gt0_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt0_dmonitorout_out             =>      gt0_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt0_rxusrclk_in                 =>      gt0_rxusrclk_in,
        gt0_rxusrclk2_in                =>      gt0_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt0_rxdata_out                  =>      gt0_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt0_rxdisperr_out               =>      gt0_rxdisperr_out,
        gt0_rxnotintable_out            =>      gt0_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt0_gthrxn_in                   =>      gt0_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt0_rxbyteisaligned_out         =>      gt0_rxbyteisaligned_out,
        gt0_rxmcommaalignen_in          =>      gt0_rxmcommaalignen_in,
        gt0_rxpcommaalignen_in          =>      gt0_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt0_rxdfeagchold_in             =>      gt0_rxdfeagchold_i,
        gt0_rxdfelfhold_in              =>      gt0_rxdfelfhold_i,
        gt0_rxmonitorout_out            =>      gt0_rxmonitorout_out,
        gt0_rxmonitorsel_in             =>      gt0_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt0_rxoutclk_out                =>      gt0_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt0_gtrxreset_in                =>      gt0_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt0_rxpolarity_in               =>      gt0_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt0_rxcharisk_out               =>      gt0_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt0_gthrxp_in                   =>      gt0_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt0_rxresetdone_out             =>      gt0_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt0_gttxreset_in                =>      gt0_gttxreset_i,
        gt0_txuserrdy_in                =>      gt0_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt0_txusrclk_in                 =>      gt0_txusrclk_in,
        gt0_txusrclk2_in                =>      gt0_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt0_txdata_in                   =>      gt0_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt0_gthtxn_out                  =>      gt0_gthtxn_out,
        gt0_gthtxp_out                  =>      gt0_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt0_txoutclk_out                =>      gt0_txoutclk_i,
        gt0_txoutclkfabric_out          =>      gt0_txoutclkfabric_out,
        gt0_txoutclkpcs_out             =>      gt0_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt0_txresetdone_out             =>      gt0_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt0_txpolarity_in               =>      gt0_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt0_txcharisk_in                =>      gt0_txcharisk_in,


        GT1_RXPMARESETDONE_OUT          =>      gt1_rxpmaresetdone_i,
        GT1_TXPMARESETDONE_OUT          =>      gt1_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT1  (X1Y9)

        --------------------------------- CPLL Ports -------------------------------
        gt1_cpllfbclklost_out           =>      gt1_cpllfbclklost_out,
        gt1_cplllock_out                =>      gt1_cplllock_i,
        gt1_cplllockdetclk_in           =>      gt1_cplllockdetclk_in,
        gt1_cpllrefclklost_out          =>      gt1_cpllrefclklost_i,
        gt1_cpllreset_in                =>      gt1_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt1_gtrefclk0_in                =>      gt1_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt1_drpaddr_in                  =>      gt1_drpaddr_in,
        gt1_drpclk_in                   =>      gt1_drpclk_in,
        gt1_drpdi_in                    =>      gt1_drpdi_in,
        gt1_drpdo_out                   =>      gt1_drpdo_out,
        gt1_drpen_in                    =>      gt1_drpen_in,
        gt1_drprdy_out                  =>      gt1_drprdy_out,
        gt1_drpwe_in                    =>      gt1_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt1_eyescanreset_in             =>      gt1_eyescanreset_in,
        gt1_rxuserrdy_in                =>      gt1_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt1_eyescandataerror_out        =>      gt1_eyescandataerror_out,
        gt1_eyescantrigger_in           =>      gt1_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt1_dmonitorout_out             =>      gt1_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt1_rxusrclk_in                 =>      gt1_rxusrclk_in,
        gt1_rxusrclk2_in                =>      gt1_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt1_rxdata_out                  =>      gt1_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt1_rxdisperr_out               =>      gt1_rxdisperr_out,
        gt1_rxnotintable_out            =>      gt1_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt1_gthrxn_in                   =>      gt1_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt1_rxbyteisaligned_out         =>      gt1_rxbyteisaligned_out,
        gt1_rxmcommaalignen_in          =>      gt1_rxmcommaalignen_in,
        gt1_rxpcommaalignen_in          =>      gt1_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt1_rxdfeagchold_in             =>      gt1_rxdfeagchold_i,
        gt1_rxdfelfhold_in              =>      gt1_rxdfelfhold_i,
        gt1_rxmonitorout_out            =>      gt1_rxmonitorout_out,
        gt1_rxmonitorsel_in             =>      gt1_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt1_rxoutclk_out                =>      gt1_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt1_gtrxreset_in                =>      gt1_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt1_rxpolarity_in               =>      gt1_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt1_rxcharisk_out               =>      gt1_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt1_gthrxp_in                   =>      gt1_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt1_rxresetdone_out             =>      gt1_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt1_gttxreset_in                =>      gt1_gttxreset_i,
        gt1_txuserrdy_in                =>      gt1_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt1_txusrclk_in                 =>      gt1_txusrclk_in,
        gt1_txusrclk2_in                =>      gt1_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt1_txdata_in                   =>      gt1_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt1_gthtxn_out                  =>      gt1_gthtxn_out,
        gt1_gthtxp_out                  =>      gt1_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt1_txoutclk_out                =>      gt1_txoutclk_i,
        gt1_txoutclkfabric_out          =>      gt1_txoutclkfabric_out,
        gt1_txoutclkpcs_out             =>      gt1_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt1_txresetdone_out             =>      gt1_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt1_txpolarity_in               =>      gt1_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt1_txcharisk_in                =>      gt1_txcharisk_in,


        GT2_RXPMARESETDONE_OUT          =>      gt2_rxpmaresetdone_i,
        GT2_TXPMARESETDONE_OUT          =>      gt2_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT2  (X1Y10)

        --------------------------------- CPLL Ports -------------------------------
        gt2_cpllfbclklost_out           =>      gt2_cpllfbclklost_out,
        gt2_cplllock_out                =>      gt2_cplllock_i,
        gt2_cplllockdetclk_in           =>      gt2_cplllockdetclk_in,
        gt2_cpllrefclklost_out          =>      gt2_cpllrefclklost_i,
        gt2_cpllreset_in                =>      gt2_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt2_gtrefclk0_in                =>      gt2_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt2_drpaddr_in                  =>      gt2_drpaddr_in,
        gt2_drpclk_in                   =>      gt2_drpclk_in,
        gt2_drpdi_in                    =>      gt2_drpdi_in,
        gt2_drpdo_out                   =>      gt2_drpdo_out,
        gt2_drpen_in                    =>      gt2_drpen_in,
        gt2_drprdy_out                  =>      gt2_drprdy_out,
        gt2_drpwe_in                    =>      gt2_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt2_eyescanreset_in             =>      gt2_eyescanreset_in,
        gt2_rxuserrdy_in                =>      gt2_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt2_eyescandataerror_out        =>      gt2_eyescandataerror_out,
        gt2_eyescantrigger_in           =>      gt2_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt2_dmonitorout_out             =>      gt2_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt2_rxusrclk_in                 =>      gt2_rxusrclk_in,
        gt2_rxusrclk2_in                =>      gt2_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt2_rxdata_out                  =>      gt2_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt2_rxdisperr_out               =>      gt2_rxdisperr_out,
        gt2_rxnotintable_out            =>      gt2_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt2_gthrxn_in                   =>      gt2_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt2_rxbyteisaligned_out         =>      gt2_rxbyteisaligned_out,
        gt2_rxmcommaalignen_in          =>      gt2_rxmcommaalignen_in,
        gt2_rxpcommaalignen_in          =>      gt2_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt2_rxdfeagchold_in             =>      gt2_rxdfeagchold_i,
        gt2_rxdfelfhold_in              =>      gt2_rxdfelfhold_i,
        gt2_rxmonitorout_out            =>      gt2_rxmonitorout_out,
        gt2_rxmonitorsel_in             =>      gt2_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt2_rxoutclk_out                =>      gt2_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt2_gtrxreset_in                =>      gt2_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt2_rxpolarity_in               =>      gt2_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt2_rxcharisk_out               =>      gt2_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt2_gthrxp_in                   =>      gt2_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt2_rxresetdone_out             =>      gt2_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt2_gttxreset_in                =>      gt2_gttxreset_i,
        gt2_txuserrdy_in                =>      gt2_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt2_txusrclk_in                 =>      gt2_txusrclk_in,
        gt2_txusrclk2_in                =>      gt2_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt2_txdata_in                   =>      gt2_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt2_gthtxn_out                  =>      gt2_gthtxn_out,
        gt2_gthtxp_out                  =>      gt2_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt2_txoutclk_out                =>      gt2_txoutclk_i,
        gt2_txoutclkfabric_out          =>      gt2_txoutclkfabric_out,
        gt2_txoutclkpcs_out             =>      gt2_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt2_txresetdone_out             =>      gt2_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt2_txpolarity_in               =>      gt2_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt2_txcharisk_in                =>      gt2_txcharisk_in,


        GT3_RXPMARESETDONE_OUT          =>      gt3_rxpmaresetdone_i,
        GT3_TXPMARESETDONE_OUT          =>      gt3_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT3  (X1Y11)

        --------------------------------- CPLL Ports -------------------------------
        gt3_cpllfbclklost_out           =>      gt3_cpllfbclklost_out,
        gt3_cplllock_out                =>      gt3_cplllock_i,
        gt3_cplllockdetclk_in           =>      gt3_cplllockdetclk_in,
        gt3_cpllrefclklost_out          =>      gt3_cpllrefclklost_i,
        gt3_cpllreset_in                =>      gt3_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt3_gtrefclk0_in                =>      gt3_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt3_drpaddr_in                  =>      gt3_drpaddr_in,
        gt3_drpclk_in                   =>      gt3_drpclk_in,
        gt3_drpdi_in                    =>      gt3_drpdi_in,
        gt3_drpdo_out                   =>      gt3_drpdo_out,
        gt3_drpen_in                    =>      gt3_drpen_in,
        gt3_drprdy_out                  =>      gt3_drprdy_out,
        gt3_drpwe_in                    =>      gt3_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt3_eyescanreset_in             =>      gt3_eyescanreset_in,
        gt3_rxuserrdy_in                =>      gt3_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt3_eyescandataerror_out        =>      gt3_eyescandataerror_out,
        gt3_eyescantrigger_in           =>      gt3_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt3_dmonitorout_out             =>      gt3_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt3_rxusrclk_in                 =>      gt3_rxusrclk_in,
        gt3_rxusrclk2_in                =>      gt3_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt3_rxdata_out                  =>      gt3_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt3_rxdisperr_out               =>      gt3_rxdisperr_out,
        gt3_rxnotintable_out            =>      gt3_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt3_gthrxn_in                   =>      gt3_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt3_rxbyteisaligned_out         =>      gt3_rxbyteisaligned_out,
        gt3_rxmcommaalignen_in          =>      gt3_rxmcommaalignen_in,
        gt3_rxpcommaalignen_in          =>      gt3_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt3_rxdfeagchold_in             =>      gt3_rxdfeagchold_i,
        gt3_rxdfelfhold_in              =>      gt3_rxdfelfhold_i,
        gt3_rxmonitorout_out            =>      gt3_rxmonitorout_out,
        gt3_rxmonitorsel_in             =>      gt3_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt3_rxoutclk_out                =>      gt3_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt3_gtrxreset_in                =>      gt3_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt3_rxpolarity_in               =>      gt3_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt3_rxcharisk_out               =>      gt3_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt3_gthrxp_in                   =>      gt3_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt3_rxresetdone_out             =>      gt3_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt3_gttxreset_in                =>      gt3_gttxreset_i,
        gt3_txuserrdy_in                =>      gt3_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt3_txusrclk_in                 =>      gt3_txusrclk_in,
        gt3_txusrclk2_in                =>      gt3_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt3_txdata_in                   =>      gt3_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt3_gthtxn_out                  =>      gt3_gthtxn_out,
        gt3_gthtxp_out                  =>      gt3_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt3_txoutclk_out                =>      gt3_txoutclk_i,
        gt3_txoutclkfabric_out          =>      gt3_txoutclkfabric_out,
        gt3_txoutclkpcs_out             =>      gt3_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt3_txresetdone_out             =>      gt3_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt3_txpolarity_in               =>      gt3_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt3_txcharisk_in                =>      gt3_txcharisk_in,


        GT4_RXPMARESETDONE_OUT          =>      gt4_rxpmaresetdone_i,
        GT4_TXPMARESETDONE_OUT          =>      gt4_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT4  (X1Y12)

        --------------------------------- CPLL Ports -------------------------------
        gt4_cpllfbclklost_out           =>      gt4_cpllfbclklost_out,
        gt4_cplllock_out                =>      gt4_cplllock_i,
        gt4_cplllockdetclk_in           =>      gt4_cplllockdetclk_in,
        gt4_cpllrefclklost_out          =>      gt4_cpllrefclklost_i,
        gt4_cpllreset_in                =>      gt4_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt4_gtrefclk0_in                =>      gt4_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt4_drpaddr_in                  =>      gt4_drpaddr_in,
        gt4_drpclk_in                   =>      gt4_drpclk_in,
        gt4_drpdi_in                    =>      gt4_drpdi_in,
        gt4_drpdo_out                   =>      gt4_drpdo_out,
        gt4_drpen_in                    =>      gt4_drpen_in,
        gt4_drprdy_out                  =>      gt4_drprdy_out,
        gt4_drpwe_in                    =>      gt4_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt4_eyescanreset_in             =>      gt4_eyescanreset_in,
        gt4_rxuserrdy_in                =>      gt4_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt4_eyescandataerror_out        =>      gt4_eyescandataerror_out,
        gt4_eyescantrigger_in           =>      gt4_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt4_dmonitorout_out             =>      gt4_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt4_rxusrclk_in                 =>      gt4_rxusrclk_in,
        gt4_rxusrclk2_in                =>      gt4_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt4_rxdata_out                  =>      gt4_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt4_rxdisperr_out               =>      gt4_rxdisperr_out,
        gt4_rxnotintable_out            =>      gt4_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt4_gthrxn_in                   =>      gt4_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt4_rxbyteisaligned_out         =>      gt4_rxbyteisaligned_out,
        gt4_rxmcommaalignen_in          =>      gt4_rxmcommaalignen_in,
        gt4_rxpcommaalignen_in          =>      gt4_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt4_rxdfeagchold_in             =>      gt4_rxdfeagchold_i,
        gt4_rxdfelfhold_in              =>      gt4_rxdfelfhold_i,
        gt4_rxmonitorout_out            =>      gt4_rxmonitorout_out,
        gt4_rxmonitorsel_in             =>      gt4_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt4_rxoutclk_out                =>      gt4_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt4_gtrxreset_in                =>      gt4_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt4_rxpolarity_in               =>      gt4_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt4_rxcharisk_out               =>      gt4_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt4_gthrxp_in                   =>      gt4_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt4_rxresetdone_out             =>      gt4_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt4_gttxreset_in                =>      gt4_gttxreset_i,
        gt4_txuserrdy_in                =>      gt4_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt4_txusrclk_in                 =>      gt4_txusrclk_in,
        gt4_txusrclk2_in                =>      gt4_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt4_txdata_in                   =>      gt4_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt4_gthtxn_out                  =>      gt4_gthtxn_out,
        gt4_gthtxp_out                  =>      gt4_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt4_txoutclk_out                =>      gt4_txoutclk_i,
        gt4_txoutclkfabric_out          =>      gt4_txoutclkfabric_out,
        gt4_txoutclkpcs_out             =>      gt4_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt4_txresetdone_out             =>      gt4_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt4_txpolarity_in               =>      gt4_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt4_txcharisk_in                =>      gt4_txcharisk_in,


        GT5_RXPMARESETDONE_OUT          =>      gt5_rxpmaresetdone_i,
        GT5_TXPMARESETDONE_OUT          =>      gt5_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT5  (X1Y13)

        --------------------------------- CPLL Ports -------------------------------
        gt5_cpllfbclklost_out           =>      gt5_cpllfbclklost_out,
        gt5_cplllock_out                =>      gt5_cplllock_i,
        gt5_cplllockdetclk_in           =>      gt5_cplllockdetclk_in,
        gt5_cpllrefclklost_out          =>      gt5_cpllrefclklost_i,
        gt5_cpllreset_in                =>      gt5_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt5_gtrefclk0_in                =>      gt5_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt5_drpaddr_in                  =>      gt5_drpaddr_in,
        gt5_drpclk_in                   =>      gt5_drpclk_in,
        gt5_drpdi_in                    =>      gt5_drpdi_in,
        gt5_drpdo_out                   =>      gt5_drpdo_out,
        gt5_drpen_in                    =>      gt5_drpen_in,
        gt5_drprdy_out                  =>      gt5_drprdy_out,
        gt5_drpwe_in                    =>      gt5_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt5_eyescanreset_in             =>      gt5_eyescanreset_in,
        gt5_rxuserrdy_in                =>      gt5_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt5_eyescandataerror_out        =>      gt5_eyescandataerror_out,
        gt5_eyescantrigger_in           =>      gt5_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt5_dmonitorout_out             =>      gt5_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt5_rxusrclk_in                 =>      gt5_rxusrclk_in,
        gt5_rxusrclk2_in                =>      gt5_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt5_rxdata_out                  =>      gt5_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt5_rxdisperr_out               =>      gt5_rxdisperr_out,
        gt5_rxnotintable_out            =>      gt5_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt5_gthrxn_in                   =>      gt5_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt5_rxbyteisaligned_out         =>      gt5_rxbyteisaligned_out,
        gt5_rxmcommaalignen_in          =>      gt5_rxmcommaalignen_in,
        gt5_rxpcommaalignen_in          =>      gt5_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt5_rxdfeagchold_in             =>      gt5_rxdfeagchold_i,
        gt5_rxdfelfhold_in              =>      gt5_rxdfelfhold_i,
        gt5_rxmonitorout_out            =>      gt5_rxmonitorout_out,
        gt5_rxmonitorsel_in             =>      gt5_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt5_rxoutclk_out                =>      gt5_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt5_gtrxreset_in                =>      gt5_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt5_rxpolarity_in               =>      gt5_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt5_rxcharisk_out               =>      gt5_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt5_gthrxp_in                   =>      gt5_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt5_rxresetdone_out             =>      gt5_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt5_gttxreset_in                =>      gt5_gttxreset_i,
        gt5_txuserrdy_in                =>      gt5_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt5_txusrclk_in                 =>      gt5_txusrclk_in,
        gt5_txusrclk2_in                =>      gt5_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt5_txdata_in                   =>      gt5_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt5_gthtxn_out                  =>      gt5_gthtxn_out,
        gt5_gthtxp_out                  =>      gt5_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt5_txoutclk_out                =>      gt5_txoutclk_i,
        gt5_txoutclkfabric_out          =>      gt5_txoutclkfabric_out,
        gt5_txoutclkpcs_out             =>      gt5_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt5_txresetdone_out             =>      gt5_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt5_txpolarity_in               =>      gt5_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt5_txcharisk_in                =>      gt5_txcharisk_in,


        GT6_RXPMARESETDONE_OUT          =>      gt6_rxpmaresetdone_i,
        GT6_TXPMARESETDONE_OUT          =>      gt6_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT6  (X1Y14)

        --------------------------------- CPLL Ports -------------------------------
        gt6_cpllfbclklost_out           =>      gt6_cpllfbclklost_out,
        gt6_cplllock_out                =>      gt6_cplllock_i,
        gt6_cplllockdetclk_in           =>      gt6_cplllockdetclk_in,
        gt6_cpllrefclklost_out          =>      gt6_cpllrefclklost_i,
        gt6_cpllreset_in                =>      gt6_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt6_gtrefclk0_in                =>      gt6_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt6_drpaddr_in                  =>      gt6_drpaddr_in,
        gt6_drpclk_in                   =>      gt6_drpclk_in,
        gt6_drpdi_in                    =>      gt6_drpdi_in,
        gt6_drpdo_out                   =>      gt6_drpdo_out,
        gt6_drpen_in                    =>      gt6_drpen_in,
        gt6_drprdy_out                  =>      gt6_drprdy_out,
        gt6_drpwe_in                    =>      gt6_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt6_eyescanreset_in             =>      gt6_eyescanreset_in,
        gt6_rxuserrdy_in                =>      gt6_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt6_eyescandataerror_out        =>      gt6_eyescandataerror_out,
        gt6_eyescantrigger_in           =>      gt6_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt6_dmonitorout_out             =>      gt6_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt6_rxusrclk_in                 =>      gt6_rxusrclk_in,
        gt6_rxusrclk2_in                =>      gt6_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt6_rxdata_out                  =>      gt6_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt6_rxdisperr_out               =>      gt6_rxdisperr_out,
        gt6_rxnotintable_out            =>      gt6_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt6_gthrxn_in                   =>      gt6_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt6_rxbyteisaligned_out         =>      gt6_rxbyteisaligned_out,
        gt6_rxmcommaalignen_in          =>      gt6_rxmcommaalignen_in,
        gt6_rxpcommaalignen_in          =>      gt6_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt6_rxdfeagchold_in             =>      gt6_rxdfeagchold_i,
        gt6_rxdfelfhold_in              =>      gt6_rxdfelfhold_i,
        gt6_rxmonitorout_out            =>      gt6_rxmonitorout_out,
        gt6_rxmonitorsel_in             =>      gt6_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt6_rxoutclk_out                =>      gt6_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt6_gtrxreset_in                =>      gt6_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt6_rxpolarity_in               =>      gt6_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt6_rxcharisk_out               =>      gt6_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt6_gthrxp_in                   =>      gt6_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt6_rxresetdone_out             =>      gt6_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt6_gttxreset_in                =>      gt6_gttxreset_i,
        gt6_txuserrdy_in                =>      gt6_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt6_txusrclk_in                 =>      gt6_txusrclk_in,
        gt6_txusrclk2_in                =>      gt6_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt6_txdata_in                   =>      gt6_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt6_gthtxn_out                  =>      gt6_gthtxn_out,
        gt6_gthtxp_out                  =>      gt6_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt6_txoutclk_out                =>      gt6_txoutclk_i,
        gt6_txoutclkfabric_out          =>      gt6_txoutclkfabric_out,
        gt6_txoutclkpcs_out             =>      gt6_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt6_txresetdone_out             =>      gt6_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt6_txpolarity_in               =>      gt6_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt6_txcharisk_in                =>      gt6_txcharisk_in,


        GT7_RXPMARESETDONE_OUT          =>      gt7_rxpmaresetdone_i,
        GT7_TXPMARESETDONE_OUT          =>      gt7_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT7  (X1Y15)

        --------------------------------- CPLL Ports -------------------------------
        gt7_cpllfbclklost_out           =>      gt7_cpllfbclklost_out,
        gt7_cplllock_out                =>      gt7_cplllock_i,
        gt7_cplllockdetclk_in           =>      gt7_cplllockdetclk_in,
        gt7_cpllrefclklost_out          =>      gt7_cpllrefclklost_i,
        gt7_cpllreset_in                =>      gt7_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt7_gtrefclk0_in                =>      gt7_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt7_drpaddr_in                  =>      gt7_drpaddr_in,
        gt7_drpclk_in                   =>      gt7_drpclk_in,
        gt7_drpdi_in                    =>      gt7_drpdi_in,
        gt7_drpdo_out                   =>      gt7_drpdo_out,
        gt7_drpen_in                    =>      gt7_drpen_in,
        gt7_drprdy_out                  =>      gt7_drprdy_out,
        gt7_drpwe_in                    =>      gt7_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt7_eyescanreset_in             =>      gt7_eyescanreset_in,
        gt7_rxuserrdy_in                =>      gt7_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt7_eyescandataerror_out        =>      gt7_eyescandataerror_out,
        gt7_eyescantrigger_in           =>      gt7_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt7_dmonitorout_out             =>      gt7_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt7_rxusrclk_in                 =>      gt7_rxusrclk_in,
        gt7_rxusrclk2_in                =>      gt7_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt7_rxdata_out                  =>      gt7_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt7_rxdisperr_out               =>      gt7_rxdisperr_out,
        gt7_rxnotintable_out            =>      gt7_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt7_gthrxn_in                   =>      gt7_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt7_rxbyteisaligned_out         =>      gt7_rxbyteisaligned_out,
        gt7_rxmcommaalignen_in          =>      gt7_rxmcommaalignen_in,
        gt7_rxpcommaalignen_in          =>      gt7_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt7_rxdfeagchold_in             =>      gt7_rxdfeagchold_i,
        gt7_rxdfelfhold_in              =>      gt7_rxdfelfhold_i,
        gt7_rxmonitorout_out            =>      gt7_rxmonitorout_out,
        gt7_rxmonitorsel_in             =>      gt7_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt7_rxoutclk_out                =>      gt7_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt7_gtrxreset_in                =>      gt7_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt7_rxpolarity_in               =>      gt7_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt7_rxcharisk_out               =>      gt7_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt7_gthrxp_in                   =>      gt7_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt7_rxresetdone_out             =>      gt7_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt7_gttxreset_in                =>      gt7_gttxreset_i,
        gt7_txuserrdy_in                =>      gt7_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt7_txusrclk_in                 =>      gt7_txusrclk_in,
        gt7_txusrclk2_in                =>      gt7_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt7_txdata_in                   =>      gt7_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt7_gthtxn_out                  =>      gt7_gthtxn_out,
        gt7_gthtxp_out                  =>      gt7_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt7_txoutclk_out                =>      gt7_txoutclk_i,
        gt7_txoutclkfabric_out          =>      gt7_txoutclkfabric_out,
        gt7_txoutclkpcs_out             =>      gt7_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt7_txresetdone_out             =>      gt7_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt7_txpolarity_in               =>      gt7_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt7_txcharisk_in                =>      gt7_txcharisk_in,


        GT8_RXPMARESETDONE_OUT          =>      gt8_rxpmaresetdone_i,
        GT8_TXPMARESETDONE_OUT          =>      gt8_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT8  (X1Y16)

        --------------------------------- CPLL Ports -------------------------------
        gt8_cpllfbclklost_out           =>      gt8_cpllfbclklost_out,
        gt8_cplllock_out                =>      gt8_cplllock_i,
        gt8_cplllockdetclk_in           =>      gt8_cplllockdetclk_in,
        gt8_cpllrefclklost_out          =>      gt8_cpllrefclklost_i,
        gt8_cpllreset_in                =>      gt8_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt8_gtrefclk0_in                =>      gt8_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt8_drpaddr_in                  =>      gt8_drpaddr_in,
        gt8_drpclk_in                   =>      gt8_drpclk_in,
        gt8_drpdi_in                    =>      gt8_drpdi_in,
        gt8_drpdo_out                   =>      gt8_drpdo_out,
        gt8_drpen_in                    =>      gt8_drpen_in,
        gt8_drprdy_out                  =>      gt8_drprdy_out,
        gt8_drpwe_in                    =>      gt8_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt8_eyescanreset_in             =>      gt8_eyescanreset_in,
        gt8_rxuserrdy_in                =>      gt8_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt8_eyescandataerror_out        =>      gt8_eyescandataerror_out,
        gt8_eyescantrigger_in           =>      gt8_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt8_dmonitorout_out             =>      gt8_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt8_rxusrclk_in                 =>      gt8_rxusrclk_in,
        gt8_rxusrclk2_in                =>      gt8_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt8_rxdata_out                  =>      gt8_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt8_rxdisperr_out               =>      gt8_rxdisperr_out,
        gt8_rxnotintable_out            =>      gt8_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt8_gthrxn_in                   =>      gt8_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt8_rxbyteisaligned_out         =>      gt8_rxbyteisaligned_out,
        gt8_rxmcommaalignen_in          =>      gt8_rxmcommaalignen_in,
        gt8_rxpcommaalignen_in          =>      gt8_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt8_rxdfeagchold_in             =>      gt8_rxdfeagchold_i,
        gt8_rxdfelfhold_in              =>      gt8_rxdfelfhold_i,
        gt8_rxmonitorout_out            =>      gt8_rxmonitorout_out,
        gt8_rxmonitorsel_in             =>      gt8_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt8_rxoutclk_out                =>      gt8_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt8_gtrxreset_in                =>      gt8_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt8_rxpolarity_in               =>      gt8_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt8_rxcharisk_out               =>      gt8_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt8_gthrxp_in                   =>      gt8_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt8_rxresetdone_out             =>      gt8_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt8_gttxreset_in                =>      gt8_gttxreset_i,
        gt8_txuserrdy_in                =>      gt8_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt8_txusrclk_in                 =>      gt8_txusrclk_in,
        gt8_txusrclk2_in                =>      gt8_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt8_txdata_in                   =>      gt8_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt8_gthtxn_out                  =>      gt8_gthtxn_out,
        gt8_gthtxp_out                  =>      gt8_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt8_txoutclk_out                =>      gt8_txoutclk_i,
        gt8_txoutclkfabric_out          =>      gt8_txoutclkfabric_out,
        gt8_txoutclkpcs_out             =>      gt8_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt8_txresetdone_out             =>      gt8_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt8_txpolarity_in               =>      gt8_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt8_txcharisk_in                =>      gt8_txcharisk_in,


        GT9_RXPMARESETDONE_OUT          =>      gt9_rxpmaresetdone_i,
        GT9_TXPMARESETDONE_OUT          =>      gt9_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT9  (X1Y17)

        --------------------------------- CPLL Ports -------------------------------
        gt9_cpllfbclklost_out           =>      gt9_cpllfbclklost_out,
        gt9_cplllock_out                =>      gt9_cplllock_i,
        gt9_cplllockdetclk_in           =>      gt9_cplllockdetclk_in,
        gt9_cpllrefclklost_out          =>      gt9_cpllrefclklost_i,
        gt9_cpllreset_in                =>      gt9_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt9_gtrefclk0_in                =>      gt9_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt9_drpaddr_in                  =>      gt9_drpaddr_in,
        gt9_drpclk_in                   =>      gt9_drpclk_in,
        gt9_drpdi_in                    =>      gt9_drpdi_in,
        gt9_drpdo_out                   =>      gt9_drpdo_out,
        gt9_drpen_in                    =>      gt9_drpen_in,
        gt9_drprdy_out                  =>      gt9_drprdy_out,
        gt9_drpwe_in                    =>      gt9_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt9_eyescanreset_in             =>      gt9_eyescanreset_in,
        gt9_rxuserrdy_in                =>      gt9_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt9_eyescandataerror_out        =>      gt9_eyescandataerror_out,
        gt9_eyescantrigger_in           =>      gt9_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt9_dmonitorout_out             =>      gt9_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt9_rxusrclk_in                 =>      gt9_rxusrclk_in,
        gt9_rxusrclk2_in                =>      gt9_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt9_rxdata_out                  =>      gt9_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt9_rxdisperr_out               =>      gt9_rxdisperr_out,
        gt9_rxnotintable_out            =>      gt9_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt9_gthrxn_in                   =>      gt9_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt9_rxbyteisaligned_out         =>      gt9_rxbyteisaligned_out,
        gt9_rxmcommaalignen_in          =>      gt9_rxmcommaalignen_in,
        gt9_rxpcommaalignen_in          =>      gt9_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt9_rxdfeagchold_in             =>      gt9_rxdfeagchold_i,
        gt9_rxdfelfhold_in              =>      gt9_rxdfelfhold_i,
        gt9_rxmonitorout_out            =>      gt9_rxmonitorout_out,
        gt9_rxmonitorsel_in             =>      gt9_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt9_rxoutclk_out                =>      gt9_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt9_gtrxreset_in                =>      gt9_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt9_rxpolarity_in               =>      gt9_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt9_rxcharisk_out               =>      gt9_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt9_gthrxp_in                   =>      gt9_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt9_rxresetdone_out             =>      gt9_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt9_gttxreset_in                =>      gt9_gttxreset_i,
        gt9_txuserrdy_in                =>      gt9_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt9_txusrclk_in                 =>      gt9_txusrclk_in,
        gt9_txusrclk2_in                =>      gt9_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt9_txdata_in                   =>      gt9_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt9_gthtxn_out                  =>      gt9_gthtxn_out,
        gt9_gthtxp_out                  =>      gt9_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt9_txoutclk_out                =>      gt9_txoutclk_i,
        gt9_txoutclkfabric_out          =>      gt9_txoutclkfabric_out,
        gt9_txoutclkpcs_out             =>      gt9_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt9_txresetdone_out             =>      gt9_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt9_txpolarity_in               =>      gt9_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt9_txcharisk_in                =>      gt9_txcharisk_in,


        GT10_RXPMARESETDONE_OUT         =>      gt10_rxpmaresetdone_i,
        GT10_TXPMARESETDONE_OUT         =>      gt10_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT10  (X1Y18)

        --------------------------------- CPLL Ports -------------------------------
        gt10_cpllfbclklost_out          =>      gt10_cpllfbclklost_out,
        gt10_cplllock_out               =>      gt10_cplllock_i,
        gt10_cplllockdetclk_in          =>      gt10_cplllockdetclk_in,
        gt10_cpllrefclklost_out         =>      gt10_cpllrefclklost_i,
        gt10_cpllreset_in               =>      gt10_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt10_gtrefclk0_in               =>      gt10_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt10_drpaddr_in                 =>      gt10_drpaddr_in,
        gt10_drpclk_in                  =>      gt10_drpclk_in,
        gt10_drpdi_in                   =>      gt10_drpdi_in,
        gt10_drpdo_out                  =>      gt10_drpdo_out,
        gt10_drpen_in                   =>      gt10_drpen_in,
        gt10_drprdy_out                 =>      gt10_drprdy_out,
        gt10_drpwe_in                   =>      gt10_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt10_eyescanreset_in            =>      gt10_eyescanreset_in,
        gt10_rxuserrdy_in               =>      gt10_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt10_eyescandataerror_out       =>      gt10_eyescandataerror_out,
        gt10_eyescantrigger_in          =>      gt10_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt10_dmonitorout_out            =>      gt10_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt10_rxusrclk_in                =>      gt10_rxusrclk_in,
        gt10_rxusrclk2_in               =>      gt10_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt10_rxdata_out                 =>      gt10_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt10_rxdisperr_out              =>      gt10_rxdisperr_out,
        gt10_rxnotintable_out           =>      gt10_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt10_gthrxn_in                  =>      gt10_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt10_rxbyteisaligned_out        =>      gt10_rxbyteisaligned_out,
        gt10_rxmcommaalignen_in         =>      gt10_rxmcommaalignen_in,
        gt10_rxpcommaalignen_in         =>      gt10_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt10_rxdfeagchold_in            =>      gt10_rxdfeagchold_i,
        gt10_rxdfelfhold_in             =>      gt10_rxdfelfhold_i,
        gt10_rxmonitorout_out           =>      gt10_rxmonitorout_out,
        gt10_rxmonitorsel_in            =>      gt10_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt10_rxoutclk_out               =>      gt10_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt10_gtrxreset_in               =>      gt10_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt10_rxpolarity_in              =>      gt10_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt10_rxcharisk_out              =>      gt10_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt10_gthrxp_in                  =>      gt10_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt10_rxresetdone_out            =>      gt10_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt10_gttxreset_in               =>      gt10_gttxreset_i,
        gt10_txuserrdy_in               =>      gt10_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt10_txusrclk_in                =>      gt10_txusrclk_in,
        gt10_txusrclk2_in               =>      gt10_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt10_txdata_in                  =>      gt10_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt10_gthtxn_out                 =>      gt10_gthtxn_out,
        gt10_gthtxp_out                 =>      gt10_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt10_txoutclk_out               =>      gt10_txoutclk_i,
        gt10_txoutclkfabric_out         =>      gt10_txoutclkfabric_out,
        gt10_txoutclkpcs_out            =>      gt10_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt10_txresetdone_out            =>      gt10_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt10_txpolarity_in              =>      gt10_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt10_txcharisk_in               =>      gt10_txcharisk_in,


        GT11_RXPMARESETDONE_OUT         =>      gt11_rxpmaresetdone_i,
        GT11_TXPMARESETDONE_OUT         =>      gt11_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT11  (X1Y19)

        --------------------------------- CPLL Ports -------------------------------
        gt11_cpllfbclklost_out          =>      gt11_cpllfbclklost_out,
        gt11_cplllock_out               =>      gt11_cplllock_i,
        gt11_cplllockdetclk_in          =>      gt11_cplllockdetclk_in,
        gt11_cpllrefclklost_out         =>      gt11_cpllrefclklost_i,
        gt11_cpllreset_in               =>      gt11_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt11_gtrefclk0_in               =>      gt11_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt11_drpaddr_in                 =>      gt11_drpaddr_in,
        gt11_drpclk_in                  =>      gt11_drpclk_in,
        gt11_drpdi_in                   =>      gt11_drpdi_in,
        gt11_drpdo_out                  =>      gt11_drpdo_out,
        gt11_drpen_in                   =>      gt11_drpen_in,
        gt11_drprdy_out                 =>      gt11_drprdy_out,
        gt11_drpwe_in                   =>      gt11_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt11_eyescanreset_in            =>      gt11_eyescanreset_in,
        gt11_rxuserrdy_in               =>      gt11_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt11_eyescandataerror_out       =>      gt11_eyescandataerror_out,
        gt11_eyescantrigger_in          =>      gt11_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt11_dmonitorout_out            =>      gt11_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt11_rxusrclk_in                =>      gt11_rxusrclk_in,
        gt11_rxusrclk2_in               =>      gt11_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt11_rxdata_out                 =>      gt11_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt11_rxdisperr_out              =>      gt11_rxdisperr_out,
        gt11_rxnotintable_out           =>      gt11_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt11_gthrxn_in                  =>      gt11_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt11_rxbyteisaligned_out        =>      gt11_rxbyteisaligned_out,
        gt11_rxmcommaalignen_in         =>      gt11_rxmcommaalignen_in,
        gt11_rxpcommaalignen_in         =>      gt11_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt11_rxdfeagchold_in            =>      gt11_rxdfeagchold_i,
        gt11_rxdfelfhold_in             =>      gt11_rxdfelfhold_i,
        gt11_rxmonitorout_out           =>      gt11_rxmonitorout_out,
        gt11_rxmonitorsel_in            =>      gt11_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt11_rxoutclk_out               =>      gt11_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt11_gtrxreset_in               =>      gt11_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt11_rxpolarity_in              =>      gt11_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt11_rxcharisk_out              =>      gt11_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt11_gthrxp_in                  =>      gt11_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt11_rxresetdone_out            =>      gt11_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt11_gttxreset_in               =>      gt11_gttxreset_i,
        gt11_txuserrdy_in               =>      gt11_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt11_txusrclk_in                =>      gt11_txusrclk_in,
        gt11_txusrclk2_in               =>      gt11_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt11_txdata_in                  =>      gt11_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt11_gthtxn_out                 =>      gt11_gthtxn_out,
        gt11_gthtxp_out                 =>      gt11_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt11_txoutclk_out               =>      gt11_txoutclk_i,
        gt11_txoutclkfabric_out         =>      gt11_txoutclkfabric_out,
        gt11_txoutclkpcs_out            =>      gt11_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt11_txresetdone_out            =>      gt11_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt11_txpolarity_in              =>      gt11_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt11_txcharisk_in               =>      gt11_txcharisk_in,


        GT12_RXPMARESETDONE_OUT         =>      gt12_rxpmaresetdone_i,
        GT12_TXPMARESETDONE_OUT         =>      gt12_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT12  (X1Y20)

        --------------------------------- CPLL Ports -------------------------------
        gt12_cpllfbclklost_out          =>      gt12_cpllfbclklost_out,
        gt12_cplllock_out               =>      gt12_cplllock_i,
        gt12_cplllockdetclk_in          =>      gt12_cplllockdetclk_in,
        gt12_cpllrefclklost_out         =>      gt12_cpllrefclklost_i,
        gt12_cpllreset_in               =>      gt12_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt12_gtrefclk0_in               =>      gt12_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt12_drpaddr_in                 =>      gt12_drpaddr_in,
        gt12_drpclk_in                  =>      gt12_drpclk_in,
        gt12_drpdi_in                   =>      gt12_drpdi_in,
        gt12_drpdo_out                  =>      gt12_drpdo_out,
        gt12_drpen_in                   =>      gt12_drpen_in,
        gt12_drprdy_out                 =>      gt12_drprdy_out,
        gt12_drpwe_in                   =>      gt12_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt12_eyescanreset_in            =>      gt12_eyescanreset_in,
        gt12_rxuserrdy_in               =>      gt12_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt12_eyescandataerror_out       =>      gt12_eyescandataerror_out,
        gt12_eyescantrigger_in          =>      gt12_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt12_dmonitorout_out            =>      gt12_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt12_rxusrclk_in                =>      gt12_rxusrclk_in,
        gt12_rxusrclk2_in               =>      gt12_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt12_rxdata_out                 =>      gt12_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt12_rxdisperr_out              =>      gt12_rxdisperr_out,
        gt12_rxnotintable_out           =>      gt12_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt12_gthrxn_in                  =>      gt12_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt12_rxbyteisaligned_out        =>      gt12_rxbyteisaligned_out,
        gt12_rxmcommaalignen_in         =>      gt12_rxmcommaalignen_in,
        gt12_rxpcommaalignen_in         =>      gt12_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt12_rxdfeagchold_in            =>      gt12_rxdfeagchold_i,
        gt12_rxdfelfhold_in             =>      gt12_rxdfelfhold_i,
        gt12_rxmonitorout_out           =>      gt12_rxmonitorout_out,
        gt12_rxmonitorsel_in            =>      gt12_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt12_rxoutclk_out               =>      gt12_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt12_gtrxreset_in               =>      gt12_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt12_rxpolarity_in              =>      gt12_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt12_rxcharisk_out              =>      gt12_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt12_gthrxp_in                  =>      gt12_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt12_rxresetdone_out            =>      gt12_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt12_gttxreset_in               =>      gt12_gttxreset_i,
        gt12_txuserrdy_in               =>      gt12_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt12_txusrclk_in                =>      gt12_txusrclk_in,
        gt12_txusrclk2_in               =>      gt12_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt12_txdata_in                  =>      gt12_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt12_gthtxn_out                 =>      gt12_gthtxn_out,
        gt12_gthtxp_out                 =>      gt12_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt12_txoutclk_out               =>      gt12_txoutclk_i,
        gt12_txoutclkfabric_out         =>      gt12_txoutclkfabric_out,
        gt12_txoutclkpcs_out            =>      gt12_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt12_txresetdone_out            =>      gt12_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt12_txpolarity_in              =>      gt12_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt12_txcharisk_in               =>      gt12_txcharisk_in,


        GT13_RXPMARESETDONE_OUT         =>      gt13_rxpmaresetdone_i,
        GT13_TXPMARESETDONE_OUT         =>      gt13_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT13  (X1Y21)

        --------------------------------- CPLL Ports -------------------------------
        gt13_cpllfbclklost_out          =>      gt13_cpllfbclklost_out,
        gt13_cplllock_out               =>      gt13_cplllock_i,
        gt13_cplllockdetclk_in          =>      gt13_cplllockdetclk_in,
        gt13_cpllrefclklost_out         =>      gt13_cpllrefclklost_i,
        gt13_cpllreset_in               =>      gt13_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt13_gtrefclk0_in               =>      gt13_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt13_drpaddr_in                 =>      gt13_drpaddr_in,
        gt13_drpclk_in                  =>      gt13_drpclk_in,
        gt13_drpdi_in                   =>      gt13_drpdi_in,
        gt13_drpdo_out                  =>      gt13_drpdo_out,
        gt13_drpen_in                   =>      gt13_drpen_in,
        gt13_drprdy_out                 =>      gt13_drprdy_out,
        gt13_drpwe_in                   =>      gt13_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt13_eyescanreset_in            =>      gt13_eyescanreset_in,
        gt13_rxuserrdy_in               =>      gt13_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt13_eyescandataerror_out       =>      gt13_eyescandataerror_out,
        gt13_eyescantrigger_in          =>      gt13_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt13_dmonitorout_out            =>      gt13_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt13_rxusrclk_in                =>      gt13_rxusrclk_in,
        gt13_rxusrclk2_in               =>      gt13_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt13_rxdata_out                 =>      gt13_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt13_rxdisperr_out              =>      gt13_rxdisperr_out,
        gt13_rxnotintable_out           =>      gt13_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt13_gthrxn_in                  =>      gt13_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt13_rxbyteisaligned_out        =>      gt13_rxbyteisaligned_out,
        gt13_rxmcommaalignen_in         =>      gt13_rxmcommaalignen_in,
        gt13_rxpcommaalignen_in         =>      gt13_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt13_rxdfeagchold_in            =>      gt13_rxdfeagchold_i,
        gt13_rxdfelfhold_in             =>      gt13_rxdfelfhold_i,
        gt13_rxmonitorout_out           =>      gt13_rxmonitorout_out,
        gt13_rxmonitorsel_in            =>      gt13_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt13_rxoutclk_out               =>      gt13_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt13_gtrxreset_in               =>      gt13_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt13_rxpolarity_in              =>      gt13_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt13_rxcharisk_out              =>      gt13_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt13_gthrxp_in                  =>      gt13_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt13_rxresetdone_out            =>      gt13_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt13_gttxreset_in               =>      gt13_gttxreset_i,
        gt13_txuserrdy_in               =>      gt13_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt13_txusrclk_in                =>      gt13_txusrclk_in,
        gt13_txusrclk2_in               =>      gt13_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt13_txdata_in                  =>      gt13_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt13_gthtxn_out                 =>      gt13_gthtxn_out,
        gt13_gthtxp_out                 =>      gt13_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt13_txoutclk_out               =>      gt13_txoutclk_i,
        gt13_txoutclkfabric_out         =>      gt13_txoutclkfabric_out,
        gt13_txoutclkpcs_out            =>      gt13_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt13_txresetdone_out            =>      gt13_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt13_txpolarity_in              =>      gt13_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt13_txcharisk_in               =>      gt13_txcharisk_in,


        GT14_RXPMARESETDONE_OUT         =>      gt14_rxpmaresetdone_i,
        GT14_TXPMARESETDONE_OUT         =>      gt14_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT14  (X1Y22)

        --------------------------------- CPLL Ports -------------------------------
        gt14_cpllfbclklost_out          =>      gt14_cpllfbclklost_out,
        gt14_cplllock_out               =>      gt14_cplllock_i,
        gt14_cplllockdetclk_in          =>      gt14_cplllockdetclk_in,
        gt14_cpllrefclklost_out         =>      gt14_cpllrefclklost_i,
        gt14_cpllreset_in               =>      gt14_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt14_gtrefclk0_in               =>      gt14_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt14_drpaddr_in                 =>      gt14_drpaddr_in,
        gt14_drpclk_in                  =>      gt14_drpclk_in,
        gt14_drpdi_in                   =>      gt14_drpdi_in,
        gt14_drpdo_out                  =>      gt14_drpdo_out,
        gt14_drpen_in                   =>      gt14_drpen_in,
        gt14_drprdy_out                 =>      gt14_drprdy_out,
        gt14_drpwe_in                   =>      gt14_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt14_eyescanreset_in            =>      gt14_eyescanreset_in,
        gt14_rxuserrdy_in               =>      gt14_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt14_eyescandataerror_out       =>      gt14_eyescandataerror_out,
        gt14_eyescantrigger_in          =>      gt14_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt14_dmonitorout_out            =>      gt14_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt14_rxusrclk_in                =>      gt14_rxusrclk_in,
        gt14_rxusrclk2_in               =>      gt14_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt14_rxdata_out                 =>      gt14_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt14_rxdisperr_out              =>      gt14_rxdisperr_out,
        gt14_rxnotintable_out           =>      gt14_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt14_gthrxn_in                  =>      gt14_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt14_rxbyteisaligned_out        =>      gt14_rxbyteisaligned_out,
        gt14_rxmcommaalignen_in         =>      gt14_rxmcommaalignen_in,
        gt14_rxpcommaalignen_in         =>      gt14_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt14_rxdfeagchold_in            =>      gt14_rxdfeagchold_i,
        gt14_rxdfelfhold_in             =>      gt14_rxdfelfhold_i,
        gt14_rxmonitorout_out           =>      gt14_rxmonitorout_out,
        gt14_rxmonitorsel_in            =>      gt14_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt14_rxoutclk_out               =>      gt14_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt14_gtrxreset_in               =>      gt14_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt14_rxpolarity_in              =>      gt14_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt14_rxcharisk_out              =>      gt14_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt14_gthrxp_in                  =>      gt14_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt14_rxresetdone_out            =>      gt14_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt14_gttxreset_in               =>      gt14_gttxreset_i,
        gt14_txuserrdy_in               =>      gt14_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt14_txusrclk_in                =>      gt14_txusrclk_in,
        gt14_txusrclk2_in               =>      gt14_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt14_txdata_in                  =>      gt14_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt14_gthtxn_out                 =>      gt14_gthtxn_out,
        gt14_gthtxp_out                 =>      gt14_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt14_txoutclk_out               =>      gt14_txoutclk_i,
        gt14_txoutclkfabric_out         =>      gt14_txoutclkfabric_out,
        gt14_txoutclkpcs_out            =>      gt14_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt14_txresetdone_out            =>      gt14_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt14_txpolarity_in              =>      gt14_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt14_txcharisk_in               =>      gt14_txcharisk_in,


        GT15_RXPMARESETDONE_OUT         =>      gt15_rxpmaresetdone_i,
        GT15_TXPMARESETDONE_OUT         =>      gt15_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT15  (X1Y23)

        --------------------------------- CPLL Ports -------------------------------
        gt15_cpllfbclklost_out          =>      gt15_cpllfbclklost_out,
        gt15_cplllock_out               =>      gt15_cplllock_i,
        gt15_cplllockdetclk_in          =>      gt15_cplllockdetclk_in,
        gt15_cpllrefclklost_out         =>      gt15_cpllrefclklost_i,
        gt15_cpllreset_in               =>      gt15_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt15_gtrefclk0_in               =>      gt15_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt15_drpaddr_in                 =>      gt15_drpaddr_in,
        gt15_drpclk_in                  =>      gt15_drpclk_in,
        gt15_drpdi_in                   =>      gt15_drpdi_in,
        gt15_drpdo_out                  =>      gt15_drpdo_out,
        gt15_drpen_in                   =>      gt15_drpen_in,
        gt15_drprdy_out                 =>      gt15_drprdy_out,
        gt15_drpwe_in                   =>      gt15_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt15_eyescanreset_in            =>      gt15_eyescanreset_in,
        gt15_rxuserrdy_in               =>      gt15_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt15_eyescandataerror_out       =>      gt15_eyescandataerror_out,
        gt15_eyescantrigger_in          =>      gt15_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt15_dmonitorout_out            =>      gt15_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt15_rxusrclk_in                =>      gt15_rxusrclk_in,
        gt15_rxusrclk2_in               =>      gt15_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt15_rxdata_out                 =>      gt15_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt15_rxdisperr_out              =>      gt15_rxdisperr_out,
        gt15_rxnotintable_out           =>      gt15_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt15_gthrxn_in                  =>      gt15_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt15_rxbyteisaligned_out        =>      gt15_rxbyteisaligned_out,
        gt15_rxmcommaalignen_in         =>      gt15_rxmcommaalignen_in,
        gt15_rxpcommaalignen_in         =>      gt15_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt15_rxdfeagchold_in            =>      gt15_rxdfeagchold_i,
        gt15_rxdfelfhold_in             =>      gt15_rxdfelfhold_i,
        gt15_rxmonitorout_out           =>      gt15_rxmonitorout_out,
        gt15_rxmonitorsel_in            =>      gt15_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt15_rxoutclk_out               =>      gt15_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt15_gtrxreset_in               =>      gt15_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt15_rxpolarity_in              =>      gt15_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt15_rxcharisk_out              =>      gt15_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt15_gthrxp_in                  =>      gt15_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt15_rxresetdone_out            =>      gt15_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt15_gttxreset_in               =>      gt15_gttxreset_i,
        gt15_txuserrdy_in               =>      gt15_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt15_txusrclk_in                =>      gt15_txusrclk_in,
        gt15_txusrclk2_in               =>      gt15_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt15_txdata_in                  =>      gt15_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt15_gthtxn_out                 =>      gt15_gthtxn_out,
        gt15_gthtxp_out                 =>      gt15_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt15_txoutclk_out               =>      gt15_txoutclk_i,
        gt15_txoutclkfabric_out         =>      gt15_txoutclkfabric_out,
        gt15_txoutclkpcs_out            =>      gt15_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt15_txresetdone_out            =>      gt15_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt15_txpolarity_in              =>      gt15_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt15_txcharisk_in               =>      gt15_txcharisk_in,


        GT16_RXPMARESETDONE_OUT         =>      gt16_rxpmaresetdone_i,
        GT16_TXPMARESETDONE_OUT         =>      gt16_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT16  (X1Y24)

        --------------------------------- CPLL Ports -------------------------------
        gt16_cpllfbclklost_out          =>      gt16_cpllfbclklost_out,
        gt16_cplllock_out               =>      gt16_cplllock_i,
        gt16_cplllockdetclk_in          =>      gt16_cplllockdetclk_in,
        gt16_cpllrefclklost_out         =>      gt16_cpllrefclklost_i,
        gt16_cpllreset_in               =>      gt16_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt16_gtrefclk0_in               =>      gt16_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt16_drpaddr_in                 =>      gt16_drpaddr_in,
        gt16_drpclk_in                  =>      gt16_drpclk_in,
        gt16_drpdi_in                   =>      gt16_drpdi_in,
        gt16_drpdo_out                  =>      gt16_drpdo_out,
        gt16_drpen_in                   =>      gt16_drpen_in,
        gt16_drprdy_out                 =>      gt16_drprdy_out,
        gt16_drpwe_in                   =>      gt16_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt16_eyescanreset_in            =>      gt16_eyescanreset_in,
        gt16_rxuserrdy_in               =>      gt16_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt16_eyescandataerror_out       =>      gt16_eyescandataerror_out,
        gt16_eyescantrigger_in          =>      gt16_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt16_dmonitorout_out            =>      gt16_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt16_rxusrclk_in                =>      gt16_rxusrclk_in,
        gt16_rxusrclk2_in               =>      gt16_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt16_rxdata_out                 =>      gt16_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt16_rxdisperr_out              =>      gt16_rxdisperr_out,
        gt16_rxnotintable_out           =>      gt16_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt16_gthrxn_in                  =>      gt16_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt16_rxbyteisaligned_out        =>      gt16_rxbyteisaligned_out,
        gt16_rxmcommaalignen_in         =>      gt16_rxmcommaalignen_in,
        gt16_rxpcommaalignen_in         =>      gt16_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt16_rxdfeagchold_in            =>      gt16_rxdfeagchold_i,
        gt16_rxdfelfhold_in             =>      gt16_rxdfelfhold_i,
        gt16_rxmonitorout_out           =>      gt16_rxmonitorout_out,
        gt16_rxmonitorsel_in            =>      gt16_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt16_rxoutclk_out               =>      gt16_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt16_gtrxreset_in               =>      gt16_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt16_rxpolarity_in              =>      gt16_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt16_rxcharisk_out              =>      gt16_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt16_gthrxp_in                  =>      gt16_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt16_rxresetdone_out            =>      gt16_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt16_gttxreset_in               =>      gt16_gttxreset_i,
        gt16_txuserrdy_in               =>      gt16_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt16_txusrclk_in                =>      gt16_txusrclk_in,
        gt16_txusrclk2_in               =>      gt16_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt16_txdata_in                  =>      gt16_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt16_gthtxn_out                 =>      gt16_gthtxn_out,
        gt16_gthtxp_out                 =>      gt16_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt16_txoutclk_out               =>      gt16_txoutclk_i,
        gt16_txoutclkfabric_out         =>      gt16_txoutclkfabric_out,
        gt16_txoutclkpcs_out            =>      gt16_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt16_txresetdone_out            =>      gt16_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt16_txpolarity_in              =>      gt16_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt16_txcharisk_in               =>      gt16_txcharisk_in,


        GT17_RXPMARESETDONE_OUT         =>      gt17_rxpmaresetdone_i,
        GT17_TXPMARESETDONE_OUT         =>      gt17_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT17  (X1Y25)

        --------------------------------- CPLL Ports -------------------------------
        gt17_cpllfbclklost_out          =>      gt17_cpllfbclklost_out,
        gt17_cplllock_out               =>      gt17_cplllock_i,
        gt17_cplllockdetclk_in          =>      gt17_cplllockdetclk_in,
        gt17_cpllrefclklost_out         =>      gt17_cpllrefclklost_i,
        gt17_cpllreset_in               =>      gt17_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt17_gtrefclk0_in               =>      gt17_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt17_drpaddr_in                 =>      gt17_drpaddr_in,
        gt17_drpclk_in                  =>      gt17_drpclk_in,
        gt17_drpdi_in                   =>      gt17_drpdi_in,
        gt17_drpdo_out                  =>      gt17_drpdo_out,
        gt17_drpen_in                   =>      gt17_drpen_in,
        gt17_drprdy_out                 =>      gt17_drprdy_out,
        gt17_drpwe_in                   =>      gt17_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt17_eyescanreset_in            =>      gt17_eyescanreset_in,
        gt17_rxuserrdy_in               =>      gt17_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt17_eyescandataerror_out       =>      gt17_eyescandataerror_out,
        gt17_eyescantrigger_in          =>      gt17_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt17_dmonitorout_out            =>      gt17_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt17_rxusrclk_in                =>      gt17_rxusrclk_in,
        gt17_rxusrclk2_in               =>      gt17_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt17_rxdata_out                 =>      gt17_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt17_rxdisperr_out              =>      gt17_rxdisperr_out,
        gt17_rxnotintable_out           =>      gt17_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt17_gthrxn_in                  =>      gt17_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt17_rxbyteisaligned_out        =>      gt17_rxbyteisaligned_out,
        gt17_rxmcommaalignen_in         =>      gt17_rxmcommaalignen_in,
        gt17_rxpcommaalignen_in         =>      gt17_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt17_rxdfeagchold_in            =>      gt17_rxdfeagchold_i,
        gt17_rxdfelfhold_in             =>      gt17_rxdfelfhold_i,
        gt17_rxmonitorout_out           =>      gt17_rxmonitorout_out,
        gt17_rxmonitorsel_in            =>      gt17_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt17_rxoutclk_out               =>      gt17_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt17_gtrxreset_in               =>      gt17_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt17_rxpolarity_in              =>      gt17_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt17_rxcharisk_out              =>      gt17_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt17_gthrxp_in                  =>      gt17_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt17_rxresetdone_out            =>      gt17_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt17_gttxreset_in               =>      gt17_gttxreset_i,
        gt17_txuserrdy_in               =>      gt17_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt17_txusrclk_in                =>      gt17_txusrclk_in,
        gt17_txusrclk2_in               =>      gt17_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt17_txdata_in                  =>      gt17_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt17_gthtxn_out                 =>      gt17_gthtxn_out,
        gt17_gthtxp_out                 =>      gt17_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt17_txoutclk_out               =>      gt17_txoutclk_i,
        gt17_txoutclkfabric_out         =>      gt17_txoutclkfabric_out,
        gt17_txoutclkpcs_out            =>      gt17_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt17_txresetdone_out            =>      gt17_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt17_txpolarity_in              =>      gt17_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt17_txcharisk_in               =>      gt17_txcharisk_in,


        GT18_RXPMARESETDONE_OUT         =>      gt18_rxpmaresetdone_i,
        GT18_TXPMARESETDONE_OUT         =>      gt18_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT18  (X1Y26)

        --------------------------------- CPLL Ports -------------------------------
        gt18_cpllfbclklost_out          =>      gt18_cpllfbclklost_out,
        gt18_cplllock_out               =>      gt18_cplllock_i,
        gt18_cplllockdetclk_in          =>      gt18_cplllockdetclk_in,
        gt18_cpllrefclklost_out         =>      gt18_cpllrefclklost_i,
        gt18_cpllreset_in               =>      gt18_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt18_gtrefclk0_in               =>      gt18_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt18_drpaddr_in                 =>      gt18_drpaddr_in,
        gt18_drpclk_in                  =>      gt18_drpclk_in,
        gt18_drpdi_in                   =>      gt18_drpdi_in,
        gt18_drpdo_out                  =>      gt18_drpdo_out,
        gt18_drpen_in                   =>      gt18_drpen_in,
        gt18_drprdy_out                 =>      gt18_drprdy_out,
        gt18_drpwe_in                   =>      gt18_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt18_eyescanreset_in            =>      gt18_eyescanreset_in,
        gt18_rxuserrdy_in               =>      gt18_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt18_eyescandataerror_out       =>      gt18_eyescandataerror_out,
        gt18_eyescantrigger_in          =>      gt18_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt18_dmonitorout_out            =>      gt18_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt18_rxusrclk_in                =>      gt18_rxusrclk_in,
        gt18_rxusrclk2_in               =>      gt18_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt18_rxdata_out                 =>      gt18_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt18_rxdisperr_out              =>      gt18_rxdisperr_out,
        gt18_rxnotintable_out           =>      gt18_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt18_gthrxn_in                  =>      gt18_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt18_rxbyteisaligned_out        =>      gt18_rxbyteisaligned_out,
        gt18_rxmcommaalignen_in         =>      gt18_rxmcommaalignen_in,
        gt18_rxpcommaalignen_in         =>      gt18_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt18_rxdfeagchold_in            =>      gt18_rxdfeagchold_i,
        gt18_rxdfelfhold_in             =>      gt18_rxdfelfhold_i,
        gt18_rxmonitorout_out           =>      gt18_rxmonitorout_out,
        gt18_rxmonitorsel_in            =>      gt18_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt18_rxoutclk_out               =>      gt18_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt18_gtrxreset_in               =>      gt18_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt18_rxpolarity_in              =>      gt18_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt18_rxcharisk_out              =>      gt18_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt18_gthrxp_in                  =>      gt18_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt18_rxresetdone_out            =>      gt18_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt18_gttxreset_in               =>      gt18_gttxreset_i,
        gt18_txuserrdy_in               =>      gt18_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt18_txusrclk_in                =>      gt18_txusrclk_in,
        gt18_txusrclk2_in               =>      gt18_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt18_txdata_in                  =>      gt18_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt18_gthtxn_out                 =>      gt18_gthtxn_out,
        gt18_gthtxp_out                 =>      gt18_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt18_txoutclk_out               =>      gt18_txoutclk_i,
        gt18_txoutclkfabric_out         =>      gt18_txoutclkfabric_out,
        gt18_txoutclkpcs_out            =>      gt18_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt18_txresetdone_out            =>      gt18_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt18_txpolarity_in              =>      gt18_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt18_txcharisk_in               =>      gt18_txcharisk_in,


        GT19_RXPMARESETDONE_OUT         =>      gt19_rxpmaresetdone_i,
        GT19_TXPMARESETDONE_OUT         =>      gt19_txpmaresetdone_i,
        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT19  (X1Y27)

        --------------------------------- CPLL Ports -------------------------------
        gt19_cpllfbclklost_out          =>      gt19_cpllfbclklost_out,
        gt19_cplllock_out               =>      gt19_cplllock_i,
        gt19_cplllockdetclk_in          =>      gt19_cplllockdetclk_in,
        gt19_cpllrefclklost_out         =>      gt19_cpllrefclklost_i,
        gt19_cpllreset_in               =>      gt19_cpllreset_i,
        -------------------------- Channel - Clocking Ports ------------------------
        gt19_gtrefclk0_in               =>      gt19_gtrefclk0_in,
        ---------------------------- Channel - DRP Ports  --------------------------
        gt19_drpaddr_in                 =>      gt19_drpaddr_in,
        gt19_drpclk_in                  =>      gt19_drpclk_in,
        gt19_drpdi_in                   =>      gt19_drpdi_in,
        gt19_drpdo_out                  =>      gt19_drpdo_out,
        gt19_drpen_in                   =>      gt19_drpen_in,
        gt19_drprdy_out                 =>      gt19_drprdy_out,
        gt19_drpwe_in                   =>      gt19_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt19_eyescanreset_in            =>      gt19_eyescanreset_in,
        gt19_rxuserrdy_in               =>      gt19_rxuserrdy_i,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt19_eyescandataerror_out       =>      gt19_eyescandataerror_out,
        gt19_eyescantrigger_in          =>      gt19_eyescantrigger_in,
        ------------------- Receive Ports - Digital Monitor Ports ------------------
        gt19_dmonitorout_out            =>      gt19_dmonitorout_out,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt19_rxusrclk_in                =>      gt19_rxusrclk_in,
        gt19_rxusrclk2_in               =>      gt19_rxusrclk2_in,
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt19_rxdata_out                 =>      gt19_rxdata_out,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt19_rxdisperr_out              =>      gt19_rxdisperr_out,
        gt19_rxnotintable_out           =>      gt19_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt19_gthrxn_in                  =>      gt19_gthrxn_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt19_rxbyteisaligned_out        =>      gt19_rxbyteisaligned_out,
        gt19_rxmcommaalignen_in         =>      gt19_rxmcommaalignen_in,
        gt19_rxpcommaalignen_in         =>      gt19_rxpcommaalignen_in,
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt19_rxdfeagchold_in            =>      gt19_rxdfeagchold_i,
        gt19_rxdfelfhold_in             =>      gt19_rxdfelfhold_i,
        gt19_rxmonitorout_out           =>      gt19_rxmonitorout_out,
        gt19_rxmonitorsel_in            =>      gt19_rxmonitorsel_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt19_rxoutclk_out               =>      gt19_rxoutclk_i,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt19_gtrxreset_in               =>      gt19_gtrxreset_i,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt19_rxpolarity_in              =>      gt19_rxpolarity_in,
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt19_rxcharisk_out              =>      gt19_rxcharisk_out,
        ------------------------ Receive Ports -RX AFE Ports -----------------------
        gt19_gthrxp_in                  =>      gt19_gthrxp_in,
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt19_rxresetdone_out            =>      gt19_rxresetdone_i,
        --------------------- TX Initialization and Reset Ports --------------------
        gt19_gttxreset_in               =>      gt19_gttxreset_i,
        gt19_txuserrdy_in               =>      gt19_txuserrdy_i,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt19_txusrclk_in                =>      gt19_txusrclk_in,
        gt19_txusrclk2_in               =>      gt19_txusrclk2_in,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt19_txdata_in                  =>      gt19_txdata_in,
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt19_gthtxn_out                 =>      gt19_gthtxn_out,
        gt19_gthtxp_out                 =>      gt19_gthtxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt19_txoutclk_out               =>      gt19_txoutclk_i,
        gt19_txoutclkfabric_out         =>      gt19_txoutclkfabric_out,
        gt19_txoutclkpcs_out            =>      gt19_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt19_txresetdone_out            =>      gt19_txresetdone_i,
        ----------------- Transmit Ports - TX Polarity Control Ports ---------------
        gt19_txpolarity_in              =>      gt19_txpolarity_in,
        ----------- Transmit Transmit Ports - 8b10b Encoder Control Ports ----------
        gt19_txcharisk_in               =>      gt19_txcharisk_in,




    --____________________________COMMON PORTS________________________________
        gt0_qplloutclk_in               =>      gt0_qplloutclk_in,
        gt0_qplloutrefclk_in            =>      gt0_qplloutrefclk_in,

    --____________________________COMMON PORTS________________________________
        gt1_qplloutclk_in               =>      gt1_qplloutclk_in,
        gt1_qplloutrefclk_in            =>      gt1_qplloutrefclk_in,

    --____________________________COMMON PORTS________________________________
        gt2_qplloutclk_in               =>      gt2_qplloutclk_in,
        gt2_qplloutrefclk_in            =>      gt2_qplloutrefclk_in,

    --____________________________COMMON PORTS________________________________
        gt3_qplloutclk_in               =>      gt3_qplloutclk_in,
        gt3_qplloutrefclk_in            =>      gt3_qplloutrefclk_in,

    --____________________________COMMON PORTS________________________________
        gt4_qplloutclk_in               =>      gt4_qplloutclk_in,
        gt4_qplloutrefclk_in            =>      gt4_qplloutrefclk_in
    );




GT0_CPLLLOCK_OUT                             <= gt0_cplllock_i;
GT0_TXRESETDONE_OUT                          <= gt0_txresetdone_i;
GT0_RXRESETDONE_OUT                          <= gt0_rxresetdone_i;
GT0_TXOUTCLK_OUT                             <= gt0_txoutclk_i;
GT1_CPLLLOCK_OUT                             <= gt1_cplllock_i;
GT1_TXRESETDONE_OUT                          <= gt1_txresetdone_i;
GT1_RXRESETDONE_OUT                          <= gt1_rxresetdone_i;
GT1_TXOUTCLK_OUT                             <= gt1_txoutclk_i;
GT2_CPLLLOCK_OUT                             <= gt2_cplllock_i;
GT2_TXRESETDONE_OUT                          <= gt2_txresetdone_i;
GT2_RXRESETDONE_OUT                          <= gt2_rxresetdone_i;
GT2_TXOUTCLK_OUT                             <= gt2_txoutclk_i;
GT3_CPLLLOCK_OUT                             <= gt3_cplllock_i;
GT3_TXRESETDONE_OUT                          <= gt3_txresetdone_i;
GT3_RXRESETDONE_OUT                          <= gt3_rxresetdone_i;
GT3_TXOUTCLK_OUT                             <= gt3_txoutclk_i;
GT4_CPLLLOCK_OUT                             <= gt4_cplllock_i;
GT4_TXRESETDONE_OUT                          <= gt4_txresetdone_i;
GT4_RXRESETDONE_OUT                          <= gt4_rxresetdone_i;
GT4_TXOUTCLK_OUT                             <= gt4_txoutclk_i;
GT5_CPLLLOCK_OUT                             <= gt5_cplllock_i;
GT5_TXRESETDONE_OUT                          <= gt5_txresetdone_i;
GT5_RXRESETDONE_OUT                          <= gt5_rxresetdone_i;
GT5_TXOUTCLK_OUT                             <= gt5_txoutclk_i;
GT6_CPLLLOCK_OUT                             <= gt6_cplllock_i;
GT6_TXRESETDONE_OUT                          <= gt6_txresetdone_i;
GT6_RXRESETDONE_OUT                          <= gt6_rxresetdone_i;
GT6_TXOUTCLK_OUT                             <= gt6_txoutclk_i;
GT7_CPLLLOCK_OUT                             <= gt7_cplllock_i;
GT7_TXRESETDONE_OUT                          <= gt7_txresetdone_i;
GT7_RXRESETDONE_OUT                          <= gt7_rxresetdone_i;
GT7_TXOUTCLK_OUT                             <= gt7_txoutclk_i;
GT8_CPLLLOCK_OUT                             <= gt8_cplllock_i;
GT8_TXRESETDONE_OUT                          <= gt8_txresetdone_i;
GT8_RXRESETDONE_OUT                          <= gt8_rxresetdone_i;
GT8_TXOUTCLK_OUT                             <= gt8_txoutclk_i;
GT9_CPLLLOCK_OUT                             <= gt9_cplllock_i;
GT9_TXRESETDONE_OUT                          <= gt9_txresetdone_i;
GT9_RXRESETDONE_OUT                          <= gt9_rxresetdone_i;
GT9_TXOUTCLK_OUT                             <= gt9_txoutclk_i;
GT10_CPLLLOCK_OUT                            <= gt10_cplllock_i;
GT10_TXRESETDONE_OUT                         <= gt10_txresetdone_i;
GT10_RXRESETDONE_OUT                         <= gt10_rxresetdone_i;
GT10_TXOUTCLK_OUT                            <= gt10_txoutclk_i;
GT11_CPLLLOCK_OUT                            <= gt11_cplllock_i;
GT11_TXRESETDONE_OUT                         <= gt11_txresetdone_i;
GT11_RXRESETDONE_OUT                         <= gt11_rxresetdone_i;
GT11_TXOUTCLK_OUT                            <= gt11_txoutclk_i;
GT12_CPLLLOCK_OUT                            <= gt12_cplllock_i;
GT12_TXRESETDONE_OUT                         <= gt12_txresetdone_i;
GT12_RXRESETDONE_OUT                         <= gt12_rxresetdone_i;
GT12_TXOUTCLK_OUT                            <= gt12_txoutclk_i;
GT13_CPLLLOCK_OUT                            <= gt13_cplllock_i;
GT13_TXRESETDONE_OUT                         <= gt13_txresetdone_i;
GT13_RXRESETDONE_OUT                         <= gt13_rxresetdone_i;
GT13_TXOUTCLK_OUT                            <= gt13_txoutclk_i;
GT14_CPLLLOCK_OUT                            <= gt14_cplllock_i;
GT14_TXRESETDONE_OUT                         <= gt14_txresetdone_i;
GT14_RXRESETDONE_OUT                         <= gt14_rxresetdone_i;
GT14_TXOUTCLK_OUT                            <= gt14_txoutclk_i;
GT15_CPLLLOCK_OUT                            <= gt15_cplllock_i;
GT15_TXRESETDONE_OUT                         <= gt15_txresetdone_i;
GT15_RXRESETDONE_OUT                         <= gt15_rxresetdone_i;
GT15_TXOUTCLK_OUT                            <= gt15_txoutclk_i;
GT16_CPLLLOCK_OUT                            <= gt16_cplllock_i;
GT16_TXRESETDONE_OUT                         <= gt16_txresetdone_i;
GT16_RXRESETDONE_OUT                         <= gt16_rxresetdone_i;
GT16_TXOUTCLK_OUT                            <= gt16_txoutclk_i;
GT17_CPLLLOCK_OUT                            <= gt17_cplllock_i;
GT17_TXRESETDONE_OUT                         <= gt17_txresetdone_i;
GT17_RXRESETDONE_OUT                         <= gt17_rxresetdone_i;
GT17_TXOUTCLK_OUT                            <= gt17_txoutclk_i;
GT18_CPLLLOCK_OUT                            <= gt18_cplllock_i;
GT18_TXRESETDONE_OUT                         <= gt18_txresetdone_i;
GT18_RXRESETDONE_OUT                         <= gt18_rxresetdone_i;
GT18_TXOUTCLK_OUT                            <= gt18_txoutclk_i;
GT19_CPLLLOCK_OUT                            <= gt19_cplllock_i;
GT19_TXRESETDONE_OUT                         <= gt19_txresetdone_i;
GT19_RXRESETDONE_OUT                         <= gt19_rxresetdone_i;
GT19_TXOUTCLK_OUT                            <= gt19_txoutclk_i;

chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate
gt0_cpllreset_i                              <= GT0_CPLLRESET_IN or gt0_cpllreset_t;
    gt0_gttxreset_i                              <= GT0_GTTXRESET_IN or gt0_gttxreset_t;
    gt0_gtrxreset_i                              <= GT0_GTRXRESET_IN or gt0_gtrxreset_t;
    gt0_txuserrdy_i                              <= GT0_TXUSERRDY_IN or gt0_txuserrdy_t;
    gt0_rxuserrdy_i                              <= GT0_RXUSERRDY_IN or gt0_rxuserrdy_t;
gt1_cpllreset_i                              <= GT1_CPLLRESET_IN or gt1_cpllreset_t;
    gt1_gttxreset_i                              <= GT1_GTTXRESET_IN or gt1_gttxreset_t;
    gt1_gtrxreset_i                              <= GT1_GTRXRESET_IN or gt1_gtrxreset_t;
    gt1_txuserrdy_i                              <= GT1_TXUSERRDY_IN or gt1_txuserrdy_t;
    gt1_rxuserrdy_i                              <= GT1_RXUSERRDY_IN or gt1_rxuserrdy_t;
gt2_cpllreset_i                              <= GT2_CPLLRESET_IN or gt2_cpllreset_t;
    gt2_gttxreset_i                              <= GT2_GTTXRESET_IN or gt2_gttxreset_t;
    gt2_gtrxreset_i                              <= GT2_GTRXRESET_IN or gt2_gtrxreset_t;
    gt2_txuserrdy_i                              <= GT2_TXUSERRDY_IN or gt2_txuserrdy_t;
    gt2_rxuserrdy_i                              <= GT2_RXUSERRDY_IN or gt2_rxuserrdy_t;
gt3_cpllreset_i                              <= GT3_CPLLRESET_IN or gt3_cpllreset_t;
    gt3_gttxreset_i                              <= GT3_GTTXRESET_IN or gt3_gttxreset_t;
    gt3_gtrxreset_i                              <= GT3_GTRXRESET_IN or gt3_gtrxreset_t;
    gt3_txuserrdy_i                              <= GT3_TXUSERRDY_IN or gt3_txuserrdy_t;
    gt3_rxuserrdy_i                              <= GT3_RXUSERRDY_IN or gt3_rxuserrdy_t;
gt4_cpllreset_i                              <= GT4_CPLLRESET_IN or gt4_cpllreset_t;
    gt4_gttxreset_i                              <= GT4_GTTXRESET_IN or gt4_gttxreset_t;
    gt4_gtrxreset_i                              <= GT4_GTRXRESET_IN or gt4_gtrxreset_t;
    gt4_txuserrdy_i                              <= GT4_TXUSERRDY_IN or gt4_txuserrdy_t;
    gt4_rxuserrdy_i                              <= GT4_RXUSERRDY_IN or gt4_rxuserrdy_t;
gt5_cpllreset_i                              <= GT5_CPLLRESET_IN or gt5_cpllreset_t;
    gt5_gttxreset_i                              <= GT5_GTTXRESET_IN or gt5_gttxreset_t;
    gt5_gtrxreset_i                              <= GT5_GTRXRESET_IN or gt5_gtrxreset_t;
    gt5_txuserrdy_i                              <= GT5_TXUSERRDY_IN or gt5_txuserrdy_t;
    gt5_rxuserrdy_i                              <= GT5_RXUSERRDY_IN or gt5_rxuserrdy_t;
gt6_cpllreset_i                              <= GT6_CPLLRESET_IN or gt6_cpllreset_t;
    gt6_gttxreset_i                              <= GT6_GTTXRESET_IN or gt6_gttxreset_t;
    gt6_gtrxreset_i                              <= GT6_GTRXRESET_IN or gt6_gtrxreset_t;
    gt6_txuserrdy_i                              <= GT6_TXUSERRDY_IN or gt6_txuserrdy_t;
    gt6_rxuserrdy_i                              <= GT6_RXUSERRDY_IN or gt6_rxuserrdy_t;
gt7_cpllreset_i                              <= GT7_CPLLRESET_IN or gt7_cpllreset_t;
    gt7_gttxreset_i                              <= GT7_GTTXRESET_IN or gt7_gttxreset_t;
    gt7_gtrxreset_i                              <= GT7_GTRXRESET_IN or gt7_gtrxreset_t;
    gt7_txuserrdy_i                              <= GT7_TXUSERRDY_IN or gt7_txuserrdy_t;
    gt7_rxuserrdy_i                              <= GT7_RXUSERRDY_IN or gt7_rxuserrdy_t;
gt8_cpllreset_i                              <= GT8_CPLLRESET_IN or gt8_cpllreset_t;
    gt8_gttxreset_i                              <= GT8_GTTXRESET_IN or gt8_gttxreset_t;
    gt8_gtrxreset_i                              <= GT8_GTRXRESET_IN or gt8_gtrxreset_t;
    gt8_txuserrdy_i                              <= GT8_TXUSERRDY_IN or gt8_txuserrdy_t;
    gt8_rxuserrdy_i                              <= GT8_RXUSERRDY_IN or gt8_rxuserrdy_t;
gt9_cpllreset_i                              <= GT9_CPLLRESET_IN or gt9_cpllreset_t;
    gt9_gttxreset_i                              <= GT9_GTTXRESET_IN or gt9_gttxreset_t;
    gt9_gtrxreset_i                              <= GT9_GTRXRESET_IN or gt9_gtrxreset_t;
    gt9_txuserrdy_i                              <= GT9_TXUSERRDY_IN or gt9_txuserrdy_t;
    gt9_rxuserrdy_i                              <= GT9_RXUSERRDY_IN or gt9_rxuserrdy_t;
gt10_cpllreset_i                             <= GT10_CPLLRESET_IN or gt10_cpllreset_t;
    gt10_gttxreset_i                             <= GT10_GTTXRESET_IN or gt10_gttxreset_t;
    gt10_gtrxreset_i                             <= GT10_GTRXRESET_IN or gt10_gtrxreset_t;
    gt10_txuserrdy_i                             <= GT10_TXUSERRDY_IN or gt10_txuserrdy_t;
    gt10_rxuserrdy_i                             <= GT10_RXUSERRDY_IN or gt10_rxuserrdy_t;
gt11_cpllreset_i                             <= GT11_CPLLRESET_IN or gt11_cpllreset_t;
    gt11_gttxreset_i                             <= GT11_GTTXRESET_IN or gt11_gttxreset_t;
    gt11_gtrxreset_i                             <= GT11_GTRXRESET_IN or gt11_gtrxreset_t;
    gt11_txuserrdy_i                             <= GT11_TXUSERRDY_IN or gt11_txuserrdy_t;
    gt11_rxuserrdy_i                             <= GT11_RXUSERRDY_IN or gt11_rxuserrdy_t;
gt12_cpllreset_i                             <= GT12_CPLLRESET_IN or gt12_cpllreset_t;
    gt12_gttxreset_i                             <= GT12_GTTXRESET_IN or gt12_gttxreset_t;
    gt12_gtrxreset_i                             <= GT12_GTRXRESET_IN or gt12_gtrxreset_t;
    gt12_txuserrdy_i                             <= GT12_TXUSERRDY_IN or gt12_txuserrdy_t;
    gt12_rxuserrdy_i                             <= GT12_RXUSERRDY_IN or gt12_rxuserrdy_t;
gt13_cpllreset_i                             <= GT13_CPLLRESET_IN or gt13_cpllreset_t;
    gt13_gttxreset_i                             <= GT13_GTTXRESET_IN or gt13_gttxreset_t;
    gt13_gtrxreset_i                             <= GT13_GTRXRESET_IN or gt13_gtrxreset_t;
    gt13_txuserrdy_i                             <= GT13_TXUSERRDY_IN or gt13_txuserrdy_t;
    gt13_rxuserrdy_i                             <= GT13_RXUSERRDY_IN or gt13_rxuserrdy_t;
gt14_cpllreset_i                             <= GT14_CPLLRESET_IN or gt14_cpllreset_t;
    gt14_gttxreset_i                             <= GT14_GTTXRESET_IN or gt14_gttxreset_t;
    gt14_gtrxreset_i                             <= GT14_GTRXRESET_IN or gt14_gtrxreset_t;
    gt14_txuserrdy_i                             <= GT14_TXUSERRDY_IN or gt14_txuserrdy_t;
    gt14_rxuserrdy_i                             <= GT14_RXUSERRDY_IN or gt14_rxuserrdy_t;
gt15_cpllreset_i                             <= GT15_CPLLRESET_IN or gt15_cpllreset_t;
    gt15_gttxreset_i                             <= GT15_GTTXRESET_IN or gt15_gttxreset_t;
    gt15_gtrxreset_i                             <= GT15_GTRXRESET_IN or gt15_gtrxreset_t;
    gt15_txuserrdy_i                             <= GT15_TXUSERRDY_IN or gt15_txuserrdy_t;
    gt15_rxuserrdy_i                             <= GT15_RXUSERRDY_IN or gt15_rxuserrdy_t;
gt16_cpllreset_i                             <= GT16_CPLLRESET_IN or gt16_cpllreset_t;
    gt16_gttxreset_i                             <= GT16_GTTXRESET_IN or gt16_gttxreset_t;
    gt16_gtrxreset_i                             <= GT16_GTRXRESET_IN or gt16_gtrxreset_t;
    gt16_txuserrdy_i                             <= GT16_TXUSERRDY_IN or gt16_txuserrdy_t;
    gt16_rxuserrdy_i                             <= GT16_RXUSERRDY_IN or gt16_rxuserrdy_t;
gt17_cpllreset_i                             <= GT17_CPLLRESET_IN or gt17_cpllreset_t;
    gt17_gttxreset_i                             <= GT17_GTTXRESET_IN or gt17_gttxreset_t;
    gt17_gtrxreset_i                             <= GT17_GTRXRESET_IN or gt17_gtrxreset_t;
    gt17_txuserrdy_i                             <= GT17_TXUSERRDY_IN or gt17_txuserrdy_t;
    gt17_rxuserrdy_i                             <= GT17_RXUSERRDY_IN or gt17_rxuserrdy_t;
gt18_cpllreset_i                             <= GT18_CPLLRESET_IN or gt18_cpllreset_t;
    gt18_gttxreset_i                             <= GT18_GTTXRESET_IN or gt18_gttxreset_t;
    gt18_gtrxreset_i                             <= GT18_GTRXRESET_IN or gt18_gtrxreset_t;
    gt18_txuserrdy_i                             <= GT18_TXUSERRDY_IN or gt18_txuserrdy_t;
    gt18_rxuserrdy_i                             <= GT18_RXUSERRDY_IN or gt18_rxuserrdy_t;
gt19_cpllreset_i                             <= GT19_CPLLRESET_IN or gt19_cpllreset_t;
    gt19_gttxreset_i                             <= GT19_GTTXRESET_IN or gt19_gttxreset_t;
    gt19_gtrxreset_i                             <= GT19_GTRXRESET_IN or gt19_gtrxreset_t;
    gt19_txuserrdy_i                             <= GT19_TXUSERRDY_IN or gt19_txuserrdy_t;
    gt19_rxuserrdy_i                             <= GT19_RXUSERRDY_IN or gt19_rxuserrdy_t;
end generate chipscope;

no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate
gt0_cpllreset_i                              <= gt0_cpllreset_t;
gt0_gttxreset_i                              <= gt0_gttxreset_t;
gt0_gtrxreset_i                              <= gt0_gtrxreset_t;
gt0_txuserrdy_i                              <= gt0_txuserrdy_t;
gt0_rxuserrdy_i                              <= gt0_rxuserrdy_t;
gt1_cpllreset_i                              <= gt1_cpllreset_t;
gt1_gttxreset_i                              <= gt1_gttxreset_t;
gt1_gtrxreset_i                              <= gt1_gtrxreset_t;
gt1_txuserrdy_i                              <= gt1_txuserrdy_t;
gt1_rxuserrdy_i                              <= gt1_rxuserrdy_t;
gt2_cpllreset_i                              <= gt2_cpllreset_t;
gt2_gttxreset_i                              <= gt2_gttxreset_t;
gt2_gtrxreset_i                              <= gt2_gtrxreset_t;
gt2_txuserrdy_i                              <= gt2_txuserrdy_t;
gt2_rxuserrdy_i                              <= gt2_rxuserrdy_t;
gt3_cpllreset_i                              <= gt3_cpllreset_t;
gt3_gttxreset_i                              <= gt3_gttxreset_t;
gt3_gtrxreset_i                              <= gt3_gtrxreset_t;
gt3_txuserrdy_i                              <= gt3_txuserrdy_t;
gt3_rxuserrdy_i                              <= gt3_rxuserrdy_t;
gt4_cpllreset_i                              <= gt4_cpllreset_t;
gt4_gttxreset_i                              <= gt4_gttxreset_t;
gt4_gtrxreset_i                              <= gt4_gtrxreset_t;
gt4_txuserrdy_i                              <= gt4_txuserrdy_t;
gt4_rxuserrdy_i                              <= gt4_rxuserrdy_t;
gt5_cpllreset_i                              <= gt5_cpllreset_t;
gt5_gttxreset_i                              <= gt5_gttxreset_t;
gt5_gtrxreset_i                              <= gt5_gtrxreset_t;
gt5_txuserrdy_i                              <= gt5_txuserrdy_t;
gt5_rxuserrdy_i                              <= gt5_rxuserrdy_t;
gt6_cpllreset_i                              <= gt6_cpllreset_t;
gt6_gttxreset_i                              <= gt6_gttxreset_t;
gt6_gtrxreset_i                              <= gt6_gtrxreset_t;
gt6_txuserrdy_i                              <= gt6_txuserrdy_t;
gt6_rxuserrdy_i                              <= gt6_rxuserrdy_t;
gt7_cpllreset_i                              <= gt7_cpllreset_t;
gt7_gttxreset_i                              <= gt7_gttxreset_t;
gt7_gtrxreset_i                              <= gt7_gtrxreset_t;
gt7_txuserrdy_i                              <= gt7_txuserrdy_t;
gt7_rxuserrdy_i                              <= gt7_rxuserrdy_t;
gt8_cpllreset_i                              <= gt8_cpllreset_t;
gt8_gttxreset_i                              <= gt8_gttxreset_t;
gt8_gtrxreset_i                              <= gt8_gtrxreset_t;
gt8_txuserrdy_i                              <= gt8_txuserrdy_t;
gt8_rxuserrdy_i                              <= gt8_rxuserrdy_t;
gt9_cpllreset_i                              <= gt9_cpllreset_t;
gt9_gttxreset_i                              <= gt9_gttxreset_t;
gt9_gtrxreset_i                              <= gt9_gtrxreset_t;
gt9_txuserrdy_i                              <= gt9_txuserrdy_t;
gt9_rxuserrdy_i                              <= gt9_rxuserrdy_t;
gt10_cpllreset_i                             <= gt10_cpllreset_t;
gt10_gttxreset_i                             <= gt10_gttxreset_t;
gt10_gtrxreset_i                             <= gt10_gtrxreset_t;
gt10_txuserrdy_i                             <= gt10_txuserrdy_t;
gt10_rxuserrdy_i                             <= gt10_rxuserrdy_t;
gt11_cpllreset_i                             <= gt11_cpllreset_t;
gt11_gttxreset_i                             <= gt11_gttxreset_t;
gt11_gtrxreset_i                             <= gt11_gtrxreset_t;
gt11_txuserrdy_i                             <= gt11_txuserrdy_t;
gt11_rxuserrdy_i                             <= gt11_rxuserrdy_t;
gt12_cpllreset_i                             <= gt12_cpllreset_t;
gt12_gttxreset_i                             <= gt12_gttxreset_t;
gt12_gtrxreset_i                             <= gt12_gtrxreset_t;
gt12_txuserrdy_i                             <= gt12_txuserrdy_t;
gt12_rxuserrdy_i                             <= gt12_rxuserrdy_t;
gt13_cpllreset_i                             <= gt13_cpllreset_t;
gt13_gttxreset_i                             <= gt13_gttxreset_t;
gt13_gtrxreset_i                             <= gt13_gtrxreset_t;
gt13_txuserrdy_i                             <= gt13_txuserrdy_t;
gt13_rxuserrdy_i                             <= gt13_rxuserrdy_t;
gt14_cpllreset_i                             <= gt14_cpllreset_t;
gt14_gttxreset_i                             <= gt14_gttxreset_t;
gt14_gtrxreset_i                             <= gt14_gtrxreset_t;
gt14_txuserrdy_i                             <= gt14_txuserrdy_t;
gt14_rxuserrdy_i                             <= gt14_rxuserrdy_t;
gt15_cpllreset_i                             <= gt15_cpllreset_t;
gt15_gttxreset_i                             <= gt15_gttxreset_t;
gt15_gtrxreset_i                             <= gt15_gtrxreset_t;
gt15_txuserrdy_i                             <= gt15_txuserrdy_t;
gt15_rxuserrdy_i                             <= gt15_rxuserrdy_t;
gt16_cpllreset_i                             <= gt16_cpllreset_t;
gt16_gttxreset_i                             <= gt16_gttxreset_t;
gt16_gtrxreset_i                             <= gt16_gtrxreset_t;
gt16_txuserrdy_i                             <= gt16_txuserrdy_t;
gt16_rxuserrdy_i                             <= gt16_rxuserrdy_t;
gt17_cpllreset_i                             <= gt17_cpllreset_t;
gt17_gttxreset_i                             <= gt17_gttxreset_t;
gt17_gtrxreset_i                             <= gt17_gtrxreset_t;
gt17_txuserrdy_i                             <= gt17_txuserrdy_t;
gt17_rxuserrdy_i                             <= gt17_rxuserrdy_t;
gt18_cpllreset_i                             <= gt18_cpllreset_t;
gt18_gttxreset_i                             <= gt18_gttxreset_t;
gt18_gtrxreset_i                             <= gt18_gtrxreset_t;
gt18_txuserrdy_i                             <= gt18_txuserrdy_t;
gt18_rxuserrdy_i                             <= gt18_rxuserrdy_t;
gt19_cpllreset_i                             <= gt19_cpllreset_t;
gt19_gttxreset_i                             <= gt19_gttxreset_t;
gt19_gtrxreset_i                             <= gt19_gtrxreset_t;
gt19_txuserrdy_i                             <= gt19_txuserrdy_t;
gt19_rxuserrdy_i                             <= gt19_rxuserrdy_t;
end generate no_chipscope;


gt0_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT0_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt0_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt0_cplllock_i,
        TXRESETDONE                     =>      gt0_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt0_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt0_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT0_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt0_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt1_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT1_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt1_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt1_cplllock_i,
        TXRESETDONE                     =>      gt1_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt1_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt1_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT1_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt1_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt2_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT2_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt2_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt2_cplllock_i,
        TXRESETDONE                     =>      gt2_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt2_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt2_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT2_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt2_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt3_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT3_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt3_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt3_cplllock_i,
        TXRESETDONE                     =>      gt3_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt3_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt3_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT3_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt3_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt4_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT4_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt4_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt4_cplllock_i,
        TXRESETDONE                     =>      gt4_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt4_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt4_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT4_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt4_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt5_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT5_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt5_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt5_cplllock_i,
        TXRESETDONE                     =>      gt5_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt5_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt5_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT5_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt5_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt6_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT6_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt6_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt6_cplllock_i,
        TXRESETDONE                     =>      gt6_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt6_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt6_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT6_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt6_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt7_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT7_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt7_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt7_cplllock_i,
        TXRESETDONE                     =>      gt7_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt7_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt7_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT7_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt7_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt8_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT8_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt8_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt8_cplllock_i,
        TXRESETDONE                     =>      gt8_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt8_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt8_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT8_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt8_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt9_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT9_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt9_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt9_cplllock_i,
        TXRESETDONE                     =>      gt9_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt9_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt9_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT9_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt9_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt10_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT10_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt10_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt10_cplllock_i,
        TXRESETDONE                     =>      gt10_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt10_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt10_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT10_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt10_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt11_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT11_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt11_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt11_cplllock_i,
        TXRESETDONE                     =>      gt11_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt11_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt11_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT11_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt11_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt12_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT12_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt12_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt12_cplllock_i,
        TXRESETDONE                     =>      gt12_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt12_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt12_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT12_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt12_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt13_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT13_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt13_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt13_cplllock_i,
        TXRESETDONE                     =>      gt13_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt13_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt13_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT13_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt13_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt14_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT14_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt14_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt14_cplllock_i,
        TXRESETDONE                     =>      gt14_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt14_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt14_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT14_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt14_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt15_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT15_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt15_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt15_cplllock_i,
        TXRESETDONE                     =>      gt15_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt15_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt15_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT15_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt15_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt16_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT16_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt16_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt16_cplllock_i,
        TXRESETDONE                     =>      gt16_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt16_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt16_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT16_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt16_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt17_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT17_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt17_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt17_cplllock_i,
        TXRESETDONE                     =>      gt17_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt17_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt17_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT17_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt17_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt18_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT18_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt18_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt18_cplllock_i,
        TXRESETDONE                     =>      gt18_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt18_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt18_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT18_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt18_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );

gt19_txresetfsm_i:  gt625_fab20_TX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           -- Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   => FALSE                 -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        TXUSERCLK                       =>      GT19_TXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt19_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt19_cplllock_i,
        TXRESETDONE                     =>      gt19_txresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        GTTXRESET                       =>      gt19_gttxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      gt19_cpllreset_t,
        TX_FSM_RESET_DONE               =>      GT19_TX_FSM_RESET_DONE_OUT,
        TXUSERRDY                       =>      gt19_txuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RETRY_COUNTER                   =>      open
           );







gt0_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT0_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt0_rxusrclk_in,
        TXPMARESETDONE                  =>      gt0_txpmaresetdone_i,
        TXOUTCLK                        =>      gt0_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt0_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt0_cplllock_i,
        RXRESETDONE                     =>      gt0_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT0_DATA_VALID_IN,
        TXUSERRDY                       =>      gt0_txuserrdy_i,
        GTRXRESET                       =>      gt0_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT0_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt0_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt0_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt0_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt0_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt0_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt1_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT1_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt1_rxusrclk_in,
        TXPMARESETDONE                  =>      gt1_txpmaresetdone_i,
        TXOUTCLK                        =>      gt1_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt1_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt1_cplllock_i,
        RXRESETDONE                     =>      gt1_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT1_DATA_VALID_IN,
        TXUSERRDY                       =>      gt1_txuserrdy_i,
        GTRXRESET                       =>      gt1_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT1_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt1_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt1_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt1_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt1_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt1_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt2_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT2_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt2_rxusrclk_in,
        TXPMARESETDONE                  =>      gt2_txpmaresetdone_i,
        TXOUTCLK                        =>      gt2_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt2_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt2_cplllock_i,
        RXRESETDONE                     =>      gt2_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT2_DATA_VALID_IN,
        TXUSERRDY                       =>      gt2_txuserrdy_i,
        GTRXRESET                       =>      gt2_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT2_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt2_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt2_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt2_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt2_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt2_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt3_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT3_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt3_rxusrclk_in,
        TXPMARESETDONE                  =>      gt3_txpmaresetdone_i,
        TXOUTCLK                        =>      gt3_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt3_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt3_cplllock_i,
        RXRESETDONE                     =>      gt3_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT3_DATA_VALID_IN,
        TXUSERRDY                       =>      gt3_txuserrdy_i,
        GTRXRESET                       =>      gt3_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT3_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt3_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt3_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt3_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt3_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt3_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt4_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT4_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt4_rxusrclk_in,
        TXPMARESETDONE                  =>      gt4_txpmaresetdone_i,
        TXOUTCLK                        =>      gt4_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt4_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt4_cplllock_i,
        RXRESETDONE                     =>      gt4_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT4_DATA_VALID_IN,
        TXUSERRDY                       =>      gt4_txuserrdy_i,
        GTRXRESET                       =>      gt4_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT4_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt4_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt4_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt4_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt4_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt4_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt5_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT5_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt5_rxusrclk_in,
        TXPMARESETDONE                  =>      gt5_txpmaresetdone_i,
        TXOUTCLK                        =>      gt5_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt5_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt5_cplllock_i,
        RXRESETDONE                     =>      gt5_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT5_DATA_VALID_IN,
        TXUSERRDY                       =>      gt5_txuserrdy_i,
        GTRXRESET                       =>      gt5_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT5_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt5_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt5_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt5_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt5_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt5_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt6_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT6_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt6_rxusrclk_in,
        TXPMARESETDONE                  =>      gt6_txpmaresetdone_i,
        TXOUTCLK                        =>      gt6_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt6_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt6_cplllock_i,
        RXRESETDONE                     =>      gt6_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT6_DATA_VALID_IN,
        TXUSERRDY                       =>      gt6_txuserrdy_i,
        GTRXRESET                       =>      gt6_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT6_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt6_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt6_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt6_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt6_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt6_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt7_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT7_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt7_rxusrclk_in,
        TXPMARESETDONE                  =>      gt7_txpmaresetdone_i,
        TXOUTCLK                        =>      gt7_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt7_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt7_cplllock_i,
        RXRESETDONE                     =>      gt7_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT7_DATA_VALID_IN,
        TXUSERRDY                       =>      gt7_txuserrdy_i,
        GTRXRESET                       =>      gt7_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT7_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt7_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt7_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt7_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt7_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt7_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt8_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT8_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt8_rxusrclk_in,
        TXPMARESETDONE                  =>      gt8_txpmaresetdone_i,
        TXOUTCLK                        =>      gt8_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt8_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt8_cplllock_i,
        RXRESETDONE                     =>      gt8_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT8_DATA_VALID_IN,
        TXUSERRDY                       =>      gt8_txuserrdy_i,
        GTRXRESET                       =>      gt8_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT8_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt8_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt8_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt8_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt8_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt8_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt9_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT9_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt9_rxusrclk_in,
        TXPMARESETDONE                  =>      gt9_txpmaresetdone_i,
        TXOUTCLK                        =>      gt9_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt9_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt9_cplllock_i,
        RXRESETDONE                     =>      gt9_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT9_DATA_VALID_IN,
        TXUSERRDY                       =>      gt9_txuserrdy_i,
        GTRXRESET                       =>      gt9_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT9_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt9_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt9_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt9_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt9_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt9_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt10_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT10_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt10_rxusrclk_in,
        TXPMARESETDONE                  =>      gt10_txpmaresetdone_i,
        TXOUTCLK                        =>      gt10_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt10_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt10_cplllock_i,
        RXRESETDONE                     =>      gt10_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT10_DATA_VALID_IN,
        TXUSERRDY                       =>      gt10_txuserrdy_i,
        GTRXRESET                       =>      gt10_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT10_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt10_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt10_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt10_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt10_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt10_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt11_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT11_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt11_rxusrclk_in,
        TXPMARESETDONE                  =>      gt11_txpmaresetdone_i,
        TXOUTCLK                        =>      gt11_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt11_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt11_cplllock_i,
        RXRESETDONE                     =>      gt11_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT11_DATA_VALID_IN,
        TXUSERRDY                       =>      gt11_txuserrdy_i,
        GTRXRESET                       =>      gt11_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT11_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt11_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt11_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt11_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt11_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt11_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt12_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT12_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt12_rxusrclk_in,
        TXPMARESETDONE                  =>      gt12_txpmaresetdone_i,
        TXOUTCLK                        =>      gt12_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt12_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt12_cplllock_i,
        RXRESETDONE                     =>      gt12_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT12_DATA_VALID_IN,
        TXUSERRDY                       =>      gt12_txuserrdy_i,
        GTRXRESET                       =>      gt12_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT12_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt12_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt12_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt12_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt12_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt12_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt13_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT13_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt13_rxusrclk_in,
        TXPMARESETDONE                  =>      gt13_txpmaresetdone_i,
        TXOUTCLK                        =>      gt13_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt13_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt13_cplllock_i,
        RXRESETDONE                     =>      gt13_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT13_DATA_VALID_IN,
        TXUSERRDY                       =>      gt13_txuserrdy_i,
        GTRXRESET                       =>      gt13_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT13_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt13_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt13_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt13_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt13_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt13_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt14_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT14_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt14_rxusrclk_in,
        TXPMARESETDONE                  =>      gt14_txpmaresetdone_i,
        TXOUTCLK                        =>      gt14_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt14_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt14_cplllock_i,
        RXRESETDONE                     =>      gt14_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT14_DATA_VALID_IN,
        TXUSERRDY                       =>      gt14_txuserrdy_i,
        GTRXRESET                       =>      gt14_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT14_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt14_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt14_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt14_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt14_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt14_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt15_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT15_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt15_rxusrclk_in,
        TXPMARESETDONE                  =>      gt15_txpmaresetdone_i,
        TXOUTCLK                        =>      gt15_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt15_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt15_cplllock_i,
        RXRESETDONE                     =>      gt15_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT15_DATA_VALID_IN,
        TXUSERRDY                       =>      gt15_txuserrdy_i,
        GTRXRESET                       =>      gt15_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT15_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt15_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt15_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt15_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt15_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt15_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt16_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT16_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt16_rxusrclk_in,
        TXPMARESETDONE                  =>      gt16_txpmaresetdone_i,
        TXOUTCLK                        =>      gt16_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt16_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt16_cplllock_i,
        RXRESETDONE                     =>      gt16_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT16_DATA_VALID_IN,
        TXUSERRDY                       =>      gt16_txuserrdy_i,
        GTRXRESET                       =>      gt16_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT16_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt16_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt16_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt16_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt16_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt16_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt17_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT17_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt17_rxusrclk_in,
        TXPMARESETDONE                  =>      gt17_txpmaresetdone_i,
        TXOUTCLK                        =>      gt17_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt17_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt17_cplllock_i,
        RXRESETDONE                     =>      gt17_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT17_DATA_VALID_IN,
        TXUSERRDY                       =>      gt17_txuserrdy_i,
        GTRXRESET                       =>      gt17_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT17_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt17_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt17_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt17_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt17_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt17_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt18_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT18_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt18_rxusrclk_in,
        TXPMARESETDONE                  =>      gt18_txpmaresetdone_i,
        TXOUTCLK                        =>      gt18_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt18_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt18_cplllock_i,
        RXRESETDONE                     =>      gt18_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT18_DATA_VALID_IN,
        TXUSERRDY                       =>      gt18_txuserrdy_i,
        GTRXRESET                       =>      gt18_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT18_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt18_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt18_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt18_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt18_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt18_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



gt19_rxresetfsm_i:  gt625_fab20_RX_STARTUP_FSM 

  generic map(
           EXAMPLE_SIMULATION       => EXAMPLE_SIMULATION,
           EQ_MODE                  => "DFE",                 --Rx Equalization Mode - Set to DFE or LPM
           STABLE_CLOCK_PERIOD      => STABLE_CLOCK_PERIOD,           --Period of the stable clock driving this state-machine, unit is [ns]
           RETRY_COUNTER_BITWIDTH   => 8, 
           TX_QPLL_USED             => FALSE ,                       -- the TX and RX Reset FSMs must
           RX_QPLL_USED             => FALSE,                        -- share these two generic values
           PHASE_ALIGNMENT_MANUAL   =>  FALSE                        -- Decision if a manual phase-alignment is necessary or the automatic 
                                                                     -- is enough. For single-lane applications the automatic alignment is 
                                                                     -- sufficient              
             )     
    port map ( 
        STABLE_CLOCK                    =>      SYSCLK_IN,
        RXUSERCLK                       =>      GT19_RXUSRCLK_IN,
        SOFT_RESET                      =>      SOFT_RESET_IN,
        DONT_RESET_ON_DATA_ERROR        =>      DONT_RESET_ON_DATA_ERROR_IN,
        RXPMARESETDONE                  =>      gt0_rxpmaresetdone_i,
        RXOUTCLK                        =>      gt19_rxusrclk_in,
        TXPMARESETDONE                  =>      gt19_txpmaresetdone_i,
        TXOUTCLK                        =>      gt19_txusrclk_in,
        QPLLREFCLKLOST                  =>      tied_to_ground_i,
        CPLLREFCLKLOST                  =>      gt19_cpllrefclklost_i,
        QPLLLOCK                        =>      tied_to_vcc_i,
        CPLLLOCK                        =>      gt19_cplllock_i,
        RXRESETDONE                     =>      gt19_rxresetdone_i,
        MMCM_LOCK                       =>      tied_to_vcc_i,
        RECCLK_STABLE                   =>      gt0_recclk_stable_i,
        RECCLK_MONITOR_RESTART          =>      tied_to_ground_i,
        DATA_VALID                      =>      GT19_DATA_VALID_IN,
        TXUSERRDY                       =>      gt19_txuserrdy_i,
        GTRXRESET                       =>      gt19_gtrxreset_t,
        MMCM_RESET                      =>      open,
        QPLL_RESET                      =>      open,
        CPLL_RESET                      =>      open,
        RX_FSM_RESET_DONE               =>      GT19_RX_FSM_RESET_DONE_OUT,
        RXUSERRDY                       =>      gt19_rxuserrdy_t,
        RUN_PHALIGNMENT                 =>      open,
        RESET_PHALIGNMENT               =>      open,
        PHALIGNMENT_DONE                =>      tied_to_vcc_i,
        RXDFEAGCHOLD                    =>      gt19_rxdfeagchold_i,
        RXDFELFHOLD                     =>      gt19_rxdfelfhold_i,
        RXLPMLFHOLD                     =>      gt19_rxlpmlfhold_i,
        RXLPMHFHOLD                     =>      gt19_rxlpmhfhold_i,
        RETRY_COUNTER                   =>      open
           );



  gt0_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt0_gtrxreset_i = '1') then
          gt0_rx_cdrlocked       <= '0';
          gt0_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt0_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt0_rx_cdrlocked       <= '1';
          gt0_rx_cdrlock_counter <= gt0_rx_cdrlock_counter        after DLY;
        else
          gt0_rx_cdrlock_counter <= gt0_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt1_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt1_gtrxreset_i = '1') then
          gt1_rx_cdrlocked       <= '0';
          gt1_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt1_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt1_rx_cdrlocked       <= '1';
          gt1_rx_cdrlock_counter <= gt1_rx_cdrlock_counter        after DLY;
        else
          gt1_rx_cdrlock_counter <= gt1_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt2_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt2_gtrxreset_i = '1') then
          gt2_rx_cdrlocked       <= '0';
          gt2_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt2_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt2_rx_cdrlocked       <= '1';
          gt2_rx_cdrlock_counter <= gt2_rx_cdrlock_counter        after DLY;
        else
          gt2_rx_cdrlock_counter <= gt2_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt3_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt3_gtrxreset_i = '1') then
          gt3_rx_cdrlocked       <= '0';
          gt3_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt3_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt3_rx_cdrlocked       <= '1';
          gt3_rx_cdrlock_counter <= gt3_rx_cdrlock_counter        after DLY;
        else
          gt3_rx_cdrlock_counter <= gt3_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt4_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt4_gtrxreset_i = '1') then
          gt4_rx_cdrlocked       <= '0';
          gt4_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt4_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt4_rx_cdrlocked       <= '1';
          gt4_rx_cdrlock_counter <= gt4_rx_cdrlock_counter        after DLY;
        else
          gt4_rx_cdrlock_counter <= gt4_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt5_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt5_gtrxreset_i = '1') then
          gt5_rx_cdrlocked       <= '0';
          gt5_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt5_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt5_rx_cdrlocked       <= '1';
          gt5_rx_cdrlock_counter <= gt5_rx_cdrlock_counter        after DLY;
        else
          gt5_rx_cdrlock_counter <= gt5_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt6_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt6_gtrxreset_i = '1') then
          gt6_rx_cdrlocked       <= '0';
          gt6_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt6_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt6_rx_cdrlocked       <= '1';
          gt6_rx_cdrlock_counter <= gt6_rx_cdrlock_counter        after DLY;
        else
          gt6_rx_cdrlock_counter <= gt6_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt7_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt7_gtrxreset_i = '1') then
          gt7_rx_cdrlocked       <= '0';
          gt7_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt7_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt7_rx_cdrlocked       <= '1';
          gt7_rx_cdrlock_counter <= gt7_rx_cdrlock_counter        after DLY;
        else
          gt7_rx_cdrlock_counter <= gt7_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt8_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt8_gtrxreset_i = '1') then
          gt8_rx_cdrlocked       <= '0';
          gt8_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt8_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt8_rx_cdrlocked       <= '1';
          gt8_rx_cdrlock_counter <= gt8_rx_cdrlock_counter        after DLY;
        else
          gt8_rx_cdrlock_counter <= gt8_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt9_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt9_gtrxreset_i = '1') then
          gt9_rx_cdrlocked       <= '0';
          gt9_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt9_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt9_rx_cdrlocked       <= '1';
          gt9_rx_cdrlock_counter <= gt9_rx_cdrlock_counter        after DLY;
        else
          gt9_rx_cdrlock_counter <= gt9_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt10_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt10_gtrxreset_i = '1') then
          gt10_rx_cdrlocked       <= '0';
          gt10_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt10_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt10_rx_cdrlocked       <= '1';
          gt10_rx_cdrlock_counter <= gt10_rx_cdrlock_counter        after DLY;
        else
          gt10_rx_cdrlock_counter <= gt10_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt11_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt11_gtrxreset_i = '1') then
          gt11_rx_cdrlocked       <= '0';
          gt11_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt11_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt11_rx_cdrlocked       <= '1';
          gt11_rx_cdrlock_counter <= gt11_rx_cdrlock_counter        after DLY;
        else
          gt11_rx_cdrlock_counter <= gt11_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt12_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt12_gtrxreset_i = '1') then
          gt12_rx_cdrlocked       <= '0';
          gt12_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt12_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt12_rx_cdrlocked       <= '1';
          gt12_rx_cdrlock_counter <= gt12_rx_cdrlock_counter        after DLY;
        else
          gt12_rx_cdrlock_counter <= gt12_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt13_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt13_gtrxreset_i = '1') then
          gt13_rx_cdrlocked       <= '0';
          gt13_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt13_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt13_rx_cdrlocked       <= '1';
          gt13_rx_cdrlock_counter <= gt13_rx_cdrlock_counter        after DLY;
        else
          gt13_rx_cdrlock_counter <= gt13_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt14_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt14_gtrxreset_i = '1') then
          gt14_rx_cdrlocked       <= '0';
          gt14_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt14_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt14_rx_cdrlocked       <= '1';
          gt14_rx_cdrlock_counter <= gt14_rx_cdrlock_counter        after DLY;
        else
          gt14_rx_cdrlock_counter <= gt14_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt15_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt15_gtrxreset_i = '1') then
          gt15_rx_cdrlocked       <= '0';
          gt15_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt15_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt15_rx_cdrlocked       <= '1';
          gt15_rx_cdrlock_counter <= gt15_rx_cdrlock_counter        after DLY;
        else
          gt15_rx_cdrlock_counter <= gt15_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt16_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt16_gtrxreset_i = '1') then
          gt16_rx_cdrlocked       <= '0';
          gt16_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt16_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt16_rx_cdrlocked       <= '1';
          gt16_rx_cdrlock_counter <= gt16_rx_cdrlock_counter        after DLY;
        else
          gt16_rx_cdrlock_counter <= gt16_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt17_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt17_gtrxreset_i = '1') then
          gt17_rx_cdrlocked       <= '0';
          gt17_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt17_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt17_rx_cdrlocked       <= '1';
          gt17_rx_cdrlock_counter <= gt17_rx_cdrlock_counter        after DLY;
        else
          gt17_rx_cdrlock_counter <= gt17_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt18_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt18_gtrxreset_i = '1') then
          gt18_rx_cdrlocked       <= '0';
          gt18_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt18_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt18_rx_cdrlocked       <= '1';
          gt18_rx_cdrlock_counter <= gt18_rx_cdrlock_counter        after DLY;
        else
          gt18_rx_cdrlock_counter <= gt18_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

  gt19_cdrlock_timeout:process(SYSCLK_IN)
  begin
    if rising_edge(SYSCLK_IN) then
        if(gt19_gtrxreset_i = '1') then
          gt19_rx_cdrlocked       <= '0';
          gt19_rx_cdrlock_counter <=  0                        after DLY;
        elsif (gt19_rx_cdrlock_counter = WAIT_TIME_CDRLOCK) then
          gt19_rx_cdrlocked       <= '1';
          gt19_rx_cdrlock_counter <= gt19_rx_cdrlock_counter        after DLY;
        else
          gt19_rx_cdrlock_counter <= gt19_rx_cdrlock_counter + 1    after DLY;
        end if;
    end if;
  end process;

gt0_recclk_stable_i                          <= gt0_rx_cdrlocked;
gt1_recclk_stable_i                          <= gt1_rx_cdrlocked;
gt2_recclk_stable_i                          <= gt2_rx_cdrlocked;
gt3_recclk_stable_i                          <= gt3_rx_cdrlocked;
gt4_recclk_stable_i                          <= gt4_rx_cdrlocked;
gt5_recclk_stable_i                          <= gt5_rx_cdrlocked;
gt6_recclk_stable_i                          <= gt6_rx_cdrlocked;
gt7_recclk_stable_i                          <= gt7_rx_cdrlocked;
gt8_recclk_stable_i                          <= gt8_rx_cdrlocked;
gt9_recclk_stable_i                          <= gt9_rx_cdrlocked;
gt10_recclk_stable_i                         <= gt10_rx_cdrlocked;
gt11_recclk_stable_i                         <= gt11_rx_cdrlocked;
gt12_recclk_stable_i                         <= gt12_rx_cdrlocked;
gt13_recclk_stable_i                         <= gt13_rx_cdrlocked;
gt14_recclk_stable_i                         <= gt14_rx_cdrlocked;
gt15_recclk_stable_i                         <= gt15_rx_cdrlocked;
gt16_recclk_stable_i                         <= gt16_rx_cdrlocked;
gt17_recclk_stable_i                         <= gt17_rx_cdrlocked;
gt18_recclk_stable_i                         <= gt18_rx_cdrlocked;
gt19_recclk_stable_i                         <= gt19_rx_cdrlocked;






end RTL;


