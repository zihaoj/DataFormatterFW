

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OL+7PuFhC190RFP7e+AUu2IwNMZeB+mjrn6VItJWaLbGVPLrIcd9f78El8TYO0Uy7lRe5ft5SG2L
QUOqGhS+bw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VPsFGy1y1wgsMAZW77DuRZ4GutmU5OkV0iRZPhYBVx9VtlhryYQGswGtazJjXA2BlCFP3RyKiMb5
GCm8MLSZXhTHeqCF5kNmqJW8oV1xNCv2wHK1MdmB5hzNibB0BUtHn7PPyTfI6OsUwOqdWZEgImnN
iStGdsiv2p7qhWC0+U8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qh6C1lhwxlHVu+7MJQcLaeJR8bmBds7YkhWQ3IKMJFLdp22terTtjeK+FkKlTVLJmgSlUHuS8hHZ
O0ip0hGAWsFlfnJ/suALOKMAuKA2zc03QFG3dPx1dIKsMvsmwfnbBUvkXNHSCg702gCLrnsYvs3+
0KhNBWo+L4FIwRHrQzZv7SoLOg1PgkoZ9CYlvjM7lN9dd/jYSanNNHUgm7iFyDqaA4mb7giMCe9+
YKuBm4YCdLJ+SGpOqhMMTGNPLR909t5y+tvtPy7R+zfDtEtEEMJ1b7kj8RGqah6/mdGh8cEqszm+
R1S8UTmK9XmWHdabqMEKEJKIcAX7TkBaZrkFwA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
b61GiEWADTXp3mmaNejvwcWhBNwq8suwg3OsO0zXUc5URzQo+mfd1gMBe+DTsL/Bywz02OwSg69Z
Esvmxb3VLofUhTusvBo/r+3mV8pfqEV9V0qauDpQ5Sjg4vwdRszVkMKMVk7zTAEPVl34izdUHywF
zzhPIlqqbmnxgqC5qXE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SRWrXFPT2M4Fcu0ySSCN8VT8Ci/aHGWte0qUXDTMhiHbKg1CY7t2TQYn8IZc7S+YVCIoxPZhDEli
etbwk87hs2cCYdbyLJxVv4RvsNUpm+MTjOU62spjCEATs5hM4/Ddzx6SJUQB3z7yUczs10IDIJwv
sknFAEmPlnMxjgjf8+x/1YFmhs7yAZn6Iu7HvrJ5qYE0wSxbVFJnyOZPro5I75+fm4qfewvcC+Zx
WtC2WQ5k1b2ynh5ZSV5V3N7qTg8VCQqp4DgeLmegSuIUqtRXZwLN/vUOUubsyFtJXzS8bdIOeAlF
kotfCLX4k0RzjtPpRIYcmtxiRBUZnak30YgVzg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6432)
`protect data_block
4KmXUDwrycHN2EiBeRO2lYBVShUyAhHkCMI0ahIZDkBww/Y+T6x3VCDKamHx7T9BOZDohxsjWyp5
XjNiipLmUIQo+yO+Tiz8COumCxen7zkL0dFN+Yeuzoa/ZyOiwq9tkk8B35doxtIhEUc8msm8hI/K
5qRxxsUKzjraSCr5p4ogLXH9KQxI0fOejhiJvBR2PVaElU7GXEKKQJnHoK0kBCiDb8y17oPPNNw4
vHOGIGhHjMIUEcQiQHxSCjI26Qr8oJvG2bFRHFCmFRDYDaHrnBoX1OAUjn82CSa/i9BezSpEET6i
0iqplmAzripd3GyuaYpyuySNgNq4r/MMoqDR6jIsVlYHOEzg8ZJOD58f0ElTMXaPuaAf6aQp8ZyO
LPs2ZP8CofouNgyTWtYCwcK9hD6D7AGhv49kJPgqTaMWLqNiA7XAAkznl1V8YjYrqBOMdUlREceZ
iqyN/eaeE+iVVkwKoWld6IQ33+0QlXl6OK8lH1I4jgoHXpuM239MaCIKY3VY/6l4gZaqo14+PZgV
x/9Qa9xyzwpaZxYXtbuXE41hVDaqNaLO67EG+umBfeKbYTOGUewR2vZfEWmMeZyStTRpDVYVwWBU
4XgFLjdQIeXUVHhd+/+ttInMd4B0jTmKKEARLHQodxQK1h+31UJoe9RSdZW+OU0EpI9Xs9tCX1oL
W7KH9+KJE8ez+QSKSf2uEzEhnvxuL5SZvTQiXeGQOlMr34Yv6As7EYaYqvvN75boiaSNrSKSxvrt
oljNrpJMXolPz9Hvoh8fCh+ISVnX4iVfxTom7QuBXHyls/ZVLVR6yUxdBAT8FipEyI3osXoYqlKc
qSNoXDddRqnW4/D68LkKWbKr6fG+Ys6Q+ZwrP8fmAi9gJOYsjkQsog9JqdNd5ABdsMOXocVqdXI1
l47ihQK3REi052J3RxbGgHBI6E0bp8PaD7gI0Nz27CJ1upT6iSMxmMoDHK7Y8vZ8Z0Za4QQRWc9q
Pea6Acst3WvMUnjfIE5+uGczzzW89zPLmBugE2FcD6l0lujMRat0vzhQ+9E8doTfds7JMtnpVOWT
PuM9au/qeVgYiz1jUOLCVPk1nyqUzCv9sqj7PHWbUqIysOYNsQEPky0+7TVZ6HYq5JEV82HpFYZW
R1Cb8PvicAmeUrfrTzeitrpnshRiFmB/vlIC+oMZxKO7F8bfcZMqw7F+CEwm0VcDJJeZ+TaLdRsJ
y2EDRTJVU5jVZZYfWnBtryMEWqMVD/Bk0m8/0SRLZ5hcFh8hBbPkgvWNhII55DCFEPi1nqKAi2Je
Xiu/5PTfZH1Tcwp+tshEoGOjwh/QLiKzl3EGY6oVYzH8CMsWWpQQtPnsNowkafTsyxdmka0C+/XW
CE1YO8lL2h4Nz8iw99BljuYf6d3jUO8HegQzDgFkghOE5+tDoG180oy+YoOFFGFtgtXNJTwqf20P
sgPx+3apHoxJ116FLsU6kHirwY+t3qyGPvAf7Xin0rNL2gwcx8Luh0mRj8lCGPdKz3gkWKC1hqKJ
skv5TC36bkioqHiVE6YlhGX9q3xmBTXmUbsmlku3k6hlGe3EclxffDtALq1yidnOJonrlf1QEGeo
obKeTgzZ1DzU75MiHzN85OUZHRVmb+Jmxo/2mCdswsUFJrTKbgSy736SSEcbBxrgsV2eSfBK+yoY
VP7JyH2zbGjo1zuGSB29nUSys/s7WjGQY8gYgfa/YpHgj1Z2fgXLq0rO7w0HfPLTxA53eLm14Iyl
RNOak6qWgG1MLZHYpJbZBq5GaGFj+iKj4YMc/THY49sJkA2wTHSiPuGlXCxL0JxZoQQv01X7N+u4
g3sCQ0DaONcBLDGCgaaEdwJohRCKbji0yhiUt+g2ye3jO6pT7uQkLKLjTKHASHAxIBP3eH4XE5vY
QM3vMezBD57+jI08lr7rTFqhzBC/6NxTkQLqQyrjm8Wg7fjMTcL+UaoiiDCULi+rsVzp6VCVPj79
V+xcDCVRiJuChZRU+whvADdJD2vcfKFBTjvn4i3qdBQwWA5Ck3hciGwUAAX9zQJ5LcI6K2elCRyo
Lxja9sHDXv+vvf1sPLjS3M9o9ITzpUFLqVQ0dcXeq1AHg8dlRbC9XVH6eG44GcHpyAf8fxNrmllg
5x65IU2Ynbfpz85UiSVSTjrLZgzwhbr9QcO5Jg/RD/J7f7DeS2pSLePEF1qaZUywQkRJ+C1BkCEe
mrXe79l28Y84iKkSK1hFzUiTp9PSzWaPwkmOg1hm6b6CrJI+uW7c9YJH5yl8l3JZmK4bvRYw7Pc+
9kMiCrH5fG8VIWdMrT2crtCxWBDa0T/d5NIQWb7RYpYgi8NWJL5TTcMyndrdErlim2G8Op3wj5yZ
SU257cqFvJRle/xulO/AalZDy9AdzDmhbvLImC7CzGeOrn8qcfECKGhfy/o9Wwq4NC8R15W7nIZN
pK0L9ia3IZoDKJ0ItUn2q/6/vqVtNq59YWgDyfJxTqV3kKM0z6weAjyP48MLnKXCsbvg9tznnmdx
LWOjSBGdMNvdQj2D14G/+fsK5CORee0d2TQ2DgjNF/H+R02kkxuiKWLTn5uz6YYJEq1RVe4XJgq+
8zBIYQLVKM1G8Xk09GnKpKmaa2wNGzPWcUJI+mWMpSgSKcMTTzwxWFjOMEsna+g3vL2pH4ZFP7lA
z4bIIEsD7vn7CFxag/7M7+f9T15EUC3J+zkqgoyHEmrUN6x5Sec1b9Osvw1O5u3DyEpHih91oq0q
HW3xZmtQrRLHRHokzkqhSspTM1g27eCEGzRs/vTFblSZiFX9mY6dJePBhzkxoHNFrKrTJsq8aUU3
mQkGWYmbZDHc32pz+U5jkR5nkPTqkIQ9Y6DmypdP5fYe0O2xl9kOcVWRENdWZ3iqjjJfm+4NceLD
wMzb6lWjFibYetbEYaDTPos3zhpwl3H2v/Wg6V85ebkhGLLJrJ4MZ0m+U+Tnx0Kvk6oGNHLFU22q
LSO2eIuIUJxqU/74s8pJ7dv1d3EMkxh3oy+UYdEl152hCpejFBx8WfqejFn44ApKT3K/HOeN+7aQ
Htg1uh7zrM4/8ik8rtSBgEYspXyQINCrh/n2U1UTnhPDnzkU3mq3MUTroOrmZOsg7/WaGbzO3CF8
S9HKaQyrp+VFCDGkwbM3tqXfGxDD0ZdXPi+8ghJk3Ha5w6S80MNsY7xFzeTarsJ7LJikMh24ZBp3
W5UDxBelE4SPwpHTQp4t24vdqwyZ4qbIvldTcor3hjqUw/8h0JMaKp8K7zYQXX1vlJ6HQ7cMLi77
g/FhKkfP9Tzu166ARRXpelB73AkI0nxHQXgSJ745vyUUdreva4Csl+e50GlgjNLPYgq1CQS4hk8q
5bYW5uIXMeAmC97C/5HzLYi0R8BqI1pcCuSwPRkqUpafBEvAzoQqtB4T4PEruWOn95WJoSeR7YBU
11pMTXYforTZ5XTlSBSuPMW95G5esvtXSxJs8FlDk8Kr2MNMD8QgwmR/QVh8cj3gfPzUVcGxTx8s
8IxxA8IwvvYSmNgxmyRKsdjW2VzDTpy0VzwzgYkIeZhcMXbkaeLSZMZT5bBN06WW16WveNAzHSNo
7oujJzckh4nkdA0g0yMxwCI3AwyGDvOahgjCKGs8rza1RZC2WE8ue6qP3T0fMOgakMDzX4OfMfgw
KoRs7VZtvHGWEjwH2Szwtxl4yE+upweHg1K4Uua4Gx7NinBCrs70yhVaCAb+G1yGFvoaqO6wJ4JN
95Pdkad/SyXbIYmmjl67R86WfUVS8FVIa8kx7a8sAX1obj1JSHufbuPN/WJvyHp6+82AxvfNlOU9
RpGeAu1BNpUfrzfgYbmTK4nSTaRsWgcXGewyyZoVTOxEJn3uFi5jXHePrQXkKigiwZVZl+rzZvcg
UmWEe7y6wziLPDBP8ARYHzds9ESBdaQwD4d85qiuMuPQL85b9BcLu7yjGM6wTo0ZQMroUkWf8hDZ
XjyJrn19j2MArPoHeos34m/ZVEzdV+DfH+fqlZ2ihrwsjjn45pPSmIAcYzcM2DmKM/jEXC0Hf42G
41syuHkHiPj4WQcXkDNi9kM6JFH3B5RtEE96DJRBGvIxwBulOzb135mnK6N5CQnXg0QUF7lFh+M2
lWlOsFtPG8VV8p6o/fd78q8pfpDSkP7Be/Y8J260Tk8+chuEh/S8pfGxjCZzpPMWSuXrc4ZJAt+4
dvmG80XeqBz+zYGwX2P80jUeZmrJTDGqvMxyaaSM8kNsyT9Lv+JH3OXV97XCLVon+SeTOsBSTJ5+
TAOnUyd3DVyX9MciLDZQn77rXhDlVJP2JqOExW+tXpSSEdXC8vyFqjJW1LtAeppgWOQJ4qdTzFWr
453yz7cGnlPK467AT62UXgcRGlHPnT2WARGvVGTOXp4pM4JGhds0i3sizC7+0jzn/oeOQnl3Z+WE
7knBcKoO2omBdjt+/AFZgl9U//K8RP4iY82IOODYm8n7gLeZjz7kXxHxjb29IyZpvG4m1EKEM3PG
oiw6iymNmu61LVaXNUK/vmTLWP0QRViSufnj5cfCnf4Z5Fr2nlkam6v7RCHolj6BTf3jDGamUTOQ
Cxc4p36BAC3ayg3Nc1ZhNpoN8IMgGgaFFwiUJo33fRnW6JOVQwdVB0+GK2lOVE4YFJEbpKO/mwgS
y2pdcHAaByVST4lmQckpK8A4KjfFuUXWW8PwrPQ57LAvfoNMvPglbQzG6nDLTDryNbDiyENF3F/h
nnsnFxEaFw8MnQxN7ihcdnfYUm8WQzzMP5Q+QlnJc8p2lwDi3UuwuOOt4Gr6RNq+r+1DFhDXwaas
vK51N9Fc+9GfwE7bwR24SMbvKZCtItHLwQXZ6qTbAKWx9Tq089xztiTGRXR20n+Esh2lX9uxY973
fpVpscaFF/CISr7WE5JEihgVls4OOCmGLLXJ5+5xiXBmh7lsDHXfZxSn3RQpf+z1m++HmqdwJW8R
D8KOm0fyFHX9Lq2libUrqcImQ91tLbjy/zyhsuZTSZpDnU+Vhu+OSzR9//38+C1bDCn1OaktYjyk
3eDoZIK6gDmIkbV6VCsxfPlwsYktd/zP11COWHhxaNnj+YdqsCqollCeSGf7/8BG9btc4ly+zbxQ
q69zV+Dep7iLrItvhnErPML49efpfF9NfI1CgynAH9TS4zplYJ1UOpXtxtO4qgMHUobu4kezQYlB
ZV9NXSe/TULlaR86i2G2hmlb5yNLOdpKgKcFK7Fjf33kHxpglgrL5CPdtzPyOpBa9y9GmjxaaO0X
QcAojAJiJjMGU43qQmbWyKl0vUt6ljUAq+ntZlwkYGK2h67uliAMk6uflr6xy0VSYbv9B2UD8h0+
Dbb9u+lXdrIYPBoAIyDFWKUMFsnGrr96v9o23bBhj1JHEBQYm5bDTpe4hMDTkUIyYq95uFfXxAVE
et+82MatgvsYi2MqlEf/3pGSQ7qkLSXcFj6CBkixLRW7r4j4i9QfYy0cJM3lwQbuRBeuMfSt53hu
mvEJ+XzvuVxEljFm3dH3LVYdtjPmorapiqiqEJRoTCygpWJi7HV2PwWXct2faNheJa5Xe16M0c/8
T/8ZZt8/tmtxIOjoVbHK7wuXn8x0VuS+8YomOWsrd3FPPtmrHpS/mQyLQQVL2m/Fh9jw+f/R6KOO
Qh0/+XcB7zUse5TDhT3DROP8absyFswNuA7m755DT3jEjpOl8ypCRh8vSWSsq6oZ/WO0joiqqwbl
Gh7G0D7eX+TE0JEN9gdU6FOa9xiWHdjoCx7OdTBx6lDqUlT00yOFopBH0TdD+Xe0Ecammrx/a9V1
t7r4ezkj0KdJkJ3rCWFC8u5F0gNfkHgmxt6TZuLe6+iF2sb8LcmSxxY3LPNaTGFUSx8Pgl6hL6MM
ezpzbXdeFCNsWCs1kzJU6aRhTPiJledRccqfjmdcSMOpZO8zrJddxiiYvDefGCRR2vMUEG8MK62r
5+Li67Fxtvn7TZ7e2qFSE1UBKUpF3AKPq20lWnZp12w2xqn5mMdeJ0HC3DwOVAVF0t/bKbhh3lU6
h7CJ6PtmiLHlulVNc70n7g/cLpMVOcqFjKdsoJQmpE/HiYHG9CnHebsglodQs4xyNx8YcXHQKcCC
RBvaNkfhbcmL+sYJR5o//SUv3lFJfpDt9zeSxesnew+K/U3zFPTNwJHIhpkK8tYHTwRSII8V4AqG
fwX2twsQgzYHiji63pKe3pZCIQJYvITDQ5DCYu5f1T+hH2rX2DmO5F2gIIdX4tnoCKVvj2kbE/Ty
5NLvFshGLM5ngmtVufWS3jdIlmezqvnWlXsV8w2GHIorKfOjm3wUycsgLsS9CtlPNx9bkUZUPzW+
gyRfuxXUuXQ069aPHMgSpqRIiGevQFiFD6n89e1EyLKPYIPOhbtN25dliPfK6szINGddAAPFBAzg
sG3lhhvuDKJzJww1vCN5RpiynQDEY8IFh4QzOxrFsd2wwUQa6A0oefWq5axAQp0vwEjViWftxgai
B2X5pabo0CJc/fyiFjnHVLdd3h1eu5AiUzne94zbfFMTAUfz8c2pOhXFQDO3/ic13hDCJFdEkZzO
u251zhcwT7F04c+0EqUCq7P6e4Hig/x99A/kAEghIQ0cK+Uc79mFSjx8c3b+crc6WeWEtBbkqVzz
wq8/tVdTen4UbKGoC9jb74fGoDKJqfI3cwPz1ZL+1B75AYmggADb2h0b0nFEEWJxF6xM96tkoSf1
V1kbJLS16ekoH9QY8K34XTzhqxwWBaHQLt53jJ5k3xwzdjxNsblOlLjLbnDjG59l49JsgyflUuAl
aTX0AVaMS41MKPWdOmlfuoiXu9p9SEvP8Hrb1Km2OgPcNsV6bjc7TkG5xO5TkCCrbwLqsbNpG+xw
1R5E1kxI0WVhtEAnnPcU+3KAi+zLLHDsFWXd5GqFSXAxNKLx/AcJhVnlrD0EF+xrK0YurIb/VVcY
wKJcWXJSb88gS2738MsyEIb7HfuK29H8aoIKvns81ytQFX6iaTrhuazF6W+7xbWO9n8GXcSZZZai
PPSUNroSfRFRfjKiUm2FDDmll6PrTPYMOAcBfTe0qhR3gg+UxvuodxPEdZeh1Rpo1NaRPxN3b7yh
5J76F0FKk5sllga9cLvGGysbEgQC8LF2gVZxNjqgMHS9B6U1A5/Cpp6lr4ZwUj/XfI1+6vxGKwTA
LMwkPfxnY7DEsqMHMEzrFRoceK8KimkZ2lEpu7EnEdQUEZUPFF6hC35Kw7BgVX/CqBlOii0zWgdw
+o6HlDddrdR35tk2LcwiL7M5ZL+FfQFzmV4EtQobmzRfyOhOOnfBY1cWrx71BwXiRJEw0Ql10e0b
UnRyxCpC23RcJqvFYmMNHJlMDaKxD8OsvLhIuf1COkBsLZqFMsB03BLvtkKzym9SqM0hs9ZlvISL
tJ0d7dRhpnY0XDd6kWtmh/T99ieQzi+QcVLGts1WzOlBCO7OmRDFW1iogMhZMuLnxuOCPCSEi4m7
Wzq8KnLPLePo0+SzERu40NlvHm8KvfiiB3hD195JViZVcrSrrNTBuL82wfcV4vrOwBcpEZy5XsQq
on/8gYBKFA4JJ9qKKHskdK8fEO9tLXyNHxQ+SdAh3cTM2JYImc7O2lhQtD3J/neDiez/8IZGr0+j
dYbvdAk9PESKt8Th8mhHN4Ph6MSHZ+jmsS4SWqmAG0OGZeolHeXueNc34dkVcee7nsNlKVhSb7zc
YPAbEy7c24o71sfMLlzyMQ7j6dXRKCN0Zex00vxWtdjCO1AOVdoICeOeGocbPAFzAtsVDmCEgWsl
eWx6SnVvhbG6Q/WUoWHjuSjSsDUHndyddBYb9j5sFW2bMppOKNEVufV5oMJj0GYzXMFCEDhFkj8L
5B/NEcd99P25AjwYU/2nyjaHvms1bYTRnUpstYsHXSf2+8qV6IgrTy9gs2VhdyWWB6DuobsgCns9
ducW+n2EY0+t0B/x97x/vRBcsGm9/28huFv21W4YrUo2NzOJuqi0G8Jgikyfuw07gFInQhvsFO4R
6zquPw8S/6LkPg/pFTK/fWi5Lvzlthz1MU6WjoQ+la581xyTsAYzVlZhmKPRhoyMuzn9+QYukXG5
NJjXPYDGpeWr6gHoLoKWFh7mr3n8f+uchWTEHJWLpux0ij9wLwUDUndR0Ufw6MqbvN3nUHZFSW3L
NxfavT0W0DR3AaqQJJDUhtTiOCsq0IXR7W9qj7o/ibvVKt07+rgjY4iwsSDOI7cKNvchrxWj6L5I
uEFaOeh7T34r9aVieBLucxcwwxJAG2stksGminhQrLi0vhrMmbgp/DJTaaq9zf52TUtMZbShOPg0
x0V6Ci62lZflJ74rlBdM8Iy2lky1K3VCO0fRprz5KDWOhS03AZHfflA1rDd9SELDCUgUHwmO2Z1R
IRQD80AzRxGkAeukp096dho6Juz7eBf+MThlkDbRKgUs8j4KzQdTSIxvcSklI7pUupAtYJXj+9zT
HwknWvuZgqDkVGtgKYH6iHHm5NM9d26E2tQlOdEpi73h2uQ4T1xO1PpkrAZuroX52X1CwtAJVypT
zsFn7ecxnOCqC4EeXOzmnJpD5QjjWxIsMm7V+xJTgZCwP52AXuxYXGfB60p047YH
`protect end_protected

