------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package my_config_parameters is
  constant common_clk_frequency : real := 200.0; 
end my_config_parameters;
