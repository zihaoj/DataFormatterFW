

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lhQ+XlBeAs0Z5+Vz9RfSdGu5rTRq72Mpeu4VrXh3wDOSCvnLSQluXHrkSmaxr0yX1qCEYyZuct7D
nj02VbE8+w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BpCGJJZWN+A7WTXwNahiAmIH7nSVYW3ycunDTe4fjrLJKhJ0vJXq2ecGIkwMaNg0HXQh5F0nLZ84
ub37+gCs6vlCBgcEpOo55XXp+iaTxZ7QX5nd7u5cUZFWXcTnmXsGOMh8LSxw7cdxvzdXsefEw1tP
bEGGRiId0N2OVAmmWyM=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VZbaR7hQAwVyLf2Yf68/MSeT/U6511x/ijlyKaGJs4rEqh46+JchMDzaLJ3iIBrbZ5EiI5uXruPw
cimIxMyoflspudGxN/rG3qPgEXVoWPtdpS84cTEyGJE3vsnXflhorvq+q/RUq3gf/7jld7ltgF9d
stYzDnzPhtg0iJ7MlwjVGr2VBWF5Q9PN2rbJV6u7Pa4wqc2IuZJ1oCvxEjxuDi4Trc38w6kKe60v
GeFSXqNUeeis4SUWQLAdyoa2D4DVhkdoW2cTozJvsWZ+Dk5lo+qKRDBbPnfVvOVZ5dCugHTWA95f
4Kr0AvOjBlfr68Mw6tJTEVAAihFEspkUlSxYcA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KaMYcm8WxLyssidacMPpfNVr85s13+oGcSsIdhyaOBLinjcNDndRo/t3USIeR/VVhJfAk6UjoiUb
4Zvf56qK2u/XVISirFvhI3nK8wHHZzD9RPS9TJnQ4G3nbPnvdDTJVYzWqF2jejq7+ZIAwD4Ebqg1
HRKkbjP4//IapQ1s3XY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kwozcJxFGUF1vRYNYWvOBbLr3TZbdDF4ODupv9Oy0ncJwWY4wNMydb4i3KeBhJd5CSTGgBmxpEUU
sf6muW+F4torQqHH8YS0oeEzr69zcsKl7f6DTLaW0x5FQcAEtreGLwK8Hhfa1p2OeYn9/aR4hj4L
QQfLl+9LadlzelUfchHoSTsC2RkpDkvyNfa0Q6BQjLEI7hJO8x5Vfi/OWcYki2jOUY0D/qA1wpPT
VSsbs9N3ODQb31cNrMkhOxImhK9/b1txt+7SsBsOWZIt15aQa3YdrUWWonDbX6BhVvIEZgec0v+i
adelZvOaI4d4vyz+3C53hfGPja/4CoyRv8qw/Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 157312)
`protect data_block
BP7Ym1Az381rFnFQNSBAu1Jqav72bH0Do/6bQ0fmDuwbMg6sj8XP4XQvfMQai3YlTk03emCvaWsg
mJ31PfaPHrCLqZnQU549N0CIQTZWM8c9qM2Uuc+9qcFYwjEqYlEV31jqV+DTBHrZMf1NHOdr76XV
89Os75E09MLQvIa4xT/av6JLiUDuW+y8rvCtohMlZkaTBP3L7Kn00TXugcROcYk9/SEtIDWhYgjm
Hd3cGnbEqM2kWVoSMTwKK/Q2XPKuJvI8u16SfGYgOsZ+tHpo8uGRWcZoc6qWHmDJMb87RZqRqsWi
wQIEQ9ImMXUK1FXUJszvXqWRM/sDCYn/xUtvk1DBz+HfIKn9jVpBZdVr7xtGVTq3r/b5+UxI6rTp
3zJbN4e6YPdnvADKjggU1C2owORpxnB+27k6DRUx45libkIYISgRI0hk3MlhwJtQa8B0iQdVS/w3
qx78cu1K27KLPdrUjt/w9CaKaSKDWUEofueyoXzARzn786tTaDYoTCMIjV6aJDGmetOvcKhkqF4y
7+Ir7WKi7vOpvxpIC9Ca9yI5kg4HVXEk93YeZ7G1/tGwmT3Z2P/hwmACfDL7EARhkEmd3kvNzX1c
gP8Td6CJkH9RewoMZx3yYkETfzlCmWVLfD1CfNuLrqYrY0vsCw/zKBRzlJfnnqLCJPg8JXUYdE76
gM9QJzhpYyY6iBXBOPkl0S1u2BrG+P97jdrZ9OTy2aarRlx5/yHLvDHeXfz1EhxwuCd5ma9DPJQE
18o90LHZacDgi9DO9uRcWGZ8++LNBPSnth9VM39RME367enRkM8lfxh2uDPDpgBQVyFSFGO9PaKF
nNKJXULun/Ws/Vm3fLRa30SfIUsfCxnF4ucYGsJ1z+tC8mkESzhBwr6DrdjTPXns/61TAcIFDXS3
vNYhfTyOw8wDU2jSsVoWve/3xD9U232XUWl15X9l+oi6TEdjQij65pn9jc51ui/yZF5uiJ0rb3wy
faVoSo0KtUpi0opP8NETNMbKjSWHpIZxNk0500nFcy3Vq1MMnc0TpEC0XF4FjTxKRwIFvAWiBNwE
05nJXmwk6tRvvJUnYgfWd7aOQaI+UxRKDKluA6xH2j/O4FqE+ztAw/ZYfAPv2p+QlwSbXf0+pbWj
Mw9rkTrDNO/LEk35MY8MwrETqAswhzXt+4lcUIZk64QhttVWBC4bYd6xF7HpO+NwLf+WcOL2gDs0
8X70c2OJ93KVKFdfwVenlyUyUMCaSdYmp3zHcS6rpIEaDSlLc6vpcbVrLaOnARcjwNCBdyGsaSuj
veFO1vqtCK5gPayAzCPPSH2XSx8187vjQO/WNUB7rJAnzqDwUNYeAEldUDj3kI5b6s2XIdReGYkA
0qlhcmB7Azo5ogKlHS/hS8tIPdQ1IN7v8PftKv2Ytc8c+0GHyJgaQRo4GvPVFnOHY55LE+5beqHN
rAzGUZdP/ZC4Y1iRPjVY1KP8cJqeEPZk+BJIBOHC+Z6ExJxlwUeWpjKBVoCpZn780EbSiqN5h46n
vxuSgZW096+EMWjQxPeJ3O93OYMJGYooMhCYPMybBgdszVWMxJGP0hR8UTnCuK0CsHa+NA7gA3th
JKuhD7+TUaDi1S8XyTWW5kdl/Im4OCcsF2/Gz1N2zV4OyAlRkhpDdWRAHvuBEn2R2VQ2hjIXw0LP
9tSdK6XSD6fecJixwacou6UnFxV5PNskDwGXasLpNjIBs8GZn2y18mSnlipg6p5JlsMoS4IKAYHX
iaN4l0ofde6b9Npnue0Px01UK6xLqfXm+QmteyDVdjl/ai/tsptXckeBNgvIfJ3TaxG7m+3htW3Z
0UAFlQAGYxGFTytWeLU7/OQ5DI+koBDkpMuiLlVbAFUBTqbB+qJBC6UDnzisv6q7r2SKxl9P35j9
ETGQRx6AOVVZc0aJDE0DAWusjeGZa5spGfJlEW23Y2yMvjPrL6Hlz/qIAbsEyrFbIGx1G+P5jUHY
9D7FE6AXWlNC2ILimk6vI1opOd8uiOG5YjQjiql8R5LvdkTvCbO3MZto/RPNV5wa84i9nTyw9CZj
IDbG78khFQ34dpXlepQAXKRBdjs5ILBQRZFYGexjD3Ak+ioX5A55nfwDSksUa3gxR85aU5d4iI4W
/D6xIBd7fZKGVullxsLXHMJCcX5FcY6EB+4WssMUOeGnjGLo7nzt8hkBruQn31vzDbt8kdr/qo6d
TVOEOm9DJ2gBgwbKtyluxlzxqpyKx7Jq+1hW09b5R3z1wtf+0wZr2z9aq6nKVFAhl45D5Az9anlu
oiZI4LDO4d7VL3znrBBEU5PjgKGS2ntBOwK7g+evWsI0uHoKzYhjLpiZnEB4YIwOhdRHWodQdeqP
l5wENChAR5FDhD/lrHmwFi+UPihHHyHCGTGUTgRvReLsUMWs3mkvd+VgdiwWRwDfUuqhTF7Y4bRI
tgspGEQcZsZj/vR+54ZkgFSR0ecmgB3oGA0U4ZvIURL+8bxzrF18XO6Fkf5YxfulRCqKFnHHmk1X
sE7qWc10MBvwGCKxGk8r21rQospr6okpc60l/9BjyQyCsGw61grDwkFISMXoHDXm70K2R7Fzygqy
fEVfZXpmt2s+73EsKhMeOjd+7YNZRTl9Yk6lFRnKv3CgA2pn9j2LU8St68I8Du3ksiVUURqczfFo
QdNHRYdIDtvf0XtAwGEl9M7RwMw6urtv8TLLAB/Yv0vqXSYz2ZHoJzuFWNw+7yBMwdFG2N2/m07s
6pf9H2dDfhWw4T5m27pH7d3l0LUP8MVcCF58IqdvIIFCMDMAgwICKAiOtNEFK7SMDv593VxOW+7x
O7GirOr01d2xxkaqjbSJM9kN00mp+mkxsmq6Fe4DTA7eyw6uuEwBb5gr7xm11DsVWPn2kabFlhC7
tEoMGpRy5Jz+ZEfwCFvTM/EKbWn3a5zSealnC/B9XCBG/NFUSNJW92MKY6JGNJhjUkRJaW+M3yR9
LmSztS2L+4vsAwNU4VT0TGqYbrO3PaHpPcKkG6BwVURWvNsoBFAllm6KYj1zHTVvES6EoaE3oOsd
ZWSfnOc891gWkcuXveJoe5jyahasqXUyDtj9YuGA3MKaPpiZ28PaWpk3QNd1ssTcbBv/5+l35BW/
5gez9cLOlhdCxE+uTrtNKeMfBKgYTZGKcMaVnaBFHeGfjQlHoV0codTRJQVefzqoqD/hZrY2si1i
ZR7bxdfuLKtx9mWLHHUxvfsnzMeq47D509R9ctY/oSxRYVqLn229hzeHmf2WkC7KhPZDb/Y5QB3F
bXRxe3S1UG5R49P970kl6r7oZPxmgS6AFMRFE4vprpu4hBVmcJDQ1Na72aGTiaM/MlzH6AnRW6h1
SADc2Dg9zJbzeReu3CCTbVZ8QqLJQnc/lAKzWZUilAY5IvkOorsP5l9IOROC/ixIolFZJlppLFOF
8k47Q2gIC/ViCeDVp6NkuWcGYPUNA3WWsIZ1Y1mu1lGk6NyfI4AZqf85Z5c0T2QXmFJXSC4EE8ds
RFtIBM8jXUVuLVpQFbmq9slwaKCw1dUqDSj0qHxrzVmeE1iO4ZG6UqEYIIyXuTx4vI3hixv+tTKT
gst0s+P4JUzfF4C+EJ2vA81ZciGlsIyQ8uPcYN5sxu18/CIHR1j+LXwYoeb0OorYQtecouVU3+DK
FbJDRLrR5tieSmQPvmHqt27K0UxCrqxedAQfQnV6zZaDwnPlTcehBFpzK9N5T6IEFRoY7ckoEgL/
CjhjPzCDZfq7qyPhbtsog40cKhb5owA46a7k5AaJl+Dl8KUdyr6lpRCo0Ticer3QL+/M6+JfEE2X
NCUmUXbOqrhkZojWJmIDFrXst5kgPd2hFB/89ej6gIK93mFMZ0+NkTuc7YCO1byUm9Zru8ZDq4Zp
SB7ezGz5OzXQqDkIrTthV4CjAaPPXCi8HjtvYrTU6Rx7Y18HUU8aTBe0fSP6JLP0Ztt7tV3aeICf
5nTQT3iu61Xl94a0E09bdycJ+VoK+KCe1ba1y+utZkpy6uuvSFfP4Q4OxTnicXQtXj4V6UpZSwKK
23spjEWC4/PcvH6gdqniDyStQUa/CKc0nW6daIzX+XrWhRdiwv9ZV5MLNiO0eoRbae6uN+XWSyRv
brNQXSdChXPabTzNhYFkENJsWSpHJqE1w5EdytDjKLmJ1ow9LKpXiO49RtecNYftiTsR/a8aKg5N
bpVry8Dps3SQs+WOI6iZ5yfEZjD8zggt+Zg7YJTo4vKJK7rgNAXkxMyihI9nz56EutrrW5zyUdte
MYiiddOSWXBVumEBjE37oGjJYb7HVomtDrcQDFjRz0pptuXLTXq6uFeKaP+0Dmj4lcgpIbiahPef
9VsqMifxjz8tIYflyRErPlxfr1VApYTVWCqt1CpA97hiV5kV/Gu047jJmyY+QP6sYTp4rkiymQR5
t8iJrcA102qf2Ud7Fejw9Lb4T0km3PmTMwjirf0yTO5GWyL8VdOw4sAuLgi2/wi9JehSwYgUVmiN
laaRWy4a4vL12jPHGVwACWMAMfAmqp8H/0ziVd3ZmaRO72tOVSO0u8/9mMAEDfDUvFJWVv6tLeiN
gqpeERCMem2GkZBCWmayaYdLXt0UWEvh7UUjKbzVMi2+EaZoj6eZJf21BJLow6i3cKHIlZ/Sdc2K
4lRhgqnOnNMVb9A90vNFMXd7jMjXMlkvoVn1d4xSV5cvavYJdjFVNlxvqN0Om3GV12MRdzKzRZ4K
qzRVVrHb8BdF2O3N+J0ugaD37e4cIMvdWaC0epCirpxC3FL2Yw/25d9s05JqeoyWSnSymuLM95wi
n53EHE/UGRIycQVStm1pCPdv9OgcfZO84M2FgPQcyBHoeE8ZHWZhwC7xgCagVKzbW3J8l+qQX5Xj
VpqYpTSBXVOoovEZtqni86sXv7QPBYe/bxsVT7GKMOhIZc9j6DGpa5D+EA+Lstc/KdEApW/Irok6
v/1Q9OXs+R56wZV/jBtLKGBLylu9xho2oDwijjIVZh2HLB4XjlZslpfJs0dIkAG7x+FkbaS7URK7
Xlf17cqUIBTF3oxl0QMNlqPbPDyG7yrxxQTEBNSHO9+eB32gNekCp1QlexTpUyEDri4hDzru0dr0
KMzltxD31tMdl7xbNvCmJtZ6LbrxnVTKqJFhsjFBa67fHlEq8Kp/mAD1cHOpIPtidM5tTQG1aMzB
PPlQXWTv+BbheglosASzd9lZym7V0rU5FkMURtX8mCIICMt+ds+0uRjt/acOXoiXvqRP0ZAOsMwj
QtJyooLzgFled4LD0+b6aY0BaKJsNwkpQk68li/EicfQbsovPewWxSLfWdZ9w1PpjIp/+x8P6UlP
cPcz2iUpk0uTcxuyp/+TC40896i47f7gtqmklJst4AHNQHgjaITADAPm54wwBjegQieB4ncr5H3s
2UJByUF20Wm8DPLS0cwN3uSoun8CI+OOeTgjo3d2xorRjOLviOTS4av0QKd3fDH5tQklwDuDxHyw
UN0k6orwCGGJDwmjGcM7aeBNHX+8rQf6T1jTulBVF3CJsk32y5gqPG+CHb+OXLoIWER5Ni32B3yR
QZkYM/ns4lX95UKLM/zfgpBTimfc8QrhtzkA+BYhnODXwpDZBnQo2fJoX/Y3IRPZO872KPBCE+iy
Va5l0uNSeBgD0eOoWxBGqag1DvQK0H9oiuG1h/ZUJPRluS7NREf29HMzp7mc8TjqUFOKDi+0OJAb
lldNCWSI18iEoyXeTPfk91HcxJhtStSPl2Eo6egT18uX67Q1rYzB69lg/dx3qqg4z9v3ts+yzlfw
ZBdnyVw7F+BQhtCAfG4BjxCKO/WF3wycQa2RXVXRSP/PWEcp9f/QPMS6l7wl9FZRH1Kd4oht8KxV
5h2XV5HXibFAaYcKzjC33O1WZIcjfuOkNjibOXq/qM602nHuXFUNNNYXue0BF8eDX9JTgRyFET5I
7/3OLy9lildh/1ABSjvV93fHdDVKX61gV7VhyBH5+pBRS4XFmZ56jypwTYDjAkpHr0xUO6tAbGlY
jWUlcbyqu8ksBVS+hHzH7YH9YeHz+qM2ZUJ/GRo3QTEGuLHbPjEIuagDY7g2kGJWc6MEDfHHcBj7
6QDULYlAG890OEBV4SIJ5pPZ9GO8OLqjtBX/j0MqwLiKzAijqAaN57XLWeEcduF41D5xoPXpHumB
nSDFQcVo8XoL9hRw2HqdpTKcl+TBbBS8NDqP4b8rEkVLBVpKFaz6KBNW87q13KbUyFx4dML14+hl
LtqBF9L0puoVYtQMzxbkixn20IOdxtVPN7mDrHxO1JW7sqYzLK59HSbqltY1oANB66595jQQ9YL0
ua84mw0YtPuDHhfD6XGXtZzED7DKQPsHQQwe6JE6Hl0sabyIAyvdx2x3lhuMi7syCjKczv23uS85
Nty4/2EbKw6Dp6rlxtrxGmM3lCGcbI2xxTbxTRjepzjOB94bQLvzeprrjxALc4fN0Iu0IlVYohLR
IV8CUUvwLSLjq2Okc4zQhYOgQIxkt2EWfUo//GYb/zMhDKB96Djz1sHBUxHnOKxUhzDEA/8dcPpe
gYAYpWh4D5OrIAVrU0d29d9qpgdjX5RPHHlcmXCsDNDbmy5ixdTXNYZ+5Sl5347ciVugTATWQWOw
eTyt1DHa30qZYK9v7UHXwFMZfAh093LgS3Yan2OuUG5tbDOmId9kIGMXmpLugaAtQWVLG1t9ySr5
ym2EuRCVArNKRTXBtjtAnUmoseYbZ5fW1KsenRzcpQfp/d6UQglmJolmlr8OO09OrcI9Y/FlLfc1
67jbm3KZLiOdcoWydhByqIFQ/1M10PZnX4BFKCdbaLDSrqfMzeEye7iZRCT+5qYC6YUD8cyx2Sw3
pyZlhk4SzhBvf0j62kHTPX+olWD5K9ofLsNwESZG2q/wWvrbdeaBcLMcye0CevLtzZdjGNRc9zkI
1n8p4OoTU4khz2VIZXeJOj9BI0HY67xjrmi/56Dp1goAnT5vYBMZi4uJ3aUHuNBF7NzwDjxzutTL
z5+CiFu60Cp+4U22Autz/Xi2f4shnagdsgTAJsV1F8wsm4Fh5Si9jHr4Rlm2elEUf5u/kNv2UzKl
1QVOh4Tsd85Br4zkxsZLg4pDk4vd0e0AesBIdZoXDn1Oy+gSDthJJ0CHpqnHiarr7ukdHJensUxq
pLLrVrJJdGYzIpmGWIrXbhI7TKEGqYnGQ+RY8W6jNxJ506rBkt2+NLVGR/ac0ugoOL8YUe5oSdC0
3phw+5nbj0xDWxejAeKIfcw7UP8HxHaDuPR+6CyI2Dw2umrAoHV0zMA/vDfzigaxRptCiAotOXzK
uUdpG7DQi2mxGEP8DR29QKfJNqVtUqQiU3EmZTYI2+cMp1xgxfTCu1ruKxJ6NFqIcNODsg5ocBpL
flTOdvRqVCc0bs4UbX2tpDKR7JMN7zdt+/PHmDolBiIe4MfHsUXPpS2iwCKqMY1H/gbG2igA+9PR
LCP211lh+pg+ezwuPvS/SQR8jyphA4hBuHFqqY6LuSt09+2yoESeQw/a+yk/FBABbf+dkAA9L3pn
tGPm5ArPJW64rdNsty43Q7Y5/1k10owdVgyuOMokjgVIES7pLGq/Xas8R3NuIeUzJXHPyO3rs+HL
y6LkZj4PtLB4aMgZsHIdE/gU4+OSifcsrBBF7a7gd1ApmM4E1WXek8xl8RikdNAC8OP555m38gDt
neBnyebieVttghKktyhNHL6vLRETG3Y+B5APcHYdki33QpYYjHCcHT/6Fi9maFel0pPzZQeaQQXw
rSIZxa6vIGwyu3AV/3CSUkFatbOYbilrJPpekp9wlYuKbl92b+XFiqAlpHndrgkA7ddihddurFoE
7SI3taU383AxNr1r8/y87PjThHLBV9J5i6g5zz9ImUrTr2q7G3SZzs9/oK/9sii6//KR1OoVnJDe
E+tZ1K8tqLBD/VIgwxVd6vv5zKNqcg8KEW1uyI1gO8/AO/sQWsPwh0JQYpwUolP5GWUCcD3OrFBq
WR2efhFMwQ3XNcO/DDLsqJ3k3b9JSz6aTPNYd49A/ZZ+5Bqm/m3A7tzM6Gt9VMGCOkNy81apnvuw
Zudb1QHtm39kCvh4Qjt08R03PctTNO811AT92i4k7vADYuUQfyA7V5kYxDGYf0MYPLwKDyXSsC4i
hjt/YrCI+aDgxiPYSqGwehgXq3IgxKsy+hUGOjJ2lrn43HScATOKHacC4U8jCvBgCCG1+rFTdYd/
TLlV4dvN+r/3ll0EOW/vgvk21U/y9ORvy/Tnmb7zusyqN+EkY0mZXgrfEkFF9OhdAG/GSXyxFTS8
Dk23PDsDjtzAWSUAJBc0I0ZQsYSgQad65k9wCvSvq9tSi/aYdl4EIFX6CTHakrZ/jnfQL67kYFyI
9rg8sBnHi0JFsCXxTDiM/1/Phg/6YRFkD/PofbLfakewS44a8FtK24oh0I1PBZ7KAjBJVzMgQCPv
DsvE1VpybHO2ZfwvwmeUPKhGBXN3MCQH1xeZUVRkG0ySbDd+CPeAXdPzro320+qyYfrmyAI/QGSe
H6oEvBKB3aKmjiuwmXFQUrsSCgdVAajqHi9PZ2qHjZo5Jk3+qDmALIvDC6EhhUvF9LUMA8Uh7hif
2BEoDdHoGmWXmiPGuTW34F0t4HO8hLGuqP/Im1RizbLrOox52lfYoU1fLmN1aHV3Cyf7nCOgjH+T
YzlNlc6N2CkBGxFZbNkOvC16gXq4TGZFcEzfG46ffb7XH2dZBgXoCWK/IEpH51k1935Eh3eyGx/J
n8pNbAJZJWLHgx/g3gkU61+EsvJo1UEkDx9ZX2xwp9rC3szALiu1snfz2yInWxLaOwRYwoBN+pqj
RAD/bNDJAjb1IjAqkwuNg9n3KiRbXoAhRUaDeljpzdLznfBEkxjs9B2P9dKW/5xAmTxUoL2+CBic
xv5UgYmtvWHL3ZwEXUXciyBOkQOU0kAaUKclX3SPgWmVPHhEjNLPPaa91pbrWWPGttu8IMY6AeZF
2bjL3q/xTTUbFaym9K9hznjmtgag+494MMnvyp4mh/Q/j0Jbt8EacC1eC1mx6fhhfrC/TBkVW09m
GzvpvQXQY/fWnRdsUlkOvxipnVND/vae964kAdUEvO1u8S2r4VJbOhgsuvsgRZhiqcNWo6EH2zdB
wRudAWLJI5Xw1sZNDis0XcPVWwQkh4q3zO8Rhdy3nxFcJnMVIQVb23Z6DAUz84dg0EtqV5r6KG0W
h68rH2r1h/mgOcttYJEry6DrPoxvj40nYDfuE/HLrpCFt4IJKTvEWPop616wBr9WzbW5iaxVCdF/
Op4KwSHr8qOuQtgzKdDw5Xq1d1O52r5NI4NkFh1CHdQR9TJqZKyxXa/C7gAut3GlfbgRS+tgMgle
thfsBSlSmM3GRfBTl/epZcX0vpwGe4wMFFI+LCSmEIOxfXBycuAGYMtTUBzz+BcjCuF/AZDlC1Wr
YJ7isuGbiy+WrUlpFoPDOvVxJhmalCS8dNpu+KU2UbQq+mhEXBV9rqGA7dA626IrZlrlFbB4mvoc
EBvZt7L8yWM+S3Pzx6eX2h9FHhyNospw79HIFXySq8MTMbCWlVznkk2Hv9M1jcCLoeVgjt4KCgfd
A6clzFQBcl7Y2mBhJ1gAeUJVVjuHYBsMhkIW7PS2VIgX0LI223zA8k//Zn52zV0mEflxnHl+AOgS
GmO58KZ+L8+A2fZerhsHDaXci9vercTL1IsLcXlQBit39m0WwVCM0rm6TVtgHk1r49P8dsX4vVhb
zeoEjPQPbqiHhHCe65uUTymoShLVkks/jJWQfA5JDSgioIZ5F5gWbbFXEvWtsTJqfLXy7sbe7zo5
FXbNLpyauJf9nElnzqWHXIAwoyJUeOg3NMKonBjJVEvjaY3XQuVkczPdi+5AlIe73AKkBbrMPTur
Ohbyz2PuD0F6NDNmxex0XPN/eYK05X24J3zc1+7iHwMDkSjg4Cg1A/g6LunS/Fic3/xjO4ywSCmt
I68VgFUut6j77Ff2u38P9YO31g6swuohMPpyIGR6YVlAmzwwSocVfbuojB0XhUGg42guo+egRKAz
No3lk4VPC9hTVG40p77hqpwmnx90ctQn3UNorjUenOaGAPMnWVvVM94f73icvKuKBt5ojFv+hnXo
JZFRv0VblirPXd0KtaUACbiuE+FcHUuO39h8VRxbvAcPXTdkEzDES+bKhParYKOsKl8m8gvKK6jX
VZxsvy49GL+AzH0FqXsLPCPMokBe4leVj9VWPju0ku71DkyzQuDZyXhWj2UM7G4AYW/YUckkkkuo
JwZA7qbRGBZ3HGRJH13hlcQI/Yba7Y+/MKZLBW8BpOCVWrHK6m91fwIimk714USYuAUUKgtG1HZl
/5wyqWzgz4P5BF9f4mH3EirThEHalKGW+2mlfOewAx124awtL7ykY7p+9H5b2TDaPhpfuMzfhNNG
rLxT3wLNuq983ByuVpEMLj/WiBauUNPbJZcfFa3D8QnXTB1wba75ZlzETKuu/odJ2Q3wFsxh65v7
yBDqtG+qQi3xV8BLjB5m1KCD6F2UDOY0iFVEslrC1jX0Rc5yuQMmq1UZmqPOH0D1Z6mroPNvnTwU
C39qXB2ltKbskdoaxpPzJePQO3eqd5VnwYRzZNXjetLW4LrQjDWQhw7J7eMb5Hla0ye7b+6hlUOe
ht5GsOYd9NeGkIsCpDtiVoQRyFlMKcUF4uZbeZySiHihVEesxfRFpFmm3mMi89/myAmKPQuqA33B
quU/SZiZAWlcouI7ICGTQRly3L9IORRE6NgHGpiHNkHU47I1C4Dp4oI9QNA2w/RkkUx1GYSQdfV4
7Pz1bFdeKkHPsqX56eUAMvbyg9XKCV5WQ/oELH2jD0Q1ZIRxaIN3a3xnemmAg6fljehUQobV6GmT
n2Ra7oLQcJa0NJNdCQvkgyHfS+H7o5kMepPjo0zfPqNfWParZaklkSuTQb+mMejmCNhHYyfFahpf
n8Hox0Nz2mQJ2KZFPUkwddzz+wb9zsNtowlKD/WkjyFmYA6zN+OkCO1Va4TXBldfvSCPhPct3D0J
AmaCo4nfaTjRLDOcigm8ku/t0GJodxf+eqXoCkA0E1wTjpwagvS8mlDeCEAY9FJVcB20go/7nAOB
x9TPkwV8aPUYPqH5lXmTX/Sts/aFpxhFomglf7mW+F+FqVDoc8kgkmPEhvQKyeMFvpghfNr7UA/O
sFqc2JHkQcsrYILpHAcuwzVFprYomoIEp/CnB3gwRDLlxsNAz8goJBv5g2UtcLWlhfde05H6ui1A
93cFMh1K3OoKvVEQGlxq5+UIuJSSe93OkniN9OpG2Fhoqxoj19PmK8uz1L5olBie3CDO6mZk1lc1
/uTbLTfClvYl8CqhdQaUmKew5i7ApiO9KiOE4JwudOKw9Jfn9oaD5d2IIeIvv7W+gCm9wCbDAO8/
W7M107U2QpUtIi60mcwqqb8dZeTO/511QPqyrmBYIKh7XRoM7cLtKNX4bLKt8fci0vEIgAKjIVX4
D+4QeuUvTkewpyXZ7VafAyDf8+3thtmuh/9wHng6SMGexFhBjKhG7oB5127zjMchN/GMeL8zpLlG
hJo/TRWuWg/TdP2/8pkqcgp9hGj3sKU8FjvBIwE4jfTlimUnuG8DUn0ZDpWulNOd25ed+TVGaA/h
BkfQrZSwbG4x6I5xNVocF8PcGH55cEPkadZC7E9n5nsGFFXlEiVjgq5sAmnU+6ZRFXxR1EG6NQW+
BaYge159yLdLjc0goQuNFVCZUWCtXcKMUDa0LE7VUrJ9ZNNUwkoLMup/JO7C2hlPz5BCRZwl2cFC
ai+T8dgUqzmflbZ8ZCG3zTs41wX+JXfq2hawOADwcbtGTbMJeX3qwCfe+7Dvj8O7FPXQ3rf665kp
LqhFRXhNpOGpWrInpiW46p30eZmZHuTtw7KkGtN6XFdvlypLVdqT78cMdv5Bzl4sBDHxW3Jzia/E
+FUTF4vShsQq+0vH4NW8b1nu7W6JyGYadf8nFXKKPUlm5kMJAQ5ffhg/B+Mcy1+3T2k1ijUhcYpx
KtvoNVxMrXkCgG2Q89ri2zCd5aosFeIlB+CeH5g8WuWOdwaEbSnWVMIErdqlOfPJvn44Eh38/3/V
vlV+XdO2tWt2EpkVHx52KUtEzuvcZlTAqZJxnlThAVOJMIowx/Zkim4vRYYmfEW2Z/t8/TaVzPCm
bhbY3Acew61pCTHuWjaz/USQaIyRf/QYJwMgyQGqVhYon8+RlC1o6DDpKq5EbdlDhSS3TPyj06Wj
Vpvam+dc1dgc4lbAum6q+/+yWOyU5gTlxW8vveUvjT9M6w12YsfNF/yqL4J31PxxPCs0FjMU8x+D
RJKL1Cc1/yYMN7+Ctp2GKhsgAthMY3z5uXaae39OYRfT5CqYy0znpvjKVeecRz1x5+UyGQSFZYly
aSa1YxJTTu/A70aT21B7i5S72Ygfbh0E73kCiNuJiL5nxWL3PcjMLr5S9iravDYxbFJQfNK+iRw0
Wg5cONqDuRKJzyo6Ncj4oMA/FmsEP0gyOJU6VMFd4a4yHtUNdyrOhWUmFhfdjSza67ngJvvyiawV
yxnOtm/8s41n0Kr1GNNSifB6OBQoUuLQOWhAy83PFpfyXPAF7peDSTGXE7LPT1X3iHvd5ja4A5SL
dtEZyWJRcQBb2BOLPBMsxlinFehW7z8byGU6AfXZYeH1ypgx7dWQI5rDZlfy5DCqo00tFrgWCjoo
xygFaAaDo6ztbYRwHpqIZgBi+NZV7+epEN1PIAs77E66PNn5XtQ+SiPbI7iZH9AENRzE/WuTbUvv
vLTf+yfjvRITYcZJugF+rZqyjFrkY9DpyTFtydtgQ5xB7DpE8mSoZ8F4Sj8BLyp/5I4zEp//xfBX
PpcCOI576fPKox5Ax2cM7RTkhNJHw7EvVBltCDkjIQ1ImsoOSuQzrmoftbKsqT95yfAXecLNQGdS
u/gI93Ru+ufCawz8TmdfH39m5WMicLHaa4jrJOPhUtJJsFSVSzAxvit61SuqwoePi0mDgn9i5h3H
oLG6OpVHM/BXfuBLMDvrXqdbfqOr4Nwga+0dGFKO6klOQWKPyW/FJGZKDx9vhV6yc5ODJNwBZcA9
tun1VF/L0VA98p1ODjQpR0s0HjDILKzGEQ0HTvUzXlllxCKQa9CzXZXSq3HYU1nWevQ5j3wB4PyT
FHjGtSKLjUNGjRpyvZbSYrBvEMA4tIehtjEc9henDYKp95Xmf5zFlRppPrPEC7j+WS96PMumAnmH
BteBvdLUmKdQH0qksc2DrBXFvXdeSGmEjS/wwk2Ap6uywyscChxYS1s8ffpxmRsu9baCe6bgfeFX
S9kcT9Ie8C7EZn5nkezYCX7YB1NHiD9KhWtX+cXXGBc7v6tSS2GJWKfsH+uiZd+a8BuVfrXHotR/
IdEtSDkhIg6AKIux0FlSsRDszGsEExt3NquzmAI5x5LsyblBo/rdvewAUI5mCpz66CedyWIV0qPk
ycrVN3kRgTsMAO9B6vw5VzKUIFKaJa9I8lD5YRuoWgvrLtphKycwyGbEsORw1+xySI+AY8chkroW
oAnSxMN4NmM6XjUmts91hIEwgBuoq19RcXPtD+x7d7+Nzt0Plp8jyB6MIeQQT4VoKnuzjBc7ihYm
IesnZLaoQSFIEYFVmGYjqwuURqi2DFy5updd2X7vByl0IkjVkGuuX3sNbtbHidUDDM+781PXb/+O
cIFFGH20k6CBflDxo31vMZVEW9msoDZG3MBp0Jd4WTzg7AmEfVC7OO75PxNpV4vRRtMYc0K4uWee
9Hr8+1AQpsf6VU75k2hBV64kZ1NrmaLpF31qADoqBaoBkIgQLNLUhqeWD/wIAMeD4Z/lvbEWqU6w
nRuoovdGXV6URkWf0jPg7MtqQJxrY9kjNV17QyEU2/nD+YUgKr8v8Vv5/gi21r7SUsvL2waIm2lR
7CZxLMnaS9nhxAmwVBHY/fRr7HrvMIVZ7per/lMUJhisNYLB21MzhYUyiKX/UQY2FFxKNORTVV8C
jhXmZysDK8b1wAfUPjnkD4hQlFBBdNXhVXergtTHgThID6cPMsCtqQU2qM61V7uX8iPTofhbCPlb
OXodCL2Q9ZhcU99ZRpwI/LXUNDNESX4Bn+/hIrCMkper/T5F+Xbp18pgjf9/Jbxfvp4ZITzjvVu0
m/btYHg0bXUA7aOzj0nC2mKqPkcC7wIe5/3nvvQhzrfVMTrWJew6ftWECq8V3e5g2kNIC0aH72KX
14w/BRr5cUlSm6moCAELKRvQp5uiEKUxyM4To0azzCnGOtFnsvVpK7pyckIJvEz07l2jEaedQOpg
ROuPSCGO0+xgmMTB8knjFL9Gla54IPt9TpKjNKgEqbu3vCLQ2YpHfgwwwqDBWzhPnqcCzEKCodN1
vCLk42v50G7dHRGczvTJZvU66sw1v0riWQsG4TM9QgHnAeDtHhAntq1G1npqMPi6QmVyBkajqF0o
MPC8agXoVR5VvrN8EaKXIUuvbe6vL18DAM9/jcA16PeToBaaRRPffmY6c1FhrCmvc6zd8z6mAxkz
GBg7ln7eSqeLjZvHV/2fDwU/h1PhqbcLYarqEq6Tu9hV0xZHay//4TwlqtrBcjbAFcKQVR6QAF0V
mru7MpraNUAL2TnE+npmylt7GKq6vphrW//yo04l/67WZbdToOqkQM54bILHPHOVBKxUWH9pWWG5
4A98trwrCczaMCok4xOZKzIYbVASRzGzb30W5Tl/OWfOdWDjFb/zZJAVfIu9bgba0v1rIZj0bNVS
B9M0pVjJ3plI39NYokGV+X+NSiUtpZuPERsaoJyBSPXxJ6N8GWZi7p3nfNUwA1Q3aCnFWDmyUPQG
rd2jSxf1fzwnCLhGHdPrVTiqaI4oIXa0qe7f/yjrQIhLqZ/LpQwJNi17kIXWxq9ZwcbLxw/ICYH6
ZID8dyjUXqlSpsE8H9ivR82MH+eS8/5sPIuZqU5vRWrHyT3Urtpn7lGBh+tFVTpRU6TCYTzhbUtp
CPN4w+cuMvbtg0TGnKpyVxmkq/ooNcFS0wUJI8ru3GNeNU5x+dGyxHFVrfYHH5xASDjpe/E7Kogx
aN2xsII8KuzFd+kVdmS3PyaWBcfLQejdMyN4cxZKdOwIeGefAvRa17OEyjeZ2BiLK6bi1gExAn62
FFQQr+h7/zXWPguIVZULZSW6JyxbXguHf16oBe8eNAgWFI7OvMRul+KDYQhHEYQJxfOyY0DKnPf8
dnd9K7sinGK3Qfsi0TSA+a/AlsfTYYcR4QYLHKRzTlo5AJNw8geOOnNF17vZkwMLEWDaYc7PHl9U
sNpiDmukP3t+I02MTr8tOC3P6dpl0FLVG2m0yrE6V302cvTU1FAsOGL7WderVvBpwXczPz3aAJrq
XPB5dhlAx87x+2EWzU3nPPP6hNpNruLzu6ieneCzQqDU6hvsifpwXNm9KRYHsHyFr/PimiqK1aHM
j/6WTcKDpbJFmZedmHtKk+5J5J/s4EBwulXxrNrCgjHf8p7mnWenhAApSJI2MNoXAdtfOH7YtgAp
m8l5jB9oJ/i/A4w3UTDQJHiuAHwx6sndNOcYXwz9We/OVthrY2qYipWpn5HS9WnTDNtC1Droy3FR
s6tWu10azh1MuYUgx+eyQ3jGMlIqiFyAG8XgDOj+qQZ3/geDDioryK7TQbDm4eC3EFwH7T/7gOZu
6rNFzP3+HzFKtMr9iBGAzVNA6u4KB1eGdEWZ1SevJ500CXRdxcrWNn87dAccd5ZRgyFY4If/SRME
waH0fsUVkJV4jT31X7Msl9zca0Nqq0apdaraWQWt5OvSk/+1eGKJGJks3np1S/bhWbtC/RC8b/8u
U1uOUE/MP6mUSvhhMcVtTNSQHL7tYix+KzgtFWsiiYEneHsgsYAt+FfJQHHX6LvbdSdJeVPjRVdt
ihktUYay1e25QgpiCGXDy/DJxEwBcmRhNAsVPBcmXdwel8H2L3hhHs+6rQZjr5N9did4K778ruit
iUENHM/E2eCNcdl3gfWoWZaUcD5mT2lVzg/JIPtbF1aySNG36P7h3SF1CrsINlFWtmOIsu1LOdms
c4SYNFze1P6zipuPnKeAsjv9ZyV3XehabsSYqsvPTbZ2iw65yIe7kTyJTcbtORtWoa17L32wg6Oe
oiTwdEMy+Y4LOaLh2F+sDVayu1abXD+n+0ZUzZsIGxBk8YGJTaZq+nPM0GgalDy4eTxzigv3vbCn
2ZmpgXNIlHbTiHZ3TXBkxVU7dyaxPXtKAf9H6K4dP6DB2xjVOTNTrGU93ZL51z7qBgn9GJZ/vAgo
SBO1SmMKN+10nbhne2oEkamS05OiyrqHIor6dYEGo153x+0ugXOmrYZ4+yGknC6Qvc6gtWo81ngF
bkGImTjWnZHx0PnLlc3KbwWsAqiy/8Ar89XxaF2A9XoFh+heZwWvSeU72oWQkVXcI8zHUZ/UCdvN
7R4GZ76Eg9mQsnT7H9TO0oHr7BHTtPAEDj9nxKYyXo3GdoQLaN5eOMcXfH5tS2aeTdbHb6keBQCD
FLvJAza6NiSFpmVCTCXJ3ffE7RONGzLhAZyUI7MuRQyWMlcbqWF6UnjlQobqD/5yY4TFaxeRI35m
PiL0GHmZWuFU+5etlxrGZWEwd3+y9wo5xcHkV9GpjsYAoVqDBdTwTVyLVsit8dKR618o0FG5O/Ml
5M+qnOblhspptOKksPZZEvekXGWizc9+XT5t7QQJj2FvpZ5Bypsh2xooZ1CgXT47D+bD4PUGWkwW
OrjA+FA+hPLuIZhU2eU6GmdE3choIGha2LBMK3pAI5YlsCVtb7M90FccrZ1ob54//sSaLnv/Y2gO
a0hpBN08byXYy6bv49Sk/0A1lYU9mSLUTnZjMsZU+CIIA2f3jJa+EP/E07lU9HuIaCCzYMuuszU9
pJj5+2M5aUvfX0DqYUNuAJN+QVP7ZTjElJRUAnfYq7Iu/JIE/mkQHL60YrDpuqzubi63h5Fia8JW
Q/I4bQqCMCou3ZZTUeXNpXbJ4Y7qCtdFrlBZjamEEiyDK9VsF65Cidpbz+laAuH1PcqKOwb0Cu15
yUU8W4w3wUxVfkG7jMwTWbPqZtngUjdILgVTsX6esWCyigyAo+nGjoDXrLgIXm6pF3Zz+aBJgw3E
CoTSKNhEhCYorVJt3Mw9v8/chTUD0pdCQ7wUbkRX78E0obnEYEXLXCl5PQroXUi2c2T3aye66cdk
/YOm/EuCJbs/8gX0X0cDkggYk6eXD0kwPybaxzYeNgQWAWQp0HCPHk/4fXrE1Qo1AkofsKPYEHmA
fBgSo5x8RNXo34O6upmYIOpWenKvJLJvYxV+VhGhp3g9cluM3cgQY4kiX2JhpEdoSG5+KxHpkoHp
BRXUJWnB5OAgPwOwYwaSH7i51gSC+ncC1/Ty3SSa0ImnzydO9CrfOFOpOOu6UP2wQ9cwj3thdnad
Da7ffIZFjO0+c6BUoi/DFBi0YyUB4tjdaeK4fwYvLakciZeS99DhP5FF9jaYN9Qu6y+3+ip4mNOv
FP/ueNmGqnFW+uldUpHxtWuiNBn/qfQ9oAozy5yHl47aUX4XJG/W2/wEfXpG1X+3yPC+3e1dkEiB
s58r1uv5SSbexRr1kM1vvfNgDYWWSYat1fN7E/0bGreEFGLSIYAGI4DoRyUhE5PsDWvBxPvElOQB
rOs7mHvCxseOAYaJk0aWjscJvbikyFENtGyVJJCgEDqBDYQ5KHKcfj1CdxD1rtxqlVFAkV1+0LSy
xavtjwIKDTpEOKWSNwVZV0f/zvTS4IBneIOjRHVNtxnrR4a9+1tj+5MOgeEUg5AuNev1rqJwbZVL
KjRm1hi7ljkp3l6VfBFlZMjCNPzksoPl2pRGQRR3fTzQNZVmfYjgATMYLWb060511kPnfn9CTcBC
nS6zAqaZjLPujBTMYFqWhDCXSzAR4KHA/PDLQRMvG9XR6XzTWlu2mDzaD7rOZxCJ8TAfa95eai+2
uSiS82ZZ7OwRstRv1QT8NvmzdV7wzH5Te1+NHVQsiK6GfvyZMn563ADseq4+9rowXTJn71ZxuAbQ
Anbyxi478VmPCBvnjta6cRYwz44QXdzW+WuaeQPW9h9jRJshPw04rp34sgqf+AuXwWz9erfHaI83
Uxg+2oPXwF7/S8yMJl8MphyRmuy9RaytDlw9/4ncu+HJNJ4WyTYqeU52pmWX3hUnWqzGb5wIbnbD
bZMpeIgI57drJ7OSOGEUNwn3MM7zDSeHAdSdvqR6L3aAd3ipQFVr2thYsfEEZmii/mo2ScpCK9if
yt3ALePGiGQRw5rxNux8zwO2P9In7T5BVwK3ax8FDWDV/p++kVmYeUM367RRHQ5l9D2te6m9Yo+B
imBvroPeD2CdpHFFcIQsZQLdRDBngDdM8bTVBRg/ytddptU1iBzpcg3IKaNlzO/KZr00fxoJzkq+
p0qG5Mjt3McIDi1xi2cqXGSlusZf/knzabdOauKnZmNbmurr+PkemqWf4kGctE+Bls9K4lqKC7MU
hRepgdUqJBEXUUvi1hivf4FeFEUzY0X2sq6d+yZGtMKUsfwE+Hk/MfKibRtjWr9F7QngFPn7C5bt
qU6tDcVJbi55ZisKzuCxf4D8UrjoHmltXwgAOaMZS7zn2HKTQ/HGjF4wHq5dG0zLlUj2SUA25gh7
Zi7fnGWWPwMhGqfZ7gSLoo0eLjvsW6eOKlPRc3AJL3GvX4nfzoowXIoTKizmmecFS0ayjbBor1b2
BBF+RoAp6aVp1GKNTt4OTIqnqOtyukCzQAR3sXq6p7mdPvQzOBp9fDaS+AvwHPX8YB+v61cGRPwN
ezcjX/JlK7+GsWmJyGN+NpC5jRgxKVWU8pfpvzMlIikcn15vUebp4bKsMnX3Ma1FQDjDcijSRVoa
ZcmprptaR82hGzct3k0FIqqaw8v9qaNXhjcfZC2tvxty1DZF9bslqeEmVzYCD+xLb1OgI8cIhHZc
kkLYSHosu2UTpVATV//CRCJGOUj1PwQGcfwGfpQ0VHTg86O1UOUlq+D0/ShInxQaJJgJGvTozSFB
3ChlakG8T/fVyMxKbrlQxHAXg63ozRTOjI1thyUQbcWSAew5W/x8gkuzbBZgGL3pkJia7DQkWRAj
VfhvPHmTHE8SE6YsSzcDSEmeNidK8dDrijld/ptQ6a0M6Mi44aeQcC0LJIr906EGr642iSRY9hGF
I+Vud+vAiM962Og77YEDUcc2iGgEQwwaodpuk7gMfiiDwG3iq9x+/7FanX/uu/VXF2Gp0T0NJwbX
L8UmW3g3bXfgWax1R/6voaDRGAycrrYeqoc2ZRastGMxyVDqh1aY9UIrCHUTfYlFJBg5cDUaR8k8
9VIVI8XeM9Fw5VUj6j69TCF4/4Sbmh5zf7Qc/epLSi1NfYF7Pd8ToKWCdSf/Db1SPFZWXAfxuyZs
BPGfhRFG9piqcjKnJbzGGCgyFaZvMFUQleHRyPEmREmyyvR/HAgUI8NqovcJ9Q39n6oYfT4hq1Fv
B97oSHNDRxLUUq57/cVlRcf816dmiZEsVHn02q294q+D7bYuELhiFmfL27GOcEMquASDp6zISSTu
SoPqJ/AiIQpq23y8Co4WpEK/MknpIf2/twQxC6PogGFEpMxRpzSzvJwLxh5OxxjTACRkU8P3J29U
nv5LHT9r/ba2hnW/xPh2bnVAzjEUOFbvBPoo6b/xMZbNT1/EjDGN0mL8SjJHf7sZTnzduX9gJn41
/+uctj0mSg5MXm+Nq5piAAHB7ixi3xpWjZJwy+X3MJv/aJA0qXeiC2vpbQ7zWPeuCBAi82TVgtwK
PDk2tjI0HQ5ZyTfxL7jxy8P5MpbBfjyfQFO9JsxRIsFlkuzqrKrQMJP7NcE2tW1XRMuuvoE0EwGu
XblBe0bTbcmP7Qyeh2MspAOvSm3+wTyc3iIZ/m1Lr8MWN7zO+R8hYQ0s05bVPEhVvknQgLP56fEy
AY7KUSML+YHmaT3DdaW9RePV79JifVXwRxMcQVuMvYao31FJ36m8yxqGFswMBhPVjRfIStf9aBoD
0Rxw6GiOUkvIOO7g8JBZdVsZELwyA61tkKGKG2rfzPTlNeFDHUv0aQAUV4XpOz9J+M8jPuVxSLJp
IQgpatewAP3CqUGo9ipVKlTTHUiyzS0/so5i5UfRVfoGunOKssMpgwRpXhZ2yb3w4eVh55Mj2XZF
kL6rj3u/PoREFcQ1LWfYKDqjyazGZiw+FQbXuN4QF5aVabLs/lbSC+ecJvEyJqHMCpthOdto2eFS
r72zxuFvJ0VpLMRhDU5iNa19LJbGhbdDX2I4uBFaEO1CN/XVd6fInWmf2qk2TrIssuYyTeCpXwyO
4aGdkCCoXi0wVBPqNQPvFoUZ/9CLiUcOiZePq5xavY6toncxDQkWpssitzZJXKleasf+b/AiQ/il
R4rlTqQzXxSqsdO3z6cI6zxY8deRmHWHjjW9vx7uzvBx5M2qfntcWg1BH9v5mxjfUNM/P8j/7igw
syaDP6a7FxHj2cRuF6y1c5IkAsdxEA3cMhVGYtOGhSFXMQ/TKri4Px0twaFwlt5uXDUSphRcu+co
+sORcC59VkThLcC4SN4WHcEPCXmzPeGUg7lYRHbIDFAVL2uJpADQpmRMMZIPR9FEdOf7ijEG/yF8
+YhW+RlzD2Kq2Zicn2KyyQEGodVaWvcF+EGk1A3f6ACXDV49l/Zrt3/pCc8Aw7vdOOCFTDkPMFiV
yy/MWRWc82N8YpCyASXSyd8B31bqLZavQq70DxSgfFvCM806cc4HieN1jDSELCMhJ3mo7ix380Z6
fUfgfs0GHgQDZV0m06ReQhw8RltPq7JdlwL07OtAZnhfGOicEHsFbwMatQGTre0rw84HdeUfwhgW
AZL/y/gPhQ51SEq6QGLiwDVuPKtf5dqNEF3vYuIywLIKIh671412cuFXRiiiJbIlDFmr9qwAdlKT
p5lScgxfm/ZQbwAVbv4c9HDy10pnOM2nt/JjDjftDQCGWvg7chOAVWZC27G7iQWovYmu/d1Gr6Wy
WfM9ylbKghNa4tpUaC6q29K+DX+Wm50Q/khpO4tfulnz84+oJYT5gzhvhhmfxva4oTm4UMDAo/q5
hYXnA8WSGivdLhKCdgD0/+19UzkLhhQHwedRK7AbiAv8FhwW1/sr0yu6Aomb21xySYwSBeh1Wj1q
YIjQLjN8AK2qUERPMAwwyEt6EcWymtXqNfl9FiZ+vvX47K5tTtgRyQMFFRSd1Il/iltSVDuw0wK6
/rlnVCuF+h+/AiPQ1m/9pEJeqP7r0bJo8HING0xd3vDG/yTgazaHJq/sKC24Dom+LVwZ7KjIbEbB
05KvaXcqZB2y+wQJzocbWxxhzeJ092KN4YtBfkvAoA3INBhi7eYIYmGZSY0PjN+XtNRuqBjRQ7IV
3x4hDAgAYb5GZFx+3i4Qd1P+amYgKUuMBeFWQkdbFUxlgH71whRWgqywoGuNQ3BbF8FAMtKoGrug
G4GKGGol/b/0uFFANNd11+rZ2/l+WWEw5fsDEUSHmPsm6H+Xm/M/LOol89+KVaavxVHR7AvsfF+/
+dDTOd3UUNNT6NeCSzrYO9QagxrSrpMyVvD7FbTDCsSP7eGJaDB9QXnwzRbhTRtkYuyA0ZkERpAn
hgpId2D9XFx1DVwHZ7VQ2FQWjD7PsexRbL/8CEJfZaVHgD4hMvH4joyo1K4S5ta3BZVJuM402HpO
aSWjzE+x0+6SCNkQq4k8EEYXyOe/+98q0q/pGVW4IyI6GlB3tsGWQtzzromXViVdj9HyybFHs8MU
pj0Lp6SGlR1e3H40aQPBc/+IOZN2jKHs4T8K+pWBzkPwOpnOMAJoPpXG+r101Y94WEuSuNqDLJL6
ZpF+TloaioNwS+GtuSaoZBoyODPwlIoZE34IEC1eq1lTJ8CnIoqzhuQUh7REFFVSU6pK0aTLLbit
DLItcAN8F7CN8XJKk2A56LBJPFBiSOOnhVo/2gIdW6bUsReSDJwdd6O/iA5mjFKbDi9tflsYLjlw
W1e8gIkNqoEXkO+K4EwvHtIY7Pn45UV/Y4pz57ImDzr1+Y/mV4Yo1m5cc7vlVfGMCdoUn3UgB9Ku
KWzaPMXmsDRR+P2w/fH0KZLfZgd+AHNob4VP2RxURDT4qmOQtlO0VMOn0y6Q4niptHAklLtAKqFw
Jrfk6dcLnv9pTiRRCZnjdi0FLzM/MKcb9V7O5SidLmTzyESkEUcn45Lsu61K07olD7mlqW4AVopx
SMurTWhHvlsRsHkZEmOPOk/iDgmkK7ZyKHKce2ITXfX5EWjiU5EN4Jhk+sZNdyQqAQMRDzFnw1Hw
EpOWAa0k2a6IbqL/s/EY72lldh2bJFqO/C5X486g4EF7Ls5gsfnSvYQ2+O8LlX85Xkg9FkCUmZ6J
nLEkCmTGgCk/18U43GxiQVZEsjOCJDWAUj+W5pwAFvwtUgr+ZA6ztoNQ7IeA/2osQx2kASnYDKU7
eT8KNCj5AcMmow6+P05EhJhCNZDdsjKL8mc3JXYq23TnsSwL29K56g0eHJXqP2zR5Tt06GCmExae
1Et7Zvwr9HLXlEHIR/rUffvxdIQxFFyHlEmn7CACWIOYk7ZjPydjvUFENDahgkPL8mx6+1+IJpZv
7znQwnV4hn6j0RAqbp+C11EorUvdjkZWNxd1ZL+Mkr3uWapYWp3M6dyn1Jc3G204iCpGFc2VUQ2I
H7oMwV971si3urXVTSbFY+UI2qMg1wWc5h6BdRW9v8CXwyKb+/2y/45B9W7vkelIy6QpZtc2khQW
cBakAwvx+qPR+X90YhoAlr8cs8w5ZBr6vQs+68GFii3Sm1rDFMTdpKqQEcymdBtGlcIcFDvyESLq
QRkTZsF1SZ+L64tiDo0zs1TNIBiLtNozK752felFjmMbgIVgTjdBixiYeEm9d2OFxPtw9R/n4Rt0
eu3jEHWjzaSBVOH3vjvwfztQ68QjYMFTNYwXE0nl9tGyBF11JTmZHDKcQazI8xfA7e9AmwFsIYSl
dpcXngqextTYvMEec4dp7HN+wZ2AN6raM8RPmGtm8wPhktdbe6OhjFZcmsNCTVEcOUqS31jCw+A4
yIQnovfLLhvS2tVbW39vMjjoTHQzOyQ/hx2JUi877hPiHNnO+j6fnpghfEJoAK3s/SNM0XotALTL
onInbPlqZLH7LADb0r8ro3s6N95Rk/nQGhwqoLIA4ps4PVkQrWL91PtOkUu1IcRxK0Rz2Uy988D2
vWBJI5bCk67RR7LpDU8pAPphu4O12pQLs0feIHsQwk8zdUhbuVoxqApETI/Szls6AtvjnfeZ7Lvh
S4fwFc1OO3cZBrxPe2LFyZ3X00GBwgKpFNhxiz6MgFr2hMVIjUXa+JK4hVaqfMKN97zbbiP7AgC/
gQqyNWCakur+3tUnz8OfUivjfHl+4FYPv0y6xif2GMKrhzOFWWE5BihfiMoIlD9Lg3dH+G5csXU1
2qmeSQm3zMYpkxkZC7+krZFRZXFS4dSKVzeMrvJBr2n/Hzmo+sCvTH5jO4xfUaxh8cTdBXNywMMz
PheRegSYpV7wu4ssAIXmuewLeohqqoHSddl8ckiFEU+O6zG1jCKlFyxhENsNsyr5FeeBn6NwYc9F
4BXKP5KyqI1NIEkEAAL7sof27+egPl7RqeEcVhvyUNeCmYUE7CV9sSV4FQo1jJ7dmBHQrwlZ4J0A
UsbwhFAT9ZFAyEQIE8YB7xLjdWnbxbbEoEu9HcdNpjVKxz3wt7K65d8d7mGirqkIRXO4WYgXrtWg
7Ov5moQ/G2gn1D8O/6FRzvu2zKLYV8LZ+ifPXogoDsCxEkPLoboMyCnbcuqi+no9ScnaFvaBZ7Wn
uKk3cJs38nSInAOqcx2VxYndecfvm3/2pP4wqgsN34Kx1Pm2tt16ITPyg21XcKYKNeRldmr5hs/9
FranLPVNKL5X45QOH1sRhZDARu3L+CZz32okLL6exSslmDKtL3v81iZ6vFwIUlYmY3ix6bfLuXUI
Zc8wTg7JL54VY2UxZVros1Q7UeN+anjCb0SiKCOx1dedCpGBMaag7lQOPRjZHdI2oNTfbOLhfcTc
3RXKlMGLTMLAY3lcgzDiSHgDk3wp+wg8WJrJAyfJbbMJsAe4F09IcVdMPaSUsvWTBgERB3K207q8
g/aHijc5Xwm5tlMEsq6CQ2FTpicNsZeIbkjUdat7eN6zruvBqbtogq1SlhFOBPL/wo8FurDdLenz
j4yzy0b/vQWXdgeVOqyvLu9pXBmeR6zfTHuIkY6QzFS8HBioQcr3XeOEgUcfcBCeMtoimS0E9HFG
30HTA0XKcgoT11OV+Y5WkvmPfLRueKrLUKUuUQDiaQ9hfpK3xdr9p/7+3UJKyS+Awq6WkX/M3r4L
/CzGvrnVg3khJIj8l3X7B3cfqpoj+4QwBthwTtxfUNPGxyk1mt4SrmvaKZ8gkLmz/i7tRGXMWSA2
Rty0hOI08Pcns0MzFErw9DshuIqaXDfBcTe0nG4HzUSdRqnZ36gZAnaGBlWWgVLA7Nt3PPUq+Nfh
yOg+4/BQ3BNXRHEzKMvaTAsk2I/C874XwuJTB/JkTxPrufYMvXLdZKJTlhEcrVK+8q0WH5fWk8n2
dZ2yfOIs9E6kMRzNevl44WfaSSq8VFwYSVV3lNbL65IO89eievHZHRbAD8hfcDQN/BmNDuTJlA0g
X9N/4IDK/b6nHbUqFO01xrYFKIU2NasBETzjEzVP2x0ZXYPB4273x6CDKql0w7f5YWAdWqxhNUQe
lr7IzpLeg4tq7C376YN+6olvu4xf0WRpqZmoAazF5mnFFhBf1u1hvRU0NTKUHNn1jpiYvHBQKO6/
aZvBN/7U1uOGKv7EGHSKP6oaP+X3yqZ5Lf7whZZTUIduhlcmGJ3Kpd6xzfYQK6rdv41BgoJQ2RhY
AnRLUWLTfZrEijRyI0tE+R9jdRf6uefj7eVCkfhpRPqM4pqtV6VN2EFfbpDOju1qkGe4mAw0Lbe4
ER5q7mzz/mYQSmwIANTdLNgco4IEkYfi2WOoxtMWtSKK2bUe3KvErMkoM9QRBDC8v8PDRPHj9M+V
k6WkWbhLTMrPiAfW91nZal+rVcvSpyF8Z1bhB20/2sysCkIxTtxMV6TGBXtCRRY/Dc3I8KSGer5J
kd30IKdIPFgQuba53EqjgqtXN/S25d042sp7dY4NN8j43xPHTois+K1JIq/46RfT4G5AsIrMTWEX
2c2Ugm+R0TNLqIlyatGUd1fmxv21acALmmu0UuqIA+NNeFWNxtWN4g/W3HAf7kCjiPvMcCvcHA21
9TmKD1UGDmJf7iZep/WAuVbA3DVX5XVaXaO2xoqWWdUlqb+k303xLREAP1iv6D7gUoIXysV6rg7V
HRFZks59QF5HbmTJOaxlfHEDsyBKHBrTunXSZIJDGxZLY4doirWjTnQWad9ij/vsiMAABUvdimb1
mzUTM5dYAMNAPul1qxpXSlzY5tNMV89H8F12/XJcGxXNOEfSqgbctGQh9yXM56ZfUyc2bt0jDs4o
IFp8Mwr4sZaSajy3gTE6Y+8ezvvoxv/jodC4umGApminyqgZps4L90SdV9NW26HI6E/1OMRyXrrP
BE6yK5iYryjPbOZ/W0R4zN/fcdZLUmOYMd+Ga0F9lyYjLdRa8TRqvl0unrIBE/IQSDlqee2dBzdf
VZQypdReGfp9o2TbBRFuUczkGHEfQ4pci2KuoCkYaCKPvjD1iqQ7abW4rJ1QJKDI5RyBrs6vkMYU
MC1nM4gmSDgc6sDbAnRR1D//s8FMriFmmpMilmho2iDJQ0UQKVNB7g3faDkfqnw4+kB1DO0MWP/y
yZjKrKb5lIqnYigtWyMXQtOfUJOI8H1GCZsJGdkcovzMcYhdLXSD0i5LQw4dhQilPnFB1IY42Fz6
ZUXGyE1TJPit3qDvna0u8uip4RFcjanKFmmf7zUwTSmJA3J3O/2xW6qOy0Hhd+Q7L1ASbm11ma5V
NFgdw6MC8IYaL+5W4Bwm2qwRdye+Bs3zi/JLE7ZkPxBoCUafuJpHw9hVtS4oH3KA2OUIFSkFaNcR
xm2yyPc0L42y18eC3s+oEcviUlp7i71iiBys600WDrqXvI0vyQ2zlp3ojRC/xXb3UhlHJ6JDqjqJ
tsa9k0weoUhtxU+LMRbXVVu6pD0tDG0yq//EBfTToB0i1AjZdPKkXf/24R5FLF7iT6BHj8eUEClc
KgblTdeShwwL/cJo0nOO355EtSSbI9o7+DZAhbOB95Bwwx+d9pCjQ8mWOVM1J2il4niSmUFJaNlF
tar6gcr1+Z4c1jaqUJkcEpnhqLQclYRBiBn9uFPL2VRZpMl1czbil05jYh2WLip8XThPJO+XI+TH
pcW0yXtO3kpgZotHvNGKoDR1/vWHQuAqKq4E7OQwliq1AX5JwLhp50MXEeVohRYDNBDl1zPpCO3a
Y2z3Q6Q6e7KrpTNZyBTuHhN3N+pAiEwBClsTg0HRGFXQcAKbJ3KwlS/JSC3poAcn+LP6Rx1y3MQa
GV3hfscAuq9EsRwNXMBcVDiZGFbYJaCKt5Eovz4oFlQHKAYRF+UVn798JRpGFlnCdgeBoYK6V08z
VM5HYeTMPoFe3w7204k/8XCc5W5F1ln9AjdHmeeKDlmRErZSNZp/LBcT2drAIdgC5c+w+F3U6//A
EMQra329eYCaJ49ClNuEU/JvjRI5WId7zPIPZkBSKlO7M/5D/MHb+MA+8zkzg/KUYKcaEaWPg9l5
/6oDHnhozwqqBTw5YXnKodpw71q21VlTE+jnKlE2C2MM6qzd37ixVaoPNMm562nkd3+jAWI5fi8r
JT4XxGKPPmpVjic0LjHODjV2ncyO0ab/yXAVAA/DAhkZQ8mKQzSXcPxnw7FlpeG1r5+ZRdnSfvUL
Mu3k0CSEIvC9WVgSe0R0io2RDpzCdLvaooIkzA/6gqbxjbgImdCxO6exifWIQMO6QGq/OQPv+U8e
tEoCJdCxM3qqkz0TpD7RymtsigPdjlOxPFP/eIJY4CMlcAIti/oOcTiG16reVVLjlosCk/0wTJFy
rIPu7rzqjp5q8bfGtRSd9NUzMUDd10fDaz44knOXJUW9hbDRxx1MaQhdIdUktvkUtfYwz41GEyPi
KKQ/UNRR73ht8mMWdOD6t3q1mm8LtvjpUZrIVjO/OsVFaJN7RYRwmuF1Yy98ryZxzsiIOvmwboJ6
45BTOecO970mnlR8+oWp3JK1uJds9n6DCpKG+6QAowMpLnfMKYCg0GwToifgUGJdpPn5gCGpwR8f
Z2rplXPZ5mZK2tB/Zw87RicUGVyjKmPpx3npY7FI9YoqiHmu7BHCOSioyU4CwYO90aDKSCs07ezY
auxrqT2AfODY9TknIVhE/vdExlRZS43dOepQHA/FmDpiIVhVvrcNXeNnpUpamxMQ0yllCLIyRTv1
aKY7q87oZxXWGlY3sXzQuv/eh+FgZE4pCt739yAKETpUZYUP4emwUAil9jQ4V++1xOyy7u+vl8fK
a/DTN75KMP/Bbcdi1FU/0xKj5jGl3n0CwAFpvr4NHxX1mPwl315b17cN0z+C7bOC2Hpz0PdVE1am
9pxCVR760vAxUTOy2WRCG3VsgwfkoiV2VKFloaog3zLUyiCz7fBq7dKCvUACge13jY8i76P2tUbc
lcDair2cGCP1MOGzrByCFYM9zmsl2irbWiivWGGQLjxdlU4Srx2D//6AaY1+PDeue5dV6Z+tiFqS
5K80pD6BoBTSI3utxqOWBCmTH2TBXQWbj5Z9v3XlFp+2M0cXOlVGtMAYkSld55Xtr6T8hM+Ww8qS
qVEIgsbdlPGh/pZvIaOK1SxYbqEcanD79bM1TZAkD//3dLE9q1F31BRuLziaASUJlkGPf+JvyOjv
Gqftu2QP1uw0IGXGXwaAUIaanS4U1sAFVVn9fy9UAE5TH4FDtRo+nnw3mgEp9FHH5yHh3X4sZw4H
Ty+0dr6kVauNBMmF69CUfwhmoFuKz5Sf7XTILVPyDzApdC/T6+eSIsHFdmD8BX07dQ13Bap8Jn6E
c2EcXAiSFDWMPorL6FxBopQfkQAbA1OKXJuSvpvb3bn4UxUZDPhT6YJhNokpOmXu8/Ul+MsAPsID
h0MARNJAcCINQ/TN5ZjyxZMXUM95zY7p9Un8cC7fYg7uZSz9Ra1Z7t8NaUH0SJyMSiYVvTizbFgT
LsEqpIgr1xL1rkmOdt7Q2lOzS9mam/Z480ZA1wKUshAnAfC6CmX6/K+ppU6A4NNBuQhkYsmfFWKk
PqGLvlSsC69cZmTcO3r1cZqxMzHHCdBpFgqT8kEO79plla8rK0kYq3kbfjSBsncytVo355c0H34x
Nbnp85TkEmnBhiftC2z/1dfM1rudTDdUxEhiX0eRSQt0+piYsqU+/lSRZbTa7w5y12HK8UDpZI/0
SwKvKC5jHEN1L5bRvNzvm/XA6VUcKvkdjF7E/QhLEkfGpHC/bcUHPaQGROX+MleQ4V8DTjVta5HP
xYgDVY1e/Lltf1tmdXMjN+uNmPNaofMnd2vOD+QJA5bh4TBi21YetOYRQ+2pjwWdIoytQVRRYa/8
Jnl4s8eG5Uv8K4weCRnWKB9Mt5f1Nz9szQyzay4dsqVhy6aOjRjwo2DMLIxsYBQJPAaje1LpoHKL
w7LTKf15w9jBs7jnXZ8X/4MbKPCmIGWaVuhrpZrLqcHgDk1rSQGO9ej5kwNql3V/mWj+mZvN7gYm
OEZMsO9Wd1KyB88uzzH+LGUKDb+IIR6DnVuZIgyr/ASKi6D2sIto/2gGZOntdNkhfBeztzlo4op2
NXRO86+buFmmmxzCiqOqdNsjj4wIqNADPm++/Zf0Loyzi/7Fa64A8OTpObXuxJtLNJmSPXmOpXlp
SZhayFL14DT/4Cgk6Z3VI6U7/8yHV5+mS9D5Kj7Jnoy74VKuIIDyPebMI4G1yTvfbMZmFF24v0rj
Ka9iozWe77080QDqPSzBMZuaFCiP2S/Rff5zm+AQGXbQ7AgmDZLuS73a54slTHQ96Dtu8CatdAn9
ZEU+zSRuaP26vDiadjUW3FIPDJhAfyzHnb0yJu7yjybNyJisaJzS568BMXSDDRq6cGmk/I7odJdT
DatrChz+9yv7FSOMtA51z8iCYZdydujZ5FYQ49Piqn6myhGPDf+QtRwteN7evu6Yv3ruKFaZkWeX
8zkgi4cnmkvd4PnTqH2PtnMQ4+8FaH+bsxeFxpXKbAIZXcwStndL6Y8gkzcd3hfFsMXa5K1ywutB
qguRgSdw0XV6AgWkW9lSvZGRvPj8fOW1iFIQTpGSzb5fIHOP88l/WQuGXYvkAVFUOGg2czBzwoGn
q9rDMvK7bHSNYMuiRvCwu4hETlEXjnWMRqzQgB5eO3SSEypxGmc+yOLyxc6JV+r7OXqYv5lI47ES
eE9FDa16QhTw2dt4nnt2MFXPhBOw9Tk3p1868Ik8ZuBA/WVuxpLUXAP7GZHm4tPwfE2BWgN9bMsi
V4qi8mWhaMWw2cZ/hp1RyN4/aO4Id4oHsL6x9BkVmEBYOgeIsgewFodv599HhrIIr0CGQsG+By5Q
kvUZ6Yr7MAOCHtIamd7QaPo5bf6PUSaVLCIeqq94M16rKycMNx0RqtobBACxfgWQGAAYe4I4IQeH
ElmHiZ5KPJ6/AsZkHgv4FPIeBoN7ApOqaBszePWKGe4YVPHcWPyEA1CSk/XCNmnpyaoY6Kt4Rite
4QHl0kYL7r0DuhBB7FczfiIjpIXZRy1xZosaGh0UYncFASH5I5jmRtwVwh8//APOuGhZyGs5fXTo
x+w1hdLzKozbaIzlB7ILU57n0AN8jTMtHYIq45rwLTj7jqdNlQK2h+tXrytCCxwS3DWQOTOsUiV6
77xJNzFLjfn4gcEKk5di7B7peAWWjhAFCxLNB8+DWZGUOCQJIKdp8ROqEIJ80Ky8TmWpW3ioa2Xm
8EJnRzg9muFQYb8eaRZYa+xg71TnahWzqleL0EGTxXXZJekdFMqeLLAi/RoU1/a0XmElBF42gVfk
pzhX7dexNvYMsOTpEXhbO2JP3vPJHZ+WpjbPpr4Csd+d/jhF5mDwVOFGJaiqcpFbahSQv9NtbxWJ
60tgUglg0V/yaOOx7iPez+5oDTztq6bAhtk3G0CkECMBDaWO5crqLAiiVZ7hXxeDyRS9zI6HHAOJ
vpIW8XaC4YJbVOs5iixQhSzcP/dfrvKlowuIecZR1HGPTPGp/0serGdk9behO+KcAzqxO1vYkY4D
IoPGKegFXrxKk47xWR5NurIgHW/yF0O/bsQXKknKNn+SxcnI8crVPe8eIR1ohR7OTjp0gUeec54u
MdRuM6qba37q3I+roEOSU8AA90XIXrHq8e/cC6vy/Bl65kkEWt0frNZ6xNNOhQL4NCUpSHx+LNSB
t66bYV0lCUnppgrvmGD6vz2q58yL42tpUZX55X6nxGNdtze8sWMFgYsqNAaUA7O84IvENjO9bjo4
pe57oqlBbcKsrOWKq+Z5iRA8ndy5TzD23x7hZo59lvyxptx630xf/Y8ZXshWaJ1rw7ulebUl2miM
1SMuj+GuQ8vipEbbsdsdGc4apCBVaUrgWRRgridHQLk22QhVW0hkbfsf/Vi2y8XaIS7yH0uBn/q4
dRrK+gneLJtdclJ0J6EGXHXYFvpICvdqYtc8ei03O4WE76rDiZhHFbf/mbYCWnJBXCvyN8F/vgZo
9KVRlMdIQBRFDEtrFHpTFVP6jjvD3nN9R8gM2rjTTrEHmTjz75dWSpdDzaTiAqEv5FFz1K2ASdJl
C9zBGt7yovoL6CjGdIryJYRrgTMnsGJnDLCYZt7L0xpHhslsJXQSaoMA+X67NI7JEJKPtUViC+Rg
ZCuRcKOoLXOT+2da02X1T5pTBQk47Z4/pnwGWwXB1N2ti1RYdwd1k1T9lttpKb7U6kikQdMl0Ks8
zIkyx9yI18AprMoMygCGXASUjhPfxLTEBKmS1KfTrugwyrUfUM9551aWTx3QqHA76vXcCMNSvOpm
bH9Hzomt0iloot14yofmhMDjwsxa8xoGRISwf73CH3dMXNXd4eZOxXdyJImOLyibTDoYvQaVsc5o
X/YGGvYCnqihIME98fNuUmrS3YIzZ12cok9fYT8ePOH8n2R1oSA5SsEbv2bn3ZhZ64+C0TJw3oHV
dRPuQgEYxl07H61qq5dZOZWcId6bWiKMItXNFKXt+h8kCT4eNtTyyAdmfAoMmVs7eiNZiJS/vzm2
sad2Fdiv4UKjGqLR8/6ruuKLxuCqdj/HHqpkf/maZYDAOHDb2UQqVPDAdnVmH/z3eromQcaDi5SK
donOhsaYtHQRSJ7S6JKh7Db1d/+ozAlcF38Q6GaeN6GtdereKX1M+x1Tk9bs1ifPBQE0lCmSGCV6
poqbeYzTLtjxBORtVhpWOGQg7Vuz+NpxW8ONaBcfe/RBf7EGqDImqEWfcBnjRaFEr1jny/rUZpNn
s5u6TSIIcm+inDV4ozV9vZP5yokhLKfeegqLrEGig9/r+D3bkZCAXqDYjIEVKIlral6o5xziP1Oo
QFp9j2DLXiJdj2WDUcPe13PePfY52JSjtjWjE/XVakThqQiItJNEvbsSl2z4LneTrmjP05ghEMoc
ckzGQHhhgzutOOj5y48/A3rETn9L4PyfYJ9mtKy1TBfuGX7PrT5h+FedpUCqGbCu2ZXcQIQO7QDb
5sJYsXU8GTn9K4r1AkBz2GojoHL1BXd2cWEo+Ybrh/5jd0SJNyRs6Qo6R0sFI0TeN7nDghWDH63K
+HtJ7lkY0Y7+MevWMIoBZgxhlAxFgoKRFdA8kobgBDeDgAc0D8ubWycTnVEx3jGu7NtsgnWMaYYI
57+M3myY8haFLd2d7iMKZ/Q97Oq/hO/1x0bZVqg9Ljrrh5sUc4NnbxEWrwhjRi6kBSfjHgc7whUr
QbiFg6xM26u1SgTrZRiU+PNgEjiQSHG/+fjfhszc+rujGJAGPVs+hPlVUZaFJefTjEc7CrxnAqVq
owWTb1yDye0/RfTlpfshqhPLd50QV4LYEBG0qA70PlX98SWhCYxqeMloJQYtJjtPzFE6fNl6btif
xDQWI0ZRLGU3E5n7Onjti5K5608VEQ8hducPkIrc66Bjc7bdNISgIeVmD0Ykira/ojDpVciybpUm
xizCS+AkL1mtDwd4gKEk5Iwy4IiYZIoDS89N6rGq2t+/dw/ww0IPTxpx8P7jJyCqXm3nwK6jgP8z
LYWeANv36VDJ9y3PMnmjl8W4KM+A0BR2QHpQweGl7HkhlSNMWvR8IE/Z4IGxQ/btXLZg8rkG3nD4
5Z/YGmLtHd/AZk8nqZ1QoGFCUV/S354NwrcEAISeu5qNMlmrffZQ6UCdvUBC0mK5MoWUVRc64Hn1
33yeHztHGX7k/eCSsWXgKpl1CGKCRXha86xR3uQVS/Qu4eeDnzIepBWgeoHyHSCLePjwGHRRTyeD
2a6L/65impN8pJFiNBteUkA3SUwyIqkdr8rvZVR08gKceYNzlaDHG4/9lyVXy7MrZknQndUC0dEz
e1c33O6cxWNmuzDDfbC+7Txd2LvamBKRRAiHq0j4qTS2vGL6JXxEnYXDuBQruLeBpfzjUY0o7qbd
tRShzlF5mLEXFC6zWnt8iSwhHbL3cz2TYkEFMFLpWyafyLW1dmat2069c1VORagCAC+mPrGqKIkt
OW2iuNIAE/OtFnAdWvID5T22MIvD7EZ6ckBX4vDGCfMPuexsNjdiEcJtzgYaKQTtJvHKDdKd5R24
4JD16UXm+d7ve8Wxu8VHHOgDL5OpOv8MvGYh1yp050QjsxbO9Vq001QG2kGD0WvXlVnRFDpMXk7d
FDuE5hLdOGYuFUQPoUfZzG4KprxKKd8JhhnGQRg2fg+Jf9YO1kYEm7wt4sbow/STf0700bnxQFsr
pO9WqHG24oWRK2uw9b/D7zXy6qYDJTvNcQITBaHkwcBsXOlQQlfx6KLcRQEQbyzvXZI4q3ORhVGM
tql6KeOw38CchMr+YsBE+v0CdvUY9S/fWkenCrmKhj1FQZrfh+MCm0Q1ZJslbTWAvZkxW/ApLAWf
YNuPUxlOo28hhqYp0Hf8wqqraf/hyef5GYdNgoN7Ky/FoP3cB5Srhe1bsFunXnXFpFh6Ii/izQau
l6gLeJOaoLD6oY5GT0YBphrx1V86FIWY4IvWkMpflVbvgfvQVSM1xZY0j7LXdv/1pGilzydDj1Wd
M1dmKfppMidLEe7aVqOp0nyePYtVMHAQDvI1dqxTDV1XhHO5sJD/AhTUUoesKVPTX8QDt2YPgd71
rDnJHyGypZ+D1r9NL/Tupn4dAJXgUg7pinC1ZAIHs0LbedxomuT39jG0Zi0kqNDO8ijvNru6JWjk
4fyEAhzUBtG3DM3OnBYqUpiltvXjuYKlbUK0ApNRWx2FyFrr8k7JyLk0eSEDReLFnIVW66fUSGCf
IA3gLtmCfW8XnWmD4fPIfLi+DZeMTv6y4AwXnapuO+DCwTPd0vnnB+a/iyzZUbkI58cYZEResDUd
kopTp6Rk3Lz2KrbI3Hhm+7sPVjYI0iddJ0wlp/AuvJc2y73Rht16LX6hHPzFurGOAf78jZYgLdq7
6f8iUtc7csT5ikwzmMaU7z5qV03Pl1cjK6yc95rLmbfrOPV9AcuiUSbAvcEOS2y/AxUT9M3GRR22
V9N2TXB1H3tHlvUtFKWzZmuJ3wHwZ4gMcc/rdL/YuAy/rTyCrTEE9CUsZqq7lO8hfyiH2UQ3qWXc
UhpybHPqzXDpcMWg5Q1dDCrKBImmA5VU8ToiKb1p6p8I9UKtcqbEVLy/MKq3GFfkf3GSotv2bgic
vQx3SldjCi7fnyY+aACWFrH1pZSJt2j45dKvi0ubSGeVmzTh6l4OdIlrQDgzPK63tcxlEt5txYDC
Fm1ixjLih++YIZCpKnHdZM30X46U/WKq2BHRYrCpy7HhQTQowQF98iw++XqJE86FDQGn3+l8RYFU
vssvBVQPi7/vXL/1NhH4GaNiPudUdSLG0CPmjH6xcNbbA885e/dU72W4Y2dcCaW0sRc8xISXb7tx
BM7/F+d1ae3f0+qzzbZ2cVlPOf/Vvl39AQx89gVImcyASx43sJtuGQeDanDMDg8fp9EftybOUs/R
mpMVg08aORydn7ecV/CyWSqelfd7AP1nrRs+7rLuB1YvyRHDuHz7vnGRf9rrK9sK6TXrn9i408ap
foHpwmfW9OtbjG32xVcqOWSi7e4v1sZgLfdFItr8b8JWY4EJX0cKAFaFBxF/cu7j2MByFVO4ZaDz
oI2MDsW+gaopmTv/CE7AcNh+qTjCclwviNTGmdYYmvb4EyS6PdEUO4fTFk1bBvz9Vv43R385K4Vb
W2+xeIwkJE74hgB2FCtO8tMkzGACXanrKYAXLDQH/ERIXoQWQ5XJxrYInFRkskoEzQ1KzoRyPBOj
0jI+XtoleQ5x4ZojgwfWArRKiUMzLFiu9b17geSutBZCj5lr5aVkVRWw7aACXNl/hb75EVk9MlVH
Xo6Nq1zt5YJRGy96njqqZqwg4v+4d8UBaA7UaeLXlvE9meTxk7KR4t9tsZylHnQKOer/L+AftHHk
sBVDCHXj/xRQka7FHy/jpoPBmmKUPMrS1ko98iHzpnl96iXNFa0TagO4jvcNFN8Wv3Zry2MNIpx3
gXfzKxyPg4CGkP3M3bGPERX582UyIZKFTYqcC+cdQfqzbHsE4Py5CHb4TsqGiGtOy+IJC3k3XbzU
YQD/5aCm2dRvnWzZot4N3Sx85uklrvF45czN6HoIP6JTczY/VCr5S0bTkX1+MMBhSLZE/N9e9Bxu
ddid5LIVUFPnQBxA03zAgIhsAgPlh+2wdMaiF5+QdwmfXnWNLVpuUtv9BHgHnMsmSyt4BghnWdTq
qHaLJ2NYCF2EaLIiiW//LzzVzA+9zzzfOpRvksmTn+cfYoaS+t8d7TrvYhcHfTELFcu3m6ZC1Zn4
gDGuShMKdXsZOEc1dN1MxFUTrvy+Q/93U1d2UNFfea5RqB0FgVfu9w7gg0Fd7A+viajarC7d/+du
RpzqLZkzQePLJh+PGeLFuN+J20xBfcvQgINjQ0FZJFf2IEKPyi2/JwT82GDpBocGG2QKTq+TuRkn
0z2HwZn4MJktQYbaCO/TsbbACdymV/rJML2VHwb/LZbl5B+DpITxn1fFgzToEoHlYAmYvEejM9Dy
LOC+DZWbkriOW0aryi9e1yTbNofkhfD2q7aH09VwXGcC+9rC4D/hfsLbNQRTivFRYvgAZpAjjY84
ZKgb+/llS929Tnu2SbidYJsszBMlLomvWEq3wuILQQ4p4t1tKDu4cKhC5xZjTMJ7orpytlDSqorQ
lVAHnsnwRD90dgRPpIIhKWBOpu6LdqH3sRxjaVcQ+ODEVw8pmpSq/NIUJ9DhHZXheMilzpsnpeZ4
em/dnb8OBI+o4syxRob4HHRGpmh7cUs0RjgSyzYbm0V7NpGfU1Zgtve7bJbM0z3C4RnesXJXpvEs
p4XAmuDXQxw9Ab5pOCMjVNy1mxjcmMG3qEBPUgeBHApBmeYwVzKg2jNqOat3BQ66gYla31boOU3P
aB4SZKoZAWnC5jlll8vvt4ecLHWOr9HcUymTMIUgOnZhyXVA1H0jWZCZShD1GKThls154SWStSwo
mk7NgUAxEyom4NZITUluBtisRoHtb6jPL2Q1iDThx9NK6rc10fUuRJXl5Q+bqI6ti0QzzWioiOCg
bOHnXXwH3di4Jt5zI8ll9FKpNlYsxa9NQeopfqA2SQzshxhGOYr+M93vgvIJVAMcIkPDBY0uucAj
LQwJdMZD5n/VAtCdK7ctRt0sDe7xZ7n9YfqFr16t2Ek+ejUE32KkzMl8DVtbgpoXjx3mycFmhSLX
7kOZGJF6ZLp8Kspt2QHdjo19kH2568l/vUx9msvGcBZo7xuB1t/yx3N8BNH9Nj46FZkmBYma2sGB
i990VSPzmoDCGuYTTtjlpptDqFwW9QVBdkA5KTNQ+4DrdvVRMejDQXE7xGPEulD8tNV7pZVjxvhp
mRUA7e6czoJDVusT78xK3V7iJpyi52QEcKFhmQ5uhv4kcznjFVeMhpXEYKhrigPbUI2pEUB9eD2i
u46yjEs/qCekzkb6zhUtSw5pTG1QL+iSmUZiSc+aonOUi0C+iQasPf4lyH8lT+hbBgIx6gub3YpE
D17wDiq6ZMuf2gB76XUQMthwHR+JuXUO1EvfBKKi1UJHBcbBkmGBIG+/tS3M+z3UdWu3ZFY7URaw
BX9em3B1YjLW6hDF83UhZ/6LEbBiHuE/jGSshfzaOMClbrVYq9E5QlSl77HQSWOMJ34eXNSYQSzF
WhHt21FczMY96oXmJVobQOj6qWWjsGojc0QYAtkDVwkomUXlHxhrN3NYQqlMb4BOXPn+XoBALHx1
LOMbMe1b/FrELAktjLd7i/9nMHvDUIzvv0HEYifzt6pDmgVytGqeVuhs+aPh6aRWYC3Wrp95ygNw
4D6ucODH4575roitNQndMECXkwIjwp8WOqi0dGNEbXDyFXzyU/acZT5b2O5OsM7WmwRiVAoB1+Nf
kXd3NCWf3Bjh3vDafEccKthWefPCgXJQ1a77dWSfovWzPJVeCBqN3o3wpTP8ce8894UrldPypYo8
MTadlWxIv58wpeWdiKuP0JmViWBGjPri8kKXkx0ULaFAKr0WVVKXQ8Ktf9PkRKJUKnEsCDbyicpp
WvUQspO2xfGMn2rL066SjQE5YfvICIZRhPEyhR7FWV0ha0q326hmt6UwPgXUR5fAThvLStZL9u2T
1ENNjHWUcIJM+L46Gk8dZKzO3fI9fPJq7HP3bVKmp3jphqhDEHc+b82nWwk5sRQyNhUSaAsbvrCQ
5zmIttUAehJw02SNZ907ZYI0UnM7JKX+C4+rae6r97jJGPcb31Vi4a4fSssv1oe11Qgf3+aScZ8M
ilGKULfKPYEjg1+2L3LSxXcD9Jop4cB/AS663DQ3KplGGHSs0WpRHz+127/n51OXdozB4czgbHSu
0ZvR0JtxrDisELYAk7YMOVWBApOsHkzbzOwVyTLDTaCdE54nG2GYjKCSDciG9jzUAvitiITYFVM6
fwX/T2D1Yzss6EHAANa0VKYnz76ObgX8epZ7nrEtvdNiurI37jC6RY6DGYPQVU6dwBCYMLlYF/ut
RsN3SUIqAiFcBAGyOQOpzAzNJ3r/NeIW4Xj6jTzDxFsU6TTGbwRvIk7PUdR8XlLZoRdmnNiSPwg/
9zSh484enmse/QSBDdcjrzV0HnMgYWn+72ORWpiJ4GYpj3bv3SgxDAiGhAH4BRre5EHEuVXI9hWD
wWQyIPnuUGXInpizXVJrDc/4+0v5y8icsBi2Z3fkxiIEuNyiG0fJv2F8we4EuSRIKz8dEFTNzDTZ
Z6G7jpg0O52jCj/NpY/GZlrs/GrwjjKjJDQPbRpaH6K1pBAMk8E8AGtvL8HJtAlVMPrJHhTdZn/W
t4sjmwm4SERYri8P82lmiXn0a3VYWnLqSPPWsDWHazFt3rzRQrqz3j0g5aaJQJCBb4BikXwvVFce
4u5wV5fdgrX4CZiiEedLusib7KmjrKIBVAFCGWQgg57FaNs4ZYqb7m1NEpn5kB3THM80QTFnWJIV
jIilqATZt1/t/zmiObxl5PIG2CdyCHL0xoXvzsaavl4H4PRjtirQzhA29sKyb6fPp/etq2Hxavdk
ShnbzpIw/6RhfXceh12xj4Mo0uUS+ofAMv0GZNJUJZ8vJUrub5a9wFywLX5fc53V/vfCEfN4JTM+
edp9NwOCQ0a2W25R3ZHZIx+MNEb9d0mxY/yiMtYM9IGCTIF0ajzulp2kqr00qSntr5UhX5MP76rS
qIaMpD2ff7YeAVlRb6DcLh5hRihcw0iMA2Fgg79teiAlbbcCrGFuCjwgY+yUDXlosnQgBANMy+zr
fCoxTZ/uHlF8Lul1JEXgOrkcmxCQKDzLlN/AoK9mi8idNBnt2HZ/2DxMlP6XUGx9owdH2SBsuxl1
zr4UXdY7+QHNLhR+uKml/gCxfIlr+40i3DkitcSxMLGVdZQrLdQRk3EEaFz7su2+4kLOg0oqZIp9
/0A4o+RJFM2trydDf75u9FD+1FeAFVdJhQpMH1xnL+BgwnhTXD8unQXRf0xXOfk4YKsNqZoWIv81
2UE0yRBlXL1v/HIUS9wAh8W3L6QQdEby4p960Zl3ZEO1imkdBNFvGu5iVEzHXTqSlUBiMZ0qnqXC
GfXgILzjy1WWvQChftQDtpYpbEfQtY/NeJNVN5HQmj/oYLnaR+jMHBMkfA+dWDbJE91D9KyRNvDD
EIQ3la2GQgx2BKcseJOJoz8KdSJSdXSYybG3/3uE9wKwnn1Y6Nvitu1hvPiEzByZC2nimbjz55wF
sT29lrqzTXCs2P90DxV5xAfOCIeKxSjWt/28DUXrRtQNDOFqu3kO9Yz7BmpjmB9d/8asDDXqwy2q
EGUJQ/eGaNx0X8Cp2/d66aLbXa9WQhJo2ZVLzbfyURpkFbEWzih844FutytIHDeJTlPn59ZO63Hv
QAFjv46OhLSKn2DDK1kNiExtJgT11UJTT+7WADPdmQ5CAMhyiscPkWnbiXqrklM9oS9ryx4yoD/o
2bU0WGuqRKnpLjWyvjd4maNRKTnMBSk1krnMRmderhB7f/UEMBzZnPTeiveZvN8s/l/oXPTlW6iy
Fw4IYcurVu/fWhqhZTkSvKFp6xc5FXY5AXNm3aeD2e7bs4EwZwmgHSYDSavZNQr4aDmQdiu3qZ/e
daGkMRGq8HcEFN2gbiCjsDtHd5/0c3zWD/Doiejot/nmYVmadaqZdh+ruAMZWJwWa2y2pboukyik
3h/3CWhto2uCMM3CWjOD6KuBiMolz3+nLwzoGZ4yyAfkhEJD1RJGGlwDLcPa2cUEoCZsPvI43JtU
quRrcZa/aHSOqAIDUDyrbXw0dSSdShQNYXt6Z9bNTbmv/wfsx5iQY0IifzJ4buUa2o8ivIK4ZYkr
6OfKS/I4eA2rRZb27TzkwTrCGqwoFrjOvPvVnHSrT94f+tvpMmR4VNi2xQsetNhH+FtQj7F1dK0X
UMbq7kwpJxySp4KwV1zZn72c3HArhrxfNXuUO0ZN79Kph9OMUOzjg5xPErumIf9TjBkgtmVeh1DB
SYz/jeNtj71+sfG6Txl7oSH4wsM7a/H11n3pEbIvcQloDu/OwhwXUvXDLFKEq6Vf3LlYTkMPrPvw
D7gT4bg+ukk0v3foucbf7T182jFVgKsF63Du0A3Q8eR0UPxtsC7+mP+mWOk07kbWoBzBLSXS2Ft5
v6mh1L0HFQAsX4ACoqevceUMcpvl8nhAMO1IpqMOc13Phe0snvbGQtXYXzMCDS0qO4EEkwTXD3cO
mvxldpSLgUmB7Lh6ZSwU0b8fjRwcXZuPDGJQzp2z99gPNvF1aI4hnXKkFjOCHkqMMiI8a0FYOt+L
xI7f+dOXuDQJPTHseummjsMwUpDHlf+tu2CyuDFr3Fz05tvhwZ68llO5wUy8/7hHVlG47nBRg+0e
W9cyY0n+8gMU4hFGsUr4YB54UaUMF7dmNVNLkn5K6rFH66TgEJGA0FOa9W8GO4JZPLXzXoWNCI7F
wmftfilVo6hebfNF8Ub1s1g8Kh4do5lVlVo7tG1aH7wuyn5P8yuN4ts+k4+BX7RlT8rUKNv2iRnK
nimzfkkpl6DE4tyOjy+rCwyIN1CjjTMxqwCwK9cr1p0jMPHb7QGsMKVaLdTSceg95/j93jSndLSm
dMXAoOSVeCqzS0ofNPiEgQ7BcZp3fWVy9ctZDYcgaDTFymeRIjiv9gJaFPaW40RqMwPv4SXdR2F/
Pb63xeyflTXyvwmkeWvwefOGziT9MKdVI5QywJUT/A6S3taRd46XMZb5v/KfQ46woFNiZCgJQAeC
PdlKDSI8BJwgMsEgg+kr8n4dSZEGcZqzLPHPWuEnXxIk8kR0hM5QhZ/zpZEPBl9taSjnfriQFZWo
xVov8bhWgeYSawzEuY16bcFdDgtkPj7XD/3gOlwZbqpQXb9aPcUlfnep43uDg8vfhKzEgaKdGOUZ
Vfa6a2MWKYztn9P/97Ti0U7HZ9ukIIjsvoLq/pl66M5cMF/4V6b5WzlmsZChIifkbL5/yk4wZ9cf
a+lnJmqvhz7iLZynSoPfbhZ6SboDZOzFdTSfixj+TQuUHQlr4e0rjF2QJuRKM7fL3nGTlOuAN7GW
SmPxPhcC+t7Ja7NSyvNxLmFGar2/h7/xvrKqjuQReG1dcUpnObJiiKH4atCI7yFQwjdbLJ+KlgXB
iL941KIKzX6V7ZsmcF9h3ZBYzCBg2hJOtfDNCrPFZIChtvNjyC77nfLf7f19lCTEb2gO0/rDaO2C
jMT8NnoymyVEd6f0xqBeyyBW9FNC9Qf+E6cT7JBEr2yUNUnO4g2D/OYnR7XxThyIBReKFQOP+qWH
y4l+MbIBF0A+LU4So2k3JgeXIyN5AN9tLbnBWKbwhvKcglH1OywYP49tZ35r9pNTQBr5JWOa6iZR
8rZlJ6wNRJxoVaP0Fs2Q/RZGa/qnmlSg1JTQLQrpgX2LW8fcDou4TAYoTp6lwR4jSpFhQ/73BKzD
ePi1/XQM2czWLmvlz66iV/fYHzTvPUmtjYR5fj+5DCfkwBzpTTugHhv7cQayFN8SRDLWkCms9AHh
xAZOiAbBV7T7MU7FIHmVY6po80njUOTJPd2cHV56/sneS3xQfGRG6gd9Q+kO6fO5VfSFTfpvQ+zq
xZOlKLCc9ezbRYCk14UouspCMAfGaJOSenqHZzeiNkWHClrPcHGRHK97Tp3nHeZDavd6vql0uw7F
4/uaz4gshhUqTigd8jw6HqnLN8EezfeyVnLqXzIIpl2aCjLnUQiyZkTCzQ/zvxMSy5x1pusPznN5
3Lxhyf4f4vhNdBRoEcazt89CSz+yGdEY2nRrHX/ieziCpejn1IBIFgZRVvQXhFcwOHNF3UgGD3fu
5VO8KlnQ1ou/RteW7Ah4ejHMOLUyitOcNinInzGdI0h9DgluvxbwAcn/DNzPv8ep1jtYG+JP8IVY
mHHchJT+hbYW+kKu8cVWO9ZwpmLnJ0cgsnfuIk3YERDMlsiEV4vCbMAGVlWYHpC4JmQ/ifKwr9pe
xNo5BkJ4z7rLBnimJcRkNKfoXuU7sn7Ul6EAJEnRceDap/s7gN7R87N4zbbCTNGPSeTorSKkYKCI
nXyoWqmjfibBQgeYC2Qwl9h6xiZIe+dQt27ym2vG74os8w8md7M9q9BxLeU8+0CUVnCeE9Q6Edev
E39K/LcCQT/3t+x2i330u6D+GaHVtTSSGGvL+BAW/ZEpfZSZJ6nW2GXksAKFB7on9q9GU43vKggS
pDKbKJpxCelt1jibCpAQEABZ9cdzNQstB6Lf96AJS+uhnA5XgIfAAg1ZE+4TfjRsIErZp1M5A5G7
jYJf57QX4etE9NoWCg6JbSzKyv4k4/4NQnpcdogI3+/kEb7Jyu+gZQRxtR+uLggaQbz7Rl7F6SrO
g4mjh4q26Q3jS1bAn5GLup5ibscE3jEWrDmc4JyjzkLW7sItaz9SpAFUxvS5ow1G+1QzkGwGNM3m
XEL070eQJeKVsVS3w3LGbza3yMp2KAmQAmTmq8kd9iraV2ygskQTSDZS0hf+mdfHAASlOIRNcBIk
UbSxntzlfP32iO8LWdY2iqvwqeJO3In9aunUBbPpJqYaHbUPR9PFRmQJvzgrl851AkW8CwPcB/xD
/p/lWdayVA5BgRHj2KUhJapEx05OSKs+GNc7RFB/6KkgIEQ1TxvzPMWYRGMOdov3IBWaUmbvezRa
em4TfYDiDWTejLbhqx6Z6TSTV+rwOjJMK4wAmKRInWFmfh9HjP/X3h/AOQad8PFh4s1Hhpvh4FuF
Og9un3F2MXSDNlqZv0FVPvgiPE10IsdwTWjikv9L6KtWVvjWa5c41mWCWm+v1FYkv3Oc7qlmXKj/
4un2utRhYEUnL5D80OmabCVFpYF78can2vpiz2IuMAXZ26ol8fJUPyhIm2qP1C9EJHxiNSLNF/Ng
9LDNgEFf8UBmKEj4+W5TKkShzwrevlRXBei/Uj5uBvPMDM/kiBsVN3p/BFXiSB99VUcceWNd9Gtr
KdcK0cekYzZBFVRb9yXOdeKxjUqIH3JWtnk7qSi0JQZC/dF0bP5rlvnJM5txhfbcQNTR7Ec76H+X
RnbJGO4Kx92ZTm4sxEXHHX7vIQSDLd32hWzfju7W46Ed8vqPTJo4EYSAtpTVSzJFHFCzqG5s8SjL
UOkO1IN3Q5zfnwjJJkwPsIdCO39e1CzoPevUpzaDZ0Kfiefb4uw4f7YBo8zNk/nIeggTTQGuO301
nXRkVwUWbmVVzrCR6AGynk8Qs07gqC+1MxhWJni2SNjdQxFoGbsDa8kkBpGt54mKMC6Nkfz1BwvW
K8Mh8q1RcuFujFuhthaP+7pPdoEV8fmjILHH85hK6f5fMGQmKgO2isBKlDbNUBfoOMOQM4V2TZ1t
edXNkXIyyRPhf/tw4VpQLJUblVFHCsYyho2DKmQ8MDH2Er0zWUX7dyyTci3+VLWSB5FA4tPJqySP
xBO+2ZRgwdk185Wg/unKj9dJXbkJUoojqX0q1Pr+KvgnmEKFuao0sAV9tczBUHdXMmXBmF4ahhjv
/P8zFFa41Qhe0wYpKC/YJe/zUJyYSCrQXxmL6eCU0CxhBeesXnT7aj43DQ6YuvR4gXySiAiLHCjp
Bj1dT0CIsgz/KDakYrwXp82JJTDWXI1AtQqBE80K0NHU0Ew8aYz2P4oqi9qiUAG8pUyThCzqYnE9
3DAFjXtjtSy9YXK8lDI69M4heeTndX5jvsCmDSKuV77b20dByEUaMxcdDtHG8o+Wxy96iUjTmhZO
HrBWt/2EpBOn3BeIbMBgCyMwVgWQaxW9onA5l8SKCLbKbGHHTqR2PYiWVgX/EF2LEIts59deS4M5
bkLBs0by8DEcsY4CUQondXUtqZqZiO4LpNvCxE0k7FC0byCkGikQVGNBdVtW851ecrY2ozmzVXFO
n8VOh/IUekN0pOx/Ylc4y5SWsnK1AJecsIrZstTHqPHacoCzsJc+pvo0fQ2m/qGNGMIwHLu+TF/5
VaXh+BuE3B7iz5pv+Wa4t5H0GjJ33hpYskoruWeNEVLjYXoy/r/+u0d5hIsUFk9lLQJ5lM38HgKO
WNnkxyCmIMC1l8gkTyyvXewIyRhw5o9nrj5Hj+qbXYU/QwzPhOt1WPieEewD2wbK649j84c/EhMr
bAb9H6VXYl2e7AMnhUDwpdWcMswTWz9DTcNBNMEFD4iJYPRID/KhOwBaSfLrk6gwwQWtbb/Y60Zd
YLWmLJcQ+czF64PRjHmpk70qTVpDRSZbgak96uE8rAB5VmXuAqqQlQGAebIEhrgOG4BUwSV/Y5cd
VBe56NPgthDOgJlsJURB8lOG74bhY1VyaeSUv0liPmXjXBSNVlQ52QVR4SQKraAr1CsXW32Z3FI6
8jXPk8XVrByexhyAPF1N/tYKOxItNrh4IzjYNIPExdKGie6K8kyqx1shxlj+6bdWbGkEg8tLDgps
TWP/up3c02M/g5kK4Sae+qLkvVQiXTanpuazSZXNnUOVDfYVyesTO1ZK4oi3pLey4BGE22Oi/rES
D3ojR1M1WUL/PZr/OtHZbq5bn9XLWHPDOQ48QQaC4UIaICtmertpNsV3GQF91Nlc7RgWV3+loORO
lpJCoNTPPk//9GCmC22wLqFMEhZsqdA2wD8PTMEhxVdZTY0cSe0Uszchg0cgKkSIxfkL2LnCFzMQ
qqvJxKlul0wyMJRN7VqUAtAnxYKhkBpda3ap2o/aAkMO/8q/DfXg1s2lWUOargkgFyZNhhUHcRef
aqSAy8K2DSDkOyQfJBZnCdcjbeXKd8xMFrwVOFkM4ZyHUDWtUniyESDsdmWDYV23VDpxZ/KWHa9S
At1P5xxhU0ZsDHmCqp07Ab8i1svArMr9Z6H6MhcR7iiQ3DpFdeNIvIlQQcVdq8815f7gyX3lQtvg
tsrEZ5obl8BcXL4Z+yknea+VPcFRGLOdm/POx0bpgob5vn5XdfGRja+UephEL672Rp5j65uZulre
8E/PFKyaoUpCLmAZw9GGquxC4sPqI8VCjmg+vWuGJykrMEamrMwIMdVYhWaXZJ9jItf1NK28JLdt
smqKXVatkDTLOuGV0L/GBjT6dQzs9/VjonpLiOJDXaupzcJsKwmfp/kVxqNu8l73gYFqVVXUnyIq
HttTz/ZVYBswCyAEqv2VN+qgNhNTRtQic8C6/RcxPqoP140JzCNMAE+fqZH2mq5aeqNM9zKa7tXz
4skgQhByea8NNrQ3aA/wjNNHx4qsUD3iTqr/Mo5cH+XHKt5K/Ip5P0bmtCEIFeud20hBt1ouvHKC
tpFEZYqBKXdDvHN7vIZct+2Ni8ojyf+Vb5T9ALiWmM/sAe0lJfmuTGlxXocpOeePC+zO3xCYUbM8
Nv9Eha3HJ0s3tHM7Ag8MvBELVKtin/zPm5dNL68yWH/035rcgIUMrSQdiMnnHzDYL17Fmq9l6xX9
v7PgM7ecNUhkxBGH1fe7e14I8W/Qdr9nzrNGF4ITkMFKCeezRxTH8nK9kINw45QovZaT4oqLMA2Q
MFw66slFyEWzu8YD9GtvsRUcw9KZRlnovFbLbmFJJkCr6vn7vGUCBkON/LL42NEzfFizE9RvNVGH
/v7r0j5QydwdGLZWTqT7HZGoyCT2jVZUCwdDYHttLLZtpqWd5GJKETZVH5IIXIHgDFykiFhdlRMW
LIxEHW7YO+hhaUO5Yygh4kawkasPogLz89l66skDeFeZZXmN2b/EwqrxDg6SFg/AlN26VzpPyREM
XHgz9QGdWZAIlDEStcnMPoBMbz8nJEkRKVNRzZff8eQ2ncDAS9FR22/Woy194hh77+6637Gp0sR+
85AyqzUa/AeNdrlkXKZGvMReBsypWCw4PPvfsjoAOl5cX2QBNKiZWkLoTiTfZ6D9hOig+89i5cL7
Scm6UbzN/o7p5mxlJS6JjQvLc2mJ97ljPxavS8d9l3x4Z4679VTi1mvlRsJNQQ0CXgrkfOR/OWxv
m+z3xEKCVGPgmvihv+l9GkwbyMhb6TFNquzmrTeIJ4uROoP/TqvdGstLuTtwKv1N5OtMGK5qEXHL
qsTkh8gaC0aBL9SLZd1Z4IiqNILd3z+a0OjYxGSqKxPLHqTWcC8y6093SO17yOFC2VFb3rbMkkPu
8QIOx0vdpm7FMuL5mfDbXe0GKpr0GW8tWzCCaXPNaOAdH46NXW2LZr66RfklZWRaiOVoitgObraq
d0quLcZYftP2jAfGWWEsd5ghiTofpKp2hjCv2mAmEvCWa2c4NK1/r8mNwL1WEtfzjs8qhRiyAmwn
5JMFc/454IRYNgIBupXJVorlbskNPLPr16hKG6g7EZPWFtpkxzXnzSESGxXeAL5s39LAxYFT0IiF
5ulznalUvFpR4Alkg+bVa+R3RauWsudhAoeEU6IZz0BEVa0OlY7JW5kjVGSsBxxAS2R1SAiN/60j
xp43w7tOKimyxwGhZbjb+pT+uMxtiwrCPk44opThZdo/3dnVAjUH9+48XjgPkew+qjl+iqhnbJKk
jf+MxBX9UcvOtk1lb+rFrRndMtgUnSRr+OVfb2JAsaajgWBS7oqTFTqb9h09xezk42RBNSGLMeW6
WarTGrP0qvRLz90/0zASaC1ZtLPG5ChKY4H3KyMpxccRJ4X2Q2qOs4saM54f2AjgbEBwBvupatYP
8b7eeD1iIyX271h9e0YSvKDS6U84FSAwyJslKEEtsoVXM1eNc82IkNfzqJO5m0PZR+MqiBPvO98i
rC8m/KCqXXN3ZhurFKjVzUXCtd0cDpRBzKqrSV6VNXyeUT0diDuzBQEM6+lv92Gt9mo5vmmcCk1/
AC5bEgU6rvkEpAkSglbiHgLS61i9xY0XkZiAQGBBWAnc0p6DxMfJW9+amO7GmLpD13wO34CNBDCx
GxIGq0o3vTD0ysqyggb2saxP7qmELXAixDOj1O/YwBJ9uavxmtvfaPs/zWJQ94xs654+0arDNSS+
GPLDtskJBUYi+qNB/L1Ya96rM60j8TkE4zJIPgB2Dp4BpZu6SbII1BrX1I5VY04ybZx3rYnCHIGM
4cGb9IovyZ0q8WSc7WtA5GRL5IBwI9bTCJgKIx/Mf1Faq9C/MABrcJmQzZQ2VsGOFQHuB+UMpc2C
BKL5rDh7ctZnygkxNproUsPjBHwQOWIhJVEALPLkSd2VQAjedLHvdSGSFgIbLwOzIZimeuQ2YWtg
Ic5db2MlHhGAgHqBw648KhuCTXQDI7u79olMDes84gaG9ilN38yuoGD9yjc5ngKLLPdsC7+6yP22
Mfgm6/ox5VLTnVF0XE13a78JO/6fmPydXbVAzGtm8ecMFL1giFSCZDI4bEAKn8z1ot0A3+xZc04b
/cVw+yDpqaRXOCyhpE1CtyOjrgjEdVN3bI4vDNIRYADvfWDc9jTN9u6a/QX5kosL3NnBsRouVZrl
/fBSTk6J5n5SLb7bM7MNA6XdUOjRI273Uqzzbv0wyEOq655TNbfCmfU+7oNBxzrvRQ4edH8jGSTF
WvP7Zo0+YcMJZAfMVn/cW6zz15vo/o/EwG33GC1fmkgXOFyG2C8COY+vghLTkcOKp4AxLolrsnTy
/6DLu7+QRME96BCqw2W+ayjLZ+lKIFm+VL37/hqt3gKKLvFXyDjQHOLvQ7mo3y3K2rWIt15C6aSb
7hNsVIhdfPriSQAkeh+4mO4Lo22qDpvH2o9X7Ypg/1K7SRA4iRe97gyQdRm4kEXu9aDrHJ3bIUbM
jvg73FUI+uKgMuoHuBxkWLO1Dn/yON8d2t8wR/iOOtSybXWW5i2y7jGcfR0seF2IqmW+3z709OXK
qZhNscKif3X0Ei4XhfKKRBWXussELsQZcsQdkvLoRLM1eY1LSEQfTRVfJPmeurMOulQrHAoX82pB
9GNlhpdzsBd4lXCnEcWriAUy/cMD+ehI4pHqIG570Ry93z1EcQt7lv0c8yAtPIiDpp0Jo/d79zbb
RwNzVstDxniUHXQ3+LGw9xsbOd+l+n5bwcHpqPKZpccT67j+pf7436jd5pIETeGwCiiaWAe8LUkh
Mcq4cUJHA3dpvEzNfb3TRDSsYJvW9MDadnlwiQ2waMZBfMUB7xndUfbmvQ0cdppuP4uaIQaC5KpL
H4BWpdGED9P3UkuconI7onZv2EoikeTlj3h0fL3SdwTpRJjOHs4N9DK2rjpsUrUN4h6f6WhOv6jr
gMk8ImHlQHKOP1mJNNniUyM2r1J4CwmH1GYpKpUPIUKdJxFbg/kMW07WqKxdVIBcnQLxKAZ7OA6i
JLO6ox28K1ajf0r+4cB1S2A3GjXNcTdqd0BRS7HYBCUYwzUzY8CpjCHuvViWqbotxFcaZqoPSweZ
Wh3x8rmVEpG0OofVI1RekybNKe/EnDc0ev9tx/DjchDwfpWhr7CGZCXHpfVs/PwTfg6byT9qKeR9
k40feRqlEuhAF/qm2ptq0iIzHQVJCZr2bw+a+Uonf+Y/UwBZsEb/LXsp3eHA7Pb0vmM+KPC6HCM8
TLO/40rrKS9nCq0+ftRm+LaGmkoO0lCjYOcvws2h/hiiBHAdaGpBQPi57DkqKcpQd479kVAJkINL
Y0T4cb/5nDBqIXWNh5L0ivwhToPJORIwk0JfFIZ20I0JsIO1/0nRTOzPDh9upPzgoXxb61uyeIB2
RQ0fpJOwLP8QRPu1DVf+JRiGBsmSmNmtR0ibH10AL7M9TgokcERSPSHXa9hWvINbeppRR+R6IwgE
1riWC+PecLsRxeFDby6VD0QQ6ynPDYvIn6gfaV0S2Llaps+SeyijqAPJ3QBkwSBIYy/TrwOH3z6p
/OEnGZuMw52yT2k0eKjJNIBGFTUCd3J0teNdNdIX7gMYzi9DoS/lknE2Bgid/5+J8A0Za2qUnf7H
ayuBGImJy0mcD7CgrTdmfXR9T2BGmmuD5aQQ+Yom8TnTAXrENAol3eW1ROK+1/Lt1xtmvFp8HK3f
UW1Vi0U+E3kKxuy+VBK/k7VidJgS6YNIfYtIGATMDdO+CUSdTRlAu9iNJR4QTu7fd3Fv8xJdQ5/O
gKvsuXyhwkv1rSfzLdG7nl0O/c0uuJwKnMWoNEaQrfEwbKoB/j/ksbpWFDOe/z68YQkblYCRbD3m
JSplb6wZYBS+pTcFf3dwU4iA6lih1Pj1LRoHr9Jom5F7TjLUwKRz59kHxhIOb/aWK4BoXdazVMVs
e96hmyu5b7jr3XF2S3ReLeCt7O9FgXemxBDKTWtzaHHRiO++fmaSZRxqPSvgw5KPFMGu2bVsqhgD
4Z27gszDG6pbuAXXgJHq6+jLNqdG8xpBc0zx/lCbtbk1hdcs/r8hhaL/7ZI9j2Cyi89PHabSiPlu
8VJ0eQzSUZ/Kz/hG5p0dWkhx+naV9lP4UNA1gduCeTBnz5oLCggJn4W9dB+goT+h10VMM3VRuT/V
gTUZGayvRh61ncBe6MS7czPRCgRqx/OKAlGEEMJCBP10FqvdepIpU9IGB8ZR9UetSete7N7RAKue
/8PGaxb+E8qlUR9h7hJ3d1X477ULaz8GR6zTQBMU6yBAbuqGast0kebNynzJ9wWRz7pGmkdZH2jZ
13do8Gm+7ZlkIdvHwYuuN+a1f1xks4X9YZV2tcZ0/2j9EbVDaZE9yG36fGO5SDWcthdFK6ljAaRS
xdKXWfPye0DRWnak3r/uLWWXM8S7SgQrTNR7drmClzKSEAAKdtQiig9fEqzAvzW7h/VV44QlVoqy
/szn8rHK/nPusNo0nUYP8b3GimpZbQWdo8uPMIvBZsoHGCewiFpmUUQW24eaFx2V0yWQ1jw8mszQ
iHr6cS9ZQgM5aQTFU2lCgxJlaGPbNJs+VY7+4jdcDesCmDWnVbdoI1F0z9MYrB8eUjshZab0SBrO
dB0ZhRCEsMqNIUqQ/v5EhDXyQdXlwDFo/nGZjO8+gaqi6vgNXjku93tOUL091pBMbIqO1wQoz/yZ
7p0Pye8SP9xKhFaLDnTy/XjpY0o4aW7H44JtwnJUe+j0amgTfE7cwPZIPWokUBB3cNtozzx2WI2y
F82fEqFb0RtcC9tceR3pRT/wE4cgqVq5FPijdsIsFB/4n5q8+KdfWjfvpMrAUdbFddn31VhCoUGJ
DrdknhwOaj8nvjQaiO8hbIJk00jVSbeaNvHeydRtugtmCKjLAahPMJfyEMXwn/KcJuoLwJ/YChyn
fD2FGUMscv5Ni9e4l/FA2yTZ5Mzz4Mn8GwqRPli7Rwl7P8rYe7R9h0P1arG+Ny7Fa/4guyccXoAd
B/olS6Hz0cAwJaRBAYCspmhN7uczWq3l4pv/Wp1rxTf8EY768/w+yzIeEg3aVtfMxGot4gY2VMKZ
pmq7ZnyN5Hb2q7U9EiR2RLoG1rprkKaJu8Dj0Jcb/iTKSipIYQezSk0WpZKKCaramJ6p2EQmKUIv
94p1Cirs2xsnxq8xtQTmrYr1wm9KeT/AOAnlsuG6cBbw5gEdF+iE2R5TxuKQIZ8j4NQoTPvkZ7ql
PIzs2W3nLaUllzyqubhLcQLjhX67W/aMbI1MvJJZsP7YWeCUFUhIK1TcYX3P5YE6XeDhBv1UPquB
h+Zk+cNwTHgKJuseO5GI3LBXZOZrLTx8hyZOLewKeKiU7B631QYKVqdKFBAiRJjj8/9GFWi80S7+
NypFBdyJkocqPf3G04SAOn0/XW568N3+nEm4eO3vCkRD2K/C1MZeRQiBK3OWNaMTS5H3VXKJcoCx
D5xYyfRE6VixxVn7Oz7MM9d/v72idSF+zkoHZle3VqihP99x9S1KsyPiMwiFON6JBVqtmCGzsBjQ
+PO8NzS/UCV16zF+A4bvM69be8c5GFI1jOmCEi5qiihex/zF87rDg6Bs+iXEezPIiwIAw5wlJQFW
CPP3eh8PiCfo1irIWzTPrjivyiAAKDQFgoB41yY5l27JZGdaJktiNatQ00R3Stg0RLwLf/vBx+Ow
vB4/KLI3jtrF9M67iw4R3s2yLM33nXtAUMEQiZGI9OOds1UoAzvBzcUYkzt6R6LMgLhAzq5oc+Oq
HM7jS5eNFkPzPIfxN27CB/oXGP1zj2RhiJjf/GqXKf0VZRiRu38egKmyRguag9UjDDouAEPFC9oA
BOMbry6VpCgKHlZ8xP7pMUUEQDmhXuGkberSSrJZyzcpLjZFefQVhiEB8AcJqzx4M57C7+4mmjMp
au90ZN8F1iGU0R3o349dWNFZDQsULNd4t+apLhM/LuVlGTSieDa5VGMjK6eyBsAYomrdw19s3BD4
I3f52sUcdbqUn/3U8p1d+A6S9jBQJRkDLK/HwBpVqAWGdhLNP9he46X3qugAm9kxTouD1t46g09u
e4DTf1wsNQ58izxurJziG9D7bNVAUwarP073tKj/a8X36E9XE/4GimBGfxkw3onGYIW5jj387nV5
nqVc0EJGOxyrzz67VRNkOwSB0jSE5r/6Qpx0TI698SAVadmNgR3JBDd3ZznB9+ddF0hfkqGryVo8
7scPwS8sACoUiVfrYlLk6ApEKDlPDjM0URl2wsoQtvfJo2/bST1c2I3NgyvccNPTf22frNYnIiUb
cJW/dAKEA12eR2TznZAYSJQDjHxlJzDNR5URTSr4gU9iKnIosstuAJhdeUevTsgAvzCBYUngf8f7
o4JpdO0VctFv1dJO4Ns5q7vJBOV+T/TsL5zK1ZM47GTXl48J2vZahnGBvGWDcwL2EA7yc0AsLTC5
CNBGAmtr+zDYuZK6j4mW2MxTmTrm4Vb/U+Kvwm56Y6k/afgTQ/B2sGVkHlWBmDFZQHtEN8UHFSoW
moXGZEG8EJN0/f1zBtnvCvMER8FZlGb4FzWMF2Gwfs7D9hVtuAQpUeKIYA8UzmjH7AHj7lfF5bT8
SYNNqNUgaZvrnLbcgnjCuKpZrUIKLrjCvRXeoiKrnQizKs0a0vtT30kB5FXbMIDIotZH5lRaptu/
8xc1IvH3TBo2j93N5Inv4VjNiO5haHJUh/WOPiMo1xkGL2ZruszxEiZXwNeMCS0fdKEGlgGuoeD4
+rciAh2133q28l+jFqIATKgnIkOU93opKP13MRGpICavfhYjHKwd2bzqwcfaJ3THgLFHCHBNYAyg
JP1lWnaqNJx+yDZFG7GE//E3SOMFasOI+TbtYATyVBDSIrYoImLxV714LYbZqNukiTTXFjlz/k8z
9Y6LH148g4Rybr/jI6Za0JTVAaf0qFIeW2A090taga709xyq3PPKsgKCRwEPGXEXtHQ1x2EU5E8l
mIFLVyeQJ0Osxqr2vQf4e+/egoKvTMEsDajaRDK8cSy5eHnoczVq0J/ZB4GtYLucBgR9v0hZ3F7v
/grTUvFtBtMoqghxeHbcKJaP1XZTXAkCoycPk+gYcFv2vmKh+fCwDhvKwaGeAM/+DFukxprUkZ6W
q0zocgkASEi4WrMpftRmSZOjpwhlHIRMEsH3NwQ5eg6AU9S0+0YDyuVJMFvoVawZZR0ZQXq2Syfq
cmNUDwqs+7YU4CeHPE065FRE2Yx3ZpWOAAYRnXz+YfkKT7WiI7W+vFANEM6eymVUi3pzK+HkGAw8
waH6911KOqThrYH/HxeWTCfCbE6z4kPgHj/ErvjxfPT2c/AGJzIjh8YTkhUwCFgQ9NyGL7HHpSYW
a23mHB0zJ+d6h9kNy7CFeL4PPKYWg8gHGvunmaCRNFm+uqyAJe013Kxu5VFKdXqADtz1QeL6t2GO
Bm3Nc9yFzoAlCkHpRRIwZc3yHCgwv92boexE5EV9GYgDyYeYQ7h1x4M9qfPHXF8zDyQG/1iCGZ4R
aGSg0MLEvp05Btc1fw/3YBcHeRqFkX+X3j+xXi0Tsu6z6xQ777YO/8/hgkXkutJT2NrpLEh6R5f3
l23ZDCDGWUW8NITWLL7KZGa6DyuXJ1ZSF/o1T01l4/vvyzKmtfwE6kMkbA3FBFCHU2wlruOWYabs
fFqvvUKrgIVRA9FceORngPoJ6cwSwYLNfPNpXWvR4HDRAH6jENrBl8uKdYbIW+US1Is6ge3QY2wD
trsYIcOvjYvgHW0HeF7BboKRj6mGqB2jDYPPHdPUAd0wmmuKwzL1Nlv7+LvVkwda0NNHbhF2cQuk
/bPa4C5fI4GTjhbX5KkNNSPwxHwQj/nrj1YKIF0wCuCUpif9v98KFc1ETsCG2E9bhg6kbm4VHylg
nK5t2ncDPaZnY6C7mR3dQImG7NetUjHIE1ZqN/TqRLmW1RvQWhRyh9DLJ90T1gFnT0cp0434W7qN
XV8zva67qZrR4LKNcbJfWrLfYLte0Ttedq4SRePjG0kE1iQXTtHRczHVSkJ0J1N4liTJhHO1N28m
AJgmWz40bnlPcoDPdbNgnU5YclvNqQKptfkznaLAtRyn8MjACYR4RhOrn+VMnZxk7oc1vEpn7x1B
DE3cHA2oX3yRmZ7JwBF8JpoZ62jRvTjsySk5UvfmQr75qoiQydhUlPkuctQRUS0jH8Z22YNG8tHG
RDmlb0VmZI/mZzkkDo8IaV+ZCm4X+bHE/aiR7DeN+OCZwtv5+fYwUQF6I512fBUaPFp9Ytc9Ihcy
L9V0Uj222vrDK74oyjDYnW8ini1EpiDD/1QHIE0Wy4w6h3w2d7/3rGibXM14uctOUSAXOU8DR0vk
EB6NxmvU7Z5EhS1tSijauCQzVv9hGuUKvVOYuTgiw0e0A9JhIuOBmy4sRnpcKTc2ZeMGDOgC6gHI
FZrNxhTpv9MGu6Q16Md5T/wm9POF+rR+B9EnEZ89YQPdnSGFVAOKevILrCe7wrlU47z7OCNwAiCl
okhUUlVfKFD8h/oW2vK5yqXWPr97VvtrttEFK/yj8+rchMW694yC071qnfgER9RWufpUH9TUKRt1
buw/fbt+IFN1BPRSSd1NH3ZHljgpuEINvWIEhNc1vxl0VRrMouiOOPfqCOv3QKVUJrQRgTen9fMU
FYPs9P8XeGZXFAjn893AAx+tnYwFRM1XlB7bHuDQurnAiuIco6wzA009LkPKI5ATEiKz8Ap5iFVO
nzvRl74/n/aOxXtjgHFoyOYWWowRX3hXsZsbtg9tY/yhGgI+07l+E16USleU4nYwvLZvdL19lfMI
QtoIEN48tvosyOobFJ4XMEvZiQTdecFbLJ2VT6TIr7O1b6yl0OXMD531YTeXlT0rwS6abvQlZNqc
9m+UqXmI+HYrv/0chxnE2MthdUPbnpOjL2Km+lRDlft3O2Xdsccw8gk2Igrcfu58J7fcon0wMqFj
9WHJNxOs/JdBDOYy7o0oca0SFx85ftdt/7uXZQ494rSdme7IPc20EhW1xe0TB/kV5AOPT/tosNl2
whw0HUan8MSsUIrylinlJj5LgYJBhbJNhQziK5EIADXcSofsPkHoVupbM9T+z2X6TlvqWcUtpt8V
zF+rjhcqxJ7PB+S2rwBs/ZXPvCxEpOeZaf8jbgzBCXxNMwT8UYv+sUIPXKA4EHIf+yn/z9q1ckS2
4w6JZP68k6FoCSXuGOCEuZbBgCnxdxc7BuBJmsDxvIpoB3+6pK+2XQ8/sD+e5zZaoVnlcPjpbPfa
DgsSGw0tKDApDMm1wveaqTFPB7NLMOVWLefWEc4EhYi5GXw5nXBQe3KcewhIz3anrubkEI8JBk++
iOs/lEQRnSuzRvIlaoUyInGFgxw2SH9qMn3OxTn+bTAxGOZlBTYyat/sEFyg8DcBNO51mqrDzemE
ikVaAOhN6dQCNkRwJ64tucmq5sw4+aY7LxqKlyVhUZPD6L+CKc0Jm81hkpr5sRGGRvxo7SzCqN98
TbrH+zVqZTQlTUxw+OcL7MejwL8E0nI+5SiYp278Qyv6TtmsrypTByNWrwRoPemw0nB9qGbKJnez
uRPdvJVIkj12zx3co4sRFXwbVlmmhOZMuYXokCTILgfXb5sQbV9QulvW3HzBuLys2skqok2VxEx2
7savqv7IOma32I5C0n4g9/ltsZV2sAsoNvgp5EpsjAvwv0P8Dza7PiDtBWkQlipszbVhd8C0NWvz
qVAL4j0BIxyeLJU9DTf1H31sU7zrtec12HS6tUjtMEYRZTB4tkBR0sjTFmI5V+S/bJZ9adVUDWIm
bvUeFhAWqH1Wn3zFK/vhdgtt1pRFaspaR+5IqfUMli3QC297kuvYGQvLw8ev2cWKBrDoPD9dfOUt
0YJN3qjxJgwhagwY+ZxPXMEuuoG6JQcv+pmdfzG5z5ej9oti1Rqa5jvHoUS9kO5Uu8lhQ9UN/hIh
fv+2/VDk10WqzADoxf5NdVG/UzjJ1PDreWGD06SG+EpY1kyKfgJV7LU7tpDh9cP43sys+WW7HOHk
cpcKEbpUgfELAI13lTkd5E/m8KDq9P4qhhPNfmWNIzYyDIgeCGxB5Mt9aAhvVka0GO5t0MAPfxIc
yYyoOhMGMkFnGsuIehIxJMaQKOJxY4tYe5zrwG/Y/sTcCETQ9QSb5Fd5aFFBTHOcf07rE0WRa8ZZ
FtTGELYXFdaSBpka6wEAYnqCiPtd/Py48grIWMQECNHNcth04kFirxVx2hcZe8/hsLYJNAIC8/gY
4Yw2pqAaTPUpJ26IahPwyvlPyWbTHrYi0n3gwu3rA9e6vfmQg8HOi0qVsO+xH/FcuBO3yaw9txxS
lTOE0hc8JUco+oaXaerdfrOXFLBL2k8mC5bXBqPEys8xRO1Cl4B0Ho972vAqQSp9oRKXYXdG3hHe
/GQDvVshMgUmmyckS/P0RSNsM096X3LShvFp1sqhOl1gGnNbhSQwz/3sjBpKCjAjqG9S/k47uM9Y
c6bFvuKr0BD1klHF4IM0TZ1hO4a89sBg4rmn9iF6sYMtF/NdfJYEQ/egwb/7GxtUUV83PyFi2hab
qcbHE8jbhYq5nBe8kwFggdo01B/zpTgI893e9pwVs/z+tpyfWTN6OV2Huehe9XJ9MQQCEPoPmXLx
CK/rVeYQE7QKTVSsh6bOHJPrJtFAWQZajWIsG3Y7b3wb0CyJMITQAuoPfTxZX4bylm1uUZRcWiJv
MDbk7fYEDHdWk9+4lqJ/T7rS1fLQzSukcwtmjaUN/SXbagJk3wzq3oD/Bx4oRTYDySAfOu71QaOy
Oxj07IOwfaHka9jJWlYgzcSnsutHQtZ/kIPdudsaNU13jRgEAzoF2xOKgHst/xA+xzSV88fR2Y7L
nZvVRwtyiMhFTglYYl3djo7FxEfOseBMJsVouw0Cv3WDuFYjIUPHz1EGWhqmNrIVjRUwBoi/ei6U
MeXrDT0Ivnp1yr/NHlA8+749htLcMKDUkMaZX1pyMfYqjZ7LE+fRIrDvsKT4HxwT9VtAB/24XuYq
IdfV5eXvWaJnh3QKE3fjFptGm0viBz7p4aQYtBVlkqy4k7uSNfW4FqHm7ZQvLJV0Jl/GhFST4atl
yGKb3HufzMajnpEm4g68/wLYcBHiX1VdtAsMZEZ7ClNLbx26jBl5v/nFR01lhfByold2vSMnA+80
95xbMlyCMhtN8m/bjDQirihXAC6qQXYNcB18WSOPbMmY2ibiBqWa3us13DKzTVui72GxVFnCLtsa
WEoscxrKbA9ruW/2edbTw52YWr4hhSUwr+ZgWw7x8yFtLGPbZFr9oVvf1rTNFwW8agQR8OFMGWWs
Ue0UOI2LX/EQDxXNnEV1kKW5u6hH+5C1dWMQcGiIp/IebeD9neBhLtXds/DHWv3+hMFIq4E5cPve
kQHdD5++5xWMy+BDLooA+vmllhjxBFDXgXa7ZeuzvJQdGtvAQV7effOKEzreIP0Ekav8SPaBlPMq
WNO9/JXDB5etheHPoV6YLr/wGQk9lxweOtuEN2btuniYh7TCjQLy9lhxzxEXprxsbTxWd8jM/aee
HfIvs+3QNpmSOKtWT/+Mc9OGVHWATd//Ati9uCYoAvtnCwW/F19GwQ5o6W1yJDazFvIGx9x4wFuF
jTdKiHhH2IR3fE49V7jgiCbf3l5qPEEdrVF61thZmU+D6Ys+9yVQNXbGdpSaK0s/22G60tDOJJh2
Xu4nVF5wARD9yJ/N/wfiYw30G9cC9llZTx2PVeVNFzgLj3VD9JOijsYwMVLfIWS8zjENr1+0HGqq
KN4TRTXMk2WFnsnAV11JCsCP1QRLNXlqZIettHY8NMzudU+c/gkAukmvpufTlD0JGJV/WOnGV2xl
VdcVJwxeCYtwuMc2klb8b2VKkGBmyBaB8j8gDSH0sxY6UWrfYD6uBOSm+wzCWQitu+uHyItGyIRO
BrVGa4T/Z2/Unjbb7nSODKS6jOn442tOS8slsMgkJxb7DvHkGAzjg/UucQ007puqEwBtDfJ+DLhq
DQ2NvMQ+rYep+UEr0V2kZvoxOG0yddWPTraKusuBVIou3RhJkGsjB9aJo74mqutVTeXq2/uYccw9
fxvDj8q19WDwoy43kHaeEkIwEarDfN/NN8LL3JQtr0I0W9BWWxGzvJE/r9aiJhjM7b6enlycJNGo
RYRCnfwF5sHd8IqoTVfPD0+HdxVxDA5t6ScxdPNYDiRfzDqovNBXXZPlUJpkNSlv1e8vcsrZ7Xie
z64MH2Zwce1CdziOnejFUxuGiG+79O/vnBrQ5IFJaMOLF66MbEm4OlGlKzF7kGR+qDytO/c6xpgv
7v4AvrX7VmcmrTwKoPGRIGB77rxL6LR6TifLl9jOEPCHIKLyjZzjZPFGsT/XMSvq4q6wGrxl70X9
EOntupxRHjLagtnKyHMz7VhaLol6tOqnyNkxOlllfQMyb5cNOZ9aBpNfc493ZFycZk2ZXGPDN+yF
NnA6LiO0oAG/TuNdivsPN518ElVwWxebs2CeQpc57EYQ0DJwc//jmVHJXwV7vm0cTGWZUuNh0T7l
1TOMFiCR7bQIPLPsoF6zMGtcjWxK8uR8wTVCCQVXM4F9qb0AzG+oU6koGtuzqaLDQdjAww0YGIzW
cgTaCSvq7c8atsTNkI6gamnjfcfAfSVDICzPfnn5AYlO/8g8N8KT967n2GWdhMeKfhaIlS2WDX1m
40AtsxOOz83usez1I7T+NZJe/jwKNzrZbwyKGqOrmri+IV5f7jcKn4uzKTlRdUIB50mgZ16sXdMR
0JSAeE9RB6MXv0mbo2khoQAJEzKeSMADpGcJWBKJyGhsSiv5zeKfyhxr8v8QZr/RKoigsGQ3Emir
05k2qbkiySzHy+We7LL9vKSlnIlSslzVLqdxC3qF3dkgzjyQnDAxst9N4tbptdWmU6E19BXOCfTn
7ZsSy/gQzsCw5Y47zZ98kKLXck+qoV9+0C9lnya7AY7nCWtonUzUYaex4rXCJTW+bsQ3Y/iZYey7
d61a9YH0bSxRvmJu+1mjpcBMv8fjfaBTwLbm3JfRyWcKjb13bPE/971zTkFyzz3MhuZRaU8QbxuR
dTWNid8FevGJl4ltdC4b7FySxUXWTQYvyXbCjwKT5+o3DXb9+4Nv5Dfftqg/QAl5ebiAZQvNCZsb
prJ68zOpF0t/0R0yqb7S4qWuvpBUUiTofmkPcn4qdUpl6wA1B1Lt+qEDJ/7zjpOPc41DyACrn6EW
Pz/LKeBwynPbJm+ZKG/y3DfECcY2Yn0vP6IpLvyOKrp9wd091p2vSAUC0j6IihaoNF+CoPW935TN
NoE0uT634slwzeQZrJmPq+QyNchF7S5Kp0XLrhe8seJ0ig5LmSLtYNYCpGaoq3Shq9OA9FDZkcFD
8UMEcL48EZMgHxPPFI5XMgs8GC6WeU1IIA48ADZBPFLZFyLJ3VsFBZZBOTCwPKPXu+sSdGwti3gT
ubLsohZwog4XcHvD99F5G1a0pXiM8pdMWDy4wpGOYJ3hjwOF9wTMzRmLmY+CDc4opXhlR0Jd5kZG
mZ1w3UB66Eh6ufy2ANEomCQNOJv7eXnaKrwfaswxCL5TC9L2wMB3jaByCSQKOYJZsPuImy8gQuES
VKphc6SvvLonBKeQ0L68o7eI+YlBuOht/td2znPRoPyIXgaPwcJ7ktj0v0x6qtjZ5OUCizmKBh66
y/zrxDGzZHbF1nxT8DjCumD/0WM+YNW4CjLrUprcL63oQWg4D8UN+bVLOvPVHlSNg598dtz5y//s
SW2/dk37ra3dPkeXXTuPa+bwbYscP6jAIFo0VJDd9XMrirK5HEV2Z65F7t28CRBSnHc1zzpAAqU0
5dqTxItkBdvBnYxadG11ZDLfPDBR7g+9NsQYWhb0XA5QuPxGHvcIchqD6P2QMsS3UOBkQ22mGTHK
XoiVRHgSavXoSdzWb9n48YyRqyk6vDsXUSheV56a3m7r2+zOBWJ6te63FhQKEMA/18YdNcV6iX7z
Gz1NZ8RIpzAQmXfcbMpFbI6Uk+NFCwvfSso8IACEMU2z1kWkyxp2ZH2yubB+hy7F9YlomKlqhjmE
tUjXpSmNkQLhycyn2BxPJLrQYUczPVnKqzz6a8UtoM2y4NtgAfemeii7+1pV+4j2iR+RiTQ605gR
Iutjx3RRhuFN5eUF6wA/EabEYRUbD5tfZlC4yFSiYRV2fk53/p42hRGW4j3fky08GS+neck91nYp
0cJ8Kn7zGJAD/8GJBzNvqYlSjf0cNyx77QK9k/M3ncskA7+vF8/Rg3XTxKDtUGf/9/rZW16CA/wA
e4wxCfY4uwid0pt5JtHrlgl6DvZCguUmIU1E6jbJMsqXYyFOVW60gPwJn9o2epByioYpIi5dmh7j
1FgIh52VYH12HmG7pIWGt7+tnUPXzhBrPY5ok4ON5tph7TzEzLJ31PYMPINliN2FRj+xl2Wh67tO
ZnvNioRXFsPrxx/nTfd3xhtdge5chaFxselTEey6uUUamtKlBPZK3so+sNKy6maM/MpvU2UvHZfP
T6c/ht1wdjzToYw+HnAxirl8tZY363J1AfTejvvEnMH8uErAfhF8Onsxat0LjZikYzyP5g1ZhYIM
Keeb2Wkyc6rGkrWkEadyPE4SvKF2wMAM1fYgK/0wP8Lsj2XODu6jN3+4uEzRed3yafxWXrBZduj2
2Y7OWGJfxNdZGh5sytm8RpnK6/ObcPf+XMoNKyXIjOBqV1qles5e6QAp+I6xlFr48DVVlRgsBpM6
Tdpqrh5AzQPkQkEVmg0pKhOWqxAxy7zQuI+J2x0chJau91F9sh+cKLT1vbJchiQu6I1SPT3q3288
RPLx/9olDzOfY7h6FX1WCY+c39ubDSdXs8occHqs/8gXEUibEI5uZk1xseOiZGtDm+b3SEVvLpQB
R2WNkwSUHIUuLm9axFwPhyyQuToQpcUTNnCyV1+0s1N9PUaMGxmB8BHBoR6iNcwF8go1NjJUyABg
4fVWjPoR85MilJBTFZSqwwX7gaw4fIgMldtKPcP4IK2/StqHuhFhEkSvnxU48VP0FeVdd9D03GRp
tP3RJqxN04f0U4e5/93FsvwEzEmJA4hamJikIWWFqhKPyjvs3+hXAuX6VYR0Wwd6ueFjy7Y5FFzv
kbxxx2P+/Of1LLsIcMTW6pLB3BV/Z/VqucD/tGkvGm0kFi5S9TGEesrvNyJlhdwLw1umeaW+L2t5
TacWDZ46mpWFNVbaQlIbQLO/EKSINkOuXALWy2TAwUmOEXNEYn8xbxwck7PeinAxLIDWAUbfVNxq
MPRL1JyFeTGdkTdVgPPxfQHQu93VHv6qs4qCY/+L/leFrQFJL2KDo0X8G1CHDqWFeWIXYCxQx08+
curp9Mvp/1oAAHUU3b6OfWKvMpLkyP/3FvVrKjFRR3pbnP8aAAv5F+Rea8V9ZoeIOPxVeBez1k5B
+qX/kJ/Nbkn9wwxRN/KPDybk0nwxZFBXqkBj+Du9PZ3hzePliCgwefPVN0NiNruzF1N0+Xw3mLyV
RL6NC2XDwDCXXGrieQQw5cU0DB3itPe/j8ayg2jJy5BF4l4rAXdaMSrJQAs0sfjS3ZVapwrwH/0v
nfdjLNxT5XFGzZyE4xeeRkgAlA7PMvw2wa/vUVgXqYbHqWFe675waJuZi8RSUa1YA149m46zXVTw
DbO5kZCT+93jDIAQXOC6OW6Us6XbI+IqmJDuExVKWqk7mUoQ8pzJ+5OK4UbE/QT3IHUn3lGJYojU
QOmv41YlRdZv1vKh65mKJst8P957K3Er7MSs/4h9duCJyut1qTHWwruOQuwtYHlZcjM1BeLeoeI1
mRXQxN8cCJDRM/+0RamEratuSa7QlYXVPT4lZd0WYyGyWHCi6b+C3JMixh0oaApZSOCQwi2XmLJf
LMF1CU76QV+t8aZQEoR3RJ0oruusGS4w2y9B7zpcXVkjiuRHLL/4sEpxRuuEKtU/fR6w2S+qIISl
Chdfr0TqdWWfFM6CF0IS/CH3R3yCwldwn50AtR3RqCf9Y+7IlJj0ppiVt4W13NweqEn8RXplHwxs
gFMRod/QQzTvqke6wS/vj+uK4YyKMn4Y6Mjw47gyJUCONDk/39Ah2h8o75jp6765Tqlp/oJvrbHx
xAL6nycUJuI6ldZxKmt11osVHwnGrPkW4hav92MqZUD6J0n9OKv76pGhFs7K1o0ZjhVwzDmHN24b
7b8Aw9MAy1q3YVpVoliHfk9v3IS81CS4/B6iZgdUc4umUBnwYYgmwL4lkcNR2uYPBYDci7dSVUQl
SxEK5FN/iMmTzeq/PnuZGeOoL7WUPQoarg1b2X7bCqfmEEIFRLmXG0wWAKlUzwFVaIDmv88A6+ye
wnn+4pjYE75dMn6GJ1OfXQR3kjI1e4uYOKlq/4ofxxU4XAbu8dRfX74t+Oyp+B83lEVqKSaZvz3P
wXEL1JS8q/WdaK4FbBAe0BXxDD53YUhWCVCviUvsiyMXWlNkcJZGHVVQ4oExunGUXHRgDfbryyYH
6YWBKvhv5LeFZFbvxYRrwyMTrrCw+dhav4haZRpbvwj+iPP1Ux7gagdUjmzhuctAIP9UeosvatqQ
cPYL1bf9nDwV5jBJst0Y2eNBY80eI3VPOARL06M5lXmYY/h7k1PY+TRKGuYngOiKz/4iafNgxIYl
vXjvmEPq9Rw4C07xPayoKIX7nlevFfsE9sfZNpFHvG0CJs1mNMIz9WWtEBriO5/F0j9VCcg2D/+M
SDaFVqsMzRKpTPOVzbgg+7vCMbkukhwhq6GHieEqdEsI+lvT3p9CuzzsXCgFIQvK0eslO1X8Jd7m
akAiJrMOrEhVldFAEbfOcB7ijSLLyBvZcgwSkGi2jDrl49+373Fl9KjSAPzrV2M7tMFOfSd3J21e
5UgIF0Dq3bpXj2xU6sbPl6ytys3fwHX6RjHNfwS+24pBv6zIV1L9+fjquWII0AKu/rnIls8LLXGc
07XYXdFde+8cw6NDfvzS2KikFzHwbccSgStdjLFZHeqbJkLgCoKTvOCGtgHkWuKOk6C+sIpHNIhM
iksHHSwlG1rpbQRPyxD+FFt5ta9uRGLMQ7eN79cwXo4WY/MgCl7uS65Hl/XvlOJmudTYXc8JwmTm
GYmb3fYkBOb2vmTmkSy75jPEgUgwtTv8vSn1Hf16DBWFs7fSnTy5XpbM+Afy7VXNa8w6v6fMRfw+
kuBViJoV1jd+Df41Jx0Uo1o7vyDUanZtZHwGM4fpZ01StamdOIMAuYn4+yjA6HzJ/pmmHokVuA6d
QTewyiCvOJzf/SO6oW6v24IUoVOSd8grlNXttHc6s0R+zTHvk/z9vy8gbh7PgftaMX7qDZjJMG8B
yaRwWylWyiijk/ZGJOR0PdvDih0NSCghGWIoV6jSLXWPrGtZpPGFoK+6QDDBVx30FawQYyH4xTqJ
t8yKmFs9MybXyI/DNBqVYfNJW0aNmDWQPxrUgIDnvDZQuAjf9IoRqglTCYf/C7P99q1Ur6fA5bGb
VLUu9UcceWKYFST2d6Q2z2dsstlUsawb+2bIpqmcjb4cDMVXRStwaUytCBjIfyVhkRXQX/aDMvDA
eSI3rCDE2MExc+uyTdkacSdaY5qE2ns3kwEOQQjzTjsPlWnH4CGBkt6W94UGz4xhAJK04Uv8BBjS
DDOXux4eLgnBBrprxhhJMpPMhjzmYz+FvBt/0ld+felTk3e10HmqkO6XvVtxqjT2uAid1NzJ8eJQ
sgttegpD63B9JevtgUiuOP/Ir+w1WxZSUGWWt1PSaTwF41c37OrNnhUZyt3ZJwDowBGOK4BIFc3A
3Oz088lhpHbH8WhmuWcADhnYC4mkwOp/JvXIxHRjlmRmVAmrxeM/cUYmzXBoOd3/t//WpDPJ0MAz
CiFC8HWjzArJlWNZyuQ/e8wOtHg6EVyDI9obxeDnXOFILE/7YhSzuG2kBat6r8Mm3myZ8wag/fqM
Ec770OH5ZAjyhqZoucCz2DjLTWbUdTicHUekB0KN5fcgzRqAX6P6hzseYsXLSCn9V/wZfh61QuHP
vsw7xCpA/x7aIvPXqmhP9bTkouIEVol23Ar6R14l94Si3UK7Y4Ol/Z1GOMT4jOraxrjJalc5zQ7o
x+ePkyixx3DAWGt8IkN0o+6V5ocmETjJ0Ds8JVt8DqFFJahXsragRLq0pkYAPNA5/ARK8yUdvhb4
HqgRjup8fxq+agu4SxNnZSGh/OAlGKVCjlHdPpzl0Z44bqTlS/geK/5gkYucwE6btK4IUU8zKOGy
sPlSJ22stpHqkBSvjVbD1NQklRlFykFknRYQzDxbAcLcxrYNx2ugTe0goCQzwj39xoMfX4UStiRO
cHFzakCR9BlzId/N38PBSvdlOAdCO8+vZqjDCMhMJg04lNCjwbIIK58hIZjTlIQwMtr7XRFbauuH
pyJnbi16mdrJOQuZ3bdeV23L2MlPFCwoPMnbp9tDgcVYWFcBC4g72ee8WS3ToMvppcoNlLl57fH9
hYo2xvikuw6w+Ot5JlYeO3ASajkIK0DY47dZNUt+oLWCKY5Q9GuydUB826QartQUiFK4cPabD75a
1I4pWqgD+dz+b2GDwfl7rgrSzG23Xgsr6AnDLbozKyKXV2MFMKR6SRoGnEwYLKj4NtlWwWvBOUA/
c7wRl8tlfBjS30PP1J19eGY25Ej9hqG8irBX/5DcdOENE5A6ZoqI7kZUR+cxMqapSrR6natBhLd1
JHxfvHumVMFWFWICvlzWSfzfAD3cDlE1Q210JJqsYcqNa167oY/SR3ZF3eKcyPnClhJDZtH4EQSN
FJveOfD+yvRYE1yt/T0yqb665eEwCanRsVCMSrb/xRSxrbiCnRANgGlsCGoz3exw9P+GwDNlr1WI
7IwSfCvQd4FYqnRDC1WdYz14hiq02If5300BLofG/yiOLw9OQ41QPjPLgZ1Wx/nzOFqf92uyzTZv
yZn+noEb6SXAQoIW7DW/gawepLyXzqo1tZV1tzYhrO971bNDhcFO3XhL6uWj9KQQ2Wx0ZDc0wC50
GmICDbCNSPrUXGC/rjsl2SZXUDVv4J9Pgz6eCTVzFu3+cYYcBOB+z6nLeRicFI15iozr/7tvjuPM
6OsaZXu54OIhmeVZNfJ1ElsvMw35Hwdfgj6g6iwLm7x+UloTuVlyf8vSJJwU1UGv+turZVsRy0A7
WOrtLoxyaFxTabrbz7T8CgI7cHk+oFKBZ3SyCigcAC0OA1xG5f+FbEHFy7qByOwO+X6PvtkF2jgi
znjUK+g/Ua97hpRsWUE8rva5oM9kpYrHJEwYOOEcoKfgd5I/DKUZLD3RK31fi42bbju0hth59QEQ
+ytrlxIeD0pH0XQlCDOn69vw5rQ1fqZIg4Y/UBsOdE4wFl8Ci3rddpSZZUaK8Dv/zsuNNRbBc6w8
d/Ef9bCBNxz2qwQr8xsTohr68aanXl7zW2NVs04LbjFAqXUE4o7CkmWpo2zpmVqUK4UEpCK64AnX
Q+IceXYkEWs4S9FShdP9HP0R499UEWaQwBicpj4jkQxhvM8pTiMH7jhLf2Cdi8bTH8XaYZ6eJvHV
DXS+tZNPamIbAV2KexKra15D+ywQsUbc6a/93Z4EtyDhtENyRtkqBHjCfkQ3bGszmxdUX6t7/Bf2
79a4cYyna9qqgTklguN9c330vAgz/GgRLKxJYEhmbu6El/CdYzDDV6+aVRPHSwWSxz64A+KWaEm0
Ra0whJShWnqqJyvuLf2WOXHeZdIaMws5dAjOgjezRLaoUYq4Ko/biYnAKuOj6/rYDGIxTE+0Kqlp
gX5dDW8SYKlSfJVRmajvwEyT88YnpVowBdg7eMjZnvi8cF5Yakv5tGUYQx3GvOsqaxH7QPfSTTfA
EO8jpY1KnQTDbHs0Pd1c9xy6elAzAE/Pll3DubXpjT/lgCCHPDtPgA5x319ITqpYivA24bHc4y8r
bu6OOpVp0ugyDBGOoizgnSHA+Sy7OGXVUlxQKIrl02DiHoX3kg3b1XAmo4Tvey/t169CxK2bIyaB
cimIwHKu3oKOngNFBTX0aZqnM5OwqEz916D1Ynr9ozvWawEbZBJ1/IF8q5kk7Z9SLT1smN4NkNzP
CsE/3rpe0P5QmOX6mkTs29LfbJuF3ye5/1Iqo4AApoG22OYMe22lA+juYjhAIDpVPjrTfBX/h/9v
JSSrHg/eJWty6yTOffsmL5jRSZnr7qCc/yf51g/PL4qi1JKDJlCPuNATcSfsSx/m/xEfwBvuyyqt
mLiIirZi1k6ceG35UbjbN0ewixe/At91sjECUAoZ8h+rYtdNG53ovin9dtPjqAVAfNrMV7fOtg9Z
RrpxcEsOXmRa5xHDoadNalg0TE4jYKH9v7r/e8AM+Ga+zxWLGgjIlAwZ+fnrtNR5CQuRK9hUe3xp
mLcqP2Cmad0o/T7iJidHJ45dnUCPbQyXsE3fg5xlI7V3z9QOMVGh2xY1KIeKHFA6ntRGPVlupwFs
nUzV4O/ewo68SxdKvUJKDST+N0ugGcAbIRSrhhaX0B5FuDGR9CIwzm3tprdQYUuaKy29JBEsaxtC
1m8gdklcqF/lLp7xArvy1u2p/6Ag+gR9vvTjzWIZR0ccXagB6iWJEvtcZHiZq0YSaDk7wKWme3tB
BWQDpnjf+VlWr6RRcZmYpSPLKB8PIyQdJ7/FYOoPWZfkVARJdhpB3QcKQlGpJ9ANVAiFdyvqexaK
KmlWRMAD2gtGJiNA+zxYtxFuTo7fAW5KToynJIC+7jyvkN9xVt27799rTiXhRSQjNeEqxZYRLS7o
3zoLdUa4wN3bUT7qumY7lB8wpPhMTTzNIBbtk8il1NRUprCK7WCPDRymRW936RlB1oD3nnJo9VpT
ltmy+O/pkCCa4HkE5KK3RrwSykAht6QRuUR6bP11bQyNw6IxfX1I6nMTXhNZBC5g79NKp/mtIz3/
d5+DB66rIvXuB39MmToacW8je4S7TAOaTlSRuhXEn0YbryHUKU/Idb3Ov1IELwvxsg3NMjPayR3W
fQqLz9hu5N3PBqJlhdNaQr+A3B/sfoilj5Pn7zBGniqOtceITrzXDl93GZ2vKRJn9m8u+ZLJUAXx
E162XHSdb47thzD4i0F6wo5drh42tKO7aXipTUTTQs06IW4wxJJsA8mNzVOZPvFwltJwuxog3krD
N0zXCigYRquW3K7WXVDbxo8NAX3E/AqfN9/esX0aCv5VDMN3zCwmj1g7nInp3emPKFmzEjkSqFjJ
35o9506ZUx4bFTxZ/iA45v/WPznCGobfuUuFJYbXrZZO74+BX0+DswS17uni4kQeQkbEhqJCBftH
evIBFFal8u8ur6hOmU5np/2LOWqYrNwDTiEUHcl/v8et0F+5Fu7aWDQ4Ap+QiwlSjbuqM25XgJip
a2TPehB05Py6sLe1AE1+JodbrCveHK0BMGOxI3W+hMd+oBmBd8fjtdgO98SMqWB4mmjOXqw7WY5T
685wUHTOFPiOXju/pzcdtLczLeVTzFIhs3bW/NI8gTFhxzgWn+qT4ZxOs9+YpHLLWJ9hRgrRJars
GEaAmp7RNHudejMBBU4ACx6OjgZLK4bxHeb6aJlynsg8pkwq1i7QlljUCQq5hExTRmNl22/usiZS
likDAz6nF3JVeBluagd5F7kbfKeZ+xzNn/UIDWD0dKkVSH4Wh6lhhs3PUtlWfp6uewvzZhjdKWvh
ogXF/mORS2qy5zqsWDqp2+GvoPoZlvWdWFhkM9djm7WfgRb8h+2NTYcr3MVpLO4rVxRmWWw8OiNW
8kMmt4U+OKsd83p45GKmVqHDiDooOoVoPYC2CB1OAyw4WMSii5nRzXV4TgohLi3jd3U4YDBRdNn3
smWJJ8eLNGL/9OOjZPgzRV+BB9kiuokeE7xihiPftw85qbuk33mxuLFYO7Q7FLReHXs9qB62FJa1
l0xXVyG7i2X7M2UozoyBG7YuFGHPVjrXaQ/BTwYttsIy4Oj3h2eTTFdW7SziZOqsWsTvwHv6ywFx
x8jQfRv9H5VdZ6GUXEi42poh3gGQcIPON+qPrmLchNal8aVFFwFAHEAlklC5jO10I3RSD4eawMES
LdFWbJEIhtpa9OfdwFdNs3gECPNaeTeHSeNAAWZdnPJ2BlGcp8UVj5C1XbT82x9B0Ce2PMJG95iQ
dnBDm4Sph5jnJin+8S5GEVe7cU0nVCBR+teaaI/kKgMFHVwfMv2GCBp5kNIT3MiGdPrABzaT+2m3
Vej7fXGQux38AoWmVRWLvwrvvWcXuP2bQ2UTA92YpSs3QOtPU6i7UFwiv8Uo73k4tyL1RXDm/3SW
2a1RomEl9YAuhI/mfFE27zri38mK8xEeJCKL18JY+BfybNdRXAIWGHTNi93U+vYjRbtkburkkEXr
YoMolfjtsalVaqKF6gBWM3vjYcXSUyVlL72BMGThRYMTMF2k/EWWU4JbBMOZVm9ZabHFSowg/KV0
KszQsQrMRW+DHNZFC+XQQOq3gQEHK4WUa5Oqk/Nx9rOfU5Bg/nFlsYeR48zc6C6NFfltfNSl8OLe
67IkvhBYQbejOaeckvrMq5fD7C3XAfntk0jiZ5wOOzdXrstsqquWCuk5nNn31VIaKFxb71IAeMle
H3jW3na9DMY/v46QvwhxcIUNTlyzpB6QHp0iWivG/OF3m/uXp7VVsx2c7ekyEPm1rROYSty8s6kM
/dzR758SCmFRV8gun+Mtz/AI2t42jLsAe9zDRa5Lnl27OX1LnHOG3GojLQ5GuArvLOX/02qLVO8M
zzlpWXYNuOGiwjFVuMWnHWNPV5HrR3KdTlImDC56byDzqCmH1538soC0QShDLgjwKMhsTYMFsrtm
2DbilJuKBYssaOScq2rLN35RtiEQ7Q20vOXmv6dHkMZjDPXq5GcQQ45P9JfeocnbsJMgsNkPuPnJ
WE2LCUrJhxgdFTx9qJLwcvpYpRwEP61j/7lVQynhL1fNqKPH6FOZ5+Mfidmh/pmqNWDo/SuG2bU1
Sw8NNZIv/G6by4ooRkSRIiw9RLX4gcWxw4LMv9AQzR428BKHjT8Cj00GFUyU+rtMTFA9LTloXORM
w3ZD+id6LqN40tyk6ETtDRUo8esevKkW/khOwxSxy0VM7qHD4GH6hMs1swZEV6plZfky2QlWTtbs
LOBgmQhbeES6K2SfXUgUssXdAN2iuSCtKoYUzWLaYrzPAEY41lI3amGwTqsS4brGAuFfH/W/D+bv
LfXj4wi5SQVO5lawlNXRRFOcIL4wVcz1vN1aSNrOBG7amN/8NBMD0xh9cT+E7Gvnk38PVttoMtjj
omcOm8HLGeEFsUgdwIcLyOov4NxTxJ4jHBv0bZ32KfA+6cTiL2ubxM4X4CuBr2A3aSCxZNiGi9Fb
OHQz3+3iqyJg1c+yYJGjZx15RhxHT2mLOv50wgtciJRAa1NnsvFgVgI618AYPCDMP4M9c8THPC2x
o9c2Tsrd1tAFwGbh6zFxMcp2SkAdGeYlba+j/Fv//uynMnEHJ4qh+l2SCTqaQCICso+yTrKx54Sl
SQFWRAF7WCOz5hBcVbHLHfz1YuTi03f96YroUp8wENVcSJRnuTQubkHRPtvKWfEXNVO755OTcHVg
upMO4WJlL3nZ54MfeKbpzw/YziNPtGopcGpjrHYkO6FjlHImH32WvcpmrKQr4wkRHK7gTfLLFHvY
YyNjnBKq+hLdXIGrh+sSXxuLzAIDRe8+1CIIFGZpR1iiN6Byd9zPNcln4qkh6EC1MEerBAN4HO9l
t0nCA2hFFtUj2UIE9DMGy7U5vQgtNK+8nyh84sGfE3BDQu+gtMU2a5U2fumI5E1RCCVWx82poNzh
sc9J1kw+aHZzeJc/aZebp9xgA492CGhzWMzon7dHS7Jh/2MckfMrFcUB4HKHFwE2SKVfPzK1jP/B
CSj4xbmPpn9kO+3lWKFDVAQuU5sQ5KKTeTiHfbFMSiIF06KpQRiqJfu4HufiBK72ZzFOS/7Sm1hL
l08tBarSHo6jCnbgbM2b2EMx/2R9b+6hUzjt9PcJ0BMIYwcHcoY1+sulQ6u5x9O48lkFdWnvX2gE
7ZByIXMJeiejT2f3RuDJi21bPdHoZ1uHxuY9RegHfEoIEGNYNGlv+0lvR9Kf2EFXtwLAr7vGC/5w
cwYUegRZKZXG0N2L6159nWLrbXiOSU/Z1A1i3VKAkQT88K/xKf9F/I655I78nT6feGErU7nbwiu5
ZSnINmM3xk2Rj9VqneHW1mkXwA6enSv2AcS70kFlDS62t3w4sF/T/7Z+VnA5HQ8cMRevUQuoM3BM
GEiF/9GIntN9BWLd7pTc+5663xafiWuHzHRFwmvv9G8AGmoulTS2qMkmxFdrG0pFDFaMBA9AH96Q
mV+2XrSIeD2GVr+cVH6zi9oAX4AjbUlATeqf2azLgnklOAt/9HjwZJNU5QpN2fFqqR8d29wXPdIg
kcbPvqokklnaUzu9LKR5nWZ5MiFufpnqK+jOU8jSSZPgNapSI4molYp0GxBTqqoUp0gCUPEytjlo
AtahaTvEXD3CZ+EI0rIZ7OQZ0evZYS2ZSyycclqzgWp9Ix571Qoh34yAPB8HMs+YeTEW9yLchdLu
Vad/rTOTKLPDQRbraDBdlYQu0z6I+/rQal/Z86e7ZDBOFrRl1EQR+klstXBJDajrdo/TWjEVep5V
xKGI2uVVEIvjtYqQjmz8xQRlfm0CNu9+FaQyPQOx/ROB8U+OjcqNadlkaGUJZTiLUvz8oCkVrxn0
dI6/Lvkt8zBXv+uhgvQVSZQioy4wCbXj+cYrWENLKC+lQKgyzezKlZCl/2uIuxyO2qR9N2dge1RH
kAKF5rLlnlxdBFCFpOF6CYFUSqQ+aFZOjtaCHiRSUcmKvcJh2Nwq9fkJNU1or1usLvc0RNjo4ozu
M47n6R1QONqNreEkrW526Qw3OW+WWpJgf2XoeBsa9tBqKRTfDb4y5cd0piv3LEXaqjvhxXG0FDUd
Hi7R53IB8P9vTzWRJY+PrZV7t8fN7R0iDCPH20Bh/EwLpdlKIXxvm3ylhEJPIdvr2F8UY3U8im56
XUxtkG0+zdd95Vdotag4HEWAOOhbIjuzXaiHQJ3gbCOohoXaFm5QK8ooioPH9LUESu1orIchHmAv
pGZrPBJmGzKg+2Ww7A9A9Gf4CbsgM9qVfslMpxJ/+v39agu8aHms/kQb3tbaBnKsydmE9M+lG2Fk
rykCgsjUviHNUCC+UO+xLmAlIoPpR8GLS2yrDxRIgC0ajdQqOJSW6/wpjYKDppMttoRHnTR4qaM+
iEQkj/i0buUIzu/DAGdSb7eW6su6OP3mLQ28jpzRR8fHE+hytFz2eO2G1m9xQ/RtxK4lP3Hd06mU
+evJcu0VA4SJ+ypc/QVTLfP5v2p1OKtRmPo1iFFqXzdwVMiZL09IsoYpWZNU8s0sdjeMZ43Ro7Ab
/+7hOpOzvniLzaWZn9vq7gOtLknTOCuQGylMVLaDwgT/Q11YNxrgmpUEhfyTR/XvCwb9PZ1arCnS
knA2ePmmxBRXeMPQZVAoMqX3bUxoohJ6Zs0HE088RLEW2RbkLeRBYSgwHZYt+/bYTJpgPMcesQmO
rqvzcZYLsYDUW6AmtEQ6XzeESV3fTE3c8kS15Uriid6doq1w8GZ1x+Em54DHdjTDyN/Yxw2C73TM
C2eaQMqhRIJE1Z3vNpMD86UGy3s2IkGS9qe45gxfzt0zgMvHo55WUWP8eBFGVBonGmeXdNnlS/kJ
roy8bdUM/YEcvNNRGpyuWqLc/jCvFLTmwLf3zR0qWmsDPbBvsLE5BsYfKNcDR4buhNZBgP7jn9/5
J8m/MI9u5OPZivUUeC436NoOsr5bdFWdyeBk0V3O+x6iyNGm8GHrStZvbh7O4eDbbBSFfz3JU9Cx
BRc1wXxXf016Zn+wYwFvWxv0CiFLuT/YXA6NHXgBQal0YNhJIswNbZ/HXHLoVzXw1p7YyQ6/iL/i
CtWwiTfOKWDQELmxyxFIWFhJkYd5t6giGsFggKsX7z1LiAl6mvcMWUW/Bhu3FcDLSOOyiOMH/GtM
dBHnTVEW1lggN9pwPLsBem5P7n2pWTOKOCm3fJlTXNEeBlzpWBHax+2f8I/ociLAgzDY1OOHW16A
/UAz1UGF1lxr0hxPTZfssra1l10sr8+R9IqqBkYPaZwKwjfYNlRTcHzwbytFyOqPzXEtO5KISzTk
cYIeavfxLBBeuRKFJigvlHubSuPdoaK39CW6UH5BACADRyDqBjLwYooY2l/HR7mOyw40stTuaBbr
gpreNEBa1ZK90Fh5R83NLplBRnlcs7peXM/T/FPnjZpl78KTNJQH7RX6zXgyfsR3qaS6lsQzhv+m
BaUFPyjrXRi+1D2ZI9U+ansFTjyyKFZzJBgKEhiXbPU25zUnniHg4ZJuhezL9jzvfEOYtMSowwSC
pr2uAIU5TCsAufzh+goGsh5FBnF7Gj+kqZRsFZckJzvMz2KJMv3qBo1cb5W8Nw7h4JtoIaRIbtIS
UEM7eLcizXirwPak0gENTlsFgC4KzQvLjJJ1+4S0Cl58BfJmcxWA6Kvwe+Ba5B1cL5CoHWxf9JfZ
0v9XDWA/HvlJNq+DSBve4SQJyppQbz5+dRZHY10K87nHXRhy9G/tjqfB23qAbb0ecSGzp4cV/TLj
XgKiSIy41mwEFEBuHcleOqokWJ3/e/B4jjcYmR12KKA7wB9b78aN/fd7aDy3QMa1B6jo5ade2bM4
Owrjd8Ma1LWebHD/8RrPY65rsZIfH2fxaBkexX4YumjkR73Jua6tYH/psX6pdRpJFxjtEffuvoQS
3p0AapRxJXXEb5W1d6k4jCakRDFB2yAsndbMGwLWaUHMNvHPevxGm8jrygtUQJAmx0R07j0IxMnY
Px4qghJ29br8DobWUUMfXZbFNPtT4wJiIqyTb9iNjb46Vf/yitN5vCmxM4GTO33fh7P9e+D/lRbF
lD1WeWLPRD+eqfKT38Wh8u/OOAgu9PFcBUyj6ql3vU4tdg6MlDmx2qTXb/1fT1CjRXM+ILC1IccI
4L3mrAdMEhsr/b0QsXxZS6tznwF9W/4HJYKle4wAJjDumz7szsL4nnUtZBTGusdt3Z+1w9azxjyZ
/GhoUpqutGRkTNscq6vWKPupqO3p6E7k6TUBExkAbNc98nBAiJ94levdpW4UWmnK8yRFXMbB6SWv
P7L8QnIFgbS+iCQR7HjYajF3PkhXLnTSpyRpFQI/LlT1U4LddLo2RJUvW65cmNEqmhS2YDfy0AIM
v8QyHvxvi5S8O+Nz4+xJNyjLZGJMdrTacLLzFejMCZlD64sziKsMjdoUeuIZrLATcdYbUORAmb2I
pONLXEXrq3ot6Qgz1M4o73dmZFL5AtkeGzMd/bfZT608iIXNMaLk9XgmxEC49QPdd9CLDxZRqDGO
xEVfFMWZHM3KdfXuLdRz2wX2a6BqTqn7un7KqGaG7OqVrfkRzjbQ1Gyz6CvHh+V/UbfVvJtKOaGd
ScCTlbJwQZa09WjSR4ChoBTF450U6VqXYlXxEKfITglyBUb92zlBP1w3mb9Hooq0WTWv/C0jfPra
dTkXDwKFvAXF83u+aUqj+PAQPP4L/OG223OpFF8Hu/xOjrRTLmVA0VY/2YVa8t4KHeiiIOf9htnS
lA03pBwRxpBSgBu4jMF6pFzRAZ/IL7VdYayVnnXRUHg40WWDeA5cT3CH1SP+bL1Go2IklNCNuVHD
9v6wIk/8KF6nY9FRiYzkk+nHDyiXbI/Ygd1lYkyOjJaU3UmTAjM8L+qXX/kt8XYkmgWDQU5uPDBX
/NdHcQwY93yPZssDgcJBnX8YcJqKFPPhKFmu3M7R/mFRBjLNLg770B0yBLz0BVNVZtexeXYADoXj
z0TSpQm27lx30HY+9D16nvJ91Gb04qjg65OT8AxSjfRVaQD0hVnzN1jWUTrdSejudgvLpbA7V3zu
jqJrCc5mtIeQm2wFp6kQvmQbzgb2kDU6eSbApg8KiL+BYEEyxRqrc3EWS5hF87TG/PPZWhgJD2F1
nu9PhHljO99YDX2b4MPq2L+iEXYNJJ7bgZTm9JjIVXWo6d4HMSd0KigB7vWt0S/jA3h7c+4eOTsb
lHLPO3GwsvSqKj4kSMGokob6t5MUrLspyoyDV7glMcCWHMPV+NfIQFXECG7NtdKB8JIL2gdP7o4o
51wx7ZXydN0HGRgPgwIzjOnk+CGO8+EdXfgZ44AsmbCdc4BOQhz0ZN+Jp4t2tWpexLBuJs069CGa
VOWEotoOy88WnYWbfILgHYMBbpzb26Z8qMQQioBSWqzaB/sgD6+sHYWjkS8AE465uH8rjLQjno2j
ChtrOnXbCRvyz/BkZ34Oqsf1+x8cRD+V+HRw7GPG9Ah00cErUNCDgcZRJgeFTlkr5BxvRCMfxtbe
rO5IrxICs52jluv2y4AlslKmOoBJ+c4iwAOOUXrjlUQ6h9VyeNJeo9pJyMrNuguhf5n4+C/5EqFX
6SFcFwVfAkSGCfRuwz2qk9Zm9yzKceQARGkobxgOoW/zLhn3bMSmPnnlA0oAhJ207rXIXNY8uom1
BBDfjWA3NiDRuPGqrBIT6ric7Pq3b3j5DEo1Hbmm7Wx2D16kfOQ3GpRx8H/9eQhMLzgrUzVyZ3hC
vxE2RkNInNGqBV2FUtmo2MxyQ8w0EHL0pcwCpe4xzoKrU5ZJgCffOsdnRMcgcllDrXo7yLhTs+DU
wjUisI3k2rokoTl38Ur/bFNebJhbT69vXU769e7WsvbWV0C9R+Xy24QxcC2q2+jiUPIpGGBb4KyX
m430KeYMHGGw3UliQdaALfHTMAVGOOKuOiClbIn4YejWSBQYWOF/Dshg2aHyFMrpKyAXUWU0uJdN
7Ow6cze2s80gQmz0LcwkhFytLGRCXM81xPaXoqgCTQuTQ59fKsJGmV48bbC3hPPaiXTmTfC+uoSa
9eBgmUqcyrlRvaPf3da9JbwuBmFqs3URyxW43lLUkDavcV8/YmDV+3/SppA987rsS2e3es1tzgcj
+LKyvBjWhFoJhPEkuaJkpwKUrQ+QA2CpUxAn/iKCX7M4FYWEsNxbpJn+ymLFUS/M2BVO6aPOH15u
ff11ewEpLs6ElKYEipPOkGVpXsDVVgy36DgnevQ7z4JiuHmKIAHdL1potsZEV3Fxkr45sZrj+g39
SjD5hOuEd9XOKIuZwfsp/JTggVII9HfY3k8xNlpb/bDyPrL20UEkTVGWsgO/iu8yqlaFlMz0zjIa
3PMl/8UenmGhaDJnBmgJbmmzRj+IWfyfKGGGltsivjQSLX+EpJP0SpW+KC5/vILxbF8JCg2DNGio
uOHeSyRc7h7uxGIYF/+aAHlBiDfk4y9vuyJNaEo/0Q/KMGMh6xR7RDAOD1ef9nSvii0nE4oIsYxj
4ZNAOf8vSHQgVq1NSkaITUkZ5sWs6iHiaytETOkiwocXuiRdoiWVPRn2DQwufzm7CS5T9JFRMBbC
xpERBV+HzUQVJu6bIC91UPhQiCKPO4NxVsKEqyZJaYvxRgjpmD0hfBkzyBhTGmptjuH8Ri8T/nSK
MzIRN/gwgM1qSVMLHIlpglzGYFbczve5ap1kjwHs9i3hI+/MmCgx9IvyhZAPXVLax8qQE/bMnrD0
hj5mbJku0beDqC59Smik+l/JistFAA2C1240PVDkQKAv5t4aqIaoa+oSH+SrOqNZozvD1Ckx/JaP
+AJTgFir2Znp+wLs61l6aGbpgaJ++fhnfeAlpqT3TppfTj/CPdRSlKJ11Rq7CxX+6WKdqGJEfsC7
xgGQvdNzgRj2tNYDmw/f+gjSv5+qaAUsXdhGnAbixIWGIUhZW+WLfMBzVygQtoqz3x6FHwb164V7
EXvMuaczBKiuZmWyLJRt2bvD1h8co+MvAKTaoP4OgS95YEkA0HWo0OCo+3qoTgwOqcRshxxq1epr
0WUBC5o5kg3snVvZLOZN9OIKSaSTPVA+VmJZcQXngDWL8vAAYT85iJPhNnBhUx4PqW90/W98DXiG
yjoLqy1slDmNGXTUB1D5D4BS36z5lOv3HpjhtfOO1S+ZC5cxVVQgtRcmP51GsqqtnoHrXBSJYN0G
4W+/LJv5SejWS0H549xUgy0PvoyQ9mS6/ZceqNDTjaMvLb+Ph5XDZLwowhF/mgXU1Dpc+RnldhDp
t7javwlYxSa1JL3smWU4IBBVDs+XsRHcrnbOTICxYKDa7v99a7LmYK/wWe7WKx/p3hTo4vJTB08R
cGO2j6dpDTAEHHLDgyaJyODr4a0xqW0bh5jBFnqpTIljR0FChCf5iIiYKpCC7YwYMaI+LWadIdeW
ALH+RKAP/lYUZ1xunQEX5ADkuQkul7zRwQnspeLQmhbAbQoqebfsleDam0TbpVOWTh8UJCXczLET
SvRVFkPt6NGsKh2ZtyJOXRYu/9JbclZ/y6cDZaKCawxar2+PHNToQI6Rzd2CntpTjplmZKyu0fTq
Uvudw28pETkPS5CiLESj+4u84hvCgK+YLIsvYmawUK1YXvHDY11RA818gOJJ0N56WisXyP8e+3cn
5oGtGPL/ge3+AjtTJYPeR2p4G4m0049Ja5TfEUIzkkjF2DQbL+I9JI8y2v/vkD7/ZqJ1pAWqzaZB
P0PXy154MiAo4/5T18D32KfYAOqGl9eKXDjDJ8DfOhp03EntACMdQVKJ9ZXbbKLztQkKJn0ltXtM
Sse9nFmZpT93GGdQsWA+guH8sN3uYhRVUaUuCyiDngIPPuDUSBkBf3LtdLMnB/jlLAnFRPHst+J1
GQO5R1eAaWt4ARpp07G4qbUfBCZZvwZMwM74sXJz1YLKueZXJ55mn/6SauUaSiSnadX4ay14eiE7
jKX9LOFcyPv8vUObyhqZEZC7erZPDkYtWlwazrCt9TqQbFRMNPvDab3XxhdgEEPPeNQSSKV5rTAP
7/wT/nia/W6kckpnQb+tH/MWFiYwdGQncQtqx/NWd3PIkR5fJ1nq2Nlqm+m2F7WIW9Nf2bMqnfmO
fKNvUiwFcx/XHlhDEK+mYjXb1mxx43kbxx423HeZfZD6vdX3j9nYUhcLZaLPpci35xf3l1UBq2LI
bLZ2IinSFO6uYWoycZqKWT1btDJ9Ldx2BjdI5WEZnoVOQIL3jIqhG9Cv3MjWjWldrRKmD/wQpbNG
zoJWGUr5y533//ph+OMWhM75VEF0Ag4lqbcJSY23xpfblQz1y5Wt9urDhR4LcDu4IqtGbNgnwhEL
wV6NxBx7KFoTEJMal0d7HDZJqXjU+7v5MrszO6cvgorW/aU2ATPptUg/PIyDLv/sNiLkxHSGv1Qc
MeyZwkNgPhPCb1xnhxxsRWa5GvV+q9yHmI7vJ62B1gBcguB15LQcQMmNAWR4BMow3Gih+DzpYnem
B/DvykN0cp8uSbb8iZeEWsNS1O3R2zRhKO+LIDRS59p15EZi1WjSvb+n1nM0PLjQvk3oBTt7MsSZ
lHVZHptCYqz7159bGezasoaxvx3bWEKeu4cVxFF6n07Bi1C3rJv9fEJKKIzotUlNCG7lhlDXRlPA
4qFvfco0kOGuEpaKhI7Q98JYG/LS45nnztpsOUpY5XrOGKbpk4eeH6XIjiHSnwBeXMZb3qiGY7Mz
/OJmzTMDdBatL+7IjJQ/5pVgwdsJGHsQ+l5KWRw2G/cg5iwpHhhhtTYdKUhm7yd8uH5DqPFnhpLF
dCSc1DX4BQMbKBKl8FqfJj7BBU0CrZMExzXsERy3VxSPQieJRnxJLdoGempSwvuw8snqlgMJny7r
8vF9FAqtrql/iBhRbNDZwVckQoThR5+7ECaCR2qX4Qmb3D6jXcnoXuz3oh/++zmnbAxir6MzE4lJ
NwGUngmWYpNSiEzJPN+NBpWueVMv11/1EPMAkz3wv80vURqD6Cvwc80jcdHsMKCRZkXfpOzL9FrQ
NEZlAcjyw9xVcAYlzFrhxLsY0Xfvn3vYgDv1cgvHCuPf+MdgLtFIy5Ei4ezZQ1pW8x4MSbHCfu83
rNrzDcL+47GQQd/IqO0JH1N0SwV/U6/8/tiUmojB8gi6ATmAX1d03aVK5l3AGYNbpWDbMh7Y4Yhb
C8ya/seXiOLQH1H8OkFnpY8wkneMifs6vdHsbPy1BuZsUa8xPsZJIBBu3HIoPgOGt59mTNrgJlZA
VqRjvbbIMEaJjXLZjQFgK+xUz665iG+l6J/ZNqAxh51WmEiKcTEv8abURAPaBmZVc+/uypv7aPHx
zBM7WlydJBtodqTpn9Z8CqVZWcv3qW7f/GVN1ImuVWJkGuCdoIw+wzTB9xiN695Zx5I60EFB00iC
TlKvTw/Fp3jMnKb7q62fBfMJ+wVo2AvGcT7pSNugHgEDzdpX5mKioqwkETjP6wLj0OPvHXLilJfx
sO74Bu4EMKHA1LLDLFuaqzlmrnFBruUtitKcrFrNj11iBow4mIpzPPSkjKZJHYJC9yygMoRkNnKP
xyyftNAcfzjbvxW/wLxZBTLm31vUAi1HNHELUJs/7jzCXXR18NTjVL9j6XnE66E9ZjQjYRX1A7NJ
RQcCp7zY795D25t9wmVx1u52XCF4jM2pzda+LQbCdxFh4lGBtzLWwyIKOEZmYZ458lrmBcmHG2Sz
16ZhbJ4mkryiQ9xXVSHTrWVI1xmRYd9CkK6iw5xV7Q1Ph+gDHy9qA7WnhH1k0/xEyj+94qRKTdnt
Pqx9B1LNx9PHqaQq1HcC/8ic9DH0vwRmQieo7JC8gfUnKOVmFo3LtnAjOxnhKjK5C0eqHDETR3I3
PkeVe9tbvJDogMqSrICPrt1QiaPLSH4LuWQ1llKP6wqxEk6X4s8uVWPxfxoB6VzprhhlK6ULsMfc
yxslTBX4vJ1T5yvC/523ae1puJonNLnlsgwl78ZF7onsoWljNCauSUklFzB9BNncWrdmV1ClnfmB
maZtQvG1ItJ7LyXk9BimWS3MhuOvcJYGz/nL7isLcUXP/B9UgalToL6QwvSocbEB0MtaDkgnXgEG
T5wlUDIFLJfOeUKDpNTFaBRB0E2DA7NWayYA4DlpZId1RwQQGQ/6ECR07bsSerZGaObV9J3vxKoL
1A9klO75vLVhYZ4U+IwUP4JgfrWFGHWzDIDB8Ifhm/tkiXP2g9wGdQLxVm470pBVH1d/5WvIgsRE
cSHIFdyUug6SJ7kNcgmUsrD5PS3fkinJtHq5Y9cj+Pvxzo9jUP0Aq2pM/Axaju+ARjGpl25TPlbg
5BF3J72VnFOCO6DLnMCP3mBOynVDroL2oqBWI+zKjwu/usGWyN1VwmG9zqlcJUz42o/7agcVUL7R
SScderrQ2I+PRQC71VgupDYr717KRuf1aotRBp0kN9Wg4rD9jzG3gLaKiZhWGRQkRpoJce6GVOhQ
bEGwfTU4o1x8Ckv4NSV1mNP3sFWAyvo4jlaq43stxjLf46IULvIqKhUiasbM8vFlXrn2doU932sj
hfOAeU++rdZjK5yOFDuTQ4yIvrHzal4XFvD9WHiX4chXxmAsj5eVjG/nEWgp1JQwH24zq7rLHqnX
BuYD7a8wB8qztwpmnBQGe/bSRAQlaAIayWjGXx24H+5TN+3hyh6bjIxT5tFULT7jQwOwYkFzJGh2
r7QhWwid+aZY7duVxb6gjW1a2gQZ5oDlliJ1XpdYeOppsLaHGqUnUgYXjwXf9I8BjDD/gkAYk7FY
Gl/v52fOkgie7Y3nDNoz7cD3Ln0YDjYNd3lqIxWhnvLOlVIO5lDlycsnkhyqoSbOkVsAGUYaFUxg
jy7Ny4bHTqlbsAiE1uLPT4oJGHBxmEAx+usBwfVE1GqQelJqa2ayojZvqynhI2uX2FzvEZ67JF6Z
pLP/8+1u4AhGqZpKEuKjICpYtbPeHzG+UntfVp7fYtYsy0aP4wD1g01ESo0/JCcjp1Ip2Hv3Cc6g
9jR9s07gLGTOX/fHFzStyDPufro6crMawVw9nJFBmA/9AOrnsCdVZB/a3xTp4JVeFY9zJ7Hg2Mxl
9mGTl+V4hA66/PXvuJt21A4kLbGMC4XWoev7u0DFN1P0+lqatjs6IovtwS4MqWgWH0AbGPP8LR3X
C7dXKc/V5zZbS9eWqQBu/zfPE67Udy+yUpI/kEE+SgJp3ISts6FzObVvt/sFoxF2A8Vp7qNpO8oP
eS1kaEYCMVBKBPQQvVNmNW71EQA7EUi0/upphzHawLyx0ylgsfP1AYuE+ZcDDa0PeKgvnKdyUvNo
9KV/7o6q7jAOYJsme0XpngBsV4I/Y/KrpVDwLeWV2zHw57O0OWKaC5iaAR9IxmMRDMOWbwixgIvp
Jp2pu7+s6GfZUVxsV+3qnRZnL8Vh8KdObWBvWidwSgwhHCqMot1VY2o1J8NKyf5++A9REuT0I1+h
ILBFG1/Fv9/VKcBcwLT+hT7EA99YdFBmPL5YDI+xRV/bzWW/vzCJCxuqwTrIMrnh5C5Qh5P9oGTp
HavuupgTaVpNWD6loBHOGckJkq/ddbpa+7TPeDgHlMQ46vs9NLGa1OxaF5f4krq1fpiuiXmUCIvj
j26f0saqx3ATrcn4UdAZepeB4gXBnOOQram9MhmcgpEuXjj0fTAMsRxmAkw9sumT0y4d0Hzk7nPe
eARwK1Iftbo1PHscGZIDJpKPEkmmhiB2T0QOuBaxqumshVaxMRfCZ1O4HXUO8IpbL17rm9Thrg8N
Xtd1bJh5aHUPzyfAMuomZJRwsU5GOmlQmmXQzLdiu0pS8p2eCiBPQifmHdmW2ur55pV/TIGJ/X7s
6p1KQ7qbn2lIkGTi77P/1hV661xxVV6Jm3FxEOrMrDgFyozRKSg/dz52800XA3CwZFSKcZEB4bv/
6mpGonbjyy+FHv8iiI3oRopYUxuYPDU+R2p+rj86ztXp1LhFbl7tS68A/8uogZ20E0kXnHFT4pcb
0a8r6dhOoPabC0CHGsRjdYhJWbbKR+uW3x0esD4PXflgI2L76z3+vC/Jk9SSmxwc6H9S2ZBnV0iC
v+U4W/uKDq1A6HIH+A/cv9P8DB0hJtlS8gjuMIDXHSul5tZYi5OKJGVtdJo6ghp4jhsc0782PzVF
SoFPnAWE1WbNTrmBT85UPjY4x8M9m78czvttKEoUr7o5QCl46ElKlbbmru4qF7h3OMe7HG6NUj0v
D5qAvVL9kT0Sm5lCNxJMR2NYNIPkntEnvzIkmj0lIqM2x5qzwgcS9dCTME6BYj/UYpxzrioib94J
YkDhetnPSd/rTIC6rpP1iIWTf1DxFawZKiV6YkglFl9EJBA6ny+OU2QytUTeQU5sEdjb9MUhGyRi
PXP1bvjxFFb/OEdOS6qUe9SpfiEj2REmMtbESNwFhqxZmfWXB5z1ImSWl88bdkymErEwrm+aRXJ1
fyyh36yMibUHScUd87SE0JnAFGhzmd7viaw3TTMbu1k8bOpwTC46bmH5n0TR9w3Tw4Q/k3lLJ4PY
kWqZa/gFC1C0sK08uGvjVdO6Ne4IZd49XzWobC+uqzTXTZvYV74rY7PMuVDOp3pykqDB9wMe5Ivx
1g3aX6+QpWXLAPX6wngLP9cqGd3OufCT4AS7KJv03Qt624HX/X3iZuMXBy+dEl6pN+JuuwKFTafm
Lr/mjB5TxfdFjhE+SNLwXY4qTdKB+zz8ri1wvTuxm8RMT7PNy8apfpMpEIsGK1LZRxYqzk4VyvLR
VWxrR2KG8FWYhPKCawi2BVR9xkihyU7ZbqLlJdYUcRLNpVws/9c3B0YsvItQzby/WqbJtG5GwPU4
pa14/8kP941trTFCF9pfVas9hlctoL4Cw61cKjlw/JgBBu2aJ3ejyHG7YpKZ9VTavaRlYTOQXx5D
gkIqBTQA4tnL+RPJPfh/onTTqYSOHUE6p6bxooXkFORXX1T9dXgVV1HlWDI8k9A5EX0FM1t7TKNf
GS9CWDacR3BXODSusxd1gokzaaxMVpjb7cjTG+oMd1F2yk7FVxLzxjRYwkATwvZTshVChXzIpv6M
IMXCg0t7cTXAutrdKGVHUmmoS7a3wYGKsgnujiS9+9OJFAbn6ICloJmlAhzzfRvF3/UQdfZAj7A1
uLCn+938g56UCqxCr7kH5jaQLnLt7r6CTvZE6Y/kVKEUDe3CJGgYaFlHS8QPaREfQBEEMyEXdbCg
9K8w6UjaVVcpabDjR3DkU0cuuWa7e/uqeJH+FIp53XN3Lo7oecH+86VLJQfTcaeSDzbSPzYdFqO4
2mvLm6wlqBpnBVHQv/IQOpie3xNAfm/pohvhRz9z8MK3U3NJ2BmWsIC/petNeADDnF9y5xNJnwL1
XIWi6VsNp88JCm61GJx/gToMxG6Kh2/0Mm+5gcTM6suXiSDqGTe+5So4dBbSTWu7iMC0/a2rlt+x
zEvTGU3ChtE2JKFWSK5xcriFWtO7gpAikubrRMysTrLsQ2kr9saWvxi2o0A/gwYptE6qTIfCUJLX
G2k1D3RhxmWi4AgAHZHFhOoXNK6UzkU4o8vi6bMgFA3Zhe2lDhMCazRgKDnCzHa+i9d6FZwfwBjK
ZbOj+s2tpPzq95cJocvEzoAIqxOv85yr7gypgPyFbwYRymLy6PFGwyyUGdldYGRqVey7XXngN2yC
u0qsxOkbE6FuNa6K261EUlV94uWXU2BjQmnY7TAtBladd6mBXB/+NRzjBR51IYjy5O7RD3CpkmHx
2A+dodURRM+8Tf5aY/4lb6WOS1GE/u1rX05ppvcHwYy15NbTEJBXckzSz6wn6ogBeaDT11i3sdff
dzoTgREkU/64hmU5WQXIEUrNJIOVb/1nKvAoDQRB4QasD6edsb+k9cWg5POA3zuuEF4mNv+8vbbW
tkeyoQHgMOmmS22OZd4+awyaz0H4vv46TCGVkT2Eem2UmOL11hOkl8EEUzdJ0YNzA+r3Mkr81v7z
5VnhsFtG/VcNo0wufjgJIdKFt120BAfVMhIghqpyzEIz9ctk9W5dWAg3tiDl6Be3DC1dNICq88EK
iise6A0ad4Pn6dzTdgxs3tEe7OnCmfBlUUtLK8Bb5NU7FJ5fxZ0WXCCdRigIyUUaPwIo0+4jjNex
5gKlNYRTyxnUVuoz3zYviPrsHDqIm0FNLrZjtI1bZaxbt5CriR9cnLbRpGxDuYII5cgA+EQT2f0s
pWLmcfy48EQk3b9nGGjiXu0CdpjWhmrgrupkJADQ7clbCGUBaRiDW8rEnMAkrmrl0wTluUJ//6m7
8ER0rI4OOuhKIgbnpOm3hNQAoxmxlUL79BfqZ8DxjnaJbtuv40XFG7nSgNp64TojxgQCbbH7k9Gt
/A44Fd60BMkxgDUYBuaBDUYYp9+YAHHahVmeyG00peXLj0/8SeLA4KvDuKLpB7S8zdGxmOmeCP+G
WeBR7RddEBITVnT/6nvdoWaBlIj5rlBW9ER/svvW/JT5xZPrMQOmaNWSjRgzywtpj9IiTGlC2G6T
XG5EWCaYyzcOmMiudtETTi4F23txafox1K5p/InpU0jWtM1Z7um+CGrKQD+kxCdTkrCpK9fP5bYy
XpU82OUQPCRJ8tU5TnUwn3RK6XHFa7u2hCzksA1dO6id+Jbo3Y+K3/zqByN7yliRnKiqNoeLYafi
YdsSmTygR3XCfcndou349qMP1ourbNFrF59U1c0WB/e9EW6cf+Imi2h+loZX/zOGKTHN0hYgRcRR
4REvfOPImq1ukkjX0ustyanYA2VTBwkCTDG4Yd1lrMQzqVlbSNlL+hb191m+P1D4AF4NEKB46w2C
yPe+pnJu1mL6LRijpAAU9UzYyABDou6wR+eYYrEw8I8JNz88h1CfXrCvUrchy9IL75KV+yWBaviR
FG+aB2Eaf8WogHVqKxE4fUYeP411Ey/PQudZyB8SK/lmAHNzZMWyf+9h5HxUuzXh8jHjwtXg2axK
s1bIAAYFtT30koIP6Imuv861Rtutw+z6dw5uoVCKqLndp/7+sBQW5OQpbdNU36n/2Y7KOzKuS/l0
PMU5OOS1J5pcJE+hQuGrgOkv8IE7LfInYDhRZg4C5ChZbIBGG7pxkG0OTc5yZN42/ZrgMm/9V0cv
NmIPhqZwD73vUI5eBPMPMnSTKWtih+KG5hjwVl5YMKigQzqo32HaKyIeO4bQdJQ/KG14uTq/u3MT
la7dLe5JlZfkZ+k2CXqaZ8vENwv/Z5X0cjd0EUEzPMZ6uHPbFoM1VpnSfkkOFllcDmjkKZ9KzGW3
oDNq+KTa41CX2En8KeCggtZATHWyyEhHGSX9D0eEvvdkBZ6QdMP+/ra/rT2gM2zIJwWyBBDvtgTs
vo89DhfAALDDkW0xV1oeoqfSmMRrvFcxzzecNRBaNij0zYZHDwZN/Xt3oYI2P9bJjbbkLVKWjOrm
VKQT5VqN/keOoP4nUP2Gmu8OH97q2Uy+2GZt0f9oYux8mXTnVAjL2Lw66mIagLD9NvcmjtTk59oi
J6Cgi/Hy+fnS5Vd2laOMAN4jV5aHnvnKKeGXlUO0UbxLmslO7rBoBZHGFc25NdmoWA9gd086B/DG
923rxJzJX+FaO9mU5E4ckJUzab3OmzN1L9cT9Wh/bysyLC4bFAizhDKBH5BMJ7JraYyAusz7IQKr
633TtjMAbrArRdkvk70tyqUirQfKd07Jr/4wKMLpkb5+zRw2Iiue18AneSY+M9VJzIvH+1AoE3ts
pVAxODfh+CksbQSo5syREWHdNMcraGBzOErUG4Yzq0zZXdCnkbYzMZq+GP8JYmb/JwbSh3YbnFTw
TTPG+aWI+nEsSN+ZXRKbDbiY/JCn43NUlIh42/Kp1YDEcD6m/MTSKgbJ5N3OGPKouvogbQFGGue9
WRAqIu6+iM+XSxYZzqKknBF97FFWZPIPXwKFFQ9VJPeFRZb1S8G0tW/U566hgprC4yc2Xlf1cFCk
YKTOu1UWyQ9nUUPAUvqlrJ2Ei6XEIYt57AiDqTt00lFiAuUqMAYiakmkuxooMiBtYX/+dreT0Oo+
nQ2Q/WGP2FXzTjhpA9CW2Ntg5WRTE4MIGlU3wleLBCXQTKaYoZouRoNhwc2F5hr3jC2KGwz8D98y
3KB49z0K3n8T3uiXUT02DspIyJGoUYHoqTsi7iCaNza+5YDeCHACfCcveAQIkKs6raF75j345BCh
TZxfq3FHc/V/Kx3dh1LSiRLLXpj3NnnpctKVxwQH/A/EqMcCDyuSMPROf8753m2Dkz+Xl7GcV9PY
trYMWd38mwa9R3KHRKJGcZ7GKJdMM7Oor2egUup9mgB0N4Kqhgm2WR76gWSq8pzHJk1np4ddBfdO
NWn1q6HLy4MSLGgEn98o0tJh37oh3L+dcAmwqmqj/z/pkvxBSwm7+OdaAfVN5y3YsMPNZ5+09PgZ
JYNh88SiFHKobePxBhu5zF0B+N4ZLN6Vde02iHQ/0ZlONOk60JgXmNygeDPjVM+psxASnvp/VB1S
AXwzKAI7lm7++ilMZt+6fe09qO30FdEsEzlEPnMWFnvtCjnFffoYRTxOXM9PdVkSuJlllT4WI6F8
z/KvAoFIo8LiELjBPbsf+nA3HFmK957aNysKI9i7M7P1bwrlRwjQbord0sATSyqj4Y2Hze50xgtP
VnS0wero4NJusRFVUZcHM/LnduCiuk4NP1FuVlDbcqDDT/v7F9GJXW6wWQVe2CiQGgjbPJXVabeK
4VlhC4Anotk1I7Hm6CxiNOvzFT0b0RXgxBMMJWQ2NjQs9KrvXZuG4w+yOzlGef2REG7JAFfwr258
l1+4izBkNdCl2bffbqoYUZPjdNBiNWf6ikBtVjPGJQxCK8ZNbIScsee02UCU4ZHbkz8COrDvSlqz
QZv1vov9ep9mghNAoIxlzy4fIp5eAw1D7MY9opGQr+64GD15DjaQsg+uohMzm7VX7yPanPJMiPob
M77oy7Hrq7fHu66GBJPFr2oSlhtUZ72Y2o/Pz8L1bDa15VGT9AoLMXYbfYoZf/ep3fUNjHw1SLJi
ZRosROIPcbNxuniC/pkoVdAwezEqBBz/j4X9IO9EgHzlDuAbr/oYc2QdlDStrPWpX3c6ATgXpJ6e
y7UjPdF7XU0L4tliF1x4Y4xuq5lGtowR6gJe5kkWpDlX8jx9C2bgn3TyVIWZVs/sokc7Co6SaGg3
ecT6itoDSiGmZBOpgAmqzsBqBzCOfIeY+Fe0GPOLUkkgkgvp9foBU9THaQJSC5mS9woXrE05aB9/
cXmfYaPGYjx41lgUeSQjwTRUYFH6qWnb9BYRxmUq3e83p4GHmE1eHnm3+3pjyGIkW9Jpx+0M4poI
AHm1XZSWOIAd/QdiEBJT6i6fwGjoqT+s5jJTeO6L8rEnb5D2SBwchR9kHQY4YNq79zevVKrM17+D
NlVwrPO6bpIpa+X4jBquU6BlSQkXlTI/qexf2/1uq8ZRgjV5GMEFMSNMww6DCIOph6ksavn9nY/8
mEckKdGVxtztgJH+qRJavI6Ap+Su49hJGUhO26DlqteGiRrJA07g5cFbjgQaF+hRL+uovJY7kAaB
WTsLJCM0kIHGV6HbyFvtP7hL3Keyj/Vc52tMVOiozdBb/4Fn1PpZMTDawKq7hRiuu7l8/XAS8R9S
sDmXT5zQUJssKiL5uLncu/8wauSU8EJBr2CDYVPhm5+H3qd8nbjtuTWLRp8n7ZCOE0NhUXZpG4OR
pl9AOBCg/w7Y8Hg4FBsJx9/7eANLIPoTeIZL2ft/279ddwf85A7D5ZJbotFpBuyBYr1EDIwN6xz2
eQGOBX1L0Hg+bZXeSCbC80fi4DUfRCURPsunw7rBYzdO4UaJkFgPQUdYQpv2QjFWN0KnrLgJ9Kxz
uLEucbCP1khV9Sx7qK4gEA8hcBPB7VygcIrW7whRVFAqYChKii/eBkU1ARtc9fT4H7h0oLJfTTt4
TlqCj+saXQpu91i+0+qaJDqOI4doDR9HdzrzDxJn5okBZZyW2Vneyu5LazK6j+HczqftlVXGePS6
N6uV/cU8IaSJp5GDPsXBCgxYh5ZYftsqHJcjNbhkBIgu0KpfdvLaJHxXVzFfCUfhCdc9RkpRHu1R
u4pUpahx3lMbs2XJV2/4FhU1UsgscEgzfY8EWjAKKRhRrEPpHkbxuM8po9xMBErOiLqb69dM/w/X
Db2G8kq+js7HCWkQXwieqxJ94D9goR2s2TvhdPd9/WFbBGKtGDrG3GK2SoIJBErIkIeY0lCbcb1T
fAQtksgDJS5mtEFxj2DKDkBZ2e1BoXCYoYaFp7yfR3fRVjz9NEryRO9V+5JIndx0YqgOawsaDof+
bnHsfuOIHt614fj1+Mjt1kjSEeHko1m/mDaWxDKFW3dyQL5vwQ0INPQFeqzS4y8mNTftc8a8AY/V
nbs9BBEM1LHdb+LORKXlRoOBNZYk16CaX9OLUXUyBiNeQYk17BCicmd2qyneBhNhUbDuQHRh8uCH
GnVCld4iumlNHv5yF9ZpfGmLYUrUc3NJzXR7TwACRqK1IC2oziwA/q4uHHn1i+D10H1pl8Ap2Rj5
95OnlMygb1NJQX/5ShQVOBf+fJ/pRpslogpD1sfMTrkhmKFvXbm/zFKwCW4rgx1nqHFGaClYUluS
VpYG/lo/w94iZmovBlQYCLmTd6QJE+9Xtmu3z9rObUZgi8/IPaykiEoYCp3WVJVEFA0elqSThAgg
dgMytSFLeEaNNj2Y7QEUpdJ/BSmwfP9ZKfz48pUTjc8sh2qTfvhowwUUBAAM+/6dtznrBlFna1tU
Yq2i7OkfX0chg+2mDreefzTK8F70UxT8+gdmkAhDQy++ekI4IWt57uhR1S+C3VAI5X6Taa/tLwPl
GgmcDaCNRAiQghDXhvyXOIGfRCo+71pV2NLOz8QxxobpQDWIAPBCEF1hIqecro0gieYOPokfIfmF
YIt02786pp8KHYJZX8hk6CUqbESGDZYQZDDG1Whb8oT1kKLNwZDDiQ1EyopYp2Xxk43sBq36msTI
yakBiCf48m7RQH1cM0gps5saF8aibtcEULZink4rFws5FweLdIZ/67CZggtA8Rn0gkgr1Q0YhAW0
2e5PH2U7URp+5HguQDFvm3MHM3DjeVnFmPacwz+HbH2zbg/czE9M1NYaQ+2uvC+J2efnUqmt/kgi
xVNjHm2oHqd+55zDlmPIDmkp+CztgdPbrK4cy/SfYppzHj2UED224Z2zz50DN8jD6wCFctjY9ftG
492fRKzKUW4uIAcJhCs0kTdwR1QTf3qABrf3OaLutG4sM2SamONvaR48TksnhS0MsduOaQtIrD/P
Nake+Vx3Pf2CB83cZBx6Ip2UDuI1p2KEaOPv1CG4wCUZoR7YrNMUcXJ+PFnraCA89azWVUMD0+Ja
5XdLZnE5fvRUdeodeC0UCL7u6OUZxMgxPPbsxQrufviWW2I4AgUQFDNKpO1E+ZyjpmgPBtBsmjy4
Y1BroJJFXfhNivZTCWJrVOEd8PKpgmIKGi5NFUbh78SG8VvpPAXYbIL0dToHvBEBqJVzpViY6Yku
zRCXcZLU0lCjucObQ4JtMbbVQKuACGZaoH+dGcx/f2xQ0us0lMmEb2DNbA8NoBZEJP4QAZ7xdkv1
H3V6daCd1ox5IsXpL2bIKEvT7CUqMf9kuoMoDhZXrX9hzSpPfZj82xJxbKUJmpG4nJCPzpHXZNUj
GX+q8ai5TIMYhQXxBxHq9T+IUtHU8Y3ACU7zu7E6cSWoQJuiqiN+lg+fNNQRmOD4Gdm0jpfZbqbd
+vy6WFr9qqK3hDhxIxHUzNGvy9uDc1rgeLq9FGtSWW0cOpHj4RwylmHW41CqtjZRV+ab8WERL4c3
QT4PZqjYgJ8XE8blzznUw5vSIsrPDL5N06gRnBkp72CYASECifal1BHB7Bga5yxRrkl7HYbp6g3W
CsyNT4RGoMmZLSHFsnaDOk/ivFcYhPIFI7/oe4m1kAS7nOcngcmR/f/juV0nv7fTKcLSR8sHB9Mw
WqHgpTfBnOOv7oI00qg6Pn7GT+vfiVCMXIJO5iaD9dHEF9od/yVFhLVMFzB9FEYvw4slQmBi87jn
xRLa5/4WxSYUc205VzDRsrceAVAF01Wht6gzTLejNwfLLir6gyBh/a05nURSes/3wC3KsfGtTMlF
sRlRgKQioDXvCwymoLuJT+of5EeCoPHDtkyKzMhSIW8jV+mVGw+XZhTrCM+NF1f1geMw/T17htIF
2ROH6yoMXhIh1U37LxwTHMONz976a8BpC+x2uiNJnN8xXN31Ow5xngWaZrZs36UD1/obBUURtUfm
dPzHjQdVSbSfZV6hvHroqi9mWqijvTEsf/MmNq7V4Xnsq+hFsO6jUVDt9fYjk5UknMa58SOUd3Op
aKvIU9qVya91pflioqyZBQ5y5JCNan9w67vXgWGQJLElMMU+qZ6mcNmPNDTYhv0jbt2QPPhKL8Ti
ZYyBUtUaEYGrKAJN2pEseP7hEbDV4mzPk8IM2+wKnEBN0ern88pDsZk8//xmJlaIXEiZnZ3/ysvo
R6gftC+/4e+PjKH2CkEx8uZ057Lc3H8hDCupZ8AA+1QEiyNPXMDl7ZG0pDqj1vpuHN5fExknTOwp
SqQWBrq5MKh9lwJlFbh1pa50BYXe9VQ8z0nUGaKMovldPJsTOudSOiN7tqvkv0tccsPFMVKnA+Vw
IcCZN7EKYXslwRyNyaPQFaDVJOI3e8qDv4P8AqvYVMpAociXmDeg598PCzPlrKHiovpatrQeQoDl
zRvCekwHwCyze/1qvWnTQ4EGjyXfCyBu+8xwWWyaGG+8wk9UeJE6a6XbeE660spB8RJMm6Bn3RrB
UBkZyjBXRRryH/qb6R8M/TSyEyrBW/hJLSNmsVuonpsWjzQ94gQ6gH9dfK6ygcPildJcb+XC7nKO
YRCVRv4SoWf6penv//exvRJQHY53ASBTP/5vQP6uuu7MpEQ/YDe52mcXnHDQaItDumBSJOb5LEay
tE8yAC/RmxSa8TsB34i+mEq1TukEIduz2r9hdXW4F5H+dpmVk/uAoQjY8THwHUhEhs/fr0263wtU
hABMhr2uXJgifBiY67yBoRSFBgwgVhwWgCsdBsSUXQeTRvBxSLOhg0Q0myTFhkRY1S/t4CyZcXxR
iIHavvDr5d7navinBTeNdUi2A8X2sHDXI78cleR6ptoKBuydhENWMxmLcTw/twQdW4LHFECbe34R
fbY53VpsAoBzh1/WzQQ0UT28rhRH/+rhyoNwfhtR6Uz1gb+1m2ZTJ12aGm0ibFNuktWA84xUpezG
+iPn1TANq0tju0LAVz/nxvXPMrLGNHq9TRj7n9fUOo2z41QwUopuT+CuIk58lCsrI2O/htEfZZBU
kNqTLSrPT4v26Y0EHkYhsCYDu2B86QzrqlOq0E5+C3JuqCFOLuXSaEe7kJNZchn3F7EZ9aUj59u7
kIrXYN/j22u5tRUxE6EaHbMUWDdY4M+SaQxvfK7hYvSh/vbnCkiGyw39OnwmuUAMH6eQqX/tPOTo
MkHLzEPuL5P2idMniX+yHlhcDZnSLpio05L+UCZcuA46JIcG4zbvcNxjIoyahGOVDpd4Gr2vJ1xe
lw8DIJ43dQZ42taHTAgfgrUVh8Gf2n9XUxKUi1X5E+Bvb63eJmiOCBZLZPAtBkdk1nPbyrTyLPiU
UnSlYkv0y6sbjXmhHyC1Zyj3BXUBrne0rE9mpTqzz4196v9f4wytzyBQkX39+L49eyr1jNrUq7Sn
dylYFJpLnR+fplx2H4Ass2lNg10qgNV+wxqrj1HUqqEP1R2SEd+vIxct2sirCYAlLhqvvD3vEry1
OsYJ53SZbuVjfZG3c27cNkWqGuMFJQ3BUt/o6PF5DH48FH9dXJrals+VTbEMoUUzIevBQuLc1Xjm
QiyJnWvCTEuuB3PGjHaiCeo4njt8j2E0W52EnfrvFzwIQ+i/x1IPEKEJt7UpbtboYJNcAJP8yOyI
6oSIegseOiLB5zAgjAFZnbvh47D0cWP7ixRwKY4ls743jvjxXNsug9QNNfDmjQc1Q+85aoRsMqyu
3s3t9aJtJLiYB6044aIspZ4iqOeiutDdWUHwWcaFBSgqyXAxO13eGacL46Lf+9HT2KHk/6Kw/yQG
WhJEx0f2gNiJnsWzjjjGXUCAJp23azW0nRNnn1atnh1TYAsIOBv3GoX09JaMbh28EMDtJmtoZJt0
RNsdrWtS/vpaFaMsVlaiqIn+EY04wMhn2OXYFl9gujMA/rtzHKSUzRLU0lfPIFLj9KsjuBcTr4DP
UXU24NkTkwnMFSo4Xh1uzrYEqoGOeJkfM89iJ4xm7NSEJSRA+v9xB2kXfQPqSeSStFN4ft5isAyY
bypSscOr9UzgwF87xQT5uMeRqx/16WZW7tPxl88EwRK4+DM2luBRClKtX1CrSUz6nsr6JIzU6T+J
PEtOToKv98Ssq6j3uVOh48s8Dzz1ADM0w2GycZxZfUyAn8eXLSSsk0QqGF1cY7TakJBZJLfyHhNM
W6AiQIaYbbpso+lwTpXolP7RpnTLX7MEFiXL1F5CMioq72mPkeaQKUVqjxdeduGUtXKQDG0CFWLP
7mA5W9tBW5Px8UTuVPCjRq5RGGbaPDmcTfBMN93JCAiDrPdGvfYqpTpg3BWsOHxwKMobTseWGs4Q
q7TTsIBMUexbyy/Ov8EE7TJXgRR4gu/4q9GnNvuOP+gAFS8+bhIF2P+Lg6tGz5/uIZeq3Pza/8ps
Fqi7D/MkWIG4ZCdjtXUPZzIKT9QX0cTeJrzSVSSRCLxcZtHLgC9ZLlY3dm1bVL38KGc/0og+hOOq
084kmrhjegctVQmXpon/KBTHXBVsZp2NuedkJ6IOn9916tziGF78QY2lFxHSMyK/IAbQNN+6dGdY
S6NWvtx7enGgcXDkLZ7Ly/KdULR+RKOgaGogqs2sV2QooJ/2D6V1ZrAaYefIjcLcWDERLtaFYTre
lmHhOVpRy54u7/arKaP0b4CHobHArgWFpGdrIIUH4QYGDJHdyaU6gpY7L9iECYuhkIXCmru9Wz78
NSk6Nx/beT1QkPTbM4KG/avn1+Z52Nac7Krsk8QC7F22pieTErVlMLP/AjIlnahAtLey+xaqeSyW
3s20BaWnh9+fRACGYpPOvxiuKzobhVMkJjuKaXmgGQowD14q43ihefdY1feC4fyefrBw0+V7yU3+
+6x8Nw1mnt8yMcKO4kvoRGVRuTv2oyDilwY7wsWQEBu1wYr5kiBNcs/XSud1Iy3zRNzQfXpyKka5
HdoaM3CSHQ18VaF7HvXcqh6GAlf5OTF2V3cHJMaOI9PVNXM17qx8C+g6ohSGtOXj6Z2oR7/CdlMw
b3mZsirk+Qn0gCWD9rIHGReqM7byM7SF022OjQDl9WpvLbWuoQHwXU3S9KGaSj/HzgrJdp1/0P6p
IuwSYYfaed/AYsvHyQzOZRyfHIlm7q/rgQjQGQvDh8YWqXMJYBf/FmcZqix88J3vmKfD1Nxazf8R
nTKpLat+8fS0kCUkbnupbQDAjGQ4Wc6tZGWCzPRKP9MCbWbc1APNYTqgxH/1L6/VQz9XwGCOpQHY
YQDSvQg8xHgzl+NtIkfCbXmLAUa/+rn9MAGiP/ZXgNiP8EUt5EqS2AC14pirvZnUJywbWT49DrrT
klU10PR5G+K7AMh01aryV1wYJeifuK6ARQiN5M2CAtawNlpj4Wyo1ctpylDuD5URnoBRsTsVYa1R
KYlLk9IlKGg/amV43IzKQSQ+11/v3YBt9LZa6w21zSKpUAU1EIEfhe63FWTDJ0NW4vn4ElHteNup
2X49FJy/sjVupvXBdHVMyKMBf/gTdtA2rGPrP0i724IIfuqY8AZieWvbdJzuK91PfK6hfusCmgQh
bjVGljKSeDkNOt8QXa0s6mKPbAa/NyG9UVfhndZpPk/e+uBUmMpB4+QXB2bdCAZj5XO5itoCugTJ
DnJVSf9jojR6CJBSxQ66/BGUaSv8ZeFLad4gCrkcrwxTLwQp7LJgSbflq2t3j2kSnxvZ6MvWdzKO
SQmAZFXi9E5TdQ+gsqTsedTvcqoAZCLr6rEP3YtKXILJ3bupO11G68tAt3ezw662CA6czcWaNUPZ
g+dOLC1s+hxPlLwWiDRBdtGU6Hun+JZuu618dWUERn8oOzbuFGoHeB74qrhsy4iaTYeqzf8J/nvu
7x2otBOGY3FtVWlTUq4tLELQ4uU8CGgZZSe04o284VWP1dGmi3pM3iofyc0KZoRMRVDTSAvPiTbn
d06BuyfsD6uqrRVT/4ShexHldN+A8tl3QhnxHa/ykWoSqH0sFNNyKpWm2OJLngOq4BH1FIuHdTPa
itMDRwvrTclW71W1XLc3V3B/9xCc+X0V7BWOp3tNhGf8pOPmNjVufgJ/YdVq2T7fLiz07phE6Fvz
mRgtLtjcUYUvPYSgOPcZmwGhQyeeOa4fQmDKZzZv4L07tcVaeD4mlmAdL28fnp9emgPweOZR/WVb
QCD9HwggIt+yGOZHbdgnZHhbi775M4AxQk/zWYO0l2EmqvirC/3tGNQELUPckPU1M+IP7Qn7zfOi
728ghVG+2chkZONMeZHRgsPbVnB50ftgqvBWyclSXbtNcKHlwrZHJ0FH4N0PYOnJq7TzgNMHG+Hv
Yz4gaKXrkcGfGTdMYRKJ7xnp2nsrQ36tDXQIhXeaLM4fl2iQWXNbn8gXvlikKuYDo0Uj8IMe8WXV
P+Trnu2A85qiZLDDAdVBR45KSCWPSZkCGoSiAa2GCYqqMpWddz0UTK/i3kmgaDLcGTTUaFHUIs8n
hcPN1Y9TSePBL3lR3aYgjDtPVx1BOofAQDS4v2Dkk91SDZdIY3DKrE8VfiKnJSWHTlRel7mE3SAc
rGt+W0akr4NDXt6Lu+SqhPeTiTYqmw94WroBOzF0WrsRljwXLDbO7uUBm6DpVxyPJM90mn2HFhW6
E7ogwhdSjAU5qsyl8Pxls8UStL/ikwC9ACFZT8IxvoQJQkHTRVPwZHsTIpOluApa++r70HCBq5zT
ZnZBNVc/dFlEySOgCFUPi2w0bzsMGlvCpS4U/gyFxlAvLqC6YXT6kBZp1hXp/q89Whlh8T/wPlUF
6dF5by48ixcFDQyjCaM0CAqo7HiDZuJdHVgHwcdQxWUlQvuKfvTJ8qSz6OAdCMeHextfrclKDMCc
0ksa/zhn1nnWmFy3PUzxiSuYv4ec9aKquI6o+5DByCqZCzeyRuYcL8T45uqHBVE7LfGiFZMAjr9T
4YRQgiyULdGv2bMX+O59ygX5WsI/r+CBC3qaSoeQOYaIIr0WEP4qwIigf4L5ICv7Vi5vIwSLolzy
n9LAJNXrc+2UjhXPVoV1eDCsYOgXpzzJkH7uJDhRave1XxhDZqpZW52odwbwUhNG/skvZUI1eGCt
BJfuBHscy45gn7P/OCpAgqa4FU+Cu5qoeH1YOObyje1aRcXeTUSy/LU3fmJZuoSZLKaexD+baJm6
qscAtJ33Pk/hc1RSvdstM1xPpXkxqhdRqPdQ2wa1G4bZnNuE2vFua2szyB63ECpoEG7pprseDLI3
9n4BPbLbTIWnFvgem/+T9ZzylH62sAH+yEqR4JWH7asg5iitCjU6VoYSeLEJAjreG9YtNUtlFjb7
gkB1+pw8OUlZwRk8CVvl7ZSaYg1egjS6K46+mVhjIz0M/Ja4eCBWQxi+7hioZnVdbfgfvc2dCjMH
92xqz6mRsoJjpczq8OgF3V61oC8XYbmFdTQJwRC/2cP8diP6Wo2r7r+Qmm2Xm9gr40cVJZ4Oslmt
zmWzAWN39ozoPNf7BFGoJ7SrsRwXgiXmB6c7F//db9iqiYfn8Z9V3GNj8MJgweKHCN2lCHpeHRHF
wvA5TXseiQH8i7eTX86ggccsKZuXVOt9sx3dDioyzh43bLmVBzFb7aGA9vUDJkAsAaQJicwQy0fD
RPq0snARTCgP4nKVEkQmTVmNXLbiXgGz3DrgMiDHrIsflHBKGKIrecwxYuoP6KbN4wUtyHXaH7vJ
SoQXWYPwl8bLCqXr24sPZBVMcj9o+qQpHv/NC4H00lFrusm6IWT25DCe9LoP4G6TcSL4bmoMULap
jTn9SeFRvZ3bIBWPCTcd6d7KDHCne/CgqvbQ757LO6ETFGnUCKlkViHMiEYfkzunyadIet2OpgEx
LidCOWGt3pq8eV6qNVTx0p9J0KCj1F7J8pP0/Ft3cmxd11h5cKv2wz7/arxyyGZBKXBDU/FIub+s
xi3mFYIMZ0R20aZTjRBljFnLEPScUbWxpsr+QlIj+6HQYUEZFMVRVzVM88SCdvS9mTo0+0bFQ36I
bJKSApWe73ZhMNj0WCVxG2Yg9ov2afhGkNKvbCOlMLBqEP53FVEDa5icjT/Tyx4QpzmqdP6Rgw6W
P6CNEEUTsDfbbaAjAgAO6qtewr11iZHAxmdmD1nESpExVhGfnKsl6hS3YR2ks8PQInFo8fl50ydv
L3bC7FWHN2Zpyh2m15vxdCdTltug9nYVO2qPUQmv+W403Cy9S2Rqj2ntetmN9rA2kuAoVN7n+QyN
ObEu+iiiKmlWeZ64xxSVU0kDfwujBqSagpobbqVjaMS+W2AnNgKaToMKYUSH2pQYRLgyIBfr6T4W
e1eZ8HkQdtiE/fhoJ1yBScjn1N15t3zmkDMq+MDcP3sicqBvZZ1bc53lp0vsrK1E6bygGup9TaNz
7WmKtarksO6jn1pl4+JUm4UqWxARUBkvl3nZ5FWdz/ibm6Rgk+EJ4+kuYTjfn5eLZgF72w9q957p
RXF8THyWDlgqqF4wPiaz60PYqa3gKQu1eOZHBZF79MSBXa3DiTxkDgVsPqIh8Q13zJYyyeV6gLe9
h5wOFPWDQoPSCXuGKQmNL1vjiVXnhE1iZO/kikufxeN0oteBGVZg14/sPMZT4PxB2agkMGNk1eKa
SRlbS7zvnRvZG47tN1bR+ODAUS0hvla/sbCfv+t1us8ETtMA/muC+kDPur6+5fwdsTKRhZMDzEaC
pf2l1ggTemrMxRNDjpbUgnaaJpZK2cIrdA1IFE5IegjiyBDsJ87zzi/Ibzx9y+adnHEdTZsAScb2
KEOXZk37shEvrLgZ9n6vziWJYSPbxzmQVmDPcuqCSi1PiP3DpjrXKV/jbYebYA7qVbB0ZWdOqtMr
B8cv63CqDYr2xbqqblJPROArwsWYXQnoe4fzv/M/HIjVMg/cWF3HY1/C7AckENlqIHrSXau0RRkX
mjVkhxaXiCgt3s1ePYeT82E+9Sucoa5XvkLOc05p4fZsQggLu+U9qB5aivMCsFtaSCjXjPXHWD4a
6Rz9INWowq/Ic8BF3AQw14K00LSXMxAPckglfrpTfyTIDWYsaEDUyVYnZI0n3O8eftk+3FLQ6XGo
eVrGcxmMkYOeZV517QqRIoyyTNKaoJDJ9rPEj7c2dRJRRzhkS5Qd+NZu9H8JHLkMdBtoQ4uGLQx2
tvsFl2NjH9bMwMEQRhzF1L6NnLfoM/ohsjAlCysi9WsN+slKhae1GXnr2tGmJeDeqO9yKwx9C3WT
hAqz1mcWUz07bcnWSq2Z4f3MfUCnTTni/3ZDm5HvXq/XMnEWKzYsZJweZxojWNPpZcUrtCQWXyJJ
J1z/+ru+cURXU7Jen2TUOajyUwXn71fDt1f19ufyoU5QvU6UuO77nNapi/nCIk7i0rZtdWfeHf/W
ZzfKoNpPjXUbOWbGXLzA5oJC8fRpAkIoeQv/o1pmGNvIJIHw57RxPFycBVinaQmPocQOTv21o8BA
vH+WDOkBTgb97x+GvgntzO9IVv+y5pfHEjdiujMK/hknp1wmTXpgLXvwb5AHbPykwXkjhoLyHSF0
GRjUO14zJx1ZT9HK7BOgnlEKmcSRhFTE02CfxtFQA8I2VrfZ1AN2XjfOEJ+pto1WrHfHb7Wmsq/I
yMRXpiR6WKCHPqGGEaPpIvU/yE72BN0fVfyj3L7SCc0VkaeydhUIv8om/kEx1FC5uE67uaSpjeCz
PfTjiZNqRhx5LKe0tK0O0ApF5wkJjdbvsUN9G2VogqXZhGEO7eAd+Vjw1RJJnmYLIHjhejHzS1Gr
6/yE91E0ha1hOZZc+PfZT4NfwZmby9EdApCbNdW+b1c1J/wIqi6jWfw520uE+qXYIscYuyz6Hnz6
FjxQpWovdKlL97OrYYLvAWMLkUQ6eh5cM3EMJ8QKrZN7/MdwMA3bNwPNEiplOeleFU10oXmc4YOE
TOIZOizgoaN5jou1cxOGFDjuUL4ww5oMod5cfWSbdEazweOPOLQIbwhIaZ1f0skf3DLrz8ZTF9Wi
M/BC4wKmDRDxQzDh0AofMmPzlZTkjiCv6DWq0AAV4iUeuIYb5CgvTMWcGXpqsrmnPK5Qf/wdON85
Yzzs90ZNxI7TV3IVntDKO7mMCivWTLjsAkDVoU6wgzcjEz/IH1t08eEWpw10X5nJb5UtaA8PCBq+
EBUACRAiWQIHCnLS10pylNnnCFOKapsu1aepETZxkpFXJ78nTfGAC9MCWn4IGhDz7TO5jCaaJO12
VvxioT345EAtmlljsHQgJbIB/vKSrkmQo9aCFp67j2QrqiTbhYMFirJTg8QBcKRmBAwcCclOYURX
4gyARCeM23RZGUcpZ9TZVjlRvWyBU0e7NvCEWPsEZa6Ni7poTZ0kr7f15d50GoEGGVUivlophy/p
izvgjqvu8Zmv2W29Ohz+qVgr4hQ3a134EzPm51WKUd08jthouHQ+0I4rQiqUG8JjMZmmO+QUkpP8
FtuoCOShSX7v5aZGXOSTVnXxontIpwwA1/jiZRRqgDaH2Rzj9vO/oVgghfX3szGuzWZfr6ouXoMf
WtdkciyAPZNriGybGofKIVjsTYAI7mqdDxpggoofhcaCt/0GrXOkkftn1rT+KLA8W20TpAL12RA4
6ca9RguzAFBDVNZYps1Taik+rDnHkVLX1myA4IGGwjnR1H/DFzcMm2B2kv+MotbtwVMAyRtCWmzY
Dyp9A4xAXRRZO86IOpcEKtm44lWtPYVR4N/1Fke4UC3YplHiNJo8ff+6kbN7D7/U1roCF1qxFuSA
SytE7NW8636RnJy2mwZLtZPzCmnLMDRg/744gAbwzb7cOlNuaag1fN//vfcUhfzCzLuxR4tpZZEj
49BbVEwUdKNdpOAOkIT+QPwYfruV6M3eiiSly/LqUxvY+G5IEpboHiht/W3QXJq8JrrZYfY9w3Y6
Xe22Gq9eq4Ib782S4whT3VNO+3t7MH2cYyXyq6CCrp33Wwt0zSXX2R0EYLKgCn7fnGBid6uWFhrx
i4xPMs/+q+Y6XxPXKEwn+GKtjonw3ycxoNYBX6DNj6M7XRjQdtQLlv01zFJ/4DK5h/Z7M0jCOdly
nxBKRnJy0aoFg0j/vncwVeJFzgFaLsCocMs45T8bwdR6bf4KzJjuUkL5EFAUZBqfdYOizw7wyNl9
lWFp+v1vjd8VqSFm+6QwsuSVz87Bp0S5vMWRWFCfP3aWAevWyx8Y5ZtWJSK+gsoYOIbu93AVmkju
YyHQsQTRO9jsSWouKhaarZGCxo5qvANyb/fv/P7bJwD81gx8BaC80Cp/PP5lRQzyDXRVnTpkUZB+
st1VNAMdf5vNig14XF0z0lvfse9C/l3Q+wqHjc8R+QxA/zU4mbwlRExhPf3V+Wv3K2R+SpJK5fy7
mHoBs+o6bU47uzKVfy6LPJl3+34YCZYIdgHj2XgT1jFAG+vJECvlV5qimp5/lyBrU5V8okRctk6v
okSiKRkRcb01eH6TiLuVifCEv5Yg4rSj9H/HMPKywbxysbSBriFz4gpLmOCpSeZ1dTKp8B8piJrq
w71+WP6ECxMwyrbv3UhZGEuP87dHjsF9MhT2+CHWyFq6gJPwVN90glf+JqFbmY0XAdMC6tceDRAa
d2vQwUGMxGFs3TO9K+TfajGdvelYeZuk4u6FjvFVnPjZrzPkZPKWR9NbwzF7nVYc3YiBqJGohH0E
ZZqt+lTV6d4jULgxp9OeDeITZ7d35wioC1Ymeh4aOMaR03jUyliWyGWskKZ+NW+MKfMBaPPkBzsw
bDd8xEJqDsrtxSOy/dWa3ngUCE/URUMvZ4cEtzTAJ7gMFQKe32V8fvthjTfhTX+8ZJlITLIL3ZN7
r/k1mX7mN9XNMNrEXMfevWBXSJFhp0rYohM8fzcr0WQ2Qqj6fTu6vYWGXOp5fucIIKziq6cEkMCt
HIqsbzo84vgQ6t0aAtZ6hPOQM8KVzkgwc4pE/9GLs++oU1b8uIWmh9IPyavNWqaoXvr66Nj0d9O3
aERThPVzz/uec+bn779nXehTPvOrb5BAVN7eTe8MWWlXvyXcNnwpPgHu/50RI9lqdwu6GlY87szN
Kwz11MgiWcWB3ItCdbpY1Sste3hkm53isD6KZZPNSiThS3vRv5HfM11JdtTIlXsIqhNOYe25+8SI
EPgAvvgQRtsWMgVv8DANNW0UuOc6+vM2PhxBWwNRhx493sJyvk8uMqHftiufjFtMP+jRslps47pv
FogRLjvppFAq26VQiSlm0oSxVdCId6r5gH/GWucFuEDDU61tyBoVnBQgbyc5VZCBDoiTwhY/F3Dz
elq2NDbC77PHE/U46stAzqavuAT1vHAFu2RVwzI9QAEPo38MaNzQ9CqEucA5kgp49bsqlZmz0g3r
qPR5byVe+z2NYyTRdoahHV2fNpQX55/KdcEGo5V8QhZqwMbIcfxEq55cYdqgBFV40rYE5IIMhAeI
O4uS3UyzOYshKaAoyZbKHQ+MqVOocIvrqa/xQFGReCH4b6OXLtFq3Q3ZnQJcXj4nO5cW9ulhP6qJ
ChpHsiRk+diy3htgr/UKhAF1B1Q6dr1uhENtPGUxyWVOp+Ogx8dkZwO15gnPxHzmEJOB5V1Ue3zz
f6HFs8E/ofFA+E0CrnbCCSO9lQvFWqVF46KWRDVgoszNuVPFzv3khI0FAqMrMPR347wlc1OzOfhi
tD/yaDNI0woaqaEcSff5dOt0/gYyf0eNqDgqeSPbMp1oJjrnrTC9k7oqvt/7XXEdL3PktNpCkghD
r10ce8TNHZ9ctRlUsceBXOC82GfoE2ntu37QrtBFcEt5V3iBnssH17PqV4F7KECg4rCLwqGysOTf
mduPMGunoNNj+IQtrl0YtqtlARpaUJTLY9bUPqy+hgCRT8O6sNj+q7wvDcdmrvrGTvDAtusFr4g4
A1fZlNQL0wBBdngB8/EbELMJR0mmCdroFQvTAAdRCCUlZyDSv/d0W43e/dj9zYzqDeND01YJE8oY
YNtaTl+2p/eG009e5dmsCeugOc8o8CsM4N3ICfEdnN1Exe06AVHMDX9z8dyEqPVadrVH03WVToq9
mKPt7rIFuyvVc/2Nae4wgdpnzVE6EyeUVM1wcx+IdCJ2XAG5zXeazDTtD5qLrWyonkY/W+PTmQYr
2On/WdmABvD/yoWst1pnsgXjLOA6qrCDegxfX2mPh0aD1mimlDkXxxCOy9A4O0ZYnWwitRYHcvUH
ZQBZiXJv30NeEu8eKAOqn3PVJKyqgbt9xDYY4AgH/cYGwyhJvCc2LepWlUExImOOg+wk7OceF+b7
oms4ENlFQ8VO231Xjy4uIV57juF9aRlw8TubpaarlRrHvINBWPLT0MxpYdIBKI5fKbAK88WOrt7R
k68DzCimTxddjgxaCUefcNwpOs9a4w267UKSJGyoSld786pRZyUmE1tUbu4ux8Lwk4aQ4IJWsM+G
Wfj3jHOZuJUddkpru0T8pj096A3wwihzV5usfsTSb4RWbf/ohQrctHgjgIXjcT2xYrbFNlqGWakj
te/iVIjr1XutaP1NIhRS33dHA/ilL89qhZ+x7jtQhKe8QTiZ9lyMkgCAEhLYb01Ti6WmwvGBjsG5
Ph2dw4c+LogXWckSQPiNbUqfi26Xm2LEKVn5t42TAl8ank65PCRrNpPAIj0QdIsE0Wa60vOUazw/
3cs3OcDrtkS0GF3HVS1LeM0fwgsUkFhU0WwsrftZnkj2qC5gv0cIanSRhqja2pSqdKukvsFGitjo
2Sy01fE7nKvg0s6oXsNvEq/ymg1xOWA5Ze/vkQwMPt9pGdLig4kV7vB/mgW93+u2rL4/FoY8krKl
wBqPCNIz0T6gRRI9qVWqg+WJopQS4TmvsBMBd0Mf/GygYcE69QsEub+LdQglZQVQ1Xme6sIY9B7J
4mtvEyvvLqp1i3hBySJAXujJVO9JYyZSu9iSL0zkBvW6meC3GDLW2jrCad/MLfHhLIjTmlGzaWfE
KmK+qKOIv8Aa+vrSTiDaLT0h2+UMXibbY6M6GdIA+GcVa88SO+QboO2rM1KsPtj6z3hfH94ab3M2
rDaLJmj3dCtD/VtuGCKmM9nm5dtAIB5W5mceM2SWW7IeiIJbwL88rbkjP65TdDYmEQCWzHDvJWin
j11wZPAytuTQkzqUMxjtoGYkaWAub7IxEVtA8HkvhY+T+kozBNkiD7Y3Gtvh+snKn96VugvbQ+ue
1tvjoRcARE2f9BBg1sxByCmNY8bigWrcpkjVW81vcWXkBUVOB7IodcAF+r5YPYnHamyY1m8awIYz
hGj2ArQ0wXpnnj6tOyChbfPHXGqSimUsvxN4XBC3BvoNayM1GHZzakOMfKEsA29TdK1yue2Jk9WX
msD7/CBKy4OvFdmx5nzvdixjeyos4eIQowchWmv6aO3zRUIHQCh5sIEjOEqfz6OP9HlIGmLcOE/o
bX9yFqijjIv9QqXQonD41nEZ6/KmxZWQAX6Ww140VYou+ENy/K+Zjp3E7jwJjPHlcdD1FQqHacRJ
y/BK0VwZE2V61dwcIjgY0Pd5aV+KVzcQJDWcqxQchd5d/iYyGQW9F5QfscHi13/9L0iJs0X5vVbk
7kNJ0JRPyRssTqrejcqC2mG0Q/ck13bNdKBEuZgl8yF6N4MQ/NcAlcpEvAtTsLmKEWa690keTVzQ
pHYGWK9MzzLfogNVj2iBfGLnOrPwqkdPw/Rs1mD4MUUAKj5aOi025xcPrYloZGd7WSB85HXgfqI6
CVogw5ZMC6cEu2sMBfRi7XOZCE3JPYEHKT8BKxgaa1ei7gR9wBYGRKEjZRe1Z9OnrQ8b2XyO9AsG
GT0O0tKSxFuXSY22grLoazeFiGUNydBXoRX2ubxz00WSv0DapFWqqj5e/XrmbwJKUXg5vkuElcex
y0VDdyz8bI36Dvk5PcZD30JY+my2JQLlm75Cjib9BlFlPZXnnB9NOJtjbUxuIeHxE3KrACMljPxd
r+TTtj63wEssU0ifEb63X4Y/EvVjIttrdCZb97eNpIUzjwlq2nJjNNLd5NntGvL+Swaojgk00V7F
kA7jzRNC2EUWAgIkQxFhYp3VucScVznv5dHRtcxNakJgufMw66wLCsbHFtFy/bBFVq/hCTuJ0FzA
CYWvNp4SQsu8dV0lAKqBzmCWcLX1B8gu9X8JgmaXkU9RZlPYON95ErEnRcZz2eK3Bu33JcYy+xxj
KnJNNsyq6mGrqIHoAPNrOaHm2NAlLKRdK1QlFW0HIcqvtD+KKrNokrYD76pW+NlaZ6vSsH7b3242
KJ5efGOrw67N7LyCaZdK8mDx3gvRrdiOT34tAL65or2MUEQuCv6apfBba7KZdTE2VJpcSsvMg5dR
4ge6dm25v5hcOpcyrEvnojPKxnq/9G6WT2FL28PetX62Ihb7/Tws7g9IiuR/g5BS9QDWCQpM/q1L
JE8ufbHecAhV1BjmOlvYtH6I05jfbCXdX/KaFcdRYrgkPHUwtHSxP5pJRqszLKnXRLv6Rgf8Wvoi
5iYYeHypiq/Er9aQLwFfyw9D63kWuAf+k2cvt98kcRZjCBUoHhcl2S09dOwFzafIxMgn6JTOQiV/
5dlSeVVTQ6yxp7/4mShVnL+DXLAk5kXiPixx58V8DFanBjsMLqW+QkR3U16jQquGFYBN8R357JnN
ilao1E5LzPlXJ/Q0idgDZ8qnNRFms+SANd0IWxFXSSxEq4qo92qLdQgiVKImPdvhwaTFJQJhWhNQ
2im4g4Rmzh79Rq4PeMgsYapF2106o5HKj0lJx9MkHr8ceIr6pKeAci0CTiE4tNaYJJR4kBFzuTKb
SQvVymWP6h8jWh4Js8Ip8UVntTiUevh9ZkOBfhmHRmrQqJWrYe1Jme1TU+o0CBwe48sz0/eeLhpF
WuRkkUlcDHUrLSMMpENYEtmvxxrRTdGmv8jbTYGZwZMmih81UGo01MttHzjJ9GhQ9qfal2nzJC+x
mv+KQzrmqBoMsO9eQGLDfjPmvGarRc4fCnFgkBxStVM3Eknc72V1rkWShYk/PPHDCwF2uIIVTBj0
hWt0NvOZNjXk/xytT3LPoMnSC2ToI6/j+mLgsiDQc1nu1Qq3q0nopdJwHRVhzRCnxuREOqjbVjZF
SHTL2cIFQ2ESrgW9trFgFEM+f2o+vhkSLg8KxqfwE+gejpqY1aZBtNIOsx4wVkOfVKTF6eV8kNAr
9+dFZ1Ku4YGA65kjLUutL5z7q47RHkHNydiTTVET++FOj/3ZmeY0nL/G1WrH027Vj5uNK+KyZYnH
ELGaFpI/RqM4gzoYPCTdIAu6lTz4x3bZG8HXDkDzkg04Hik2kqIKTofNlQr0jqKKrbjq1nfvUTUJ
W350nXYusgRkYyOScqiHM9VvzaTJDCjPVSShEuO4/pqye3vKrrAt9Pk3gdY37wXk7uRbFjkKuB4f
IqvR2TaOTN0fxuYtzzVWE4OxVN1B4TE1oZEaRgbL++J+SOt9h6vPIn/kZtRX9M/17FWBsTYmABXU
6OX3PRRqPmWNLJXtiadMZ5pTpLpieP2w1ynJfoqFfgSjTO0PbBEc5oKjLk0Qe7FWvSdldH6DRY/B
cazXa2P8VbgZikc/yp6V5xxXBO7bMlWmbIrx/iHQodfyYpIxrZQagE9EvPZ4yhyWWMXVDhaFEERh
4uhtxPMRb/DbCWGXJPhLEMu7K0sQg4o6UXPou7gGp9NxadxlqHT36HiOZR4FP1FIbGoMS4k81G7f
jMlK/Wma27xqR5KV/oASMBg330aKZJknpnwlF9FGrluSKPxSo8oStqGHVBp+k4W0eJ0USaHpwZl6
kjrXobLUxYxTg8Tp+vecwW/kHnfb5ra3Nlr+0e33YqYetm4zren+H3QOt0a/7X4+Ieytqc2iKJZP
XFf4Q0ImRLE+4DSoT5xGCPDfddckDoo38ZZo4YrFg0iWsIlOGaTSu/AknbYhoJur7FXA84j3jqPy
kh5EaFGOXgMkS9d0nMKDAMZzvGBqN0AwX1ZAwEzfcQpkpso80+S4uU8Rl0mw1vWbb1w/ByKDYiu0
0NX/e58LnhUwZletGRhFGVWmbQh+DgqNzIjCz7YorLLyYjJ6mt7frBpMlFejmGdOp+i64Ztx448H
3QdgQI//8vVNM//j4f/5ZAFkr92ZkS8t3kFZvyApfv1G15zgn7w8KijssXrtkEm5tdiJt0Go0zad
7uRkeBmmbbqw0QQzJUmfuIIFzwToBwZ9IEnl2Ag/Za/oH2ami42/os5z1WlpJcsXkr7EViJ3CIzP
GmXMSjPtsXyqQoLQ2D9XEhrTQViNbCMFiZC9C5bLNl8iEdzjAx9/5BSU7hb8ye3e8OEVDGe5sviW
iFiwni1R0aq9glQ1/1fRSWWmA6f8t3mkGcQjoK24tIrOMLkYaSF6lgyzaWaP027ma21SfF7zQpV7
OUQPkOrlZgo6eV+N72naWV7u1u58zyqY8Cv0vGzthxxa41i6rKqVH1kvmFSUmacq0xMRHgJ1wCLk
IJAmMXfdn1911iTGKSy0GV3ErC71hvYByzftRZO41tt2L9nO4WBL7xTLYmleAk8DxlRKDodAd0zU
C6RA2G0YEgpND7GIWsuuEAnYu1M7rhc1Q72NlQ1AQvBsCYSNRzj0YT0HSIr0tsejPbEqN56If5rr
a+B7CJmrJB7ZsDsfVqBzfeoqDG3M+a/BdGoU4FRyOSVF4RBbYo77vk7Wu9X5KnIBEfZexq0vLceO
Uzl8e1W8Hmb1kqSCWYj0x84zH/jfIF1A7ou3TsOxRN4qs8MhP4hDKwdvJ1wpfhqULy2QpR/btq+p
EHNT5LjCZkEomTHty6l1yFmsaqPJI6moRM5kHjnVanobGWC04CC8Zgnz21qxlUX8NPiCuF2l57sd
KIyCnn6LK8TMhe1LZJ0aNdZNgCbvQurF3H4RRWqDMae2Ys2LCc6cJLVg2ehntLIIheZCDp6gHdjc
3u2u+/xyElv1FlvWfV7Gm4p2hHxhZSXu1x2fTdgrZeiMHUb2nxTIZ1HnD61CRz1s1DLwmejaBsXU
MXCBTAv4n4UdU5+ei7ZsOIgko0Ifr3OTYk8YyfXa0HuKPYsOe35GkmiP7I9MeHZey54RbOBO/1ZH
4WPho8KmL7Cnu+8Oqc/V8iVzvaluiEMI53zKN/mS/I65+5IZxKOvKtwfcbDdjcMHyhfbuFWdDJkT
3IUd8JuXByDSJ6N82L5ReKHI2qvMroNZWEg66r+PpUX3Uy5mHyjA1eUGWLr4W6nTPFXVoExIPmdv
z1VQ3iJexN+0ewk5G5a/9cOjaMuE4rFx/kgqsGmFb6pdJzly1CaruUiieK7hcLhSao7t6FUtPk14
IVddai8am0jrUQLi43jnkJb66SPMBlG4XKRcuDEsEUH1LisJRgmmDL70g+gfygIVdU5koWPQ9ets
W9eW8BwsfSxg8CJdPVKuYDpJFjZ72ArAsBqZesuIOrwyts5iM1eezGOiIIAp1yuFEJAKAKLc50OD
Z/iby7hpg8LzKK/mVsFz+IKJp2o2ukkECy4N5Q0dpOa415uItcFZKHu4dU8bc+xSK+G0zKoR5Mei
iu9TSpSWnFwyqwUi4e4zJjwfOiKplu7JMEdaqeufJMUhxy5uVI4zb9uGMNgELQ5wE8GVNpSTy6Kf
awa42ttXhZC//Y5NXzpoc3ga9nRxrYwiHrQmfEVXGEGB4q9PB0ImyzTZuycGocAw0aNZCV3gq/bL
/P2sC6qM6+v6G7Tgul+Ksr25as+NifMb2SOifLMqx+ymVM3kcGaIf6UG6b1QZdBakRZjF+cbRbVp
HrhVLykipQ3KliBSjztpW7knZa2R31zUUl5RvXyQtGgKCRefVekg4KjJ4yq4I/bllcJrdlgbaskB
XjqF2jaCpP3fgDGw4eexOViI83OV3MPVtPlC1WU0Li5INfVwXC3BD4Jqp1kg9r08iuGcpXqzrYfy
yzAaor0PxPskEXUEBTFeZ4tkuXDScQSdDBK4eGwc7b3bUbnLxEdMYNTbuLBodKej1a4E4qjdRSWf
++o0DknxRbvxVy+CpHDHVDNW5Cphwa/cmlsBkhfnNtE3FSrvsOPQda51dWu8wo7ZKpTUqSyF78jI
0DoPHspTCBEJ3qZvCkOI2HpqiAlcs6FbXL0fdJuvQgqDQ9bfCQ5GayCnzNvqrDZ8Mi3ADI3YAQQ1
0m5VlaDVFw3I3PBfYx3o+xDeX8tvZ5H6MUUrpGQUoUtqsapDrmJK27odqMWvYaG5UxY74Egzm8ny
zm52MCreTwxVgn8w17rza2Xd/nPkAB0Q8GgQ5ZafhvITPEEq2gtYIntx3uzsmDU4r28dr4slbHer
I2cjRi2E36AuVoEI+/of6QAzwSkbtpu2vay96Mgb6ccUglnDzKTEhL59mzmcRcMZ96PdEaZ5kKhT
K+3PGwFh1QY5f9UGQ6gjei/5KoFB6FBur4/q8WAIbigGasvG+hObTm2q62Y65/6f6yFeE2UNSHd5
GGnY0nVKv8vexEogoKuv4MojM4IcTVg1xFbVI+LOJZj+yPlfQZRmmHx/zyVOkckqQD24AZzl1Opo
h9fzJMBqKUdf/mrFmjMIQCJy/KDclJoJCPfPepNGp/TI8guyL/p5t/bSPVONhZH25ujpbczqvmPC
KA3u0XFhRm02BcTw1SZXQnaZwOW55n8n86CKVdbzEOuObOgRTWOqaX/c939D9SsCO2AYzB0ezcmJ
VHeLh0LCav7vWFfcY2hpCNnf4LihG21eq6txMqVja4yihcHqq/ug4auF4wBhrMjAULRfHwl9co5E
Fdo9O+stpCtPzPF3Rq6M7wW56jZfWY6sBRcr9eEWEUbOiCR7ER6DENbPvmQga4Tu7s0WshVyDT3g
zV3De4voReCQ8m1GJfhaz1a9g6SjdtJhJsvpjbo5dCZ4StFgVQdthnPrEn21UvZp89s9XmN01qK5
6f73th57nzDFDzPtmDVjz3XVk0lPDkKir80X49bF7/vb0eUkx30RwHBWQvWKKsSTb87aruqcBn2d
beaPeCwT6nqa0kuZMqyZDvqiqoy6Hq1debd9ZUd6H9nSPiNnfK/5Xoc3bOsgAbTlVdQFrfgDdRPE
am5nYjAiI/rAL2yYW82RzLkGPjKw1XtPYHty25ZQ2Dg212AYnyCwiZlmo6EhjATjuqD4p2IgF08L
ELFy5DLdPJQAkXgsxEa0YGBl0HfBvlt5ty7jYD4wPsFaN4F+iue+8IPy5T88XLTS1ord8jfmIJam
eKzYwf1iXitpUuTQhF0Qu8lMThqhWA8yzHcIPjfkbUJ5vmUoYBlrPaSdOTNkNeUsHk60VPFV6uiC
3YdpOlrzXhN+QInS1v0ujkUaR3fuDMhKDpyYfJRoTNOug9BjGTVPyLrI4bwGz5LF0W5bDYXfIpgZ
R2qgGWZCEVbNTMmYW+m3V/aYFonmR5emJt69m4exlhQY6Ah6o4SwveDezo6EZ4PAA0U2L56hdwPA
O1lQqAdTZQ6X1TCBzHG9UlAYnYY9wDqVU4VZTaKkf61LDLDq/aLwLKK8337TXA15KhutdCMBvUZl
pQbm5PAyUmLN7ExxsYjB2HqQscYNwn8rhk8Ivkt5wEJF+YC3d50rpc3KMY0Zxg/QRwKwh3Zo3lpm
9WiPK5vAtdzhnan1Fs2rUr8cMVCo8yvqJEXTVRu2cqQBerlP1jZJWOExNwLrIPjA3PZb9X8GznDq
6idYFrNBIzMeCQFKfPsPjYfHfD+gA83Gq3fk6QIvxeVETm85//60jqYGUsbw9GUjAf48QHdMgH/c
QRYAo0opVq1G57mPnuQ2IZ/aFU6T/LW2dx8zwRSUHa9fAbELP1n2aNximlwrwTwJoIuYJxG87qOQ
LQAy1AcZpSLhZhbUIriUS1pP/gdR2OINsfS1Eo87VM9LXAXaWgqrz9x/k/3YKD25bVhKks3dgUcv
xdavyMun/hyDKoBn1AvMeP1ChQTL1WhOFjYXlnhh4YG4W2Dz8kMb/d7D0q5jFBiH+EewPZzCwSV8
gURkVB4ndXCqXVrdU784I9erQ+S/Xlu5TLOTJ6JXMvYQZCvDo4JGhgk2iHHDJmByJ4OdM58l7+FV
ioD/xk6S+eTbziIWrpWBMOh2kUxSICs0Za8YCbzltZwXSj9f1grJdGC0neVu9vy8383F9igNuenS
5Yrirn+zi0rYrcyEyQyX0tN47baXPoMzeQRe+/yCCwOWOT3ovgC4U1X2K8p01VdKnCFSG1gQtCwa
Vu/XtrOV5u42kDTTEVi9YQ+PO90dvNiZEu1nawd9NOky+gRwvvLKtIxokPcv02eBnrjTCQKpIusy
a+cGmFvxcYy+6IawPJixeWWKE4BYhITxDpGHnRQYWnDX1tz/J6g5slBKyp5ZTT2Xv6jvOJlyeEIr
xPBoPoDO9y+UKd+6tgVtJBs/X+kw/P2ca+RjNZ6Md2gVXHo378DXba+u44vt6XVh66R5eke9gHtV
k8okbXW2a4CE/r17to+ieVt/ovkARTiz3JSde58/sneBHlN5kJgooZXeCFYVEWPr5ERdqcXUiK3s
CC/4+YDoOxTthNxQBVLOKyhWZwS3ET8GwbGmW8pzsR5uyDPyk4xVIcmNibU6K0e/tWOe34aobuxV
ero5FX9yu5zqhtn3XAyf86fmhiK8nTi2SBFJkGOuJEJVNZZYZG//B+5QyXTIx6LBHiKOJfAYL8gZ
IjdRCvPCogjoTy45frAcN698qFbfJTY0X1xEJHFFD32JlZAokxld4XWK1ZNHCumkZgvNRNfgIxPV
J9ZfYc2Vtpa5KCp4NAZW4oI0IZ9mqqKqBzb6f/ykyIVD3/jTviQKRz/GCC9HUmxD0GFKNtfVDZz+
ERb5f8gG2NocsNebKjujq9JTVdR/AIROA73Xtm6iLFM21dbpS+jPJXEyab0k1i9Ez2m9IIdBwm5n
1DeuOOqZMJPcDNWyrPe9bkibeydnltT+Rmcey6d+1R8PEik4LUG2wkK8/1OYaqVLtoKhvHrHcfy6
TxjEg6QijMUV0gyoirhJyPa/nTTScBskkn6aiUSSGGsaudqEG+NnZzV8YTA4BCCoFemv80SOX9GQ
ohuGrMkOxf00KGFzmhYJE+JHStbSv0bW2iMZBSqrvFPzh7jYvMpC7ERXOG4nLji9EGes7HINwWlZ
VcsyprB7XLh5WhOBlduBDTBt/H6lkmEkeXhoYJAbFzpEaOibHUZJScsFyhG3xKOxneAgxRYBc+VU
vaxL/gkIqA5E+JgFSBCCyjv3UeeCdmM0TInnalRPMiAMLhbuMsUT/Hzjl58zTTsU6k+G2LDZg1mC
4R24wgRBAGcRh6DCJMofw8YMrOzIfdJJ2K+VoVFZ2329TbiJ/GUkLZxS+wx4hsvmgrI54PkPhwp2
w2W0BXnVy7c1w0IC2bcGffjwV2yI422+5jg3bZvMnyKlohtgm8/uMvls8SdQbvqVF8f7mJ85xVYh
zSPH7rsCvPZ4cfeXCMlvIax7eSjvlo6N6+UrySmoIeXl+m10MmQsr31BQszDlwQlubsYkzz3dAAa
wyOmhZ/8KMU2He8esvTIaoigBvcIz4eep2kYYZZNRFwBEunE90p//KApoTf8KwxpjwB5w0PZaMh4
efu00RSmLlcf/MnA648gStaEVLXhLBibEHgrOxWceiphBzWRnN44VpfOssOuG9B1trkJxRrXShop
3Ij1/Kw9G4sCQe8qNi0Cg3VxRxdpWVKWEPToFGTJz333vwyXNbYUBPvBaP34kJyNifmnFevTl3br
3J5Isml9EZhqB45tvctiAtSpusJ9yYaAC+XL7mEhHL25MrYoG1DCCnZPaybuJq8AFC2Bqqx4xBnw
nL9R6ofOYRGLLGQU0DfSLv+2kvfA9QQ7SFpp2+wMmj69FPegev4ZVPpFimOfn89JQvExyzgT2dA8
gdD7EJUoBOwWB2XyTtKZCNbVhVypF7AI0QaBMLGd2p8SKDGEiRyfYU2u79Y810PdyLBdkEMn7EoC
7zOn+dMUhJE7Qo8Cik4Sz70g3hd6hIinuDM7j9IOVl+br7n9q8jMJeiLm++dYxLSCh08/iE5ZCgu
g//fDmMYr/pa3n+IvyGyw4PgjwqRmwHAp0R0DOUOKrn1jyP51AjBhrFAkSTbhWQ1So8hmbrLdneK
bO2nPkIiIAMOeF4kMCylB7UQGNCQ+zFDfjmXG6ghNW4tWvo7FX4CzBDaJvuWQge2QfkotCVKs6fy
qRXa2Olvp2Yn5gStyM6SThlydj11yHJ0itQ3/yOJyPyadRF3ApIasgcwnj66stB81H23B1J0vUqt
pAilMWDnogAPxrDWb+LTUbijgFSV/oto4PLIO6/+55wT7YOPj85A3VEEvZ17uAgE6MtXtvcfmBGi
59Bgr0QCY/jzC0ZF4/Jnrfh11e7RcJpT9vsKq0qskEzjTI65XUqc/oLD3CNRmkxYMLCmSBQ+CYws
qefPtQ8cDd5FXTRfH0s6iV3Prgkgt9Lz7OrgFT6c5OKO4iuLYtGink+jWj+LnVTdK7EuQobK/yic
50oertypcGZeWi51wWRwTJnWLNpPPQmVL9+JdEAGMJJv78oaN9sxfHXeDR9nJoqqaHos1FVkH/Hz
OgmLwkdJdrqE9xceT2mkfYFIrNvAamw7brcN3pSZzgGGdDy2wGIMpbyfz4CaPANEFTICQRk8RDBU
uk+AY5V8fm/gNZ2cKWrCCHK5bGkhvB8XjnZeLJYegN8VTTWQ5cl6jUMUyocJr0xf18J+zlFs4XUN
ADs7rznlKlTuSIX8zxCdXvbOYw4G1MGJBSgIrFt9LUbJINqKZPyLh08x92+Zi6PYcfbgREiGWCpP
O1NB8EuTDmk/1xi82rFWrzKwqQJHdGxxlmWBwtORcWcIOJvzZzNwK1ThDYciFgtowi0QMhlFsqql
NpQrzKq0UCz9lCiP0jOzep4iLiKR5ATb+2l/cNx/N4UU9G1+oHXlUFA3+8SqVvbNKn87rTlUk5T/
VkPcdLU7dnzw3FFPZnEYnmKtum4H+Vpl8S3x5Tie9lS+MY3IfR3TKDcBxz13I5OP/e21H2TIIQEj
6rtIwhpDSD0qM3tzmDwmHhgd6B2lvHY9kXo/K37CrHhId5k1NS3ogxahyWjusxz8+4GkvkNotvGq
KDnCMjZX3oDkDssJQhYMbH4Q7+yDhowLiwGFVR1NWWosEF7wx7wQLcG3yY/Q0/Tq6r30H1s5lSkP
iNCZoC5ef4DqXYhipHNWAm5jHV2xwOPGI1ytrx6PsgaLKRpZyNB5zcBicb8ATO/ISgI/02CNTcKc
9fpHH7DRmlCCEN8hu1mYGmDDg1sfGhXC0h2Zms0SGVXLceOgkRvIkjpSIgO1SAFt0+jgBjldLrIN
D6KwT7lngFE1LImg3IRLWvOoEZ/JPMnmUretWjjOSeUj3XsEa6W5WieQ/Op85kY4Jj8RHBnvaWBm
64mkD48jM8bPL4azSgB3olDL1vc2meRXvy/vBYZNyzU43kKUVmisNlqLjcqF8+cIb5Fr5Hm+nxB9
uMlpmeXAlv93SEiASUoFrh2PYGo9jXfl9YU/t4PhCP92qbAJaJVIa0PkdRlh2LExAJUmVvvW5Ozy
yflkqZlbVF9h2pmPAEijf/kzPeul3UDx+DyZ65tk481FQzdzL5eIxBqVF+eHZM87qMumXXuKz9Xr
MXkFI9k5hX3DwHKnkjG71VbCl1Eh4M1nj3vAoCmzLerEvKAVSzjH23uMldFVx5lDuWctAVbPZth9
AusDx8KRJtzRKwoADbh6PtSbJcCbXBVq8y0t5DjpH5gOlSmT32M9ZWWzZfTvW2uDJRtIL0pP3Y9W
L1eXWrMr/8rJnjCEVhTUXsja25/356kvY5Uz0H/BGrnqSQyVi3t0mXJsVJFZpaXIR/A6QUxrXy5V
MRmwERR1mOG52unDNbt8Ch3zSaNT7gEDu/5bgOnvrKv8vY+Tubgt2va967a+WaNzZn1UOGHKZsj5
H7N53Pw41vJU9Z+iQULMpjQZGtGDjxeN9FYmkVI1vzRROw3EAfo/uV6u4PxJmWPrs8AE+XY4/apY
aHfYhakcYMbtgeMM3w4zTYvl08nPgQl/k5jmb8xc4vMr3zA0JiL3+eTP/nIU+YRmPdx9hhbEL9uE
P25uTZRHnzzoc5IplUruM1VzZqEYu2wDV7jUS5cCxs1khFRJm9sQgyXYS+Cd6mHenJO/NmBBFE0S
wJToxIQmUB7a/8Jxsj8BesqOSj66Szz7DTCNCLx4oy21dwFqd60I1WQxF/G4l9GaRq3XVg4In118
FPY0iI2uOd88Dekk3T2bjp0gqUqD+frRzxYInQyyxG4GhdtFjq7gEoY3DWkKk4ShIDSg/b131YnA
zYTreH8akAYYsu9T2AiRjWbk02A/EXuLnkbkjC92D2P7j+a74YtexFnjsUF/rc+qDisReJNs+WWl
85EfsKM8o9m0oWfJl9Z3zN3GRA/4tLtlFGvp8YQ7T6PXiwqCl3RGLQWyvRt1Rnr4V9jFIYJ2TG71
O23dDEoB8RtoiM4MJkiPi3BtP3U6urx9kTU/lIjD1sLl27vj5MjdPiYdcOjV3nIRgZrJ40oTMYUh
KkasApouddBZc34Lwr/lRI0E0Vd10mT9PdjJu/9YtZe9+yyhSWeSOCXarAbLsRwWi6Mso9XYK1+O
E8LH4n6H3IFp98NZylEuBW8AliApRFeU/2wSOR7khTonsbrJOa4ciZYoD/HfEkruKDOb0YYzoRee
OezlzK8ouXqJ/YtMhWRTOZWFxs+Ft2NLhLPs/39zsyRsC/py/FmVDjV+itlequD3pdaK07654PWp
ae/0M+YrkoB9bu2c7fGievgWDF6D69y2bcsawYRgHiDR/I0sufWQqotrjrbCaSPmglX7JjiA+lXF
CX6T0pMgu3LZSuV5s+hR92pTU6e0ygRNojph/NKofPUV75EhrlUj7n3nslel2dooL6bqN/Bqsa2D
Vma2XfWIh2f0R6ovLqYz/fTNQs9ufCUzv7bOUBtRLHpoY8LlFzU8UA24cSadiRkuGEF7fTXFZgTZ
pkfMWhfBhwfElyipJtRbytBvQqvXjMnqt/sKrhC6mkKUYyDbHGxC6WZ5b9qiIdiAuZDrpKC60KXP
VAdC9Pn/0oRO84wbkajtErhToRwEH5yKW79sOQvkCrht2mBBs8PeE/7bpFo64NQ6DvrEgVQQ10Xq
pRQnby22G41JiJGosgLdV383Tf6iuiHcEbSBIpvdJS9H05H655cYJnGvlcYdiQOyLWu9hpcDGMR4
8XtXGLFRVWZhYl7K9pqyiJVl+KFneZ3XAq4RH9elSjV8rHTAU48U++a47VHjxenOvqp6ydDfRTWe
Q43FE8Jbg7dwSvSp4nLHxIA5Td02ADb5cRAknR4+6CvT9uii5XrOtFMdGEL09kq4cB+XJlf3M4p9
F3y5ADPCJE7k56ZxEyyyKmI9krgjgaBSDcXkr91B1BwQXczlB6xEtwo+Pwcta7pF3ut3P5UUphu+
tT7YgD9kzww2jrdEEKUGOZ1ZXRwThT7eQMPgzAEUwc/fiugh5ukst/C54dh+no7Odkz9wE55tf7a
ig/UjVQxnKUVzmNqtQIkkkJGb9vO1t4NcLUOMwfUTChkXiHZadU6cZ1NdctM5SESzhUIZOtBj/nc
iEhe1A5rGnpZquC3r3feSjwW5J2P/JZ/rR2ctM3ZjKw5wSRoGC4WfxJAcL9ZCaovVT4/lLRCl8/8
3XHMHgkzU2E53NMexfBqs2jGguN8V2XUsENnqTFvxqBpp8QGESUyJGCgjex/3GszLJKHSbPCITrs
kdVwSw3bJxlTWGTXeC9dygZhqeP+uYdyBWnKKAd0e8bBVHIXuYax+c24JAYtViAZSvRHqepwwzsZ
iEPMWvGKtKPq7EPtluPSWhcL+64XrlrVCAuI6agy7xVi/1jWWiYBAFFKq1+zHfUaOyHBLnMtocTO
iatUEb+5vNGPuvUcCwviX4jKWyDoMs/kL5ZrlHWXtJq9uaMk2PvKageDu66EQUaNpZj9HJ+gl0Vg
sI5LuGU4l5kP9+7ONwol9JW+xu8xZeEjbLa41k2/qK3U142asUq3ZUOZBZZpjAk/W3dEdoxLEPYn
JR17HXQYUaqA7Mf0KvcGlQzB0dV5v8+2dMSj8NxzpBeWCdzMVUl5zs5hH7pm0Enjw7oZgaUc3v0r
3X7d8nSL7oe7j8dYn+1Fjb5cKDbN7nxLa/C9BVatwsCRrEVEsGJ4w+X+8g7WqIq4Wv8R9w3XzEGy
YAUXYULffv9p2ZfKMCiwASfxxfyJDszP3VSyirkVkOD4eII/LWhVgSJcyZCWTTKaMiXUczfaXoOe
RnAdNcYR+SVKf9+HT046zJmcmV4I3QXmF9P5PZwD9aE4doP4/boDM7WGxBR47tr8KxnDwFHN6rV6
bXRx4aYGgFojsd/PHsNGLuckV+mQZzJzCFx7zSGpNd/sswFc4fvuc3Z/9x9Xfhj/qiA+6wRwEpI3
4r+ugFUVKnL0GhIVwyams6HeAiAqnkk/1PTyBF16We1pXjwcVy2j8bG1hYx8A+TjQcFAov/EVYK2
CdLvt8idKIDb+xuDOCSXPAEao8BFGceps0vYNnrCHTAAHD0/6x1RX17wHVoCAJ9IrBMZ1yB/H01j
X+oAPfWRiLuzUQ/CNdRiG96WJaIaMs1kdrEU/4jkzCeFr2aiFrOe+FvfET7aP/AiBN7Z49GyzJU1
kHNkpw7/B5BdRBGqvI1JCGXYTP5p8nazAi4q32Q/REes2bB4w+wi95v+KP7gir/AiZvtmPCffkF4
U5SDuhAmNA0V0L0se0Tqqjx7ZV/SXlOSOjHZQCeNfKIQaDGe2/zpalY4ezWhd2dMXO7YjwjjwbzC
39ZlCy0toyCfb3QLX1r4QlOXZ1znLfCCHqPRkVk6ytEx3UfZDfn3IaeRd3WawYy4Kb/NA435Ae1V
IuYndJ+kVKeA7s0TivcHGfa2UFxPWIMA4lZ3b8BjGPK09oY35lo/RkUmGf/I87VJb4B6Ti9YVgLB
xQuVBQRmXdBf3EVJrNPs1ojxKV+AZXuIrF1ng3gTaWYxg7Z7EwrZQn8jhPvQxeJhN/5R+BOjBF6g
iVvHPZoiiEjmMvafSkTit+Jz0MBNX06eWALhANQSuM+FA5BR4I0q/Uual+HhIFH+YUdP4SVOIoH7
MUl4NPlwQ1VZ2jxy2D+xGxRT6GrgP4PTIet9F+d4ukJxyh3Hei8paj6T4+Ftjm6fbEtmeSjZGYcF
uFr5q2gKIPHyNbcUcMB79r6V61mxQkry+b5T6s+PajbDS5sLssD8nOYzEkCZjxc/DChBXoMmmXg2
fbGvy9yqRGRAVcOKB3DgScRI3f+Z0Wce8giGRarNlIBHgmdZkNsJcZcXYqBN/ih2gAqUGxi/YL/x
ZuZtY/2FOm753tVaOSRn+oVgcyPdv3Bt8CqK/vbGRH4xA+nJy8UuXYn1vPMD/7Vsns15SG69CMnC
Zhdtw93/WUFfoX3QbEoxFExyX++Ved9NK1MVIr0Gs5tq5qPuCZdu9/9mGvPLfo4nNnpMogKQYb0R
jRZcFMxPYXfc+7i8iP4hu97se48Crt+KkQo59zE9C5K+pxUT9f/BSNEVgWfc9CFEwMfrPMo9isJO
HtF+yJPrnESyLu7CyaV0ElIWl4A8voZK9DUM/a7ZEYwzMeqZ7oO9Q4lnzcRy05TFbCm/LIh+JnvU
dU67DJpCz6UrH6+Z1C+Xaayh/iwo5YDElrYrHNBGpj450jff7ipXhGYuKtJ0ZWlDM3L1XHTH9IkX
EbLoo4z5+W4MR7ZtmXk84n6QwMWgeZGv5wM4BqF6WTFTwggIblF4RKl0g94aGx3Jshnj4HilM3dh
35x5mNjsTz9PR9lXjpER1Auopmnw3xxwX4ATj4c3cxs6/GYbe1BjtKmlPF/db4+NxO2eXDkQG9Cx
No/8xeMSSLfDa++1juXcBwDp4SnaAoSYQ63c5RI9duj62dK2c/4ucDfdikXjWHQkLQPYvI6FivmN
IRYyk+Zv3L8brtQUncUPekwnX64kugvKOwSa6jBPOjs7CUgt4Squj+4zTUAZvFNG9xXOE0ojWqPH
Qp2IORz0W/AegQKdJF5KU9sIpZJIJePSmBcxVNFvB7+EuiXoq6mhRJOKv4UgeHhjWxX0WlOuXYtY
jHHFMdowpD41YpGYUyljSy32dAXU9vp2RLwjdnov1r4TRs6pBmUXqEZhL2Eh+k9vkLEGPHKajybx
uiQndnFGUNLt8Hhe6aNSd5BTJOhRYA7Mrmz1rth5894QnUh0nN4gtfGYxhGz/j7w7xgmCRpAh8uu
mmG9wrrLzyYLv3k0B2pEt2uopNkwhj2KZgzLmksB7w/iOqx08vbbAWezGfqK3atkqfhaKqx3a600
SoJXbRWMxcq69SEUdNU4fwLh2Qt9UXC0P7AyUA127JoHc8l4mZppPuslw/fvhuoUqxY4qo6E5Eqd
fT5C0GL/2vpjiIXMuRP6yURwmIC9GJZFFQk7sI04KFrU7xnxjhNhIM89ATQhLsReD3ApIIe56oHl
AZBgB/LKhlcapWGrW/srvxs3niwYAypipP8s+/9hbv1k7wqjz9dFvvuCLrtmh7imiobcJgtQcRTp
qiaWtmxziVqk5dVfNAHnzOBQaXTdRJH/oACLYAhlKwbiucSLpnYzyszC7MagwkdmTM6+jw3a5q1n
A/ncACnqeLVCl+vlwE0DCdzHjcwW+0UeuQyaTeyIjm9S9d+p7W7I29OLpdGHQMk5fm/LYMq6P4JJ
35VTXCvD6Z7XVfjWcMCMysEJhxJgXr4xlsd1IaOSvxMQ9/PtvmGtnhxd1zd25A/lPf3A3GmqtYec
6y8sBypMgFOeEPGI4ExmWCOY8AVlz2PUJzAa07XuAOa5ypJhwvfl74t+G1m9fqhb2RV8s4IkOCL5
agQGqEOk9KwgjW1gzaHkhrXf9gL53KUMDN0iG0+z+WFYHEWljK/33EU9D28yFat89oDdOmAfgpvI
xHU0WjBomyYsLxctgCn2eb52Yy7zHnRT6WZIvwnJwnUFwx0dW/gmhKMsi/GoCPsvlSFne264F7fS
eXsZTWyviV/T1N6AjqeVe6pHkl8nTBF7rLfnQyy9sir22yJ8jJ8dK5VGdnCgSVvKSfg11nuB8jnF
zvTrqYZltRWwAdpzMACsG277hJEJ7Cts09BTkUd686sO59W6aiiU2RLVSXXLeoNXTLNchFKfYQkt
YQmjYxrc0Bc4M6z35efxQjXkLt2q5F+YQB10pIc7OIFRodvQUCpwbGyLVZ/AgDo+E9shjNgGGgK3
tPHnBY76zGCNOk3oENtXi9jHUoUywQrtFOTQ+cfRDB3Wy5LjrF6Kx2RT23yQJ0QA+9jTijFs8XWE
FaS/WKtqjbszRJDFF7K/eWhJ4sJyNUPJ70rzS/AP4tbwrEXAmhSlgIcmme64KkqhgBE/vhWey39J
6iVVmfQGcDewWfzDg7swzTbPkpd99jfRxgKDGX7tQ0DybzJojUk6msPMz4smPf/owApTamyPeVRY
H1dCd6+JZRnSkPqqUofOXuFKrR+QtH/xZoIVn11YPDwrYSHmhHRdbghZb1x1wBXmgAFCHQi4/nm9
ugtNEzZfnReBqxHwIFUXjPHRO1lzULR4YES3cPgv8wiIe+L0yLmks9n4j1FmJ89EkTxAJr8PpWVx
ou5k7CLuleKw/d1leMoSLkpR/VdrCld8G9d3DNd1auCIf/K2F+4KIc6UgGy45WJ0u2ZXj2xmZss1
fpZ2UP4AMzuHm4QBzD5Njsk4oqhj1kh43+eK7ldLBs+yXd2vD4acIUL+aEe+pP/6Ju8gGGMAnP73
rfblNw5LEjkIKPF3DoOl2mfCg7JMBZMHk9mwqYZoITzo+6llJvbkZcF7mvI0GfgqU0nAqv+AMgpO
7c9DpBi5szj4dTkG2GMUTstGEjQKsJiN09LMqWCrdO6BFgQIUPJBWEHn57dCxwoMn8IyRwxueH9n
wgyYjtW6RAduSekXiPxhvwqPflVbX8hmS61as3SfCHYqy43KBFrIFtXfKay5IFDngM/M7e6Efdpv
I0dW9Etl0NW9sqErNBCq7yFkY0cUj8N2iFL6fFgbkKPd/UZJhn7pzXcu1codIPb+wnv5RnFM24R/
C/qTwGMUsjuOcNf7PeUFc7VKeyOrnLQoWy6vRgmfAPiRqAeZmtmnYCrZN0Dt8rQdqog1hCiy4F9w
XGfhQgETSlCyz+YWZ2QJ3hcMDW9yVFYxQp+uyvM9yGPt7UZAVWiarNn61RU3aj0qA1zmG+URlu0L
H4ZgSqSnosv2040KwZoxsKXxToaaX+qJHd47oso+qiOC4Xv2Z0iuWs8iEEr799mvwxxiOTgkrnww
e0LkcPYf7nhH1iXtlHoFJ71dLb7xwry/GsIkgXGg0+u0PGVCJJlFxzdwzuJd/mFD6nYi4manP1g9
sdQ/0LdjUYiSU/eWMGAUwql4Y8duZm5WUAaNqxDwBASt5a4U1TjE+KQHwI9FdpYRGeRbPK/Ifpjs
WxzyZ/0VAC9otjRhUx+PpcBlY+mcu+2fPf9tmJichwgkWKml91meps2IvRgBO9bJmO+cxQGVTjfr
GL2nnzO3zM/mQiL7bJ3yPaWpqvEiCqNoc4XeLBh9oPChY5jBpJglcszilYJSnpn3FjpQya9PuNIc
4081jVsJ6yII1fCCUI2aaQpc5K5rFvta17vTkSr0/59vAzgr4IcJFcM/Wxm0M2oNWlbYh6lCIZfU
zrQveiApo7Gm6+dQj7C1xfltJKcbXA1FHhb3zUgG62Ozt7kiU9eusntXfryyDPqk+8R5VhgQbT9E
2L1pKdYYPAPZBxNHvtiQWEpeX0h54VhoyEgoXQkLOMSRR8UVFAt7pydY58lMz0GMZI//uuO0p+Ge
ZUvJEtYtwE/KI3dPTikQfDLcrZu2+tfpOuassqO2eGFAhpZry8jZooJ4PccMmS1gpFz4AyIF7JIb
ch3mdjmO1vcCdXwXcjj+KDh5mjcFIQDlYUwh+UWLYmRHORqaDJ1MWjyVJae3HGaTdKN4CzFH5pzK
tcYbFJHeM6PuVlyBFOBGAfIge3FEKlqqtDAkJ8PIy1QbA32yS81979hUN2kp+LuSki1dCX8VYCWH
laK/BsjmnviT1N8JMRFJWBF2L/3eSYUJBJFTmHARfW8+BD0elyxAdHqPFRXzhOQ7fzRP8vU+MYOg
Cfc14r/Wp8vTWocozm7yVDxYdzr4C11dorw+DWKn87XbWfhBXLqkPSA9q7NQJWRs9CZM501zJh0f
aC1IMJQs5skt1WSeeCtZxOaWe1tYZ4Or4wdtbbs//4PfDXqQXnersImp/ZBNQcdZGIxhZtO5gzOm
IhNHfTf9uMfr/sC1I/vK5AqxPbHRQdD95bHcAlclKpF8V9TLMEotPTncnf3viz+41M0XtOZ4ElbI
9cTXplnw+I27toZ//yH6AyEJmUe1gheU4NaN4xEhzJIEXvI/R/AQ44ZW3lLBLlBgHI0CGNi/dTqD
S+35+meVEqZxeLLXnylriWQVIUMmWkCQAJj5r65LeFEqOODpeFao8gLcVNveOR5ZKRFur6hJGvfj
mnOBeLcmttgh+dawklXJJ2SBCgsKreMJa+/9wayZE80KNFadkJbn3Sgra0nusQW6STeH27fkY5C0
dTgSo8PaTQiiHDnnTKLXq285MAawatL0nUsQULo9Rwioaj8vqRiVxq9DfIxTLP+2bfKLMNgW0h2D
2koDcHsw2TjluxS59RFWiiLsLzWWLvRHPN951Nk2lhuDB0NoW2aXcCKIOIiEPX1sQdbrLps0VNMC
A6hc/b4bJpI98Gq/39AptrLPOAXTppGPx6f2122ucAy2AJTPwbmsW0hNLc0NR2KSwroLn7lb0wUi
E8nX2t/ORlLtn/zoUt96Oy0jTWoHD/SYMBFzkYB5rP8TNpGJbqs6fh8VNwdDgHraje+IUoi1iS99
AMEzp50AzVlpAK/kWSGASnRbK+cyfGRHZDG31CA5bwKYI0X5nmWhRh6vffHf4bQqz4OXy9eWtKoG
7LkMQOPJ8lAsBlZQXmzTa25G4s3el31WdQ4mY3fx3ob30wVBiiOo+af+94biM4LvSxEXOY3Jw7rK
86IRpms4tTSCjl38xj504uC0W6/WKrNF6AbZQMNbs2uYAEQsGiEN+0ihE7OJ2aP9QRWzcFrtCfab
oNyTyEe81mda3iJ9SuPRqkJbrvkSLrFp2ksqQ6mjoQI2OjgozSsyuFEcZM6R0Z2cmZXLHBw10cIw
RWQsA2dg5q6kEMEz/1hUc5wTNxQyfCSqwwj5IiNQhVv4UpQX+CqMrz1NDl9zhO80I7EhRhtmHAlO
TcdWDH232LGz5UZAfUTImNSFiZdtqotgOICzi0JqZIA7G7ubnfCCRCb/nAkF81Z+1MfnEsZeFDbs
WjS3Ve8/bHwGN0uHTATkJEzLAZYeeRbP4ry/KGOerQ+nHEXKrQzF/Ze3UNFxmYyL7beHrqxb5FQ1
t8hwl82NSFuTUAXs2Ps0Ea7o6rD7UpOcLWuxf//9+jeHF0zCc72E9D1MtLiAon9kgRGT0WwIVrPy
3suQu4POkzNppYA5DlYml/C3e2LIB3Y3WWgn49fZkvHWg1/56w+/QgI6jJqYyZENotoOa75tbrgR
8cesJgbv11nG7f0Dmfzqf1xL29/f0IXqH3AoUnwl6xyqkoj/Ms3xk8U8hV3Q1BZ5DJ5NlDMa/UnZ
OTtqAMGlRyLh8XkPKpnR2H7/t+mjnA8eWtr7jIGYIdnC1oUy+GuVHVcH10UczMC08XUAglw/OSfY
ZRmsBya6Bg+pcGfhBCBpIloZoa54N7sjwteCZKqAexg212BQriigs5JUIUWAGdXX5zySdd3eAaRH
XXFhMEdT1cACeOWwkoDySzeGsuy2axzKaNXOqMp/AhjNEqRVhnNqcN6vOdAiijaqhdyxZA/ETC8l
TfjZ66xnPARsuirmWlyD2ERfpyVAsd8Bp/j/+W3yA8A/SY3dxkLmOEiRDFEkpAcsOfpKm2HyStdR
NVki/piMLRo6VF0ew6VKhKnm2DANrOF4tiVuQepHAwwmyu9ZUEjkP9F+xlEMOdG9lSMrQ1Rixlvb
+ZqtfA2VIq0KLtCTyPfGTD0X83LOuIl4enJNkiCLRcrdxWuYed4l8+wv1SogNbLasItzyluc0wdo
6k1poZk/UNLYqUHC2yb2NGsRftPtlrYC3r+fZNLdp3wbPPwvDWp/QFzFHBrzujC3+pHqjNwBNwOn
Df3v84Tl7raZl7nPS8x/RNZF/0LHiKpSufQe9OcrrVsAHUi2pgpilzUL+0RCGFPihNsv0mjYS0Xg
FAInXylQWAIgOAPPlk8YxNOBPXKCNPffDtprxRUsx9S8BGHDcfEBMH8nlS5/rJ35HvKWe7WKqixF
zebVr172zr7pQC9lNdahWPjDN+E1DzcYf8DzRxe3/I4CcO6iqaEwRleSfzdItf26IzzgJG+ymYnu
mH0/1glNC8J0zizTBXgooR+KX9H+iQFYnLCop0562FzlHdg0RBLL+8oGc/yKiuOLHxDIpedgxYRo
qU8MUsmgXkYjDrEzUBh5/SSSQ6dPL5OiWX/h74o2T7iV/1qb6u3QxZ+78wObOR5X9Zvm+RBBPw0z
xs3UlTgmh1V1jNEAREpJpTKHJ7adIzu2O/ryyESyDutCGCxLkd1te9lxw+qH5DN0fVjMkf1Nl6gY
++G7d0OnI4fvpgW4oK7zMlqinLRqOsJw3RLyHjWbrIZc+gkrx3GCmosdf5JEh5iTnih+imT+DlUi
vs3pGzkHG9yLBAOMc9z25XNg5PyKbCo75OF/nXIZeOmrA9TUAkGgZ8woPVYxhw87YUY/ePSnPp6p
UOR54RSsWTi3n9Ru9Fkc3oxh2VZsYY5F9B9o/bDEFrdDOW4yY6chjaD+4dehKazGSvvMYU4ipZuh
YIu9kzGrFmpxazYW306nuODqlL4Npg9U1P1OPmnPtKWAMF1KmOj9H/Q/ZWO860YjenXKrKFGgI7M
THyLwqc7tTb8wrMGGTbrSj+6L4eO3lVszfPYs+AJ3PAlKemSzgh2sQsM3b2feCRA7HemeTAYuT75
JFRAJZ1aAbATxvFS+tqIkgPCLjZBDzsIx55gHRV1CiIMhrQ23U+jh9YdekLzoSyW1BjyYQlij5do
L0vxG9jN1ir/qUTLILqtWdP8VfX/rzBR8SJMZLLnNOdP4xdYZf0H2np+bTohP8PKZbMO2A6ok+Tq
s439AW6tLtKwjQqZhLrgVjqD4NpB/9DxclQ1IEzHk20OjIhK2oYhSyj92L43XFgEaVI5sfZH9pKT
WwORMs7ZBVsT0M/TWrYUlHy5/BcQWtW/636Ufm1oDotjM/PF42vuVCKkydaetC+s8nTgRGLwL0eK
vvqD94jVzBMJ4S9mW0dKtcJyXlZh8tPI69KwgZ88V/NpmD0AHpxnqLCZ7mktAx/jt8P0KH+QMx9J
nZdu2l/PuPp5rIRCjn1oq8JQc8KXjcApT9zsKZ1zy7lNPrKx6aBk/c9xjVV9xJojrqTa6qrk7i/q
Y1tD9aDPGpEjTn1Edm3iBk+2bJMSewCTxS0QNBGTpfm8rBZ6b9ekLLrT7ssgXH3Ruo94094ntmXZ
P2yfg2nquZisk0Kf2K8IA04BOgox1C2RP8wwXow7t2OYa4Q1FtpSnAQQ5phe5ubMTll2PiLQkIqe
FnNHn1PLUlnLh9+4DJxEWUvEOUxlxm/58lbWil3MwI0xa6sb3BTE7r6CHO4HX8Eu3ZrtWcfM9R2w
kxnDL8DFy5e91S9xxDK/rWTbAc4MLPGwStHI6KV0yEO4Abj3+JK6Hp5sKi8oDBksdxYHR+eroW2j
J/BKJG3mX7eYCX6YqeRVmpLTmP1DhPLevPRI1vwbyFdQMWtAqkvzE7JQtbc03A7WgHFQ2iUD9h4c
B3liNOx+i9GK5cFKr0g4TaiIk9m2ZCk61wTynNjyln7NjjhQ7atN5ukNOclR3/wXe/RklfUm/KeN
TNct+Dz6l7e4Q2OMWMJWrCwRdfZBHgDpSG3JSpko67V/M2giDjtAPknbZs1wDZPSuC6B6tngc/Z/
6Ohen0kN8simasa4IFEcRGmgJbvQ0HncT4I3g9mZBCtJSOrj5Q9vwry86YydaaG3Lw3A3NJa8wjI
sL8IUQ41rCeU2lhMTno2FlIbe/tR3OmcLKIn2UjPpuOCWzrboEIaurIoaYri6i5naGD67MtB3nIo
0RLWONq40a5rxVo9CldzxoSswdt31ev68CRtjFmwinFOCBhi5wc22UNcy2CeJECBNUTV3cXrfvTc
Afff/ac7H8Kcv6WGQEsWJnQGbRh/25wp3VwDQG2xoN84l6uYa1LO76gBkTce2Sc/zD3s0c8FhlGk
IkvPp+umtVi2MP+a65SZrRlyUm6CVS43TjXxthHCr/zesxh7KZlR7EhY0bRQ7mA386UeDzWv5Uu1
EZvfphNhiJU8kvrFPH7sASvuEfxxP/J1LZRERLQk5QgmHC+F/XgiGv4SCrmuv3qpQfD/5sK/SOv8
BYde4HfCYvMFmEe6bEUEbqkcEAnkHeSf/7zfFzdZ8u45fWzpVou3Ua8NAspAQUyO0VJrkPV9akrN
Yi62No0gFNuowL/D+BRUC7ambXGspbs7AuNxCp6wAUKRQEsFb7QQq5Adv41YlkgNWhSGCG1DaFLP
jq6Q7KvoZTRFWpDFNw//7Js5CemsTJLIhjjQttj5cnFThhF11dSFPAcdKP6eFKvzvzpGAcW9Wvgi
zQ9sU8XoSHO+mgnoB4ZRYrU6emjhwExpZpyneaoHdIxgKoy6hYh4n/sKvDs7/aky20lPW0JGrPUK
Q8n6T2FTNXZYS59vWh8Z/RysRKneoVUR4rfE92jy9TpCSO6lrBNImbyaoC0dztN21I/hMQNZyDAb
IF1l5/fqUirBkUsIHFb4MWOBESnfaMCuSXb2/jsGp0u/8RsuwXFbhzsNQCguZCJVb2VwNpioKnnH
ia5uPy9qkx1Ddxpxqkb1yDNhv361i0I2zNxZ+yNArN2lWAaKs/95e46gB76l47+oU74XJrAaqgII
8NdrFGftIxeMQDUhQxrwg94Nhm+MkTdERvB1WBXViKWsYDwomH/kiY+Xpy67dkUYbWRYTx9E5Y+o
+UEnz+Xvsrhpqg22y9FfW3GJxnwGH0bmen9+0DMB10Wf3B7DZARJKPLMSwDtCcbyblIUrM8DOi+t
3VJH4j/AUuVGfCKtOPsIt8U4/aWjEDrUGgk56vZHOg6yEeVSlEDQ1q9LIl3QZZokvl60CxL4ibi9
5zH+5DjqqyKLWSNpUbJ+oi7J1yThOAikPuqvN3qy4bCiCrW02dZgZO3hAaRksCD/r7HKXqJtMCI8
ukdewxnYmOI3n3x9/smwuY6mjJGmw9RIEKnkeThMzFwtreQwV/MWaGNl93ZSURtvocZhAyMVOUBs
MVfVTvj4SY4zfOPOYkaWJ+lZCO4lJe+ntVaxNN8BKSQGyrP/85ElnitsM91al+EIMHxviOwK4wpr
5j5x9VYu69lAshENIDZfTahIoU/5ksYq3a8EK1k9H4ETCQxANHjKDQL83Rs4iho896FMxsXvckQ1
omW7zO/3RF4Uw83hwS3t6I27NJ6Vomi2vNc9xeC0Ya6hGXwvgJcERGhvENBWdHguMPIt3U9qjGmZ
ALol8BtmUL0t5DQSLwGCB5fkBu9fRF5PwNwQolfvbPg4RVPqpB+Mzk7TdQt5gtVCHxEL1V0zpECV
paO+TBgIU2hs8oXae2sdkjKQEdkUhqLET+UJFPJOFNrttzRdhvdnHV1MkBMrzfM4dA8UCOJWLBWi
C906Gj9Ma0gcZTzp0PVuzG3OM+GTEB6RVmmsY7ONAh5WwVyYBHYh0Hwjuj5xmD5mK6z/1yDKMWDh
bLnqqRKU1pAy7cZZl9ob0Y4TMbry1KdMpdYpaNJLVGep4vCBuSYboTg12sOzlXEMikdca5hRLXzP
o+rlp17lLf1JJF9oexxz3Ef9nikZ9VScvr5x6W98+dP1YMwnA7QM6bA0cigUlxpXs8IK5VEBT1eD
Jvg+6LGzy/OWbT31W/VrsH2CBWO+3CLvc+UymPBBQ114/HgqRet9DuhHlpRZ8Dn43Nn12/MiUfk3
sYU47su2d1hD5eOh5EkNsi5wYlonCexUUlqCrEHwQCNtPqaHhwWDvmvIJzTttiG+ocNOcx/wk6QC
zF1czotrIBm3Zrd2AzH5KJnAFdaNjtLOKgPqHHIqY9gNbDlWVz1pRrYKumOlMUhjAzI/izxQwc3X
aKJKkCCiXwO0OfPcXPSNRofOLAKmy9djI6Dkm8PbfULp/TLoN9V561Ts0IEbS3jLNqLFI060JKy7
k8/RuevaOo9qWR5fc4m0Mj2uCHYxQ0tYlU5WiFO0CV7agFwMMpnwZKaMflLIRJRAYCd+Qd/5TzTY
6sgjrLx93M0NC+8/yJzBnKNxUCX/rCNcLzeiUF+pCAjavBCBt8sCP08NZ8YsX/DtR+wXshZ13NC+
qae5ee7NgFXw0NsDF8B3lYltBcxbP2RKIdQD1ka6qH2cj8eqA4mBg16MGQaiiugPCgBJU73hZbxw
+tLxMI9fB4zqi6Xz5G9S4nvlD8XOq0aCcO0mZjMi6X0M2NPnS/+zw9YZAOHGmLhEf+Dc3AUDB9Uo
4HRKf7hB8JM0qPiOLSaiXAeUV/EjiPcNTH8qtL+ftyAnlwT0j6xMuxFaxJhcGz4SAX8U8e58T2pR
pHGhHUABeRNQSohMjkX66mOUwClIyqrcHSd62U70K4aM1pbdBAM0dvYQP02uIUvhQseLHc0xQ7so
HOE8gzKcBXsG8Fo7VyzdoLKaaF1eR0RI0maoSEG0akRtU6QvV7tBe+smbiOYtj9FGkC5yHsxnVHc
BHmAcrkPfAdvj0eo6H4kC6Va1LJTghRUNW484T3aKQmKlpYKrG6OazhYOtx+bUlNtYOHvY6sBRZl
qD33dYceuExd8nyt6XiCxGtJv5Y95cezakYE+AoXULhhh57uKNVZi6tRHDIyzz9GAJnfANpZ7q4M
YS3jOeJaWUamgUW/TcupvSIvwPUbk98fFr5b/CkTKvhp0V+m9udEIykv5lRg+Cg7/Pys7+lilPoW
MakvC2xjaOWJ7TFehTTSAmdZ8BBpCzrraaIu4vZntKb03rMYzIgvK5clV9keUz6hT4kY8Np/uzTU
ACT4PuE9zrYl9gIqQ6HYC2Qfna6qVrpU741qjtzUNtCEYt5TZjd34aTIcQQjF2BHCFz7O/PlG23t
QVpb90u6QKL2k/gGIYEi+HuwizmRibpeL8sQC56U92XWxnbNdDp027+KHppGDNQ9UJyiErne+o7e
yY9/TjOZRN0Fkm/f+XWtLCb4enK41jBtFaA0sCTiyhhfJar0s4q2cD0GJsxQwGb8HTyTk7n7D75h
ujqskk2EW/hZ6BtgN0gCgNSPiYja+XtyuIvcuFdyynAxwiL5K+0v4IvkChJBs8h9DAy//8L3zBNF
TAXEBwIg37LVT6cF3u5I+YMkv9cNVGnBppjDj/ndP8GRV2sVXVL2g4xNMcmx4es00mgEqatcWkaE
mOn9MgDEeRNSqeWfYXjbA34r1MO0rKxIdyP2xQ/O7/SJp/NVSVYY88QcvPfzlvIAeZko3ol+SsND
yT/57wTEVaRRi5CneSMzx4oU9eNj42ByLCB8AC0orCuXuk6fTSXvUpdbocAs978FO59sgfOM4mG+
tTeUcsXh3enedD2krNOtPHz1AVvhv1qsOTkgc6vkmLfLUpOz9LyfDI9DW3cMR2pApxa9LeRq/0c3
Sg7dfPOwqN8vnwoL5NDSAXdVMg67obF7WTq1VJLg+rtOLiRAvf/Pj1ufKEXW2UvB6HAmGKPyL2WP
+HdYgqqFRJlhY6IVBMtpI/abo5Wr7yG6L98+ILb68oWLiB5tE7oYk0wepwfONu/QYUnspjDlxsxL
Or6kzgCygFKgAdozbPbWFbi8raSyZ98UVPMldhibR4IB3tETEmwvvayFqHgEtD/FMHz7qSDXm8dI
i1VM6UCo5X2SZUyZ9TpBhG4Jj6BODQZlRnICnOAuM7FN0QuwZDx69Wxx1P331hIdrEyCBQH3YgoB
O+BHFEAaZca1C/2JuPukJtcJxpnbWAZlA/IgsRAsVqrmMJBlq358M+eGFxJ+wLFLLi8f3nED2Vmd
aKzSAMMxiksyaK2WSSHMDFiKHrwLTNYAuONmdF5m3DjC3LPb4wA0mGEqjZJTeDlyOAyWaGAV1Pir
haVqJDOFRSi/HgiYFO/Rgv5UDl7aQ3p29nl8L3XX16RKeIq63UZOPa9m0lcl8wuOi/OSqvzrS/FO
h/BjjnSME4a1mlFxTR6QWyIPcE1ybARNPdsm83S5FuUIkOeVbNlfyycS0+fU9TptUE4TUWVnRn6t
9Yi9E3hsEK5Xfx6pwdErRKoupRH2x00bSqdHjnSDJkmAlcJ/FSIuhwzsYhY+a12G/V8GxVHZLNXl
BjQUtmw5oaCxzSU6wO0s5MtP2vKUgxaRVaw3xwIehffAY3p3oBS7hg1sGgnUkERQ4IIYyF7sphle
Z0Jw4bjzB29/q8yRQNmdv9i9QBnRv6/5qMYw68HeJzijn3OdhEbLFLtHBMCjOF62KNwtdfxTp12P
1dcz+02hoUek7EX1f1Ic+xOdlcxEeayH2zgaFWS2ZCGe61R/3yL16Q144HMj5khBH32li07eg+CC
ymNmqilcJKZnBBostT6/uH/O1EtWm6Iy2KIlkesSm+BXpd12ZoW8Oz8zo1V43OpsHvanZKfumjd8
aohCPjnI+5B3sbO160/OMOGvkdF/gVgUh3RqkO/vxftNe82JK7nQMUjgriE34cw3BauWxnCLqQP3
aHMT7vVCinb/zsmP/fw/yJNNqm0SDc8hdMCISpkrNKLdHD5gUaf7uWtQmWy/h0JgqZ6Dvnr47Ff9
/lLeGT6BuQRZ1ijOq5kDlGmgoxS25WztH1iXVrfZ1J5J2H4kF+IKeEn6AjcVqn6h7CobeGKc4Y/r
EOrzL/8GSpWRRgi4GnDsYAAnAP6j1qIf6ZKNQhdXaCZgbZmefl6PuQde+Rko7tDFWtO6kQbtuS8e
xBspDNSdjkhQam8cy7KsLzczjdFLUHcZVR2PtFEnd33gHUEDYOqZs8dWKRlQ6n1s+1Z3CKcKw9vq
ryjqiuN+xJFUP9x/QqJigMZEdjjnC59qsV+TpLx3YZiS/7LbjSpphtUjwBkMf20YRLC0W+SuCLhx
pOsvs1BzBivrtMQ5s8NrXdMI1mgqm9wgB+HwPCQhZoE5VLQbmwDJq0YxyHcqH1YoGx+OZoWI9d5/
DZHkuAHNeXs1LH3LAIJ6wHcVrlMltaMMZ+uSyMGxKgk4fdl374xVvp4nsiqHz64xAE/RgzgGEZLI
iknxFMLHtxeALNK5ZfMG2y3PaRZ7D5/sc7dm9ocXZJngjmfsG+N7Ou0UAVwaps8EnYUtuiJQc6Il
PF53acU/NPpXWcjZgs4LY7bQRtAv5Nx2hnqduvHygzjsbw7wxDY9Bw+AeWMltzqRWIfNkCl3bqT/
9lVredSU3ULw4R2Nii9tlUCQJCl5V3PzB5TbZhk7ETAAngS9muWvtyBYlAdNRGPGjVhDJrIqeETU
49Pj2m2WuYX/aiJ11MBYcgjmptd/pZMPwhOymOrjzq1QlbK0G2A4Redp4rFtsRQUwyjeaTQaOJ2+
Z99PC20uwqgLI3eMB3w62E9y3R12w41zWVBflM1LMGmbnQiyH0sV0Eunq1ljLZ6H/1ZqRHbw97PL
krk4Bpxxb1f8HlAcAaTa5WF7XAxGG9LIkmuU+r1+QUoT2n+27gk06TI4nn4yFA9U5IGGRlwJQzWS
210N1lNwTXb9Drxvq3KeoZfubHbCMcNAkINc8X1rygpoWbmLgsJfC0FOkMpz1GJMP+NOVY4ENJDN
RBdBqq/uDXo9s9dCt4AsaK64roUqmLoys3kQ55tTUhZDS87tD91KgvEhjXd/i+LhH+udrNrSZe3n
19OLJZVgW8bhHj1g9uR7kcH/YT0AOWrFK1c+qv277deOWlDJWbgk5OxaKAJSlnFYrYLpvlHyy3Ej
ButtGlebegbLza3sGMDQ6wn79ZmcVgUVbJOC3sA06lqMqgLS2S9sB9wuHAgQ8eqDAHTpuWRMQUoK
T6WF1Y3XrSo2KdRYl39ixLRjTtaC+yyIdxHWrsyblK2fTHFplPMRaSnPrFzpupxvT3sfsoxloOLM
S3az/e9g7zLFqs3OSydo1ZVm8/zBRLazxg/X3v6UhxR/X2llLI9KQUJz3SLAM3wcTDfyhvjFPdJs
yWMZDTotSnAuLilrZuo2Q6W6FBq5B0/kgb0DsNsTABbzVtIoTr06iEOgc7IVTSMckNXOZ9CJi7w3
cmiuGaByfq33jud1JAAlw5xcje8UU+q5gOgY1VOTWOEFh3eSCqi/obGndPiwKz4Yy0Dfm3Msi61+
lqgZcUrB3MMAYQFWGz2orMbC0j1LBFjSLuI7HAvhvMYO7EEiDohJgGtaydbrjyuarxtoAJppl6aR
lv62HUyKtFXXQVT8tE96etVUQNIr7bUp3oSCkG7URGKuAv72kUNjzDAFx0KtoGUzLVy5oz7gOx8w
izDDCvwJCIMb/vw0RGE8b8DRyPwZ+Q/ditwcZQeIxkNEgP8fOvm7/bvIGe7oExUxHmQ1tyOsQUtz
rN8fvClR5YNXe1N3hmNdb/BSoXi/lKR53iuCZEiU33t1MtzeRfStyICg3NBCIz9JNJQCbq3OSWh+
dFZizAgFniL6gAvg3ItmFJb3MItZnnC7c8I9QJdlcZBc7HdfIU0uvIp/IVE99+VGlaHrUdn5ljW+
rOkP3iCxA+m/lSAM5Y4F7wYa7aycj5enjMIvqWfG0orTqqbarOXNYu8h1EKWOFV2uifRMMpHX8nN
RmL0WIedJQB0lXl+f1W7N3VW199EiPHDmS76fajgQULjdGYeNXkWGXQhBMBUDetDfTWtCUo+zCrI
IHoHfhetOZgiSOFKZ8tt1gnRGwyEWtJlQcjqsOQTZD0qNF3nWGh7mm2gCP3AxqbEvHg+lCmpt3gA
hQhZQpnmAscgHHeqvo/r4bJzwWLEY+7d3hK9H9H6S+hGU9BPwb/nPVdNZGiH0KspXOrwWpxluA2/
etbxvKcQeh+yxs0wIa7wHtZFgR+nFpGNrOU0zOUIKF2AhDKtB/BQi+IpMwQOw4cZGaKzTW67hHVd
po0wrE4PxSiLzmc4uczcr5NJAtW/1Rfw/k56lp2gS34XXCwtIIJOLVCmQsL7Kq0aayXWOuWjpZPh
OXI7lwpdn38Jvt8pKw65nEU7J3zn7BB9chrUw7hqMlqylL2foWwxkIlR2fC3M1XtRW9irf+1XYeU
pmQlxFLLQfPOjCfLyHZAkgduolAX8L+5IFEKoyDF7m4urmfmR0bq6xZRWxKPROEoz+LHRkVsskTB
Dl0+O2EJGdQ+RJEBo2ukbIH5Wj6FWIWb/xURMelzxnm3Ugnnu1Bo69AiMT2PLDAiDD2CS1YaMR+D
iafEW58aEOuD7Gy2FkOQFqXq2ux09qMQG5yvMco2EVkJ9gXycICOwFnEeyZM7BS5Ow7f5KvRs2vI
NRBXqsCj5/THoeb/rHMUJaZDIXj7cKQ8sEJ6IKSRN9iXN91RqMFY97RIPdxM94h9rhY7ZKEWZUvm
4s0F/kC7tOUjOvNcaeP+UtOGYKTJSXK8FGx67EgDzi1K1Btxai1NYlD0pAKUGamSnFcEqXpLt09P
wLzDawDEUNeMMn30/KlX214hCHsv/lKeihqHHMWgAN4M1F0aGufOmVHPrdsGT3azBFF6jn7Sg4L7
9XhQ8URuQvgZFSfRV0rC8varL13KEu5IPZlZVOyYNchcwjoCsjqfYht0mabT3IfGEaMn6kkZj/jc
ta/Gn/g0Xigbon9r54auYP46WAoY1gm172GdgMbgVmU2WtUjYax5pahFHepMUBGn22wpwppxS8EC
mPjBLe0DPnlKCz+eiKjUhlfDOLG5gTT1bVQ8Y0JiC4eJJQ9hLBlmu1Sk/VFsDpCR5wr03TF+niWq
5qtBuOpmizYCiHIL3RbS6W4bN0REqEkYikY7CerQQmCdyfYm9ggbviG8nWJqUinYfEswPvivVxni
BGCfSqlUaiATkc87XgHafDkRKC0BD+sQxwU9dvTMYhl6x5nSLs4L9FpEtQKZxWDTqU9DdOXEjJDg
0vDHFk2HNGxZGStKUf6UQyHtQmOj5eVLhZyMPyo6FW2h4mjFEjj2kHpSHn3wkv3R/UzCTqmIqFty
fMa58hd139yLbTMJaznUa/1LvQDmx0dgM7kmY4D7pf3JjoVeBWrlgTZuLodOyL5JNF9l5Gc7aEIa
LkZ7uyczrFhMNNbEHK7gX3zIbU67LzOs/ubjuleRbAJSgiww6M0LNgEKTLR4KPmOqtKZAfXlWQKQ
kCHArxbYlA8tc+Xzm+F/WsWF3h64l1CWAww0rqkmD0faehjDwQHl+jZbUrI/neHpm7NbaFHMq0hc
y3WvQkhg3xr+5BwVea+mKV8NfawlRzrEAOnvIrzIbYlrudxGERZXa8/tKwLTGj5yyKCmQMEPJFXj
Ajeu4QsKrEpMa5exiZUCl7Ich1NMVvTnSEFb+1sQLJZ55NIySvl+y2bBOHpxKfwMRsqDgnY/F/em
2LqZROpUQL/7N28BaZbr0UQp4o2XCKBaxYu9Lo+rVwnYr2QtNr5XoSpbY+YzE0gYL7jSgguJIh8i
kafIgXnMCoxDNW4MPGBfEOdiEsggOepX+iGj+Vs2/sd6WJe+5hO3wcF8ume1ikoXXt+Ggo2TgDEm
r4mIgbMX2ni8TtGfw2aTto4vzbZvoO/h4FNmD8H/y9EoGpxzJrqnb7uvFwqTynv2qTu1hU5Fa2Fc
o2bsJD2UM7XvVY7xbzdjYbMHCzv35fjkAF95J2Vi1E6UPIxA1+8E0k7ZLahWqUmN2PgVrG+HGF7m
of6BvnHMcqnJKi1qZ71l1mSRyhrWkB++jy1NaC9/qZBFHSmtSeDLogiPMB1tLOynWs/qa6ACCkTO
r91UGFUH+QJeqfWBCqKFtuEl3vEdAOB6Vp2zbBl4ElHWxL/1QYfMy6Uonflik1Wzm4jFibAHxxN+
2RjDYAKS8Br7MlpKHlBWaNMIU5zo7m536Hofp0MX+VO7yqCoqSo0ANqedbEU5dYipd1pUSyRS/3E
zcEy15VvobNTqXJDYAPjO6ALivURxtsQHiBaEqVkwcGDmpEQABqQIaTRY8lgbPuiV9lKhuUOAr1f
7rv7w/eniQfRm2JFB0VEh8nBI+QzCAQNQ7/Hd6LgV8LkWAjaQOom/khGj2JOhbCulkQhAo+ayIf8
7A6m/QWCKIsTVces82u/ZGxrxy2kngYD1wMQ7YQd4C9pvbgIjCx2ArxtjfAk80hPNqQmlFH+WWn5
zwP+PMKlZlCABwUIhIFA0EfAKLUMHmTOKPMyin1SYkQjaRDb9B0nLOKSkCd1LOVrOCn8/oW2vz/a
HlZH5Z2quCxMkAhMic4qtPSZuSQe4XwCGkpt9zNu5m0LF3aAZyLp9isOPTiRW+J/BkPh23yTpx1N
iMYM8uX/qfvdTfBg5xBwemFMAUbwZtNU8jjDsofm/gUb1nhS2UQj9L3axg/y6YgIPYCrmrsy0n57
KZkmFeQH2Yq8EjrEUv7VAwQ27nWKL9iuhsoXV4lJRXktMK+H98k2sDMCecVTPAHH3gvuCMVaVSI3
khvqWDKUBMaZKzvtDR4QKCHzlgPXdi9e4cuMv9oKiy4x6nBxY6kdVU4ei/5d7IuJ2NoRQRKA5Q3F
tOkOsxJO429jPcUY6dNiKO/533q9W0VoYFq8ZEvPcEn5JD2EfxP2RdkDLM9ORjrn9UI7GwYnTVkL
wPin1UqBs0HruAtSfBhPAy3/dMzGs6Wffof2TAtLzgCnrqsFLoR/tZC5dtZgdQIDTorWK1MRKB14
Iz5THrUkcIxLRsKFt0/l5c/gkWhLBP6at8bSuTIOpAwXROL7PS48eX3Bf/fltPb+B5ehmXXEHRcM
28+QU4QMZpObzfQD06L/XIV7W2hUXaKFW2viLMFNCmxtNzrNp/EnmLOyRIYdCymi/VlnOmrxqagO
zE3mFEdm2SWyWRM43ufj6w/TNLsWeqZhEJkKSCGSXo27FK45n+s70fMTTh6A7MdXq3F7YapLnxid
WDINPzVtjvu9OZGLh9uzzLE8k/9Jhuo/wgHy9QJFQjUGgI3xX3a2nKCs04C/tBuhBINbc7XuAAh1
RAmA64LdIF5VuX3VsIB71ydlzcL7k5NPiwhvZt1WDOSSfiI/fBFCGJl//PCMAmZgmLgfbW7Qfpgl
5bJxoZnNdFpAUcaxmHvHeZZhcEMlsFgeaQVEb4lpCnd5ERvRpL0aN5L80gLUhmhuZH3bUu7GoH1G
3KmZ+qa1/VQ5F9FzTkrrmxdqmFW3iJNh0U9AY/DSxPoW/8cIH5W4FSN/ifWcIqHzBNy/FPRITuAO
LPHq/fsamIv76AM2kUmxSAYw3JYwSSoNp/05EOdH48B2CsHvuv8txi5wGtNZ031zskp3wJCL+Yrs
kAv6NnQ2RS36LzK8cwUrm3A62jnpFqa1rfqd6/oYt4a0mfcA0Gq1lShUkTt6DeEMNDlca8o5CaRG
aVHNSaa4NC8G/UY1ipx3pbzG60cK/FO/raBTkjXZH7kuLGAfYc2oZOUkSkULdfXrwjDFj9q6FhJF
ob7zkck6k4WEMpPGhc9xrMPHhs69I4kJeKWfXjCJMlwH5gtXTVXCMqYOBn/ODX5/l270la9FMuxi
8I3fDHV5sd6wv2kjXTZMiQcP2KfxulM1UXWv8rCasikan4repAnXYmUGfGm2Z+n2Zkegpbu3sS9M
3W99gxroUCo34MlfIjB5H540T8HUTQTLM3EbZvzXWqvyye++CZE3MZOZgboTUnGRg+75TnZR6dbW
/UNqMUQUhxBKLK63i/IuYhIKuPTszQyy5aME9DHE1zrjnCtsfD50Fbl1xP0slkFWF/bcoVxw9PMN
gOIK4eqpIRITBm6xs1d8SdC2PotFlsLgkxVCB2ou0F+wnn9UjldciTG3pNkU523jdV3ibwzrj+Sm
J04aYZKA63HHbqUknax5hF6+c2gS1EJ9aZLuy3z8CU4N6nFN/k91UXGmrgWHFhqItiWTEInrFQQ1
4Ca0yRnqxGQZ9zwHQuv8JyEj8SGgf8jxof/aPOR4POG2TQPLOJmslQbm/PVYfhK+0h2o9kt1d9gU
ynNZQzTvwWIhbseziu8pXb1gpXp1l1+bxRvIcLe5kJ4HzXIaY8fdrnFdTTrcGx5fDhy5djm+uioY
xynay6VgkDEz528a9FGWmxiDu0UBwZL6bwLn318uaUJqYtQUZt36qhIbMS8ibT5oiwAQ+dzYm0HH
qmqI8P10GMkvWz6vYdw1eFqw7xZXRqMazLVVu3K2GIjjTsLs8MVlzYgaEkiAo2Gb5FfruPQhmNMM
ZZAdCa/I2Ztb77nRM4VnLduZ+0hv4SCOklr+mYFAvht3kV2GVAr9H/NgGB7lJxcWfQXwt2JKeHVU
qHUuQBmlfFuRbjaKe0slF1nu2c7ka/ynUDegtBRlfr2vfL7OHPkK+K6fNWSDSYV9eSK/16GqbsZG
T/UOjrgPblR6VhHplAJumY63EelkddLvGtEGBOD/K0inHLyoXwWbiNSCUI93X2oVTbsKMKvGE7GE
/Pq+HJz6k5kHWDR/iloSp3KkkAMvTwF1RoGFGi1KmFGW4EyXyHtUbXuOHcD+cj+THWy20FIhicQf
RY+qk+BWhpAoXY41d12XTbENY87xMuSGa//rbpsvUyt6Tlr/wgxudIg1Kr2e3WMFmABdUgxPy7z0
I8pw0obYzd5/fziprQ6XI8ynXstNvJW+RUAteTuEsQKcpFbGEZNz7cUiNZMT/56BtDZCPWRIVhKT
2k/NB6UvDNlWEpLyW7/qcEsqy4T4XLUvlzW6XcjYzZQdvv2vX0ylc2tj53GBixAB2N+Kz+cLnlhf
QPUvOOhG8PWnqrdPgB4pZdBho27Id9Qk5nIDJYtCGeIM6qXSIXw5FrGJq/ev+LcNnoHvNraBsAp5
d0SLu2aQdn24sJMzas+3q7QlxiNmo7XqFlFRJyusDb0OR1PadbKjAv7wxabQ4ueB/02kJa1+M+Y8
wFUg+dHojjMgEkstM6viH8WOD2BH9s+njHRHPOreI9ufaypEEqcc7XF74Vf3qxk6Jgx0uWQWTRb5
HWaieBOWw2ZG7fzdtEnTdJNdWhe34I9Km2nugM/4pxlgFSY6B9O04Kd/ezYv27ye2TauKjs8He7R
OdIpz8dQ3Qbc/teEbTdbnNpqnzBLhDGeAXlU9vqhBXj1s54a4peqXdlh+Dfc9Xk9pSJ1zq8l9XuP
UuFlqsJkxKxCecdqfNU4j65a8CVaCodYcmH3JAuffw80qInHG5+8iiBmGXi+qI8ON3gNrSl+ZKFg
nF7rkET7hk2AKglkwnPikaYXinY8G1DCOg0vxrRkXQ8Y9i9+IO65VP9bRfcdx8GraC1YDmXSyeDh
pXPM3LPtuvL2D4BLseDYQ+AfVI6pfbF0WbJ29zRdB/f0JWuiOXBLZmfI3PJ+X9ZM1i9yvYCj1Vr4
Y46Ms/W4pxfG8ELHDzycN7rIOSAnnad5QDqpZaLmJFWkn9TLLGbMvwplv5gHUeYBlzdrJbpLTa8b
8zz54Fh4UAfseHMRWqcB9HJisOusU38lXNM/tlBxDG7Zy7Iq/7EO2Z7Q4sw4xhteiWbWP6BQv9kI
G815bVzWzLax6/s57itWkAOvbK57Ips6v5hDvOdhxDU4De3LKznmCSeloOtJYEAyD8nxJ2WDiAfz
7V9WTiqOK8wxOE/6vpF06P4sFQ3SD4ucjiU4X72UGQ3wWdaafvSyKhbxKNgTRx1yR4QOuQom+qBN
+FGwg/XmJ3GOBePTOB99OBCghwS/h11uak3srKF8LrOFD6O9PN4xe9eHkxQQQDTsg2zw8e/5ByS+
xV+wj9y5dVuDS29vS7IvrjEYyh7kr4go0PkgSIiT4RTT03bOjJRJIyW2BBj0NTKAdGpu8RgyoGWJ
CxIqmflsKj9XYvRls0IP4aLs3gjs3jyXJPgbLT96CpsSs0wq6CvettbvcCMmY8f03DSzv8Pw6up7
0t/xHkoBXeUQcCmMYO2jLaP4hqqNsmrCGc1MZKzVjs/imXabFIGLehFDCHxg4FIuQXMtr9ZliaX7
4nT3hOKaEQEWhxNjUJcRS2GiTXXT/ALHVxPlkDNL8ljwa1y49K/R1U89Bj6j7jChYDfr4fVcrM4C
VuFWWdY1G1uhS7pn4FRU+7cyKn7igoI227119oBXtDGS4TWL6QbzRAaQwdBBsKhiXMR27/IrMssp
Q24rcIZC08fmB/2XAeYj5cgNfDcvPns9DVzbCPiVh0RMA3xXXF1Tzy7OBH7fnovsziPOO/zlQ1Pj
b8FV+nPOlTirCIhrWx01ySi3AAnEo850CktvUDRFLPrLIEAfPBibG7sReQ+0uJE/LNSgOwKV7Npu
vUFzu4qctemXfAxhhhxirEkYiAeRJa89O8TFw533Fr+Eaa8IRxchkzBifiGf/yx3T689SZN673Tw
VglRDDFR9V2Wxzws6Gp27trA8KHKmNVqOL/3WKRXIHPO7X1PWLB0XUNHEPH2HNsdjwpgAbbdIhtv
YtNz6bJkQYrTAGcZtASNw75L4DjbexlMF1PZqHl+O5Sw66W8+GAQmqUaQZPDLEwZL+5Cqwtx7IN7
/D7VEF+wB6ddU3ZYGV0B6vu6CzdZTt/lz3w+uM6a2d43N7i27H22yrNIJWjDDGiji1orT7GXOU28
rdu0MYIewqkU83yF3GCYhG56tMB99sG660P1XVc/8J/A3EpgpYfmwpeLNF5V5KuyScakb+hyFsVN
PP+iKI3qL2g0KVPV/DVbwCLcEkMshkY3tVGzC+ELAnyuJ2iNEuzrQP9Y11iD+Ivfmobtq26bJDf6
x4q1cXCXjx03NNGouCPGLmkltAdNss/rPLQ9ZRW89l7ajr/8/YeR7pTEq1BXauVvBES7Wi5z4F91
t2H0oTL9SmU2XWIhxvaJVRHMFAq337GMKsXL1aSBc58Rv6qDiqt760dJrL55i3tEVGxBycY2veLT
1S2HuBufeZZLa0KzhkHk8FwqxuAs44puraHQb8NOY0GGCSYjDJhxpDLGJ4lT76Un+UQ1Tg+FouhO
Opg6v2g5YLb+U9vc0i8nmEmYAcS9m2AMXLzPmeAm4b1uzigmSOJRE4/eFJ1CKDpVXHBsv/QM6psJ
LCWhXy9S4Y5phjnbQjtv3wIO5jjvPnleklMU2fB7E+0W02Gd8TYZslXhPXtJHCGVK4EwiBtzrc6v
/Ch8hCvoUZcSr2vx2mKnppBV1iQAkwjSIB1VK/73e2KubqOoRq9CtaECdq/C+wU9bFN+AzJnGdp/
IcwgpObQL1nnOSON2B3L6cLWvTvuSHTIYZ7pVlA/bd3dqS7WYKM9JktGuLLEnZIhXPIbct9PV5QD
byatwzcyBU3sWf1Xsh8bucSYDRiXF5ZOzaIr6bJiyuQjk9lKqFgg9Hr3afxBan8PeQYq+kcfeaaI
gNBBOVK33cd7y37H8eFyqXsyPqtV7Xb6deel2uFHQmqUg8ZFbZ20/F4zfW27F2vNKv2wJgLOaVpu
uXiLdx2toc57ZMxD3DAnSAHwDUzDlNKRJNYo76k3YN2UTtBz/a6VMw1FQ9qRcOMAB5lQQ4E19oWh
aqu3NCGHO8vyVBXjFiFfz9RG9pKUfiDTcd2TpWnvH95pl/0/x3NbFBD6CU6g+ySS6IuYOYOVNvDd
a91rVXTubkQpuTA9lQF4+2HeeYy885bLlgvCJkRt1Y2l2hLmVn9gFR3X4iAa6RVXR/QqGJ6XXkAK
LmzZBx7hHPC8DnAjc0MG60J9fiLkvOX4veTmwrXRiUpQL5j4XOnmjrvSu/ddkYYNVPchUNmx32Pu
5wRe66k5sIguF9wRt0UvIxV2Lbz6j1bcQU8TgBV+KF1LlG1QXYgYNqkxRDKdhpp+ozyaf4XBljwl
WYUHuckqNmac5154oN5wWm3Flc/w7EAr4WUG7dXyTLzY4E1UAlrCeUpckKP4v+c+UJ/mCUPqFKV/
TghI3rObWImwaRqLuf8SiWwnpuNYSyYepOV2Xh7vA5ZuAR6/W6BrrZbVyLlTOlxxKcqy0KN2mvbN
rk9cPIRHP5vD5UzRe6vT905uBI6yE4dB3dHTZxxLkTL61jCRF4hkJN87OuM2Dz3kYloQ/xKt0K+i
aY6Nh36Vdlbab0Aftpk6vVUyuWzohptn9v20e225Gph+PpziJXnukoLD5R5KZ/I/7W67E88kCmQT
QzVnDJ4wT2Mzo3X6PcHOnh/Fs0ETYAAfXoy+a4kprnSQwrLcps1kJ+LVS2kyUmVHvmdOaYn35pyn
+LHrX8glP8uOC1NVj0NOztrV98rbAa9TahsuBylDHWjaF1tqqmdZPQVEkJ7SiyKPlcPHfkcWxcpO
r8QnUHA8dse38JESa0g6iZrW7l6pQu1b6UF7NMW4AiAOZhaAJSVsi9rXWTwIXfUPCJx0ydfIWPP/
jJKgRDmtR5B7/KkTODg13O/hbTswRErjurpMC+ckfUscCyEKe19pMgCzyhUYbi1U/xHxNBDXJHql
3LL8pkoaxyQGwciOInwdtypC3F4oznvOpPYsi30OpstQVbgQez1Ib9XwMM1SlRP+7ypXVb/eFJKg
kaFY8pbITFOAZfmpZWjLW2jXBk8Zl9NskOV16u5mGFLBV0bO2yNFziPGxIALm5xQLoKO57UBIhWZ
FbFawzB6T1TctWwwfj5SMH/FqGc4z6hkeAEGYF8udTQp+vQ8Gj+RVkA5RfB/5PgAz64VEDWJPvdt
vHFWQpHPW1pOJIfkzoxT+hOAgiZu+LjrQJBZAiLOy5qxG7VCrKzYE1L4hvI84fE4niFC2wI6A4ad
+qQQqssHsFWYVDE6G113zow2q7rgjLUyQwNPogbMQP7d7+Ff7fKnkM766WFBZGpBRD114lDt1z9J
HppU69IYvpnJl08MR/cG4MhTnO44m1e2pMgWstxqdkMjc9aaCGpsrnA5lipUspp8IEvAtvGQBEuW
15yjJikKmCJ/jsgBSDuJ3bxbj2QEiLmOBGYCs2f30LvEvTKtDvijEBvsZKQ+nuw+SIaYHKYdIYnU
eH8/Fw5xvgZ+67xd13fLV0fQHr3aWEg98ghrtEAd7+Mq0RvIEmHyucwrD1VA8Xb6HUmMPuOR0qbo
ecU+DHFXccDa/WvaFOfrTutVDtTJRuaEYhWomyHdChvk3rABFfNvHfgnUwVt0FLMj69hvrWLCKHh
KhynRdQujBF8upRwV2OgiXrTPQuwAJbTkQA3Cnj0sYrgtLwkxofs2UMvfMZMn1H26EYRee7q2LsL
GVE3l2qzjuAo7yvqjToxoR66fxogH+1khB/TFIwtY+Xy6dEcJri4BgvrkwuTCrvtZLlbhGATA5a2
bFYnGZ3e1+NJMMVei9mkV9U0VLC8HBdrTweWtWjTcv48529eQBItIUptdqUZOjA8/xAzuS5eNauN
W0cVjNKwg0ef8k5qKgMIB0pgs1/BvpfswhbQRE/VUEpEmBDcT80A5fDGj9kIHsXWQ1FIJGUGp00c
FRvqVfUKgnaKRLrEwQX8r3MMXHVoZo9L/bzrhLewq1carVWhGrPtFnqnBaXamDreCKRl6DvjOLgo
qV2hxcCnVP0I1KlrWTPjm6mjuWiOXdCNf1aULOziuxZlizCi76so4O5q+FsoLeUuflyb8+GVDtsH
DHMAPAtoLDG3kpp13IVqCoMzdT266zV0a7AAgry2LGPlWSeawW7bwdhhuQBDf5ezYN3NgOOF08gK
ruWNg71vTaOXEkHHGQ0KQPUGRwP2C3Ff0009pVcaZQm1ZGkjIBuT5xeg6RK7ibbWiuT2C8x21r3n
jcO+VY5LtSRpDA2VbI0FozX7fL7qPZmW2woI3BBWRcWT8ok5ZyNmRmNo1h18qeNoah+ZMG2vpoSl
AdA1yoRievNkm7+ZlCHH56YK1UcaZ3cqhAdVdy97cP1ehNmYn4XLDdWiBYpl61tg3ye3e5Ypi0uD
L4TxQdhvRhxvJDEyNSYZFxUPYMS09FNOljjIkbLu/F2NxE0ZFkCxtPNjsvS2+b2AEXEJLZ1c2W7w
gQ1M6GLrDUSjW/GojV165Pijsej2M8dj69hHHcwCZKRdRuaKrZaW+W4bJBL/ENAhVn4e11Yxbnvf
ePJvzse8DLrb/1wUlRNFCvnwGfUD1cr/yKdJMEAn9YOQFsqhAMwhbwZDkQNFCYd5yMtBN+a5Um/4
cXQiUBpHTT15G4zl7+uZfrQ829G4GTHQfkuNMapNySVucVl0Od5R3uFVtAxPzGRGeSjCWI4Pw+1J
HWoPlRzAadk8Tb1YQBu/s2/hLNiWJfveKK1ef8TQZiSj4a2p6I3cUOTYEFL4dP6pPMePgQduc/uE
q+ZTxmJ9rG8mg8gaaxs5CLqiB0T1U73Fygq11ikBsawuixYLOKuGhL6qD2zy0/Wt5zYOV2dj0tP7
VOp0Bt9GXnd8EcD/Sn3LYjixdAdHKoYmfryta6wO/xSC5kRo/HxTMky4SInc8GzUipxCUyTvvBCY
GPgStlwTQGcJxEZC6vF/2h9pBWys+i2eCwCZAOSedfUSXNS9PkXXfAGWkC4qhBztGLIA/LhslReD
wl1X6LAg/NgWfl4XU4Icsgoy4/nj/5aSMHMUqBPeCG5bBoxAhcG9/XHfes3vzWJYq9qyDxkUrJoO
K4zH4Auvv8iP5rjMFNpmO43mkHWYRFS2VR12EnQF8DboaTwYIoUKkWCtz4OiC6hpv/LfnL/p1bR+
86o5+bD2r3F36hju3TONIFoKKdff1wDKymXuxJjt7l3JNpnOpgB875ejpaM2I68MhxlnUy9ey9Qm
cGpZGUSxpsOUwoFvePTvcLpLxlHUQN0gHgR6v0Ms+2Rp+c6izPu5ItQ0CA4w9CJrAz95T1XK63ug
A7yVK8GnrbmHL2QU8EIZCAcxekbIFHk3A0bwx3TUFD0vC2bZP3z11ysF2q6xz+rzBRKqilAkL9LK
Te8A4r7bfla32u35/EmjKuQ0LL8lvxAaXmszisarE8ELwcVF0R2oo6zlV3EOvHgXEON9Zn6MNn2X
+lrypimB4JYIOUmV9YbpDkCWrsS+dsWOy/jiz5ZVvHy/3Eg9YyHb2o2qzK2c0grLa30ZFsdRopd2
OSx1QTaNdLue4Qzr2L4ydyPvVI9mKKdUk7KuHN8SDnlbW3LgQLaGutkyr7/9LTOCT4CWi3CqUoKS
EVQHWRxO4a55Qzc6ovKDajiui1kOc/Ha0SYGx8fk4sCpMYlb6PP5D7k6enJvx1s4J00enroYDl7W
DzDNSEmtTBnEm5ZBqoBTosII9H0X2HwKShx6kGb5EIOJX4j0jhM2Odzlu+QZe4u3NvJ8v4QZhtLl
McBskoPI36XPJMxdHsJbbGZB8ynU8GrCNOmEs6lvx8DMLMZPKx1KEPFJb8LW4MlGtAV/ifog8hxo
qR4G0Qcecigvb1AR9AJZGRwC2CHETPnO9MDzx0srmqQzuVJEmUbsbFq/vAQqbfk23r9f3JuThBhZ
qHOyXz01DjlmTHc0SY++OqyLuBorwdaTedxsO+X1CX2syKCrRzw99h5D+3G/AnCeUkIjMfNqGHv7
vT7xciGAd86Em3ntXKfNM1CYTZuA2MygBxaXFAcyoFx0u8S+zAjCW3/4wipvZJxbjA9+7Y+zk5tR
ZtKQNL12y5hakz2NJS4xD9buAItKtJDg6oCRBJo5km9K5cK6iBbLGBq8njIhwo1gXmq8/Qj4D/kS
PmDwIcMnZy/UpGaqnpgDxiSGfaUzKP0hfC+AoTIrsP6ptLJrx3LQZ6qgycs+TXekxF8/5QsSZzbh
ccIK9rh5QLFzF6LmK/wXpZPjdhz8BsnTrbJ9DES9egmDonZdGrTtqMPzXsZ1g/HHMOq9NLK00XMQ
kutS0TAme4RGCeFW+Auz6JJkXr3aHLtwFF8iQtnfvLwpusoda+BAjz6nRbz3FoXn1ZRH0vIQlDEY
HzAf2xYdwxqKPw0VHsOHYgIwQHZvhgWaoz36sUrDkNsOnw6alFIwoJfhfmJ+G1wWNbIdQtFqyz2t
n/4c8xgs3ZggIRkJpDPmWbWKVrBbNtjhjI2OV0sHgGBFTDqNSH1Dgsvi/UAo1tHc5HObPyFfLsh3
lwBSkPptjKkRRv94h2xLpggyZAfMBAKdo3loIfnHZlOYr83/MzGX/iiFJhqL+lVsMs/y9Weie7Zw
53fibtjpgVwNdOIadal4pc0xUUj+RDYhWYiIO0y0MaOhpYPkkd8BCrLqTMWiFv/KA1EGIf2B1182
BO+ol32PxprnmMmv3zIK/ClfO7cSFMuh5PPAALricA3kbJeI24ImQmYjACAvDOrBkyIOvHyXUcGA
ydhKx6ND0A3nYVAcotozTYYzO9FjZUTLDf5BMgnp6bBNp9fyDKKkCgo/ssDVOUKpU0Jj4gojDeS2
F9EvgZ1SpPb/8nxIkazJwKv2hFqoWWaMuBWVEaQWXVvY2n7I9MCRdGZuQHNdRZX7imqDV4GMC5Mm
CGF/TDE5L+CnWpeiuPxHTpKSDOkA6qT2NPDJh5PD/FaU5Mhj57D30PolgJft19swQ7WJypepIrYv
W6LGvorXtgGDNwhmjnEyAgFg91vMIx14KUd8CRv5YDj3U07JRukjGmtLamwMgUmMjY+qTdTDDQFW
ENCJUip4WcCPOKqUyQ9FcB9QylU3dtD6nsjsavteJGPlsop3GbNPwVZ9/s0nArqyfUSqX3LHoY8C
j1EOABYRMCnld/mCSQEHapbcSeSESTG83V9oyh8XKI/3OJ4yfcO7eCsKHNjvJeQ9/okH0TDoHl6e
Qro9P6Ziqhz8CzDL+OdLkK2X/En/9xdrRDhnC5dxXp7GRvSACaV7AMa652POkgT3c9ZClMFI9c8m
nhcQHVU/pSu+EdoUmAz8S9I8oWRgEDuFiNOoHnN4ZYyOntKrtD5W98iqTY8c+85tn1ln/lwuFkYE
mwORTA6oY/3bqqss7OO83PWde03N9fZfmOoAU46diVWQqICd35wljqq+ZJANALu3USToR18atcwy
6qDF7ttKiddsQUCBMs93LCCUKUBZKr9qyNinNX/G2Vb0IyrrjHWab9QAjjercoHLJhItyN0PNThR
fpEEyZ7kvTB9AJF8PQ/ijjm8nnpgF9nZPV5dLW0iLPDSkZu/nCv3sQkb3UAlFnwIdZjVyTBHVW26
OPZ0Y6hg30S2yLtEYbXl1ISnyes2+Y0NZt/oFotKjQs1BAO0x6+AksfMQlFTFE+OIvga0OfMtNHF
c6Hj3BoT7PJKsTvAS2FHLrEKBKRpsIttOQjaBwFCe+CICSXlwtSD/L0NmeUqNLGIbPxrSXm1wQF7
tgIk+Av1uAI045rSco8+SdAyjzTf8xIHEaQFPZhSD4gB/YBD5MnHnc/OVoxBGyJaJZljbNnwwqfD
Fymfagxm5BWQ7SClvm4d0ljVrApd32LTWWFrva4zAYcj1bVQ0iAWNqq7EQyb9/aPBNiC1bWXwG0S
2H5GmSZ0RF0BKG3TZNx6egfjq4sII8crZdd4POIOKj2UP/vvArZ/h3BJe7z+t2mk3E4vi/L0zIwc
aBipFARLvxGbu4CnFDYF8NeSrnZNDUdJvtNI2KxpKYWVmC4HnibA9r3xHWYydM06ILDAdNuUauDk
B9tLi8wL767KVd7wc5rTXr9jFf72x/bBIoOPmctYU7JAuQ2mQsX76mwWoY01bE1DYGVx/xydPS/a
9VYZZHMsSdIAsKVrvBpxlE48wQYtAplsce2bkOI8widHUF+8U491aaW2FspMeuFNS4JbG3pzbLLL
JLiYyuRIiC3+z6anvxj3JBGQK7uWjzVKy4loLEHO1ZU9w86aoqyjbM+eKv3Z7gYmu01ldwVfwOpW
N6p/GgZYCp64UZBk5QpaG4W5305EEqvmu3DtM0D/hKyjvKR2MnPFZJM7qb9gtXcrNWra874IaCrb
/IOkHMovJDLG6ehwrFWOlTu6VBeEsBR9aj14feef9ZX7nJPCT03Ih37DyKF3x1+nKHg/UAyGIndp
7BvKCdDnBEwAg2QuUBntJMI0n12MkLR9fPrYcHCflWwnyHTBbqSgGG07hQ15ivHAQ55sTOxydVcd
9amcC/MK0XdCQqNU+s3+ptPPMxDYys7Uy5u8qbx7ZzEOAdJG7ScFTaQPc8YnitD31zSqsgx0PSbR
0h+tEPVRgschf2BciebArmcwGQC2+Ixf6cLDP7GPgMrtut4kPpbWpaYm11SepYtF01j/zsmqi4tY
3/UGbVYGsE6/eQUodqrQFVVUHdRYJV65zP0DkfkbHj6DjHPrqSy54TIj9F6MzutqaLLOEafEqYiY
clXZQYLA0/Nn/rJi+qsosAPRg8ohlq+il8DtTrTQeqPdP2z3FzyCJ74l8xmJ2xC4/RrFLeYnE/+E
SNlR4gx5JsT3s7QahMOZVjrhocIW59HZkdgnFp+FkwXJ4YaET3adjsmUhIM1hNly/8DVYzlvaxqV
4q5H75JVTCGBxRZLNbBKUH8qidb3qCpKxEu+gw/1JtPx6x/6N7WhteHR79/xvi945xqykC9MyF9p
YYKGi3PEdgrB9Zog2XPDTUaXSoKfHna7v9U5MIQyeejIoxX7gfK/7kTLftVZl8QcGKL8OtkwiraB
El6anNvU8JNjcGJwsaLnS4op/JcBSzPItErQK0clXgd018kpusSTaeCdp+vKBC7RuXPwbDRB8q1A
Ek3IS01wQjbzf6YozkRD3BzTUZUXh3mRRGnYhqkpoMDYvQAiVALxmHB7tzXbdJicso9o1Hkx1ovf
0H34v6r9SHVy5XP7dV7Gc88EKQ9WB6wB7maHOpewnxmWIUaymWufCBndHwhJn/xVbtT7zKHXkpFV
+K4AX6hght7xUAePSEkRVIfqvM7iX04upON6dE3cYw94IQ65ZBVkDbIKA0IJ6xgo9iofnnHKT/+R
X/6uDCDcy8CwBOwTOx3Vpj3K03TWtGl5mRuOGw68nMTi7c7e7g2T+r5wWt4hkbYkluRE1C4oU8n6
hW3LZ0AYDPQzVbkV0AV6qgdqyvrpP/AnQXSP/idZtky2imwsbG/r6P5a+8pU/zQKG6v1MKV7OjVN
lkNIBKVkVxkCgvK/GYsHmTIrVUj6g1P6WPNd1MdwFX3W+oI2G9DhF/erI5J6EN/ogEPD/OSHF2TC
m3tFQizayiETCg6sNjPaf8GR9X+Ts7FdMLInC7xUxs+qPSDaFeyCk/o1AOWz/p2RRTCEbbSjNA64
qf0D7YHYWqogbP27iP9x/N1fVqmJkP+k1yvb8k24VxfZDg6zr6eUbDfRDS9hLsBVl8pwz8uyQEER
RCqfxSj5I3QOEfDrUIn3MCInJcrqHxYB5M95TEmoZf7Hn8VFW2F4i5faSpqdkli/izoOgD2LBZtX
DVhXpkLsaTZUJYP8DVjH1PzoLz5RLb+jURsX/qOU0Mo5lC17SVivVVCl1zkY7jMpdkQfsQ+jtw5E
2zGzPjCiZgujHnL0xrs758evkEQ+kAql3FjgRAXth9sjJUkFHgUUPmdJnNTiH01zDOb9eTjGEPlb
rumu4QJYEtZeJGkoO9dVAPjvJK//nYg1Vmz/4WEWKiI6XMNU8aS6ZKWS2RpxELv7IVdc68D+VUep
/PGixgkof9DpfaGny0s8TgbK1G1cx1U5s9caUbP86dlDognATdGDJqnDcfDJIeLVfWujBRsdsMqe
ROYF5pviClWRDLXeCDA7VL0CV2QF8YUhfxKPQDbejWJ3fJb2KCsPg9hr40l74ERWjy/dFq6b32Bo
3fFxmaHjc6MxcBPBP5c2eXSIZQJNlLcKFPFeOGhsCUAhnxs6dX/lUhvOZ3oLToyrCYAWrjvfQi+U
W9O25a9eRrM8dkBgpLvhoc5iomWFWFKgJZiAL1S5uoDF6QRAZRv7qObV4TZkAaGhPV8bbZxlbI4u
i5QRQCZCYkrdHOAiQWkxw6F1MMHUV2eqim6JVPHMy4a5gFs/30hWoHcY8Rwy2ykpS4Hc+OyW7ugL
+TaI+rdp0TXmyVhEI2Hse2lKw+qoK9NJGgGiVQ52QkJTbnxSdGC6/3gM3mXsCwT/3vfpgKwz154M
FsMNhb8vCJ2TIEdgmAoEJiIf4bmCXF4XZf8nTpHzBYCScoFjQ1TovnU7VEBThkljhhQnUdFQT2FS
BtGHyO9KWpznEjqUMQ+GSOqJ0dNbclU0o3iYuttbbK+4Lsb6vr1vkSdbgzliD/9kyh/gUAuT5QnG
+9xsNn9y7WGnhCR/XMJqxuYxuuQ3NX6b14v0fLzVKU6KZQFatMCWYDQjAcX9TEQwBE9gk5/38l2P
9gRf/j0npBaYclCDy1BW4TnKg0f81nW0SxzYYFBmfZgdWU4iNh0M2b+RhnB7UcAXI7kQ7BkDteOM
KKENm1WPtfNgMNMpsXCGJRQfNi8nnJ5NOEEjSdNSqPSZ9szgas6Gupd6SSX8IlNmy3ZeKh60fddH
ivjgiM5Dq/OWWUOSG53KGkoSDicFq1j3Y1I16yGFM90qO/WyRywsYtTuZ2QxzjAvKjMOViN6e7fd
IJ/lumuaRAEeKGRpmgbuzAPJysZ4psFuCjW1AYHDukP959HR2ltSrSDh5By/AnUjDdii97s0dcdH
IvmnkU4n8K4lZTuSM6odz9aJQHNLhQ3GQAllMzC7lVxkIJ41Y5PIkFC8fEFAmmD9uMeBIh/T2emF
zQaNJDd1ANhzOJTsNxbjfq63lsGyP/iuq9hdyR5+Nialq+spURSF/1hyEELG2koYEyuIM0EHs/DF
u8VYEPlh9V7sFiR9S9iUv0pw8/qx61ESBjnXel4+Rl28Z0N2xMqfq7zN8PNx1owEsl9+o27jR/pQ
Xj9FvKgz981OTCFsWnGXTz5cfIMyqtINVOcK0OsHOlCF5I7Hjym4HdT0AiMPLuErrHdMh1jTKxUg
pZFMWhkp+iClv6r5Wjw3cO/Y+bZAVN+Y1kiSf8ppculoHAAWV6ujgFeqNw4+adiFwnnUGVYPYB3v
k7iAXHn8J1jsTqgCK9Qv5eRav+JbTc+7T86ObkLj5lrAr0Uvy2sevy6WdSbBCpsakRcoYAXMXUrK
UhtuQqIV+dtTXJU2LphFjjbmJ8dxz2Wz+3VPIcy8uWjlLGq6VViL1srr/d6nUBFr3trZw1gnCeJ3
LjU2opuWznlI+g30WsE4c2EtZFkOCm5hE7TNOt0ZjZ1NYtDrgNpAZziGSi1epkOnPUjLG44zsnwp
nH6SZj0t7wZmNE15I/m/S2ls3/jFHeZ1qnF6LhJkkas12nXMXge3xZcQQKd5NHY0O8rB6Kew+1qW
OH7kmw9FaYsT9OawEqbjW+yi84zFx8/evTXKBexCkBMskdpANaSF4ewfpbXkYiXhUXXq5WYmw19+
3Hz99teyAiCLF2ivX8QCZ1EBj37606L++wVvLH+eqZ+sdV7sulpRImK5Ey+bmFrGRudhU+q3N3WC
t9Ip7Urhj8IAm1LtORHdjG0SExRd40YYiDK47UlkG4eP4NH9rOgOoB2pNS3cO/c/2L8BfvTp7Etn
qisrae2IJNGVfSMTvP86DCgd8hTfDin4bcpHEpiUoqS1+WdfcByvEsoO44wiTrxIDxaKXUDFNetd
VRZpnznwJ64Y6csLC1fZPiJ8jghv2Z9DxK55cksoF5drRu03LXyXUYExmq2Rlj7RwM5oyv3LEJOK
n/BHCxwjaT0NRu6UTeQFbWyZuL0HizXWU1J8Clb2ouTGiWrixjvfVg5JZKr0bnJzCB6iU25uOK2s
oj5jquJcuNCdmJYncktLhJbeyu1KcSJ3vpXJVWytgavm69oiJFpouZy/i0uoGPRkFCRGyg3uszxC
1tytVRSXt3Fmu9wHo6wyQc3LfBe23/qT28TU8nVxMB2zUGXQouxO4fV1Ss/dKCHGRIW3gL1LZBiR
4cR0vNDtHk3qBLxy/i8cFUjTkfaBSJXE6eO3yYJGPobfiJvGxZicZPOLwQY4CQKnunYjkClZgZTN
xMh8rwY9FtmnmQoScpe/Lu4h2cpL1tI4cI3DKmt3Eih3P6hIwvl+HeE+Nqjmsdduw/yTxyLAIaUy
d/avQS9h7hvnEXKyjzFqatO3W7cpTyCTrPe8fBQ6xiTaZbQObqvj3IhOE39JsFUpGxDuUjNFqqk1
Kt8gj1roMa2PyY8l4fundPJ1RzTBx2ytNFT4IX4ruUwD4YjOWrj0G/LpPGW3q/Xcif2e3JvTQTl0
xshIO9K0nAW85EUAexqya/bI0HMvs78jL/QcKiaC3lLrVOaSijB0Xeo4qRHC7nJxQFKa/XHCNTWF
k+V2fO7m9+x0rTGPvZv1lkQ0rKnW/hMjv4TMLqB5XFy2u6fsevlWvxo0F/04Z+J15wVKAyXlCX80
YM4A5Zs64zq7E0DNDwLeThTefWkppt4SQ2mNaNsZb2OCQ/xVsCpTYf7aZfXOmK07rsfwM7rf+DIH
iyqZywJ54t/I+l8w3LaXeU/W1grzGTqXwU0cOrSEkYGDItTxIecvbbMucRmfX3izyFhDi+FHW5Qa
Jx1kkXw6Hqhwq1sdL+uzK7fon260goUHxkKMcENIyQK/NPdiHwb7OeaMig1x7nToZF0QPDXnttzp
HN/EmDKrPoBwB1TmNGqODMRmlVLH3O39JPxenS4akW38H9sCK6FaT4jmAKNj4ISiq59U4V2IkXJB
XX/G3GdtC6X+jz/XNF+Us3SFXJbD32481aAYoQfYPIs5FSBQcz0vZZyVCpWHTmIkqckI8SHwJ+4k
RkAztPmotVtxk1jWXlVPQ7gcc42AngCtKUrdtxutj0/sFws9XRBqQJqrJ16/FkkxcfoulCvoQMhO
MxPAw5cU5MCn44poiMGx3UlpF7RxF+l0HvJ06VLY67Gc6SC+81PneeVxU5F8/H0f8zMu9hTbhdI/
+6v8AL4H9yCJTJ4hZz6Q0mbBMUsJlyb0alITZ+LpXJHZzYFx+VERTt+8qZlpzXotPWaazKR/Uc8k
XvfMx33zBZSjJPZhOp4cxlEauNy/q4aF5LhwuvSn/rLd9u4Aodn8kZ1/rvkP23iiNwfD8d+I7oL8
zTV9jGZQAhe7MWQc0SqI9qqnRANWMmBBnv/aVFYiC7pUpolyemF+fkg/U84opEoJ1Obig98wqaxV
ODnjtHtPKDbd3v/2dOjFJ+1j5bdJR+yhhSoEEGyE7qyiFOkylop7UeYsOcD/0wPWBCK199EwCzVW
sVsMi6Pb2uRHTyPrOxvkA3JK6R+qeqHleHY8jfyPrpZgfP7tR51lTvJPs/SrZUE3DdnLsF0BP3PL
enoj3/s6OJzaDd1n+2RBIzQsEibHF5fLYFaslqSYcXhXUsBZzTxJau229qas4Ue5Xok6SdkesF+/
FN5hXZdqWM+6q8CvUBXzUqEbTkRsB+E+s2V129uHsOl7ghD3LVzCO26L7ojNj1FH4ma0eg790nq0
UODuJLh+km7y/Fud+Xr6/pYv2wzEEOxoekY2/dArcmcYG948SyC3iPb5bDeA86O/3KmT1wBtral9
3H0PmPBBHv1ZoExouc/WzlCsy42Om3uJh7tCJGl1PdjxvkIh0LtdviLGorI2gZlge4SwFTrA9N6V
nuLV/Xwn8zeVWoV/NPAwNjiEqbfPG2JO/VNq9UOWLEInzBrOibXx+4Ij51PTFJpC7eWwEx9KAwof
JlTB7LGvM1YrMnM0ZtNYttSuICu5nyI4KXPNRqZM6sK45ekLzlCU4brbhG1G6axYIpKwR4rYmK17
Y9knU7JUtJ/4IS/bJA4XqqLAA3VUSVCiUE7FKgJwqS5NPE9nuAFzVSzEOK+LJOxEmgZXPFAtemJp
KPDe0Zq0hLg/GbCr0xd26BLa/mB9IzqyYQFrQqAjhLHORV+5B2axIp9A0Uq6x9lHia+I0G+D8Iv+
vAo1Q+QhBAAlvrcG/YffAKvCxtOYFnNbVbI2PMMge2pLDgk1ZTMQ9g4gWvNf/GkhujNpXJ2SvR8A
yst23TnEU3s53LlLuUAqzm9tz96lFLKZa2nMAEslMaRgcX7r0pmsBfxTMKIcCLziRhvRdeL0cEW6
MS3vTZ2o3sH9/brTl5c8CohoWBL9vaKnTJlu3f6AO3GIR7HMADDmni0942pOTLop9IMFDCUfG36g
Q0uMHXo1/Yvh4WqGpy4Qs+DOgWGIjNVOrLKn25sk+/OgWHKJgSPG/7FD6Xfwln2do1Zl8Kyk5VDI
AMqS+a41eNgAsBHjXMw2KScijnB6BcRIEHgfLpDlV6ThWE09SCtP8H61mIY3tQH2IgTsMP6gDpY5
Cfnett1cdy2CLxCFu8EHzTA0CsbFb7mJY0cZe6bbJTAtTdZ4JSToa882I9nDv9SD8YrVY4UETNZE
EU3RzO8gfxz4JVCbSsWml0TEqcv8tyI/+Z8bYciN4GrqR2Xxl031iqzG2M18VIqeLkyYJPqnQSWn
mBH3P7pj/8CGoYzvwiSPr22pCxir7nEYtZJjhnq5xCadvp5en65sUPhBWVDHsi9Yy6rqZIxVPA58
JWkHzsGztcDOhq5ezC5Wwxmup0iRgu1iRB6b33Z5QAR2PIuX8bd9A9z02Xt4cEbqSe9xX2dRUk10
7k1xQJCucP3oOs26LtGXYQ41dKP2NZVnyl+6F/wk8bwT/+MApa2Izm8mkJnL2VJm8dTCncWjzHPc
RJ0aHe97yAIFRuK3z34Y1e8C9TDHzyVgGc0a5613TSMaOYju5MvH7Ft32MoN81kSJIxb6+hN4wDV
SFRoj3677FhJD2Qr/5baypGzHkomArnsUzlxVi3r3cUJNydYDZKHEADPs6Q+dvxH2oFYeXshG+sQ
S4V1IPxamA6DxmbUbvZK5algeKQV7/l0Sj8EU/pN/lLBcd9L4lY0GoyeievxqcoCCPjaUUd/WkGw
a+61sLWaNXkx0oeIExfTplm+doxZm+SP88h3PTSjQ39QwLQtzvQ8pP+6nNg2YjYUsvdlchPp5XII
S2LHMZEvveEaupZrDE7GTkWs6EDO9VI7DeVkgJh/kOYv9xmP/xbR6o/oxOQTLOzZmRQ2qCzFVMYe
4exBr1nCpETRPbDgX8i0FCLr+0E20jnGGuzUbI2fTqnLpaMMZiFwf4YIbIVuitJYBxofpCZlClyi
cE/BxofubNWFUwnlPg/aqXLGWXsC14n/yhMqLvxafKkFJ2RM/ofV8JrPdVTxrH9AJkJVXphEQ+G5
tgDo0l+g9awmMzBwPTd7q1M2/8tI+JoijiqHLKJY7Y+kV6rVnqqHMcY/4yQW3M7e73sx0gUrSiQ8
nceV7h2JjdHN9Qw2fwqQZNLXTTbkJ3ZAZUbEEIT2l4C9VQKiq3LJCc4IKr3GqbV7k14HFZ0a4Xkj
83/SE6Csrpe6mn2O9pQby1n9vExVYcqtbWhMIl+NxbqIYxgAzpR/hP0k0bN82HllItgv1RU/PDTL
qKFTPA4CQRzi/YbwXFb0dli5irH6AhQjJWF29tmtSzxIsFHJciXtZeGF5TWgYUf9Oc5hoGSM9NBp
UX3EK8Y3jCYaEsmo9oV/Ug1slJueZ2iuKxEJr6Ex5E7JZ8ITlY6vA2ILdZKUTp58XSm9GuE/dhGZ
wea0W9K4tvn2qFthKO+Seuaq8WuytBpJ+yBe7C+zKXo1rpg+rXjWigWNQUWC/sWGcO3XwVk9yBeH
LOTF6C56OmgVttS6iTkwznLJgYCIVo9j+ClrF6BNGDjvK7HHUJtqxjqc9DuXzakOjpuXdE++s5hN
4nsxCDBRmGZ3UszLkCk91XPZ7757p2s0ZkGuhUWNrHPFeJJWpWbSnmG54JwoEVRSmbZlbtSwr8q6
LYGv7UVn1jWIlaKzsR4C6RyPPkGPkza3yuiQw9mkgflWTz9bIP/QrQyRI641+kDKVvQSTjUK8Blg
urAg1g0lnHB8W+qsr4VQek3qyGuixexCikVWbsG5rQu1p8TLms57VAvGuZbOgnCULmxRI/aWqpY4
ELViu6TXLp24Ag9uW4KlNibhjxMgkIzBtIdQOUGy/UEmhKjF6IBvxtKHwIdOqnSvFouYOxnPi6Ig
P5N7gUyVCyx8SlUnnzxCVtQUwiYn1GMzrHnTpbCC2WCUDGsp6f2BZJUdNeFckKiJyERrfYwtGJ52
63IU+Ou5A/hha6ypP0lzgLn3NbVKQxeR1MN/OdqaehRbL7T9i+TzZtbvwM3EJaT6H0FMsZe+YlSn
ZqRhL0Iz+pJ8OccIHZ/jZ2SJPJtrtZ7oMX19G+YOFGSOvTqwp2TFLlHi+wNiFvixPKzYm4ab6tGP
PEO4dEtMxsYlG8wLX5S9WHW3YPSVUzoboYGDnOt/HKALDtDEApuVVkrMIN+VNI8v1EScvsIcVCie
7XSjSH+MEDTq/JrJpSShA5EJsydqU8b5i+3ljtgF55qPNyQ9akSNcs1k85I9PiyzuB9TPXbsATcD
li6T+H6Aq6KLL3A6uG0ODspPtBKIns0K78G/RZPd6VKfOapouxp/gPxrojV+Q7ns3d6gLU5ODDnW
+hdHlvuQ4NDXHNS004r8m0KOdmeHTjtO5ty4ES9YVQac/CcKMQaTgpzxbvtradNoq8lOntZlE4Uv
HTlqx5Fridu77FkY8cugmtY0mdlxg6R5YUZEeAhNeLGpl6GWHZSS/eT2Ch0xb/TfthyFiboL4K90
F74R7cl1xIoG15UeY8g48JqQOsaBUBMbh4BYvP9UtoopIhWb/emeYieJCHL0biAXlQRznqZeOj41
2GdBp3+43P5nC1XEqn7r5AXqMhUnwwbYjOGF6nAwGZWmm5R8c6DRpZ3ZiFEtDNXwCQMD/dblTkRo
waJzEtON9w9MuxcKqD5Mg13NPpICiQB5A7M1LfY+ko0dF0nMzG+GCzrS7qIb3H3Lw9umlepkDrgr
FF2Wwac4Tf9hzos3mtZ+NkvMRmFoUtPcSXoT4DzeYpWrXzaZA+hD/V4bVyO4dejkq/nWSWG5tRyc
cUoOytyYZ/UJ1Kh22bOfuB72MWXa8wLfBs3u62s1bT6kEBNKUGxbwszVaG7FuutQnTPRHzEh4t3s
bSBf+4wrItJDF2j5F5fK3kMhJjJG4ROsJEXzFTDs4cZs5pIu8xjNpDep10x86mO9e35MDnTfUTLo
kJZEZDxYhKkdoWce8rEyyBNfhjVEw7xy0YmSbEoObXV+bv47tRyjFFXjeFnzLJungv8k+3XMsJTs
HOidegSAVXuAigBRAuvbxTf/BIzAfZAClaiMeq66+4UNPkGic2vQqqQm53lt/RYJt4SFCzugCvFj
z97dZWLh8H5XutMLOtwyrMkhGIv9P7G5uVCRqSbm/KuCgZOg3k3JJTQ8o4qLA3budBQJMmV3LfAy
rM8XVEBPnfb1dPwbwSeXMuRLOGTNdj3f1hDPZLGvf+djKFKA2hO9SWL0GMTb5EvksP3X+4XNp1ML
y+LReetgOw3r27KCWjjnX9vHhPP/I1FN00HiwIMNjrUwxWxdSVy0d19X7H8DbQbG34eot0frbDky
ul9vDDH7TIXf/xvBkPFRl5eCHxyRafPkN9LDfpa9yT7GA7rsTUmGwFi/WgdleLu6hiGnIyeiTk7B
xOXddClfCad7/53cajYn8TfeYHNhMvubBBHcnN/phjtgkShy4EGMnpqMjYqTQJW97V0fyZvyMFW4
w0AX7aeRyzRwYCwfijXkwgDJuHNZkzjWils5blIo3OXoKUz+6M0NaxKjs0nfW0w/pOJS9z3DZD59
eZsz4f8BI674CbAcMTBaQBUtfK5a012x0oXRfrwLha5fQAO3QIDy1io+n9zryqfYMQex8Vt5cayV
zTJlRmn25Cn0CHhJ2UNn/zTrby5BEtZTAYtEUMnZ34HPdsZWYfLPLDcCPKaSrNSX+qFC+Rn/mFif
BGxbcqwfz4eHRpfbkHsEi+oEQp55KqaKeJyP1CbNQp0RtcYA6t2ntURy/ToNmAmoiUxbxqJ5Xx6i
PIGbcNTur9wU/wGrP3JytvrVZD5gU1TLEX0GFxQlNoxwmGm16sBm74acflgHj8k7n7JOXHNVXL9j
hc+jTWS7dtEiZupkCfWWi4K1JBgqLea7ihj6rwNXAkOGccF0+3tlV4ntd4Beab8kbyslgcoPLWOh
MAjBdoHEQ6qF+mwgxgeyIU9WJDhhXuXsvaSKme4lfia2KrPGe/CIJnWZCxzYcxPKue85EI7nbGb2
bFMxIFPHv6RTQB/qGjTdB5ivBJQLEUmIeNfmuBKy7CNalwlTi4OUFStSNl1lNPPmtE9b6REDvaDI
hWwTyfVbKCujrWIKnNP1OZcx7v+Bj7zrjyLoKFmlSQndDfTuEjHe2BhB8tEAV4U2M3QXd7awbDWO
LWvFS0aZt95f91vzXN5OX0ulfeXMxH+55vMfvkxs8G5SKWCCPtFlUpSrF59gtIwLHzmiWEUq8eFG
WO8QzLY9BDja+BklFaQH7Js4L3VjzNrFV/tPLisYbn1KQ58H/eOjVCpjWkn7w8y2McH2tcSAJBiY
jWqbfXKuO1ae90YFAQS27M8jsaSvWKe8W8uz7ldddGhTC4sbscj/K0/yDLldBNPxixBtjzTzqtt8
3FsAjT57Zqchwre9ZMQl1KIop6Wix6f2SPmqz7QOfRU5crwRJOAzqAWElt/S9tuBO/s6JfChMWdf
v+gnSUsabAmKh2HNlL5p8wBiHeXqsgeAZud4xJ0/2h+ODuKNE3alhM7AnHEwN1G7E/zRTPbJG+D4
zlDVUXjpxbZllO5Yrf2F6ZVAYsUzMTnldZFO9l4GU0m8qj+2lfwOEH1f7P53Rkc+pkzzOE05ZdFS
o2M/lLhXDr/KaAOv4POgCUnULWIDwaJHEYc5UjKeVgI+bLmWcRg37iqDC9f71JewmNDQBdrlLNNL
DuEKrFg2ZddqfKxvDOEzSjdo2s5ja7prpbob9+3D3gKXubKGRNYsKqivaiwAxtm0QNVrU6h89zIQ
C0Yc+as0ZgXFEyOgpgCsJ9fwNrGq0JGXJvXvYK7Wm1FPaxwfnBDjeOnzMlL61ucPcKSIybQOm1bm
3c1qtVoB7UeXtOQRfrAiXHYEaaIO8xiHbgi+ynWhI+P7Jag/v3B+V/0DTw0u2nogSN/smFvFa0JX
xxe6plYjz/aGoEzgzo1/IKRv6RzR1CyIxWVW9995xVbN1rMQdGDUgJGZZBgYus9gcMk4VvVgUHZl
b1rbvipXBNTRkE2/xtmm2/dAAAOK7ePrAtu6ni6Pb5seJM53HV6sxZZuI1cjvtcCrzG2L+vZ6nnx
dpx7RhnOpXh99duCE4kNbsgQ6/EUcp9okdjml4DhwsYJE3xp/+ddhfWJfmdcw+/PcYz7yNZSWpXr
qekNNrlvY0nw0S19MMCcZcgMiilLXg3qT/lIGOC9p3tOXTSfeYkB394/8+JBZrvt3FC3O+VwvmG9
ySJN9pTCsZIpsSXTIEANv2f01arniZVrMqIsDaMRz2BlICyovBKNUgLCXYG/YPG6eBj7MNmg5TJN
GaTHXGTTBMZvMp4jB28pQmDc6MGfMi9pbxO2KY+w4wpHrYGHAnndOsYC4Ovb3qVlkg72PdddOumo
wtI3+F9io6Y0eu4ynRrv+cqVGBkBy+oIfJpFzOM5cetG7tJqn0hd+01tY6Zklx7wUP0RrE1SJJ46
kOu4P3QUUe2Qep1TSBtvARYogwNcC58Zf3sT8rd5jXZ4FUxwzPQpeh79b1xwBC7GkEwgceIZ23nm
BnErJDYFBFUBdZN3iZKgBhd6JRvyHXhecsWjUkKbO/3vpGO1KH55Sm7b+C650P+NgVmxwZs1RuOe
jmfSLy09O4L4GpjxjFN0dtMjR2frwSfVnjwCV0e41nU966sY28jJpW2RC9sgPXJ6Y8ByBR7gqFeU
NxfQJnaCh6am7dYmglAypd+nEhkR/yRV7xaig7r+/O2vE3NBRE+HUkEGz4OKQXlGaJS9xWqCnY7m
lg1lx0WmNOQDj2YG92x1j2tPeFAgdGPqwNAX8OQ7pVEa4MeG8ihsY8M/N/VXzM+nK9PTH944oFRv
KmlZG3tcbBMR0T9THl60M4xJBV8rGHAWnc/+c/PC725meciuY0w3xm5zgJ+NI4o2npZn9pVCdBbS
XF2XF0K4JNPlkSVzyUbIej5RWcICdQDB45n7Di5PCAoQZHhKHhfCBM4iC5IjD+fD2JlGF4iM98bf
hF2iY9GOb6g/BQPsT8vPYk08tfDdtFwVuh4tg3B27jGfE25/73HaGSWkCVyjDJP6aO2m6G4fGAFh
jCedDI6Ir30tiD0P5TXyVL9c0wndAtB/UzNxAuk/dYVkEbg+Qthdg4ieUmEFgqoRR6RXGmHvwfBX
Aj1h1/5egY2POfDD9IK1xJKDW+uopDvW6pbqMUjVK4XB4f2q3UkUiXhWIZ7XiA/WiM3cNYEIcts7
jyldwLBU4uAEPNGmbam7ArqCS53KJRvDT0O6Lvid8f1H9PUjpb6tr7dx+96s1DJJbOxf2hh1nNZW
YcY/kGXbPuMK+QiZ/HoEH32mlctSzstSeXbE0Q21Qz3t6FA2ADjuENqGJ+q34VsWg8ACRslMtMlO
msyXFZkqTQSogH2JjMrQT2WaOV9ajN7KJUgkRfzOD5N8tQ+9xTOuturpy+Cvg9d1UBIDmDZI6W2U
3Z868iaz65cQ4GtY4flB1dbd5vC5Zf1WnOE/nlQRGLbSHrpiDAJdHTD36J9GzfbzjfGtKqGIWSZK
7ep/MgQRW9sTFo2cQl1hWekgwPVX1naUBZH767O/9MMbZ9aJjDRERFf/4TOyGiJioxH1hIre+ebD
/MIs8Dryrpw54+MYkP6o5LG18R/3V2vr94zOb9i26Yp26nuvG3sUCMhebb4zUb2xSCUxzHKUpYjR
ekHZ/MpJKq98KKriqHT7ASLaRWOjrwK5NKu2PH7cFU167lC/JETxlzO85GUBBF2Frbz0sGHFP6qr
5lN005aEM4lyJLe2IHLYa+Yu/zaWZl97Fz9PkDr49VlmTvRmXq1Ru8TtBBuHo+8oyr7LccDF9NlE
Gr7t9iwlQLYhZydcravYqy84u3spmVRcgDY74MUbY3VsolI51mcJ7Pt9/kjZjxqTKoIYq9Cw+ecl
TvFFRYlQe5v+/ofqbU5ANxIuta3cucmOwH/FMsiuTgb6ud1Bjj2Ac4eZ2Y1TypoYSNnpFoU+xKDG
qwU7lsC3vg+WjjtrbqlVPaycdpnd745g4SJwiS+R9+nFCUCwiEyifQ8uJxxiv+JmU3zJoAUhUrFA
zgCyk98cBZJp+Kd/PM1EJN/MRj2h1NTIE52TkIpSLAuyXWqS1ed/bBYOQ7cu0S67Fq1U57Tyw1Jg
W4tmiUPN/MdRYFLMXReZOgQ0PcQ+uVifRCIrXs885QYOVVDeTXJ+mbMqGyyPliXZmfLWH7Lw3K8L
d7yMQHIIMSE66um7ZQaM5EFOrJRURmXQwgd7FA1EeAg1ydCGMvWMUbJ/Goa4sPlzo/EXGOTxWrSY
g39O+SsWeanShyWbAuRmm2SUnTcuSkFMh6V7wRRnPZC4pH85/dhN7sXdM7mp1qquzmX9IlCvw4UP
zUIl5/PHQBGmsyJERbN9lxNgArVpGOuZf7wYvbTED/t77yQUMzqVqI8s1tX2GOMD2p12ANyX2F19
UctyQxqpNw84y/zY4/SAes6tvUeSTzNB9dOc7uQqv6xIYcHtZqydqw2SGUZyAUYwQ21s21KDE7Al
jd7HT15XjUf+dpzNEqeqkmk/xWrAIngr9/M/2mougoYF+djWeyQIUlzCB2E/7TGDw2GUl4A4QE3p
XdLvhKEkzX1WLOi5XqaD+fiMU4OGPIBFUuTB9r6T22mWbiN9L/hvk6jAW+JpOr2FVUfj01ZWJbOb
TcEjAEruBUDk3wFQ28p1SCju0tFgmSvTmc7Gjk+A7yF/CRiFmXoZ5xk+updS/RO3Rgni1F9vU95+
TowY2uo39vDlW9mnjm3Yj4gY19kcrg29U5wDRShmmIgekEZU9Uqx/8RHU7VfYYw8FHlz97bCyfco
jG+Qk0YLbFjtokKCn9/IWufnXQ4p/JZcK0t9ZbaZGUEZNY25tDgrdsV4GFHgjgoMUvOeqlCfvKiY
ZH+kWvjn6/ZIjSb0LH8VPHJCyOhBVfaT9/Y8DRzn1oO2C/NhxvTr6AnrCKQO6q/IoYHgR0L4hnkH
/6rMy6ZEwaBH9afnejPhLr9jSP3XLwVO8O5HJPqXCgqjsewuJodQK/mtCmnKrpMC/1CgkrsuyM7u
LLMWnwXkDvNL7arzy2Wi4fClrZAD+4EIzBI95EVDkyBeBHr9aS8r/w3ZMs67KzAds3hMYCRS+wNe
qEHGSl75nk/2vq+jCwhE/uRFYqGunvXkRJHpeVUMzWEgJIA5+b9nhc6UFG+VMkdBUPHgjPQbiMfa
XuPfs16Pau2R7TxyrOi7UGP8Wvm1hXZW4yr07lJEexP14SAANl7yj7kDnP9BxEpySzMuL/P4enrC
Q6TDnQPjzWWKPD1q4ehD79/Tm2m1KGToKyWbyMIsMr00YIBJ2lHYof4OnFlv7bF0CBcXExrxpm1Q
6JtRUlqKKH0ZY6qqMF0BH5PparDZOYdt1RISgmpnhfZ1Zypd6uamGBSXPV3gt0rDngK+6GxkHM4I
Ob6q4Dya/qe4QGHhEzBmXM/6u4QJNPoSH9FI5KcRlnI0mgRHtZvns9fRjxzTXWoh8JJ+DiSJ/LVR
JWxYit761TcBe4HQI30p9ML9RlmXEj97URnEN7OaQs6m3J6Vp2o65JtJcSHh/KYEpo/ZGavyAwLa
2/PkPLpT6sDNc0T+sfd6DVo0HetixWD5XjirE43dcNnHkFdJ31uh+Bh/HtAqzDnsXOWZSE9SbcGl
LKbcXsbgwZqJjB9DVa0/17D7fOx8di3K+8eZJYZv1BPV0upWWxUdW37XEa0lcKDWdL82suUwkQ8A
sKA8Iy6gBk/R6QP4utpd1p/Cu7M92xfEL3Zfyh91x5RdzucbUNnTUlbb+YgvlzogUWh7xeSoV6LY
Kjz0t0DmjiLWZF+IH5HlcuQcaAyMEkWa6hextxoxLdjNEzU3qzz7LS3kRkWwZIuWrUfnD/M+oRnP
LNu7nKeEq0EuBq/+FpHjdjhbIYhp+QoplF3ZM0GQ6mkys+WSnZ4Pift9EnhmDhYFNDkLVAQL0TbW
Yikih4zTDgcXpzunUfyM2AVt/jjwkOBUZfpAm7D9iOQlMpCb1GgAaRL5/0oJdozMFL2EtIItCpda
cYMwu+WRT+J8ZjFOT08+TCygXYMfFTa8CqvDOynZOO4pQF4k9QyEk0X0pNNS2pge/xm9q/wgsH5k
CVFXsaiawPhfpTqjCjsnvPzoAUWkDpzz/wD15YDpFKnNcUfnLJEH8Dw7Pa2xlux8qFLnXrG8O6Ol
2kxHpNV86jjfGZtgFEKjkYwRp31Zj3KuP52dxNe445T50nHyhVoX+SMdcSkb2bebnfjfmqZbC+0G
dmjz3+o5gvEp+jVmRKosKtJ9I7ktRdTQ12bHuErZI2V3JjSJs61S1BjJIFT+ZDBTZGkF6Cxn1upO
2WRb0lxGWUpUzpwGmgmLku2h6DcTLN/vyzyTaHyMLsAGQjQU3I6ScM14cc+p87oDDHaB59ZC38Vw
gkQpOSbH3tfbCUgXGklaXFDB77NkONFZK0I+PwdU+S6xCZKlmh3Fhr2fgjlriKMXC42aNF71XTee
xGfZUS0PTYtTfR44tPYdmKDU25Df5oefCpWDTwuIQkkULZb9FN+BTV0U45x78o8TK//vPUq2f9W4
aZHyQxa59mNq3m5J3UXe+K2dG3XOZ1HsJXNyIVxX9+/bw2eVOjLBSNZoDSYQYvPjhe74ATletZoc
KNkQpPq3fpZB+LnzxvZZIJE8REbtwiFMgPxpVARtIs9VSMLqnGkPuZ6PyEDzTA0t7OBxNb8upbKg
FC9YUESbqt1m+aSEY4hDSU3hLxaWNp+Na+bK++sAfHrUkpTwzgI/kYqqyfeIVksJzQ0ZnNgay6zS
8kxuIawwOc7ywjhkzbbwlpweOjFZelliDMH+HX+2pcc2n6Z9ko8Uq+aHz533wbsa8Itk7Qr1iDHl
fP2agKtQBrLk5LUOIDd5jWZautXZ12poszSVaOzCFKNIBV+KBYVmG1jEXQ6/nAnVLguncFl9Fjpa
OxdXeWJcY0I+3Mo6M62Vr7zsZxQHcA7SfRb/0hWQxAx4szp6e0hWkAT3CaEB6KmvLRa6D039tC/3
1s4IZB3BmaBnAX7eMnMCxQkRnmUZH+6w8JGg3siosso/ABX6IFxWae8GRbe5XiyhV+o5ShGuR/GV
xSkrCKQQpm1KckV+I8XI5lM8JF72qIdKGel/TMuOSGsp0fOxnqBvN6v0V7j3pNy8LA0f03iZ0n8Y
FQQf0FRU1/QTItscSa8BTjpIpdlUmj5/VaQ3uHb2+qc0fm+IlXoofwl1vON7VatD3iv80Sy4oX7I
fnRIg96E3EkPeTWclRhKt5oIFlYc+07p+fsaWvTgTnDvSxACpKmjTvz85g32YDMUCKxEU/eMgx7t
pAi4aZtVbnP1O1ELQ0C+ANDcooTR24uuz2UW1X6U/BEhW5bcgtXOHVFSDrRNOXkbLEwazXtW4Rx3
UqygnhBU27M5BxS6GpBUpT9zzPOw1R4ynITKtXLepK1YuikGQ8O3eiSpugojrHzEdx4ZFkCDlUFX
j2CMgZ/SifeqWXUxipeFaqv7xgDnTALwMce5If5iLIlmnx5NfpnmP6bCIyNx2QeF7ND4q+IsteZ3
r/ADF5GqxcSXhR5QBJKxniQOFO8yXvffc/Da2LL66RBuQKxnrqYbKZu55Ob6DZuMFjBsWtRarQaG
w+S9kRd1vvicoajSeFa+e+VHtdAMzi4FBbATmFhS+gEL+dJX4R5AGK+1Ev8jWzlfAG9ju7h6umO2
ywOlucWuBM5V6ZCqJ8hJ+VG2rJB2CpqrGF9N0hhQ7vJ2rNIy41L/Nprs/k6pNs8p79f31si3T28r
GkXCeFOSMi8PgrEwUyr0G2Cvgk3houxnl+c6CmqhoVKKsVuD3Ft3cRh8zj3tT0P/KYvovtDpe2+T
P5cYBIszqj+YQYEUoYTakIt872PVsdfLmlR29izaiHlZ43dXlPdThzpQUwN9xd2Eod+q0TMj0osK
JjAaETagheNmgu+pDK009Lg9GBGWhnqCSjnmN5KLhvod4WzyHR2c1wtJULdEyF9RZs36Q6XmNKEl
4jfc4L1B+wVeqQ1N2aObosj7LlzsSjqSXvlrsa+yRvLX1mUT9otll7WRU2lZmmHWrWyGKIbQ9AhB
YccYxoWKYza1ZZCO5es183YjFdt1Fg2OjDqxnE9CB1DNH6BBMiuzu0W7g/JuDtWkmNr11BcVhfp5
WddOGEtOvYHHoz/9V8QVKBNqwe1UZExqi5KSqg6pM4aGhbnpRCkXhzB5pbsb2hEDgQL4VjL9I4iW
vEOCaEjUciIBvAQMdeQP6W39RvBIwlftXuUXYiyfducH8lQSG3JiDzf2irlafeeQNI8vqd5diYZs
fZg1Vb0H/6cw20wxObpZ5g64JWDjlW/gesdVhDtBpu9LJm6HdXS6n+CySABisypUDMzGTo/eUXzX
Q2y5v5FujkgMdD3/UPhHDDaJVSTEc07fmQ9ji5HWT9ElhB7S7kAsu2CX+/uWc+4iQ5JnnyHZoWjc
poI893gEFBLXyg8r27peGb9E3atseVRcOnZGNUOyFCSrbFWRfi0SYTnjSAWApDj5x7XEJR8Ffuxw
pp9VmDpmehr4ImSrG10AqLgPjmjYr60VOHA16luWH6KBR+QCAqCiEjWzupMjaCa3DPuOT8KMMBAo
2RNXbutyVy5xPxnjkSLL/XKSvepZDqbt3pVuMOvzCjrcbRhQJpQb3E3y4shzAnSAVejrq09FvIg5
v6o52MzKiJlnwGk8K8xqkqExXzGqX8qKbTm3o0WaxO1MJkbCPJvsRiXUQOLPc6vI3rekZ7lMBCxK
Y8Ooo5tNeft7wAUOMiP+I5pXOEVvq3uY0yk9u0JXmkZPjqHbVj8AzNe0ft4on6BlARJvm5vPKyTj
UKdJnlyqEIEzptH3FNsETF6aZ6E16lO/yIk2p5EIqnhvdBZxDFMkOMTPgnNTJ8Nt+wudunQVCiAg
JUtbXvGBDXqnvMHqKwKYHcy8su1p1X2GfH1vABGrRO8K1cUmuybi9iSbf88E1R63Pc0GeD6yUM0Z
uPe/7pekI4SWxzSAfF1q5ZYrwk5pSs2P6kl7hqsqaWeB+Mcpsp31QPPmJ750SHSege26DssTlzlh
CY9PxGioXC51NblAP5vAWyj4/uPGzQ9lf/l+NQ2Dd/5Ldac8rgn393UDZkq0IPGZbIj2PzpUeuBJ
RBl1IKpaBK4q3Mh8NMl9wKLzEJFCi4mUYkeynAV5fVUTNOE8cvcBlmIT85su+JT/juqDbq/grg6h
nB/fJkEs8uY+xmt4ayi4VoZkT/c9BoGR+JjC3EDBHuWQkRwOUsB6t08IQxhAqhlANHAMckugqYMn
qvvBtpDYYeE9n2U4hsdmEfVWt1sNouysuce/Lb+hKfgPUKLcTn8JHs9IOmXvJmqbscDIke21Lohy
Toh87TqaePlqV5CcGFiCmoRnif2ExenijHDa5Q+eloO0C3dWc3gvPB70GfScEO8+HXbuGsAZSBnw
kkFwP58Td1unpADcH7idt/jEmir8fcltW04sD5hPScI9p/MPQ7sbcpluqQBiPTIdsBswLeZR6EtF
eCRZlNVDBD/RaOuNwFtyCEnClD2CUGfDsAR6wqcvdvyP7OgucSQjKZmlxmSkfqKmgPF3Vvh+PA0N
NiPTb0UN9YhxTYhs79Pg2ou/3OaKUZDgLYDyu4bNNXg+AHqrSpM2I4hja5KeOiSioS1NnxxnHRxc
RF4ZJCxSRymJL64ISRp+T2KKnvhQruIF+PSNwfoflmyDQGoJ8CJIL5zFj1nCt4snUw/v6USC2kJf
OvY0J+gS8Bvxnz+QdiIE6MLS00b09OityaCjmpDcAQllC8sWcfKFOGCetfjsDDDe2wM2fv0GLE3M
0tpCsddJ4sb8rf0UKwQDCvslQoYw1uPE/FgUwmObur7WTfG6vpH5sSZ21BkP5vbb6CVZIjLTPoAg
x75Oj9O24bLN2yBIAW//3MBnvuMJbeLsj92g/RK9qnZHwc/Uow9ABf/DHzZEaiXw5eKZnXyfKd4e
sstNxMAxLF8Lhqf6FFBfVV9xYuqEHBlP70Huuzlcokzzl7vRgtKoc+y//kvnu51TxrV1oySqDKYL
mJqrUAOz2bXbUt4lQieCXj7uFugjfttOM+IRVKfVHee/4spOpOvbUpG5UbfrbZUE398pMRDPJvbj
NoBolySDrp5pPR2PxpjtNfqMEaRvrg8tmv7v8Ic/aN5sCVEvAcb9fu/iSBFBjtLSWv8ngLC3YJQU
1wfoLUw8mD+EN8r9/ewr0vZ0Z31fEwOB6tfqU6efADJrnTGLu6S50QC3QLM2sT8MtBGOFI3YjHlR
ZX4ylXp6zULQgHuGRlqdCQltetcRRN4qffV4D28HDRYyEi4B0ehYe8C930cAQorvgfcoPRZ3NC2w
FX5f8yJrOX2bwxh7clSwFONrsH/wvdBIkqfCmkg9HxoAPyVVuKtc9Tk2Hh+z/WqEP5/R8jl+dleP
OUoBtaMABqO4/RMYHoGXA4hs250Vd+u/5tI39riDJg/KfBrLihuTS+Ye+bFvOJSFxDnoenTbKBZg
0kUayXHjmNu9NNgkHNazOAXdTZwQkpCB0AY3IqmmQV5/JeTFLvvanfR4PP91J2KOCmS9XsyFkoa5
Lyv8sZuqZBTqEewEci35dcJgwAwaq3XSKzY/u7QV2toYIIVzWtyR+3wdp2zQWEo+UF/W07anMFvT
Wkk7R4sjn/G3VrWCOV8eJref7dlQc0s/WwKt8t3WCAnivOzjYA+4Ql1PhPT3j5h7eUYywXxLjl+v
DFhl7gvE8xI4sWHB6S7z7kv8/2ezNhAlh3eCbH9yBHP1a7lwIMeqj269XDwvmxgNocco1l8pG/RZ
FXI8nZQSIrfbZZ9n6K2Laz6Am8pBCewbVW9HToIklx7VXOpvtbI2jk9mrxddFOmcTsEjkbtPbcJM
YMNvhouhcbZ4ADcq2owEmXrI2k9FAPtAOPuyQHixWKUXMKe/LdYw4z0e3rv3aLyA0v7I502n3wg9
R/97eYCcoW+EhSWiDXI9Phx2jtsY4/64sVWnT102ykx2ZuOXSMJPhM4ArINAnNjTczTZHJWG2qic
Yx9wmU+RS4YcNJeXoikYIvs0hwhq+0Kw5ceKzHQXPP9NdkZ3r8f6TUnpNyQRV6qxG7Iobs5QbmjH
XxTcT6Ed5fbpH3ljpmKuT9tL5p5AcWZhTPqBIw6wZEwwJtZM21wQ2/DJqBusSzsSdFnF1knLvqDB
nURFkipo6ark4N0fVfeE3jGCwL/yXPImcq4bRFTzCjHd2F0LEjg4eFqckm1ntMIFrTN2vDMMxoh8
XHr3z8tHEY1hTW4ffXDbF9QkzkOFQwbSbPEl6QQ7UAXKbqd9UNxg+N/vJMHE1LmkNZ3aIk+Bx4jY
oWoV2HgF8Zp8/+YaXhTFjLiwGDmxAr07dnVf8foTPizvXXNPaIu+n5lzIpnQw0mmVtRBpTmcD4E5
1h4SgWgSY+lbAl/8Y55QtxPp6yYCpwCTX0NROzHjxnV9OZOWRX3MOzW0hTReROZ7NFilyPm/DdmA
6J431DNJGINgX5NLojhlHVgo6FXpD0QP+qRT/1gTqOwsyDtIEoR65qm0JOC0wjEcwxVUA/q9WRFV
YZ1JMiciDke8k6eNoKosDyw0qF11ApuNc4zxSaQOFEyQrr/CMqx/u0N/3RsNGDklVObeVw0FJwlX
JEysifQExwd232yX0aYU6sjmZh1me8AMSswf4VzII9IySF34mwTzekCmfyPfNm5li+niVCVdnO5C
DfliLo0be5ylTctpHDvkpi0iCzw7VTjDOXDRwezdf+56cQfswNkFNJ67UXQYN+7hF7fCiLdH+toG
EEyKUI36AIbvu13irT7rGvG6l9SCztBNdg8coCoAj8fwmRdZW+34EOklBtNoP0d2W5BLdcUajP1Z
t2TfZA8kSn4O+7Vt5m7x+c++h5WpVGoDrqZEUH1Ax3Jx/qYijxly6lo0qUU76KghA9RsoytPW0I1
zLQxbSYMWsuWBOZkx5Bo6YaMR/0iiV0vAizJWuC2fkUWlE1vNYFfYnsywk8b/e0B7DNXVnMjtdZf
jAc9Ur9lsY4DovY3H3rQFcANbPaRQoof5h4Av47Ckme0KG4lCEwAG75HgU4ZhbdR745/311zhcna
sQ5NjDHSwmO5Cw7/7AR8XoDZFt16NiF3dVZ6BVOjg6PYcYpEO2Mui/KrKNjG2W8MHr9GIzMMcM1x
h3iVT4ITKBOL5Tr6riGhgwtrIFLSRSndTk+pvRbRE0fbBqH6gM11TNi0BIboMvb5OUi+KcIUAbSU
AgZRPBV28dJT3qOdV10nNAZrz0PTr5HlLneqfuJ4owZ3YQy6r8g84xNPhqqQJzzHKEcgDELzaREy
VK+fZxPPeVvylFaYPoo+l63A+NGcP0/AdflwaJjEMQdAnPzs/x0rGDGCctGMma4S/PUKEfRT1u7+
utEetJs7q90FOoPzkA3OSbn3paAZk3DjSW8XOUIdNeSqFrfTwFUSn3FIMqjYrJTw7UE3bKhfmgZu
xx0hyy3IjQGh5ICz0mxd+hQKtRNwgLxK2fE+fMd4KSTnWrBaKT/kKg6Sk6W9xqcFeBB4VwXlCNG0
ihMa/eTCD5wDRkYrZb52by7T49FeIMQdR+FaRoh1cAgTNA/P1wpIDE9xSZZ+MKtMGB+XVVHfNsr7
G05D9JSS2FnmvVGSoHMKdh1j1EBZ/JeUq/Q2NFGrE6GuZJg/W3yENhjmJWyoNkumOBr/BfUZs0XQ
Ou2qVelEPABP/U4fKEit4wOpn9gaFT+j4i3NQ+YiBA0mQtfGH6A3ijZzY7IM932vG9SDgMez0JtG
DXCFrVjyuFqPHW9kIOXNh/7bYBldyzH3QD04nJ4KH5Ae/7kO3Cgq45Vc2xKPUWTRVGthjNqgK7MA
jQVbIbKIpj8xmhrBdGwxGe9lZnDt4++yRBeJZbMvWDQufDitKGVfK6bds/IOCGnJPfuHTTD97Z3d
aEuGYRqvSpTDue3xm6S6S0YsWfvnH2cnI7RPQ4GCXyln9x9fwcuhOfoixyLZTvFFIFCtJ6DNkcrd
ThG0lU1hllopZI/nCm2kxrDV2gd8tdGkD2RDvCyLMaFeTsNppfNgJG3jK30/xgnACAjE4CxfEtFw
8FzCE0f9GC3g5n3FnRg3Mn3VSDuf8KSBOrWpjlItvLMq3NhcvAi7yNdV+UXuNHXLSaD3r4FL6TLI
ZG0LiB9tt+FjR81kq+nPYtYhM+VaJGjvz5UYW5JyN+HGsXIRmKcE181Zui7agGGhJP5Yg2rkPjJF
PjOxBeaARFeqvoLw/5O1jnYOrt+PBPlFeT1N1ikI3Xwn/AxhM/Ey/WOlf9IbADkYllIrOjOPAMgO
70WtaeIhoFaonFkBpkme3koAi3ibi+kzq8ErIMyqThDlEM+SWPDNimTCdDANKc6Jwmb8PNanp5f0
S+msWPIsPW5Pe0T2//Bhce4mdtJvrKSEwMHvfuiu890AoCWCPgjIQcGxrJ3nSfr2op4U4DCy8AgI
Um+3X1WIGxEbfpYRYMJ+ZYF1edhfvQ+U/CIyhFQkEisuM4NAeUJzwwW/fBH1cZwRFnMg0Ljkf6Nu
gpYQXvxywRJdHZJVeDRKF14lbZXXRc6D4n8zAGRGDLvsXeFQXnqXims2VVQa7dADTmjTvL46fZ1O
2W79McLSw78O5PN0xB8cxrgzUL8dKDTcIIsGOLXJGF1eCLWScRZtsNRzE2LrtAH3W2zWwIQu6jKb
1PfQc81ttG671t65I9WqhIEZURotHSgzcTF4EhAlWzmPxYhQJm5nlv+E2WYfCtsZS2lLBrZVP7+C
D9CpYY2o9XBGED0tONLxWus3lnOjTBCHPb3rI4XChLXrvkxkP1GwF5Zq5N3sLjVoc5mwAY2ExmlS
69fk1b4iFy9Wh/hW2PTXwycSen0HAMCd5gwtV6JjrfS+N8Mtmk5eeoE7soECGD2bnggX+U7uBENr
9KxJeO1m83VGOR2zlzqsJGX9Z6/zsVB/bwEBvQ3ZQia499WBnd8Od8vBAI/ZjabYPVw5V77cXiCx
jqSxjExuAnwwhWRp8VLlWhU6v/cf1udhNu/L69yMKsj/4sxRQ0rEDlVmzyRsLBVc74VXIBjl4RpC
KyXal8PpSziHIInb5jwiO3bqdD/b2Htyr5ielaSVnhCZacuzaQOk64hfRqPkUiNNRUk0TOAa5iKA
toTr4QQ40xnQkaMWKFGTuIquNbYMZQR3kj3TUC27vT6vEUVL0aO5uISIq+vESpPhMQt4AxcZXzip
o75wHNx8K3Pibg0Z95maWxlR77xyIztqbV3kXNzKH1GaWG1d240odr785dE3CWVoaHMBAYGUc+os
K8112cqgslLxgDEOR8fEV4RVgKD32LF3QYuAAQ5VCU9IMsGnpLOPbObSlIEvVicEyk+VV0fNVQnC
PyOk21k03li3RzXj4hXTDVLEfM0J1jiLOdYKakzkLy5dSN1Xc8b4JX2uINbra7xIByk4ww0VgzUY
R9hBao2Fg5RYDQxjRrnRhpkCfYpCXvtwCEAe3aX/zklzJMDUxYGpL9/Y/6vWtpf91AgAFOEryfAH
POYPZIgiSq11gw70X2hoRit3LWGevo1fOrdc15iaVno+WYOqh9COQ65gsKMCNb4VLBc9bIsNber5
pbbSddCIbcCMmz+zgP1re9yFN4W1pi1uA2qy2upqM7INKTsYPjP4ZEu+RueM7OmiI2jHN1Y45uW9
+IbBP7I5Z9Tmshe+e/8S9wKlCoymEIiTV/POC6wSF2zfurR7vCrerBYTHvpdUQfYBtF7rLSlk6iZ
IDL13t2RXfVmzIbasCaugevIO27mFfqT/UAuZPcgse4RLBTJ9e1nfJzcwWsq0wZfivUF+IE8CXut
YamBuDf+U5GdbGeV0vMXPj+2dx1tuPcRi6mMAUp08gNp62GBEZTkEceh1CfOxBxQ7lc2UNVNJcin
f/IuWqC0KpkLkjs0gvujx5usknIpdw6SileUGFSLXsbQrMgZcnwtSq4iBQ8bdb0B+qU2kVdK4zGF
f/bXMMoxLxOC5wrLSdrECwM6/3XD6TmbDSa5Gbk9Aigd7HULsMF1JGgGKcg0OlfxIuP7Ob0PH2ll
ykoU8aPFEEdmZ0d4XH9LP8J4EtByTJA35u0B+zl76f2RYN1kVUd91FfICHV5cMeTdDV7sD+d7hBs
x4c2/7J0K1JxdnXRcgt8Ownz8L9AY6D74gNBRoWE8k631V9o5Rnsm28s54iXh82bC7hS3zphrE2J
VS6MBFHq3rEyU5V7O5dRD3JQtvwEuC0KWjxLlnk8DO2xJeS/WduT6z6QeKpQh4oAX5b1djVcJQvh
dJAUcTqRGXwRUrPo3E3ybpyR0fglojydzOYN0TdyYeESPPtmTk1rq2xWXsfNJMiG19zNZ6mIwca0
/0Uctk4TVYlGmKft25DYKcz4FobV8TYuKlo0YUR5NMhtIkObWnuQK0webPc/9FwgoCBR50Bnvlef
s/o2QS+Qa02OKDKfqOcoN1FYWCjcobLCL91t2yg9cM6pJ7b797rxJnLSYc8eFRRIr+ioaWfZrSYJ
VnjUGTECT0srZM7u+GCqynDFSXm9KFSsh88qM+2C5wYgYwMIu0Q9MdQbf2yWV7OFFzJkrONaGtm+
9f7wRkOEOTu/h9NFo4bNRYk6GeNFas/uhlj63YvY4AEpKDgHaQr18bXr3omTiOOrJHkAFuBZUFxK
c5ZBOSrTbwKs73mXpnJ2I59Lb9U+pFscB3n+gxpedxh24E/C8q3IG8nKx6nmIWBnmG3BdziOeYTr
cqlXnzqHPhCcLo8+QMX72K4MWYY8IxKA+tjz/bW5cyW+PuSESpzlKJLUlbKm8csQnQ5k3y6USLH2
/X3ia/fWNW3j9htVSKT1zpa5o2DSJNxgvN9+z1KLUN8P3gpjBMFZEOhZthRJmclkQX3rzfW9Y3j7
/hOilornVEmIS7jeKO4d+aF8mTSaqh2kywCaUy4ta/oyIQKF2ZLfU227wazsFghfEkvQBJA4SreB
6/bEPrJTGdBrFoyvIXlRrf5wI0FrRM0lLPStAUJpReCYCmJdGYGwzRGbD99sXfomjIeSkW6Osg9L
QpA6pr7IFXLE/qHKj983Q21JFkNHRHiGojW0tk6CfK59DAy0mcBrhqG94Dg+mEhyDCQ2JRW4WDgS
R08KDmrj+6xsj4dsm6AGHJPzgEPl+P83EYMxsB7HdoO3OvAxz1/pBUtwtSB9Dp+0GoxeC6cICaSv
5zt8uPklBN5tARjOsAVFNh94HAhWcCP3CN0YkBXTBXphV2WJWJhOXJd+Iq2HnVXNB79DW8ORrQzs
HmKnHh5qrc6kQfw9MKFHTcSBjErkcBtsDrkmeA4OLapcZbCx7m7w+s33CQqSv643Gwb7GpQ7CVgc
2vhhjaTkNaPZzgW6GT/lj8WOJby5mzFWy8W6QEp74lNh9IuelLcNo5YywNCgd2wKlNRL/al78ICo
DIbyH/RQ39Z9tmqUSKBmLv6xrcuOhPIj2dzLvFjp1LlcYDxp7F4uBkS9XNErsKHSASaIdnd7DGkv
MwTc2u/sq8zfAfWRlja3/Jdnhi7MvAOcCNb7+8ukhZh17B2O7qGJHHNJWOVid4T431fo8hueeq+3
Wul+pb0sEUYzvQe6pNXbgzPUm51+XeSkk4FIolU3Yl0TBQDIevR/+oFV1jxE6wzf/hbCr2W4LydR
c8YxiRq1YHzHQzaILWwOdom6neZj2nYT+hgZzL4w0ymqLLci0NMCleXVGqTGHzOeF2+6BSGihEw6
m/jfCqqxmzRpUx05gcTxinHYOZbfJU5eEjlSwPQRfKgejPMnPHxK12hbytYZri9EsJ/Z7blOcB4z
8NLWgRKGAl9AfQHgyOv6W2TR5tlbqCuACwMWtMaK1WfW3KN6w748feGsPHc32Kdp5OL6AKQjmRcb
KduCvcnLSqKs5Jz8HgVkVUVneeUaG+AtxybWaCgphhKw9D888wuho2JaEqALO+X8b//ZG8wD7q1i
nQx584QnFSDJmEBTLUQ7DyVoAuEHm0mdZ5d58a3ziQ2BPPpssMYKOCznYbF9TOZrf/CqoLYagu1c
PdzKo7pfugnKG3B1ij81o17mPxKT9NourlNHWRahmePcE7QfbP1DbBRR7b9pCregAnM7vX4i/4ji
HwHyPzu9vUtW3tIyTBBDRvNG+gyGRj3KTDIyM7/+sTIcCJBIMzF1BLnXmT4Bn8eecOvlSVRs74/i
aaEgEICeM6YyD7rWJWJbQm9C0Rvj97pYS2SqhR583C6jmIG8y2oS1vEvu9zc4gWOaReXcqD6KBTf
vz65X01aV1N3CsmAYhRs7LeIL4shz+HRGBmF/UhX/QTcMQPknqLCzndKs2gqjJ99sEWbLKZDoKhp
M2DDpg+NWtO9+7MzdEjLYAOfVWp5BiHDfLRBreuOm5DXwjSPf9UoL09zb7za+EITZIlv7p5EoOlH
/B2zbEbbj2zv3QJWnoPCHEMOrRIFvdbmPVzblAjrvxqVJ1tdJk9LDjzSKmCrYDcWdKuskDdzuULu
OBdIIdWKhi7CljU5OK+bkplNdko0RP+lUTHLOJyqLvMPvQ58KRMf3JaEjkhxcBRYJumm2HEEnA9Y
5K+/ryD453lpmZIRBBBhrTH/gURhE0qJaduDSe0/lJvUPbApcixgInz1KylV33XYEsjaB66A17Ce
gPrC4TLItP3foFn8nQYFetJPFhm1XExaMOk9O8RpUC5PmlGdvkzDZk6YJu4hcixiCOSJlve+8jg/
0sbxJCdqcSKkxlc2T6Xw/cV01PfyNygTIGbDXPNjvp5lNuemO7/eWEWk/wt4Ojn3UYyeVvg5mGkf
jSnW2QrMraemUkjMKpj/zXHNJoTTf+VRjyjzfrYmjcrApyYaRjK/gGmrH3ytsi8lvuPGyoGeflzd
SUt7WefzrHk73/vwKz4uvkDNFQEEFLEMXGidPG4uibTrSUj3o9LreHyQJLLwMFwI5elC14WtTiqi
avyeBp33sfDA87AYHa4f3MdPpN2uW0q81tV0a4gsvG2z0JpigSakYY4YSRTpwcGyru91aVMg+Oaz
wSGylSqVx0Z3Qilx12Y9cuAMZ/arXmsJePPZGOSeeOY4OCIy7xuEoNjHrIlaaoTD3MM/m0ApFBQo
zwWkhCdejD/UVrviUdzz7FME0OHZa9EozeB9sV9cVvORyy4IaD3gPWfL1/FS0W3ojnRFbR6r25Wi
rhb0Q45BzA/p0UcuAziEKwu+dI7ZeIiAaw2sp2F8TCPo6Ja97sPO+jgtmQuFbl4ot6N4CQGBguMD
PkHeALw2tGBN2IFXmG02+sstePrQzl+7wUlaj5dtbhzm7EJBXykEfwK3IEM6EJH6f04AU5RkjRu9
22FJ/0nJwkC0NyE0IIInbwrElH7kAVFlXWdKhvAjgXBxAzVNdjI0AhBxtixbX5a2j0Q1+juemw1q
OEp4hIbgAodnZdBS1IIaZZZPIDTM6KjAZDc05Ft/K/iWTk6njS3erYs5k0+mAlrwUnfkiTjGbeRC
mj4M7WdoDLE9w1Nhvbbx043bWJmiw5strDgzKGowUaLFqIM42++qB7pCe42Cn2DM1SWgKBzxxM1q
2CRMUJidMPc8Okh527TV0bPBnNzoakgOl+cMAX8dClxjzG/zBZOBrtU0WHxdxt5OqD3KtA/EsaaM
0jhbBti/N4YazOWsqPXYEsfJnCtqqpFBIUtdHpZPjw8voT8BjYHfAAM08WGcOPM41kpOLCiX2Rz9
ldzXhzbubGY5gPwZN2AZmIoYSchtVxSQXaXcIQxQnXVXyAg/fhNOFv4fJhOV0CQgQP2FnJiV67gJ
z8/0cc3ol0heHm7KEP7sHZ/JWoQAHqaWRQs/qPZGQnWG6bF+LD2odrUL3XrnMZj92J2cmpAc1JA3
nwgTr2mY6cByEYkEOAHSCWKb+J/jYmtPV4YMAlt6Pg41SfCQAKXoNsXjpCCYtIKYinvvnJxUXwFH
a4i709lOD9SnA5UTmeUTsZd/Ww+XkIwwbf7unK5cX/HGe0i3Dvk/Os/jTuXZbGu3nY0Prpu5GaG0
ShQ1Xay+xqrQ+vajXpAjeA3nvqSxvUoK4OC0BSGY0HWy2ls2t4JFxlvJSdxyyDSMr57xX25OdRIZ
DiHeHY9EwlOPK3epTaVEqyTRsy44X9w98rOYwXwarrW6y8FDIu1EvZqK81yXZNplykcKYfXmHGVI
HO5HrS54JTf062HXJ4L/L/fwQsuL8EnMNqAber1ftUGOu/eTBBlD/slKigvGhLUJoGcm9cS7mv2V
A89ZC2iex0LB3c3xxLf0k85okXfMJGan1lAp4Ek+z6NpUEywuGbNje9NtzV+1F+BzYQ30oHeGjsn
2FExiZu4mVwnEUEtOlr8QTTFNeH5GSMnZmrIv+uK1iYzEo1Ci9l2bjct/fiQDlU/7mavDdBkedd0
mIp+5wgAiU87P8u5wG/YX8Glx3T47Aqfin1UVUoiIndSqv4Xow2FeOkf9wU2XQMW+BbzrS+tzYu0
i+SrR4zSu1oqDZjqQ6uatGVLd1OCcsP6aYw2RaVA3qFicw8m40lYJGL9ELj9nFFiLpypvyKYvrzG
u9OHk1h5VfRMOJqq3wPxTVcmqFUq78eBD2xo6KYSZuPXT4r09NcgUGiWww+WXW/5a06vB4FK47X9
bBjMprKG5Zo0PHivnZYTIIHGRFFtyRVM0Ok//16kEEups1aZGyW6MUP6kUYCa2AVs6oZot1+cJ1W
2yBXf4YN+/iTi3770428zXH2daabZCcHF56x6C2aLvOAeHcqbYRB324pNUe8sYQNjLyNvaJtP186
oLWhKIQJlW9gsPXT9gNmfMZuDX4ATtl1AyVYwUCPctioxl40b4rphjvpIe6F5IZs44/4ROCF6kc/
CEjzN2WHwdJjnMuQVj/+lPJckk6XAefpjN3WgA9yV4TQue9zRTZP+NYweO5MsNFpefGDq4Ap/MJK
HFF9Qfke2/+7UWnaRYWGjuhGdwJ24BvwnkWB/XyBUW9ajE/lhOndLdx6hQgkhuDGYOtlsvfi0azp
gDGZC0ON0evcN/kxL/HoxqEEZFmK/+xICWm/jKudx0uuzITiUItc1UnKydoPA6y9trwWbqHZH9/n
QVvFQobCKFSd/vmQ3xRy1muQtluE1qyPltpcNb/KMlKOhQYaGoI9FnkZ4DqnUk1aMkcxROB7IWYd
oqiiz2GV746gPys+reZzB3dKvyYz9RygC5aXuVE6grRPrEXd5+CHwsm5YfUb4PMj0nxz7RlFWJr8
MARaXI7h7DY9PWIBEkVTPWg0svoXsDLBr1KNxFRhdWNX5Tx0Wfd5XvRk+emx/+eMFLTDwefGUa05
tpst/o4F4V4cEzQOiab5tZEBeSmiaOaDq4Q3bnYuYsv6JmA9wxn5vEQ8Iw0X6dFiAem8jUQyhwFZ
eHCcTWyHdY8/Ck2LCw2cNH8xLG1UZ689n2jIOv1wbD95NNkMj2eZXnsr37AOHgJODxFOSjtINpW7
awynmZsg/2s9phUIl7Wth57PNUiARTJx/EVMqy2W9sIjZhw2g7r2tNtVI27hV9qY9f7tDtMdrFf4
wvgoAJDMGWOnqx4jEP5NvL4mq5M7Nq4KvEvt0OymMuzjnErmGE2r8CD9pcHbIHGyMgo3Lu4M78sL
aYK1gJ7aIh3wCN5Xh+5hLkTnNMf1yfHqFn7+QHl/9YJt1T44ze8t9t6s8SzfrmUTjYbqvzths/Pu
FT6NnK/IVztN18rGxLyA+igUiDlXy0QgE/KX18/oHbUoYbIMNu4LWGoFf4mxC7EH3q1RzAco3pcZ
q7U2K3CmnECfDPZQNeNV4Rm/jwxo7MpLkX7fG8H4la0ex7FM6ZqmZXTrKZOhuC7A+44MbS17gUGY
5W81wReig+BdRCir44zRszNqaJ/jEl4Y4XKSnTuZciE6d2AIXP3OUh2qDVXIneh0zUvfZ+1J+iNT
sa3GXXXreWaNmCTzodHxhpM0PrAEXwDrUrAJinK9R7Vy157zB/7MH8y2wLCl5kN7ePyEtcIuCGCt
psF75hYhYkbXrJi7IpgvAXBSVDh9kO4xJSMcGLDhMqnZDl3f3sf55E37uFVtgAsoG48JfJ0HqRzj
8kf6plulcM2ufl54ubGEazxXEG9s44OIqkMGJl2sKDedxclMxqAYp2N9QWomKDBbaGEzljuvauXk
D6tOQVPAYGX27o3PzroL2K47mvTRAD0KquiyfaD8KYW+VOGhvKFnevEFXPjF3QjKEqHgOW/TrZaH
PwxYsGQbOyQ1AIhhMpDWCkGlshhgneOjUojCiMgxbVPjRYuERMr49rub8f3cgSVWAxoqjFO+fXft
gxHJvHbdxq2yPbh0pv3fjIKHcCpOm0IoG3luBfCmYB7u1tEEVeDjEJXvQHx3LJO7fIGtVUBlVLi7
xTqC7Hh66PcT1zZmRSDAIe+GWh3v8lHaFkgNKMGKjUErHW0noN5Yg6DgY+VFNlAsjX1kKjj5XHNF
z9j9BLMN4AuE7zU9ZnHZOJuRP3HtTru0xgIMC3FPuCncUBuH3tkoAFD8Y+OEs8Qp7lpuaVoZprRa
EEM9yJa5UNQMcB5vXzZDERaalcVSNZP7HUVKjYz2B5BS/YYjaSOfpDfoNjV6M9L9CoJWj4Z4D44C
xy0Si27IW3AbDIMnj6ecdCOd6vJdKmYumYTRmMFgulW9//8i8dnWrrvBK/+J2W2eMC1VmUIJfbs7
i2GbU/QqOE6wbNVxqs70KLivkMBdTEcgE/As9eg1dtnvg2indTgxMOO0kxuP72cmB64NQJ3U5YWb
c+ipbQNw25435wmQ+kcNGEeQx5A+syUaDZigZW72ITVq8C/R1Oa1HxaVr7rvC0PcXmdSrRPdf5K6
5G2ZFA1PHPhIRZrWPNFkw5a2+SRLviqPzCvnoKLmkvyhJBDsv+hwKwVioxzNUrhIMYCIFikh9LsC
ZrFmRRgpSPkBq/AibO8XHGI2Lm4w3geCOW2FZ4WKZ+OwRepz89ofrznlxhWQh2fzaJswaz7fZOFN
ixc6Yei/S1fMfiyCbRtIY09N5KbaLSTv+4fJFFjLzCHb6e4AvSXyLqI/aVmTSreMEl5AwsBi05b9
oE7A8SKmnD/fT+PGzsR+RYLX+AQ6F+DsqKMlYEdlsp8Nus7tFlFiFT1sJ9DTXmmAbau5IC16I5Y9
U2/wcQjvYZIb2QTl0UuTwO82QDaZ2ZC0q2Iypa5Rdst/NyvGqSjEEIHr27Z3CxdPO6u8uvIW/WD/
VlYzNIpAqfLWvXWlXMRTL9x+NRhEgN97dmEmem1/6H2EvtiCgF3BMv7OaOez6E2T2C/pZLDTc02m
CQ0Flw8IXbRpy2Y6tq0NwWEa2PRyg7pZh7PpqW0acJOEiadvruK7Q5eIyIjlK7QosKJTPrni8Qjn
PSrv6Yz6mIj6gRkFwkK6Qc4TDjPUbyxvIWLb0oCxDDq3PZJRKlqm77i5+PGoEYPFqIP+atzE7Vw0
cSxMWH5z1NDnRRNE+aiW25wl16d6dj0KfOWteiKlbr4wncU3EBu0C2FKnPoEaBqZR+kXDIwOdDEh
A9SRbvkajqUSEQRd0I5WtZ70fN50IMcLSrqKcjUvoK8U21INf55qus80TCPG1LR2pbYRTtWhRD0p
7nkBv6uk+5a1SfgMTtdXgPtq+kmmax4okODSUk7fFb60BjZo1pT0eTgd3s5oZH+fvxTQPdREQPlz
amN79UCVaq0DsmhqTgpKiM9AxGH8xuxDA2JjkM7CIkTt2pJN4+n4IjKRrq4aqxWU4egLgFyB2vDq
9eh4DU/8EG/0SRHTui7OO37yCwQvS8fRpx8e43FR5ncJ1xAxr2F30K9T1htFb0BhBuLnurPqG91B
q7r+Obmy6quhh1C2m16pwujs5a1K+lgWPMZ7BScYZYMxasOWZiDTXwU+AC0XJdXMmeHJTFTHo0/e
EyOuFK5hCDdxX/NRTF5rNZ/GAjbZOfflx9VpdMw/KQJR6EWp6hwJl3N4qN2ShsuePopig3kLjN88
dCfd3ggnb6b2I7cypMXNz6k0ojCGz/47dj5AACVpV/vJgXCRz+WFBdONsNeuEit7zWsqf9K9AjO5
Vp/N7E4ej8s0XeuJlO3cPRnttAf2RKPCk55dH0YBon1wOAmtr5+088iTNEsvd5UaCCVr+wJk1Ktp
UYHZmVA2cG6hoCFEccsg3SgEFEapmGVVkLxIHjC8Qf2ujmClaoJ/WM989/T1QZ3ShgSKXUhDntCD
5CbYwGyd0+d3D7As3XDu5+xEyD6uGtmI3fm15Q8kAqtVnAFbOtexQXPOB6yveznI5NEZd9lN+bJE
usBsYUA+SrvqgmaoIBv8Wo5x+lDH6MFsacjBpSReMwwLwaVEG2Rs7s01NZqwKrHS3KU6MO4EYNwc
YXmKIM90ZDEfg9UZj6cPujU95DAcsUxRAXMGNiH2BTlw5RjA0vkEMrcBU+dnt2EB4oyQzdHFYA+f
XZoDbNR8cDr3I2QtXBAEtEHusSSH4dJN7TraCXBh5mdsfl58jujQ5xvKJNEuY5u3uAU79Qhb7pIY
DcYN2tm7Ps5qcbjRXvjcBwM0VZza/d0xutnfO5vm22oQW0TuMEwD8xTpmT0zUhQc51SSdLG2rp8J
vtECm15fiiBE3voLeGTptWCWnuoKc8hn+tn05qL5IfM6SZIWxM5D/XTsYESFF8NpcoKE+zCMkNKO
Uk7bL1JJvVave7/OYYCJrIcqZ21wPGWmfqyG3jRkOtjjVO3daZZgu2W+3B42hpxMIh+wAatrAfNF
7sqT87fsvNugHi71wWQheBy5xV8Rnb+aBjJdZs6/7DkF3KLRnGtPegH0K7Rtyebhkgfv/SGT/y1t
CgzgOmgRzYIDHPO+ljBYb0kl5HPm0i1bojNdfxOe8GqxV9WQY9yHfJX7qK0vqpOSgq3f2jd0j9R6
wKlVQA33K87QxpeTcVEZyK0aw8rzwZRyhm7+0zEOVauIb8TbmL4iRmtGyZMcZE4FiuvnvbAUUj4g
bvCrRvvb7liIRgXTV63wkB6aeNVyjigqemECXhplmnSK0gbo3ZgjUtoeahB2dUGGU6xbFILoZ14U
0uCwUt7/3DSbEZBlgGTBD3QWCH3ZgjRUxXdlg51pq7C4H7L9tEqbVQ42eMQCkh8K4KHEPLpVTJwP
gcY+MbwR2JRG7peTjeATYeFpPl6H2VbFZ+Ija+isc75KA/YWrUynPNfMK/5Lk242vu72HtGhPJbN
tlYmXzoYrzAWetziKrAHr4yB/SCWa7M2FYtl/uL6ctpKdGQUUjtRtW8FHYCHF4cyIEgG1wZk86c/
O8yXynthsH1hI2yLjlfEgzTNcHms9G+4ITmZmQmdjU/LEuSe7Ipf4HJ5ZyxEHTrxsAMgIpHIG7NK
J7uJdeoxtpW+TJWZ4dZpDXVT/MAo4SzVMYKa68TVAB0/PUXummw0RutDa2eNkIlyIUCf13sQN29O
KM66aFfuV2889KShPmdd+ISpoLt6eJdjBnPjZa4Lrnw8QVCY5kKsjePLg5zl2pv+/n9ZeYQSdZXf
w7z6MlSNRi8zgNxpRE/seGcT7d1fmO8FQ948nCY2SyaHCav7byZ4YJZwp3mQTrNfe16RQoJ3fnyO
m0mLZsnYVcj6G0Z0jzZedWn7DupP7g9lD9krL7vpwQWG3lx/n+COL+LXjg2t0TiCiIE1eEpSdUsB
h1zqh/o+/fz99RnsOB/F1cXI0C59huCXRc5rj3pxEwi9jD8zoqsTLQY30Qoxs+ciL4tL6qHHd0lC
cp9au3aVchKsm4gdII7TQFfmxigJ5aWQAUOtyoCy8ulIsUPIvMLYwI92TQdsLrNXinHJt9Hwgtx9
jJxXd7e+3acCm6v1pueM5AxT8FoR5rvQ46r4UnJ+Y8UqhHrb4Vh1EBqeeGGPxGKqIJpJFbRkxfR8
NGeUa72lpCwl5GPDOZSdrqez/H//aycghBM8FJkiIh+F5KZwj9RU3ZeFBqhO0Y0kiskglCvWRbsk
nKunfY87YxIC5XPemfmlUDDIcr1VAhSqnwlc1RSwWSJnCpnHgyCJkLc6OIHGrFRjv1pQHWNNNCwX
JRMAF2Huprp6uTQq+VikXg7Y67xDwIosg1/kj5ipH2/QQPZon5lFjZYkWaKNtjE2UdXDpt0niHUn
3zwgIcT/U0r2h6e/qFh4ow+UG/Sn7H4N36a1vK5rn4LvphOJQR3F88XU1OYz+6EdFfrtwSCD+egA
U97dq60dRWjqNoA0/3xFitmTPuqpO04ayM+h3FkpYmW5TgnrrHEMuHWEAY79UdFwTS38gDK4u1W0
Y3FBDckHGLBFIVlsMEn48vN0c2tFscunWcQTxP2nJ4x5Di950+kOLKkWFLT+oS4DV8nGoC6Ngvrf
J1EOJmpWjFcik4KT5lENYAXGUCRyqYY/VrWB3xEH8JhOt/jZPk04RYEZqrUtDEOW8fPfA2qCg3MP
TmwhMwjqP5mYBTVc+b6m/imI7c9otw7uIa1ONcV1tgvLM2yXoThWDx3bhqBttlEn7Ve863Eb9EB+
ZQ4cbyghQBpQAwl0FTwejCZECp6qkUt1JXBZIdo1CrUrj0bejX0Y42IdoWA14ewtM6fOL5oA92sC
yb/7asTxJ+3qJB387dmVX8HaItS/JzKa1Ni4BIlfuAiz8CX7ulu6oiREFBl4LzCsVOuAvJ8AiFKb
eTGN4jVu34W08cvTdJvg/TUKdyy5GTjP9tnz+MT8ei48QIi03i1QdPAjLz98QV34A2regR/5n/dR
j5SousphPzHYJjmagNCq4I38tL/L0y5d/a5FKVut8t+vymGxMC7H+oGXGspuGqxqvV7TajHE01Pm
DZabA6o/boHLxAOXILdOu3TS8Q9KM3CWpSp6KBwkyU3QNoxfCE8l2SgXZkZO+M8hY71nc5/iTGOu
5pMp+L0iwMmEswqzVRmXFcUW5CI+H4cMUA1y3QYchstUajAvIA8XNDaLyKCXRFv06RqSiyxN5yZC
LR1rEmDWtJpCu1RGxkLVVOwGKGeW7GCGTF/JKX56iPJ4uaxTz9Dk5zLdogmvf0+GY2KVrCa+fY8B
U1EvI6DX/pM4cqr7sHFlNtxv3lYj2pzPm1gPDq9dBAC6NcqfvR5/Hn+FQJ+6JDfCPK14HRFK/SrG
3+T1aNHKCnIY5WYup5KDdUL3a4eB5Z0HiBooV0rxYeH6pp6ZAsTiZ5ejqIwcay30BFVyQ2D8L3Aj
QkCaInJxfcmIeYA3Io39KiNK25jyVVJoPnPWZ2IflEMLt5yR6TpHKp/163ZYiufkvNngsK6UXG97
FmJ55inrowEXdJFE/1TNphPa/ToJvzVzd4iCT2NDmyxUpoWv7lNPicAlf58Vipw9vapzrqHQB6HZ
d59KNKDAnRhAy7KOtgImniBT8fcQWrEbOGXaqJptrg39FjjTobos6HVQhgSuxgZZSW9mvVUqd9wT
pf2msyIrQvdPQdIELIrhg0l7GgG/ofd6UdugNwhthQs6sE45oaS5NMEzicS8ffMyLYHhvuhL7ZbK
NtTuo2kOmwtEcNI3JPjRaYQTqFlDNAoaCgMmQ0Q3HGRTXcts6EPaDDj3gY1gGt908gorRv/JMj/s
Xo/jC3tQDb1VysBrjgekoTpQtX8pcDb4qUKGwGYWYLH0OfrpS0n2zmhB7mlykKazbxcjKhsdpHqJ
iZeYE8KBNkHEFhYRvht6CMznDTsEVcaJHAuRDen8SQeBJBpFf5jEBdumoF79CfEMmOeqyZ5LC2SZ
X5g1tfy/18fc2481f6iNpxdw50wHu5FxNNaOI37Vcga1+WyqxQv0Y26ErEP3h7FC1aHk0s/PVhJf
uotQ8A+oYT6R9nxKE+TkXtjAmTUrcFzCIFW3Wj9h0jwBzU/AwJFNzxhRjoXnhfQ42QWXubNtbH7M
S5BaVpWvm/rBZixBX2ec3/pwLGYEllTrRJDKYPm6dNJiQjm2eB/uQ+qG2+v1DXL37GeeGvTFyROv
cvEMN1WUBhCL1sIUeTcP1aU1WlqqT5xFvEwEDOwXwOsNDEi1mL9VY3yoikC8yvlvb/F0FTS+tjZh
ZAym+M0OT026Ms7x8kWupHqJWC9yUi7VXD2IyjGFDgAa2Yi2kSAY2ONiH0ly3EfABjKmH6jKjPtG
1dxTNZgSgYP/NOTVyjJLX7DGJRZwdWkMtV41bSNjnNf0h32p7p0MPXEJDinc4APdFbfFGKiJGmqK
QKm634XFJpQqKP5E3Ca9MbBMrOry7ftLbwA2oOk/+7lhkMLWMCuFgiPFWZolmXRk+03XzAwf3O8W
I63k4vXFsaApCDSX5swoxMZzGGp4ng3ZesSqImsuIqP/gis2dj2vJVpI9IG8CwH1VWbsdghuPu0g
QPYO0U8CQRUF8JHXM5ukTogX+2VwnpwIkewbsISnTwgz09G3fyiyWpxjsJlaTuqNDkwkU+CeQwNH
KyexJVYzS1pkwnZ/EQkYINgJ6K9A3AoFO5BSt9+uJaxioSHgZhB75aNVT2JubTtheIHOto1IWR87
Khg7/cX5ylatM7R/YnV+NtAwZy7gIIkdzEexgb24OmlEAJcQ7KwXsg07sXLeKZR8Lqi6dekL4Ihb
zEXCTk9hDBSsNOjW3NUzX/KK/xTNisQjXgMtyrRrF0pFeT6RgUbjc5ot1Hyr4RZaXcPa1YBzlQZz
KRgfHMRyZIKwjYdDiCB1g4QOy9au3QsBP/sg+sVtcEy3Js7fXoVTg8QeqUSkhG83gS8je+CuqDki
KrlwQw7oUXQ9XHS0bgZ1xL7IT+DByyhb9Ov3pTmP5rGhGSrUxO0YPTUem4YjeAP0dyY9X36dwbad
rxtVbTfpvhhLpOek8uxjp5RPbQ4SZ4f+mCV4cNzirM3Ww9Oa9AWuioRXH2tLvweuDo9LsUSdu9mw
E77epaCAO9Z4YqRYKD44dwqZoTPuAhRaJfzxviipOfMUk+0qI7w6xdzpQmo8VtzQXk5COpKNeAgz
UW7rDeOBKfXTfOT2QF+E83xmptiTmLDty9y26i8RWrrzhO2qxx16jGYC9LD+pJehUNXGKh15A6MY
+EVQWh7OOxZxx7LJJK5SiLbE0g8lGk7RzWqWvEfn+iTqBiGB3sHCJ21TwZ4T5MV9Iwz5v5+aEnoj
lve3PnpzHkb9h3aT08l9Qfrts+t4OabIkwXXc1OeZ/RkAEbskBtAVo4MmzpRFpzr3JX5MebJV/o1
9cmPk9gtgNc0t9pLkXH/0c8bgrlTYanISBU5eHOAFp8oXeXfZYtDUsrVJE407LGDR7eiBwS89eqK
LM+HegnRJ7YYktSFe52XqUNfshCxjAbRp0y1XnJtcYjWwzXb9wQ6Mf9/9fid+iYAzXTi25q2nPqN
N9UQcI2pFQfjig1OO4Nd4hHLE+1X+FJdKXpd8U30KIY5lwD3RahxvP4YCzIq81jhEGWs8Dn9XMnE
wsKga2iRXyIluyIr5KDFN7k1EmgZq4dXhPaaisOEgoL7ZxyeOX/LcF0rMchgHljESvtuXdvXq8t/
aSgV8etEGS9pKb8YAb8EcxubIexMlY7PNyYjJP6+8BRJuZHH4ZhwdY+P/n1Cfd5V7yyb/9mIyvCj
LNtFaYhl8+BhFQvIc5OVKqN6dLUIU3pf4X1OhY62iTUMtLvmowMhpctZT1VwYVu3rpdfJ/YmJxHS
IlQC73q+GkiV3pM1DxluU+rImp9xt6WGepJAIVV6ETYcUxQIdaTuoQsOLtHnoI7x9wKePZvDm91U
kpKhokIpqeEYO5aBPF5xnfLnlMSY2xvofkJU8J4QTp1dF5Y5tRa7i3HX8iEDUyQhhOMaJhAS2S9B
ts+ZFVSmnlZ2YNqLLDEfSScPVtlipN8zMa+oY+QhtFsdifTvrZbyxSxC3IWoJDvv3w1w/T1GQZeU
6bFSNMVtkWNOdqO7hb7TvfcyazVAU/E6gMVd4X0V6wuYYCR7lBO9vR4v6TSTI5ziCvkPn97EKL92
YUkxAy/YWlN73juj21YaaaTixJwQqC/XPLeWBN962X9z2pJUfQfsxb4cfmOV48rN5ab5335Fco0v
vrPu1WgdiQvjes8bjLm2gPSn6dut9/4G7O0D3gYKiVlahKyRjSzO3pI+jI5fD7EGNVLqF3mKPEHi
AapghqO+fIOPCzeB7sNYL+7TKVFEVoEmWYz0vvD0qdxTuGInHrP2wa1C61YuaWoPnoFiHK7sRggh
V8wspw4NT8wuxFesjDnxHpMz7KUQbPJJx1rvm70crL32Wxtr0LGn8OSwdhNnIPLeZi2GBKiHLIzR
cRJveVkHTqJYzcpog7hsz5Xg0uFDT+vgEOg2rrEflhVJUWvIzRkeBnCUFH4xAgVs4oH6yzSfR3Ik
g/xXIbGQ4TNF6spHLzLhiIyt/Pj5LQhjLu25ylJToj/tuBTiebcZG0RISCsyvE8FxkU7QcspBsKV
HGo9Is6qBM+0NQShhWUbT2ssqPipIQGNe1wigcxT8gzjXf+qxbMRepu4r4B8l4xO57xUpIUBKKbW
8/p42OgdGDFbm+b5YIjs2NUHlJyYI+F0XYkqwet2HmDpHAnhhbxt7Wp87ZZinSLcz9HSaplpA6hc
mCp9cMn/famfeYH3eGWsQ/C8zRaZ7H++paxcyVRrqlDigy6LzBaLrMuVn7OviGDdvCAk0TilrBRZ
O+dlvMcq2ZsUmvIwTzJotgE/b57Rk+BClfky757QyBvo1Q045MY6SG1mNPDYfcLKG2bBX4J8kdgG
T9ScTgHtlz+h4+gHFiQ/vshJXHEN8y0ExsR6+nNCS0OvpVrSQX61rvojr7FgqURYFO3o0UAolbOr
/F3aDIpAcCELYZwfnVg0ymkuWM2GccAqWlHI+WGm6dR3qsZVShaopXm7tRw2Gk9VuK5ufM1amJKZ
Ji4Mgh+5e0DykoNQcUg/sPpUoeF93jCBO7vHd77l20LceaMuvZLAmcp1O1Af2+pWJ81TCS9ukuQ5
nLDHqrIUNRGMGTgHdjpXVhHCD4RyLpVMjIGGtiM54Wx7Jr4UsV67JhoLjLIULxhZtbYzsdX6L+JO
8h/G+ajNOOnZdm7U318X1wPx+cUWC9kGLg+vnRU/4uf0WZnGueiLghy8UJu+BKSH+f5J2uhMfrXY
GU0TJfeaW/Rn2F9QXjfnEZ+iZK6+6aBg665go252bVzYccjcwP3XJoQvEwSRuwSUEkxRxO4pj1sC
d+gsNSUfGjBFkIqwIPqC8KYtPdIkL8z7Blp30hUM3SV1p64E1x9EnpBKuzK4B90+Dwi6BeJzDnwo
D1SIGFkAN/HL3skj0urjlTGGoDp66EwJoSlHVEj4asFnBALye1YuUVe47nXDUh3UTFpwEZ5Adece
n5CXH+XoQZqwvT+be+9rZUqLiIgxgKdfoQsyZBlrcWl6tHQXYeVxeWiGGdP2FkVjQ2WI5WRp61ET
K8B4nFq7QpOlWp/n3JO4jFxBDtckArs9qSq1yCVi1q2sHGm5ZJngDHwTwT5zT/yDX5Q+ijq8kZyI
BQzSmsC26gB/oxeBtt2psM+wJ5Kr/73HGsnadecqa0XIHf2weFUgpke4IeZdvMp48kE0aJNaJeXL
c1fzOPGdZksPhV54EqZPqA2/8I1HSw9HVbjOzHBrLNTUaYHf1KzhyGnAPl40MfAFkd4sIXbVfsU8
NKdbFQPuzOAKhaz6H3FXDuOiYah9FYkQAQdva8TBqFFA7n6uUnPl2vLrTwbST6JoSGLdovAz6/mt
mD+HWUPDwAEvdjBZMWLRIvHH3BqsnMA6dvgKOGCpzHisrcR7VVbxmgO3dcBm/M2EgyW3Jg7hW4dY
dBuzJ1Oneqmh/oqqgSQqs2AJKXkVoo/CQOJEJr5zOQEVEzgUJiiektzw7NCQfdCcgegOFXVrGLku
m+02EWVZ53WPepuq44CRaHjR4YL6ZGPS7hRrItsqEvCVjj1qVgNrxkHHx1HBW4f+BXI3qGUaAnfr
au6ZYUVQhfXTrXquSam1jqySltTjpU39+1WK7TFhiFP7USI83qii2BlSTF3zdxYIC8Q82FVEAlNz
dCdxjL1B3RwIvZ+YbrJi0whC2/SzebRKspfKeDb0bO43kGMjXAb1bPnoftHZWCoy9YyfkEdtmO3L
4gp6xZdZGSNUoPlC8cWsDNtNcRbYsP8Tt9O27G2zijhmmHJMQuWT57gLlww2uamNiG15PECknGyX
nMCBCJxtmcQiL3bdBpqOXkIpfpHOYf4Vk1RLOcj4TCxiMULdnT3qmC5RXEwv5m6Pfm+D2MFhg0sH
UrhnwYvAELTzUMfgBx+9I4gxDuZNMD2PALS6k1Xgt5l4bcNPF4t7poqRrEcRpOJcUeHgzCh/u3a4
l7sgP8xBVV/QhNOxi3QqVsi8JEuOLNbvRmL70ifNqoXhb7Jlig4zuLChBD4lMEOI2MxyYydyGBY5
Rvd6lDu9BSVT517Xe0Vs9uenRQ4+lQ0d5dSb0Slh12vGbcugcQHzugzhdv1Lm1atSgIoVfdIRSyY
qeGJwiv/+Q6GS1RHj0Fl2RgvA/mpLh7wLl0zEA/MtLqYk0sE50JPPdclaGyZl83dVsIVh4lhA99+
z7S+n1va7t8Ss248f1Gtwfaz+S5l4aBjpHHEzQXByZks8X3QGyIsnGiQF6A+aXaX4Ywc9m6dSHiZ
xsGHzBgMEiCjbNXpJHriltkvzb/iwL9gqKpagRwjio0jCNdik48HT3Xxz+ZQK8L0CzvwAWTy8P3b
lztfVPFiOvT7kJ6DA7L9GlHdyRp9DPW0tWQIs7HDLtJRBFBCkGhgZddAqHq8TW/J3ojMFrHIFfGF
uuiV08CBSn+ZYeqJzKGbwzgkISh6Pbbbe/7385YVo7Cq0gewX+70qU0QsXLSZ9qlMAJEFd5UkJmH
wAY1Du3FUOLGazDUPU63q15lGiO20ceKFIUfDHNk1mkJ4YDuy0R/LtawC3ovXDwzZr4oxldz9YNf
IlYcslBK+ffNUkGoXUncaN04tKjJFEa6qqUbAH3Bugfpfzw5QfBOqBa+wZqJLdMjok3ciy/nzwbw
2yXzk6VECCHN5iU74nwHk8ftlgjHjpOOYe9PbNTnb8fgSsu+OeS1LmusB8KIy5dDI/gt11ZAPuJx
IDHEGFpMb6mnCqhmL7TDf47dLAPwYrdCQeanClZOKvrS2nKyuD4eCOfdJPAknyrwKXv30jONXvap
zS5Ckeyw9jncwujToEjA/bhEYF8lyN1+QkIAEfTTBCZVP/gDf4KMMSx/EwZRxH5/OuO6ZMO8GksZ
Pqf12MKxB1+pEoe+2P1qVRwzK0Vpx8vuhTGPWrngoOw0pfP05kcCav4OYbSoOASt6vpy46AfkUIr
yKXR7BSvBy1SZ75BxxFE9HIDLy/Qozs2zrB5I97IlMejIQ9wRnc6gwpo6E0ejnJKhJ03of7xtadv
QUxzjWDmDZUYdaxx2G+O3ekEz49EwoK7I/WZXmU+KeGAZur87Y2zPNJoJ9evleHB5st4kPalNX6h
pS/6A690QKu50xGdbXRXw5gsG32RZ0zOp8U/Am743Vex5byElDzPYPuKQFMJoFkO92gVXOOC4GQB
lxnnbLbnhO2k+dlmG7Zney2IqUakvvVsUPUNBZVjoRDwqjigdr+t4y8rc0LopyAdl3mE4l+urlaR
EZboOHfd3Z1m0CJCjZoxzKS0N53Ru4Dlxru9ut6o2dbpfNgaHlZUvQnyi2MQCwHWF4kAaL7bLBma
YpT5Zw/WiAH1PaWIkOzZ6ePJHkJpanyGuhOdSvY2rJu8qbVJGjGsjPFCk/t5HqzNPCMwkUwilzPb
DMMG196I4j+CLkKCoXQiRHg9EfGxrD7UYg6kj4AZZ7m86e2ubbvkA8KP9Mr5zNw5ylkdrnfBs7p2
AIe+8LsSDkNQDOnfQOLj3K2yMMZ6/vyLYC7coizbBrqOLzb/SRKDeVb9GiJXPw7tOq7zJKEUlu3/
HjNQklcRQF46y9+Ad55LlCPR6ZdQ2vqdsK8D36V8i+Dn5RAvNEPjQ9tZ6F1Iiw9HdaW4F42D8KHB
/LZVt1J9bjEC9kSABLYZeAyQsJAkTWVZiwHDHwN2RAg/ZLSO2bwsaFleAnLyUvjqZuTwMiD8CN9M
QdLslCgYDITEvgudPqyebdytMRROg0D5jsPovhmcsU3+vZCo/pVt6e0AecTp/BxIHLJnltsTWZf9
Q2E30/qfMwFPJkfHcobu5LFYOa7QXPyvcVeKsuXT6+vdvo+MJdghZ2y3M/AIQ+S4kopW0DWutell
NtVQwAi4yWms8G2xN88oeWyzu1T5ttOWnCDOznCxEYgwVNdyjXiDTgzdb9VMaD/4lKukVEFeO8qj
OwuxpJnze22kLoVzEzYj8PTLo5yIgYZ47WZKF4i6haVyTjYN2mqcdTEj4WEXTxRiBkjUx+XTrh4R
yGoZzo0cRT++eA0K+H8pG/UhEhBLyc0iK45duvBdYgHQleNTchtnCulFIOgJANWp3xejsw1uyHFb
j6hKAMioFwQ8eT6WOTsguB7yhzmeOJT0SDU/E/zkzzR7iVACOxjasYwh7qQ/p1oXdtom/OZB/ULA
snHMJsRWcVBeIEq7DxALZ9TABnjXuj6vXV5h09KZYS+Sr8d2eHA4ij5wldf7+UYQKNijfBCbtBkh
HuUHmSgpebZM2ny3q3gQ2/CUj+Sl99B+9x04QBS6GdHJrX2ydoj0XMeY3up4/STwR8qiG6UYgNkq
/M9GOHzkOnogkxqXm8gKTht5j0EpKRj8Zpnnj/JifVtishnsnS2WF8O/Q/ufCJ5rvv4LH6zf6u0e
HDw3l+xLGX0G4/jvCTsN+n/5YjHFMFymIc2zUgElL7VUhMb53NJubW2qwf+3QmW776tgCvl7aiVK
PSGOrwOqKNbApjOr4RM3UEbMTMOSZQ4LfmYHvOskreNfcFlj3TntTjd8pAGlcV0MMzu+IwDrc8+z
h7axzP6xh60LoKkhBwJeq5UEckNTLY7GvyDU2wAitr3d26CthW2VNCxWXu9sx/70268uT6hoAqKL
8JEFxvmrPe2XdGAr9av4PhOuh3ExQI8mVPCzt3vrIQVbpag+Z9IEx3UuXU8jrwYZoviFg0FL9PFd
erPw4+4IQER8kUO6zmDLfYe+gnFgQfer46pNHdbTs1chlWNr1v65dPRJT0lxnpONu/qDfYekwXGW
Jn0Q4mYTGRzoOpIyQKRB58EKr4LZGufblnHCckSxKVcsQM1jX4Dna9L9uqpF5KcSuPNlRkJB8A74
kBGLIWR4qv4Wrq8IKV7MdpuslOBaRvtKY+7iMXWyNdlZRG1SCYQqp3ku9kOOSBCG+GipYu5i8w91
ljvC1MOjOPXIRpSJaYQ8KpACxXb4/BI7GqfParMA9JSV3ddEu25A4giCX3D++8/J0cMd3sIxpBmX
SAM+0ezkF7fJVq2KB7IOM2vNhe8yM9fVxzAb+HyJEIjNhAav6WrFCe672LdLN1KwCLTNYYbDQWdY
U/8LMoqErk9M5U4CS1whTULpgxfmrDMucLQHp+PbhKgtepNjO9ICYgVhtoNQBTcP8wX5G+/IfvxQ
JNDYgsy+QFBOsDSrF/mUtqEwvtc67FaBarozuhzY1UHfn+Yat0lU7KfctSZj+MrfYoCHUZ9TQFDz
RGrwliSMglTVAhgTBLGWRuwOtuw0OABJ+W8AeE31JSvNPPGqSugXHV+o7ylCaJlYuCf2yEuyTMJH
R72mGNpAvGw3f9+gTwi+SrwEqtaHq63yBD1CwHT2YGwTkv0o1iO6mbP1PMhA0amzcUPuR8TY4VLK
va99kl9OWv9GBC9YnI9ZzzEoTnbkHPGFEMc16ZM+zQreGOqPRSD/LddL9hb2spXKs/B4hfTqJnxv
IayHynx3if3sjA+QE4gddD4I6O2ZYvXO4nVs8NShOJGxGmq6lD0UCxB+R+sEkI8XB1qv9gqBZpet
AFfQF8yJT9skS51+/hDt5xFPj8aDKYYIko7G1vhgq2AhrT3HdGUDffPqnQwqFlGE/cGoK0YlR+OH
pcSNapZpY9yHbyPmQLz6T0TkAb2zwlpC8+I8R7nPm5topTjvQCpcq8yEoODYOz7KSOKf0hRVqHQ+
0ZcdAqJlTj4Y99gDK4o6/TiDhplf17Nufl6SvblJQXD44uHkqCvyGkxKHCknAv76T1cHfmjf+bvF
G8K34ddl81uSjT91GEVxQ0xGw5/BuC8CvAsF6IHAykkgTGg1kqU9T1qhDlUaly71OzPHwETV76Ao
4DnojfszLVjdzWHwcGypObITRy+dcuwufNXl08UFOAgrXjqKlQO24s8mEARVIb4u5H3Up9xvbI5f
eZFrMCcUnjLMP43wQ3HM+2XTO4PdQK2zYsr14fGgYQPnkgM7xkHedU9RtLev2zq3uRS5SD9mymef
FDe1Ve9UeuEDL22wrw92SBPZlviPSIiqK+q9giK03QB4GrFyj6UOp+QSwqMKJxAFFPuAt1oaf3I8
e8o/HaMnxvEVXQrqiVHJLQXPU/oOUr8AmQJcCL72pnzw9YDxNiPZnlUlTivYnkXAFOUKHKWL26kd
mXO23qmkMqUeKF+YK4S3BzLla0sQUotEyro3fAgT6CFGj80+JaKyWB+ILSRI8/TM0w7asO2YE6NB
bKhPrCrYWDddS3PdcnBJklrjFT6eo5ejJs8LShRVITEMD/nAw2GjOBTiBjfndsCz3fxfWCjF7d5W
qb9s+DcsuKkkUpeSzvaQZaJe8b1DtcL+2lCd+uV+93KV9G8OcwXId+fvAgWZ1El/zP3TaJfQzPzn
K27Lc9hC3t4O5C8P6O+OwE9kc2Q8DcTb2NSnJshPpLgjty53KeRcbnP62kme7WcWbBxcx3CRvnfP
E8BpA7h0p3PhbCmZeLHMsE+2rTqfM6ycbk2wiAJwNz1fGn41n0W3pwmL0xkpoV63N+F2aZawLmAY
uKlg8bqRdjplCjCBpLqtOwFTRLAcxGar6kOIJn6SP++zCYNPAmlI6872AuLM9Nd/5KSnjlHfoRFC
SdeUZ5vI+I2GPfVDlJmuo7DndAyCBBEvv0odE5jVWwAH7p3rKHS/vD2XU3bLb1WXsEA81KuQGzC6
CvF4ebIlbkRBEC1y+iuJQSHfwNVp6o2rAsTgHYqrVAvBK6k39Afn0EnLa3+DP08TGfbzLUjvOmun
HDt2WmGt+Wt3ZqOg2biSm6/vlABRyjAp4VzF13NI/jWXoWnvln8FgiNm1EQuzebewnOnS5vB1zD1
qt4o6B2Pgh7fCrNCYS5RRKYmq3N2rXQD17eA0uvhu+r2vISYg3E6qarZ4YTm3yeLfgCy3hz05rbt
vb09RG9GdPdeyYZVFGItHfDS2EDKSoyKzwp+RqG+0W6xWgCkW6qrZynRrC0egu3bw615JvjUUcz4
+Cu2Fuwy+G2NbJpF6bidk6K9hzu8UOGipzjeMeYZPKpYGwZmkROR/4OIgutNtmnosMq5BLaV6tuq
/Bdc/kiRu6DuCMNXSsOB/emI611twX8BrpE4yXRwBfkHH37BQqpbyv+2NpunB0N8BL8EYCXS8oi1
wpZwyLKlSRxQ3ba68oWsM/3PVyuY37rYPj+bL4VvQ+kEmYk66O+PZk/gwUR2phrUBZaNgwBEcXs+
LBviF4UGNg95KVY2a5A9K2VMDj3hD00s1JBri25jKDREcQDm/BvEt+C4N2VLjNZxYzAem/FT1TUz
/gnTCbVBU6zr93NPOkmv8E+/ajZdWI3i8vkh2sNSsfhPKW8qs6RHk3+0Pi5wboY2u3MT8zabfNmM
p/CflHmk0wTxpfTa4UWsrmKrFE03l+PW65w8MhzduE7y2EU17K/JTzBJ8vPdcmWwnJUlSK/dNNa4
Bcy8tXZ+4ynmV9efvwkw+vGIENtww1gRoUV84H8qz3R4RcBkLV6vEH+FpRzB9duCAIr6AHgcbKAj
aOyzpVksRt+QImAGpMXWKsQPrW+B+XrAu6lEUE0J/kuM4cf1WQeQlG1PWSBUnxL2vojC01iOkOxW
qeBxIkGqE8dK8DqGTA+FBg4qxcIDvhkfAGbEAit/QGBHgZLs7Xj552iesYIJBrdYkCOHdTHEdHNv
dU/sK2SdgueLpbXJXMCG9y3yj1K8NB6LghlUYa+IMFfmJebaIzG5QHNEvfD1EmF6wn8wHfQIoMUz
++fC0kFrbrbMm9u73pslA7bgbrskaijKSSIcLeLKnsyKsplDu4cQYijBWduwxAzDpgPXk5tDhGKO
12fO/kHFaTr5Fod5Q4XCSCxM7IqSUonGerFosMF12OuSAE0tWVhPxJZveVHR6Kz3Am7dTBQ3E1xD
6RbxeHANH44ORpamG/7wZE2AcYzIK63WZsFZxBEXn4gh0C8EgOEAi5Z5iE27MYuZ+osn/+We33SV
eiJ4y69PWXh8e1RExU1i/gDMOC4MUkJ9/JO0DsfJhHKJOiP1kdIjaLXuz19+RWkbPmTuz91i3tq1
050IpzEdDzJSsNEMNy3M/VJPVZGcmxhAGcKlLQ/jkajv9njdIAptCoBjC5ESDxA5TzoOJxy3M8a5
7iSlgFoUjQjranVfLqwzX9Pu+zAzlrAzOr6ZvIxPf0y7q5Wjpoc3rpl/1VEsZH5QC0H/bN8GNogA
0ebjjbpemCFfyJjaB/JI83JjmSkDnb4PrfeXuw47NEjPiAU0Vf6WoVR3vpnfAQVnz5tEJgz2RauG
9fMf71xrAxjD/XOcsXWwLw+/lTRKe19Ar4/wCJjD8GKj9jRoFgT1/Vdp/81miXj52a9uUpNMIl3p
Glf8HhrCof60OCdYrIvq3igAK0tRO7iw8BxHuLVXXfdgavS67KOlecj2m08QEdoH4yN0/DoBOBUU
Iy+OCrdQO+btKhStBTdRv7SBiIFT8T7HLC/6exApF7itDhEuB2yYmLJOETUobj/fpmavZ/BBaXSo
Z2G7H6uEY6ZXS17eQCkfOhfVxfS6x7TpbO5nAPD8QbINNYBt7TsiRJH1nsSvC3vA/wCzNFRXmTXv
uytvz2iU8d4xrQ4aIpIBiC4nowZBJMyTkmWqoLkW2l7xMf2XtTsU4MJtuwhknsLaC5EpKevJDuD4
fTwKbpucdHFtVwHXqhjDaLBEfXEZVenGN5N/97p8hWvnC1Nxp8K2LACWo1HhiouAlXbV/XJGYawv
lIBwodr33RhITRqMDYUhL21J4TMgbCijQrPrK60Ica34BYDvM3zanzpHIUV/nI2O1fplfFvFEPvd
WMQXE2Mvfck7fLZ1llXSvtpw6wiqJDdEojd05OFoD0BW5VaVQkEbFSdsghpSSAsYQTSHTKHHrKoT
S09dUcN+o0/qDEK/cHCMFjUwB+6pOzb3lqqkkRauuRV8PuXl/cNFVYuypjk+a5acyG2Gm1iugC4/
0c0uqejug5y7DkTwlfVnbUF0RsFwQYQg/ByZOq/QrK5dqOe7PFfIdkNaGAxsxGeXoW8RApLEWhtb
lX2VqbJyJlWB448KYEvXDi51FMpSg9BvmEmL67asz30yk9m8ojG7pWDPktOOzGUONy6GwFd87psa
MBDEKlGU27mrQERpqnrBXD4JUPkYgZkZTON2lAhxrllI+3mjun0DBJC9gD5IPI1EcZKqlvhvGt2q
dxNRs6/OlkWKIRIYcblDCUZfS2cBzimF2YZmq23FYG0YgUUFGkFfQK9qwCMHx/TIdIXjURz2QIDy
qN5mNxSPp2JMW1bPy1T+7cljKhl5YmfoMrpPzah3EtsJDQUNJa91TPvvWd2DImC0nqoqKjp18Jnm
i+nPBdXK4CJW2j0DsaOTxGsTAIXLeDVX4MnurZmNZT6U2lRFvd5op9YFIuL9jMct4cJxHwca2tTP
uIZRwyrcc6R6/RJZ4sDfTc5D3UJQ7B9LIIEhWFxeCScfZx3+xUC1rPECSpwcVcOa8Ljbw6aDe3MD
68OnmostRQiGDhQ4849hnqKK8YnKlHh2Ni3FqjufxRlDFDa/eBflrH2h00VQaJ+ChFywkbHG9HsP
qlRBJJaaAVlSa7A+wu+PCBioVtxfRNNP9B+5dWOwo/7VMl/i72ly8JkbHK+yDCd/YR2G+1+Xg5TS
eJWAw31bQpiAbb8drGRLcKRql8hMVfwmypHcXKGbCUpvZ7KWxy0uwNw6CnQFDlrtcWbeFKCziPfd
K12001dCqeGBNTG+k3TPthEdRWQTBcgqVuP+MYnBBmXagq04u16qeXmO5KgzOpQOZ8ZsniDH04kc
jPtNRnT/OZJygKCXwlZZst0O0+SnPfjQfjylPZ36nfqNW1EqR1KfFbgJMD+QY8BsH+XRTU6ywkVa
yDRtpmkxO7cvvudrBGv6TKRb+mclGbXuWCnvxmhL6BrfgyKJtSR/ydBO9OrHs6l3tSZ/AQ0fs+me
Tax0pssGsIqoWeQBrxufJmSG4cANPH/JwRptLwA/GIXixhegzBQdVDLuKyIMzc11SfYw4odpnUnl
tDPM2oZTumNZqZ3xxz+wmshaee1CbaOJsCyw1IP7EH6V7t9pG87wuih6fBa+Z+KDEzh6Nc8PEXqd
S+pWldM3UGm1E+WW2Cui7/CwQf0qq2j76JS6wOJi0MQSkc8kLm+Emud8AJ7xpMbOKjkztAujUHz4
zLofftDWU35qc7++1jCqN+t2MDbIpqxCm9znTenYZ+Q2hlRkbLkl7dZBBzDLiz98TR1xWIsABf3Z
BfRgY5gWWnH/Q6oL/VMeJfUrhTzLHTOQIzbLI8w43I0pmNTY3Tvv5wXNZDY45B+eHDwo3esPN8lu
vZQ41uoEE//X9uaMw+5cZarOO9SAcJZTPYdc++Qfb8Jzojk26rWr6El6ftu0e40Unnt4ehB2FNkY
1AM1IjqivW4Onx8wxOXDQb0Gdea5/1pUcfbERMg1qselnjxbkKBRVr6TsOkR+/pxmlwo4CTHIvQu
sTnNuc9yn8axeuZo9iVnJPTf67umMc81cjYYnkImaRgkecurcCPRDTmvJchD7KTt2f3HCbAxk9Al
nuLklFq1r3e1otNeSRM1rjXxICRIvNQzqs0lKf3pthCV3szLdxCEodhHJz/4EJINXkYfLL6JqKsk
6Mq8DSSMSYfH6sf9AWOD4hHYXeJHVoQ0JKqiZNiW9HloSf9LnGki2W2k1eKV/w7ol01RS6Ntpkvy
WM6ameA6ir08FcZyBJvZxMwa/uslUbsdJaBTfQtP1lQkkfJOSYAqonclPWiQmUhMxk3dXCePLDev
hhkOzh/6+Bu3TBnSWtbB7rFHhNeq6K6+GlYIsAamba+02BSNtqLigyQ7eI2/fgYJZd2tFAE7rien
nIkqeAcxoTHX7ETahQ7UrqY1OeD1hwAz8I1BIBlVcFLeD9yU3o4vw+t5HDB5Fei6IKg+zgAohIKZ
P1PcvPTz98Yq/TdZzRihbb6Y/cmHBAYLbroVtJcqkrrfNwMiD4lbN0A1kU4vmhgQ491APN4qE/VK
NzMV+CYokmSTFFAuKXCCP5NCrBAWPB3Dowk+YrvmrrkJwIUfkb21RliSxgONWsGyYVf01GT9spI/
Vokw0kXKhfzg0ugHTuVsXCEK5YxutHuHe3MxLXzAxXCc/JEmHGU3++OoMv6vGpqKyErXKH77IjG5
TQ/FohLAxi41CR4cTkdbL6edK/PtCAJfTPy8zmr4xRYfzPwMaYtYUqYHTTbA0hv6RZzLJUKg53Bg
7OOIwsOLHD+VjHiCyfJW1WqIegb7wuX7AtSsgeTCBSujuafJYjUgwpl8Yj1QWoKoXSkIqurC0IOb
wyGOW+qrU+aTrlkzWSc/VxHap6GaD/L5raPLC1KjF5dmJTYgSgMVwFqVBPiZqKdJ7hYV7LmuDeEw
3f37gv3ae2u5S0wd3a90uKnkCYReTGvgpgibJUmp/La+cfiubjvZa9s6u0QxjD3E9bzLJusqwHhF
vBH6vSbO6+DerK5kGyfZGWggCQEwTFGVmdiswwOq7EQGMy0a3Ppad7y4jTN98gzUBePjul3KdXC7
KVwAmtegV/RZKWufYTZqwg7mx7/ht5zae4+BTcnNVbigbycOoptZwuaAv4kmi1/AACWLgcuPZW6J
oUYS7E4IkQTYf2bzPCjVxOEk3gLfYa5Fjw9WYY31LYq7If8NXuj8YklQo2RxTO+AYKs57tYV9Qpt
dPvshhY0AqYAUvzcHKCmLCDg0MaFgXurGCv4aGVcg8FegVLk+LyVnHIiJ8L67a27us3Xo/gtEmFo
ZRTl4NRMUKlbPgH9d2uXtiL75b2KxJVOrAlP4rYKfMztjqHEZiXYnCPMQyyj5wyRBWO23wi5L9w2
TorEQbz1+qiLw5ZPi5ycEPza1mNvhpPTWX867nGqXUi4X+7XoQKT9y6meXIGdzcVJr+9ByIPKVmT
dh3jnRMSY1nHCfdlebOWszm+ERm9pH7aYpTTWanENrJES5LvszwfqAfHNXOZkbDQ/teeb38xqZyL
qd6JNwy4jGLOP4WPRelJcI9OQuAjpJS6zsduesZ61a67PUge0yd4QqjA/EE/Feinx442wiP4+GaL
HNKTrzCdOrJ2JT6jva8W2eWAe5ahstSisJaVlwjgQ7R6SvI9kzVnCto1e+b3VYjBxjRuCqirBU1N
5ipgxjtGJPaZZIqvRXjTnihouUFnOoZoyFq7efzCE/DFrGr5lCiLal5KJhnz2/yG/I48igAAQF5R
vFhXz0e+20tEmioNeYPRRu1HcttkO9sL9XEe4IZfkF50VaQwFSW0D4znZr7ivhzodE1795+TzMXe
uA4FbUb8HfeiGoO3YPUukT9He9Er1qk+FrNSAZI/i7Yct7QaklZHQpSdg7zXBwxHkIgKk5fIWhuH
jiOiJswWUox8aFOPPWLxqdisdbOcJL9/ssK6KQmfySbWdXZzr7I2mG7NbgWuSDrAy4qFu86xg3zW
nnie3KRH1BExBmIVgVFZ69UyYzcRnuJc0TsewR7zm+fsEAsc/jbM+by0l59a7mEkVU37zs/5+z47
lYuAaHKRFMv/jafw3q2I6xHg6dWH3j8Fw4HdNNbtL3zlZq7QLS7PBTyL0701soW1dLXcUYruqoZz
BXKqEn7OrUtpsAGkSyjuu29+svifdZ7gUxgKXtRpnmqRzHto5bmfz2uz2RFoM0Wq1UeThZnPdnqf
KcUFQZP+vBR8fYeaqQbL7IrpqB9MpVVSFJPT7rn+fmJ+X/th9IBNYPApabV6tGOyQcwRuIhfdzMx
yOIp+bIDd6rxMSS0YlXDHWT5q3uepPvCXwRFB2CpzvTBcNNURCr3zt1wK3RKeCuFTDCwyYKJ/AEo
zBTnzW+6NG/vFyRKB7dkO77AOmWiVlnnv1mx9lzjAY3AGEZ5Yma9Mkhrc0ewjbq+bGj2M1nJK4CK
oTL2yidOvaEn5ponG5dWSaW5diHW4RvHyfh+3fpJJeIsRPJ/lDeNgjyuWEczWacBy0sIBOUaWUmQ
W2mIkNoPHTer1o8/FM0/oN9/1GaUTs8Jua+SvSX57KS4/U53NvC9ajAisPQgpYQN3Q432nXlOJrU
OpXaER2Vs3wCHpeJja7nkbKt1RFI9LahsRneLC7/+/14UuHnR8JLjIZkRYxAJiCrX1+SwSqQD/t4
fC1zcJCdhK34uquEJlTL6Vq/FD5HADwaCpnkHlCBYrgW+g/ctYEoie3a4q9d8clYyLV1wqZhNl7g
8mBwRSFngGABVpUW4AxFwX4dJtSNAsB0CVI5Wu7ulQpXuygtLbZNfx02a7oVr07DOaxkcekyg/GL
kXEvNZ0TN2S+L4CUwQOe1yoOwhnK++byiqgVUSUl2MffqoJOIgCvYTUs6mV0tfkln2NLIy1p/oUt
wqvODJWs+C6a/53cZzbqgpVTt49m5McFb8yS0FdlgtZ5i9RykaiOzlG2v862wgJPu0glyAhDKDC/
99ZR1bznY6vzroTAlMoqqdXwUkOBmqCAwL6Tr0weAIRe4LWWnixw4bbrl1HoA6hkzCiMJ6IrJlEE
XhOscJDnESI3FwnmPkQ9US7nsa0eXBSUaAW5oFfBO+3jCPU6VPzuxoersA12WqmMgFBXzrv81eQc
WrEvEQmXnARHavUuy/JGfPT8wofKYtvCQmXVzJFdIAiL22AB3GI1EDLu5U0fUBJNdsgj75n7DsZB
v2TvG4Op2Y7Wdsz8eS2/LzMVHXeFgBYzqKoLvki3sKk1yNU4XSbfFadP7qJFuy19+hUMvg7GuZMY
WtBYsK4L2k15AqWsBL+xXgEZE0geYcCD7RnsXF+LMJTp+R4CtLqoyp1ODXvqIKGKQ4BnyhpUNFnE
4siTeYI+gbzqSd0+apB65jusFV25RK7aYgTqXdqltZ7Rt5ROXvN2H208LX94NwrMR/4EojE5L1hM
SEI3s7SesaS9lw7LxtCtRshleBETnFz/cZVKXWrHpG/32HlUOxLIKF0NAJ6HVPnkOZBzx9bwz7YB
/pSfalK9ESXB54/yU+iIwaqX1n2irOcalyDhDqzhdznT/XhVBJrxjoll4WxN3+AeuXVqS8NKsONF
K/Rw8zEv8AVGpzsYEbqkQGxsL4W8RguCISjt7FqOJDxOWjsdAb8pU1OQr3Ph0PV7Ddlbbw/7Ex8z
HE8v+00n+y/J1U9V6e9oMfokjuTCUWd3tLH5SxfKlg+pFBYHzSixekis6KWJUYKsJXuLbXQ+wQQf
qW1rth/VDWTyo+tyWejixb6xIjCOrQGzhT/s3UVcZ4uaL78Nvq60vl+poJIZMn28bvLjAtpuAIfv
pMCa5CNvOMF57/gLVJ7gtcNFuUKnfoBfndhH22Q4lMHkUYRiDdbJxry+LpjBfmp4Vk9YBfQkkLIr
c2TagkWlXWxih5jinjvFffW8+P4vT9aCzU9n3FsUsFdQKIBHpcts5ngYey52meY4Ubwg9gZISGXB
T68rE3l4IWbEL/lSrOi3A+6w861NkpfutUDb5KpzK3ztM0OIRHOcgy0BS9iWiUp5AQfzxfi9kiYZ
jpENEEmJYXS9Ewg6tZFcM2XKHnuD5+A0RDcDuZn6qGB7uOOtJSjhpC3Wl+/ZC5vu88X06E1ckLKT
sdCgF0TP5fJWsAyysGV12LLhj8rTynlx7ND3kmWdporOg3DkjGcYoL/6Si+oiI/6O4oueqyARzMR
2Swh6Zo9Ok35N3RKXqu5TgPTfYzmIPjI/etCQ7iI3z39Q7dzWzyGglMLgtog1O/mwK4mOI9MvFv1
IVD8Xbmuy1V+Bd5KB2HTTptDFc4XZTk4v5328qZZs+KCABhV/ulFtTk+gwGho4+nJgH+oAIxlaOA
bp7z1mlW701WFxB4hXJHetac9s/xwN8hn1AEtnPeN9TIdRZUUMiJqbEe6KOSGKLzRPd1iHCY370S
QP64l8w20ohcduDFBG0GzmjWWkOrcVtRsKpNsfhmcAwVWJ9uSawl/1BkOI6mBVfYoooTXQvyUDbz
aD3nRjMOqR8oykJigPId5MquUbAvimQ2bU1FsHCOtO6QmFqcK3lgaOnh7RGwvwymLNgQcXOEoN2+
29NczW/e55LUmsiRrycW5pHngSdCww0OpGNL6TdB9pCTxGPZusuBz3BuHv9jhoFGRIiONMb8RvH8
PGdaM3a5qVF4GgvoaCPSS6qZjq/nqEjQYp7kAhN4MlwBn39o6kLdMvO6KigqWwtWQIL4IwNSlhrC
2//Rhb+nAuJ/bVlNC3ZomuZZmk0mmIr8ygcEiOXkR8FIxJHJ38RFFoUZSptw1hRssgWy3voZpCSV
GB3EclkYYVHpVrYHxEjbdY43bhB/0b2Gcrok9VDjakzLRTrAPlGqAahYRsECgpmCqOQUUZJZKWcn
UvFRx14seLcD8gLl17h/hDiBUMme0UZ3R/FhMwVjcmTPvcmNMjZOxhnsOIp8ZBr1QNTrEeOlYOrw
sv7YhcsAybhC6Qx1b2eaI4xcefLPlvyJwV1f7zf+leNHvWX+RXwRyWS1YeJlqekTGKHwFmPkNE72
hZ0obWJVVcuBGJuraCthdED/2j78kpe2FlO3xv3IZ5KWSsk0XNJsCfhfFyf3e5RnyVaxvbQaTdH5
ANFPqzSkixX9Kk5EOGf1OTzI/LszAczIl2i77V6HbDF+92jjGZN62x08FxVbolsX8bFld+u1SGGS
WlAxCK+meexp/pnRfsmvUGMs+e1vd2Z525vb/+3l/UewUuHnXm93WaGtyl0qt//4YDnhn2UQRSSB
xl/5T/pXDFZ91G8eKKJs2k08F9GUKyD18sW1/37h5xHP7HVOzxnH0uDoyJ7RsfSQtOlUKKNnMuTQ
FXEqdA7c7rQ6INuBQW/pkxUjZprA++7ZDP6tOwtm6IUusbBYnNsaKDjIRrMIgrivzxNU+4oghPtk
L/78pO+PpdMPyUtTtPidZxH/KvHB0amNP3jO3IA+dgm5geP0jGso6rJG1jRMkaCDiCYJWenWy5JE
SDr/iziwuG9adbHRqyZMAtvtTVi5/8wNRKivhnMXi97gPUhx2TkQk3jqYTksC794r4CvBh4g7jOH
So6JWC0jj3UYVm8X4s1L+rX8VV5zeboxMIwiiN+eDik0M7IF39PKENKyzJAWOp5snPJVB4fn5Xh0
/+tMnE/ILJYH5J+lrjuZXIUmyIFPhvcqlRF35KF0pJezu+3+6/WbZmoUvlo7vWD2bH2EaxkuK+0u
iYLaPECW4iXCyM/FSZv4SIvqqHHK76rslpZidvAleO9Hn6i3oRQ1NRB0x0ahJ5CNit3czhUA2c9g
kq0rCDPVME8RBjnd7jrh4CJiNpT9q/LwLxNQhz9zppeJce/Ic1Td6Mx3YhEAKzV7EMdYdd2segMv
o4wInuP8gcn6EFibsVk8dsdd1rFxSQwS5JM1po8CYjGadCHUMp1GgxGZn1jT7PlPh52AJHdJua8j
JAdqcJRVW9BN+dDGjNup7+f1XlpZ3qRCKNNGLc5TQVOa9iMPrYGQ+bvgTKSFJOyYrpyENRbj5KQY
fmsxk3OYFA3DbZ3mrFWJyddQjh1ZgDN8NBplL5AT0Uv03ktHU1KwBFO6z2Fj+4533CYBM87ndVr0
FUG794xo1aBgu/A5Y7PZxtqx5nGCrJAONnOVGDBk71zNlaSGRhBLL96KilY2F+YTGtHIwKrQPrzD
3G1aPFW3MahMgU4uUE6susfKpY/YdPf3tRvcfxD/bqmi5Y1XKTAwkIuvXCxyvp3JcUk5oX4Lbcph
a2+cuA2JNfssBKxgHsi1bLiwvgFp4ubyioYp8qGOAcKKbdWI6Ctspp3hD4RuqejlCV5WHLVQTy/D
L5mr6pc9o5vWNp8/m7AB5Wr6M8ol1LaqkUXC8L8LCYOIH4jkmWaAI0prDcivBBWlUEqdxakF1OpH
eqpFZp2Xdnf4dK4UB8yJydwASd1HF7NGpcylVl4AN4XnFUv7/IwnRDhGEvhg3CzyDrthXeEDqKKJ
ABr6W02mZbhz+N5PixATt8hhXhU2ELKATsWBphbKHqonJ4EXp22l640JjOw+sUCO1qjPiNCE1AAi
NbWoLenSCMtP0b94Bq0eeHP+NnqjWMf846Aj/Zrt7PafYa9VL3VcxlAub64uR5sPGYTnHd1ET/t6
Akr5ClafHMp3bakHegfZ/LsVId5r3RV/FnJ0LGc+L8hsEqDtH1LZWnVjQLCblns1c12Fpx43K16W
G7wNdehhvBt/N0iMSWnd+OPFmpA2vbkI4kOKGU4eVWq5t+0xvt95vRQNZnEF/0+DQqSltcT+bB/q
Q6UO9SOoLNvpqTo6qKI088aoIIEYXQPQXaRk0W/Np7/QrZ4gNXOYJnsQnRgzjoPQAVCiYY4kv1eH
nKzaxDSKYEPoKKUwRc4RaDyBpFCDaSls/Yjjr9MuQUaqI3WJ4ylXG6SMDgLaS7j4a8uXjkrhJ1Q5
55qkXcIWcTPX9YXb+ojnHax/4CtEhE/8fTvqXFYRsWIEx2w7eaRItJe44ze8JMLRl+hJqz0AbOpt
JUWXVGHZlu/lGtQMjTIa7EaHJzxm1pKF/yhcJdHsZ2L2ho10m3e3dWa8otGDZflFzAC2lpiUROb8
nVI1Q+mCHHOkWMrWxYGejDASR7BFlm5+iXrC3VEJKtXVIiQ2PmV681y5mMmwUEf9NWopWYzqn6aF
wYCqlUuwsvnJpbXXrVNEwtMbqEZaz+aqY3n6w4HKE2yOwWx13gfKOCOtZmokEDDVmBA7uDoVyaVe
crkaCa2VfOlKCYSzywbqngHqPdBmdUU5eX47XevQ0j10RS+5rK7Fp27OQPPf7oeMRBGYy0INkKoD
2EVcZg+c/lxLUbChNzkEsIQW+T27bBB5wGLP45VcRM1YsOxrp2XconOBo6bKfJ2HlTA0H1EBqaE5
QChiC5Z55brclaYYUGoiNXt9QdOxPyBegkP8YSoT+eCpDhQ+PmmLrnvT/mzx/XdMF2Uweo6csCZ9
lOQ0tmijUc0mpyTZhl3BnuFRT7r7lGiwbbZ5eFWy0nZNOPuK/fCSM3Lzkh8OMUXMQMHpRrIfxIuG
bhDxV+weQkpFWlNtvoIum8pBlsWuWuA2aea+VJGqcFE7sB2JLuHy+Y2NwgKI0XzDIN9zovOz+Vxq
MQQ+ChYCIty3JyniE0mpszZCvYrsbH5N3s73sWP+V38bEP5UqqSaJy3fGdUszmAen1LNZ3DGjDpA
uDQTqvOvQNr2TepXRIa1rarqI9YbCA3gaukaRNcxEcfn5CisHSTUswnVUZGSpg7+0Xxy0VLocQf2
ABYp4fbQ4uVGxn8phY7i0UzwMjevqN4j1iYzRWMjSvhCzIaui3i0E02SXjGK4wvgd0YcjZwtg8xV
e/tqurPFnxX5MBGCnsgrGK003rB+r/sRA+m96lv/tHsJNuHMhcA1u/Gn/EuC38lMhD/nWqDRY/Nk
DuxeoRKoYGwUsKbf1lczVPTXkFQmAuKkRuFSt5Ha0B0G3LiE0m1+2XiFReSePIuuMHQHtHarAYqq
KGg2Zb5gUw0KafCAn7c47MZJdJZOwcaEUW+rrVqVj68rX/uFw23llTtHgAk0ZMsBY6YzX2rBrbtr
l1D1oSSRsuxT4JVqdpC8gDoOGxspibZdi2fwmLGg8GpKZlVnTMWmaNaepnhjnKfmPVwTzlqbKwZg
WY0pGVfspfbRYl09Iu+laochHEili4voFRVrsEgcRIlmDzYr+anhtEsbucl4j19pgiHf5Ay21FZ6
X2ow7cQSUGPQvy9/EoIGFHNoR1qbk2xpl3UlPHV2kYYUxFYgNi9M4dExWT04+rg8Xe6xvDLXDqbk
nZXsr3c5Ln5UVjS7Uu/4qh0n2jK3M7GfE5gdn9aE0yan90/q+bGyaf4xYtmUVJ/Qf/lkhP9qteQQ
v4slAvakn7w5mEAlMd//KYOMupF00ys/zOib+HcJMLpm271ODiEJEbnSnWZJfW4HV8AakbVP5PBe
6qsh6tvfTDGnV4wh3ICi6X9pSNL2Nrk9hQO1Hni4YvvzHEaCL5MYhScY3ezvHgNiQlsKbzy9uYNa
zNBEvj9nN5PrjoQv2a04E64LBlYLzu8Yhkf4Wz3typ9GXa7uVX5ORPC3Tc4iV3m/O7gFwffB1f53
AnQB4TtsQQy0G0XLkYWxSSLMGAsigC1azQ6J8kRC7dXq4u8/KRwlErk8p+wxyLVzV3Q49VvQwsdt
mK/eDKuyKqZ9MCAdJ4PxPn1jFBF1dzEBBAezOelQaA6PZVLK1226sFwL0Q37+4YtVINzAhvPkfro
32PLgt8P92uczxujMqhug+e+mQEZxCfubPuR9+1UIQrW/r9F2b4xBECc1X7OE6+fVnPfYHdB1G+r
aDZ8TzGmVqUYRnZnXO/E124i0KQmFFTbPkpqZkdw1PpzaaTrRxeRokmmvYy3xS2VC64mIxjp9pqf
zNSZzlArNot6/KVb4LhFn7IbBkw9FykT4eGpSZ3G7ov7TxDL8IrOEmCEF5k9v8EyuJinNwehna5m
+OGUxA6antJG1+ctQ6dVGjCxNxbnrhG3IEIWF+XpDb8WdYf/2jVL2UL7jB72n/+vhXhpMuofYl1/
0vVaE5PEacwHpvA443ZHcxr0gK4+af36j6smSQW118GryzqBvCUzHKPLH65scyZNR3KrRWFwYSjU
mdT5JqwwNG/TXkGqSsjdtFTbh9RE9GABpFlci9lXfwWcanPcYAkHYxrkho91d4//unhS2QmZ/QWN
zGtqIymbyRyvPnpqPRM/3BDHXbSblmdzRqGF2R68Lsx7zsKrHBwsbmhepyBnKb7peSI7N2XhnOVn
LkJgCHucKUQ1lcYyEw6L2md+AgIz3jQnF02CQuGUfP4G3/XgRYcBHks3hDEZRzUMiD+sSloWkAWd
6GluiUcxGGxH2E7CLedsAi/YxxYeL+oLJoe7vtABu2cnGgs3agtniQ8G7cDlOj3lTNUyxrw4pspl
8FKhTP3lq9m9VB/X08uSqAw4Y6p1u/Egm+viwYoFBB07YIHYIs0TMJVEPcSJPJfd0yXl1hz/zdQ2
88TwOboV3EwZ59IAygnMWpDNcs9jT8b+GKAo+6jZtGXjEa1ZshXMTjex5jEq3kkTTjJa8JdFd21q
UUXLiq5MogWVAZ4aaHDZFlWwGnuR+chO13s/yhvdnF4rBR3jz75JLu5QGch4Scz553BU6rhg+zxg
G4WQZZKCr2/ynkawrlz+I1x51w0BTvXfDv2lZzhMlPoyuBOc7BpOTWeE4BZk1t5PwiW9tTURSIEm
/RXs3PdXDNDrSXZBS47a/hVdUAzqCQuA0aAOuCI2bb1HfleFXo/StigQ+CCvhDtWPEgQwr2ARswc
mQ+s4RyxIhzsCQfWKqie1+BarDjjf5SYXQ8R7BrZBj8M5pdtJs/PKPucsmfJBcl8UDrxlUCgvfI6
dikJHgEpunLwKCgq/97J5IEi+Zd+vzqAf3COkBd/oMnfxiBUTsqwC5GOjEV37OP6ov7kI8qPp9iN
6waYWZ17Rid+uxIcj6b64BvCpo7d/pnpUTh72cL1a+7ZJqQl8VQd4A7MzVWGdVmZirGrSmfKAugI
TmLMq6k80buOI4c8Um2wAmyrFSqsqN8PRWqia/VjlIdN3Jih5DBE3HKLkhQ6vSNsfXey3ZzE8du3
D9NSMRiLXk3j0d1Q7A2HhjGO/fsRLMKG21xfw2o2qieeX2yYouEiVJrDvB3TAfVVsteHIGtmJsTF
lbVEEUq1IO5P6Ah0sL/XOjhvLURK7GpWRlMxaFRG3FqkM36/A0XokcULYGlVXaSszF3CptpSPozd
sIppCtDVCU1ut48UYfhr42pP5hh6+Xiehsuf5Ct60Ch0ctU3ozuORFpcO1gTRlsgynMc+Ir+NtAT
9DvKQtD2GHTYXNWLq5d7gLPthFm8Bjp2FRTcQ/Wm0jytVcdaGk9ySi3eHGJX5facmCwJUpLmbUoy
EmGbA3RplQfLtaDawiPqXRz8GAMrvtqawLjY6a54xNfLOJgrVLy91bdcxmbQgosd97GjZ93NFijY
RXxEzfPlF4oGd3WCSoDCR1kQWpl7iDOQ+0+uT+PZ1+T3zLE7NZi2Z6N9rAx2KWhtL/k/4TdaHypC
hfAKNrxjOe4PAokX93qymZHUzIqs3BhqfiFqcLyuxMJPKX+ph8u0DoOdkFXKzBti1iCBSSzAwtXU
GIH46zSHrj2i6kdSGLbOj7xjrCFK8Z3T99TJB4xkB5o5z8YD7qkPApdrCsP0mjjvJBb+QEKGV8na
VXHswcCY6OGo94iiFEY0n31z/qvPFmXZm72A5cBAjzyS49nfOwZZWdhu/Alp2utSfisx2QFuy6bI
97Kgc0bHHXG40k7NPc5dcmI+/wwsmyjqj981Rk5oH/3lzwNUEG4Ye2gBGL+aUNeqvgUWvo3BBPLJ
TRpcRQdhlAcrE2gHh/9H0f1XdK3s+eZWie6LtdIp010EK4X8vucCzzx8oUuP37AMtGnaN3a1dx2Z
eTtm00+Cc7gtq1SyEtshHhqXcP2GlPxxJsgjH8Lr9VwQqpRIyno6bOw2YXm/1x6UHEbvGXmMlqva
yI+eVufePaXJ0FsVQrNo23xBhI6dFh+//K7ysGJCM7UKrGgikWBt200KOZV7lyWKfCvSOEyIguZN
7r/drqo9bZZrmmU+TzN4QuSdCe4f+oKHXwaHcgJWoeq4cusmCVroUC1Z/oigaUcxtSM+Gc0AVBLN
s7adi1dJCb5X8HWa6ptHkaFcpOdHw9Je6XK9IaZmo0t7zDSjQ3XwY1fFJ/qDOzsRY1B/V4nq6/XG
TmD1vR9ib0ElWPsd7iVSl0qv2DZxcMugi1Xh4CeN8uZw6p/4fLv/GqTkFuFvr10mU9LMYuut9tR8
LBGTEN35LIoZ8kdesfRQRs4+RKvLSMamELsu07aNloAWvQmGtwfy1gEOGzlR9+Inu4Bi3FwIqJYX
4D8sj3gW43Slk51hxIFm79Z5sqg4EGtNq5X23IaCTFqkey+ywC0gb4xT+/K90pRyAdp8S5PMEC4W
gAeDQOSrJd4rZwDN9/498kO+b+tEwrEffdJzJFUDgPTaPboayF3XEPMAQYzq5iAY5EW9JcvI7Bpm
Tx74FVLdRCZaNQIYt3+GV1mlTIU0eg05tR8L/O3p/8z2tLUdfv8KkqmNbNb7A8KsNipi+0eK0NeQ
fr/f372X20Iy8KnVAJBdyIGm4rNcAUjHwagAZOQt55XBXJf5huX40vU5YHk0B3Z1hV0CxNhybDD5
rnr+lot2wD7wz76Somhky4e8n1CkGkmkwx2/veO+CJci45mTwu5TAm9r1IJ92wQjw+wMi9wsYexT
bIhk3iFCleewEPTxhBurCbZBQooJi8GnXOxE8hZduur1EpdaSgc000wrZeSkJrd47lJetcz/gUze
p0yEcdLqI5wZwVBk96vqSn0maElMJzPeGwy4bzYq+d6hutG8tASZwAxcGANyZt5ACo9yvs0z1o0a
zwAHVne4WDYUwA1Hfnbutcq/BgOdiVhQGUCYWyX/YaoLsRqefRK4Cmq3cYJJEKDnEX/kaQSOwa7X
7r9JhhRqWHRmA0sPOaXiSiDs9smIcjh/lNI3gajZmdsbln363H/YlGM8xTQOdYBbo1v5juNYwCEo
a8GRS5LmoncKVOYBHBR08Jej+Yln9Q3BG2aKPM66hJiINclZ9eS9UEmFdJ3H8Kbtq42tay3dkHbI
Qi71XAVIzYyS7j07RAixyXZVbOnNaTmdb+iLl++cySkBKlT3FQ4vWVqWm9tcfOPT5m4yqMO3r3xX
Wo0Hhpkot+P3+2WCRi6kBhXIHVlvZPP4AxVSnmmh3J/g2tqWK9ie8gYeP7QGUQKkNsTwAwcC38Nm
bne5T45TEJxWrDzzOQtpoMQPgOU7nnlyXfGx9cjqRV4a6pb92RhlkUKai68Q2qlUYIGbapkcobjc
nWm+AlwLQyjgzSQ5KY3yyipTLW7fYXOxiVpEKqR4CIkTdI1+bSQrb7lcuSTOYIZ4B7oBnU8noQqr
Y2MqAfegU5wBJnvfaJA3/pVYda+0GwMcZ6ALAg5bSLW52rirQ/VPXdDSl1Dz2VS43gr085A/qHQw
GcoAneYtL+/KOCUUuITUw0fyxzXxWVHrCog8H899BZQels7TIAvQSRF8goofhAwNDGFNAzlmZtqB
9vXSNFWHtJEcgu2dbvfs/Ofwfd1AeNLoG9ItQAK7C+bPRLRB/Zg4PaRtk+r7GAq2+Ktde7BuJfW5
VbYpdZ/U3BsFnyIis+9lF/xm0CEQkWtrQLQ+6zXCZpj3NJbKVu0tC1Q4dfxFiTXPV21bQxO4Zk7u
UPDSYpnghDFBUTnwS83nvsEFp9XEc/WEnjSMuBOD9oiOdXZ2V+RsUqZvaoF9lX/YnaOIuwFG4BZ6
zPgEkVTuB9ad1eIOscnv7R8yXdy+eY8/F6YYkUktd0/invrFQOy0WjVpLlzHRU7X7gwg1VIDSYgI
H2X+OAjFLcfSB55aBz+4pW3AumPpbvl9Z1y0wNoT21RKYz4WL/XCrxbyeG+K3Vj5HJp2h0rPUJnv
xh4C157YqxQ+X9OuqawlVAyaJl50oALrq4yyRJtfcjzR4xJGWjO0H5oIO+juixxwk6WQCj14UYz1
FyORJh9EqzOOYFW6TAX2ZY1XV83OEhOQ00iPyns088c9TGJzM7ky81qY0H9NpbLuwpw/r8bRrpz1
6DftRny3o5zHNXudxsuGHctiVcLywd8A8nZmN1OaBBBDqygVO68gj3/9APdXmiPlOPqVjKfL+w9D
Kb6XO3k82rsL7BZGeD5ziBh58jRhqJcXRWUFUh/Cb8UGMdLWwYWDP5W3g7TGsFjD5o2+O6TV9/sc
UtWeOMBGFn5BjWXbzgucRjKiLTYXi7bPnfDvcCgxXzLHWG968HdLByGztDGSpZXjiQmwxjKcwION
F2bypiVLvzf41i4LMJUTawn1D8IiUZMxUhMoUGhX0EHOprBHJy6w3nr8alpfnnGpMNcuOuU2a92k
32lPLV1hbMAzDJobKiYfnrkiydjYYNfvFtWnXLk0oQ16tW6LoDPMsZIYYBi+KFBYeohOKx7WlB6/
Mn3Z2K0Up4w8T6hQc5vhAk+wnrsOQR0hMBA/zLjGGDGdaRXwjyB6yfeSLvCPWi3p0Io/Epj0cK+D
QxN7E2C2DlrcFxrJpMH/LjAMKD5lvqxlZ2ciVuO3GSOJBckPKMKyKbiIUKsxDSVyubDto/F61WYU
pmNPV/TKqAsIdgdNMgp/COwUX45OM5sMJltqXYZEiUeLftnGI7hszVabhkk0yi0XNjEV4TZ+d9jl
2KoolgcULbIMvMgoEhWFQXr908KVdb5W2Yt7xsv6Gk+FdXGnc8B+5tbvpC1kty9kC4zPXPnGkS64
WQuhT6B1ht22QzboIoZFr9yyKOj6DUA83JJpNz0U9XsXbg9LbO6NwTjOVRB79HDOi/FV1HnwQX19
Ap1z+eBHzWsjF80/fNkho/3gqf6bT1FeoC2PMrsmiyMH3c1aeuRAfT69Hal1xHfEORb8jUhRw8du
bcpLYz9AnCDcqDYD36z8jUQiz8unNIq66v+xvNzG7R/IjgUyoRjDUtNRcdkKXZj8yIYlsbYQfFjm
V8O3fA+xvqqvap3uqYJ52gK67S2ocyP97cGmBhAVRy9Jn7rgWC39O0EDZbrT76ssq+7TLYdvXpgw
WeQkhD29DTMdOltuHFke42WQCH2oYYi0JX3FidwTACO3SiEM7i/5ESrNkxHOYn3zEnYD68AvGTM0
1Mhl3t+wpNnLPZ7VlJIFp/cvYv1GLywj/NUqsI17WI0nYzkcIJUl/WlX9HTUcB+K7VkFjP+mtNOI
9N5/5eXkoUlNyno7TYmsQd47EYrOU0aep520SM/DXb34sAtAoFyhNbU/voM0hTgQojgCCj4zPQCj
zEyISrurPdQVsVHELwA03gakLV8j9ZzyLpsHcn983Y4YsaIiEH1ybOfSD923wv8vxYaGyECZ+5JA
HWMSwt+rasgHcCfkMuzmkAn5ogvQ7tgo30heU/XxRwKPCCVN8CbXpxC6Ivvv8Ro3Pk6xvbTPlQ2b
4pVO8FZpp4FxX9JnNLMuQFugqaYvdBJR0gxDskDlnIUCa6/HY9cCrKPKT9Lf2HXLSplZc7QgPiym
i0kEc/rSFmm1vRMGtluojwNKUKFPreSjhuiAaIAwxlE55tgPHMVfoE05O/958lyX6pRx52jasLJn
ckmsvnrr5neNnmkiWi9E1gkDcqDJTBI29uwcMyzd1pYamIHGbI+ghnbvtYAVk8AyyEAYJttp6Ioa
ndlAb1W8w6iGZjsdeuF3sMN9vvvbRo4VJQ2M26ufyfmpM+hanVur9Dt6MC2n1QZ3WbKVws3tCd/3
LUSwq1pQkXUZe0Ajx03v2GG6ee6sA4nemk0zw9NRSjZks211kZWhtH+Gy15B4lmvv03jZ7LX8QnP
CAnwhV1pau/DO3knc9fScoR7RNQThF+5CHEon3DIMzwR4744I7Ujz5M5p6o2kIDAGN8KcnnhmIoV
zIwP9jQE/BiaYNMImUwlAlYil+GINWWXMBbPI7aoWckJO41b36lfn80bUmiWhAXtTQpL6ydqcM/o
JSg1P3gNrbLWdMY1hW00bE9dFnCfCO8+QjJ3zgsIuK4FbGY9pW8qewEHRdBVFUdnNJNUv7/k3OSi
qiEXSvXmxTEJ7O+1iwV+zv2ifVvPpJdu8YIQW5AC7CPAft+N9pY/dKWyWt088C0o27kLisE1GnsK
6JiubBi0KidT7nnG3x10S3ucUGrfnG5s/HoGDJ0O9RQHCWC8Zw6lp+ykVeXU9KreSF4wHloa8anE
Q6xWmLCvNhCMLNPq9sJQRZaobe9aAh74XfS5m/GqIrU5wp23ZivQ/Uvk0aJe2RCcvPJPXH37Tgte
6ZPBfxZTfX7Emfe3G1caqR2RAZ/qNl2btbXC/RoQZ7TuNM9tn/hBtbyny2yLmvV9CBv+n/Y6MCJo
U82mvWBLIdhqDxBkbhXifj3CVLZ3MJ764NJugp9fY3aRr7v/psweVR+MIjMou1cL7hC/4CIfEqux
ajgjH9pCDiCxOglimg60hQWhc8Na/XyKqRjHskcgJrow1O+WcCsnO1J1f2uvnN5P08fd5pfO/DAR
EsjDjKuqMANGejapJIEFmxkXOH7JzNxpkPyfbZHWZao25GzUDVw+7DFKA1FdyvL0mje3N3pCdJd7
oUQk80q26/VFEwPqYbtqBz5Avhx5v/OvN+jBYfszl+oZN86lLnb5Td08M9/jC1s0RIhozGFr/9Z3
etn15m4ljUOVLFGsDDJ5E+uMWaj5H34Is8NNX6YXaHgPV8JNHX64ClZDLYetCthpw6dCLIOQwRez
mWjuD68JLg40IrvLuAjZAUWp5T+Cj4aP+VnVYU0sozNDb23LfjqA/aNVeRywBo8TMgX62rl2tOzI
WdBiSkyAvqrABLopuxm0FMu55TDT77Wh7LVejCDqlLD5h00KCnEHselrqPhG7O8dEXnrZsSLKflv
QmKmD4Myq0lsqJgnhlmhr/Zgh7Bfb9Dx2qhzU4lebM/C+MLVA9frExVCdBsaUOo8PZxr2UPYD1xz
nHcrYY7YAXi7Z3PU3xeaqMqd+sKvKWcKR/YZo+7PvdqVZxZPbyJtzr2Wr6lR10KUpMERpnD2ineP
vSo+c92JR2DR8hD1eQZ4/u4H4wINTQuM78O/F0A+kZ4x9NMt4NfuT4fCxngg0Mx4zbbQlyHoQx0L
CoCY7iOZ9CtthAUnRd6RT7oqW6wR3Bw4Uw3br8dYyNebwGZUGHanL8KKhM0/xTYjUaoXm2zr6Dyk
f0NpROlfHMrpLP3aX89nOtHEPYzst4N/CZC7SeC4V91kWgzcpD/H3Pa9HPeOAcIDORamOZetdrj/
Xv9nUYnyPs1F3ZTCy6hPMQysi4IC+1URyFvO7kB77hjbMUxd6jcEjN5qEP6XqJCuSHvHP32yon4g
WLqOMExNR49PJyP0OcOqq4l17quFT8yjwV5BjGSt/880tg/6oAeopmtI0cdZ/ZMcj45fTaghs4R4
4Tp0fxojbrU4vg/JVradNzDrWP2rdy6/PKeeQg9Hk5v+by95xipBWnrVxpseCh7MzP9pM9T5BcYA
kpIipQoE/DcgD52dxjMwkErAndCvlaKWv0fBBjN5HusJHIj2g37bTOUdE64jhoU8XjT+lgHKDhdb
WlOq9Zq/NkJYAaz4//Bl9sZg8vhYbUWmJGK2V/YZVkvaQhtfgAmWPz2YxOGsIJOILk95d1IqECHU
lh/o8nP86IoA1ORu6VUZNt3z2jN57UpDT8D67BueslIudSoVw9LVEpjyXsSfhWKuTgvsmYw8v0Sy
97aGSHWNStqs8hCkUxyMdVfrGMB+OewrPP8CnXc82qE2AoaAlcTbB+eHxFxFEKEEpGiJU1xE89xn
HBKjlaN9eYnMOKDTQmAowZfibt9LIgHSqiV7zO/rS0CVQY7aA1oKFvCNuK1bGNKzHGGMVvTxuoOW
NocTht/EWWruIV+XprDnqPWsxNaqSsw/qtZqNyBIpmEsZtAw5ohGTeRoK2/wenlW/DhpKlRCAylT
h8I2YAkGLYDhniqbAV3faL+0jgJxFz5leHF3qPqv4gwSkjzQg/nT67xUITZAjGW+pQiAhgRCZrXb
985e5psA6dGsxk6WNmlQ3pRjVOe1MBLxbZUF3aIukTQF/jRVRKg5fsBLOxFPJtLX6wvdknf3LmsO
dTZWmkVxCa4ryTtK1itlMMK/kTdRKSX+vEfb5rNffApgkUbPC9a0XahjxrLj9kRw5S0WJ0fpR/sm
lTIiuvKPiCmZDUPD+erVgWk1QyhshstKCbFR0hctEVjuflPDaiMxYehtvQ06p6fJrHyJv1iWCoiG
2MDb5z/xFmywjG9hg6+kjdcCPe9zxcFw2oEvDeDpgnSuoWV5m+A2fhq/MXj9M3BwWxIjZ6rFtB2c
s+U60tpeK/HbkoOpGTLvhnfSixbpUmtNYrFFhYTnqEay6h0cTI1j7EgE7zsaClGPK5s2CkSo1X8K
bBy/0QyPWYYXxvIR4JbijlSPYehAtyU8HEFBOnWvKr5LX+Ub2nM8quVFpn2TrxIJ0RQgX49cxkSo
+LmvjfOlBBFXwcYbClex37s9AJmb0WH1NKr/oVyp8EZaawz5QA/0duX1+X7EaOmq02W5vZ17d4YF
EjxirVfUg8bGEVGlA1pyozOw3gspmYmZxJNxrLFhcG3LtOvDo9dcQwd91zsIxdP8y/zm34rPAaiD
eZmFzmVoJTD67jxbAoDm58kaB3sLZG0AABQaB+t0C6ASa4FLxhiuafjCRL/v7d8Rh0WonT53tZ3s
JrPs7iW91BDKRRUnUY07yq6caUvcMv/hROxWANQfQrO1HsN3+N4fORibG3fffxYMzU+vEecIeLx6
vmuarVeGN7MaveIHxSGUAcmnGSdFUUGazZLpdHmRDObGYTRRK+/UphNqWxtAHMQvzKypl5vaaZaB
Qvuj6nEgx9SDCp7bRZfr2jj6R5yR687dZauAm+dCKuQDsOXZCPA1ft7AIoBd6OsxW88ME/gbUqPX
k7IJkvX9cZ7pqgdggaWoE+odl6PhGo7Den5yOdmnwaoEq993dtCbpmzsRJplzfqSRS9l+1R/Is76
jrwQP+6CYaPxJ94rHiXzLtILn8X5P2XRPBQvNjeF/H3k1binrqxqyUpdYXzE5HcFcE3FCyv6P5Jj
d3a/rf6d8NfPCOhfMXKvMXV+fD6VVVttkp/5JDs4If1NbMrpj8ShvPwkh90S2DjS3mql6zCyDrQj
GW6F8osDL3etM9qkkT9Vd4A6TfsDbLQU+Fo3glD1ifbXgoi+twLz2OTT9UHN4KnZ/hKP9kCK039U
fztzBT0nFzR/YB7YIr4JhlkGH1LuImeab+i8na1k5HQBDFGWuQd9/6t+PzXxn0Kyrdn8pkLuLd4b
Ykc1i+E9Dfx/1gVe35hR2mwPENhjFDno4Ap+alqUR93Ta9fbXALB4+QASnM2arxM2bmqWWoSFEkO
Mg0gouRclczQ2egIpMjyChAR7smtSJDSsTheeIWdNk/H+7H40cfKflFhBmeoATKWQw==
`protect end_protected

