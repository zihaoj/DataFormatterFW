

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
n/crKkuvxtVNYWfgisE/6GYjSzF9g9fB2HGdsJOT9O5wSjq12v6FMaUlD59TMUEZpTr+/Bb9cd+8
veM8c2v2iA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OWGsJPD3/DEM2gr7s6C0VMwHhyyvICHT4ThnW+pWsMA7b2hLKa502Bjb19AapmV2/RQfvnuLOi/i
611PK6mddaudBWp458lXWCSN2vlmEQ9ylT2l1+h/msF0pH3OcO8G/zOujtc+LLe8sH2p/DqD6lU9
KVbU+IubVqTBYzDXyPs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Unue7WtjFePi9ibPNeVwg6/qEyfqiIC6cVVZEqZ2SYPuMyu9YxP6c1ZJ8YRi3D+EjlOB/Fu2QV8K
UtU3Y03v0jmXHYdPRvvNe7TCKdwTyLS+HJ4FZKgi0z5aBTQTx936ml38iRpH+qHmDR5L9n4Q7f2Z
LBLP4dusbqXjmjbEv/1rXeOa5smCPNByeZlnLjugejfb4ACipKWslrbExDb17YQT/Kyrajd5zZ0+
4zyOtUEVEValJuy4cmSGQqmp5RvIqoA/iI9dI+Pd9vPoo/jweFoO6DkZIKElW/HmUkSJCdIIT8pK
uXmUGsJs+MdUuAMTciwPp10k01Vgp3L1UIetTw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tvKnlAI5F6F0JFxQmEAUm7fNYsolxPrPmYzFHyc9XVhZoYU40zAvIJ4IW6Qsa+7NGTePcYZ1rgdX
1j8Bv2d71pUYj8z19+K4acV6qdRr0DMuOmbmrCvhmu9uGkGVvwdmIDz2YPRUnf/xU1gjoqj3i9s9
dF8XA+wk4d5r5spWCY0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l3Nkceyz60Swqni5TklaDjQbMBZMAr4VHU3mPKUNk18dEnIO5YQFbIHmViYskq2te86WICthxt6R
zmfTIh6MWckD6AoFyspypNvna6zT4+ioMCxTLhGHCmUUwqx+RfR3Wc4PUkB1n0nY+1dHRWoJDhp/
ozzSOejfsp8uDb2Kazlt/YkEdi+VSMEXMZ2sjhBv+SIc2fkJuEA/RZeXxxdEv7l3jZjCZkECgPSL
+BEGG/MOE9twcjcMMeeprXVpFu3huS47589iBVYIyiOG4X29CX90MXKrPpYiEmRCUkpIs+7IasxK
gcgEJ7ymlZuezrJrTB12j/+9BbpwqqANA4SlLg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13104)
`protect data_block
VLIH6jt37kKCsJkzaJBsJxkZf7Y6HhJurDnJywE87xDr1cEmYkY9HvPOJ+rZd2x22VeMqyo3teXH
Yhzjfc1e4E+fTqcKkADZqPlr1de4EVIF04OL+0ZzwMVhGeof5J+sv8gUp48OEnVZcElDEki2NdVJ
lJOGvvZt0nzouYrvNpTB6xzBv96y1T+GvPPrHryu4EfCv9Xu+Kcm3xy8DuGYJ8VxQnfXNXHmjJLp
yM+o7Bh8G5UC1YUjNB8l/1orBIxk5rMLYZveSUQXJ8EINqu9mYo5s2zWJyqNU3nt5uHLlTev98IS
zZ4Nz4eJUdI1qtXX9h0mi5qDClIVzhAkEm2Z8flGs21hAD3lAXbq5vq1KPPOVieecKkS0epfqN3O
21ltxd43Sy/khjstASc4WXVhGFU/UtXroeMuV/jVkQwHzHy/s9/ufiIhwVXJ4WX2jsokhxZ6NISJ
94M+od4nozkRMoN/auuLVeWIutgUQoAmop6QObtD3vw6LNfbot57WP5gBszjBsMdHf7k4uN7stc9
uXObExiCId6dfEI+4kyTkmzrqj0Z8vqOJq3P6XEIlRjQDmjl6WxjXqb3XDcmQZAlyi1ieg8rD+5t
bpxNlGwxmDAIZDJH5DcaC4fYZFUNUFtUJC9fL/gU5U8/9JDzC9gscSKtPMvNIClJ0BQvPGrlquFk
+U3rrIkeBGPZpdLZ+cPcV7gqdK5RVtHBadaqzuotXtQrBrGkIzCKQo1cMLnucLTSCvxBFM+xisWY
jWvxuW67cSEvN+P/cnPlAZdE9TPfrHl1Kkm8t9zqzjEr3ab3HcXDx7WHVg97X9Zre+O25/RxhA80
nEVJM5C8dsCovofdQsjBOXzEif6Bib6kffJpLyLf89p4pUGUD4Csg1Or2MFTJVFNnlRAjfswMn4O
yguAlHAgC/fY6SY2S7BOE90BIKjFLZR86I1uZJNRUKlxjEbofxV2mmbcH96J+yVEl3EZZ+NniaQk
BJPKfvCA6UwlJYRTGzNlz411riceI13m8kqm0T7Trhym8BlVaL6v/HAN0xKVYb8zcTflzeHH6jVF
9TQNrfM7yIhDY/nTBpEOPt3C0PJatQFBbe68Wa3fqDTmZxiPY5w1cgUzQZUee4x7QdJ4hLFPQuI2
rFOEFe2cACl+yQLMN02yhohLIr5zycwcPmG5VY1wYrPbF2U6afEzAI3O4+QZSiFcEexuUBNgtalk
61smLyh+FvRHFnkn8rWKDoIQn/aeOVE+lYApanZ6qwhWkCewxAJan5vGh31xxj27M6LKUEl8YIFE
satVBiTrReEMeEY6qPQ98CNaVHzSXRVBvC85GKeNBTuPadEsEqZm68/wcqhkgfs1Y5C+uxMTcQKV
Aj7KqCA20B3yDfp35LtYt4POxarvsIOhoMh5nAmausyXHP1I2E0VvvzSbWSHjbLjDIW03ZXJ3G3h
wLgKBWXRmthxajPuujt3beJsuXVuONBtLzGFu+mcQlLi768kNht5ZN/XtAIXpsZ4GA5ufODip8gd
a0Noim2JdGYyUAoqWlgybGnFY/7YHAvbMkWCraEqpKiZv1quhmhOOz6Lix6u35VBSKmTfJ8ylF1u
8o6AiyN0HK61j/aajJTsgCRIuNSsRAhvY9SoA/PfYeWRvOoQlObmLY9wpyVrprexOn1F+z6wNNJc
Dvc/gFzCp0vzhvudx2QheCkKN4pkg37hO7SHa3cFpNRs8yyJMO5oXaJixHv2jWI9U1FoZU4H7olf
yNOOeBAKIXh2LusJgvCISD5QpQ0FJPGC+IXxgbSnfCEw4R3iFQSD7Ax/A9VoqdQpnYsPkv+NXlrE
iGfwZMcOonn48YjKgUwBPpZoghH8N3DLGeJ62NeTiqnQtMw8uPlejxhyQKHyv2GN1Mrtoaf4PE/Q
MvacpVkgFtv/E3ArPiQCc963qyzzBwgLc5SdCnS+lbVyvT6rFWu6v+IWO+rJOuTRplM91b7MZqtx
WZL1Ft6CSIqLYTpslppTDhI+kf+yyeL+IqzhUTkvWJC+mB9esIqMEAc7w9mRz/AnAYC0QO+cTQ5P
HMtiYYNW6OqsIMyii+MrqyXcgW4IZiWm3wHH8mbiIi3MgT9BqsoAgNKr5MoPRe3VblF3acMYkIli
G5UJQOvtcUi6xT0DGBrV7WkM22F0sgytTnd0CRMUsRxhzdYDsdk8aEBd8e0sx6RA/OPFndk+ua+6
xfipJ/1KQyR6rpA3aFQlY7vXqdA8J5vFUnGX9fZQSygsNhluJFjGj41W55GRmzbJpqL6KHbr5Rx8
Onji/VEiIauJB+mJmXO81RvNOxi5cCyW0NXZmR0wIshLdzLVrRD1riuhftUn0yoQfudjsY6uxEhp
LNFLUOT120qMr5hExTfD6LF+iYFzvsL2lzz2DTG0ZoqkJdLIvqErWyhIUFZgdjSEphdBfvzySEV7
HzBCm7XF02ZVvxKxb1nysrfocw8joJBtHBErlIfBvez0GJlOFIYRhzE82NXJwhUUCvyddohyXMq3
qUeiVc8MJqg1acQg5ksFXxlsZML2botyJRBjQGjQCs719l6tJXjzWRu3MWCFMICx+2rvVW5+SGOt
uiIcMQndgjoVmzEALOzcc46EqSZpuZH+6VvpRPsc64KKxZqomZti1rOjszmg6RqGJrsILXwbGU3F
Lv6v0pty7fhEWK1dilfB4Osmd1S+eHrf1aWg5xYYLZ0iE4xjvkeAQvkPxgwqvBVmy92x6P5KNVyS
WWzbwZjm5qWEemY7fbaTwCjs1I60CqGntKOZS7+La2ihOcuFtqo3rlKvbPPd7gQR3krysa3qL43Y
DCqP7/zFnRsi6Zl6jcmecKX1kBxxWnhpXAvnual7Vzfo+wZ/wHAQchoKDqNNmFhc0JpgZQjo67ci
gsb5lPEAmvPA2hv+WonO9opYTxO6MZXNuQpywppnBRcCAWhT7VC9h4yGAc+cPGIv06vIXpKcs21W
dkeZ83OSLUZje8QW9aUzJqN/sT7qRejJ05vPEjyHU9ElsKOT3WvE+aJ4Be28umGEfPADtoiOio8v
AKiNgM9Y+WqsKUTOEXEBsCo84Is34gJCuZXTs25l8ktnEx8nrhV8e4GoNKSmr4AfleOW1309ctAp
55m/esFRJQgjuORrTXLwxsFVpLh/IxFiEjZmMfuvOI4oVxmCDQhOpFG0Pfer2awmYpxtElvgAXUq
BxrTp42J2QN53sErngi/dcwOmMp9MysF35Dlc8GZ3k8/9cX5HTQ1Y+pTMmPX4L4I+fT+om078JVy
lD+FzPUVD4IRmFyMOOIykzOyzTKFgaiaGzB4GVkjDRqqyGShPtTUk057QsO5zRk3Wu0cDIfaQ/4B
jkUwRnsKENzjNXgj4+owT6O3RTNR+X/BzBqye4AfwsvaHWSLEbRgHPchVhzqnkmJOCq7TPxIbUzQ
E1XLZxAmM9BE0ghq7ZJlYJDiGNiuKpCKZgVEquwYGHGUWTiqmKD3ZzJZdgniRGBlpIK0NSvZS+Ro
JAdqetpJajD7PGViCEC/xv1VV2XecXBhYwYDnx21KzA7dDNtahUDq+R3RifJNF8xJo55gmY9WxXY
k6NTAnxMjpF0b/7lX0BlW/2UQtQlMN8QBAi+vUcUHILz8cTYrrMxiE7+H4ygZ4vP8830Qs3VdZc4
oGcvCdQcWqOPXi9UMLnxaR1XG308x07dA1OmNoAY2NHpHizFY0eV1go3QwkbPUeUb3zmS4qvPIyO
JytVtiX0OkapjOFz33jQVf6gXPsHT4XLHJUThyrOnESe96jhFZ0+qlN4BfSzS6xK62X1SI2O0i6d
LazdeggvXRA/1e8RTTnRFoq8SXbFeBPqn7G2eLvyXelgoCX1nJ8n7JSZkKkQVHk9Arsc+yIvhb6E
RtS4dbiXoY5jW6pzCoFWUoEiLrOSYbtJx5mEPxP3zMj5PXJrLTNvSRwPJ13+y2AKduZVECeV1L7z
wvCx+nAsnEillZdjHhH/aJ1IQRFY/gmnJ24VvZivqcF3YHb9XkBtOOyroxRdcf06L+90blNMDp1j
1YXwz89b+fQF+9kumNm6qjkVROben3yalW3Os8iql+zGllXGvj2Qz4ipBW24OaiBZ252hCXC7Fh7
UR1qFFer2emHSIEFClqz2yIkrWylfewKo9mMRI1hmjZv73JwTPYjBM/GW0PSmVRpsltduuoxG0UL
sasmhYlWYJ5m35C/Ot1WKFh29J+lF8bj0u/ss0OUxatJkMnk+YnCzjvvZ3CDZ1J3iqWmKGvpPZFy
ZPNspZJUlZr8LM6GZFPDO/nkt/m+Hz4R+MzzoWfaM4qGm0z4uWfW3UrRgGLHb4VEFAVhxk/9NWge
NxfUq+JvVsItKmYaPv/EI/P4+TJcBvVnlEQ8k/ZZfmw0pXR5toEZjDokvHMjvanFLPY2OA+rT3aB
63UrY/+fPXMwEtP/G7KfdwW3VNNS9BePu8kow/A1CdSwk+y7Z++WhsNjmU+TB8D0VO+3WaHvLWH4
N1daQzLEibJNcaNGpikRwG0YFna3epHxwf00RW+EJydy5Q3TizOHhTddKPOLKsr7vA0FtEq7BsHL
zPa8we1yDhoHQHc25ETQkLbAWML9FxzRR3h11uNjZ5zRZwWEPNpX2h3/k7BoIXoYTycohvQ3a/Ly
jZfHi4UUz+DgcVFw+z/xz3q7QZnqpo7ANb5asKBMkVN6o+gQD6yHjOFjrYQMjU9QfW+yLunClcjA
BOEH0dxkk58suIG5BLnEw5t6+kN6WnQqYWAkL9QN990kXgaQ4jbYf9ry32ShcNMl2oUgbtltNai1
rkbcJohPkVmf2Ow/0g6mvs8nBaWuKjOe7yewgCiK24ZO52UIq3HvzMOdUSSclVjXMB+CHS4nbBKB
qRz16Zb0WeU6aJG7I2hn9aWlqF/au//LDspWkHh25ENVuQS8Sgh/ICj/WrI5djj0hExgr1109igu
5T+a60U+Lk3jYVPBTCd0G4hyYd3nEtpvV2AK0RfHprGVUipLCSMRzpg5LOe+JCDo0MGTEjJZg9sp
Bz8yIGk+URrAxT3C/JOH6KzXRSJDSBZUqSPwtPFi78Vt7Hs6nG7swQdbQIj4Zt9cWx3NApQHQE4D
jM5jpYJLa8AvH/6MtBGZ9f1j51GHG0qjb+Mu8sNSfwtBqGPqKZE9tcxyHEN/4yZXujmL0JQRT9i0
nXwHaLMvb+ZZ30UqAEJiOsjc//1zfacmpq6WAEoiuJ2YGGk1Oo6keUjAPDb+toG9/72eaHsIhnQt
l3rjhyc8vUEqAfpSlWqMG+fWO6KWg4SSQZNBVEuj4iVExkwoN4XnITcZvGpxsv4YbDk7Or+goT6f
6moGuPQYzFypP6N5RYzEpLkgAwy1FyTCA2/Nylg+t/6/SP9tLUULD/CzT/I2TL6Bk5fhjDBDPpiZ
h6huLSuvS2Tc4iOSxw9l2A+0NXNmKk5AMrjDT2zTdJG751BmQnjxksT0IxTKiQqffTMfGr9Q+x7m
cuVraDLpl0c9vXHDJU31L5u9+R9ejxX9ien3JiV+yTwa4iuOxCERTf6OEM5v3fSDV8VJDMIBLzGU
P88E63OrX2MpNi8uAmJhXDWb1DkFifpC61YUHrxVLD+ELTAR4ws+laGmS3bv6NyfhzCe2OsbSEiI
hprawzM1dNPcqar02MTxYY6z3Y/RvbuFa5XB9IyyX9OR524Z2pJ4BNyTPLOZPDcS5UDs8vvlZUXF
PJwuuTtIrdBWbaJRfexcaq7TAAxGmZsO1zI2UGpW5yPgOwD6G0E9WXYp0iZSkeF/9nI3BD8qCFZZ
pNR4yJEnHkD56DSbUP3pforh7MAobCtqztKqxLbhghMEIEt4p+xbXfwmH++uIt3Y0FDd9THeyHT1
mV92Aa27x08/TUKiE+ZbcYYGp/gsnv9bCRWzDX8cezej4VFzbeAI1nN+3CJ5DSSLyMyl/xR38OCV
mBUKZHVtZu4TkkVPr0b5SWe1Oz4j0LkP9ZA3SF2KUB16BcLiTjHM08D9JHvjO5KM5sOfi/TkKgF6
4f+hfWeLLo7uVzlbvanqw8ozWxeG/uJmq/u2fuCJUsVN1bgmeqNDCbWIbDcBbxqZ2TmdDMYgcxHs
Yi6sBDYbKWZTkj0Jgkq4qtbbFM0ExaOnfPBhG7M+JtRYgujFXZoET6LJxdtZxpkX3o2llfNTONfr
gmr6vTSkv1poX9iVDJD79VDgLySBJp1lngkM0yGX6dSqusj4yf8llarzUsTOCfA0Tr1Ni6c3AKSF
Ud8W27zHvp2xGkK53rrfQP95fgGFO3q4QY++7FdaFXFFhVsEbLaEulQvgoc5xwO+GoNzyKQEoVda
woGastud5WYrMekkHMigmEmCn4kU+ZFPqcNKjiVjQDCqzxJMqsevqjM0HTGuyTPEdxyW2ysJCvQ4
TAp9R9y0EG2jScLG9oAqN77EJULpBgtkZyVCsWAt+vIU8pU5U7YfHBJiu0TopiyA7N9YThaQFxYE
BLgVey4TxTcZO+RidtV2kdYczI+pXcYLScaUjLiFma2IU3RDadMRphPRiery8Z+L/WAR7ZTAa4L3
/Ni8UDH1lVNUrMq1Wx6fq/K3JpkGNQQIrqjRn3EOnf1/3tvufFH7NPwMmi1SYojKPlWCal4irxm0
qHagHFdnshXxr0rNVrteD8iKlDfH4I42BdPuGQxVk8otJYazPlyzOOMQmRL4fuWAgruTrvsdV3xw
37Jo2RomWtUAVScbNlhD6bb7VWSd5q98HTcpZLJI755XUrRS+9CKFqxLIQe2mJNmD1PN2eHhmlXX
UuI8kX1IUD+7s8oGajNlXKRJf0GYNOUojsBnEVPv+/zjtuC/3wZDntBT05dHD2rZ92W9tJB/hHES
vaImGVyFAbNzXNA5rrQPNsPEw21ByHK/oo6TiQfkBN3NEjmp203GLqLrnzYgKBCqcwaWh0tKfp/U
VNS/fN1HLTVIOzg8nK7ctHV37xsswczHp42bCLIBTqTocBEtBIx2YSL9dEnq84Wgj0oiAN4jYN+1
Wtr/54tFdac5eKjBoVE66jxdPHplAtzoSX674C6JGnZEu6ObNJxNEs8401EyJk7xViboRywWBGuC
SOh5pLTeBart9aykxqggjWHUNTKe/WESuouaR3GHNoCG9iTU5w/CdKVs6zH7I+eMNI+YtV7nbK7l
Oqkgj/OqGr8nbiueiF4HwhODfTfS5VPMI7lON6fIComyR4Gpgu9gnXxAxBHI518hUIzQOYx7m/v2
PgN/Yxy0r43AeXXHDQ2sE2ybWiRrUPjRLcP5MUw3ACET8KIA6UyAgK0P7/upPiOvmrK1HmBAx1cz
/sj+AzHjf/tuVpiAtbSXfrTJwmLAX5oAN1okVcZ2fCJO7aawDbTxhF70k/Vn7xSmYDQvexcBpF0/
qpPuMuvHgGb7NMZCbIymxeilDMuxYaWTFb95pngYGGbf0hkC1TUDpVvwocGvMeLqpapWziqQ+uR8
GdXx40cIqFY+1IUIucGax5+0YRwDCUtrfrjsu7ppMjLG0N0S5KJlOxzaEdm2Uh5cs4tlGSHw+D/w
+8AMspFRmqGVEKgVnedNxGr/4H27pHQpwJ+PrLtcN+0XQB9/+td9atkQrDaMqx4hSyztMafDfynG
3nMj24BCQxFvedxwOFISqeIJcxf/SyutVwaQlGRd1mgANMFOrYHG00PtJ8B0MkuEyx+V81g/reze
EmCBX5sw28xHPWKSSCC8FTazKqESYjo8hxHffP4SClRPJzrkXkQXuV/ZAIPZ7hW/nWEFONegnIcl
+49F+ybPMUu/e+H6AV7S3tJezo48vT6MGJc+F4D1jiermNAqeX0U+LmxQ+uAAzQ+zUQ1YuHq5nib
GJ9Nbm0uEzO3dXq9EQ7Tr9mA64VGHPXaq5PjLuiMnMeWztfUNjA695bpMIoJAEbOeGQXIUmn5CjW
aAWCOYNc6Qn+DxlIGmWa8WqfEjyxulG9pmcbvObgH8Y8R5PCaHVfYBJYu272e5ABwYBjGNZNSGAr
zY7gJZJm++pkS24lwZjvSMDNofMjaSV6DYEdzUSFjB0sAqygi3g41cUMxG5bGfam2iOvfsJuJofR
rMojFA869n6FvJaN2AFs8INGvix/+w39wj0gCd8I7INRse+kg8AtaiibGOhIDUS+8kMOdtmNR8uz
8G6YLSzL6kdOTQ6XAZ3GpjS06zlFRNJyWKGnaljCJGNlmAvUJ9F87p6sCKRGB2nXwBbaYuJnGe10
QdQsERQ7oIaAFtsA+hOhLx3LOJqwbjptOXM0qaCmyBjrGZgzCSsYcRkt29VpBmPC6u+Yb/cd2G/4
PWgJ0cNVbBJUQ0F+S4OzWJDmURTMW8VGzc2LZAyUPgpNJyCz4Zk/WV5AFHNH1Hyqmq1V9wGOiuVF
bqpqLDCOfNcQ1ZrZRZoQhfvq6ll4WSnhNk2P6qUhIsgQchmvf9/IBmDYRHOC1TSxMSCNZmYk1EEy
jMBaDquao4J0bcdh2sQHPNTP9QhGIFAKvLLFopZnb4pELsTKMnN8yK6OvcnBr1mIFOZeO6PPSivf
18Uo5POpvvS5ThFrMc9o0Sj/1tgXDFj7fzth5DAQv7bw8fPKKHlhyGnXYVaztjSUlVFk6wZkdbX7
mpsH1EMfvHbdb8gjO2l3zYLCdALh8/lkBR2uRBWwAconzid//z9r1uVgNg/rAueNJhXYBsQWrEFD
htiCAFMWttyLgDQ3ZJjsVihSQZF+yNa1bEIlR5LlArMLt+3taMapz7Z7JfVKtNliY0LX8o5f4/0h
ZjKJwZiiVuX9c/UA3E9gQnNA/TQtRTmNRZD+BYugG93rOuwhu/dMpFNKofdJdKd0GXz6uxwwtMUs
0aNHEVXVHC6jYvPEib6h6s9AXKSLsY+swpqmu0QU6+Rk5sTasTGDwt7r8s9jOjKaCeM8J51amULL
0tYtKdMmqd5aFE8VbxutkKD7KgxId0CbeyDmP9fyuabzuposiL32gcsgnYbq8F47DwZoxbPM/lLu
gclhDxK7K09z83kA+ZsIP+DrGr0r2OOgOtu3QU/FtYgiOOru6A/pTtSzrpFaTeSQnJYM2cEPubhJ
NXJ+tjOZHWwcU7AlK4Ch0e+N4CN5SgZz4Jq6ktv74UmEhFkMAObx6V10JaNHPrQObUEUll8iegLN
yF2BHSDnHbVqnAYda3owcuUtzab+p935UsDIPPbmg9oXCmbdWiiLdx1hWhaXiYuqUUgCU1QmQwpI
MEaGZXefSgdwlOUC+ONwBXsn+dOuMz7JSHRsQqa6gsxUVqpotGcEIBoYkS5DMuLolmNz9nxpi/Qt
xlGN6MCd5QCVuZyAb0Oig96FV6VvsoyXQjy7/5DJWrNnmHajT/moKiZCGw5BSq5gSA1aX6Wo9Xwk
hsCIi/uPOHp+BzKHI6ecS+cVV/z3+Cct3lmSDT0oeHqDJJgo/dzQUfBClmW4IcPm2aSIfB6bYqzO
AXO9fCJVRLwxZdPEPCe85lh4pcNuQ3v8xlxE0LI+tXQxjRp8pDs9SOZgIljr1l4YR1egZ6oULN0Q
evmFm30SIqx6xK7g4oFdHISkpWpbh93IDrloFMxuDkDT6hKJwyra/A7Rkgr/2AFwgXYw3lnfkDTj
//itJJ2f+aX/NhpNoZgPlRCIEyMdK8R8T8WW8nqTcSAYRdNub9wTMYJogAAuhig7U6fKBrhsrgAc
MO394h5DL7DZnqgNc5dr8Z/Vqo/OoexGl6RmI64dg5PvCNRIqxzVYc5DkP9nurn2foqaiOXbHs2N
3DsmFXzx72mUJrtMUFEGmoOhGbhkliZWkv/VdPJ0DA01p8wzCg8oGwbZFmypuDsYTT4fKWpNTLgn
yzPqJDAgEgI2HNNcJl3p7BkjZ0Cz0zE0hdcwh31WULNjbY33UmJr5y51+u5z5PvsPq2x8dH4GxsA
iLdCri5so+XO2gCIVBAIQhrIEj3d/UDN0xhfRiz7a7tHK/fswq7hVkLRXmJusiSjFcqFNZHw92EL
UpvTUZWusWaQaspumP6EPj6tXa9SgaHSc6+2Um4DHMeqKBZLT1iwQzkUh1CM+c9gkokrH60/T3Ii
7BKWy5MfM7jKC0OCsOVH49O19sY7hWSdB1toWioAqgjWXcGlm2NzOfoGPMXxEdb36R3heB1C4GSG
BGht5ptrxFnyWykjeYj1eGySGNSxou9SeQgBM3A8c7pIZcDqYpV6vYr2UC2RAiZP/coKZefqcvjC
g6PzLahgyramv0EIcuNm4MMl+xB908yWm1FGRjk7CYB5+E/uGjHWFeIh2CvhNuecFW4istYTFkf2
wzuXVoeHvYKEXaM0G9YExGrcOBtgYr4CqZ3CSohRWt0C25Y3Xe4xI5teXCR2T2zVqFkl+UyOJiSE
D0hnbSMRqylRwPcIl1FNfd4hawTU/dHTFsdb87NR3m2tn9R4Fo/adH5saWHscjj4z1DO6sYClRPv
zp5DKQfb4AYgPH8QLiIwG2CoTgKGBX1MKtkHIyTqvLMHniSUURZBTTFgn+L46Ci92zlgGXgUrvbY
8G9V1/V7wGyyaQw040qRHXDoWe3IzHNAzNnY/yElg+6A64hT5OFlWGu2dm0LOl63EzC0OKKuQjYS
FpPxnX392P8KxnHEYKGa6BP2KfLsZr/ZMj5pnNXoxV4fI90F1MkGXTYLyFXJ+cQx9ir+fOTaU5RY
/Ap3k3J4JOONCXyjkEF44d/09bawVnW833FaCJmGiA9tVljOEgLAJcsCyRWnzE/+oZ6LYLW0egUv
6KUDxhHBWUdXcwT9yL/PaBQ9eP2OiBK+aJKXd9pR2npGBf+4sjXxUWLvgohDFX66857dERf9rZv5
+zs/kF4PWg4+BmG/bHxr0QczbZgWOCXALcV5SpYG3HDPp0iyXhRI+EJSIUPTTL2up2cs7AQ9+xCh
sErajrM/FRKKBPNgBbvqc/PVjwPlGNu0SH7xu6Ul+3c5f73zf70yN6L9tsB8xltJgTuwhVN0Gj1e
6+DrVQjbqq032xPippy+Kw2c9aQvFmoAeZnBkL9ktngK6Ism5BCWdli7gFABn5PTzGMercsLwImf
4svnTewN7Uwsv+oithDxN0GDpGg+CislX0QT2gwKTlBwWSY3QnNval3MwUL+oKqESE+epOqQcKy5
TT/8Ie6jH62gGWoMnVS6phyH9BESdhPdeWsrOo8GBr5wvz66EuOsGtEXimg+wjpAw/rcF3xMG9yT
xNwSQRsoXoiisUqIvrUSl1n3xot77W1mJMq4S6yjj31uc0tyAMgK0i3x9XTA6y3CPZLjrzGQegz1
+k1PThzxhSlvC7rObJ4gmpo3H7aSjEb8YePJnnxWikOFKn3QS494l59/dy780mVP6Q8mmhHO46A/
uOa8A/dbLF1Uc9fBZTTBqgH+yYx320j6q6s0Yc+rPfhwAR4cwGWfdo3Jq/+z1cpWVYmgyiPYxViE
/qu/J1hLV/xZHktQ2gAAZRpuGxozsl9pe5vZD/Kn48VnXprcJbTe14iDada9FnJDcbdw22WJM+Yo
cmia8GrACG3UVfCwNrLJqzWGgFxs73tyf23GUMqj+S+or0m/rPEvc9QcDpegnmeZbZgkGYH3QN+a
N/zg2tz7B07yw1b3ugyoXdfbviANUPBTVQAT6+ZepZmlgtH1r+kYT49Wm143Nm2CxKrkL17kBrsu
5Hl6ogzgVY+JgTAEm4UI7WmjEVtzGWM1D4w/QsdgbHMt3Odt8MQKQFh3U4DYTln9pe8hODv6w7/0
9EMS9Tr1WuCrYWod3A8+aYup77+3uUtWTV/PCPqelSgL3q5TtOEGJCY26Xe1/KCxk+6bFqgh3+tb
k2L+WGLO3x8goWUuTzqGaQaFMo84QX0jaFb2wvXnYCgMJbiJdvaVx03puYdsbZBFt0ddnH2aNbQD
fGYyz+DvOJw4JWBVmBHUZ/P07PG98nx/EMyJp3XgmjfoRZ8TFiqiYJdMXpaNZlRAKvgJfpyk1m7D
bj6cCTU3Uu91HN9rjk7/dCVWTf6N0HFcgeNycfdc+ZMIIf1G3haQJkDbWWycidBQyUZCtv8IXqWZ
qNA2Noh8g+mqjy6fWpZlojtBmF6THHFcIG3eUW5GJBk7mZyXGZKTVBDAc8kfahOS3eXckpNb4w3x
AN/N9pTkwTndfIqoWDvkwt1GZ2Q2301Uzq1lQ/5fDQF8xB/EkcSdtbfAgPYweoyJSHmoS7qH6wkN
rA2+e/wd3U2G5mn/h315gqnIoHPL2PGi11Bw6HTIb7LWIs8GP4vCg+dzoQodBYKhMZVr8Ai/Co69
TnKDN2cgs6IVrjVbcl3Kow8sROU+rQpgIy1XM7Ly4VFexcJ4REhDf8kNPV+OOARv+6DPXHzZJXSS
EyvTiXqL7skrcRXzy5tODE2dofvw+W03RXf7JOArORplmBOef8j+4tk1m9/0y+ii5wvHBMwFSPd0
psowgHhIoYm+OZiVx1nGvFVpZV8heuOI5vcxeOg5qy/6+0zgi5bZkRhsq1c5a7yHUxLvGy7D1KfC
jErYvqxEG13HOirWviybBHpEiwI4NvAXGP7HU4jAOtIqZ1e1Jd99JQc9imDltoaGvZ2tL9pk9eta
XtNz3gFvtID49MA5HphsV+gf/VlsRVBSj+OwQyJyAKF1nlid+SQZnWCEHI/JrR9JHnmPy0bEGhFN
S7xKd3JEWnQBkakt+CowzqO8hZs2tfNOJyNPzs6qPtSPgm0C1yemDRgjdPzYIVTBm44ZdT8PGu5s
4mO7NPncO68dMp+VukDkcY3aSgfRDh5Z1M2Loh/dReJh3DofKIoW/fwjBVmINr3Tj7u10Hbw4g/f
tKr9rUU6bnBsu5twfUbym9+XdpmmHjnCIk0jNEDLF/XM5yHL4C+X5GreqgCsRyGn/++o/9XTTq48
MMaVY0l00AV4wQwc8Ks7Mn5G1mVTfttvsnDh8civut2YEWtSw5AlwJ82wBjR3wHnhOz2Gy3t61iX
ElZ2ICNICIwTQKQcXXm6RWs6dNJJVYA2AwKXtU28nBm0wpT4aC9VZm+OHokXgJcfreFDjnVsdXz7
HDMUnBgom2xm0hWkIaZR495rYOyqeLxBKRUUVv6KkR/TRXVWElqV2JE32X4aifH9Cw5V5eXdp3wQ
UzkdcvrMFeTwznM6tg/aNibXSwU89h72lx+tyOTqMuXxkdKum00pcdqgpdTQ6w820K00euyKkbyQ
MXheb6zZLzLNXSwdcEUVlYUMlGarvR5FGU39lu8eBWNsh7WPALkWVYqhh1ryC6jNCMXmI0tSe9tZ
bq9YhxrOlmVX0K/nQdkxCk4yr1YnuKylrkGGnLICSmkN8keEE9bmVmhKQhV0Wm6Z1cU7CrrXxrbC
F8fy5mJeLTr9dOjWC0e7qamEigQC84hdVF9eycLymI8ElT5/Iq9alXtIIYtAWnc0xMLqX4bTgffc
y66G6rQK9rG7iJXY2mhq2IgukfRH/9eip4FRXgUQbuOJe47xHqBXo22k3Vjvn4VA2KLZWUTS+p+D
46MPZRumMsWuMR4ABIkgUBRKaiFXoM4xpEiiZLa/j5Sa/XfF8K7e0LMOY8CCH2vMsQL/lMW3FUqn
pgqU54dmUlUli4R33ScBtZWJedtXXVNuFTKN7aF9HBjChMo9+m8v+SiZpMiSF1qknqkAiSfMSHZq
BsqXgf0OZNSmFoaEFSoAVlUqCReT7HXx8X4iQRbGHVLbgJG59ABqwAp9uGqORAHrGLg7CFG31nZd
BQaLzrb+lUF+Paa+a+uAZfAl6f91OlLHhPWRcpE6N4Y75cmBmSmS2mXTclx5YDtUs8jOPATPg9C1
oy3mKrvuBqBkZTHQPZNlHYNsnuZn1BzU9iIkC2qlX1zUtpSeOw5KpKB1IEk8gjxVCLiF326d2F5Y
snMaI5Tmw05yFcMdOM078VSafx35GWA88EHOp889s33kJIh9VJrFWqodtVceYLaVD59Rshdo1msf
YQVCbMyds/87N7owKeENPxihHWksHae77QfGYpGv6xM3Y6d1Ly/SJwjULuzREisQ/cnDG9DptaQp
7O2kpHHm/ro1VypcH0GoTS9MxPkP91/uoucmEBX6EEuSgTePVWuHHt6lEk9gmziUmj0+YcxQPlxw
FfolvMcYM8TZQFQgCRQCEX8Nqnry9ySpQEmBq8MsXq7nwq/BopkSLTTsMs6Ds0EKFH/Am2lsJNtO
fryQgeUgvU8G++18J8t5L4pinq+fvM/jGh1Oqqt4zYccof6+yNmVTiG7szg+sPxwZjqa+Nw/e9EH
9HtHyDy2dmOaQ5hGUnL07RUOpMqDa3gYq6mlExBWsiA9rOogq8u/2AfspYFOsUVN75EOBUhIsdJ3
dlSFwfYabd7zAms6PXz40po4eb0Kl72gu8HGHt0ERae8w6NqjYeqYgWLILxJ1ePGvRtH8IDHzDKt
VqrFeVId+ieg8UO9uVaBL9iT7bRERHFhPmjTb/32/UgA7kVMAjBtjLcNdKmqWCVRQZBcgERgrz0W
3P5YooFQR7oYFMcs8SDszj6RnF7BJWB7c2WY2+ytPNUOQVV5FyQy75OEeOV/+Hn9DN2DpPYcI+vx
88GQ2/JHVT6/mGA9h0vLHVLGWAys8pp7uk6PWWhvZjW7skXk6PFsOVK48kUF9oZYtqjFnzBDqzRH
wl9uHGqxuVRhrh0l/3m1VU+VGmtKK8mRKDtQBu/vbSh4cuNRfDZy3UtYoXhHjqXcsykIKdaAFQ95
/h218HYrGOvm8MibdoOmsE5C+FVGhTOCgLvPhHkK0JW/qtbai+OcriZ/1oS3lykeyQkDagQtIhwX
HILI/joJTv9CMlNpBtkRjU8tS8PQp2d3qEJ/G2pYVv7ospdVqs3VM8JCUOGGvTVeukcQuCjZ9b2w
TG525qWlCZuzEiXQzChgIRjGs2yqrOwuGZOQDUQHYfyLVQ6dmy+yA/5lhJ5PhgMysi3FR2yHh7QT
0zNggC6MsH1MEdKV48Kc6emcrvffbSWmIJj31dyWPgh7O9Uvm/Lez9C7GJsLL8H6q2hBINBC4SPr
wyeI6ROelXB5JF9vPP9B65az4OgAt/4V8rmxibJITfNA65RaK4PMvGkRxzMJQvx+i+B+uR/srJHY
Qel/vR6AdZsFGff6gUrV43XCto54287eyGS1foW80JvchWkN+w1x1mCF4k7HH8FbnoMDqZzhqsHD
TXD4r8LTqdTQlM7zKtQthH3hFjDglk8wEc1o+wRQq3loaYmBojz2Th9u+oFt232+Odr7WUdk719z
aIRbQyyQkeFGE0qfAVB7NorD/yruVi4w0pXOtWi86Hg+2b51yzZBHwoxSsKPWaJZWUHmBBw5axKo
1duoX5GYsymIY0qDTYPp1a+dhpvoSN2NrvIr1D/InDknxNrAl0rfq/Axkzhx6dbopvVOS/+lM7Tc
wLBXB6A0vojsZz8s6w6SaPkiUbDRsAwGvvNP3Uc8VWGQpg87ZikEWpC8QjRyplkYAzrgfsiHxhBG
nxY/RYroBV6HEDD8oW6BdbPqAu1yaTh3ddOjozZ9VHJq4ZCqZSd9xw12QFVkAjede+kN/g/+ONGZ
J/AGADwCQaaKQ+zYukIGGHOIsqvIG3BJALIZdVuUEgGg06c8g5kHX8nDIsB7fYAD6pUb6Zv7zr1V
5Mi0aBusSePyYFiX2JEAv0gmXOnacInmRbUQewOfBXjWQPyEfnKRmT6OvSJAR8EmEPQKgYG6TI0P
7BydzKbMlhF7/M2IrIctAn4Mqj7XThUVzN1UMnjKNCc4JRV9q9tM/1YaArEo/Pp2He/INmQWHBhP
ckboEdzS6mTUqbS0zPKIehep2em66U90YDojmr2RVq+SBs8Dw7EEk9cnB+yvEDhCYMeOaa73FTBa
62OkK5FTIdOVm959pq3EVcZQ0xDOdzV77N8IXbL0equGRb9sFZ25oeq19TG80VmpWIunkzpTgYqg
fgFo5PTf0WOzjX2VjE8/R8NoKjt3Uj/6fj/mI8zYunkiM3Lvtc89MmCmUpYIHu3yydvIdPHKgvzj
8SA2VDDfBCs4xysuebkIIBnOehH350nes2mhHSSQO84L4c8VdYXi0PYreVSMDltvazA9H0QOljpo
Qa2DVkXumDvjt9zn8UbwSg/V3bxEw+kCE0JjxZPDbxlChC56qqD/JFqICrvWYdp2aMnP1/rGgaeB
W8okRnGYM4BtKD3hyRsZj/fAU/chNozJhjjxivEEEWSjcwPPd78qbxGkRxwKhWfu+NLXS+5+nETk
4MJlGcLuNleJaR4LceQRYCT6C5Cjeb/wlILzRufEex6nQASAHVPtZdz3tp6bjLzjTJjCkCh35mHJ
63ViI5bfbdj5pyvwQoLByfhA4BGh8T0nAGTK17FZtT1UUFfwqMBRsb7xxTXN6nwXQpfWq3rsHUsD
evEdR0ePCkB4/CutnlpHKLU2EtaiKLDgt+Qr8OQx1roWQugI144vMO5+3H3z6iNV4dgR1sk5uQ4A
lPq6LM/1o6cvQTAFfCNzN2TjYn5sbeV5CJliBgoyzORoIysjf9ra55QJIcK/re1we8bFjLLivnpC
PyyjRYZXjOZIk02nKMM9BJ1bntNCO5m+DyVCC6iYZ+uDXLCUIgkwvB+VBDYbI/ehi/b+jl02ri8e
RF8qe+h8DMosBtdJrlPT2c/bs61KqTwsDfvuQ6GFc4V6sKLUyZrjom5khd0ealM9X+de2txXjSlb
yyL8fwbBwu+MQkf7Bpbo5afyKSlq/fp5FoV04eS4Ca4qz+/cyoyY4p4EEU9qgJsU33zkGGJrPQ2z
t2K6LekVrsSPcw45StREzeDRtDJ4yu737ylk9aBE8EEtmw7PEs89ax3dRBPmKlEvUC9DkrZpI6je
l5FL0AW9dFJjDjcX2Xccil/xlZhBY6Oc5FVU8sEXbsB81VME6fQiOvOkeERnJt2WsqwGd5CGY61D
yvIFKDTKamWmaaa7hJzW9xvDC2o8cd+SxAAuyf9UTx6dZ3KPC/173cVEUBPiZyeYvNXGNEH/nBd8
imJqDO9TUSNtg2c89LxHL+r/NZtIpXBCRDh2jxDtRYQKANsqMIbLlcnCgbCljKqquS+6FyFcGfJx
5P0KEV3GUxM0Fvlq+kD7nAvsn8eipnRBWzcFFX8w9gge4pjPK/kMagybAcNOVuixh0gbQ406hZIc
t36v8Ir12atELx5VHTHDEuab2ozohN0WWMbI7wfLcNw6z6/uPut/zPeQpMhyrJXpHqeCKoLvrIow
iB4cxIjEP5oHLQ/ikfLO+yuIGi6ywf1z7NVPr9/JYpm1xn3Zc3MfSdwMOKLVtfr3m6kuqjAp+p3b
3E2yP4ySLuMnoyDVaGfPeWA/rattDcgv85wazqjkBc1TgZyciyMDxd2zOE06lVNFfsmHe4QboK3S
OBgoO+fxqfpFkMYTWd2X/nNjQymXiltZfIWdD7b1B2E5JQ2GdBe4ZN/XMi27Mvqh0p2iUtNgtrnX
9+1LvVzR3IKynocxM4F+AKkashROm/ddA2AU6kwIF4QPsCaWpCnWyICGBksT7ZhKpgQ6
`protect end_protected

