

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
M7PDMVhprUegv3Fyo3UCFRz98q+sdWzXzBsmWEeglSgCqLz68TTTRxBWvnDiWAxjiyH6QvFNzftR
315ukCC7Eg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kOgZhKtV3+N7NWsGkFLT2AxL8ecGf0DLJZTGo13KVWEHi+SNlvkuewwGVZMeIlx4yyHGX8ePwo26
SRLmDgM9+rtDeXD9e9hBwxmtnnCEG1UEc6bZPLup0hwACOabm4gs/W2xqnMKS1VQT33K1lFP9il8
fPCRBwHZ0/H2ByiWRio=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NS9817b/dMdt81AE0ON39/vmj3/3YkjtC+zNieuFaA3d0UmLPh1GugDsf0S52nkHSYSprSY1x+xU
sGJZJzYtFZHlfMOPJHYQL1LxydjrVfo5xifmSodlJWEHxxyXMN77HhWoj9GO2TrZpWKnqQJ4OGzL
c7kSGUKlyeitDr6+aCXZ0qH0Q3KK524PRMUr4LuJUXij9PsZNCh8GaMEGmyJe+fUKobusvByg8Ck
CREKugpY8Q/BdIsEf5r/Lzkz9untCOSig0QXxV5LPibFb5JSAEUrc9gQY4adaK/4s5spUrQ3M6bk
Y6F9NPIkWIAhizJPG6DH7k4HzeI4UTGTiBH/7g==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TnxnnsTtq1c7QSaBdESsWsSrvfig4iom56Hs3BPkANWSL7gztxeRxR/nwQ9Gt2ttX7MAFBJQt/Zy
fLfMaHKPr5+9L9wJMwfP4MGXLmj27tMHZ5+SuZpy3zVym2gn8UDX+DVnvxdMjLZ0cp3Q53Iw4hOC
MzkprG/PmMZNCaij5b4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
r8CDojp4wHpYiiKuiSJV4RjmPUb8RaEZb5EZm1UCHrPGSOyGQcJsd9eIuLSpNq09t5+db3UNlMJT
8Tz0JgVCpFINctYw+eNe0Lt6MzP8qpyYhGt7nz8pHrnCHjq+cLNfhelFmn8yd0GQt9pSyrFYqm4U
obo3Vls+ebUBUB5Zib0eqyW0+NcLghZa2vOhKBuuFM9Q61tTTORqXHBjPDVZqVg3Q4n2Ovoz0FeM
k9VdcUk/aylJpft1tEhYPbQz9QHQSIz3XPx1fmLW+WRkMgd8ni9FOzUsQ9WPjw45KmdmPXqSk4hV
pWftsyXj2ZpKjn2Oiz5HbMVJjw5e27YgRStq5w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62096)
`protect data_block
Qlg3ZPndpgtX9hsDNPduYJGW4ZrmpPOnhZig69ukS3F1cUDEDixy6OTadOcaOrggjAhNx/Ijeaxi
GXo1sberYfK6K/uh6QYF1UzAWv1Ow5cq1cWawcwTbmG7sxIdQyL+HvB6E0SKvEVYQJ0mH5yODaA+
Bwc5UJkIrdN2BhfcutauSBfLJoyXwapxAh5BKYLf16P75usdgif4hASwd4m+seYkGH/SLw3vzCd8
NkkvuB3Qsc52UYTFnKanygvgQAvSLuT79ApLSaAMdkas2lkI+umcAjQL6RTj5EutIq0/VWQMkG7y
lmE9L1OUXso30YtVit95CUrHqicY0oPDNG+ZnoH1KMNiuUSPvYvDYfXmJtksNLyoIJ4zgARToMEi
0wjTl3h0z9wOaGaMp4n0T4X+eUGtZa2lpXtJFUbB8tA1UkjlTQol6GceggZH4SUe+ySanAR2dA1m
zWMa4kpWUPIghnxdJnaLwBtbTn4dceK19U7N0uRQwTwb8om7llknxLH2Fnbqove6Pa6QNx6hLiu9
Nve2qm9KXYKyP1TrJzRroGhQOSBi8btWyvCcNKlEQO194Foz0R9BXQ7E9UZZPDyapBMeZNLwMpzs
KDKu4VDth7R6jolI4mYvoAG2OlJxaRQ9NjSWByEl7tzQvUCUTbc4VFhCsvdznTR7Tz7GWYye4fo+
QvJXdQkyPbrj+VbjyHNDOM5Z9R7Py4B4ZLYTIG9eVusL5Cf5NXUHdT6nvWE/XdgLkjBdnLtXhqqN
KvK+kDP65606h9WrYT+kYu7O1o/LRbZwRLBJjA8BeCM/+WkeRUnowd0li4qXPkAqClGG2VMFn+Uj
pEh/CLgK7RZIZiKFss6FOA/FYqOS5Gr7dHwQa/af+tKAXGxovUqO2pyciBg9EUFUzpczL5kKXyXj
vNAH6MuvDqoIJmjaXbxed8s649u2ej3eJiHZOyn1gBeenxtGL0tDYe294TvwVCT3umYBMOAotr/T
1zQm36kzAHwrw0lPY8vnqBEEfUbea2/+ghqBmdcr4uWtmXzIRl1iJqBCt1eCokTr4vmJxywj3yL/
o2f65mJ+LKnCVufbN4oms86f9V+527w1WeRZVlzf7jJo7v9VuP53fbRSNrLjqKKZ8vZOqEGz9+c9
EqwW60q/BT1hO6DxKkk0BPCcVUiKOvEeF1GMnk88fQxSjGj9Q2oVDMGJGFqIYXiisxWnQyYqPTm5
YmRpT2JxtCLSLlpALyMT7pMSFnVM2dS0iEVkJyk77pJBT9kE0b5/f5Oyke4Cl/E8yqVpGKU1fkdM
SN0BvOqcEjnDSN+jb64dQm5CXpHtTGidESbrlBRRvJWB16z2aohLZ7AQtrPUQ0dWyNdKhWl709eR
PE0mIqRL7xWdM9Pw/F+SDKxqkP6DFQ8oeusUXtScg6anscG6dH4VMQE+dZWrccw2TnGaarBDhZd5
H9scaXYXLXgk16pqaMtCRrToKmPmICRS3dod2Q+4K6IfT426VE2X58p/aX2v/2fPk4H+FqXgXcTG
PvtnEbK6EZccm+3RASbN+ekigzEqGcweU+C4y07vdpNzXcNb7Q5EF0u58HTeDVpV0A6lVJCafQyx
Z73NnNKXZSsTZG+xaw3nb+lP+B+wSr7Np5o2eN6psiWvOWnf7uuGOYnw+8g1NI2iRhr8dQv8JYmk
XyxjNQgK7B+xTARI1/2SyXm+7E70wlH0v4MR8+aQl9X6HfKJaC3G0zf6FYlJdpxs+1L+P9u7IoJQ
0+Aw/lZFjSTeGvBam0CSwMrAy02JBuPf/+dXU1NqsZxqTu5HGojQrRiEZcY6pcWqCZ8foziEDGeG
2YkQvpy9NL8uRqk8zR5/k90LyZ+46mKjGoCNTBLNKY12QcS6Hq2rVu6JRPZHSoGIS1Gzm/4/nj2L
tHtZ1wggXqn5W4CWY/LQo2bskw6VpNcUPJ6dTnQiChL1SAqz7HLqf0TJ28xz9Bs6o7r5P1snDafm
X+Jght1qmees8dySkjDdpI4qwHMIKW5w9tptmQc5FgV3ppo/Bb3FQVzFWVexqgA6QOuthSkpapbV
Yg1c+9oH9/cPpGfZ4c6XamLjAx7ryQx3oU2m2x4bK5aFAiQNXxTKcOQ3ocJGOD5xQoPu8FFmslxD
d+GeS/BGVf1+6kAQ0oh9aBnBlGwr4Pnk3U9rY1P3S76SBjXOkz/Wfnzg098UggNvKtQAvo8swb4Z
jaen1ni+7KZ+DuOZ3pxRgdNCqVepwfstnytNVFV9FzEN0fGo+ugrGlMdciD8uV3ctvwqRp2oQ6go
vOFRZmF/j9It4RmGx3t5+6n/ySSBkybMfJXMwq6irxH5sIWx8oAxpNorZcCZ8UDLfsU1HTtih9G3
sHjt3ao7Y1225s8Oi+VyUhConZPEwHTZCe1C7Ghdo2WMZFp9PuSAh6P2IMNrYwzjZfcx7AVDC5Se
pmikX75Cg7kaukoINWrydhkTYKwmMaePAMaVBoBsPi8J1Q2OP8ZPtK1OmEffQPtZdfGmGdjIoJoX
BQa8wni9vwv6t+ZC2FEA+w1WJetfnRTF15Kan+cQiJ3ZnXvyZmxLzq11TYi+oDuPFGGSSa5MZuHO
yxPvLBZdE6EyYiu2AfY7wF4dkkCQ9kmETzT0kfhLaD35DXPpSBfJScKyX4jvpXQLAnlbYQw9QTvG
4zdA3MYPVc3+35Pk1eRXf6uJFmfsk9xYS9RYs3Oz0nCFVZVVxmlu9+KD0BVPD4lGcNhYx47F2CgD
U5WKZg6KdR88T3wsakY7B6v3ZSvnvJvrTnI+GPyuuKj1goSyDNv0A5j/Z0S5C8fD3JLaPsfCAwmf
MLRTW2+zqxpecJeP1lih7g+IptdpKkKkRQpq5iwYc8w1GGWnqlmdXHiG6bZq4LL8FsRUQP6a35x2
9ZwFzokcAlvQKjDK1bmbiuD3PAmFy2dWdSpm1Pepg8nfAsJ9ZtKOYRYUcLGEb5fVLgZdwZZRGWgk
V4oLFjbPPV5FnbTDzh8/EfU12SfptU+gnzGxW6sJjY3QiuVug1R66iz+MQ6Q0q53lO9Y9bM0OHZh
A2i29qcyZKdFmPdha9DCPz48g59DAVe2mv0hUNYQDGmvq5Ts7qI1vjV29NLMSGuBMCaKNS+er0ZH
1RSpowNVUeTbGUcUBhysLwRf9lFrJtzTFCQ6D6LOc9yiuGWtcITPHMMZBVfbpKwjS2lOCtyoYKJE
iBFdKxiVc+I/q1IR+uEDuTIrTZ+ZWEiNnm2bEjq3Tx68C6XVpLXe04cVUaGYrnwM0yjHmUweP/xQ
eNG51MJ+xHU7k58rjTyDLvCpcdJdIWSkmSzHMcU36D30hSRIYviMduSPADAoe6N11aOgSuSeIbOX
lsFyOx9dy1ujJPFh2mxislZ8+0dM7XlwEi38WOiBFILPkSORxoJxJ/xfCxRsP3FNQadffHzjlEDV
mGbi1KJ3rw6gQhG8GKfr6dsaasv+j8RapYCOcmh82YT+A8+S4T+Vg6INIP/Ezy/vi2b9+HIZyvWv
OVGjpnMLQHrGciuuHFr3DNWBGo6hY6/UBvtzIjsnUV18PULfDsvHjT/GM97p6c9/4T9x1tR0Fd6E
JXS9uLjbZJyLKUqroqHDkKmpEhzpM9sfvgVAOM2fQDM1J1qVdwTwtDtmt5qFfMcuT+l1E++qHmMe
Ozgc8MG78oI4tcrgEZKUsKp6MkXIJnmsxfSfu93O336SxZ33lD+sM5oxDR0Zn6JmB36o46FlX2K3
U70/Wk0RvC3ttm+F2ni4Qnqt+9MrftnVd8K1YwwlD4QKbjcjCy30Nzzoz09U2zvBgVsey2x5CZoB
PGUAjal2Zi71VeYVoq8Lp0n1V91o39QCXc1aY3UxQzn4xADoPKd99oKISJmAN6+3PUB1XOVZBQfa
xgsVkCn6BZWrJDxVaFuQqf26mxA/qhy5gSlMNy+ghSHWkqjD3sB+4AwibRDfSQ3H6LofV1UO7XJX
R6QExszTP5Duy2/NY3EnnI2zqpBIh1oKoMSJGxeMhFKWthT3judw7m2bRc8WDcDoMH1GvM4wswlc
WgIS2kssZEKMSlVHqNs1oh4xBzOCGco4CFi+2Cfuz0NoNXVyxDtyg7KLm54iI5XOgE1ODSkQl2OL
Jb1hOQcKzmZ85as76o30MpmffBCMHS1gT5V9GkyIoHyQDVm78wYvRWnop1bIaRFyJ+jE5Wnx3POx
yNIc24KR+mt6WoCnyaPT9AulTY5NhtkpUd6ITe6QzanVd4YDhGbX42mwZZF08yMfvR5JyH9f0jn+
oqazTES86YOn+j4U7+v1s11I1pVolBogAh1gWtseYS1sVEN1qxYQSTugelb4VCDUIywUjX14rMnH
jTHDVF2vEsArby4SHQVXaFiOXOn8FBm6NkZMoNNahTb8mHOTZIERz55babBfV3X3xq7RdklEIc1b
aqhUkv3Kudy3pof05rdDWPlm49E28ycwN6Fxtkqdmad/xpZnpRzHNGpVWpAaFH+J2XFFLNOl0tjM
kFYVlOfRmXMwh0nW5ajZPc5cM3nr4LZWLkdOATQ3Q981cb2kCcE6u89FUbCzakz2P42RdYpD+jkg
oJSKn5Tlrgb2amhspkc3QKHaqXEhTHJTlHzlkXMQ6svemo0D9/fOByAsUFdjzS8fB1qVRjDPUXir
4IpmLOdMaST1w/EG8qex7pGgDCZazarLS+YCeJYd/iy5Qp2+EiwgbfDqT9bWzHYZPuiasFaoEUjM
KcRJ/UuJN3dlz94dimV7hu0gKigCh4rT6Qdboxmwhpq1WMah2gpjLvV/LZMQCtucvW4ZePOETcFZ
Vv6VRvIp3KNil6DNnOOGixRb/whllWVCVEJn9++DnLYzj/D7zmUMpoin6TyRyvUsvzsgFM2jRBYb
PxG5MUr7HXe0OADm0jfCgV26xJ1xyVFyxVgnhbs6QLnTnxqKTSy4oIKeXxyyGO5DcL4KR/iKCwNZ
l3uON35C0PETmjCGfA+eiRu7+gDXCYiZJS8BCH7LEFEei2vwByqs/8pwyNXEtIWc6IyhW4rb+aWG
SSA+y4N0jQyK1cP8R6RfDDnClQ3pD4dVRZHYVPY8N83rJZrykp4dMjQ6p8KqNTayM4v5TyMOKfEu
Lb+TdBj4oSy9/XO0vPaeYGOxhJhCSAp6OwfD5sMs4BGk3FieOJlh6gE340c6dZWe4lUG7QRJcP77
1zOWeYXKaEgrrNXuTdRCfgMF6z+RoH6fIbzElROyMdSbCVefgtBPe7Ry8qmDPJSpXNCwEdsjEioj
lIjcYXFQ2TcBY746CvJA+6/uPhxNVRR723VzgwywTDkSNx+tw4MkbxM0PGvx+FrkW3wKh45z9p7R
YBP4P90N2YEwagOD3g6745A1pRE7XWW02kHNDCgkKkodcYTqj0sYt3A7N98AU+KzYn8jftQU2C7U
sZ9H3ep/tKr0LbVnyDfS5lIDvZeUkj7kL0jJWfb/9gIF84y9mpfDJpJd7hwTEOVW8m7a3puWxHlG
c10JPbmGKtcA8TAfbhBEOAFNZ1FcGdLgzc4V1bUATdtZr0p3ZF8kZ15ExKxyq0JccY2NdNEBcf2T
yuAU2Ps15udQ/0xTm2UhHKPro0DC0pZFvYWtrojjl8jGS2HjjceQLb5JvkyOtTPwWg7MOOBpGnKc
RMYxBC16RhWSGyhiVSjFZrUGw9kRzc+wnMhAg1U9mr5sIVEhjg0ium3jfk+6q3/QcGTfIG5WlAZ+
IlYB36Ugj3nizadaCFUVh45FQCDbSThcYSdEKuX1MWxv/Kr+C/EStFYuXmYNb2c6SSACazyi25pF
GMkTB+bCTlFlTcTPCsRV28rb23Zd+PYCJw+7DBh3aa4bUyEXz/qO7Tjuo2HwdCVGFMfMAW3H9+ut
b6mY+dpacd9JeY0reCjfuoHQrmQL+T+GsX2o+XMEXQZleNj4ajrQBRyEKydaeBXKNBfMKygahbwR
dNXM2htU+2aWv/kPZwzHeTDipE04C9cFWX1uLku8AJNAvBx+HiNKXfH+s4qGhdjiNvHj4R4PrOPq
JhErBim16A82Kbe575GsBq8wHOiS07z4f7DvYExVkDG0aerocnJGzMfZLseI70tz9XHYbVOMkdPV
C/jWxCPKGqd3lX9g3ahZ/n0fMsatgdMFwjvt8dttmWWVtghc5zTv9g9Y2zVU6yBL1U8na9Ij+gJp
2uMgd+QUKiL2c/mufXVdTkhv8efbizyNTKtodkJ/QR+kKJj4nOcpNWk6nMlFFNiR0T6oZMSmWMTj
0BEXsfu/tA7Ld7GxlTg605viC4h/2y6IGIfvZt2fphlbQdtp47pHj9hhuP443E1GBq+V3FZA4OKU
0gU1bqkxvtHGl+jfRp6XriC+/Ispb6qJJz6BiadXtO9pc+IZU5uhQr7W8iMJnR5J/+Ik/8e/yM6q
1DFwt1zI2vCWaXAPlwDt4P2fE4RV2UVkrApcMWDOq4PGfqXRkLO4p3Onk2+RaU9Y4Dt/ABTl134g
gS2NqzoIB0BtBoO+ajnCPtuAeOxwuKtfDyK66EKtdGDiCwYX6EEv5DHmK4WgjGqOVWfY7guNNY3I
XqpyUPBBVvfSuinhKt6+OfSKDFPhfG/D6Q/7bWXa+cu0preQTyPgtK0XShNQ8RQl24xfadzvEsI4
aCOSS81fU2gZUAtjrJ5+nBe8u9s7quV5ujm+XP5PDfj2KscFYjgzhpIgS8+CLyIkyfTul98R2srL
GERllPWS65PTlp+AUpeh8QBbSZ9kP/Ve61GdvE10/GWtwmwGuykZvfkOfriEqEnx/6TcoLK+AC9c
jVY0C5XP4n1NTlXujZprkIM409Ef4mFG4VusoNgSb34nDJeY46pAqBJ9hHcgANy7ILLh7WHUTKCW
FN90Qk3j7niHwU8vPfnqH+eR0vLb1scKRaAcnzdJipTv11Ayx8BpatDamBgv7eKlXFAXdPskgyMR
0RZIdxVfmiwEo3kgQiuesTUlNP5g0gn3GFk/oXzb+2+RZlFXbPwCeu5iyYmHaCMAeF90U+qd9Nd9
dPQLEcjaETVsAjzcHAPZYobKUcSEjDClWWjQbKL1N8Ge185Yo7n6j38ShOwUpE9wvW9J9YYNgcqi
6NytO1klXTz80teRqOk2BhFjY+aBLRu4fnnd9lxXYYlRf4yXU/7NqHFVafrBqAPbVCSb4eQvJ+xB
Fr6xYLCKOA5DJfi3iidRU4vI4/ZjM9bCTOioaOMr0YDBacy2hdv0wALUQpIr5hhyGaBZPDbPhbwu
K3AZEMxaJ7yNKVOCdLfvmjhGp08LyRHtHyjmz2IdF7IQ8E9cxR4lqGz+f07V9YLts4zXWzjxO627
4DSCum2fFdssMNJ3AAgnI2qF/i7+SDdkhco3oOSUJ/9ZyJp1oCPzyWszCTJZP0I+4/o2N/JP+8GX
DxcjRp4K1MYK8f+o04da/VXEj3nUrAG7yrbidAdBMYwUwW1M38RY3WwsXJ5ojkVYHvM9JS4SMC0C
EVQBRyvFxlPUFCzZCnT19t5Xbd1f9HUH/siJiFHvuG+DsY/PIg8iZ8tmoirqZnS3yZVTFgEADfuQ
zmLuxbra19e0Myqz1nGkZFW4ynto55Fx7d9vDftUOBEmDlPrvKC1nmYRmQo4F5yrN+o0EkLz2ndv
cg1M1fV+NadPpDddetbbZVCfYp3nrpbncKU3FllTTT0CVLOFOofqPXPZVjNxzyTXzm/KCmAZkBdz
VnyEVwXr+1GwL9We/6CD6TMjnwipIXaSNNwBU9OnjDW700iMa/PBp8XME+iRiYZloiFkwOgLsFtc
78Jb8ipPSw5ZK3XjsPbxrKxJ2H7MrhKDkbFmqXzKHB0CcsoXvkvpLBlFB32KUD6rgbc2LKXCM1cH
avOPdwh5ammpfdeoAw11Ep/h6qitQsngTLfN7S640SrKUctG/wntnS2DMmRY5XT4IepOU0jwTRYv
f7J5C4oIxn6p+iJxLaNR9tiA00NJDds25hem95QSUKLcm2IhK+zHaa7MQDvGCCsF/WELT6eoq1q1
4FZPZQkQN+yhLE72PXCtDxbMit43WwRYxjIBckjVbZsOiZKCsgL8lcmXz/NbcMDbQFW3p++InHB8
EuXVtMhBSanAX6NLuLlnIFnAOa5I+Hg7VJ1E+JpOtLGBH1HUtRADH9hBIMz8Nh0VYYQNwO6+7z+e
439BI8/sRYMnObEHPmoGoPmm1GMnPTomtnr9biwlUGC69ThaFZCGH+klhsWRR97agCCqCAe3awjG
fLuB8MIrv2mOSvD+OGBYw3Ju+oomeQUmM8EiyqgIcWKEBXxIyjSnKaeQC64Ib+tMOxm8ypn04Yun
8i+CP2B3HVb0ULf6NZFNPy0T37G/MHLWDgDsi/mSlY4mIxTyeSTX2K3hafj8TqpTDteiZrDlftaA
4xpUCwc2xYnA7R2vpF1Ey+oiPY8RJnyfebTta2AE8DDV0HPLu1DY2H/3H5qBPI8Zs6a1ryYP5Nh4
m2hSZwv1pBbS+Bnu/l5O27CDELw9uMpq5OU8y15D50C8iSW7cohsdfvJzi2WzuTxnjOwyo1Cpj+D
LHdWLdTePBeBON8XGM/lnYK+IKB/ERtGqPOz04JbMQuLsaYK32iaG5ttizZZYDilDO3NdfQKH4/8
eq+z5h4qVfPZVt6IVjklxD/uBPtcedU/10FQ9rF11mFAt2oMep5EFk68Fn7SsQcGt+1huO7DFB/+
QKKht2jZB+CIZDaAeMIFa9cBOsiWq0po3pu9y36wgdZGknPCCIxglYrKI06kaSHQHDIGqjD1r1IX
ir5WuVKhK/rGnPNI93nTcxrHjANkd2zbJEIwmr2+XyT5bnuIc0fdfuZCigyfWuL3Zs8uBRwpfTAh
O0Mstas2I5W06IZl3FkgpoNFejUTRHnuP0pzaJ1M6wcix8qhoy3zXlO/7VWTYBenC24CkqCqCx6F
6Ba66xnG/IOQpq2ZwmgJrMgyXWUxxBukmOxdaXx5lqxOUzaT9zi4O4JHr1ymgm5fhZ6JCzzTwTPu
58M2aEEj4hCb5MEAUpsNdP9GeumNvrBxjrMP5GhZaAIoT/6Ue1PkUQi/y9ZAx0Isund1eOOLASPi
xL6CUUXF1dvRZO1rLsPFrxFxEJqodRlQueevlYxwv64o8Dt57bW69kfkC5Jd1YTu27Njw0Zg7VE+
jfCoN9819WnlJJR+zkxj0qI1LUBIyIE8YiD/tu/Nonq974LSzRznYnNp4PkOQ3vU7E8PXOJMBQtW
Yrt57gPYKN5ET5HkzM3+C+v+Pb60RsmmR3NQvR4w/zBPtKEg/2XPBumSqCtZ0ie5ejYfnpsiJz3Y
G2jZnTriBUamJYUm3kkRwsLM5+F5aMVpGUQ5daCuVWltrIX2N4iAFaD4sBJ9SuU0i/BdURh9Duya
pLo93kWq4fkj1gjdgeXIoqzdLZwP/ezq9yH5sON89eHw5Lu7jZzFjU6ev4l1tsjDOuD+ppIoe58e
8DmfjISjsF7xVnceCy4zsM/yx2ML+/rvflXFHMDjcZXbnocwFwmvj7uF0at2W/EyYy+ueCrvqfle
3/oRsWKxLXgaQzF78RphKChskKHPzDTqMIsHcQ3VMCho0r7tR4PETESxgElGyGuTUvNSrS2j6eDS
n4ffp7F9EJp9Fs3Mfrj9zJ8nlF7Xnc7H7p8NS9wkMzCI5P4ZLn7OWoVm6hmCtDsXc2hxLQQYbXDr
ZVZLYXsDUKw7IDCp3owvqQu0QPebUWjcxIip+Whz1LWJtgWtmn4Cb73uQ5RfaKczdrHACZnnPk7e
kohmNLL1fYqCEbQxHkOzTIUuArTdNQgwMYlMx6276S7wiIinvYMPIHqGP2qMAUpryJ9M9L8qlwS8
NxL+CK4EtkZ4xu9/3FtweiPbIny3XjOVtu5/4OKmmodijMVbO0PzPO24c1vEG017JXDo7Ir39QBi
cgngjllv0ZXOVGtvTx2ZyxcyxTEWkhtf/ZBdqMrjuwd1UpJhdDiap11pCUy7j+1w2bAXnvv1PXwf
l9gjKhghPd7Pzf+iAsb6dqYVcW+uAGEOFxw/FYfzNkvKG7EQaRxMEKpL2lSaXbhoQOH+QQkJL133
wUeLa42xCBD5p6D2ULUq/lSj0sp3ecTbOSH6LSwTxwT552BJhC/g6EazPiCPhkRoVwe7B+4foBp/
fhUMc60ZUnXdXUo9Dbcoi+3vII49En2CYW2XSfVqzcH952KsB+YGNziDXONpLZEBp2cSFK+DEWaA
o7vMu6zvnQBENzGnpODBOIBmrGhxAK9LDyudfiNoixCLGTE0hg/6u+MFVAz/WSPW1VHy9ranJ20B
E/Y3APunosgN9DAOhE4dJ3NmTcStEmBq7PDOTZRO8GMgI9iyk3GI9OaUkVgWXr5UrtJKwD5h6Qrb
e7MfrDiKVtgg9gWWjHlCj8hjx54KZx1cBd2aIduTIDJxRghOZ59voxFvwHOt2dyFqaq8RXrfOUc4
6tYc7kpGyMwYBstdXHe/JEmSmmtureZOeY3FlpLQlWH0MCHBCGoeBExftn1+fOWykBjPx0AMGVV6
7kuErbfhNi4okgtsVy1nOE+F8Yq+VtGiFeyw2nhBNPyNC9kzoQx5ViW5qMDEh8mEPHMz1HQeNNf1
nmFmSSAx/vzQtvKSKw7gmnsipXtSRXuwSME30H2FO6UjAxWZjjSs1FJ3TotAI+eL/iTbBo80iolk
E+NjnGKqW8JoLV30PTGWAUI5i2cJsBjbF1Emgm/jC2vSPNgO8UMx3Rr9mBb5hc8sRaYliVQhMmR7
6RWamRiUwuTsQLpmHWnT8/1yepPzgCUUwOU7qoJpU6ut7Wq0kLnlKWxVy/DZ+qXJzz8e9k4sDTYX
5KTYfdjX2GqyyUguG6RZL3d6qjbO+PEP6I1d35fi+90OU84fuXI3h6xWnlvwiyTcrOl5wrKkqHOq
mug+UolvPAoIOcbVI7v1iGEhAtQWtx9B5G90CPFglGNewMHgY6vCTgEo3lJcbFtVSj433VAPjQAV
qa0W83d6Tcd9r//s54bHcVdm4z40ic44GXDzcf1nyewlgfHXvj6CdJWQufp30AZoxEqAmtg6KdrH
/n3ipATKP2DwikQaStNyBCm2lk9Wa8GtOClti5re+YDqkVD1ibjbOgJy6vZHspOOTa0n9JWezmxy
hSaWYb5F2yQgPE33BNk6B1p/U8yjOqQ6YjSbXUfEFIDvCHQo4fp8ZdKAk3gHBdXUThWvJNFbepCC
NbweHfIMfNODDaaPJD8r3vmjqB+xNdU5Is3LWG7DcE3UC4l2D5sKkyWnMlC8hNDQf+35zNCiSPRG
0mwVjII2mZf98euC7F80GVm7DMQOE50vWKshN5MOz94BzZhncGinjTs+IK2vbRCi6NZ/t/aLTbqj
iR/ljYFLIpV66f749jvrXFZw5Xq0Gi1zbjo0G7JmPwcgqbr3EMHHklvcuwBy9qbDYidNKSW/qhZx
uf+8SkdpyVwKlqPWCPTH8HaBODE5ieeLNeZ71ktUoN9mDKPgzp/leodhjilN+/kTQOs4x8y3/OtG
p7LdSsUxtj/JbBo+mX276XyDnSkqa6OavA3W1mwpfmz4XlZYX+KFDzlsU5U4uexr1zKWRwPd6qP1
MxUuEXahPLDuIcnaE6d73uuBc/ewgpQbe5Ah1PrQZGK6P8FMeCQT+4iJ+kOo0GRCkv3nDNtqaRrQ
dfR+ubb9VPcAlfRTCeY48+eVjmiJOif68ktVZOlVBmeZVtiDpMav42SlSY/eJ/mv3UnEpMY94JNq
gaio68KirW55Cufb3j8vJA5LaAzXYxN+FIJCTpSwqlsK4M85xEb3XLPEyGEoRrIyQXrGHbC61R4H
LcWsklyvUUU1yEmgRCqVytH+SbleZCPk6E/rslABz3iu9T/RR4u16P9W8Px+rd6i3sbCDLrAJ8NR
avGmPKobcDgnIqlKMIU3KeQxyJecbIOEKc8JcQlIwNKjWrM/PusmjjGfiGHPBGaWlE4VOfoh7x3C
3oj7uRsiJJ9eab2SgryissbXGZI+NSfn7CvwnfTymREa6vijvJi1+TDdWYwQXepWnxfTtfEUgj3G
Kjgou0sql4GBUgp6+JvFA6+FUCn5LjfWgXT8kjMlJWCemjO5Ahmwo4XrwfeL/oTuBlnkcANbFBkw
fTtcl3ITft5yp3e8CErId9c6tPS2Ws+xiNEDtLzYT/G7LxFM9wOlU3st4IM00kj2uhOmBNut4HoV
jIgrqfZT/tzM+3WJ98ZpIi+KTPs8hbKSqtow/rQ1cRyLWA7lnoORWA6m5u+JSFNEgfk5uNzelhRH
QKeyYX9vrFzCHeyYRuJEgN78fduEO+L7A31fPS2yJ4SYgmzUQol+jCTqVn78iqg4J8lWi4bWlZ2d
uD3Cg0ipLGAnLfY+l5KcuF4ARTLXYygjeUVEdv/rPUtYJxcIw+rqsKdAQR4FfYpfMAheRLMPZFz9
s+oDKIXLcQwJ/vk2cPBOnpz1p0Gp6f/Oi7wQMOCODsbJKGouex3XCX2KqSrG+I6805qIp0mVrUE+
IrKuqBETbuld+a0iHDXm+RCsHPx+oKuyHPB4SFAD9Nfa6X+GSkp0ey6amZ/Tw87+fKehN/33Qjxl
9uweio8Q3MPvZrgmrk9nBieXTcKLsdbZQi0++zjd6GCooUwMxBJt4CnSMYYwTKbXyTXTALXcDNsl
0vBXjnRXws/Npd+JYEzS1s4DXccYx0Jovq4a8XdsvPsipLBfq2rmGvkfZJq3T/e2TmSkLmKGrRUX
jkph4wpZxdeUtsDKbH6ZQXiBnf/6/6+A8xQFV4nOFXB+el529kQBLZHgRVeOwHLO7BcfYsdSje3s
fdNYv71dliw8iCybrlCMhj0OaYQw2bZNLFQirrbuhbYKFv1t3shBM2475rblPC4R6BPRzW2LXV/c
0TZD8L8Pm7KHvTYJp8iW5KGUM2bKZtjPSivtgvLqrLt30d8hUM7pmuIAJ3zB1fhOgP5uQv5/OF/p
0TiQH32HlZ9os7FRoq4NOSeXBgX3MVK1QiBEFoXiS31//6LGeepo6Zw8MgiCn8jAfNmPo7AXaVjm
wxtI8oPH9owHC8d4s4gq3TeDUTRtvMOy0cBeRvDqUCsjMucY1Jz804KuQFrmWDxAha2KRGblkDPX
tzidxk+RqXkr7sZEoXmxlvlAMuMe4LEPIxtAHI0nyb/UurHpncWVq0HVxkKhAK54IvoNejluDvMp
q7fd60YGOsE/IzhcsJhaxHu1xvPavuVkG1SKdATtcVOX2a33p+rSlVR5TeWDGdf2MgC1hvqj269i
AWYtmjpGRLb99p3KqnqL9qXZpmgT4W6dchgI6Q+Kw0SgGPGfIRsSf1+nTcV2mruqHZVeTFX1abHN
ul09czO3G4JkGe9jFNBEnC+UKS0+8iNScom5/zICe6YC2Wo8Wao3dFwHA+UB/gu3Z+39rt+2mDni
av5/9RLhD21nq22l1sPz7gXRoYbpJxInCt2Gs0bai5u24YGoZn2bw6iUOsrGJ03yQa3HYrJjGm77
fCWeZW2vbmzBd7TXtLT+IT9jGR84KY24IZDWW0QAMnN+NRL1OPwuGf0ThOqFBfTn5enGvqepG1FH
4m2lKX88s2c6LS6mWuNW4mV5x+0Hw7+iXW6Sys0jDIpqjRm2R5Yveol70Iy1HVFnRGvMEPtlNO68
gFl605OyF0ugbcAVMk3UH8dbLpij96l4SMGjEIe3DlTXGlr+I+1WaaDo43oihroTK2aLjgonc9H4
+QsMgJHu2cWM6mL3oRPCg5jezwpua8LF9TVf92wsGxMQXfkfJ0BIsqz1BGdhY1PZ8TWEnBsyd1OO
GkSI+HIjd+hywijG0sUfAPZiI/sMnBsP+2CzP0pnN+uZXZExoLGKjH29PvUKdlHDWZoLBEQHslvn
rkL5bsw/UsTuFPyjP17UcZ6rDFk30b39B4Z0peXgUgBgHXBMt1LmLjXOxFtUb61tIyk8uFPuuYrb
9+BgrCyn0e90Drz4tKMI76V4JdYstVs+L7QbYZjXmKxGmX9jpruCvxm17APDfbj9wK+/5FDSQm69
ADpLKNx+VIXIg2b0HmYYEXZZUhPQvs5lp9WUFOF8eJRp/ZTY5ahBXQtFN/rr3BjTHSMXH2zovseJ
xkLy8fATpfsgtMVj1bPoB83RDbj2MC2to3oYMZ21SGohIRwTpxZ7tjYqgugFDolWZRBr4znA4Pod
vJj4XIb1tiA7BvYwdDG4InkBpiUwvDBtPXtnw7UV52RqLTEJ57q1T+/euhfV8VpbmaM0QhHs4t5z
OdR8thzKMC0lMlEPDrYVs3GiGMno5i4zLKlCa6bUHrL+Ch7pIk/gIaj7VzHXtdukRp8ya8u6m5wt
1V8LI3OydDVSu+hR64ihREn1yl+efMq3h3BSceOGdOQmdQNEyompZKgKEAiso0BURiVeaiVLxhS3
BOj2bUhEKchWmtjRk0JkydyyIk+uHUDUJ63jevBIQD3amLRJjxhVEkQYP2w5LgQ9mmyRIaD6U7l4
c0q/zxmfJ6XeQRFSbLpmn3AM422iE1u+JFHL6S8eSDKUvfdj37X/V0Qb8A8rL3D+XlT4l3wQCbEu
YhiKzqEZYNPAJSV2HwpWsQuSV6HWSBJHbYHO10jus/i3adbmq6tky2T2Wt6n/jlBm3C29vjCjiAT
NizOkQRka+H+hBNhYrVf9aJojSpK/nkfvU6XovA50EJb141Ol7A3VTV9PhmQtSSurbRkRITfMmJ+
/U9BxsjfpryO+P6ZHipS3DtYOS58b8amrctJ8qEj6fIcUda4AURefMRLnG2V75zSPUGdIs3wYglP
ZNwe89GQsTkD3vOOS/RTw1lVPPLbCdiL6OSEiD4MWkWaO1Wo6aWoVHz6E2ZHdq5YUiXOFVo2wY5o
PAAd9CTSEQXCZl7ZuWK/n+RrQ0V3uoMBt4miZCovOi6brjXtW8nSxwQIJRvBlteMkcHHhUl9dJq+
QkU1uAEzCsLBye8wPZm1LoibZ7OYOCoI4QjHP3grkA21LCDwTNy4GhOb668ep5g+P7RWLpFPYzx5
Lnwor4SMborUIFUsiUBNgMD4loip147vDIcDjolZT005A7dB05g9m2a7qhefDkoRx35oqFbZdEGG
NwTjtk3MQ4YdcevjWaRt6tOJhD2wNBHh+aXjpgRlvKAnyDGDQaMPz4s7e9BJg/5tTB4b/bNtQkAn
t7sm2UK3rLAVZesmNEGegv9/v+hjatp8vVM9p7v7wJe6HyqmIHWXHKb5m2BJ981u7mW6LC5tGLZD
XEtQ2Wc+1nd1ZIchs/h33JXF6qXua7V1ILQycemBbawzlbllMb0d/lXO+XIjCuIVrXBV/ppYYthU
pRUJ8l+CxdddEITBy94+BvRG9S9InTu29huVy08+XJzRrkKlwumhWfnb/qybWv9UgoQaI2Cxoeqk
1S3QYQ/EWUWsLYr1YDHfzxmanvSuYXpThWWewkG9c3x8wwe6Wb4i9E3C0ypHOs+8t0ufi3vPiBrF
/PoZezPlGmWwkuljmdKyCfUmBQAxOVKsBh4r41Y+k4uXJh5WCT/QdMP4Rm6BiKkeubATKjWl7p0N
ST/Js2HslMEU9uVkpFdN3ZRl8ZGuAPw+bWvKRKn2ZlrqKZ76UUc6ZkYJyLoPNpUMQpWE9MmU7X+n
sEJ2mkrzvP4Thw0x31xCx4kx2YRtTTM1qMSQ6GAygPWmy9ls0j0W4P/cc23QkG63xGBLgzLaptVL
cBV0D4oc8+Nn3C6/dvTMCNiWF9814t6SyDeLJ4I2JSRXe9L7rU8ixwMgQGiHBsBMKzhZVfoSZ4GB
v56aB7a86MTaJMNsv61Zu3/9QzvRuV/mJCM5bRODkX55eSPXbicr6YwMwPq9zxWdGUshjDQr+7o0
ynz6vh4C9JZ4m6Lux+PcOUrUNmEf6oPPQkukWs9wgYzWFOx0VT7i/4HMH+jDTmXHEYT9AqxGoQNQ
vXeqzU0yOKBmkKIWHZED7bc6Ac6C/Geta/Bt84YnYZipbvSSegu/Dg0eYzzVgy874BzNVq4TitVC
3YjF8iPEoLjitwuYBomkgotA6dIJtSC6FNtwxXp36DCvV1ka0K8FwfiLHM8uQE95vF+3TuULgh6Q
VVc/jPZH3Skj5A5odpMUfH/qXhOGKPu4J9ldvF2QoVoB4LCkp5y6OnpjDBMon9a4qbgFOL8/Ezb7
Qlz0+uH540kvbzy10N21nxLJQ58JjLl/mwO0oSlLBFCwIk7hVEHX8stggxRGBBKSIqZm5/XayDhi
987klYF2EVWeq1xp1goSN94n865PpFabxFsRBJWMn60R7kAETgFeFnqEzgE87GPCkG1oeIR6PLBp
uWOaDWo5NzH8EdFW4wQapySD1cjogh9M8WGrONkb659jKL9PJQTVX39/EYHG5fWyB5RWapNlkXSu
nemP9doqw0ozyG08JTBoWLo0qYyamN29iwsr/iY7xoOu8J5OicyVT8Nn2qAjIrRHuVDYUqlYmZZF
pbrNmDQMpraaPJ8Yb5SQ+RwWBcy1Jel1hdAywhsLk425XecNWsAWhpo4t40+TwhFsbJbh1Wp2zaB
hE+U9cPHhJ2WUa7JTTGHZTDpHhqkiUjIV3KrAHq40osufixZ/rOT6vZfd62OOlika6awh3cjsCvn
4d4ycNNkyDQUK03CN6ry9laN5iXwyYQZNTIAsKD2avOhUumdM0zWKotd9I04qLntzw7YdQnNZb3p
HIWIbYhygX5UIr5VYm/ejKqC1f7BSYngSwfnfNVdDtyZqC6y1Zf0/hw9fSZQMOExC+wFZJg1C29g
ibsMOjklEaF4YROdg9tMK3rEuTB8JF16dKazDMtG7btEd9cNQm1XGMGwLwMyRQsxuNEUaM7pmM5+
K1HplGnXCf3rgLe/E/jLbhGckfx/BtS4bgbu2vq4Ozd2VHJy0vcibu1UeMC6vjrh1uXWwdcJv4uM
9q2p6c7HuLgqCYoxK7wNRiDH+dKrNEhTmRbJomRB8M2bNXEPCSHzd0K+/fMndzxExoiT/83HRNVI
TT8r7Bf57aNeWB6AoheJ9NpRFHsyY3oeQ5tXAE2lYRZPFWAtUuzsZGLs42jRU3JRqbgB8zAx1Qo2
Siucp6UKSfow05e1wsng5BOO97LP0IB6xxcNQYYNXgP0zJGyTuGkSJ0plTBQfcbJ4GxVKkQzoDSC
AurvRBKJ0GSqQ5063uCrVQCf0FQGVoBOtyUJUgyDwH+S90+xLJS92/qJfX7L1lVPRoV6CX/TV/wM
RDaAWbUPn/FAZhGgj+okshUuhr4O1HVNR9sM3bdz8D25wzhn3M6ubGkaZZJxchgQk2sssNc1crrB
AtIzMkIQR4tTE4TjdbWAOiWZ9OO3fmjH8E4oqcKk+4+4Zg18pMMMbZDyDcKPaXefBYSIYU5mjqtC
SeFUT3KookgdJ8RCvSqsRHsu4ZQdbefYVNg6BaI8Yn7RxPkiVlXNurH7jh04nP92Pmo6fx2vTQ7K
gKA2yVXOgrEYvZIVZJLsJXw+KlJ7zL82bbnM8KJCSSqlADhZ6zKhFKEeiMDeTxOxp6Hmy6hgfjDf
/yNwrailF+Ar9DVmgwqzyJjNyQCfJzUhN5JQ1wyE9CwKw5g0WMyQCXQKmsCLdnpf4i7piMmwRhmx
XTo3SgxNeHqX5YgfSjGTgyRmEiBwK+dx9yTy23xITB4NPy5w5Y28i1EOBPwbxqIu+z4Xwxe2lk6/
1MAdbS+CcuBN9QnX6FJjfeLFAB377O37X2pOzRZVkoKy2y8m+X3I7Zmd7q+EEORXXY/as3P5/5oq
9zAFJCGnqXD5rKR2AVQZN338ASqa+q1wfIq+d7XO1PHVgKYWFTXZUFXwd8u0Rxq02sF47OeOJ8u5
WkUcUPjJOZeKd8ng+8/rVayxmMA/wXK4qHs7U4E7ycfQ8aPViYojHR36f1PnBtZuieiLkavIGvjK
evCWmMbA8MvCp0QjtnCbAt2grPtbi0utI89vN08fqb9cPHhqs+gmYXkGS+BSyaMP6lAIr2M3Dyg4
VuAzozBTzebnudEku+cQUfHJQsdHjmEbeq+L0IXt+oj5fjfE/QyBaNeOR24G7fanC2lOcTQFY1LN
s70jsZuvMj/driGmi3yIFJDhLJ7kG7W7BSG4vqUS4U7cPu5v6Scdf0/O8o269WIESxd71KvQvrQc
5vAZvg2fAEyK0N/FlLhFmNnKVebDrABYxepM+AIGjVaooi7pEvS056UxvLYdcAajaAKm3UH/pPaP
4IOwJxtEj9/kqWGngrwGRu3r7Xo6/r4SXC4YOFG8M1H3mCXeUX3zqoXnwIiV7E0tYQ6vz1Rl2232
m/kX6Oj02Uy0D/+RR4xBPvhnsU+vzH0dUZDLKwXyIQ5YDf57stggBLo4XuTfFB7StlUTz2KF+7/h
zp8oKfB1d7TJ8Q157v8ZmrfTagngGMgY3m0+s8ndLHEBM7A5Oq2D61JPZqo0c2WvxO2WzFfS7E5a
3avLl6WcGzPsju/Orm79vACZ72ExisYg83cumYgolrjc/wNbNNrA8u0aXQNHi149ak/7dFDxWg42
UnqCU3uo9cI1KmifpeolPkz+SBvskIw2thHY3D7LEyBcV3+2uD1KGofqfOxG/IwH/dzKnBxQLJ2b
/eLCwbUhFUZKqUa72FpHueKbl3/1OPaIaqc/m+rf65QZK7yNfGGBjXLWBISK24Ir5fnPIj0ER13C
pv/4esJmlAAib0Fg+qYUFn+X9VXXBs7NPeGrKUlVdXLD/LRPNU1ZyoNKta0M1k9DByJJNVdZwAJ1
HZ7/8DgmQ9oWy2w5/apbvnPIVEKgFwZNAZkMan5w2na1J5+4lpPCwTNb8fQBEhBYWNSVdSjJMFix
Eb80v5Xsg/0bhwtrxFEo1+/1N4EIbH1leRLV5A9cX3qRgzwsVIet357rn+mezrogmHDsGARkbXdO
maSpxe5Wc4GuNfqoYHwk/Ph25y0JlQUb99AWzDnVrTmsFwPdsVN8TGrD/1UA/fbOCef6pE3j4sTR
Fy1YmCd1ep92QO8NBLB0K7kHglPzJfv5MpkGgoU8SnVZ70e5B/YMie4cnhDcgFxbxG2/rPEp3KCH
+wlKYFyw+DrWwXlDOOQqTQKe06Iv22+53hghFXrcuGCtZSxALXkDTEsrx1iqrRk5ceLWix71FTKI
LDN0yrBVWg9BocUQS/E/suh+/HQS9f3yVd+59hcfJBVKUPFAlHjhufbZjawueWailuOPNi34jk/O
heVkD6JqqurxOvKXhpL2RWMXtmppuCM/bxQBKl/RjwmCBrWGK7KEmoHyKNxEL9+Jd/pevEn0TXBT
ZA0s3uaa0foGb9UrRQSWVWGH19ELuxJSQ6oL3cG9ChdJxIUvWZP3+2zWEZhQRmJIXXBNDaVuhgyW
HhInPJYLdZY/0wW34n7+7fdyu+M8k145HN7pdv5Z6TX16dvGXK2SxPpp8CIeDh82wvR2t0Oycro7
vOUrryZTs6dlXBjq0nhM1B2hBNyHwNuyQAkBt78cFwf81FXokIQV5wQak0C32o6GFwPMVQz781QP
vp1XyLyTrWc07PwRGKP28Hu/xlby8mCKyfUYrDyM3lodcuOF+nfDCIXy2ZWeBljYlls+GvVVEphr
9Vzh4kvfpDMXpaoOggktnDXWpNn3XKWTVMzhkj47Qp6fbAKCZ+xKpmOkQ9nDE1JbpYPLjFhtyStS
8uF4xTnVOy63abOaJMipjUUfvXH1GJ8x61jc6X1WOS/Oe0a1DoIFcDIdXMnZG8Ty2sub9rVjrE2H
kyyd3EpoQZ1gZ1329hQh2JWOYUrOSZJGuybHEdB9/wn9wlS/L8/jQQknmENBVgeMLhFQvwdqvl5J
0hh/V+lXPpcOuhqw76Cwnv7xQRxsrlks5gOhcLJMegyj491OEqoVohG+dOZcDs9kS+6+T7CBI4gR
n+dV1HomOJLoZBzh+/BckKO4aZ9WT+yne5HLCdIgQzt56t6iNhc7kaMyl+9wuwsU6xNoj5zcv+li
uuk1z071N7IK6YyS9VO+ORIkOTCdsOtCXjp5qlOD2kYK1+l5ChKyEj8pW+QOhCdPDA4V4vydRYbs
/t02F/1Kb634PXIQJw9JjzkKGMuxmynZ7iMjfweA18TGdkkpWDdu2mtku7h3OtJHVmjgl1HhDIMU
kikyy0Ewu5SYFPgDSSD5WFkMefITCEsAGdWajCjIROFqTuUdkmSbbUVFWAPUgnopWRe9D7NFiqzT
TCo0Q126ncrDS0JydNvo1Bfaa6mdHDVMNawnl1UyJsGNOWgBU5gNJnwoJjjaeY4SXeufvtLlS06w
87WvA6za/cDjRu4xh5HaTMYY6Wp2ZvJkGlIp1VrZrHrcS362yPQZU07tylPNNvsnetJxdAy7J6y+
zd6difLYAC5AYPl7ogsRjz+/5BjHqelSUvquFPykA5mY3llSy0tGKxEtthc4ZTKf6DrXEs2jZSJS
eZa7T8qLpsHZEnLNoq1KRoWVXOgASFdeSyHKSRA17pLxbA1CdGtkfl9t1CfXMps24WtgkUs1tfZM
wubGWgYv+E70CmccQ1qbj8nspKEAWlt09XgLQ213V9pJx/M9bIdDQldfPnYltqGU3heqY8BwcvTM
+OVTD28mUEpdveiOcbdMugXlLRWOxw7ueVimOxsmF0F49Yme9kDiIu4lwVVlzgHEyW025aJBgd16
Jy1z6wlA4Kj3mQsbHQNlJvd6Wm8vxYOCNH9ZPd6t8kTWfl8m9uGS5MfusuInki4J6zkElM7bxLjV
ebLHDfyvLSPpkw3GG///HIMSP8UDvalXlj1wlaV4QrXnVleeKO9ospxV8oMgP/+lA2XuMYkCx7Bq
YDNuu/eEaC2DnhJdWZROvLEA0hjLKN5L8Zycmzu5SwEOKrN0xgWfGL7upkUTo20HZ+vd2ut9kSRG
tF9Mf/elTPo6KqvtHsTW/CbxVh8Fq51sR0oMWEYjX2zkdhGgco64so0l8pHK/zgHg62Awhbh7lOi
FqN3EfR6b/wN1jMC507NSo055nqZLfq5/Qk6WKxMeAGvXi/Y2WxQZ0mhZop1dv7wyCd4rXQ5ReDM
uCLIAE2KGhOaMjSH+htGnumetYZV4oIYibFaPDxNyezdFTQv4+ySLSPIm0ZMlUBwq6/7/SgzSiKe
MrZ5pzrpPsFpSm3Bdf4oPKwJ8eVn4AeQ9RhGcOTqn8aOEJBZIEeKEkNhYhrpo2TvZfTygs9bkjZN
qSbUaYZIfJaLLhtra66nJVFC3Scedsomb0ftigYcpEUFLdFRopB4vsDkMvfOCn4OGX6ot6/T5mMz
fH+fyzjXJ5oKJFq5uh4jfFKA7Vl0zVxmanL3BOzvcpWqkctoA1N/bqcb9jbgbPJSDVqI3ehDQksw
6UectXdPjbaZL3WfIINFxNCZFbIye/mYq6hB6aMbHTeItlk0s9RTICViKyNTUHZBFWviOfIz1f5m
joSo3ZbHaOoHP5+osd/NC+iO0835E9x1m/h/IUoccGspB0lREV23vcRph3aDWN8GT1geJ4LtMmFA
beas1GGV92BBoxdy274p390HzuFrAk1SK+c9WF/jotPz3Xxg9yofbrRNKxe1eyd+tdBuZpi91ZlB
ODEodk0eG1lHQupF1icPUF+/vz5ki3XbkulOsTWpC6tqEgbDn5tyyICCJ0EI6meFAB8QhZACgGqm
rLcwUOnLUPBnPZfOta5CF33Qe8cQj9/YnEFORyrAKFF/xRzQObYyoWKo7JyPK/uHuKbSpoRqrOc3
87NN+PRAQ1cwYLQlmlKh+a5OxOF1jsp6eu51UxCr8DjV9Y75wxBjLzTi2CQpXnLvvDXVC/OpBrWU
dRv+g1Ha7sDl/p97kLTMV+Q3E4f9Q3C0ssGyhZ2BpF/vee6Ku1oxs5Aric9i9txY/5qkDANESs4g
sMm51oWtH2KH9DHYPv7yBUvC990dR/YusPBCLtZ9/6M70TsNuPIXFbk3xzCgvdpLhaUryUP1whfe
dp19nv+IQLNlQKEKsBCUmajv47FauvF7WnweeDjIGQGtCwXeJAM+GREHGgua+G4IOf8hLXlnzh5+
yVz5ahbI1ChKh1WBxtWFxTHevCv4/EqD1dJ9YoPrduJR1kQmZd0kq0edJURlgipxQ3+2pJLFU+W9
aMVjXePiLSpUNgnNWFT6ELqGv6R0jmbwVVnVJXDm1SN1zNpAS5LYT9g2TNvTGruQQMHtmPsDm64A
5yJWhP8mxi2GICbynoLypFxO0cx9N112Tau3wxN9TmogIJpAGM7xpmMtg1unkg4GDjCalq6V5l1I
4udDr7ojN5hshqeki3A1zgv+sG625zacC8bTD2jh1dRUdmvKTZkABIAy8kqmdjgRRUnI6l6BdJQw
w3qP5qBuSYaSH2SUDgzNorMBS/JJ2G4bTsoYaUdIZW5eN/X45QsCHzezCEJpedm9aFoJHRp4f687
qZb8+JyFsKtpgNJgiU4UklylNh9fHhFn3L5FtQQQ9LKj0Ub67XPUjTpHqC6KMDE5lTpxQSzAZ2Yu
tZvz0Kbl3iDJ6MtYxBZwwbZLjNQvwaPbja9b/LAkBUMqMn3vQM8oeMxdse/5zbeWUue88XC3Sh0h
OY+Ouf0aj1M+gnzBgKBZlozh0HXBwxJWmiIPjBSy4PkDYX/A6499HnvyS/ZaxTPGRmww68/dRCQB
tIX321JrrgJ2PPELGPkzTBmPdGAumw+Axj0cdfIXjRaNpsV/xQbnmNfv9LsgZSJz7eqZ11WLU0hx
7TKCzcfbjrCVR4NIhRjO+fakz+Z0uT+yWM48u1rgg+PYSw6vYSiMTlmXpJkgEs1AYmqEHw9wCNmH
ypVbof7x00+8gQaybmSmtlodiD/VR3pqF26KrGLsRFoo5WsT2IWf+Ijz1EqF3WRO3nmVdsND58So
cfV4xOFCtwbjyfej2soRSoc4W6CeeXA0YO5Kex5dl6KRlRSXu28fSw2YApUiQ9g9R0BBlbpnvw2Y
cGbcIA9vlG8Kv7eoYSpM4SyGeMUpkqi8Zl5Jx72Mk55E0mR4Vv+LENU1HtI0QVgYGAD4pSISTZUj
T+4VJR4K42XzGmI3xqQA48hq4Sse4MIz0UOvhS0nY8encgVB8VPAK0/2iOayrFM7x80UrN02GQdV
0xvj1JDQerL535plt/g/nQ7fyR36TZP/LBgKdWHMeymshvWug0XR0EaVorDpQ1L4QHmnn3GSaX38
Sfdyun6xqqo7XfyUM7BhVhd9SnyzVckQ1MpwuvKnqK/g0mJ+iJtioxGMtw1hQA4ZiZ0yiTivm9Io
DkXJwXHMtTjxynvQAGEPMRm2tUG9ow3f5nQ8fCr5sUd2FyHrMDSi8vvfkxwiK4B4VezfgtBrdlF+
6qBJgdpfDU49DNeyUkojThM45fxOXhW8ElTCtYCYqiPYd69NVFh3neJW9E8lVHo8yDip6BQe2Oi7
8ioQVlXubTJailMKef+eXi8sTayN+PrZf7Js9n0K0j98puonJxxERRnaJkvW27R00Qqx7uAOx8nE
XZW4hdXI8mex0es5me4Rv9VAlTec5N2N0wbifwcT18QcVLvJmOrJcDRAXVC0lrijse+H0DstB401
EendkDPHTmOtrLzhVR2c6rdXeQT+DyjwcbquXynpCtzwHLoXXg6FMuRs+WdcXe5LLxZ8kEJyePPF
yY3gIUdvhwrfGkhnOSpggNEnEKfo+ZcJaCv2owjIx9OXip9NoYSAfjpVt7Cworw1ZatcizI/MZvV
nPhqmNCvVvYvKlGkLH7MayzQlLAkWcavucxhQCEXqH0gYK2yO94/kQ1sJHqwXtVrtfe4VJe125w5
cKS74MPwwvypj8oLYS327X4vE+b/n6s/G2pDc0VG4BAL3Si/SCrvBvX9dGwMkztIHOru8p9OLT6u
5qnQTyQlnEDpebRkn95HCJJ0VLGUJlRtkxZtPhhFmLjs2xcSxEI0eSRYT4KBpMBrUjWcVtmsYoTz
jyzBi9Cz1Gk7iS6wH0/figyCcQHgwqYa7iS6TB4wOuwQRpXFcLIV3D0Di9NZFLKlgRyy+8R6s/tS
n6B7xmWtzQcydClJZBDFIl7Gsdqpx1qevuhzbCwoTHN5TwKuD3Q+lNW3BdOTo5+cMSBnImwMNQ02
mpVa5gnTSrNx0Nn+sN3b5WpEphn05zCKAKAngq5L2XuhxmwmM0ZHz+YvHaKM8+9hLTtSNVvlYcc0
3XkG2GUsakgC/dpB4sjViwMqaiGHS/lwzt6LrhuU9FAmwYSYSlBm4tChr+d1ZYD81T5fA0F4EudL
N1Pl1Qjsdk7p76PnTJa4jVdw+4zpSs1QpjylJgA+OFfaaQwrSU0vtIpd5hil5XeOnHSEop5Mfe7y
C9JW5dny6ViazOpKnn7I2auWdY5a8oHkxYY6lGSrSw/0RQgJ82Qew9GGGOSxEOxb5fltlPJzbCdf
yRhjn9JPDuuLDz+o8vH5zkzAtGMsBI79eCyBhThT6RmVBAs3WJTC6Tu07tmwEGbjQI+rcSz3D5ra
kbzEVcyefG5t7DzTQ6sID0o1RwrKEYFrZAvqcNHSzxfYaNkKIZz6VpDY16MeHkP1GSSPH9YEIq9/
eAk3iexsOX/pER4npE5MjFo/YWD9iT4TCwRAn2Y3QxyD2UBYvQ95Eb8cMFEz9OZFmavb8f3v6HW6
u+H3bVMYi+K/S7IwN8ExFxe4zsO7/RnikHgVv/Ykal2bDNeRedE30skhLFg195+/XzWf6SQMW7TZ
om8DxrAj6dhvA3LxTXNScpqCy6oaT4AnWFcvrAeJFOar4n0Z+2f9rKSf4KEusb5gecqwUDKOyBQW
T160vpUyh9aYXF76RAhom54x33CfyFSkfSVmOBDFs8UfTaaqT1Bt5y80RtCnZB+ftkK5NZRBR6Ak
j/or4zxzFMiqN1M0PF9392RE6QzfYBZ4byKm+Rzc3QwjYVkiWbMO/2rBQdrlcpCHstpCXYv76hsM
rKQQfoJjNYz3tg/zUEy4+iaJrv8azaNGoiJqKVJvJEccduxLM7b2c4OJarXJJ4q9RaRzWLRnSGx/
A6E9dPVasVQSLzu+aUkdriYWrUZseWacYRbKwxGTsaZ21K1ode+1QPuaFSNsWoRSBI0w9EXFvwdS
Uwnsw+nGI5GEVd/V3qN9mBhgub4kaLywOS/aFwDbjSIEjoydWauZXXzLxewrxnHLBbMOdBLSQRuT
pOOg573J3gdQh2rGI4m3km95hCtkXfHr1gT/X4K4sT6zFfDR5TlUewwtEtUWpIK9mLZvGtrirfcM
/ry/2PDAIiLZRT5VQEy/rnWDrhh18H0s7AK1s0qz7bywWLDRmHoRO7FkxHpKklLkneujPw0xIrGm
4+NXwjPjATMi4I5x3vpO78rabJOsdrXD1Xjk77vbRhNk4OlCOV+bjJgbcIpF5E9Lnn4CmYueWBHF
m1sDGQa/DwM2e4lqAgwJ92XL9wQGX2S2w3zZrGmHB++iQOQdNdSswjO8lQTIT7UH8Rmc8POmswen
rX25/x2DmUSzcXAfCIW4qKZ0tArXpr1+BZsn0MLNA793cIZ+FQexU7ae1XQnBJWfgYCzZAk+RxGT
OTaBkKE01OCIl7tMLfqjR5ZzCtAQOTkXoaA3JTMOldR7Elv610o74MUDjm1i26o3lxNlB9VtT/4M
iDdtI/axU8pebyko4pBX0sWsIAAKcHYIe0gxwh6ebwa7yInblcRh5Dd/BpV1KatrcRK/r49THNj2
kWQFVc0nzbiYJLH4B5MIQwKIDiddtaah3yos/Aj/8gKtjR/G5pgT5eCu9QYSXbvxR1F/haKpna24
9tltdbzQ39WNYaorsp/rnN6thYJ8KQ4WskJldmN94LBr3OfD7XwtlXkkkM5prD/16InNmlsX2spM
qexc1aSkPRyvLWdtUBpNqosW2YHdVLv82NDap1VVis7puMxVgwP6cVR0zIRNrw2itZR/mhAEJ7V9
PxglX2vZTZvVKR+gtMqUxYg9SfN7o3A7F/OIHl2svhYUnixqD3npj3ev7VozFaYJNObfnacwkuIo
qc3IOS3ngurtpE0j4NnXRwy3B62BC3EkiaQiT02rZLOCSXE4DhIjXhjmCWs3oDhVowtyuqiGuDRb
ovdoFZLlKtbBBKwYr8lvpRTg0q2UKR98DtzAqZ39372oJYkYfuV9RHBPG4tQ09h567fGC8CLAMx+
+AM5dFbtJ3bDF7vCgzWCV/zRFgnt8M3lE67eKaXSOS3WVDpzEZNYVlZ8ocMB89YONBPPrGbzsrGh
18TUA9Zd0U4IlDFsUTKSh+TGPJxdE4vq1dmpTcN+FzlpaoQT1HYQubf1b+guA8xup39wkiFWlMSp
DllKCjhHLCpwLClHgupX9fM9/WOEAVvNclRtnlkcWRRiE40XiruWoCAN8eou4B12nk0tQxWd/nfL
4goSERI+jmwgIslrK3/Qp8OAcY7qzCb1Qam/i2TvNv+Hb7JVVGPb4Vf8XtPXe1p9MnlrB0xjGRD2
dhuoJXEADuoSDO2niTuPbawxHfltvrYn79CjqSzzMnRa1sKzbaxUDw/IUupkkGl+D4PcJbPaVJ54
y2avzF6DdB9Z6vzfwVs5hkOcwcVBe8ohCFgsfCsYT90NgnDQNtVYS3gAEEwWLv266MKfziPP/z+Y
2nY/yPqZ9sDCg3o49alf5PVhEc3EkVQAO/uA9fNOuolNL5TVdEAvJUIpYcV8QzYJKHmeNM++YTB2
WyW0rR7kUsc09wZtGQFHl19olsnKsYbls+ZBIC/70nwGHCNwvnoz2lSwQ7/guItfBLeCng0s+8od
Onb/PAoG+gp0cRrtTZbmEiQp4XysAC7nVju6bLmdG7ZRz6oqCrT1hSx3KV0FuuUxJfJ8J8lkE29X
obf0mnOw43Uv70G5lnww/Q4nsXCZEWofbztS7YND04TX2r5o5NlHMwIGTTku+ttSmlVOb5DAPjxM
kl0UbM6gx0LtUeuSQqGk/VlP8UU+CYCZZ32zbDdrKcCkULYybuLPfghCOp3O5t+FusGFsaGMz11r
+RUd/LR+fCdQC56YCckqGvolNN2Vp/jNWxO07XNAdTq5NmWbU0YTugXuN+1cF/UVAwIkQ408DuaU
ncDkun8velz0wckxioamvxMSY4j3QEDyJYeH6uQgaA/xV01UFqCh7UylikZoLcOAoHfaCMgJQQar
qfdpDBCuD9Mf8vJAlAa3epsD7/uJ3oz+wAFsm8QOskEIGtZ2PO7dRhDitw1tzu7sBd7bPos2wwdq
yxqS2hlpHC7rs2TTC0JVd+FBQSZfenZj+hQFG22CBfLXArN44VpUZUD52B56DmqB9GPJ3cjXMd3U
IydArbtA1gceHwHFeE1nvJKhHVob5anhp7TGo4c5lL/bQrj91RZyiEFO4SS54nP0JeYkMfIbpWLJ
9Ynfn44oJNYkVoRKfkQsc67Od6k26iqXn3YcMUweWJZrBJ+IVFaA2aWDi4Pmpsl7f2qwj04jHmr+
V2tdrhrLmct7nC3QjBi4tWdMo+zjbYqTEFVXVjexKb1BEHcy4ByeT1kaVjNnzxyzICG6T0geINwV
bElkLJJTSM96iWnvVpstMENDEfPoLMxb0CwmvVAS0TwIVhvCFN/Da1SuorgTeNqr/S3K0Pqb+hvk
WX/7fT5RUet5qbyy5j83qtENVrXi/1mBxVUqI5o9Tbl+MChOYwgUNjFzwh0leh205J8GPfuuBkao
4usowz6SrKY8XzYafDtxyclnsyD5uzNCnuHArcRjlz1YmvImawNUXr5uKcX67wrE1ACMYq/GW2To
RVJvisqJVKITT1w+BNAWao2PIXy4aAvK3Shrd+sOwt+W0SeVMlCs3RR4IFcQGo9IMriUE1a6YvxJ
MnacgIa34enHmPnPpIkjkpqkp97ZmwEYynVMg6VbSWzyPPAXJWJDuV8/q97bkikxNlOZbQDqHGid
en+N/1L3wOGnOTPC/+NY7I/gYIRcf8qhW5czEVZL3/xygKsvk1TGxVfXzK1u9COUnlbOcyXUJH0Q
lnoxmH8HP1Uuo5JV3c3LxiudLNysBeYwFKZ+02F9e2l77Al+5fHYBMrsn+poA4CMBszEfw7jxN5m
FLVIjPLQbpa7hvsVmKa/6l3V/TbEWOer92AXBygEwlYIwmJ3jRz/yI5Q6hZmWVRGPtY1S/UyoFWQ
403vkPAVNuHiU3cA66z1Woudm5qag5/668R+WSbv8kJxNQPCwD5pFdVWl3B0i+ex60BcYt6RjxzW
lgKsvPi1gIp4UPqhn15+Q9Jbgg4uABV3n04eJSdf8v16rdPWoxB5TIqwM2cUz6BUtytXI0jAfbXJ
iS3Aaif0ke62v8Jloae6HBXknj82l4Z/rz7dWve/L0VGmRmIUJ84ahI2zM5YunuEHLgcjeP9ZJWN
om+viqER8dEouRJjFSeBpvqLbutLGKzajeDiWlx2V8y8mCZ1VOSkiHGBYuLpOQIJ2X09vgezWwqB
QwKTFSeGOf/vLW3QBtTmX8Ei15Ph+XuVER20meBfOHUMa6tFEHyZgZ/k4b5/nQMe9EiVawvY/8+o
md4O/4PM4kxaSJZaFJijqveTFQ7Ba6XQ8fYaC4Zb6jmfROAr/43e+VW1JxO2kFunsmKcpB+IR3us
QajpWJB0UW9viP4s3WTYlVPWsdhr0Yktttplogv5r81puORLZTspm8aASqjnbL0/YuC8vfsz19d2
WUrVdaEPj6YIrZNvIG8UvUdG/sJemf6JZ9t8TyZnF8f6ck3kQE/RPGwlPgD1NJhM/2btTbHLaAuk
PkxXaEomFEc3BaS5IKLhw58rrLXrXEzmaLQRmeTzfnyNNtZesJAuwevpvPB/ZiDHiGy0ohX8Il4n
o8IvRmF72pcNx/qJTRKB07YfxyKbYG+V8QaAZdaV+pT6P8jgd1hYDzv/T5ywaaZDx5sNZYjdxbTx
I7lAg591MY2jin92RPue4eVmCr64cW1665MBlJvYd4fH02jz+Yy166SahkRIoc5QqaiqfR7p7noF
rM3/eBuYvNcoFbJMC0Z1cVoNJBFF4KqF63Zy9CiYz+JXHNfTS5k4ESyc2Gk+ZY75bn68I9YDiiSJ
qLCCocaqgGrCpyY+rqbwu5/i1cixGrXDVVAVxZr+0+PpbGV84Nt5dIBB8egunCrustvzTq3bW0yz
yd9NSD7aL4T7jhIE3iL3mJK1YmFArPbHJ7x9ulYLQiPAOyAXDE0ShfEdnqQi/KcQnxqmttGeQFPN
PupY4GB86nRpYtDnZkoEcwELaze4JKPxvp5k5upc3DdtAD9tkO31noM2tKMWFFXF6g9TxlsagSjG
z4sKhpBwHsx1uIGAaXwpcFJ9fq87uuM6rzc9Hgs1t7pMiCPwMcnO8NrqdgB0Yn86HgvVH4+DlbUL
RLmcpU8BqBQNwFmCIKIy8TcDjgz/0HcdTGgplBi/ua67sLp2QmnHJXKk9sMJKqRqcBMA1c3Geb5/
bewHAR2c1CkY0M0YY5jPdJAHm/MNhugPkfHej/4WTC4zl0dttxAMuxNDLO8RDLL7Ng9nghHM8JD1
7Zpb8YfmTWfuEUP6XXaybdWvVGteLKE7jUDnmGn199Nau1DHL/K5rmM0SAcO6Z++pK8j/WoFMV8T
FC7RJ/cXZrJu6fbzuG7CqUvUreSVGFlG/7hqdfn7xMLtH8Cw/NqmZxd7PFJCNirEu6CNAk8mUvH9
Hj/4YP6cJPoeyAgCZL68KE9dSXCr3eK1TFSFiH9SFKTUspRaBr/zF5wzzg5ok+ZuhiGWA2j/lH/m
VTlo6gsIjcBBv7/ty93AjJx2TUicVxoEhd8MMujsfBnn/EVfWRB2UwSrSgC0MMC71aIVUiZPobB8
wJYifxvIgmEzVWoagvF3ri8Oiah6nL7ECt5TAqI6s3SP4IjzjcwPsmmkMjsNwGqlnOk0hNV7GebW
2VBTu4lNvy1RbR4FDONM1+vxE6DOcWHPFYvQw0ddss8AWVDud99n/zR9enpTGhR7qr4j1/5lx8Hi
YohYjPWyP+dgJyAnZFyC4Sqm9AfaO8Vjyl3s+ZFwLPDtK8vqfaQJdLURJKmdDo5sGsUD8RRSKFGe
21vs1w+mCOcmcrvtwPy0GBtMuFE8XnltbrRH1RN2Fek7yRg0p1nQP0rm6Z+G2EHHNVW3OaREginH
85Piq++bYe2jo7/x32I71L+GnY4gUCDO88BxuM1MZGBsUwS7JG4j6VTDNPeZXH/20juFrbPrt2fr
xjWqFvXodqGvHGd5M/ziYv/dACfSB5c7GD259DhraLNTqdJgFA9XG3/7xCZQX8e1vUGNfBoRSbs4
DPJSNuF08bBIgZ2O4zA7l3gssGvj/2Ozv+IspKcC6YzU4c//EUmEfkQJBPEkAZPl6sXkiTMZBurS
WZ8tWbS4e/la93GXtDazUtl52Yq+xb4DuoIwhjY4rdytrro2dvXmO7/KL+8RSgNWY/gZoXta4Qnp
mlqYAxTS4e4M/7iuHW08/gUfP5e00O0J0NVkJSn5SG/95RCJf/kxgyp59JPlRyuh1FtudDv1OzC1
anLavb6qIpUF3j/H5atOzWARqgiBDpZo2nVbSEA72aC+zu2ho/acgmf1eBYLkVMaQ6RHCoxxB3Iw
XVGEDRVx/1L/3tWfLynuc9p0GVMmebybWR8/lWxsm/JF/A2qBUFr0i79pMwIdqBiUa2KmTHvvV6k
FIZiWOIWp4ewB/J9wgorDB5/YpX18sZc7EhK08smJ+ISrXz07mhf/3B2YdQlMtSZEhg4xa92rLDb
RdNryaGuYu7aRn6R7Mn4KcJr3LGAxwBvgiHebSCM5mZSzRTX80bcIcIn1lWS7m9zY82nN7jpyamD
m9oJy6fE/K/drULSPEEbHCDG9utlZUc5n/z1RMX1zRFOmkr+nVmDEEDvEZOV6rSe//HDOn3qy2zK
qP60bHEXWiButl/CXRNiYFMP2/ZVUDgB8kvvCSUa0InpI/iRcj/XNT880JfyhNJ/vldPXaSizuoR
FpKPmh3iQdgFrfZcRR444xVC6eJgwAmc+frnz6VCdPzq+EbrZ7Jop59BDuRN2z7dqhusXH1f14N/
bxac+pf+Xn9sNaiIaX7/BxEkQCj/2BelDyMFcjH4jyhZimmldFRv+0wzcAMV+tViFA4A2QGDMMJd
1s8ASQmhtg6BeFwgCoCtHR0BNUY5A5Pin4py3wcFQXEJj2ZNBPO/BC55RbN2Zp8kamsAxR0CqV59
zkH+vyONXYlpePbKYZALwx5cCA62evUQdwJYsHiliQ4XyZnvpF2oif60fRpMBnll/gcGyiBXNvEg
Fe6W6jU20WytTFXRV1itrKZ4wIdBssc0/eaJYyHObf7lLRLOApQpKQLPNGgPXXxfkuMpFVU77hGr
ajPYCLOiGWfwa2cIfzMOabOaQxntLQLhb9/cISVHgvwnVje+74qyL3nniMEX0ky0GVP4EKNbzm5F
MDVXoymMk+t/tfTdS2K4PhAUIR41zf/x1nLvwz5oLD9mWgEv31ibAHErcSM5I+z0Sttuf0uETs2A
H5h9Cu+CUDCqiky3uCCdEctD+70fXBSsx7M5FiVj379ukvP+fScBNbi37eS2bj8clSyKhSg+/Soh
panIuws6E2pYjXYl87L/73WUDpoWKWXWjyeWVxjSphaHYL/guQ/Y7PYoMMRJru2y+hZbbhUzgrzL
wwG7MNd7qLCvpgl6XZMT9YZdgcBpLv4uD/31fIKGkP5GeWLXA3pEbrJAdB4hL/n653vyQSUyybaF
mc1SE6EaMkqP6M4nIKLmid9tvuKWuZEi2XwWJpa+qaPjSlbCic3nJorlNRN7sJ+CtwV7TCYFNRWR
lZvTRdw1LSyuSfYfnWXHnmHSgf/OG9a/Q4ySmDTeQIug8UsvIeaqKMYv2Ol+V4Tl8oHNzl5kCsIb
0MVirnQvg7JSS1zEAJTv0iO0Xcl1qUfe5v89qNWGEKQkcTcgmLg3mZxcowTS1PN0L/MCFKbdjHqi
MyXTxYfACoMKkpkvFFWghCYeJs/1wzred7aq5xd60M/rRy3oGdffhr8+odFm56973tW3vmiiGDsz
cXfVyR1BqItQ9x9lpwJZp6I+v5hvXTbuZ4nT55VtzjFABmvKMI8+bL5FnEDAcDgrf3t12pwHpjfI
moRpsY46fLRAOHKlCTPZRNYyjFP/gKQXV/KwZoOsgc6j2FsyPj9qo11/DVjKxKqZSg5J7sEF5yYh
C5hPMY4rjOCQB2d3X5SiiWKfUB3diBjgknGA8DTbhFAbj5a3oGtqiBgL3ZItXgm2v/TwJIO75ywj
Y5/iYv8rSaayf4xfNsIO0rO8b2jEZL6ptV0gCBBebwvuaBbLdFgCer+kGRRyko09cK+cY6jrIWni
z7FGQnQTVwzmHbsem6+dhLiw2zq+FjEwN+kbKKFcIpCf9/YUYGWmP890igvjkUxrvlNtNj5f2wGS
nT6nx2JQ+YaNzFIZ2GKUwAU/WAcCWzEVRsy9yjV1qbhIaP7WpAyMMxu2Z7RKU7/apG8ndso7BQ73
dU5ngV+CnoEuE8oCODuoUKSStxc/OGRZrd4PNE02kgGxb1jsAkL0gfpYZjeUhoiDvnx+Ih77xUrn
uE8PQxmy+0VaDSaLmLjl2T5mw+0sBZ2XEmQ1LVPoMzuW0UX8ZCE+fNKJWLRuBPzF2s30Kz3NfX1A
SjyWeQ5JrOaFGKlD4N4bcgyZqDafLoNyvxVGX0Iy8UO8ZJAG4WbVaeiNGzZeHQXs9HSzqQTb8iDe
yBlc9hUFjW+yLHCs14h/7kn1QhGEmxFYM1OcQaIWt5hiti8zzcKUIhqZJlvGj/K/Jp/XgSJX3nMW
xnLVVhXIR0A/AUgkdDs+u4sJXD1YDvRu+i8rDN1oCfjeiKckcftZcdfEZZOs3ysXC7MP5Rux6zYa
GNP2S5Ftyg4bXV3/0fxjXLQyJUxIgiSYJdfks155o+Qfjxverjuo8ipuLgh8ksw6TwqcUS19Zwjf
4QUF+jB2+hr5CjtmHbtNi6zxacgAdFe2bFD4WKUCGeu8ttsS5FrmlXAe680RZ2os07XhMg/t+Z3T
Fp9urADuWBBuqeeaiHAMiJ7jqVTtOFN10n6ToA2eyGMZge/ItdX75ZAMe5Z/uaC+a/Q1V4Y8Od8w
yhH6oxh5Eg8EIjc4rRqsRA29021MlwEngfFQfGJgSb0vxtRfERw1hMPhpAkEdvAM/IEQCAvfqFly
xD+47EMg7EvYFW8SwE5Nxizm/7qvL9DqQjjaZKCm5Zruo+iAvl5SXqlGrOf0NGRyfeHiPnKVXZNj
0kwlEt1vaLAG9c2KOqH3ePIecwSyF4l8W0HUKFd05Qn3u24I2VwhAO6eWWZmSjioaQQGmkH4m0nJ
s4XTHOBr1kpjS9mJ7iR/DdIaK5vsSUFy7XP9msSKwVzbm1ZRUFtGtey910GO1bf5HJStnbn9QQ50
aI662h+hGuApj1TN5wlOIU63/74fgWtNV7GexIFctb2KkPoOAI5Dnh+74zxd2a8TkiEUs1Q3dtG3
ZhGqo7DCnR7VBt5OOXs5nQixAvIis8H2JcDA8LZ8AEZTiM+nTRwpjjpeOyrh3zdW1C4Hc76f85q8
sFFpETSqvB30pQhatpJWAgXkJaa33n7LIYV47vXPdKAev5/Spuq84ghcRPxVGIhXfE2qtw1L6//t
HCuRgo6oQ40EfmTgi0Sf2LmdMqsUjIC/xzQruhZY1x5+VxGwUxrgoXtPUI+QW/AlccnTdHnuNO4S
YF5c4xsRg48n0xKGAwxma2ASMci6oD0V8tDU9fnjU4lDzZsZ4pjQmCtVXmh8IxbK6RP3cuambnPz
Lm3+Y2S8s/VbQzDqMqT1/uDSQe3MZZHjVp0Vab4jgmhqnatYKKh8Mc9+08iaWb8Vg908VqXHe6GK
VjYFJ45XvFF/GrHkdvoyG9Q+nMkoAKWJ92PgWiurRveDdNkayKZ2G2a4l233bOq2j3bWul0rd4Zs
kehzYgREow2ITeMeJEAfzyTv2U/y5sRglXlCywFZ/IC9HxFPsSvAXKjkYr1JyoOGKfnUe/Td3C1I
W1G343/EkPfwPqS/U9lMcBNRUVmuVeXNtJH5mFNyQhO7oNckd77gB9y6jnMBBGeFvlzoUYgQQy4h
u298BXAaQcZfbTKyigX/0a7s5LASnPYpoYZFbkSo9ppMVmIAtfMqoGqwJlPrj5qCvIQtVai9SZng
Ew856IaniRKx18lgLYsbzGBr6im8qfiffJeVV7DsGQ/I8LZfKKYFqlS/Odn8iWRqDaV2vAGSS/87
k9GaXaty1NhFe++GHBTnqB84jc6Bi+x5ym3bLHV24WUSMW6acDCaMfEaRadfAf45DwH1YNnHAhDW
BkWOkD4CkWsAGmrdelyu2DOsvjUN5n/TA2j6MkZ1PoPfj3BXyEttzVE91eXwJ3DCa8dLcR1lxeDs
/wnqVQPY6nrkf+HV8cGdofvOFmKCXrUIvqrTgIPxazg86DRrw9lmJii4jmtUt6zEx1O8CYjucpQl
RJB2WhFxBqbY8z6zy2/LycdYkHUmneaP7bsY1mi4n+hQiPSk/n+qk5a0Kpa/HKfeNS2i3dVNW1ix
SNeN499RTq4afqsC6WKwp0tLpOUHbQagBLTlT+m1IM7YxE5ywOyHWaG0VarVxzp+VE+1/ii0SyTM
6TL5NhsJVX8jqBlt08aCVnHxMuXaWbcEmYKgekOB6LdQGmgq/sooMKSLC8mklQ4t+eqxK/l8zYjV
F5pW/8seqNyEtWwD5i9XA04anQSLIPm9Ld65ebr/++/uhGj8CfqxZCVJlalLzLxvQk9QtIODJrUO
HvAvffPG1M9uTZ9UFOfMj2OnL6Xo/6xrQRQXPtH7OzzFHTmkVmS1KClSxvNT/ky+rtsiw23QUI3t
HQbMN9w+XnOnRwCFveVCc0VG2R6BHvEDCuH62rA3u34Gj9cc5fpYodMFGEn1iYBzY4skbU18l7ZL
17FEalIx8yHh/x8I45ohmpiRJym2i25gzqIeEfifcWZkIk5BJi4+yDNdhf+2xj3L8S+Z+4vp3ddH
VQuUZtE4CuMhX75HzKYA4c/gh4ArPjVIF0+OPuJKd23aaKqzRyqdBuYOM604kBbfdqiDndKnaIWI
F+Uo0SIZBAt4stAJs0CjwHhRf4N/Pdq2HiaD/gbWHi0pUhTlF188xfXx6L+TfJaQ6+9JBd0Q7wh5
7zUJiIRaastCQZQHL/OyKdhqi7aqu6ElToaLkqXU4Pe6FF+SiVTmpk1oLe9xCjDF4UJzFFrg40IK
qZBBfoOEZKYIoQnaxrrd4K4P6ebKtuKlpvRkkLq07FYfRWNdkqqp25SZhIPVS3MVHoBS+cDDvk+j
bDZcRbil5nu0N3pD7SXrm2FYpElc5Qoq0mhkTLoogbG4pFhXsgW4Y4Z9pYkdbXfELQ+ve0YunEZU
Kn99cw/4r+zELO+SMPcB1d1Vsnfjk7lelqX/Ns+XG2vZGD0GoHGTWWWxS0JpAfD79k5eGn+8VTf+
CGkLRjILPfn8GIl1xB6Kn0McKG7K1696z7ppsDS5PuyuEbluoeXsmiYlQjpsb5oEmCZPBk/VLsir
y+7va1J6z6Aw/dk6oPUBM7503CscJI6XAmZAXwq8bM0tbc7iOPeSmuKmd8dt3jpaiWdkTvXfIM3l
acQfN/cdbPD4Ik5WnUvCunlJSUNCdBJjzl/rfJFQ4CfZ7/G6m5t1Tsbd87h6OHkwQzZ0jWIU6X6Z
WQfYH/lGM1OqgAcLa7RAyItsuBZ30qxzXeW7IoQZWN1HdaCU87b9cSpjLZpjEA9Jh4JeKkt7Ucb7
Byp26GzdhzHoYQlaqTCegtGSrz3p0F+1z+ub4Twe+WlUo/FqO8gJkdw8C3l51Zu90GnoAZtsZojc
rP7ajKXegaDugfeQ6PhzDsqehlPED2MueyvhY+ZuYBw/IaOpdF4SOtte7Af85fXaxSg5tPq6N2Sv
vEy+KUIz8ECAfB1TP7TFGKqxVipf2MhCOs5u9AQJxvKfjuuk3DecasNzhaSRoYCqRZDaW2Uw6IPm
97gRQuUYQWc3t9yO7sx04HkQW+TXmvWyvVdqHW5FjrB48pk4Tcp7aerZ79WIGgLnPb2o3BWLcl/9
kWztLgjAvx18D3c5mKFvVvGFnCpiDECltMtSj+yljWoI8zgfRyojQWgT+gudRVojjzFUFgg/SAph
PPHNF7+N0ZCFDyeFO51/I8i1pkLzFObshe3653dqYqplzclsyOrU3ANPzap95VP4zyPw+KdjP2Gf
yXvbyQI3B/HID+QAJ/elqGwTVYlZ2VdS1XsxK7HylDwxMg+NU8JhDdA7E6WONmJrtgnpmFNJjwec
LBgXuYl+J6oN2cAuQTGj3AE2IbpS39Uh78agBT4i0cCe8vsPm10/UhQ1o2aRZ86pa8D5yJM8dcIx
S4dcPxOjZMDPLF7GVgbhZ0jgjwbISIywaqKZZnmEomyqt+ZmHnGGy3H9Qc+hPh2HRX6L5H7iBssw
GtXvEV153OMRpBYBB/D/sJrwFIkgGiFs1FCeK+GucbQb5Vs7mpfF+ct1AERhr+UfpHLkF5vT+DCv
RldVfkuX2KUwswYaevlJMbfBLUdwEhldxj76U9pX5TZNCzqS3rWP6ZYcpw8DrUcOERswuCcgrNN8
WQ3O7aFlBb5ke20YHWGaMvkknf1r/toiJQD0puwJncklAycWI1L36H6gJ484R+RxcTZuUJCA47Za
VIRDoQkgN6Y8DIBj2EkLHcOvNkP3guiwi0mvw+4FK/7jJp4fECFLCP9wl7fRydJYee2Na/ntgOHO
UkCpmipbdciYpRP5nCn05a/oXK77C3b02oeBGG+9w1I2pLUu3d+jbIwkzYuZ6p/+0CSVqwb/RKXn
Y3VnXGuWlixjCJBE/g7ashfZb4Ip70+zseIbvrTGVlFDpgoz7h68hpMRnGuW4V0s79bDUVQ6uSzb
wj4qiLZ06YXAwCRZKjkd86PtOL/OixcVBBNWfOWQIXgXMfV2sq/1yiqycesXK8zNf8oUK5DuwBKh
8cKnMsepoUAURM3haSB/tiC7ZBaoWVnIUxJDxLxh1KAX4FKo3vDT9dDuVsdpTFqn+nr4QKnxo4d4
v/NHjXKDkrt12yVahRA2pfcwP1O2puSQZlqEzeeRJ0QJh6Y1zip6X63ZtAjLD9BsW60cOHoROjDQ
PZzIiZH3oMqJtMGbHFhZC9MCKuWxkrDs3W7N6EzU++ElQhS1QYJbeVhPe88lmviV9AT/BgvIdOif
bgUwOV5fS+26eMqF7gSCpn+pp+ujEHbDKHk0axvYWBUNszzkfglQ4chTk/mbL8EMc+3z26AZnKJ7
hct7+Zk2Lv316Zadu52fKT0w2XYhCYVByoye/SyzeGLoRzbaekP0j3WyWapDnSedQHuVsQZ5IQ2Y
28S4VVXyrd6VCMfh+a0BSa367KdEH0Ktyvc2zH4H4ErzzXAcZ39vytU8GiRcGj4XSqiY/yq6sa7h
FijEIg1+QepRStlbDTgIDqh74RKk9l23LvuP0zlfl57y2EiUxO6Nme/la+Lx18dq+5soQotaSURk
e0emrZvBXZZ230Ams37wItO7NbOMW5+q8wkTsbeN26jTyaJJTBABykgJ4xx8pmdEEKkRplq+haqx
JmbIUoDiM7//aKLCI7sJT5QrEUT901mZOhti8fgCvrjxlc44Uejk1LbDQ78c79kmJzP2nJiRMiz1
+q1ppzOYfl9G9ZoB7rdCrwiLB1siybFV+sfisJDsO3e6WB/BXRAhJ2s8j9/QcQVZyLy8BpYlpV9+
r776Iyu3g0QiHdlWuSjOTIUTKz8eyXhnMEkV88vkGXvt75A3iu+4mAENsrMwXGP2wFxpCHDNH1sx
mJKESg3zfCBHCSyNIziRfLzLhFLwTdpb/uHHaUc21hOp8rn1oc4Vrz7eBaGCCfIbOG4LhHDN//4O
IHcRxkfmmdvCbMkhiIdv2w3PA61hVJDSOUOh6+MgCXYdQBAqu+hNXcRWF3wa9jSPxheIvFm4Fv5i
TJGYqkGh1K5ukabczLhYEF5wXYhXCv04aFvh8PgcmGwOkmPqUYQaTiL62WM/hSToNGN65utTrZXG
5OBMlPleIJsAqnymIF3NH9c2pzNVFu4cHKN9Y5iAYpfJ2dDvsWn3tfiPYVqV7Z3DizestKDnnka+
TQye2ZzWi+l7afoGOQRRpRQnVv97CtLHX1WrgD/3rKlpaWxiqyx9oYur/WhwIwwCaqO7UNdtYLzd
X8+jPDz9kFwJiU9PSPJKeOFAdrHNhytjbMLnbQRaspOhxO/1Rxh04/c/pagtyHzhsrFC8E5z8RnS
0vXp3P2f2UuM/3357w9Re0iZRMYqhMwF22tzWw6b1uJlv+UnwfnoMQENzX/vfB8slNA1mzk4xbZB
b27CT8V37VnM4SJ3TXek2gTRlm+bYXIr6p62r4kB0ZaYYN2pcVqZiGIvYp2Uv0+zGWQ+YAo2Fhme
6kn5HfqJuoyWpk/PXA2+h/A6xqTCXYYmR2k+sklSjpoz5HPnV2Myh/UYqwV/aoWtTJLMkO8fsUN7
sXNkKTHPfg+qgULTmwIUznQMQqy70bqS2FP6U6ZR55WP+sDVkGQmXYrxESSe2XR6sl1EgYmY7w4Q
vFxfO+xGgGG1xvcHR8Q2wbeiuJZeoeHEJJLQoBMVDuCuQbLMJWeLy7cKXaC7R4lH4jT1YUYTxtmU
q6gFd+AmT+QIWjwQvOOh69TWgFxuguLSHGFblGA2rx6S3NE66hlj3c82HiOA5g3XjMHb4oZQMH4B
bM80BrX4obaaLzDWFt8rGEEh1vWrfKaND/BECs6crztPqVHi79CN9jTUlh8jlvVgDk75tqbU72Uy
3XnVT3uFM/otLlNpxF7q/HByRGj7B3SvbPGT5Xmn/P0nKlq23+Fb9HLEukX6a8nu3g4h6lemOqM0
M5NitYRdBq/fQ1pstcn6vB8rw++LEuAp92w/62m+N90qNFzZqi/BEe0ZSys7jrLAN4KjWQzlSpoR
5k+2p3AGWJBecFBlrwVeOLavOpJ/68feiBqSQzgB/TwZAt1u5YL1NK7ZgspaEdhk4OveIFYTBEXA
LTlM392oUsihWA+cFghyO1daLq4TQQRELf8Ktx/yWDk805Ik7Wqcspa5KA6PWi++HEHiuA9czgFB
xnaqr0bxQmfa7C1ib3TOfxz6zUgzZejNmsrdpy6eL8Eq6g0e3i40ROBxsqZFrvuhppDmGG15l6pX
Ny43DXs7m5/t2Kd0iJt/FAWUDDhvzRIvc0n3YY4Nd2n6ATxubPc2bYRPJBFeqTyeVP3xnBZMaxEy
6Ql0cKjAAZAFhB5rkWcS3FpndD5dRuaQPMrj7loiIjfi+pImeFUzcEj2G4WLx3Ct+WtL+nyK2Hql
jPUwJEnxGwEByrWuRd6Giw1VJFDZNc1pHd9gaWjXYH4R5uVkxiY7e8w49qibZdEBSeCcjmds9t2l
LQu6FazogRQtBxzzVBBVlWXiFOv0F5sGxwF2Ff51EC+5iSBKSs/PVJvIeksEFK2ZTadcRQfWZyj+
nHVUBgJZSz/3D0yHiG9QPZsFKvSaqPm4AA+CUCMAN4FHwqFrolNeSYOSHw5SW2e/P52cpTJmEIHQ
gWKCSgPN3DhB3s/kOXgZGC/SQ5BcFP2b2aivNzGbCixR6ROHuX8pUrfPTSY00JlVvWaanW2oEFJj
EhxtDSE4aMRjsboL3GBGBZMEDm1/P2aTiV1lL5MJD2wbBsQVh2rCZI5ZWS6KbHM6A3X+L3eMePsM
nFATDjx6+jth65qGiDNQqzgK/vxMfTJXcFNGTUEKp1UMvMzfUBWHI7S+ipx/uwq+ccP4Tz5pTSK4
6osmugWNwj7jirsky046VbrmKXS6sDJnYRQoU+l9Rts+qwRtN/qqCeypb6XrSt63L2isLed33meT
43qzH81fOHJzhwzon5hqnC7tFvMU5as4j5pK9+pd3ZwwuFJJ70CjN/6SqLASoa7dZXADfwBpT9VC
JB4AS609vCgWJBlK/RgFpxpg8zLERz4/gOdkA8yPmDo3a2h/f0TfRd70rHMnhMi1pz025Fa1LNs4
ceFkhkFN1Vv9mgUrGvjFoqRl4vF2hYbvCHOTNm6SErRJq1/9DScCxkm8w6qPavfvpk5P1Wgk81dQ
J+rHdOR1uzqHIBsJ7fg9GSlBD1TPceH6z9+WmB3n3ogkMsYb8YEyxaDWB49sBFh9ponw2rw56mWy
k3fcIRzSURZWvcoPS9NNGlptEaEQ64bL1LovOXJegY1L/vtOUP+DSs1HaqNUpPA6i3vDlK5k7mXz
G9a1/XviCXX2lpFS2TU+PDW3w9qNWE8p7EUdybjqqIwYnk6FgWt8zOf5w2dgQ5K1llChK0LpWqUm
BkShfdpQyzj+4SHUc2ur6+GhZiIxD3qqn3y8/GXcygfc/79EYcLR9ntsxiLaznugUGl84xUQ+AMD
c42o1hkMsUhrOkTzhbCAlk6Ky0YUDQ8X8X8hwzys3gHW1hT+LG2NdwdSSPfOsAASIFrh19mTzwO4
hsCBU1JdSuoKanJYhLsQbVVusFTwM5qROoewMFuRnETk6unUWorHrqOykL36+ICBifBjdrP7GzyL
QL6V+1jnFtYGsPJBhEndkCjUisRihfzD16oKokCpSPOTY6mcy8iGgGdwy44B47L6kCkAoxGpJwwL
VA33nHPo11L2bGlngLt7Daf4AsH6hzKgDKNo/IAoT11d4W4a32nyobwHlTq8/Jo0JpGO8/uKg9IT
Klzi1Mzw43ZsWeXRNdt2wLEHimlQfjWwEY7g3QnjxLPLG0vP1NqNBWYxMU3mY2uSKFMOgx6i99HZ
338n2G2z6wEWL1XkX6QeCAbyYFwG83/jdg2uikssd0n8GGztTmqfJzcwpLVfv5u37dES8eVh7gBQ
rD2mmOlKrBpfMzkMs6T4e5r7BpZmfQ6gDNg9ZqeM8alCbIa2Y7I+Jx19iTj0QEoo+raV3PcnrNzp
HTrQpkFDvt5gBiSpyHIYklgxMBX+5/Ocnn0NUbuH4xEnUbEv4IOrPXqgQq2teaovRah3ptpr+i8q
CbXC5LKwCRWTd9kLn9iS/nIhd9uitu5KkcmbwbrUj1lejiMxBFg1tumEuKP28RXTD8Z1TJ2klc2Z
vXQJD5EYJ1lAF0x2dHbuaz5h/8SOUg5lh5CPUXj7X5L6mGmw6cI6ptU8cSx94TG6v8EZE9K/rLYy
C0P1lVa5vdE12lG389r/DhiKJKhrHr3UTJvVzd836dLIGEH7VOm9CtllExBDLvSq+1Qm7zRiSlOq
VGtwG/BhasW3pTJKlGLjoiIB+IGhAIsGyQKK0JoUxqL1MsMomxMsnGLtuP1sYVPh5s3UgkDE4aVQ
6ea/NIMobdQMnxmq1YBHBNU3vXDw0ywdlP0qty/Rln8eFEua2Laa4I9IsmIXV+singAQKO7miyZL
LWf2Tkgvzeyc2WHiDU+2eNdahhcIjnWZ+SlIRrqQvmvTG2hK8Jsu9/QlZ2C2DE2/M3Blv/NQaUbB
cNLS2SRbM/6jRV88iu390D07Iop0csyIm8ZqQ8sdHil6VVq2pzIYlq6HslzSIUS18GfQvUG1FDkw
+enqP0FCUWJmBUdF7fNs+oy8z8isKROTJK2oE3UoUJgGef6QLhPfgajGalREftqIDzXv/wchb4fI
pLAt45u3hAiM/PblLqTXKwn4KpGZT+T47rlts9Uy4nRECH3CGa/q1trvNPYrRJgD0yGFImvndxrA
FgsLXwNH1Ckrwc4HC8BZfiQ8pvPfNKH/YyBwPCgTH6uB/VNyrted6gODlO+sMzEzzKgKLOaS3pIA
/jvgB+iRB5ksTJByX0zD2Ut8GDEZq08fZtdUxHp+tHfU9zIpzRzYsZ82pVyeB8/zoVxfhuVS/QZc
DCpxUeOGWK/3+3WZ48NqlmBFRVm+oFyNRLmkLFhV2I4VUnieELCMz3gBIxGDXJQ8LIGbb1DwnyLy
NAOmYE3Te/B1VUvQk2+SEfCvxOWqRGD+hLYRS/+wM6c2+RGyiZ+83jnOsH6P+XoIHyeuKEVKkbxx
NjVo8NYwiP3BrcuIr4eFOhbmKB9UbQHztHmpROadXW5PqAtAUyBZezikEQKConAwAlmhfauGupNX
MbcgPG23qpI9WQ7Uh2wp7ldXdQKlWj7GY9rGsELmeugXILu0sW6HYlIzsXrYjHhcRx3z4H2+QzQ5
YD7++ydHR7lY2sDYDUD6vcptTKSWxFngrZfUUB7chRGIO3mrHp6l9MKzyH/5dA/TBmhA2ys5ZzFG
7Ri40FgUmmm+zjqpdxZIkWywoX0WJxkk3uB3BLppbBu1ASJirp5nVxr2U6SxJGEz2yZLEs3gHV9c
7ffYyo0BAAPwZBTVMBKiiC7anEgGXr8/35l/VNtzt27HKGczvNVV+BK6fhJ/GZq4qKJ3OveaebVc
6hUFMoGn0ultIjiTpJuc8n0ORxFhM5FRTq9Pc9cFxbptjHZdfjEE61F4An0fRIJHreP1PbvJBthb
qUuGt6P7d9LEi/vMDvxVkosofsQBSUXlU2t1l/P9tVdGkVsZ+BR11+2xvBmNwBcNljYiIhmcmi7c
y94QQIXZgT3GHOU5HxuDNt5HvQwd6cllJ+iTmtuHh10K3w0xkz8AihyDn7HO4hjiFfz9BPOC62vk
mYZWRWxvb4GVpeUmv8io6Dw0X8WlE1xcb42eG+RBYLbOXMymM0WKmJmPeSKO1ay9kaTkrk3MdOwx
rJczDcEx4QauW/i7+13cv60I0klcuinYnBfZ/KZeH5HpAZivMpr6kDucXZ6mXBGJ1qMusqq7h30+
1A+HM72biYocJfinty0k31hXbgsyVVofxwEFhQbb/SDXaLWLXGtMeZ6kcFeUXOHODTYBwkyeXU8j
iTu+vbOW91bZSfNtfgIfg5xjUjRPfbifWu1Ne6+Cxyn1/C349GfdTl8arvbqr61lX0vugGREGbjt
5zVicAHqAludzcqWwM7xkB/EPhgUZ2Kmo9JMSNbTUNjne8mLSRxPu5PfuKRmvOI6MDFKcQYi4fW/
SgTPQGqUrUB2xh4xZogAbeYr5cPCYMQvam+8lz5HTbahdPBA38VD1oPGNqvQYYccwDcDtzRh3lDP
oAIf0KVlhDUThhSojhTDUJGxbe/jgqgQj1KkRPrGC7m0IiwU6ecE1mek3iOfx9DS4hj7E/RhHIQR
11LhIj1SF+TgqQNxHzWuokGW2Sp81+QWeYjhAjRts6AyDMmO0Y/+L/vhlkOSteZdPdyphCSeMwRM
2OtpcpGCz4qtdSdNAPHD6ZMjNEMWjSFrWFSBxFJBrHWBs2WXwO86Tu42HUmXqJ9gTF60yYLo8+Pi
98xz1WR8WBUyjMBToPN73rqtepIMqG3E7NgCsa8YvDA7tb6jtsCkjSloirmTn+aoxLm2QWBdJJoY
ygnsuQ64RM0jKf5TPPTuCTJ4KB33hshsHYjutQsJ5ymJ4OrXpDCDQQNcfEL1Wc+0i87lK6ywA5bw
WhgLX2348jhz0pwqXLj8bFai8APbbrwrItoATWrsVzWUED5i8L2iVie1cOF8fLZG/pLDrOY1htEp
HP8VtO3knDYoCswFqnq6cUphkFkGlwAkohdZOGAU/018F3sTm2YcjgKff1wBXkCphsgHMaJugLsx
swgNnDLAnlr+VEuozdtgCSCL93Fz+B1hcsv0/x6mBVDTEE1PEXu2RoSGsBX5dkiu3slB4il94sQ/
9e3F1B9rVgQ4fM22kE+YyYg84sohlwf26ne4dEP0gY9TigapiSZoLgYCP0vCvyIyN7zhnzPC6Hkn
+wHq4O6d2UgvkRyb/sKP9yFUZXXuKcOV8KnwtHsRQu1AUhIXlbYPhOxfe73VVgWI40i7x76oeVOK
EH+fgup/Wqy0+IHCAFgY6+tV28HY9tl+ArLAjgko4FdNGf7XXbIF2TyfCU3P8thtbeT5/QJOTTEt
PBrlNOxaEKT43yUyY9rCW9vA5BcTV3PKhnLLvl9NF02gdnuqP+iCPabM+U0I/ZXbxYeI7AOYuYWZ
nmYAbM9mvtS+9QtcGyeaAVoUs899wqeQsS5GE4LQB4X9YppZ2Rt8CXggkn4JjZejPw4ahYDsmSCM
kdATW8ag2MIJvhDbcCjGx0aaAM1B/cy8ej1s0MTH+yb+c0slolYzTTzPajgwQSKwxWGzowGz20wp
CbukANFW5c3zWVMHIUQrtJVASxNVpKHkew/UDL7VZLFJyqAJF75z7+49pnpc/b1MTA3XuROGX5MI
bhXcXvZYK0mCG08Mw7Z3W1BNS/culWTG1AhusKLw7YuNp1XhuMw+f4FobiMf8+1utjIV0s3TsWlf
clTbBVvAsthvWs7+98LosrCakJbeHsliEk3RGYj9vCEb4Sxhz8QWUjd0nKbCnR7NmcItROikYdBD
TPJD0t0xQhWwwZ02p9vOgza4PDvW5/nY7FSo/TOFOpnOFW3KI5AmhSwNYOKRhumH8673u0kUDeAK
0ipbd5Bh+fDHPFmldd2DmTiFiKvEHKTQ0/8I0zt4nlWQufbr0q8PGNugGOJXZUgVDmIyCYfHD9RJ
fYguk6e78UzrYo3k9XfbM0cYmklvcHHgBChzUhXFX0y0QXMgZcUEBwsfLtLdjJr7JOvRWQM4JDcU
1DVkksoxADkEJfAt2vPbSIigxHG9Ku3gldHEGd5RmYRHwhCRLMpmC70I2aMRhkGTXoQC4jN0CL1I
ol6zSWajb8YL5pj2g0IRaPFSI0AmzN/mtU+dQw51VBzo7Wgq087wNCDE0jYSm6Aa6v2JIUUhWklC
nMqqMm6temy2RcpOhvGPElgYt9vHuMw1k+Lib0glJTJJO7XlAdMIVK6riNj3F6NlclvnuNu7JQFI
FVEyG62WjU+R9AXmMpYA3Ta2QIok8gy/pvMxOhKBXucSV1ppBZMuDwVQdxvVnsboq9gpvYBlyPVa
DRjhpgSbv01K5tNrM8dxUpXEqFaVrxCQ3EioaB3kqOgbz9Y2mTb1a+Pbyrp6qBU6loWkF8Z1lwBs
E/yoLZ3TdPIaicDyhdJyVJzzN9vJn17ox3y6G7lC3MrsciivoQ7Mi3cBsQANYMq/Ox1mDHcABIN8
TkQ3+Cu6umVXJZ0qC6N7EhAiFpL+tmvVWlBHTwdYorF/vC9mLlMoKib1oavwWBWUl//edc3UCoet
gtGHMrZJQUBSii+FNjaqjcuaKPHKK05Ct0Rm/IsccU+RPGzAIKYNEQFYT2Mia8MGfDSv9s5hln19
2WLGju8NqRjUZOEDeMBUo7Z3kkQvrzscegiAs2v6CGp/MjZRo/+DtvhZQ3xcfoVELSSDFgB04BRz
78uZtL5ltRh/jxqZUmYVr2teiqLXH0arodkaMpa7R/C+4Qr8/3Seuw4lAzyTSY2tM0l730KbBrtO
+8Feulh8GROm8jpVMnqpc5DvCfGABbV8oGDuXtRf+YhJkmvJwKTZYf2ljmGnjdhuo9oNWiDkKIqq
wDuP6dlbuG+oYLtLx2BMp+pVjDAiN4ydLuL/71GgP/BN1w4BeiICx6n2Kix2Bux26cgtO2So3fM9
FpfRi5XAtyW+RwJ6VYFwa4AdFPng47EDtG/FmwQqfPtJHYF+dcjVPmsD6SZcdcBJcbZ37YrID/Qs
JPvyVehshBgoqUmeV/RmMe4uV6cOGwP3UjkLGJbfw1N2J3h3qV7sqYIY6nln97mcu7xi2zxN5eos
/tIbfPUTy1pob7OQfVsupNEIoMRol+CyCDp/veLLolgYDPdhck5o7Eu2Qzhm9tV0To+6e8VPUNF8
KfYjodDiZKo6rkn5Dl7rWWjQDqHsaUO3aJQcr82cNGLuwmc7dy040qEMT22DLWfi8ut29V/fYJ0f
tJShGlp5WdxDmSL1IDVQn1YtCZ2maU+irt8qHuOvRXqn+c+YeRMlwwI98GavCWvQceKO4SGA5wqX
B9TfjBDHNZlVpNGpl6sZ4Ys0WaBdINrTB1o5YucQa4u7gh6LwcHTcnAP3dXmA7prcmx32zubNhXt
yHyDzaGdYWTX2JEYhGDwCPED7iVbk9eDoQZc/3dHGNKH1l7SCMtVn/eDwJT1t60yodEYen4Y4JPi
4neZtbNffhUIr0rCxnAMSUzZHJUQFuVJvAfSYMKfE+iOvxvBOrMgtqdFmrjv3DbeqByWoCb0E1Kr
xZRF4iYnBUK02/Ofwo+Ibmk/Zm2oUdaHWsCfkqJO83gJHmo4CCwkF3qbm0Lh83Z8YSJ6MWksfbsN
Z63+zl5fVSWXAvGnU6uOxKVCE5wIoZ9iO4Xv9bfTlWBAo0kKiRtDieo/GupUdCZJbh/VHZB+kToS
b0gayQupUZVukYut+XEvSSDCrf2iJYuDvf7UHw1gHOqz+a47iNNNPUtICjPTP9DvvUvgDmGCO8Cf
XcOPTg8OoFGk0AezszCEfgwniUnYv3qU3SocswWlctJCpuY0zVLPYbfdrUsvmyugCchXQqk+SyWa
1Ei43yXiW3NKirEWmJuCPYxWjh4iRzfYhZy0Iz3TTLda6KPnQ+BDr+7qmdj3u7nGYrTvKL7B2r9K
QR4Tmox28CcxPBpBl2pdR2rfgPGZqn1yjpDN7BjLE2F0rCSPuwyy2VXsemAhTkHZpzS6YTGBOF0e
qmGAOUUwhRJ9vlJysN8HzOQOVoVkR30rfEyRfTJ5US3EkWO/WTMeYoDsraJUMAnwV7Bx6yd+n0/R
jOJ0WGO9Rom0Tdw/c4KkOVxQtOO/7siEvYNvzMzuPEZs3hNIeRK+pRgvi9mYpMT4R47MUnWH9t7Y
Bt5UPZ0k8kBqDhkSfM27UanaPfN7iO0EUfasYoESlgDG+7kz2VTg2gz0cRBPo28XJTSa3TUrg4Tn
dcTlzfMQ7D5SaIV8hzzuOr1HSn9vH67KFcH5XYk1EW0FWGccrD9ttyOF9ScNLcKJW3RJkbb8Sph4
xWVOPDUwvBSCwulYXGZARtXgYcJOPWCd1fPqTvcN2hHdSu5n/XiJsjQfwCjbqpPLWUQf6HQ4BfS9
zpg1Z5yc6mTqgGQYUP9jtnu/QM/Ypj57S2VcuRNN9rDpZYKC63C9KVWwTFYrUv/QPP1Wd9s3VvOJ
LWZHE4kk68m2zgQPZ6piTurKUKV8Pf3GGIi+1a2Xv0tkD/gx8h2IJbTDXWHAcgjCkzEQsqgC6mG8
MH+R7ZG8nJ/yY84oqJAyQb5FC3Mghnb8yrrhvpXMoSLUrlANp3mtl3VdZF336Uke9iX2NH3xJH+x
LCot39esnzb6hmlOwfyUgh7YWjjdBujQUzKZq2FvF+R1eNOJah5MQ8Gk/za2pdi9mW+4BOqJkV7M
XUmmNErM/UPmK3D14YAJPyEZA7ne90UhXEynSPD7LHFw+dYvtV3YoK+fHOurx8KrbMr8Iz4ibV0E
bAnygVhI3H7EVXBciUf6jUUy9A3kyHEarhWGXifMEW3QcvEpLicB+SiYGDvEiT828JhfoZgg2mCB
SZ5XVFfACcTranGdsaEELUUuL2pydw9/r3eJlGEMUrP9ncbsANeDX0zZNBKzfW4awY+HcwChNwTW
VYH2kPX/zQIIYpamkXvQmSD0D1Ljx710g+EVP8rPYV87ZjvSRHuwwA3cCI4jrEEW1hUt3wkfYepO
kzu8c6ibcfQYb8AV1ZJE+L1fAoKzn5ochboH6QOL1xmymZTW0TjwMzti6robyAFl5cDzsQv56wLr
5AcPBDxhV6K1/f6oImtWP4L5cAlGk/tAzcYOz7EtI1b+1CqK3/jYJ6a89W7tyOsEIN6ngU6ZxMUT
iyWkWzrETporle7hxiFwRgGO7WCDkQKhF8wLXBNU3G3DxfuMpRgcDubYIebvLlK5tQIvOQB4o5hB
eqob+furt0zXjxlbygzxnxs1aubngJy22BVySA36TwiCrhMGH04CActw6sHa8/ih7wX4TRzPjLoF
yUJ7mkqixDFWXEtJk7pwyYOT9Wbs3QiB/kcGbNLYARnKVx3eBnpRGgsEQeT1OL0mztsrkU5Ov5VN
N8CAkWXHwy5brvo+3f7HYZrZrZeylBmw+UnQ2pBTjSKGzWQPXvaysruUK2Fh01i5q6It42hiahGB
gytIda5XuXACcq97u+txGzgOHkzR8EvnmVeNzBt3DOGSZtXKJFllkkIoGFoVKgXS2/GOZrSmPF1B
GkQufHy806e08DAm6NM5tgF8Ej/w5HwpZZSd83pW+7C2Wwh4f8E32MZlGG93v7lKp69E/8yVQ8yA
xb73tEMMD63jxFP/qumIugdQ8yjk7EKXoiDI5yKGVS70LDhfgx4OkUlIeUT6hwjzLEU9WwYEqjWD
24WtrOZBQsb46Lc98/nBmCS0Whjr94kd9JhfePYv1UdQNoxFMD8Uj22CN5aJObGxFaj2rGAMp4zc
uTEzzCuEsgQa1AqVnBxXUo/O86Ypz2y6EZYQSUikMiUSu94FMHkQ3p/VRK/B9Zmrbe5sD2RWQRA5
UrBNZuEG4hd5p6GwxoToWemOimVYkZU8gjyZb8oImzW02/cz4YqD7x3hWEq8z90Cwd1XHrP38feu
2jYg/nIXCBDezZA/bh5p94oXGRkrIuhbviwMkB8tI55UWhszg1hRWjpTh2gueLikuUJtmlmy6nGm
DynQg1SmRxlVb6MGxBbbB0kWH/lWYyvgeqM29Gd2dhE1t9yNqRW7vvmA1rvqpQuwVji9hz4SZYog
oFdyhAvYuw3rZY7lK721SHMxNtkUaowpsBkfn7hAbozoq6758vpiJiI7h5iuZAgdTNQm1REsSFPE
Vkd4UTGN7lPkmRUyD3aUmfoLgaoHOz0NtLd0Sm/arpO5xKHytJICYOzA8Rh8V9zOx3q7DHGEg5AH
N2fEv2TJ68pv+/XxuUrJO+UVMdhk0lbSIy72Rj42RVzeQTO0ewOcPZqvxQGsB15a2/FZdqDuUZdM
aB5cofYXBvrTbh2b/Ei0WLSFsnAvej3S9d8cUd426IQbmLRb6tydoCDfiQrurt2qchc3dKT8BDgT
1W+dRy3c4KZtAgz61mGqKOAwk5mM+Xzt8gkTJeqagLYfYZYoqYlUf6o1wXP0s4IYk6WDqBxab8ut
jOObJFQ/j5HLa5DtoxTR+RrMpVKes1yVInZIF6xP80SixetxSgxEpqI8Aoh6TCN//wESDKSRLU0I
jEKyZnzIGkRSuPyvpXqLb+WS6Mj46+k3l2oaoy/9Z6HvPmrp2JFw4VXRuymM1L/6W8DQkwUJocm/
9155umrcBOGQwhsoT4efPsy5l6NIlibVXQXpWZWS2a1gqNKmdnNeBzldlmIWj0lOuPsovQpzn3jM
cpMV9kIuypTQnZyhXX25NsxxybntZGudG9ooogHlU3m6HIU2lWKyfrkU1zmK1lfNLnfVm/WsR/QI
SNNrGxay+dktWtwySoyV18uIbdUPGZ3LJxtC/UfBBI5hSY3KHL0W4+Stan/TTUJbkccwxQuGU+eV
NZ7Y/Z02XhZA4qA1vlLH3hnjUjhwQLyFXscWGjp2bE78qP3+ZUd7j6ZF1Wgk0apyQvC0VdxqzHRz
Yo1zsDs7x9lGqimO4X5kkOxHSv4eEaMNCEtvmGTeW+o8pmdPsUq6VwnodbpotCcI6IJu1S2SEeQv
oTSb0tnlC8oULotwGghoUwjK2NTMXTFER/V3u5/VIV4dwZuu9C2X5wlcneZWJIh0IOfvXnofuecS
fFXILOro15KzyB9B3sjt4KMPSL+jtyxzDvdVhmr4qJoMht2LeZxfCHnaFF0PIrxIpx6gIYexAwsk
MlHMhIWBwH098UFUd3bepZPIz2UH75kjsPGmILQreWGHchN/GJ5GE/dsgq4jaxOe+yBKMl/wNUdx
FGMHuov8u41M6ta0elchwL0JFCOf7+gZBiYCOSHHeRDkg+mEqwDu8RpEFd3jq2smMYDQMBKEu+Kk
xW+yvOm6ehDWmSITo/BXp94qzJzPTXca6GoHhrz0i+JmClxzxppNa2tKKWeNGEYawF3iX4iQp9he
KQJiJcDXSuDQDGUrtOOIlH/DP9vK27TH7Es2oFBIPBw8lMjP1VKEDXE4uwFLsUlE86SuV8enLslQ
p5zLET67I9YphIm3Lwg96RHsdzTD/17nIDmDqeif6YDCSUXPflEp9jHyySo1DwcnUhCpnqQySfWt
EsPyllfNdqPFzHmsVspDS1KVX1ohvMV3CO8+s9fNPBxNx9WHUaxeFn0jyjx15SvRF5sg9861IDNc
KOPJ73JodKu1fukMWIr9NxavgTA/YATGeID71h+gdevs4L70LMEYBThb211lR4SgsEoQHq2E0Vvf
5MOGDJFZEzhS32tQzLqzgIuQNWUrCl1acBnW4Ys3RZklTUUpNQYTE49J2nRZzjCadmXLwNQNKmUW
XczNGBMnnBED/Y7xWDaHcW1S2OdzqHCOWi6FxeYAIIfdRNJxs4neLRX5DZVPQqr9D6lY8r6sgzTD
nebBlkQnA6J/rtYPjZT/n4ZuiFVDcHYTFKAFGPzwPB16/lONFrCTE4bW1HlcmAuor8WtVUqX11Ib
78aEatiWctX0GHzECfiyDdlj9eWeRCk53EGiMoU8gZScAw19SRoXJuHYb3LzjAQJ8x5b2ZZ/8yuy
ni6XhrhJ1/wlCbf/cYKpgFmpRJ83J7ejpy7H6OsHOSJfilpseSwo1T9pXSalBb5XnCITfJPh1/jB
3Sg9qQ4uZiEF/37cBI6qV+8wa3g1Dxm6On1tkpVLF2NIcUYtFdlp/vdA8T68D44QffUywffyu8Ox
RCgsOKccYVfHY5xDRNMKBRhipezpS/bk7XehC9rOzqJAhtKp+n6QW5cX6eK1oP5rWhdP3nks2mBv
DqUtQk+h0gitmbycSQlhJCnKx5BCkSNUVkF8ZR0jsXLqaWD+CYBT6lHNkqR30BDw1t69cRTRO1Wm
mckLuNG6zgYvRtHarVQ18fivQpzOFgQG+R78Qzl95xMrCZlESINCIYXaAlW5tAM1hrW+Y2JMEcPg
o+y7+9NcmDK9UOx4JG3/QSI6CicjvEgyoullT+D4N7qvUChqpL8ozPcdCzonmy5U5jKPfuAXUpzG
lXuaaVARmT+tKHsk876u6IxRqpVWz/8QyQnau6qW7K+5FqyhV8x0qHedx3GW8pmvZjzz/c++OwdS
4T1w3niGMN90XEbEqQrHKDRp0ddbDVaWAvB5dCf40GA662pArzOYw0v431eGrmtvBc5sg4xWn5gj
8XvjVICMFlp0IUYHtmRVtrq9FmrRKXPjKhTxdm6hXjQjMVbnAuSOcn7oy/yIkbR31fOABNl6licB
uPB5fS6Ispa9Q7grz+ihNybJvWjzPG0/cS4wHFOZjbevzBrDBJgK5ZKisCICKFLr9BtEqSzwSiKb
YY3Toos035Lx+G9puFollpemLCgl7fklrxbHCA5vCm+FXvds4D5pLMmV7BcRcjynxy2u76lDvPGj
gVHFUXPN2hhSWUcxNs1X7bxR36+KT38ubDRZ6gW5mYJ0ZjHV/jdekbmUKcL1ze4a7OFUwdbtCvZt
s8fHYcMaNIbH5XiGXN7aQZqV53pgJfuvC4QqDwL16K1BZUK1UDk5KvlgNhfQGgkFDVCB/trYJzRy
kE0lTg6TLyi9REDlZRv6R6eM5tPNDfUrYmTC9XXdqcTMJNJU/IVpPP7YFrsO21MqdydSm9U6w7La
i/IfNzvFSfREnorTkEGiTDp7zwdZYIIKS7qBeqQNzM9rXGev4qyGVrFVG1IqqE+cWdVWHVeMftSX
IcJ0H6E19sNdUf8SbhAERKAqsfcvPpx5kGK8hWRYmwl90keAebh+XGKjAewMf3FmqlvSSY4pWPrf
w6hHhbgpEed1HOO5Kqm3l0aEdUuRmcF5tbHKEjbax26V1l4/fQdKx29Mpk2i/kOQEg73PZPubUoM
YZz9byWBscZ9KuapYQ67TPnSqDo/jAcUEzqInuMx4ui9z02fP9eFIWRu855dMXRq2OMFgWYSKtmM
tW9YP2K6yMRi2jUYOi8JFUNBbtZpEzWIFC0YtYJdp0yMeRuZfzt58hnjN1o2dQRVRZw59XPdrDwx
VyxDT3Qp4PZRpUBwGdEG+WEWke6rjFc6zDl7KFksvr0xZa9+Rnw5bNFQuxo/Mxjxmn7iEmSru6E1
e214ks1JsknPEPJvDIlDpn13w2PaPPeIA43srar9QF8o3iehPRPTaWeMmUvgKKPStWqU8wP4uw8L
09GE4A4/oa3L3/unnyrr8zATKLUJzV6o1OKYcufSbDAvHM9gW/mpgJdJnQGx0skUyIABoNWSerLs
of8pYrp7O++O5bx8BtfbjV/exgJdXFanDX2geXes64pTeNHF/RRWsOEzt53fddkcfJHk7zatOQ2g
N2FZxZp1E4TXP17tMW4/r5+tpLxTSJR9jVIATjB8EwcaTEKlfxvYi98HOQ6VCUmQWg511N5a3zKW
nxogLTn5wt7aEFfpqvMBybQGgftdejwFHeMajvcW6xOYXGRYmM8bkci2KCtHykKCYtc+j+moOzRJ
aWdeHZeXQ1nIbAfRYQw9G3DK0zCZHSeKX6r2TNijle/APJFvvxNnBM2t4pQ4xGfqX//zrnx05kgh
SOXk3RCS1pHNSHbeLhCyc0SrZSudt7TzWkA3AV6GWtiTijlyBKxXY/0lW3DKQ0PAxhn8U11S9kY0
D+NerFBYYmXi+EhKFd2zPXU2t6gunOD5xT2lOJi47uAcoLOQkiCS69knfyUrv4JhnMgUjeRa8MGR
TOWB2f3w+YLxpIS/SjW7x1T6k7bliZlVHjTzz1vU98Vd/LIDQH7qMGK0aFOmKCZ7AaSX7NTfjplm
Srb3LiZzhrGRGMcBGcQNCg8+nll0kKRjZ0CkLjxmnLmeUfBaHO+BTXi5F3JS51PVJ/l38cMRIy36
beLBpFytxrkGur4nJ/72OTzgL3WBhu1dVlk9g+Nk+omGxnG3V+42P+hcBsosfAoZhsPHn4QuBswL
pFZuA2w0y3WI8lVH/nvjHLkIe2TwXnrldkb8lj4EBi6RZQDhmnrcaMB94Y1l+dSPYyrIfHKuT14k
9af6a8P1UXwUZtLORj4uxQ+6LGhxBOIAjfL4w34s5VPCl5kzWauw5JVa3EXcUwzNmBXmNPwviw/c
JzCaPMZK1aTezNwYE5TxUJgDEmrg+QgA1eXjYX7bLgDsLmPhCOaIU6zihzfC/9yPOxpbHyATW5qq
qRowxBHOpWJ37Z6Jh0+HHgkar9FmOlAm4tArpmtZr3OfwXldqXHyPLIDzCHPvlEsxoFzz1HUczyW
mNYoJk4koeb6K3KfVcY2AdJG2X+G/5NOmaRbusMpLgh9eEhaCr8+HNQRa4lul3cN6qHPiO3EM0y/
1CblY1oyYP4EsAjRfXIYX6FMFXMHggI/sG5JkbfUgZ2qhy6i2rC/V56RPWUMQ+Hc9bac5rdzO2Sw
MV6ynu9eqvPvjJ3BQwaBowV2KQf+pWZuPDoBU80ztLvDN/fBIVywa2w4pOWpdGCbKSkc/4aLOBMz
8dShzawLVKN9jUMu2rTeAYJT9pee6h6EjOc0/5DEQzX5SvtwWuQjXkb2/LRjropDJjtn7Wu+arAT
0g9+MmoExGT+dJyI28CbcDk6nkyJBWXI4orwwu1Qp1oknovTtHiO4W+tQHHJdtTjy6u+euBOzaYo
fQNHNTj1M1/WYXjb4qxQhNExdzeqARKUuij6vaotQVp4QE3JravS9e3pJgauakmTp8+xTxqRvHNl
lRPaBQcLIIUGiTTZaPBVdn6p86GDpH/CsdK/l3EQYFekxMnAtW8Jh0B8t9cu0gXMyruZ58Yf0OVm
T9wQzBgxs+2G6D+mDmemG0yWgdlO+ASnZJEP/ddPeVNGEIQr340dm5gFR3ZpCKbi/LkG8l8bEgBQ
izyJiu2V5OIgR3oJgD0if/uJuVJDhTHxKnDHeyvhbDbk7oL5QIf/2s1bBHBgoPzxFkhQAsrX3yb7
E5zSyTueKKH/VVcnQgSIYzkjgbbR0n3eAPmNWT/akajbLV6q+7TV8ddmEjl94I2WzFFPRkdEnQNj
WM46gp13jBP9NK3tYMC7L8hoUycx44UiU8M5V5FfiBqR4ie7vPrjpNYTTdQrHiG3JA6cu4z+HP9r
P15SubtOrkTlDm3t+Gslx3713cj/+jPV2hhvfDYwcky1Po5XZza263Rkfpij9+NJbihQRKUiXMjj
kUF47rtjufjf/kUofds72Jlaq/E93NUiGqW6bGNdcK6iDc6+bxv8iaGV0b0cLwhlsmpGDpTDMMm2
nfrt65iqbGlZHj/vE2iX3ghWmah5E2kcc9WsVGkUZXDWMtd9ZIxDW69uFPJGNTBTxi3alJxvhF+m
PkrWQwypHiTJydGz2zYU6vNeqIeqZ4AYaLDYule29d3/00nH9NyzlviWVFhAdEEf1WiDRcCg6TYl
0Ox0B6ermswWUGNV98jxJlNXZnZ+z0rm+aD6Un+KFRkS7+z9F1k2825Q6nqQTXFcomFKXbbJpVrV
IeR48XdwKOykwWaZiIpPVTzu/L1tY6Dz9jjZid9HNbso8NYCIkiWYggyCSGjtqBS6jSXrR37XPAP
wh1I1YB51XWEAUFHCM++GASsNQJpLUwEy+bBO1xqS9VZqNGjDcVNDPyE/VNFuMNR7mvTyaYd/6Fy
xgoCc3S+dHg2bXLvn7R209dtHntj1dxTNv+DuOut43U/50Uaxi7scOOAMfWCCbvqdXcBlF4lKcs4
5D76Vj5BctK3WliuMxmCCDHQvfG06skjzBKcFpSt+CEGhTpq5VFu0l7iy53aK0IPmh/vQvxnsqt2
x99iMvqZ46YLNJBUP2kpQVgS4gIt8A4u9SVDGiW/FzQCDua01wMJ5Cey3DYmMAvbGqHOQ0lbBTon
qQMgLljZwmd1FX+qlYBcOvR4PRupdH9aGahziIN7sukD9u922mu9/+kuHuxV2DsIWk6eJorCsKci
svnpCm7f/LWakELAXoa0YIDm4UeTS+kX3IFM4Bu8OcH1VC9yq4lEK4wW2DtTNVpKD+h1hF8DGov5
99nWQyo+m+NvnWgRDINqP/saBJBl/+2fISvtTRVAiqzLSHXzhlUB/vUnc3XiSKf0ZT0Xvtvg1oDv
3SDcrgjgq/D52T05/ptk7pwutWBydJabUCzq/8Liv21MAqoU0LjpxDJOfmy6lsGSP9t0ap2viZv1
5/AVh2Pqm8IKAajuKecXhjE1F5i+wA/VwJgftkWf+VofCTWaIxpTKHGSVvm96LoVD6KTUtKCOgP9
y+FkbbV1Fpqi32GQu1Bs+6XyjqZQ9DZd9FRCtMBxEocTFqwjrr3SHQ+awXp2yGOU09D/Wn2Kfp7q
Q7DSE6bJAm0+C7MNedWFSNMJejYCPy3HOhl5JRSZ7klnQm1oOzV88MrNPT5rL+r+Zud8o9uFV+z8
0JT4xl7Fxe1UxxfjgUvFkVOINwMUkd1+q5A/t9TCR6lmKkKc8fJ+ZkXRCP0d6EBNjWpmhyHwSY2v
4MvDEEWdrYsxvuwtvet1C3kuRh+w+SQebJTwETo3JAkCMxsiwN6ADxWEe1HnEqIGz6mYKdgtazNy
ujxoqLH1XibEvP8cXMzjN/+GhokrqsRhfjz3VzzTkXio47gswigQtXs9DO3FJRDVsCn7SLoHNq6O
R6jXYh4rfQoCkUfsjWoUVSeBYbhny8WHXcq9fBmmamko81GQiTrzK3Y26PiYi2/3ry+PCYQWzHme
PXK3uOoroJHxg1RNj6ssU3Ntak/MW+7Wt51twN5R3vwyGCYyXWy7+p1pSf049K+TUt0lAEiwRCXS
pkeu0GEx081YdY4D49Nht+R0mkoSfsXEe1YmCvvBl38EUPq8sURYRFd1lLzUleoe2dFcmkH3I0s2
5oG5bIOAFg7Bs+98tdZbz6e4ZLkCXH3sGb7b6muZhweBFg5ognkQVT0awR4WUWWyKKoNAiYhCEcF
k1Ou1zkjFsKZrUA70ATVPmJXrCtxaZU6Slj/OIyrh8HZVTlEkeMkwJ4Wy7RR5mK30JxQtoXHubQV
Os0UuCMEdNf+NGRZrQ+XpPa5lzV5BvmihjnoUPoH/aWCWx7Fd7z2ExQ4lFoUSHdvqcXZOtUKRIs4
YwAxhQz8c+E/bugEhEgJzqja8r8FbmhucHlA1sxs2OXZy4FbozByP34q9wKvCrjh7w23+GkwyWUO
hGvsCMYdUJtg5pwHw6W/xeX13+LQrRJd2R0lmq2vHh3GboMKCYQaQN48/EK4RFnbw9x+V/Egf984
KCLUs4NcPHgfZn6RFvCPgnIfm9AtgLyt6Wgzygmuz3Pnh89RjUeqP16eQ5XFpaVNkN13vFMYXCyL
zDUp0aia7eJGQwvZVYlpPC3+08bY7F9wyqzpc5NG9nyQgVxqW+TawLG+mg9Z4glNiCuDpxoRSyYv
53/WbD8WbTrOUj2RQMa4TnbbCNvHGA+vnBCfbojo6MfoPR6UTsAjj8+AhY6T/LqIMeCf0UK6w/wt
2N43pk0g6Jhcf82ac0JEIsKBhov3kVsPnOApEBRvtkwS152NWyLHmI/5MczU6rnq0MKzuBdL6IOd
xSCEEmDdo2X3E149sUWkKJKp6GksQyhhieuiXNobZwSvdtG+LOeiEkwRSCxXYu1ReFOMxqzJC/0e
GObUAYuoL7VP1gg7QwGoaqyEFB7FuUPoo4J6YfNZNEYSEkvTsgdagBVQRyFV6a+KZR2s/3wmEDCy
z2KXFbtSryxZb+a3TVDG8L/TwnhAiNWZ1TCRwSDx6sdcwsSYlouruKvUcRkfKz6uWt5eFKmwCA9k
El4K8gUhNgr5WPxoZTx6BobUdng7qUurm83aAVD2YZ7lfEedQ0r1bhHs5JkEkFcbEytAbcNnf9vD
Thbk0EXlU3WR65rHxTTLXhcKbPJbX1qQS+HcqgEA5KGVmkXBC2i8NQFzklTe3skMp72686pASucv
uadKCBlDV1txzHHeQ0slWVnOZ96+scTOy8zrd5y/hiToRGuAakctJonQgFOFFr0LCQjh5OV1UiCj
almLCxSoMJgtfZ37HtdUTvI3YVHQ4qkMdtLvvN242XDTqDX6aON9VShYFOG8DE2e4qHgIzhTrQUY
9cOJvFm9/B9wzeSghNWKem+f80ARrd0GlbOBm0xvkB6Om6hoOS0du3WW5vtN/dVP9r5KWIvo7K5e
ZOSG1FQIR/i7rD/uoyX7Ho7bbYjQn5Iaj2hBhMSRTZYT8CX1ZJ7Oh+GxHQ1uofZU34L+nZSrthCL
MGchMP6Nj8FA9cPeByfDyfoc3SGe1266MLIahz5smN05hmm3JjV6GniiO5jg9Q9f5v/igKau+hDW
Pkeq9vSI1+T5J1H2hHY84h/H1wgqJ8p5keSsH8jmY0d8ajeIxGdqu/ojNUwru6F1KSLWxktJHulD
bXvnTiqfhyJI27fPaQ4dlWdqhoaHwen3aZrul1tAZFku1yuM+4/ty2q5idnlzSWaUvHYZHSxpSp9
RJclATRZyXfJD/X+eZpggeGOf23U9j06PrbB2tQBco1UfS7hjCAyB2GlOV47liqMIm7fMmxNB/e9
Zut18JV0O89Yh2NK5Uyjo1il2XKUwYcuiMVJiVhGk7pwj6nXUyZ63yOuXY9HMyY1PdkGU/0Rw4UM
SQH2ILdxO5WD7W63WcbmHnzBC7tbRuMauDfJwAjKJnBulBtIOa01Evou69do5urLttNZ9evRP1HY
J9+sfvg5PCjwBOdD4mFh839OMbsUvCtk5/loAk+qPkNiIJdZSMuTakof3rIdQFGqRQfxsXfa+Xrm
5ZZo/KneioJNWmA4CegeUraoV1i9wRcWqOiiD0f+6iTObrUfhbP8qOz2WehOZ7DT9P8Ur+gwiPSu
8CMWzc+6EX3340qo3nu0m6inUpBASGmtwiTlCMXkmSwYdjSrsoQQAW2ZegXOIIH0AEQ0Sp4nM7zR
L9kqp8WBrNt+DAaj+aHJnIEPyVCb2YqSaUyo1g/cJhsrdWmtofn3TP53S8NMZZIMb2sOaMkjaB6d
MVMewmDDLNwho2bR3NynRLFUhbub6P3l4288XUUvErGCCedTVGKi2uq1msoxjJxVGS58OPqSWD5r
vkeP4/A2T4Wz0xRLYaoIrPbm7oz/3V2/xT8u1nCsZkHFK5XGEqxnkQuNI86GoR/091yH/rfABjrC
SFjbERGCflWO8fJsrUD1HeonIHtoQPVSfSJ5MLaYTcfdgAjYCtZAh/RD8Wbm1n5AUa2sQcVkkwvB
W8A+3ZI3pdVFyiqVm4RS8rfOZAME1wfptdCRoRz22Yf/I31npFe6u4ZgP5ELRgQRlkmvRSVkXlWO
dGVdX7IPrB8Qp6Pjm0EIL0pgXHLfe17MXIs6AXCGQKn7H3P2YiPdDMy+LlhkFzlHFQs/bjO/OEIz
715j/sTaf1PW0Yf1YOFN0BTNTvZNGp3DbKcRA3i4zxaWXOY2WeptYB3krRZvOPvvtvupMQZQInPF
jYFk2B8HyfUOwMsl+3UYFJjIsiywasT2EGnidyCGIvIWkE12/Y8QFaPbK6kWKoPTNflvyRfZPXzD
4i2dCB4L2Rw4q6p40PgexZ0EpotiOgXDagmeoCAyjdjEvRvDLInqDC/d0Npmtl+cFlhlhlDTqY5K
QyVWIN7jIbLkuKqitDkiyTLgodV3JI2cuvfj0OueRDdGGtxU5r4ox3faDbFJKluQGBOS+zLIr8wz
dh/7zC7aYeKQFXhiMXh1tzNNSxi0B348dmtzYHqDP//SfzGqLTHQB+QoFCqncmBWQgPwCmUFSNLC
oG164OZ23Wj5CPjHPAT0ZyXZw8j5UZIoesUJ/5Q6cd+Xt2ZkrX72WLWCmN5FGs4+huJKnuW1RmZP
wx6PCD0CGY2eV1DWY9shiAJXuO8kvHoiETtK1NlBL+H9KHSAxvFacSKprSDGAVBANu8O86L9ICNh
rZu+Do7FaqcRz7Mrn7oAjGdN90WxmrknLc5SbVzL0/5sX6k/qhS4XMZFM0+6jU9+H0ww4W3XGBoB
3ll///xrfs4wsVDx7yQA3GfNtIWRgV0w8WEW16qym4zIsAnYXnqDte49iQS/dM5aO1kpvIebEKSF
Jm1VBK/JHOcOA4SE0Z4jGjM7y6DJFbx/8iLwIHa7tJNrGe87ueejXQ+lgjXUZTle7t800KpNmWss
/T7gVYs1AxZlSvtCgVgHVOhrO7PnioWZpP54JL5/N8Dm2K0iLj5vKlI+S5QJoPrtIRfKL8weQcYq
JlKYcMGxJwV0GNn1R/O5feZKO0//CDqgRqCaKQhx3swinWqpEuMNA7PKX+7By7ddQ2kCxmFtIfbG
ZFqTe7J1IfeFGHv9qjFNhnSS/Yow56Fv8BVXYlfv7LYuSqFIdX9WfLTIuvmhnblhHDHuwFI5EDvF
5WbgBAB6WVFkVOfmhfopnVNzCQFlPc/WCopqzoQXvtqo+183ElD6n9TZ/dac6mzX50VChVK5rw84
vxbIjOn8YhzMKW3EBoxoJ8KorsTDhhZ5+kSFCaqgDdocWqfGg0FLUtAA5DEfaucMlAayv2p/cst2
qGRhzHt15pANU1dZ4PvUlbACQh7Z0q2l360MYR92vRPHDfraCHGfvcgPWFiw6wZWIGR4gTYuD8Cz
VkGo1tRCVuCScQTWHDO+x7ibghYgQ17P3UGZPmHY6LRLSYmz96y9/AwrlhJyzyLgnyh6Geq/9loD
0xDAXWoQhc1A7vQZjL5srQH0hKDAVEgkHBdhwjrZuDPG9j52knWLoA9SKz+uvI1GpnQ6KpUX6N2d
z9l5EQn5aI3V3cMsfid0XrtoAc0z6uvBNg+PsHZ107PDOm5ybQLZkjQNQow/bsJX3lt0z/tSdJRs
lENWFzhc2TxfgOXbVsfIknvHKWHRbnIalbs2sJyUkFqPg/K1YKgkOw64G6ygxUMC/kAfFARYneWM
fausjk5gqCJsY6wv+M6/QLDPcLkiWala8U6o4zWWCJRBTXmZU93Jy0NXf4n9gBauo0kivm+oB86S
XkwmRcelQYQM8VWeH0PoZmSFjSWuzB+4auaJiwccpIgptupubE3Z4Pwj94SeoJozS6hy/teh+viA
EUtsFWvNKWzMYEjhKt/2ipsBlsncaXyD+O06Kr3OvsIl54B1K02SveAcd4OIV78ZkTY6IRCC1kDQ
g377YwRyq6L16etAuDTVcXnYZDk7hn5kDZLqRKMxhfhCaxLbc76XrbjFYEcPLA4MsrU1XD5iT4YO
vffB8MGVazhk2DCRAeoAY/Kq0Q/2iUVxC94c2Up6CX9rVq1TjMLag4utjnYq61dSpYKH3StZWh1W
xuOW92B32jXbEyGYPDu3OjxN/UrWnjfbRl1oR2lNy+nGpx/QaKWNSD6Mb8IzuvFnMpickmUIQk1w
UYikoPqZenAZ8LWqV80Ph5ki20HpvFLEiFRcSkRQxGz+MUNBmKQOmVlD6YA88WEi8EVwD1HFz5jW
9doDtCIdd4LQRhJTuJUG3Cy1eq1+ygfybKOLlHjgzgldFNG/mrmxVSzbayJfBmubhMu7Jahyh99u
68X6botb4xSd1xKnYs3UuQHVvXNi2qv2kQup1V4c0XKivkGE0VKV3rfB6znVJ1A5whdtPLaNnuHr
qCvlKDbC/E6vrcMe2PKmQ4TnZi4MGOheDp/zdWbpZnfx4St5OCKCy8ropREoUUKhrDI+G1O/SFZB
Aga+SyOs+Bh2V/AHJogh9EpfZhDNEwKfoTKeaY2/hm3yLDE0Fptv7IBQnfP1dtQDZ03Fdy6m/RFf
hVPELAnBweh9URdjpeF0BO+5Xw9hR9NKKEYwJrWtRn1ocdz7yzrLqdgD6qP/uT6o4U/tCMlIBLxK
8yKOwMxGKUOg8RAUpPQKXf5Wsc7T6bR+fTwy+9zB44OLOFPDcBFD+jJnvsUzfIQa/kjmWMObnYC9
J7+JX3zCnidf7F2ZdUom7675OgzupHr3cBslthPfqLIPc7DOhx4bIFRoTKTwPmD5EoyhEnZ0awoh
z1ZbHmwIpTc1eJb7/L5Djqaz6siffcOguVMehAD73baox3lTQYFr7SAochfvUwO6CKeGN1bjP0yb
rG4YuzReQL4f8vF6QPs1SRSQLDsuEZEO5Ljoh4BXitMd1RhbRACUdtzyF/L64unbu07AZjnfsu2y
9PCruk+2SidZHDHdacQtR/VDqZ0HIbmUaIjCTYM34sNQ1Nz3vQnDgswlKGUQXMCi5Nc8AfG+3pty
We+EuL8RSzsTN57k0hrgwCMLIik6VdZPiqJLM/19CmdNoUN5ci7XUjvpehOmLFG72EDL1lQXMfzz
o7JbMmx4DpOZd7ajatkANe2V9bKQ0Syy1S99pks5AaNt3yETew4aDmkl7bXKUJUvD3OPubb/LuCN
IT5jsZG1A2Uknwq11es4wa3b3IzlX44pouZ8eV3Ja2z5rrhD3vbcwm3iRFuXCKavplTP3S28CFCb
hncKd9Nwjs+iS7twENcxEXGkhpmD3VS9vQAaD8dbYLq7/kACURcQNY+K87KJ2jYdY9qAP72Pdi8U
TROABZx+TUsHo8dJ1tEJT1nQw+BXrAAtrmFFmcjA71V9z0Z/leRKtsFTYpBbWEmUSKuhhSGtbVK+
XqPQymfKhDPBqg8Ko2JkkPC7EHtOUq46Ryg8VuDIhTF1QbWaUD1UQjlRNOxwYcWAtnzZeDUDhOP5
Jn1olHoeokZiM7EyyefHEgFMZHEap+r+o/TqRycpJ5opNS+s9kK2GhbNdmCfkPhshwmhNqDLxoaA
bIdYuEFY1uk/G2HbFCcmRpLoqqjBsqSze/Dl6K4Qc9Agfp2acoZclF5K+emuAKVpj7fHeda1/J5M
JDuWuVLY/1Z3Us3v5zjIDhM2oK/YYjPiI84iC4VjSxH3QsMCWgP/SaCLYkcn949F8PppSOk1s+r1
u8oDGN8WgE7oOoFXEF53Iis8aKalzhcX6qdm3e1B8iUTFQ7BWla3yMB+m64ZsVW4imacsLqSi39K
w/FWDGFtn3zD2bOL5zssofANKQ3DZIDLIoWo0hvra6yD8zxyzTUtar5WsgbFrqeK3cIg6kbpvye6
1q6WnSSt522h38ccDqp6q93HKL4OPF25ODKmU57p5CsGd5JYmg2m3Z/02aV+sO4y2QjWYyQB5GIz
SVD0/TYLWTaWMjFxQ5OFEVZ851GXKlvukPPczCWiz9itDXhquA100sEHUg8wFlVDNfH1XLCVyrrg
4RkkpJkNJVmqHfxr2OCyIDto8qZPd/tmAK66VTQL158JjYlqdDPB1NW2INcY4+8RJm2LTouA0CVb
ZM0+tiYPCWnhCzUmdLIpjuaKTuEFjRrHqTkNhPVA7P4TgiGPYf6NA+ZAjyv84MPXjyop8raQMZra
o7eHNiU/hV3fEWyUgyM+dSLPbr8z1oFNWx/iL6yDEj0HGZ1OA/0oaP3qwdj5AKJx7cSR3rENSJsG
/I6LtWX8dbodkLpRDP2UCpofG7/z62nz9NOWf0E/xAs2nh0skzNCP5/ddh9XzT5K2VFhQs36wqVP
GZjZn8Xkq8f1wjPhxoDPPMrJ7siaenEnqzfHq080WQ9YqBw09TPL5WlwM4NObC2qWxRtRln2pA8U
Ls/2TUzu1+a2C9tamHFyxXztVoUSUW0/XlLUDSfcUGnW2BjNrp46mgTkQkJ+TwZrb6gUSqdKLamL
9NelWom5y+2kVvVAjqqa15aF2gW8bV3A54XZRrUGLtW2GxA85ItFp7ZEGm6f/SOI84gJIV4FcAol
Xd0LElew88RxHPC7B0v9bYUdhlGCvbl85aQ5mCInQUTgrZuwNS84W85CHQ+t6+Q+vEA/9Oc2VVZK
Y+R6cspD8kGAWjTLxNxj9oSHpoYPR+x8j24HN90fCpA9BBzTzUe8IR3PNDykbUnMHWM15CEGf7m+
IFat2yhyE9uX46JBwscOXdKmxS++c7uTUpkdzYpNRApqGDAQjPgk6uiTrBoy+wS+s3SI9Mcsf0pt
Rwo5fUwA40Gh8gKzRYDD6j2BKrgraf7KbpaLgMNivPrYZ/6KD3BDzJsVoggdiYipieJS8NwWkXUy
BuJoqJnFpvjfWN1nBdnqU57s6NTdViKG2IKM+u6/gdAZYvCJ6nmKoiVGd+S/SYTfS/UdAjiSOoQU
xEpBJUqkDLeHAHyfK0c+zbTRQIgkp9TSrmnZVSnuZeO4LraC/asbB7HzGhsLcLleHAGS8zUdxZHK
MJ4xId+9tkTmlvGRKhOUx6A8ZlAhkfF8eOvH1cMBmeUVh5Z3NOHNoXyNnKNZ3xXd4/PSrfE4+vHj
NIH2weadAlJDhgEXPYeF4LzL1H99lynu7XjBEJuzOK2gb9qqXyIOj1ZVhsTPDshDV1Ko0ODCQf0w
Bsb53NEV8Tn+AdazZWdsLxLWJSHEMRCeEjW91DwZROWf+bNNHFh+9W32L7bVcm4DXDPlqF2Be8QI
hfQQwVNjDltXKOdHjKSyuzNnPPC77XCK3VFGj7yjxVRve2YKMK1ECwvwD9sr0+4z0KljIzFJoFYO
SzVffzCNC1zF7fsNSxqzYjYMazgUS5+P5jfPXPxPRXPAuXd2NY8hyIJOYKlZOlv8aUng6CiE/rXD
njME1dCjwSe9VTwXxxofXzpoPEdVW+7hwQFOpRs2VXTCDe8/B/M0LMsZQ5rjXojV6Qe4VJz6pOul
7wIX/yHT7SlNPvAEYMdy3yyyTPaqf1ET0AUIs/rz/N5JLWqf8QMDJETeK6CGfhlxOMRiyqO3BT40
+JX31AepjhPM+kdu32ssFXXEzGJ3GAw93rGJTuj2dVK3pFsq2DC8JsfvahLYbAjf4cIy5dwsbT6/
0m7ezmC58oDG+iWGQ67PqYwfyFkwKV2zLM7Rn734w3K69m2KNNoH7TuQZ/0+4xGm1maL0rwNBo6k
kitTxPXMZ5724XhsmoINW90UYvTP42/hqIbLD8nWp6Wz6lL95LVx6cuLolLKbUz0fl5VlNl3ycCo
8ULWNOg9XBb5IHNn0oOLNQdOG6a2Twu1rRnquIgyZcCiH2tDeuhJBqiaZRSFbV9I+9VPnPsXBZJA
8R5YFAH8uZklhgY/sZE8tgZEnnGAFahVL2RMpVnNHE5eRpifKwZbAviOJq2vMdx49eJrC8HXU2tk
Exa0RNRDv8DMWDnmLDxWeeolpIw1FH454FjKvT7rMbiCQaec4sX4PbJG4sb7wI1EJRYZkC1vBonL
MPr817qRxlHCAKT0Ji6w1HizzQilnu47xQ7B5d2x0pXy0oC3TbMOXeOF919F2T+chpJdtSPcuHjS
Ar4B/QUGRWEXV5sKIScrLkkGwTcL2FsWSgGlYt6jreIpgbhFg9Czba43B0kyXgKbUtYf/iX+x/hy
HHRKwebkaglMCKygTnMuFdc/JXyiu/19WXiB/vuOIZQoteCKymtS2KS6x5twq8B4EjmHRVF8A3zF
eLQvUMJd9X2mypRwfCEusaVhf9tpa2JQF4G22D+U3kbnddoHzWvlwZ9Bc4TZsYRmwqBAtJoITBbz
bFamTRMQGw6EGtHvLIQPvaM09Z8yHVV11se/d4WMbky0MHep7VRSp1G0niWx4DdffqPK/oaDQlaA
tJoPr5hph2qcmspvzIPCfJvDZeZzGKe4RWia6AsmbdZpDhd6RQQzoUP6rHf2giYzenPFthwNFRsQ
T+Q+fpRB7o1a2bpt4k65Dy19w2mSxjHXIADprj+B7QpC+6vPmIOZ3Db8qFb3HyzaH4hS7x8HAqk3
21suQI0WOu13Sk07tqcQZXm/KLVOEhjjtxtTA+sRxhzHL/DC/OHm4DVqC5eCZvqWgbWEridxMuwk
3LaR+FjdIWCyPVyIIrQJb2wKb/fbZQGLncQLWTwbVbCNTyy+Bg2jMIkH1oQpjzh+VsiFalylr7JE
yPq9ZijoNYlmLmt0XHtEgSzVPpFMq2BZLRWyiZPDn6vPgeiseNiluqhMFti+s/CihG5g+UTi74p7
mE3NRkcHBQ4OLB8ChtiEY2y0AI8WQ8xCVyBT57ftDtAnQlzVVWBEaB/QHlKulMxrCeS4jD9RNXUM
PMo42/rxM4wDqN6S8prDPEtw6iqxkimk8cAOUOuXm9iDB6OP54373nqW1tppHzurJNCK8Sq4Jh0F
BubORIEAwJ/MLFhdhf0PHXTE3ldE2XJE0CmjtkbeGR5PjU79Db0kOGcZSoTDeIQE0Vkc+tN8nf6w
E1papO/S1U+shYq+Zj2BlxaG34w0PsYOrVnMtL1V5muecNX60T2L0/Vwwt1ZaRFtCUz4EfuQF2TJ
tPDVPDY8RXrj4PFfITJ7k7Vogc5cSNwn6ccPELX3mkEz3LyI6NXchfC7Rt9Vn8rdPfbo5RsinGxE
zBr63LCwENvNQPSolN5dzyOlJX5k+1+2+CHPsu0AijcsW9JNxXtvWGpyts8ITrixWqxaLG43Fp+K
ljuu9HaaQxMW3BIATtlqWx+39U+9xS2Ssca6Mrnn3QjRd5orcrDMfvUHivkPCbPhXeSYACcvlWID
gpr5h2fzGWfe7ZqJ+GLSyTFgl+bJjeqqzjrk5+z4qC5C4M3nNE+xRVg+/47wiKXilhR9+f/do7O+
zgl1HPdwmz5vrsKTUQmBaLZEhkupkdsigMACyqyroeUaqSVdL4yRmXHYhImrHhbUzJoOHm8eYIVK
gVnHM12byRsREP+p8NK3fxvNdmxI1hulIjUsidqHtmIMVdBev3kcQ4RVyjk6gozwplL8UHCpdfHS
H5xbP/V9Tg426agaiWOa2xmjmQ9iMsbYygzJOOBQ4zsuzegix34CwKWuSe1Z9RCGadWFHzfHq9Pg
hhJ5iZ0UT7z6oYOXJixuiRUzzQNJlE4bAeVmvDYYtRMxg/iw9hzt6LCHLkmwOMEyVnkxSLDKIV2j
ViQHE7/VA2kMh3BHnNOSlqn9pE+8v1/sGdDODlMD2T7M/DESM3cdKL2Lhd2LF1GGOIkw/ubkG5vN
tuE0xNe2XQYfq8IaE4l3hi1ZqXdL887qrd1Yi0UPRzHQqS4iTI4+mqiaBi/8i/5aikU9tWJQWzAb
MntTIU17mKifLWYXSoZRhIiq0tYn9K9cplMdicBPwmKy3LlFjium8XZGxlzVQimTGu+YlE2yIJe5
gsp+5TNjszDvUbz+yUFx8R3Tpacq1r3Thks/LsoayRqEVjP3rb28J/EVz3dl4658ibEKmcaefMvw
ZMFGQj9pSaQGoONCVe7hceycBg2/a2z4H3iKVQH3Nzh0XKk1n0LRZUjjXdu2xElavTAk622x8pvu
w3iJlE+/SIOcM1p2yh9BcXPfP+Wq9aZGe5foGq19jrUxI7gMqERA6AordxPZneOT24SBezRA/xnz
GFMClUI9CHAn3DsMfc1thNmiYD2l6Iqf+p8U9r8gS0/NU3bQwVKEczMxUZ2mDCROjaorDVBS28HN
w3figlL4cnFP3M8ZeraFMDck/UILotTMqLyOdEXlUwIHVnqI61hIyt8gnr/ceO0YIyZy5Wd57Z8K
leWKXwkoQwxG0NMvpfgQvTkDq1pYOtfY9ZlqyTraUQ6stkzkpUlNxI7IhLxQGNoaZ9Mac8IPuMPC
SbjOIyjLuVsSjwh5KN7GXqqbWffMsbRRwliFkXNO7tImtSF/0avMUKhAYLrdr55/HzlY+VRKjKrx
tMHkvVi3HBBZKgZX/FGOQmRwdNg4tRIVpSvwpgmToRTp5Qfn5jEM8oq11y1aV3oY5ZGo0shx98+4
7JFL7DxFYsRoys2mN2Hirk/5p5oiQk9sClRvPSl/VC88l8HNXraNdj0uMhWSaYaSKu6hOhliYXeN
loo1I+htDiDJcV4XwRCkzU/WQ7bkFRFrFnmH+JQU0BrtWzGBNFdt2XNQep+2pMyW4U07+uKmGMSh
Ct9q2EU3s3g6XeGqbV0V/ysIORebGqYZGrr3Mz6QapMA2HK/Vx/1AQ7ZJJdffQKwlMD+L9mLoDMy
VimfoH8BmlEcpnw7qc8qVoAA3jH09EothEqDBfVaJ4WWMNwqeMrTU7AqnlRBLsOb7HxobyYCElnG
tnEmiBmk48gdvYx5UjjOMIURhriLPSVLzPuzKMH44jzrej9O39b7TZJpL659+EuciTU5AY+TCwG0
+YIWTArVXF8xa07fLsH9sk5vNBKVeEfr4pIow6B4cm89yxh+d1Rtmlicjefpm5T2nH+g0Cfc3Erz
FOJOhrLnX3Bp119RRCclewcJpu9buBcD3s443t+QZZzlQwQYRpLAY+gsrDc0iXpRqJhGlbvBZGa3
XhDvthsIM7mAFO4/PtuxmuktKjxg6iEyAw2R/nXOvJr12kJF9m+DPw55OK41K0b2zsri0MjP2qQM
hPoNCLdmS4f0rClf3lGQ90lnFYRsj/bqra4trjurd0LG78E01ebMeKExNkyl8AcaPlsIboA+E7OS
iLihgPfgXUj0SePF/uh5mncaGmK3hJrE07mbwBLXishOp4u1Ufpq2HwpG0smq1lH1SlEM053mI0K
Fqg0nHoXTftS8tuzP8nFCriAbTXaz8ADfj1g77WxvSvrw9tvm326jCqPXHXYgUCbDgU8WFuEtTlA
w0eqZIte6Lz3f0S7HYt/sYJ6xEr5OFHPyKCg3/t1FCvdgqnGOIQiLIP5IsWBikr0W5U0M5f8r0Oj
6jjGlZQqpp+r1nGP8eJUsP1U0zzXS1LjaAXYZUaR3+EvbJhycNgxH3omszdB4SdnKeyVAJkMVl6u
/4AUZFI+FHMKmOEf9liCVRsIZg3pFlm2yK0sVVEtZX2EKvrKEhbJ8a8ZhY0ueQZnCpzK6H/++OAO
y4pewpLLvZIY5KhIl6XuFoVJoqqQtZwiRqX+TZ2MY6vXa9DR13KShPUce+HA0VDOWDOu8tfYeaUF
XgzQdmiK5lFQvQKcsvX/sP5X7god8uXXvIF3PSXd706O+GWrvlDBCCgyobI0W/pCuBnz3JJA92ZU
YLRbdrdgCXVnMk21CrbDYSpcglHJyHIWfTLh3r2p1D7c9yZMXcfwbdDrBnBA49z2gbS/7vs7TIKU
nA/JLpwcfmsd4MKJkhywF9xvNBULgksDyCigzZVRF3n2Ex3MRO0wpuSC1BNlShnUSOMDdkOFAlw4
Mw41Il8zarM3rf+SQh28hou6M2oD8/SwLFcEqx4rDNdeyUHNL1L/H5iASAaM+5SnH6F11IMpyzJQ
e3hxkh94YHG+hVVUmNO89GolnPul6YjxHTjbJ6rxuUL4GuF1bsxhNlbSN2s1hodHBqPj6yZ+jjKN
801TmLsX96HKo98SuTimmxvg/LOqkm0ksqsYkYY4kcyjaGlyJsEWDnoSoZKiT4HClCzAopqa20ad
nxJaKCnMv0oqpNhMH/JJno1cvcl+2qKak1OjIyYaphYeaJjlVkWOW+bckHzImCJhgZ4f9qRfYgqI
YT16Ti398fknDPvW5VE9pYtEajUT5z4zw4QbiG6Y+GP3wGqVObDUv3VDfXE5VFfhD6dcKzsaHmpG
UMPb/UDV2zKA7nCy0xEyYstGbFUIv9HOg3+Fim+thDMf57UHG7S9hZGuzUuf1HBfzMJE8ZjPhaSO
7eTCml/VgNTbymLrnSWmw/lgRrMCK/50PFs8vQZeqYCh9v7EfkZjj8qIYprg1LzL3G6ipHJ62+W9
KWdJdMhVOQ2gNn0flu40wo7+YCRLFojZR+nFYGo1Zy9LwkJxNqdofdgR/tFXE2El0CbEeQzRlYFc
YFYxTfa4StbpB6IFtYATZM961hM60S415S8Glj+BHNQ4QMahXUcsy6TOsvHViYjQux3wopEiI70D
6jN7TPX4/xgoq3SNXa/+vUtYXq+gCETo0YB4OWtgKMIuJmxQ3XU+DzO2JDCvdN7gLMFlN89/Vq97
7iIt9vuhjNBZUTUUlyz3IpaPZdV8IZHNDkKfytOBOnuVelKtf3IPHQrQeFSeV/tNGaLDyET6kVU5
BF5AdryP0/sWiHO5W+bGJYDpqeiOMwK3EiI1C2UExMnyAg/WKuYfzWLmbdD3h+mh7jpqCtTc3Bat
SAArTr8SU9VVlafR3L8ywZ/wfE6HVCsa6ClMExb+YlV6ST28EJs1lWqF2s/QU5ZZFCdN4ywtEb0d
ByXHyY12yJXsmr/t9E6aeOTl9QHuqRDjAa6azU3lOn3mZ66wUrmulBbgUrf7MK8O/tcXw0E2ET/u
GYq9KvZs+HMO0gBOLJ7y0OiM6JkSgX90oxDfg2j4BXj+RC7IO9LqrOspC0Pp1649rbaD8Ro4Bpy/
VY2AdpvY1sw8+t9ytfpnjSULohSm6O2nPkj+hFWXiIjALqVNzOd+SF7M9vcnZPoZFTvPo/PKcIBd
j/0/JhsFV0PPJ1EhH49eh6vVma1G/BclE/OqGdkzq9q3QFvuA34H4hZTXmegtfBkpDx4oYTKxlHk
QexH3nfpk4qRK61s2G2DU6Knguzy9VwGnCRf3z+nmRea7N1W5A+N55sD2JbFAd3hiTP5L3NVy5M0
mGCfUZBL4924SKPj2abMMdH5CVHsNwWfOkf6B17Z9OHeOeZXVnwbN41lgeOzpMIMBXSlhI/y5FOW
1JClePQrfCHzQ4vKpyN7r9FSFsoNwIMBxJFKBW1X5AYp/ciS/74WQz+jECIjqV+5DCIIYoGoMTPe
uPXi1SYoKQENQKyWvl1FbNd33K83jbK8PczkDzDR1kEJ6BB/wNHx/xD/PD0z7zDMQZoGi208sriT
VDYmVHAc6W/VXKQ40ZgsGTBt8AUVEy6wJB7jeR2KGN7Vps79DMcgLFOoZBawYw5vtPqq5qvoap2J
ui0rXi2BPLUN/hsNT6oHXPgFJU5aLzgWKkkXRdfG+mKZM44LXWyUGdhQbfDUtw4dIoxwXTtCErYk
SiYjjKACHSLm4IkBap4QaLbs4y6sWdGpuEV8Zin9HjG3887KjVYuTFTt3gy5AxU74pfpvhRPkxMV
/gutAGrXcKoA9j5bTGMQtF4LyJs00gfmQZSHh61PaX1jPWl7UcC5Ri8znC6xJbazqr5m9hLP6N/k
6Malx60Skbimzpj+iYaq6OBYDoihFOJ/bv9IGw5h4AXISUd5gZzwFsEBT/ObN2746N+hO6Pw00U2
9RjmH81BDt1+stcr9q8e6s+oO571DONJF7obU8Imy7ep1Ml/NcbR0A0mx3qz9VYrAXfS2RbyWKsZ
Emn4tEe8qqxWALL/t6JTtSQsysRZeR3qmimbqByTLeJM5zWqYLCW8vG13/gVTZBL2bXkJdbaHcN/
vP1bJniDFnp2Cd0/AKI5KqXULQuYWnL3h83jQiFd5OjafzcN+acTEn97Qi22OUa4cs0xXTd9xgnE
UeHLwAn7CT0WkmV3djfm2D5F5kEAi5ozlYU/MPvN1PPHVQ07ypyAdhWAk4ejBDeWW3VDG3gRpx5R
4TlIU0B6RJ8xn0FBqpX1YLMPNSbTU5XRnY3XmleIVBMuKSmbuVpIPGlSz849cSrelVW+mFMsCRAJ
91iutlCzNbrgD06BVErigAk8JZXKz4LO6TSEaGiHLfh8qnwtqlmIzpwqsCVzAACZMerlzreIAt4x
MIl1RTgRjBomnSmLnXcTOkajsmXVx6GGjRlx6RjAj5KQwE+ElwAapLzS7rG876OjuQAndAemuoU6
0oQlg/DMipH5hOz8wNVMhX3bDkjtC0WuajL0vokiJ8xX6Ko8LQJlZdwq9fYWoSd7uhN06sgK1Oby
QUucrpQFRkn4ttZzDQtKwQhu1JmPojgVyu4ONNvbXij8m+ikUHZvwaHA3rH8THv5cNCkiMV5HtIQ
E/P+XHq+rAS+LEapHle/NTEXt9sC1W1wk7gclO6VLBhzG5AzP2KY3VyQpIUQexMI7YXUQmtXOsOq
8yDQMyJWx85LtKX+HSiE0OpS03fa7qAxTB6QsLA8PnZPaNq3MiHuSa+jAz53kyZ/Fyx4PIHVb+vV
7RWwXKca5LR73yv7fbT5e2HuZLXE73gcHYSSab+Zf86gXOk50Jim+V4oBiVlC6DP87ZEzj53vuhz
zp5gNNvVTePgEmxD9Wys55hRXD6ebbPh3eu2I6heZG1iO0mNQZjk5N/QqLStAQC9+++tJjYSgMW3
D1VHX622qAqlZQef+7gvzinIM+Ma4a4ll4p8vC78bSFRuZt6+kErevMtqidkYWjjx64tBe7I0yfW
OP3SJOzHdPVgMUJXw7CC/eOaetQB9RDGkfVWkAIFSswc32baNW9ot6/MXi0WL5RntkPpJgCj/4P+
XSL+MrpXFlxgIy/r7wvSmzarA6AoXsH9T6t8oym2gn+1z8yW4bpRzS4eAcXlgRlpR7Pyh0K2Hx1n
XVek9BYREBGRj8apCVKcJOoTDrfCOcMiZbZ/Nawlujv8JK989RuAHI7qENjllOGStjmxOyaBskCL
FDfAwcXNpRhbvmtULNQeTistqqBypU4UA3I/d17OaS82BEj0brQOufG9r8uLAInhfm7m36a3SaOD
IImDUwf8MzrbxjCv9broKDk8fbvjbUJfAFydUe9wMn6+BL22IjlOg+yH3Pxz0SLYtKH9+QQpYhxv
aenpdmKCCwRrlIodzM+RXNn1/8eCJ6YXIX0qTSz6x5itrAzeJDQuSlGZGuM1AtRqSYLmmELSCw0d
8/G+pIsIUav/zWRcQiT3jygfgLsZELwMiH+Y2w6GlLj5brgpB/fnPwmHn+puDwXDZyjZ0JpHz5VQ
LljIozNwfmneVNheCdwAeAp1eL63W9S36qELPrM0v0gMs5Ad8VfxbVPbRLbwPs7tTiOt1LJz0Y4B
YTsEYzHfqzcEf3Hxh5wMBWEimrzNLrX1FrvmB4KJTAePJA2ZBVFvw9d/hVsNuHxEzSEg0hSccvt7
X8THH/Y7n6hgE5/dh0+4kvVtQrH5yzHnxocGFAUi/Y8VqL+7xHv46DDOnouRmAEsS/+KzY/N0o1I
nvbmE9bnWPZQrCRAdFuPemA98ThrdtfjF3xzU0wCv8rqlyWFdlzU48+tTya/JpBRXqAhdhfKnn8j
gIR1CqtInLDQ8XG6PkHW4+jNC9nrlvek4f5jvUUBRWIfEdpdHncOFBAc1YVGQY3kDiBxAQAJe5hm
fDeU3OxEUs7MTdMFxLrltZL73CTS+EbXO674D7PLjqIpRbB927gj53UuNkUolp8cC2CDRA1qBlvl
nlD5n2Uhqzcdp7171TSmonNa0sVVfx8P4mMCxctYrbkVrGbjWg1qqT8XIhDdFOmaTXMpZaF7eL9I
UVZVFJ5snsPSY7NspOFZo6Dh/EJNwUeTA0Fm+/LEzd1Yh4CDYuOFHo0M8OxQYsLXsf0NHSeiLalm
r6f0trRQIKA8REXitO2KNfY8HEE5NPUpmUXzRLdxaeV3rDIuML+sp36z0Zx0bPD57+s8mHyqTxtT
uIjtL5tZ+4DhsgW1CrIUWDrIADwG0Zvor+QYNp3q5JrI4xPufCd1Ec8WgicoZE5t1bjVco/JNMOi
1bg4xICizZyAfP4a6VhoKufUVNsbB4vIjEW7hQ1QWbiQCs1fOX5c3lxWnCYMFh4NKkne42vzpWKF
JqZBfwnUfr4jIcSpZsTqDk6bhI3fYAEiJTOjetMh2Rxn5XnDNqNbeIKgdsBP4IwSbXWRMwYTBBRa
iMfT0NlCYMPoMRfD2vXbxEGundwJR52cF8XKVOIvhDgwx45K53jt9Wy4H9EOALIYmLnjdXi8Cwdd
wvgfxa8xUVBfP61BBzBsGV6RsCmXpUU+yu8+EvioxmKpP9TBZnRy6CmAlnngKYRyNpqddtu0E4xO
A1IAUKR1+Jp8K7DZRStYN7bZMaRDx3OqMx9lrkRvQ7ntbkXWGrpjaI9jOvXgqcZ33mvideqIWei6
xVzdx2PUcFBZv4s/ueQbBebSKAqoLQcXsnFSqyig0LDFvw0BapD/dqH4eJrBoP5d9DNJdkxtPP1Q
Zgfkp95S9paPtUF5hkUKZTtU5AMdlMh9cLut8lN4Y7Du3bNaaHEipz8pB3Lx9FvVFuuKeIWCTmmb
13zP1oOaHzUc15xM4XUu/jGX3ieJ2EKV4LFh9kebeBbtv/TgakDXxdmtMtE8GByLS10kVRtdj1qb
WQMJSuKIZx5TUNguNDkAOAFrGwRw+HrHPgwSqNJrExYo9KKw1R4Rw6iK6RCnzxfzgLDzvlZ+zHU6
uv4lC6R49hR3U1To25IUugP2zt6jwO8qx1jrhvRiVz9ASMMg6yl20hSm0Y8a3M6KVCaZ1hO2GQYM
wb9gm7ByV2ENSn2IHbexkRIk6NAkkBhFyxWOf5TwG3VDD0y6wGmG1F94lH9cvP2zRobgNMQdQcE7
ZJtXJJbjbJEnhFXDkzYBkeliMChQvYpqK5LYix/LWMDtJo8qlxPMBlAbu3E+FX8QCmeSy7CVDoAJ
1iPADL+CbdSi5qX+A+BtJL0XVWTGTKtB3+8/LJFl4E3VJTuilJko9c1LaMan++JyzRIM3kUTD2oV
V+Bm2fp9U15e1lGAJBx99LlCtfoemIxAi/UwQg7+7FNwe+5N1foyeJ6jFYL1/bnksgri2c5VJDbM
mjHfIypn4Jy+OmWZTEW0tj4rn7F8lz2cZ7iXKKzGVp/WeueruyX7r2fXvwlsD7j72AzdoBjoJwIj
Y/zj/4VvovUvImyU504UO2QoPzO3Q5LLceCP1DWTyX1hFWMh9nNqhabtn/2Kye8f+7cjbojVQG86
8G+1aMMiY0/5Q9iQupqhAQkV72/Y/vi+/Bo+RFucwUcFICsOv/iNmVeVfnAw5SWkuUaZJGJxVFgJ
Pyp6yRMiJ6Du6COptmYN23iokGt0ZklqkQyoyKdHZn/X4RFBoLj9u6zkRtIZyjiG1QtT4rBsM5Fj
LZEmlPjqI4wTYKVRkFgc23hvW5Tx2JQmogkwtoG6axML04IjKBRBw/joYu/Wx4FAHQL8DPBBG71A
5CVc5ciUuTqZiFw9Y57rWqveqk2Fm9LksC57mPVhPL9moZIxEsWHeDIx2txzPoSMd82xJ1BK1pAq
vkr6QrP9Kc80GQElJp09xzVwjWRKP5hAmBqsntqNtMaz0Smqwh0AHfnObkB0AOB2GwbjEypbquLX
tIM/Yf3V+d1EFv25n9D4pOe6SuoZBP6cZQAi1J3nRsklAnB1Q6IoNVQlOF7HHomgxhhV+zSeIPw+
FX2sNratXj5VkN4wxei4vX3OePYPLE4gfV6bS1bJdzDHLBQlXpt3jHLyPVq5tUS+7S4AjfjbC0Vh
RtJmKuVdurXCEVdCZLFSsgTfDT/Ghj7v2aLg3RM6lSW4oCzLHLYWLcVv5SuyC0DcMB6n1xtjF2AD
ll0jn3TAXNk8E2IrXm+LdQGOXLJDP2BnSI6l5ScEg7vyQPBDJo235lPA9cjB4WQVwX950brrzKwi
cBgLHraAc6DGQGbObY2b287CH/7LswMbF0I8MdRxtkgEIiElt3AFHkSfQk/KD6od+twzdWL3VW2T
MbqklKZhF6vKuN4eUFgI1ZWSatY//0tf5plVrcNiYxDL4VV5RVA17CoqtB1BqQZ9x6PrNYUEOmfb
OE8goZab/grkGJLkM07QL5fV+sclfCjsyJRoCSThZrNywmAbHRfVwLJsdNBG6tYyV4a7VWrVdjQo
1z/6XNGdFx/eaiBlMFsDjaDExmUbIHB+NSqr1kcqp8ev7xUmtcHKzUyrZ6FTfLkuqfnSyr6vjPGc
tigMtoLqNvjpGGIKpzDRkGe22qWy+QgBBkvr9hArceNDtn4XsAZN1ZX+RW+ux4BC3k2rQAA8oelX
2Xp16V5eAG2xrdJuyNZujEP5YtPz6VSBy4fP7MgN9HqsBHOiJL1GOrUWH9Hy/NWj/5x+wXpE+F0D
ZG4gH6qB97/cRaK6/TrsBeFE0+AVB5XW7elH4XadGrQH/2bfZCnB1gqUtn/a4IITk93hjZBsCK5Y
RGjcjlheG3dHXyWFmVD9PkXQFzn3KfSy4AYLa/SBy9eEcIderCx3lU9IQXNNsjqOXGH4Wlg9DACC
Dq5ITmexPZs7CkK+Z7z9WI7NULcP6eDyNKAdkZBfQJnuRO9Uw90VWzsLOkgMcEH3tVffWepFQ3fv
o9jLbPYQn3Z0Qq4v5eS/rVgyVvrZ7DhPMwp3qFGRqpr3nWjK2UM/OoTPQQoxDoS7ezgbhsZBrqJL
WH5XvW/38XVGtLwTp7dJ+kFjy+Q63Zho00bpFs6592dkpccHgKXhA5fZarWMs15ZV65gckijTjQj
lTOIIfH+T4fGduMlSE0AeJxEjrUdRPlCpEyTXIpaVy6uzgIoBoLa39WFndXNJMQ1mviuhOdExvNb
c3wLVaLJ7rTpiMxaE3B6YQlpn4LWdkf2Mi05/h7tT4sxnNRKJw/BTBBzptWMgD7mYz4ed2LiqKPU
gjN4wr1BJkhCTakhQ/msVMEsLqLGb8s+2FjwFL8/94wSoQjA7r9dMsqqmwnkSN+MS9dZAbzq2VKY
/cmkV47B3DK9XWoHY8CNwm4ThrfRUhUa3hPpfo6mgFoHlLi9V5PRYhLIiKbmGeMds3Lv1hRysgQH
wo0EN/a2qK1hOoT18xyo+TmXovEUaKQtvbvRYmLQSI1CHPwXm9fEfDdBijtGEJY9g+/zxz7x//l6
WA1eY9YUSxFn2cTnAVSIUgXp/gpn7fsNtZL8NT4J3BgoXnaNlNlvL0FoAE7JqUYLgDgILISib9PB
ZTPvK2ZfuivhH5ilhO3CVZsWeD13Maz9MwItySd1xRWurhqhtYVKGU1bXLynMdCPWzzt5s3hUo9d
yrbUC0x3JFjoM+Kaft+pmsj2kPUQi99dGrFXDLeypHPM6D8a0MM+OmOzcHvALSITHQf0BIPTOxal
IoNKW1Wh3reluWrKsZ/peKsV+Iy1OaeGdgsMripdQdagGR5i9OXk8QcLWVZCIFVMjnAsgA1JDHtU
ixz7S+qVZrc+sqeIWmwvTMGpxzQt+oFh/yGa68+O3sxrcqbzfyza760332lY9iWimMrng1j5ZbvN
pnVwlQLIyL+15cCNAuUm7F2zxRSx5J9JtAvvnV3DREggMNPo+jopWqbsRVtwhiQaR7/TUfRFesrO
P4baepBF7Z2fzRGAKmUJn0t4cBxnUIBBhqfRSpCC5W8Gozxu29Rv5GZ3K0cHJ2X4VoED0D1f9Phk
lfVm0ujy8oqIh9ccPlqiuLQ5lOMVUKMTVbE9aXuGNsrgvnIlPsIaQln+hr1QswqdwQSaeh58hFwO
bC10BtjDL4cW9PPejR8lHmt3XAlvtCWiDSBKpozcv7gNbutgxCuMpUKuw0H+0j+qbX/mhT1C1F/E
ckwWN8fokMdHfHta0SByaS7kPHPMEzZD3qIRYl72Z2p8mb0qk3Bbiyld64VrQmmEu5E7qytztHac
Hbjdd5PVWFdQVW+n5+yHRZdcz/mq4rwAI9dOvDgCF8xiDZ7uwyjK+RJdqZliYTECM1d5NSFjFViT
vH0F9ccJ938/+RMusZWXQbyTxB2DE/jfTbHCNmQGRU6Az0vYya/jPA/EEGrMeRYf2vzaCwP7VX2g
msQfgZ2sa2TEbFNcBsaHXSp1nsHv15SXt3M3zgss5xyhZbiAlQhh1biFndv0zB2RLc6Z4sRuyNmB
cdSJ5CyLeU9Jv58xRp70K5YJTCO5Iyfdgss5Oy+bLqJ4ZHydK6wC+A/zi72sdD6nCUY8gI8QjNFx
dpm7X6HGCRH9L2V9AT+jYw2LU0h1U+Bus7dg+lCbg74EVTjqoKeTApmYNiPlQPrGimb7Deshx2T7
X/4BX7FHVLvj7+Ds5pKuDnWAT0/HxB5tDd8blF1cGaQ1V7N8pJScA+oBIisWL+GxbTfEVgFBb0iA
SV4W/S2XrSzV5bwn4SkB4v6uJeMS3k3U0+wBPKJorY57iTHkyLXCDY2HXDFVwQ41mFeq4cJuxZju
RDI5qbG1SrI0s2U2lcqtrpnp1l9xOifyaJJyg1Et/egFiImz8J6iGVomWSBt7n/10kIAzZsmcJW1
hdZ8Y3n+NK7H/8kSFHCGeaqD5eH7exnJ7ujPw/H25Me/te5zrk5bK5jnuT3NEslXpFZkUUdldL2R
VPaevFit7fHEA4QLR+YPm5cnd2jeK0f0xkIygm2HXwmJZZlegfsewX4aAay+MKJpf10uCamK/cMH
/ipnSQk94A5yV+vHUyljmnCBM4kcmDJtQIK5oIbaVS6az5powKUzJWZ3jf2BEr+uZ52MmF6++h6J
O6Wc/cKOVgmPiSfuA2frjYQLpYzRryse9ll2t/wG1RxQp88M5gjnDPlkEeRwiqUTpaO+2EmUSLbU
kIEIaAg5NHEvbAnCkO/d0WapeGF74eoHLwtOi1iXH3UBlPRH8/SAUtV7pDLFM/qlzQ0WS27NgDJl
/1vhEUmi5MHlhbgeIvTRBzxXuq0uy86bRzDRLLaIFA4UkODCoR7pFdFiCzdmopCJiyUu8+XT2EZO
5Ddo3GBisMovrR4ge6gNA4jxkCVYJ/3Ov/GbOEHZvc5eRqMC3142Qi4vAdC61IzFhEPp5tu5+7pX
QKIFy+G227rZCm1+X3x1XlQJeCP0RBER8B/jK5XkH9xylFKbTWf1nlXLOCsOS3y2E5i1GEnS2xEk
yJrlQDIUMfck9810LyQYxfPvgPHnE5QT/zxdXoflQ3oRc8sVQLQkn5TUAnRZ0mSjQSjg2Slao+Dj
SGd+KqVXjQ2ZvNw02wEnx/BmKImpWxoRCVe3aptvH06pdfoYFIKyKruVp+brjjqHGPSeLEJwjmTD
tqynNuHSj2aObjOy2H/8C4BOvPfMZQ/7eFmNw+4MhriEqJsLQqd1jPvZinbbWdKb1ou++cepw3ok
3cWwBF6mVgqBSAF4uXnjiuBtZ7XKNX+9XQJtqi/Pxx6hbos1QD5Wi8riGKzD/fUGlRMCnzWXAoiI
Aq3ncKnYfqOlBxFaGZGXY4/y3kUSOIRMa1EUxiWpm7xy8EPqlmKrie0S9AzXOy4nk2vdHE3qCmq0
CjFJb6t3kBHaXj96+sq4kpbq6bTHUsD8SbubWG9HxfPytmKJyUWs7qROp2xr26f7SmfaiikWImGj
52dSUYDIXjPOxDPly9I/fewIUucsoxFtUBlC3vI7YbtXoi7LyGjCkW+Zs+ZidEtfsz/A/X5yMBl1
jVjEbf73nBIMTd4kLLkgtog95VJMSw81DklsFRiC3vWCuDndqBg7MsB7aM6DAvv5JUOo5Lus+3We
rrWnVOWkMH/1Fe93qy3Lm3ex43EtkINgIHKB4xfKwB2dBN7ED9G9R4fR8ip7VkSPtINNAlseL9G1
TYwdL+/sRqi0iAAJWt84vtkMiHAM8V1u1JAF7DMTRbeJx9lumEdtZptjXCfmdLdKTt14oUyylLcY
QnhmSKUHNF7655W4AMA0VDYSOkCJ4P9xj6T6/+NOqWSl17JeieaafL4uoq3u44NNnlNdOi1YX6eC
Bty3GlAd/9f3wKW1iDcLyWQWltz092YbA4fXhVC7ABPhPqIaDKNsaXruoR9bRrrVKpWPryBxHP1+
C1ITLd4RiMA3o/aGzGw7aXjkReqn/KDaWT2rF40fdbjXfi9CZlplktp+MmEmWfdQuD/4ldxyNvLx
ZVd4B8V8PbiZvz33eQhr18r1c0oyHzQc4ewlHoLsuFbf9SVaF/Zb7aWoD+BQYyKX0wrSujpGUhsX
ycqRTvQn1/jCppDvxLMe0kgb531K/731aDsnrrpCr80Qt4Aua3LvUOGRzLS9dyqYqGqygCeT8vdH
JMQQqPmOHpH8+GYQRDv4hDLKjU8Q8hTR7ghE66+xnyD1bJpJFpF9jHVP19GDOY1WnylCMbBf68KM
aHoc3pXWnmuwahrCoJ6kIFpm44xbR2XOTOlN0gRNuB7ovAnEPCFpn3uF4bu/klghjv6hXLnWril+
0dxXoNz8bryLH3gA5JDjarlVCUUzABR5qGrGl0DmRJpbBzw8rU9Uevqf9EsvDV8kSI0B7ZdfUp3d
ukwSVc4dpKu3pNRysmi6Mb0K3gLcAsPY0nzUl/lfwkSjCumCk6On1939XHFz6v2CEtpGMKlleatE
YeOXv90pk7Z6jg8FshBC3E0xNKlNMe2ZryYMn9ryOUp6rocopuu60EtvemcMSDNFaO8i9zWZkVN2
cWV1ZDISzuBfvruxbV18zhle+QKtSyTQYhOtSFCyHmiAGqfBeHd2IkDV+FyMFTDsXGa3Bz2QqqxJ
TGduoXaHnt4xVfBV4Q12dAvmuyYA9BWJiWSoPrYg09JbLJYZ4LqU8Rv9m3bZy6dx0uhZvQv3bZYe
egAULBpz40HJNf/Qr/mOjgMXGQYSaow1o9CTk4Epk5Fqdsnikl1Bmxi5E2XubQwoJOmX6MwBds6M
xC+bB5A8qo76IGj6ukukz3F6epi443952shADiCf6mzQ5kB2xZ8A4SbFGmvNHy57VHAKTxCCnJFq
oUq7iduaRO0J+s7CqKy5G5T29OkXDR0gRxegPl9FriWCQCtnJreieEO9IH4s3Lnzmv+ntnXPiG1T
Z/0YsvYDJaAIfxW4uqBsbFwGQv+wONwVTTIuzyw0NnrQzMwYw5cZB78Aq8E/aBOBFhnPateqXafp
NNSMDCEzkLYs9qDRb+6w6YRjierVOMYViHbdcLgDbDbRK8aoveqUUSvPW5xbZqjgX22WQGQVKzw8
O4rKFMtsb3WXtABi8YSZF17qoHjZhznd39ur7WcQKjruRl8dybgqlEjrHgeYS5ck/PajEpJHbJHW
QzuXQafhJuaPe2mk3iaARhx+rXp36RP9RBBhTHW6PVYhvDx/sipwm0EgA1dfBwNM0jvlyYWkDrX6
2jvVOrdl+RJkuBLLTfbkmm3pjwT4/lEphDJpbiHMdl5cB/JMCNzuwvhiwwd+oXKqnOQ7tGys1av1
eVb2UCeEkhQt06Ges/tSZ3Gg7+Zk9utBlLp2/AYWzvjiDgewmUjot4hyCJ6L2BFF5amRT12TjGv2
Uh7lwxt7qY6s/PX8JT8pDAIUc9iGoIBMR5kg94kBeJbtWDgxFQ3yUY//y/w9+dQD6VwHuZH4w9um
IP+LNGL2eZfjXeyb0+ZpDqO16sb4EVIO1c+jO2BIh/FFaA2ie32OCMSLwp9p7d38TZvuaPZg4c9k
wGta4YcB4Q3ebkjgv8NjVtnOLPpqqiGENysxqtsm7ckYozz1U8Ap1CZNismsy/TlAROoSLXx+Hi6
7sgGRvH4kA2R+++b23RvP7DXwY2HIWSFDqq3tFPXGqmeXexoHb4+Cj3QNxyUxxg8vB83tIDSrewq
R+J+Zf/lIorNYKssZUaETCCDfC7en0fk+zyZv67R6ix8YCH2LharU3vBkLZWdJF7coKNaqzmfTkJ
A7AK1cjSjjJSyZt9GkT6zzark0WXVsRK6ctXFYDZ8sIoDADZEyW9bZldLqNBg0njcVj7wfGkWL0P
x76iGDUXt+tiTpDox+frrxPwOWA8YolpnP04tbAKHSTsLUgSKB/ue86wYqbop2Hyt3C4KVO6swl9
rQ7yeiyAq6CbRHfb3IX1oqdnmxGXi4GloRL5mrt8HVNtzvLf4JK0Z9Omszpj7/F43rGh1y/BI61i
makuE0RxeJMkNdxGCvD+XKps/kFYoeRk1sdrGy1LpiA3HvFQ8E5mBTMU4ucZuua+ytsIKWhjv0oQ
FBcW5TCsaA8aEBKQhN8F3pS+RHskH0TnT8xsf/Y8M5nHZmQXCUygFIWxEF8rZ/6YCdHjA2CjnP2z
B+9HPBjeOC8f1DA+lAWJCbxYtkL2gQtoJKfDUKwEvgrr54fwJqXaNInbj3kZxjH+Bzq5GmJ5cvnr
web3cwZq7jk1qWtlsMZK7gBpvY3uv1GpV/dG/lfjT+79FjfshvOd/4X5PgtBEQjYRjgT+J7M8I3N
jbpL1jN2GXU84UHyBTnCCpjzK640AfI+KecXgOQI3Opl70HBnhmr4ZkqPZKLlenN1Vs9pPGUuIa8
MmFOHXe4urNRx4zHYFmC8QmrEdSZE6kJnctDa21wpD19Ed4P8OyMaYeOGqNp0+UbyZ9iP+xQRSg7
z3ABL5DEXHAl48a5zygOMVFY/oQ8llMZIQeTGl6GZGfe2QXbHvijQycRt+31AgndltNvBtY3rcbm
S7Vf51ZwbS0wb2GTJpTk8KaiwrKy9wjYF+c7GZR4+9iD9xiyNG1osg7m0NrZoVaKMj1t+Rlv6dSi
07+WCLPjauw6YgA9b0oys9hHV61al271n4v//9Fh8j6jcE9kKWxSSNMDSUniWk19Y+EKETW7vn8V
mdPWgj7LBw2gWa+fb4aI42h/jnBT10X8XwVpE3j2VsrlWyEkGsTguhZl38EXk6B/+K/Cop2+xB4j
nF7mbF9gO7EVlbJWJuNg39ImRc2EmxSRSWuTu8WcCOhM3F6eJ2SftQeRVmMXCISzGkNJyrC3MzKa
Ll/9BYT+j0g9UTZDDc45dxifxZXm0oEY4itDjrQX9bM9xklaA/BQaVCwOuiU7Z/7s46KO/i4Auce
TZBszeNLTwj6JgzLcxG0i6tScZGvi1ioQtAlV7DAC0rmXXWGLjSgYdce/YJCUHIyh1J0KcMtJNLA
mvTRvniTXOGUTMt+TUGDRP2pz/MFsXowO10IKrBVNypt8qdPHdvfsxXHh7kPyKsUO/loQTowc3Z2
Rer03cueH1BLr53J9idPVqR5VRnrMz/qZf0iXh2NXIdhbVNRvLhmqR9hycaBloefDzMFoabi06nQ
OADHSHmqkMq/5GVrBYKqd3i8oy5tIVXsJbxlXI5htJHAjioUwBayD1d+xMG8Gjg/770bQ3UurOy4
RWr60yjcHAeJdBy06M7RWTxGZg+CVAZSirxGWbb44b8xGeAxw293ZJZOoIVRZFh7srqlJIsfm2qV
g0hXcDwaYjlbMTggds6p4muRCFa6En7ZLRv64EUehjUKWT/ThZTkNZm1FN+mTZLjVopjAFqd3Sx2
aN/PKHuXD1FSVmQ36MjYLfKsyw4nuz1MpL0FxO24LpxzbcWQ3m4rtgBcXj/NiPaGJZMCmAbTsmDW
bvnhxg6ywoNYvSywU2+z7qZVCpqD+dtv1qWFiZv/b+KkkZbd68ahfzOSmvjDmL3OGYfEga0CvDhY
xAYYhv9Yj4kDBL/H+UcSjNLb2OoEg3IMLHYFYpZWXiQmo0nH7B+yKgsQhy73g7HBX2LMP9O47uce
Yfo2nRxdQbYrmmUzv18I5DxFhmUiiOdYjHH1jg4oeLpRldrJyF+N2CYOgO1mDRUy559BondPGKGN
F4ihh6Ztyry+Hpd9lr4J1S5X7GOwVCn3kHlmMKix/JQW5CxQAb/X7YmcLDupMAgnnY8tp9uEYjAd
fm18PM1IxQ65s+bRqCfulOVfKE/xNa+sEK/vPARZHuL2fT7ZQVgwHPD2SPD03T7A48YkSZLfVwm8
/crYCGfynHdGFMhgqyAfp28tsyPuF7wr/Yn/k20CZZVhLMT7AOeNyUr7ivHAnWJclYBZB4nmt9DS
ZGCh+zS+ZeeL88AOQA3vq2Tk7NDDQNcDtJ3niLQnglPBzDceEJ0RJPKjNdZgRZiZWGQczCdclo40
1sz1ftqtCruM3YGj5YIS1JZTkCsi67eUtT9M0AmGMed2iLiZSEiG8kUJfosquqDw1zHT++yuSQrd
NRkTiYHN0ackZMeZNlxYhnafq6yOO8miJh6i50QxsOWOMtNqmHnLlwCBYk1Q/rwaM0HCGWS/qkJD
kcC9C7HhfNn4qw82ABPca2ll33VLW3risC+r2rNubqIGnclPro3lpQyhUuC1p/LIcko/ctP1v0km
bEPbqKHq8aBBfkgSvGUYPKjyz2iWBiElYyfVKf6YiqLPvebfJTB6giKBUDVefsucGxtfE76fKiS0
+Z5MuMQBlwKl70dNC1k1r134wGred1wDf6WH7YCi4/o4SOIw1/qwQ2YZTesNu1j7qAP8X7c1yvcF
KHxOrc2pXeh4b8VZraOQdDLf0ItjLPh3tD39H88CI3jzl6P9eGdr0Qz4QfU//yVvZSnWulAtyJl/
noG8etxkj0xWwfAwIdxmKzawuESlHq8uvnKtrUC//KNn8z4unKfV27IWsEtfg6xVbC0R5E4jPoIM
9iZ4WFvond4tk3CJnpJbbxZe0NO2C9oo2Wq054/HfkgkFSC5NgWMDcSJ/YJf4amRcj/Y7ZBa7hK4
ZpzSKMm8U3co81R3vwCf1M3nqxpPb3c=
`protect end_protected

