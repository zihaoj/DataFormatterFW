

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BDznumM1W1eztEWVTvKjiMrW/yR0QpBvgUkowASRlDF8GAWZFC9GGmnkJ5VHp3MvUvUaeihdVeXW
Oa5aZPGGOw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HY72OWgnzmDl7/Gp0YBSCjXdWXnXwGe0nqTlZ8ZTx1RabNWXsEL58Dut4EPoioN8cYxnG1OFX+eV
ry2RjsTlOHGV1nJURc+uRS2Tni0+zwGLpda3vAqh2Cj+kSMeYs1p9/N50zg3ombi8t5fY7t+hig2
nTssvVb7qFJ92IylQpw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
imSFK2hCUfblpG2zlDV1ZPRhAW7A1gZX+Bab2Ck/1vm5FveKXaLcOgnRJ5Rn/qdr6L/67JEUomaY
IPWOFSNM3u1yP0HlB01Q0+L2RY8+1XhUJMg5mDwMNz1gJJt70L0fsHsyzo/frvLG5RqkRqN34MZA
HvVDnPgJGPgF/NnTxhYJYkedrjnFlfIyC/ncEZJD73VfSgenGMOvUf5EGz1ji+M4tm+ec5dOVxWQ
gfVvYfOSuGkFvdokultsw3Xo/dLCki1S3Pezk9d8xRUrCWxy+Hdod0ay96OlkvmMyNTLFpfoY09Y
kXTrf/oEV8BZlQX+/HJlNRXGeVktu15Wu0Lrgg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JVQ+pDCh3zh3ADzjmHakrTo3lZ+0uly7pH2iyfQcD7e4kHZJ5Cj73qHR+fDaZeLL/dKkA8u3YKh/
wbrRUGnxY6mUSUvz+zDwB9zw3T5LexaSqMnrx4SufD5q/8xthrj4KllgycqN8KNA+CAhKtGKvP3l
uP2NSsHtwFK27y9rAng=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ydr8Zyyeie64n9LQFWuYsXtLyZ+C+2YaUB5ukT8402/ILmS8rsTWJKz8WTyC/whqfjJPgcyYFHfh
8oF9YO5rq2/lXFzP99CPFUu6v4MGWDgwqaJH/VCfWseA0uUPIBUaASLog8vNSPjKCxey+9sY6jwD
nJHz49GhvGjVrsjitQX9Nhk8Rfr+HUEaz51GxOCXX/sshVKCmHddXGOgHSmTyRYtUG+9958h/c+f
vUhp4RMEm4SuyqTf4NvEn1ew2X9buRQPbvkdxauvXYb/UuqvMzItAWALg3SJ9JKOAHelZtrhuGLq
E6l1+VeLaN0WijEoi/WEV6PeoEf1SJJYa/wcvw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11664)
`protect data_block
iFEuig9V+Sh5T7FPWBB0skc9iiOzVufb7u68Apik49UtQhI/2trVBKnUTsin3tU5SwbangYVcIJb
N/KtmNi8t5hAIw10vKzuXFqqn/2dxNABKk8D/CnEOlhP/E/88NEhs+ZRFDn1gJtJgOahGKv7Rtt0
+WxBu3F6uMSoGwz5qZuOpbrUh8n1vyK3qrJZvAUeH7uvlqHaFrXQ8ZMBBJ8RcPgA0+vx7w9vTEvX
bNfgPxmh8TV86aAPyRh7Kn3Txv5efAjAj6O39O2ZNJNRGSwqFNBtKVJwhuebPLGMhqHVXpPcMvDd
3Kbd51IUAd6SGxGkW+Kr1UaSbejOa9dPkBOd4II+3vT3yRMVyq//+GVW4fjfKP9P7YcmUjNh3ph5
QmcYA38Etz5y/7+U2crSYum2hTjzm9Onbpz5rUkIu6oumIvDv6VybS3S+HXnmdex/pE6v0sl9Rwu
kvWgZMYw+QzbdLzdKP7Q8ZukclQFtsiKgK4DdaFjhRkGHReJCccAdktjdBeTCIk3OiV20OvpO7S9
lYQjJzZA7H3HCzSIOS4j1St5H9P7RMifvOfuFS7+Y1gbFnVCnTKr2ivAtTPsY7nZmqWkRdrQZw51
dhJkERbTXTnTyIdW/73sioq4VJ7qSSFGJ+TvA+A3ryaKVABllem4kgn1UMNIlnPLFDCTGwB22Hj/
84lkDqrdV5Bv5G2RADqp22hiItQsMbTY6/nNInBoqDLilnQ6jCDxCfhp3UnXFGXfSsdKc0/BZ91J
TLAEHR+rILsTEAfGIlsVEbnkIkUd5eu8fmNM9HAiozDL+Q36REpMmlAT4i4mYXiq+CYKnUfZ/Jej
wb41uUmPiBqS4hSJ0j9dQ5ARmjEl9kdAtpN6kBookzBYkOb5wDr2VCI1fjmAoEgediL8F2r+i/xy
JTmNQVZok1KjqwNd+hO/D4HP02ww8GZE9ekW2noekm3w8kLniEkKOnTeMD2vfq9L0M6kOiKAPFQN
P5iW5NOh9FVi9U7fKw8X+8W5gm8Gwe0TvFicX3gV+ezqdAeUiNsGLUF/RIulvT704uHGgmzHOn6D
lZmpnht+jbQC2kwf+BnFxibnMh3WvAfQjhRNuhuqTFVPiV3Jn7JDEPZk/luPq/anXUbwFiakPr9J
DJjLzRtmRY+cZJR2ZUAwTw2qAz+giaIKZScApczTwS5wE8sbpwjaesDqCi0fs8G86mQakc1LqfrW
Rmk3m18hQsoYvbxKy5/W61cH6Mw6H0gTePxIsMuE/DDBZjXVlM2qS/ojMskWwRw8P1Ma4H5Ed7Ib
SJKFw+xVZwe1zpuU9nuPgYEvvefvllhYWrettR8d00PKtNt3UDa9TIEB6ThX3WJtfRsaFvV+1rfG
ARyn4X3RC3bS0X4nLSdJ47EkPslwgO8RSe1+Fefd85AgMIDSvlpfhLT5fzCFHsMRaMNlHKtl0PV2
LETDGRcIwV+r8ipCzdo+2MRJ8gotrbuB3vTawoa6jmM9fGB99l0uljbsMXFOK8NJBYx9FuohzKBW
CfK20Oh9COwL9j0KQif27VYEOvS5H73Rj8TKFIFduNM06eDAUjGhIhjf1eR+DAoU2Zb7KsZ+dSL0
6n/2XNRQju+mJPTlZSZytQVbI04unEGU1eId3Pvcf+lI6Wy9cIfZmAJkdWhs1jJbk/JUgMNDIlJS
pYKDwfwiR/Ia4+0DtRi+vIxpgyhBKsyEs06B6q69UxnVEV3jLvpLRoZ0K/wTf0qbeyWJbkLVnJWV
N9vLg9X8fckNRPfeso2C3ZfY4/yBrqzSsZTow4NVo9ztiid/eyumkLHAavwzeUF2ZYq7cLsiHRsf
kXWr1EUsnenwyyjVwikMBYHcCdt3y+BRN7rj6rEfQVysJCdBWKPwauyUp3RHUl+cxj8gcIzVYQTe
EiKU0Qa1uisAwbFqLYcVhCbQ6yoOpTJUBY8O9Ye2jvxKhQjAd0lvRDgB8grBtKZ7an9dBaFxduo3
wNmusC9CagHVWptxKfx1/OJ8be/oFMZGArrPcd5bF6lcPy5m+GXfatIV9OMeDit9ro8i6bE36Rev
fpHm0VqZduaq5sTSwpSfUuFeCLqqQp7eM56Pajs2GgC7hK//oTn4mVTq8DxHYu4rTx2AV+/cQmdS
K5sefrBEXRVWoFnINnf1bhNYA3ItpqEC1jt+nz8qFCn+jdqwXBGBiI7+xpOaoscf2f2awTBYEXEi
CvcG7AL9FowXPEvHcjQ5EEdbzkTpW5pU2UVVuWFBUY3r00HrQLcfFpl+7FnYEsEJ2q2gB4yh+rOR
5bTszbn3UbOvxzNt7HEJgaQJOd1H0V0pAdtCsO4/M1lLzZY0HWqDLciisxgODuLL0EWXmFTdD4Pk
Avhwah5u7MLH29zINHnwW4orxAuEqfCt/9cvlrk1jLtX61iIJSG1s2VUdMD0idPv4nb5dsn1L/83
1A1tuOqzeVPJOqoGRJDg6ucLJrA5jLWJz6tBjQy0ljDoPTVyfKsBam5jPaLllxmlHEo/VQqSaE0R
ugcdJETZlYBlq0MNkdjz2A2Np/+zW8t6HcLJ0u4odl0OevsrSmRFOTC7NDMC3Om7K+xkirgXaRrG
bkIH0MyZBpMRS4j6nIvIdsl0X4VycHJPB+Ii/hwms2edEW8UdTeQ3rJwl8eY1o6qBiDVs1beJu3s
9Hk/jis2ktZWa6lZR8vADjKpnd4xXUmr6gvUpRTAwmZqsb+upyK5MIHUBx6TZ+LZF30Ldsov/ajD
toStlYw+Mg+HQJLqssWO45Rm+3TfM0Zt423MM8faiC8CgkBOKm+xeYmbm2cks9g1LMsN++JKPDtP
GBgR3hf4UkZC62TwDX6WAnpIuKHdIDAMsADlg5ciZ0IbOVSDrUPwVAnjzyUUs2H2xjdL6nV/GkHC
smZeu3IWoDq4Is2fOAA0UpK1U/Rb1wLhIE88lNxmWbvBxitjJ8FCiNhr2cIT+lan2uYaFa8bCR6K
+XJMi2w4ztoXIvJVMiV/RM3+X1140dWCjm3Z3FCHvMQD2bFkWzacUgBGRvNOCcoDMRMiSAbDnD/u
eKsvVy07j6Y7l8M+nkb0HMOY3P4RoqzxdytwyJ2/1dIl+OOXy7DpP3c2fGhHRbk689Tmwge1KBrz
21V2SnhxtDVMX/lfd4iAtOB3OI93BRYyFzlVnroOkF478EaFr67gv9SbIKL2UJVReD3G0CROOY8b
EKjCpbZ3FpHayPSjadHh6XR386KizdXi27JCYSeej1QxkNKI5ry49Zqhag3tloFm9ImKIar4N25f
/UpzH0aU1WXNK0asJqHE4ji5nX1Ep6Xq0VwKraITg5GKbcpTlTlRU5zw+Nbgqk6YEyqpxzm7spDt
iESvlKWtCDFR4g3JYIiblYG33HYPBdFK8NomMbBhMjROtTAoG6J2R4aQSE8kuWAG8PzNfEIUgX0B
ciyMxmwU+qbCGDsK7G+XQ96K8m+z2vEs6bqD8VogeL0K2uutQjHcXMEnQIhm2SUn59dnrOXAJysh
ZgX9QVct5LWhBa2e26yDgyhkDbLfKsMiTNWuu5HfgFJzb8Rhclxv7dSBmPKx37k8U9oOPdKGPgbd
5bfcBtt5SKI+QO3PDLwG7MkNa17/Q92spFwZEbYH4GVFzrDxU6xnYt920lm6bjZQfP4i63ahuYUX
yatzIdWd7NstpLcc0Qb/RYxlZf/ndV68jmSWk9b67InhHNQnBhsXNz29yhOFklVq53YOy8QN+0VU
16+XDoU9lZzkSH+qfsC8aRcdYgMuOl6SHJ7XgEtmmiDrRuJ5QgRwhynWNIKZj7dMhBAdl9aK2GKk
w7iujIk8jvQmivRLdRx6GZS9HWp+xJg78IUpoCP2TPOYo6zF7lXGq9Cfp1V6tKmu/2bOleavKWHj
hGqAuhuj2mbARQQjRdhNXCXGoWJLIm8Ena3r2xPDR9N0k4nRvtdTL6E+g28Oma6YUR50lF0ZlTRq
hK3EXqvteiGUXiJ2ssx+qpuQF+Sek76+TT+aSUjVFYMSfjeTMI5+F21+R0jwkde1AKi1xYJWhFYE
J2lfoLfQ5CGkR4yFZMIrM8Q3JSIinPCP7i+WzxfRuaQrNFxSfxYdQs4NEcWZ0vJxYKBeKZXX6JiC
X3S4aLiMtPVw85x2f0s95llFCYUNLCXG8/WkAPoSovqnSpcjq5bGnv0kpGrM/ujUTfvaX0W5zh/T
cdYGEKM18Eick6QS9BGKLO+CK/wgsBCvf6sSbfT6BB+wzQw2IsaQJMt2B0ej44+BhxARumnFGuf+
Vn0feDX+wPKONjXZ+qbiDxjxT5gT7Ob+rYJL7anHlGi+K9ylY9yMwZYEBumLeGbV480vtD1KEtw7
C5bT3FEUeH6tLJlE74EpoEmxwIaqIAXItmMtPpWPZwHHxkJ3qcgxX6EXVjOPKMfU9ZtPlV+9phig
hiasm1hfL1cvJDV/ZZZda347yrSuF/heDp9WigVFFwrFOxUBBOzmnMYXPJjKvTMh7fs7RgwsKxD/
q11dVoiDX46/UdQiYwPoW+Emsa+A8CsqHaiuljDslTeX1gKoTZOxfArRMGlrHQv63yQpsKU3U6e5
0Zn3hcT0kFPOnCDwY7R5BzdqA97ilmZfEVap0cECKQw8GX15e5G08nUu8T7399yETrlHfTbL42g8
VtDuJYq+O/p7YFwLWsi/0vvNUldN2pXtNu3DtvsBalYphzcGxDqEcLFLCWJ93qdZEaKEM0eJDaHZ
/ZkkTm/iwV+uJhs5QQu/ktHa/z598MdfSdkHdpeskA2/Gfj0M/CmNhTIX5TvexKB9TqNhVn5lVzB
toNAdDl7HD7mqhzPWWWGcBr8ejpfmqEU9HjUl+wc1YVdctImfXS3+wgrdRCDWVqglVRsdygF+CnJ
kj+AKOr8zC3dES5J0fqcJfoO7LEZXz/TnonW4lscC6Bx//GJarSBwb65xDjAAaSf2Z/PaprTng2C
ldW5nvZLd2ByWubZuDyq8RBVb7bE0Lz4n0yHm0dS7WgdsXkzB6A1A8NkLtkcKpi45iAKd8bOFZFH
Y+M9g5hj4JstoxFYKie1FwaHrTuOpA323U5I2IT6Jl1jNHFVf0fm0a0XohX8d6G6kG3ezf/NCjog
b7Pt8xPUzBSGKuOlT2n0ZVzJG4ejWMc/n2IVPCJMWKEcRm9Sj+uoLYNHQjR0q4oKYDzPI8OR+fNS
rbQqwaf47QhAOnwSuzj9HP2M0jFLsLvxGoPgKbvRIEU4BU53T7t+Ghs2TABNpUeBRnpbyO1o1huE
mpJVWFDG3ivywUUUhW3VDFDskqo8KtOxKWSqL75tgDcvYdyXxBF3AsiKS0M7at3H2AoEFG00qVL1
Rh35W8qAGGJUnxF/gZY7Dg2ipZfTgJCN3D61X80NVvcm6qS0MVqE7CiyEhPzz2HcfbalX9zU+pUW
BCVCN4564SkCftqc1h6J3YdJbQsqbK/eNv8jbelYdljahnVfmTPr4RUl9Ii22NO3HdlkxnQOtDZY
R9RtA4oux7lz312QgVY7ET4VW0lpvSfg09WIw6Cuj3luZzu0/88u+l1eChIyaHGVbjehRCAdPRW2
gl38tTe6OvVdQ25JriXPqXvMgBInwPU9nBErd2Hi678O8eXTTxl9ZItGl7mcKAHl3pcFG/t1Olmg
8tK996MBBnPggO7477AyQMVq6yA1/GFlqkXRYtvShv+QFjZl6nbjGeoTRSCH4mIO2O8QFig/TGuE
30wOEyMHRNysNHTwQyz9FJW9cZkfa7p+Kn4DrpiGOZs61BVndzkyj1tkcuRQmxCGLtBTiC0J1/f+
Kp8ylDZIIgDWWf/OS/r/vRLrTO8Cv1szEKHvhaZ8XjyhNHmoH2ge6U5Jl+Z6RLpl/LVfiWfcuD/Y
txIExxRmpJe6/hc4PMttafW21uwyKcL/IPAeijPCWbd5qxedZzKCQUFq5NZnUWiOkQCl69v78csC
P1R8V0cRkEQTKgpjZsCJbsUvonDyIL1kTfmXL8GMMrBZKFEZZiOkppNU5DtJFznfx8CPapmUxIeY
rILTuDsjCQ0RJGOj5z3SzTkrfu+QOvGLZFe1D8Mv1c7PcxYqhaeG10cUNmpfHfx+QcQQEYrzyd3Q
PueN24/5fNuR/Ov2g563lu9JeyGyPHCiLgg4yTKFAJwK77b6CO3V7Zkok6uB112kFqCBid3yrdbQ
nxcFr1jXiqyj6eimeZYdGUtl5BtSLR4gl2+tIpTuP8xjUS/MyncNU8w7Eeykn9mXnqth++WpT4qo
pebULnMfJiMf0/F6S2tRpnT9r3ywRuZjMJR2yemCDrgRSv2p9PrgGfBQexu0G5C1PWgB3VVSn5il
Q93F0kZbVgBNvJEM4A+CohAwB/KyoFX60xe8LH8zkRXR5snErwfGxWy3QLSDPO9BAMFxnCUJeuys
fqxENYM2Ff6Cg6km2wggvvsshhckGGeBz8SG9lVNoaoeGWLbkYRNEau5iWLj2cSbDjQrY1NwZb2f
ej0uqhkPXHYd/mUJ7j75npAfAuE1POE8gL7BOHvYOjCoTdZHeeGr8akXpWje+YGspdDQw4/k8JqE
BX80UmqA8enGAYEKUeeYAhNrmssX3ENQkJq+MKHG+/DkLxxpkdRguKB2cZCuoqTDe3/C59R31iH/
efsVE9ehlbtiFRtDu8MSpUR4eXlfACzdolC8jWY3vfpi+RpLq1yqCnv8jTJLNaX7sWfLm4kv13G3
Pqo4HA95oFutccFYwCISiwxdlnli5W7Wr9atz+ZWCFRS6aV3KPbZ895bj92dNF8WJjKSp31mVNPZ
obTRUbzqnGRbE+ntCTpCzkDBxdEderx/70GYtpN4FdwNxYDLTTcNOu0d3i+shb+CNdbL5v2wbWbG
dle9sabK9AM/+D6GzcggyJ+wVorxHYoOoVlNWggP85AwROQvMn8DB/uUTcIhZcG82iNazL/wx1mp
hHC3DjnSlcJj96BRdQdoDqwamewkzUnUFYOqLpzwEQzSh8D7g7f9VijxkZ1IrfJrUPRaB+kX0dHg
wi+gY3EfRJ39SbX5jkXgE3puHSv9PT0iDBMbI0SR4Iz6ZhVKkfUGfw4t3uIFS3JZNGmZppDctZna
WvBboqvv11H89HXCBMZJDVSGRtaE8or0Ura3HyLgseAIHoMLetAhmqMwvuW0jVxo7ItUQjSaFDva
GN9gIDtyaOV28OD7v4yPy4ayWW7f+Q7JTjsPNv2Zb0xpDn+9qKFLOyiClIno+/HX4zUTYs/VXia4
Fl3lFI5FkwSoTsbzleOcDfEzQ3GRMoXViseii2vhZ9mkA8SdvpJLaeinnmbCfAYHlwxeKG7iCEAE
ICWmoV77sYBKWa5m05yA/8pazM6t/SipYxR3Y6hR6td/Oy/fnyMIXVvP7tuh9A9yPhWkGBRkZ9q+
EUehtP8tHH1XBtHiB9DJTJQiFTxHIkaF7d21y+lQkOYzzswNZ8sGhcfCLnEREm+Rwi1qA315lfA4
5idKbp8+lhHc7H1Yjv5lYU77YBBUinKKrh4Zv7vC3sBedvAsBTkDZr0nvVEOjY5C3fVzEtkNjFQw
PpAazDh8ONGCPFt+XMkSt6QuoMyliZZV3fWhaDBgBG5fxALcYBNvqAqt6uhYBINOmGVjOVGdCXQ7
I5z0rNlenIgku+jhB+y7kBrosWqPcO0UzJdM06QRXp8oSuc7Cv6UZzDEYMxKac0HbM+zmiSLFET8
mfn1ngG+hRXS399gEhtJcRf82q1+rEOVEQzfD9zHRxgiDJLHWksBywRY1coKgs+CqmBmhdcPC7O/
loElVJ1H5m0G0cgn9hE7n4Tt76KXaM/PUWuCL820h/uw65f2wIm64B1Rya+dM9n4yI9jaYn0WVhp
m5yh1JraaivOPFC9IROcg3ZVq0y8Cvdtm/bghblNh3XEPXoXdUkFv4lHKsqtQOzw2WDbftjwyLgw
19pDHY6ldbWyor9mT3bbpuSab+KE1wv7Hw6ZJ01bKooA3old991hDL6MNyXIqIcqs5TZ+MziewOF
uFdslmFDSzdtWoThtA8w/cqzzBLSsjdmCmfpa9YwyTel3wgJqcUIdGnziDV/jczKChjEe4ELRIp9
oR1+JGEkosNOUkkgfVS6ZSUA50wlo1Nqkr/FXx+YnkDpZrQg2hZmMM/4he6ccZJAbzA/W980MAPg
vWEvL6ZJw7ANjB6Ned6hq16koAJvLwPJyWv5xAJZ0TCI9D9BnXAdN7vygpjVNS7+wB8+UZDF2X9h
2H4Mv3vhAgpGJO9pfqM6qtF6WqkaK9QADpb40Op2XXEmtlBZ5oKaXBlMMGItZH7VIjRrMEYSHTC9
vdWkJqUmVbGkuPVfJWDW1VoAlPqjFlgwrh7lTxPZ1iPgz78XaHOgkiLvCCGGmgaWyB5hx3MYSRYO
XsL3ap/uNdHbFuVMfHp1NbuGYCiKQmKc9bgvl6eYB/JgjgPZFVFl5h5rC/UqI02EIk9mWpIa/mhB
mALrD4YZ0EAtd4eS2+t0DwxJ8BVyuzRM3FRphppIdMMulMxXG7LmYB4g28HrGMij3CobybkIeQY0
B+pEJrI3xPmw1Ruzj23lWdVFe5zNSv4YpX/DGJVfMwQ/7+dI6UXDkKRWWBj1GxuGvXUkF/oxNFuw
pRzBjnKubUvPuuATrGZKikxFqxLlARCWjSq4/F2hmRwQSOdlkQtfV9KMtgTJJtM7lLhTm2uzNQOl
SR5yIWrrUbEjYa6PI2bTPNBcR6DH9WAKbYMQQASF23q//xKK3yRMYvT6Z+WSznfkG+/8KrmzM1nx
ZVDS20mlKZM7tPtmDHOhv0cXMuXJWex4kro2yhkfGs2oiGtLvpRuTkuS3TBnpDd9R8qiyhpGFRQG
s95flUInyh2kdHnc1hIj6FnXFNcH1YLp/YkIBsVTxwQDQKlQgSUWuf60wXPCK+EMkKixmusuX6U5
Bf4zJFNaduTMKcT8sKsQcbg51cxATEgN9ob7Zmhjy2QwNLGGg2kM16+3LN3L8Gr8Vf86KA7rBjjK
aLGP6OgTYl6JT/2CE+cscSFWtoxF31KFfcUPc3gGCpT3CtjyliAVuc/zXRYjxdqzQiWwENB6uJF/
qeF4P3KUV+ne0Ixl3BHM3BxycWyXSZpgzoQqHK5kiL+XmWjFPAgoiqn86q3L9DKgArEiLduwDT2T
fTWmzUrX42dfaCwc39KZH3ex5q3oPH0d76rVOpqQ67cbHuSwIHLgP3EP01pB+sm5N/yOGUtvok37
hRrVM4TaFmTIxk+eQmPPy/jwVQL6Sbd57CjkTrIgXS3os93y34KLZnIkDnHtKTQHRG/PQRJaP2YQ
Nb/VzBMrt0zJ56I2zvQ4wycheKQ3IA9zhvOFj0wApOl5zeJ/Wi6BcOKvjClm4uTaHMR9Fim2Rr5I
wWomSjnCJra4dBPzO5v5vt2EFrclGxWp6t2qNbX3BYrJx7n6BWoHuN8ZNFkN5ZEKA+Y/bOTR7KaB
eElZUfAUzvAgIyw6T9EfJ98MCGlKu/aALfR1RX+P/+Ea4gQnwxHXAx2+XZ3v6Vgb6Diez4yiTfsr
FhUl7A3gwHl4r4TWJSVkTsv0MfBr3pMjBpMeDP28SN9aG9Q+qFaD8VA/omVBCmMgV7QKdjCCjo7w
zGuvmToQ0ArK+jAT9CYqTa/trRQVHdWRlJI+Bsv7m0QSq9JLjwc/MZHLQtmEicfIzVnXzZ+rWr6J
+CD1WodCVxirG5T4oAwQ39Xp6H8mVIqvMTXN0zr98dd5T8+//8hjh1/89OGNo/N7LqPFhlmCco8T
aEB8UGig1EsEUguWexMNM3Ywdbp+9RCwd/2fAgs1ad9JSl8DhRDhHUqCIqGseovc1z1m7Cfa3VNN
4SDA45NtGFUYOtBGq9z2aQXdVyZGj2WbSk3X/a2E3T7pz0Z9pLW/IEswzouTBx/RqAkfDrLan/WY
iOouCzMuDSqvphsScNWSQUp88+YlhiaugQIFyOImgEiWBRdGWcVEj7aAVx40Han3jnWXb0rmgnPl
lrR4TzY77jDGPmd19XHzFcxzU2hOpScCcza+M2zPElrh4ORMIEhCVLOxlsl1UutlOWVBeOSCOHkS
YRmiqRL+e+NPs/zV1S3aEz2AKTWywV9WAxvr1dMca1ueixDok4eN17aJ1GULQaDbMPO5eb5GRRIv
OSultKhR09Qcj5CtSE1bhPV5jpRhKR80B97I3++T8hE1JrKip95vzzNb/3fLt85TPPvGp0ipq65c
JoMHH0y/lLCHH2YoSNV3roIQ2TqImi9VJfL3HcwHejpHw/szhRU3/ZwhJ37Zw7QkVVBHR3cfF+j+
6jBxchxly1ljGHEk4lQr614Armp43wCrskCZdosIZwuXNzi46687bFfZ5qgJ37ZQvfK9iYKxOfiO
NDOpBM2qbYieC/G98LFMsw/Z0SCk2G4jM7hrp1D0X2SJQPw8Yv6F0YJWyxcUNDI1EdjJnRKPlRW0
LqDvV6/xR4zG2GLTuiW/xPGz8y+4uUE3U23NOYWYSxBLas+TaqfMw0CfEYxp5syyRtCGjDR4gFTI
SzomfqqOFLe7k9GiDAjSIFezn4VCo5LKsY8ddv5Y3KimWPnWs3gYDlgJS2j8BFprF40ghszJea+p
4TndKlif9GjL3dKSDSyaEPEono6/jWhPvjnDIevrCayu6njDz0wC+u0SySWc0UGddjjcscXVGh75
1HqCN3DecNOQu2ZzEVrpmqcar30RI1MJKjbPfhkxmI4AmV+YKT4YQU1UKqTz90WowQrVSZu+IMo6
gLNwb3g6iS71tt3leXYoxEmp9AJmxIIgr9CYTkSAOcnhBOUolMMdbcFj1hcOHZP9Hqh3dqB/Lg1h
HMtOh7NS2RHKbsjJdQXXQ0NtHEQupHOnzXxnv/ie15BOm6SSPb/sFq9F5WHQw8sZBwVvIntVtjyr
VqUKebIZsAj91q7HwI3xQzjeJ7vcFlBaUm3bS7qphoGWoFMbviXN1EdEKppzHOc3lvGjKR2DxMEi
5hfQnXRtSMsSKxKez3Hml847udgbechKStL7ozg99TYXbuwBXr4cVM7ZLiiGgzsjw5i1ZVM1Pa4d
HuYV1zMbJhnuzObrXBfS54iv/2yxJn4eL9oVWkjcmn7A6t0HmPCKNkEYCIDH8mV5Tg48vdNiq87E
nCrYY0V+aPudZBsYb9QOw91EnUh2fh4ogoNysoShOimGRoJ/n+4FEg5vQQop6unCGYshU7B0i9An
ftx8Uic6YXRlpHdZHDgI2RI74TIqu45b04C90FeaehP3pZ9/rNqe0rBQF9s6tIaIZC9vqUnZ54pe
D0zwYRvZ4YPG7aGY1WyU1L0ZudfPA8k8wUohYQzVSaB2Q4z/8d8g5ByRWE+tgf+eaaBgsE1uXTga
wanj2adTYmD31vhLg2534l0ddFcn7eWOJb4Csbp6vOvIEuo1Q/UnpUfjBDL4mAA9QZCEnX6kB2k4
xWxTKkHNfFOg3TP1wouYVhfL5sFa2vVVKWyXbQcr59kdYvEjdYsTWx4mIrVasFNqeUkCBu63FYvI
BJRXPJYXQeDoZ8gPAmWHykp7wfimlrcvf3WvxTbR0qQtDz7YLlT8rcApgXd88IMu6vRVFdtWg6+t
PmeRZQIKDv2c2qY4QtXNiQh8OZTFlqJkh8HfGoWNm9+tjqMBqibYIf8KUHcn7hrp9PQKrEG99CWh
QF7n9FBn3VgsMrtZ4ia9Eo5ktFTGF+bNcHmfFCOGsEdC8uCGjZ6N0nf6o6pS8mcxipxlWx3+aKbm
TfaxrkiEGj+l2aejOQC6F0P/XXHzLk/DiBiHCu3R6h6wlJYR2F3duGp0gEIFOxArUKsWHNiZdRIN
9xjDjqnmRq1oStiNn3RkLQJjBGqsEzHMuxeYJYsbQC+fsFVzvX9BAkWer/umvbdHYbArPwu9PetR
sDTcH4MJpTI9e2O2RlTcnIzT8+WYuFGnMX/DNhWIoBF8k10eCXpPq9Qsh87d7rkP1ijQ3CjvWpmE
e0B7cku86Xlk4/aBp7q0Jiq2Cob03fHsussTw9aocaEQuvav6BIDQu6gOArBZFRAMsL0wlwmZg4F
RnWf/frZY4Fw+81etzsCToZJKtxwBrJGmmjw3Izw8Id/ilTkuo1mBUTiwxh8WSIpwQVkTojyjFE0
wGUe0P49iD2pqG6cRRnAKYTf36Aaphgnk2vUXspBQS1PI6hTyjgPbyxzsdAMr+u2YrU01ej/PrVn
fVQIkWWza49HrqMZoYHWDiFjgNGWKX+b1wf1cGcR2VR4a9soGOU+6NNjKgu1vCClig+Tf/m5WeIX
swFzf3HKOdUeQqAaX9YqkQInQgeRSXz8kYaREsA2YjWDcELOSTryaeBZf8qziq9s8QqM7gYzJbZl
TCKkybidgaz8wdlnuOnfG1JFIl6VuTMoNWqGK+Kn80WAYKFxhw4WiJRRp7ddSBEy0zDiD5h1JRKW
mWnBPWfnKoXlyWrLqI7iKTNTDUZt/pHIQJLP1hmkNKtsFY02gvuDnOaz3R2h3qyyVjDVHhdwCJQY
ju+3PB5jm6HVqdxTRw18Pl2ObeVbdhkdu5PBuYJlzW5m5QDAolUkyyw1Xh4vfTHyspLwuPdbT8Nq
UPik5pA9Zl7wvqBSAySRaGESfHC7cW/cPc4XXq+TkbohgpQM71ZdlPwBcISFCZ5SfGvnDsofhfiW
k7wFJBzs14mjkUoIk4B1JzeImTttIpBfIutYybbe69f39A66hFLWNpg4P1rn3Gf9URjkWvBPXQta
pseHtm2+ya9sUSzn5+WrDYF2R5bROotbg9s29eZm9nb+8sF6zOcRHJ4/L3255MpeAHFXd1CwicIN
+qzjDK5aMRt5f071gwtesCXAolhZwAbZgY5EzOJw/nxV1e4xxz6qum/A/xbGdBH0Hyk9WpoULiUn
S4AUQ3qGMktQvPP8agq1olaDwTkGzyO8R3mDj+YhwuJOHyHPAxtcXKAKV/toYpO22UJu4IvMHE/5
x9duGfHhvEDjOdyrlHkcJ42lllWLDbWCPKkgJRW0iBi66ElK75oP823wlxuBL35qHg6Xg4ZagUYJ
vMKdJv2Ygftk4iR/wZw09yPflpiN1qdKUP8h44nvLvJl9aE/FpyWaacHEDJgvkfqKg+HGuYt2ats
l6t2XilU+E9MuY3qhqayEc3rklyhYa03ysWzgEFctA91b8idfle8mU7UnJNL14avhl8EPyNUBYUG
fhVV/+HULDqdtApvTxSv+PkDnowHKtAoPEHERGcKtyvt0IWL6r66apP5xSysfriuIewmdu/A75o2
RqQTZhfP4UnoeSJ2ti/gr/Eco1aadGwpK2JtnJV+bPSuwgmoYIgggvC9Dq5W/RFYdPBouQ8MxUg7
CFBzDxqlyKBXnpwZwmIEZ1746VWjd663J0t84ktOUKD6X6jV5Ds5dHsy2bB0+ekLkAhVY2v7Rkv4
lKW9Pf17AG6ov3UsJvBGsueZZ0zTFbRyDTEsSq8JzVF0xFf60K4YiuImDhS4oZ2GopQRdM4rOdEq
d+7AweW09Nj4tXxohpI4IChZRcUYVJ3i8Sh0K17Klk8Y7neUOStVcZv4C8sb7FX+ZJxcWnkGT6sW
wxP/8Ijkw/Im99lH9acsvigFff1hZ8SgdrHOLbquruPwdKiJIFvUtm6UZq7yHiZ+F1Mz6YT9AMWl
m4OvSmgNfU4cCP7168xl9wuOzYgAphSGq/GSErgsoH30fCs2NOfTP0hqLyf6GC7AkFoteZz0xZnR
1xsqG+pccQnNYlsFDNLfONumAiA9yHgbUh83RFKdoVRqKTrTyM4vIRUFPZWIea8I4SWHj2w0AaLm
tfUxDEUu92/pB2MIQizDArErI9uGf2iUcLHWin9508hBjv7tr6Z/iRnhMtFiqgyJ76SN04+9cMUh
ufZVDCjQ7n6aIWplzlD51oQYCX3v34+bazj1MfyHo/YOAq29L1AwYTwQDmoWmJl1jjYCevXXigPi
Y/V13yz5pC63DxSwZ86E7QxoxbCzaHeOYB6TreFZ2Q1TWGuCAfgJS6pOMtITmJN9eEDMKjxH5DJu
JLq4Td462KFQpRggPTKshA9vmVi4E2d/EFhNiE/QBM7RADsgFp+AeXrqdr3roLuGNjkAqiJx6p55
TRJvSj3P02tbVtlSXdWmERmUPIVg8GtRKzqY5+MNcReyLaCLbL/2F0GJkSJvFNhokGF13XlX90TR
ziBscG0tracr2HofyRmYXMeVaAscPa8TD29K/TnevmuzfHrtJzoIa+NlkBqGGVzE8J88fKkZkFkM
fzD8laxDTShoQgVgQVD/LQjSZdhu6ay/fLukdDCpfg7R302ZY4pW1u3r78h8WcdEPEolSU3pUzh9
nxhguguIOmkse0FRadCoMlkIrNTBPRRTR9CHEBLXpBpuAYLeUuLk7GtwGOaN/fA/VLAaE7OthAAm
L008UuYWPfuO+F+jKNrcPT3WBbEhCB72mg0DZyCvDH4ezulYnAWKTy/wd6LlxtTmvWnAsOm0b+xF
xgzSSMIPEYuj3dsZHN6XiTW1awPKIz3ppBjRIWQZ0HmJTzIRwASXpclC3m14XR8bAqOFXiU3T9Em
9oGkBKGWegGQRBvuxDpHpHQx2RtqjTxBihJcsMbMBRb4h8ORAKHJ+vBsjfa+QAnhMLBxqmsPC3nc
S5sofhFNYMqXcNnf5lGzrnNOy818BHWDPDbOHnQz6upkG+Ty7JpuBmdXy2+0eMUdiAt2S6lk6HRZ
z+sTx4PjKdbDgtlmv5MrG+U638A5HTPyW/xrYz2vIfmBBZ7awtKHz77NghtejneCmJk0FWCrHtur
Bw3OgWCBtLXNAmiWzyTRqcoC1tBu0/9Xmx3Bu95zuazC4lv9tvUgZTyXGYXWzFK0FFJpIvc/Zcw4
Jq+oatOfNNwqmk1oD9S3arbPzptJSK4tjU+YvQ6r1do2qiMoxz2LuUsYSsdeRhxv3bbvCeTpHZsJ
s3CPf800UU8TDITTyCC/wBp8e8PLe9LK0Ks1TF+OoynZTYAKFmB8Ofs09ShRK6n8SF7ARJ/iXJd3
skJc0AvQWGq+1cEjLpW/7jK/TUCsJ8be+jDa3wYLg2pbq10VqN5Y2/raQc4EhRwE3DoyaD3PDSeT
eLOTZECqxZcnMaVW9ZcuyBI5RacrOfnyoro7megbvXX16CFWMxRIawZt+L0Z4OCR8drq1kXHpsDq
Qo2oEii59Y4nkkYxcMBTtM3O6Jr5o+/0CmuK8LBMkV6mUEijdWMMTq9/Ei/35ZpEmsViBRQhzmIM
iMZhsVVFPyuipIiSRdp9KfqEbbowJ2QSc70RYDqG2Zj12KeH7+pxF1wORFlI0yFDU+AOonnoLFwz
uCLXx8gLTfPLcpBCdmHSKfN20BBflPcvjPR+qECd4iiEmPAojdsFAUY1C/2yMKU3Ea6bOtYJwGBX
QsTwXBBeHzxtAW/HQDH8Hm3TixgaA+9GQUf9QV9In58o1ybeGUVegg7Lq5CngyYSD5zfT8rJLAFb
C2n3+0pz8z1cqqusPyJJoE+PEGZgH+U80LeT5ZYDJqscIbPr3Q1YavtjYUcuYPi773eUaGNHzStu
AsuYBFceQbol+GRLPks308jN03328NFnbDYMwhLaynUkvP8Y
`protect end_protected

