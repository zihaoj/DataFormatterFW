

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IVxyk7XRM4VsQcD0QPYws4xsTeDPKdwWYfreQJ7l1z8C+G+JAKZ2psrNI+b5ecZ2ziPH9MBGr/oY
8XtzCKmjJw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VO3Jpo4aYF9TyVwyAUb3a/oDy8Yhm9ea/9mAjNtuOBRL0qoy0/CWzL7D+bc1SnZvEP4BG903Ildl
dM2y4TNyVTBUaU7Cz+LzZfu9kCPWnmttlx92LcMKLNuvGUMPXmV5jr3PzSFEvoDuCinMqNc8uKFO
Ux/aX6fmBD8AbQfpK30=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qOkimDe0rSU5f1zKvoE8a4lZw1WOOUxh8wtTIN0ys09AXuQuNNCdfu6VL2Xuj0Xus09sBU1FazgW
XpQHuw7XcozHRlnUFKPJg2P12yPJsLRkOqUWtHTUXmH/8s2RglOoEcmFeX9FVh1IRMdnp+D/F4GX
/80OwH0Jtm4eUDa5EFkNoIfhlOG4JOG/JCsYRnsAoZAbyHMEk6qPxdOGDrYzkbA3CMCikTuE6wOm
0j69ZgENzpWR5aludQDu44oKZqgkdMKNm6Mvk//s2aUOTBYWabbSKe/I/+cEp1tWS7+9AAmaVwO+
KwmsZsNR4Ztb6OH4hCq0936o+bycwR0b+Wr1VA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4df1QYXbx3PmA5i1scwSy/ZAJgZ0wNtl21eeCeUI5h4IQD2UalJOUkc5a5UR/j7lX9ToyF2yFHzK
L4EoH+xXm54bGihfoaTvocQQsWhCDObbmBOtqB6WS1/bog7FNgoEObi/E19vJsjPSd6nCCdhglZ1
j33mJRkZed+lVziTR/s=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Rtu5N6w0tnewss9ZQUyM3gMzu1D5Ba/+qJO2rdGgk0QN5Nm+4TaVyiEXzVM5DP8z3mycaRD+z4HG
QXarW6RH4GHKahoLlSY8cryjSJRWS6D7/Z1joY2fgJb8apydMguGWjRZ/uW6R7BEimGxB3Xuon63
ZdpcvKZmoyvfg0kjAjor/DxtP3SP6DKxH3BeegGQKpP/+5EmCrAhhPu+NA21340wcbghotvyYusJ
ErSZhtj+1FLwV2sO7TUt1etBG8nf/yETDQPE7Q+zX+BzOktmY3tIKds/9qdyDt6Qb5WIxLMyaMa3
eyi0SGAuZdeDtK8Os3w2ajEZI+VjufruVqtCCw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17760)
`protect data_block
cGLfFxlv2Lp+HR2FHlxMDn2S8l/DwxcDWalUAnd05f9BKBWt4wTEiisBex1HaHwCGavQ0CSiKNly
58HtSMx/B66pbmmP50FCcN2hlTb3NyJ/YCsXIyom06Wh1z79WUr9alb0Loaj7ZhnjgU/pohtlXO/
O3x6t1wtbSybBMkGESwtd66Vld09Dg6AVz/Ahzn/jEcAJpmtihovJfjd0F0varXsZSLFatCBK3xr
7HzwtULLE0dx4d+JpqoXaK2TH7uvK5KbINUUYuAULXgylS2VFY1EftxuzJyVg90QaZUZEyswmDYn
AyiULrxXlnIvOXs/tD//z4IsXPTJJmB5Zy4coYtaElMNPqpsIKrCjgtvRfAhLt8JWoekl7cKq9/V
dV3yKSMnnwkmbo6XaI68fFeuQHXMYn7X1zZT9SogxjHTvADmidHFZ9+OlUf8HlwTv6rT/jGDe5P+
+SyBZ1muMt1Lla8CJnBai2Qh7uCDsvwxFs+sL1S9ABmdzLcYZ2jOvqICN2BvxJ8ljLoUfP3wjFCz
u9P97/wLkQPFORDgsVUym7TpAet+HM7bZz2NcREy8Wa0rojCXAvPBOkguWkaf1XV8pN1KneabTW9
pDVr3vdzUABP170GQ40kdh5ZwT5WuH56ezxsWTpl7U046qxdUX42w6Sz/5EQobvzCP11e/paCpGF
c0/QOXGl8CHKwLkvv7yTsbNI2Tc6sa4EAcDVmtMFJ1Dm+Cu1UmU/09MXc/GKWtaXg/85hR65BmSE
qur1ZYqwE6P0u8ofKzldM3WKPZSWwJzicH8ZbFqI8w50bBuMiNNi5ym55RTo8d/fi8Rte6sd0Ctr
jkSJIG6us2bqhzN1p+b6txKGmZNDfsCADNUkzm7+YeFir3XkCdRiN6yBiAeBiNsR0vH0Ol+7GRLJ
UnustppT9inqvZl6XIyNGZB8dRsUmE7QYmZ8ov+eTiiCyQ8pezXln6hdU5u4km/IsAUY9MUOcyw/
zzgSZmw71AWmRgPx+1f77vka6k+zDcpYfGCN+q+1t9iLN9VCQmwZPwYbWBZxTpj1+HeGLFrvS3BX
H3FoldzonOngAXfhexz9zNGCAGWwjH7QEfFUKbfBrM4F6W2l2q54GxAQNRDayVknsu1jpMv4f0Tm
HHAGKb89jt2BCklzCoemr2rEYi648DAdwVpeTBolDNlaks5avmtHK2S+Mm3nPLlgZUtjNhb9vI08
USrmYJoqxbyWdodbBNZo+HxsIFwhXC7Zfi1EnBZaj6yLnSQG2FdwLHXkENX+XcGWhIvSeDPPBsHk
GmgzebZuz96VQB/AIs5bfqVk5M3xYSSJGWVSaeeYMwOBkj9ZNZqrh0ppLJOfVie8q3M8FF9vbqUM
rpZiI/o71vtvuc7PqtDSxinNfNQpl/mWMTW8IxlzLTfxk98cfKvDtK+ngN2FmfBPKB1y4nZZvuUJ
TnrQZ0RVsYJXM2JScjF+Mz5/wM5GwIgQPmhoapQiC0sP8MFZI7SHckvndXEgeXFF7J2XAjuJugQa
e7mRL0ImDYd7hHOQ9OEPEKYBpCZDJWkMKb5F3fjTg0wT9xrSTkO4f2CACfEk00XM9s7NU76/pWt3
b40XzybY8snKA8ieCBK/tp25/kVsIt+VgMax3wdL83yrulNrWW4tzQauQJzkmSib6N5BypIDLHD5
yLkUumcKWonSHysX9WLc1K6whLEUUb5BrvH1DjftoE4Pvl23Toj9sdnU7MXlI2CNTCOEdX5+Zqvp
tjK05D47KOB6KY7X8pspNm25gTgA5FDAhai4QJWmdjP+Y38QBz1HaZoNBVil0pOXwcsDbTk987Zl
cyTqOI0ZPl2AEN583OomVzIAsaNX3Y6uM5vA1RLPCQzZoZliBI2+2jtHcod58rNPdhDlWIRo7ZQ9
DBxuOdiMuGe/1EHvkJa6ShG7R8PPru6oVCrCQwZ8j4LNBt6EcqOOaXlWUGhEN+6x+1TeGklMdYIN
7XUFFOLg7tl94XJGMwlZVvbJW39/BPEBasKx3vG9ZV5kzMJE65nAwzsH5OolDtN99oCCmQ8O6uTk
a3DoEDLthx3EOYyNVzSTG4OkE+IXrezUz8bt86Z3P0MUqIGHc4Qe4CEkYP3qc9FbO5xo6pMe+GLj
MaxL4fne7Dpuh+FM7W7CJkM1K6GT6QyW9GVDLn03bWlPDB5EVxh6FxNwQc6c0WtX73woK2FUVTfj
ZPzC4BUxgNrr85gT04UzCw3N979P1357pAgkKVEdB2CbdfC31d8dP1kLgv4A+WioKQFza5EgnEze
xIf9CQcA3QVdtriJVRVb1RXVTHod4fDqpCYeR/LCx0tQkpALC2GT9LdTMgIyRJztLC6dbENoNMyb
YeoPp8W9VlCKxm+jvK5bkj1yl/GrkGcTZ75zUmBKsqw5TyfoKqoUcq7JqxnRrxTewuAfxOtv3RBp
EJjk0OisH4YrWUasT5Je5X2+jmeUXa/8eUntFHqut8eUYvPwt62w2lyizl5uHCig1XnIwGSE2q/z
Jes1/8b5qqtK/I4Luy+z+NhIOPWIXLn1KebBlrl4f01aImj7jYMWS5m4kdSgthOt9jft0esenX5B
ChcOYnZkC2oewkNdqXCsmswIwPGChwobml3hZDe0kZqi4U4EvUfmqG+rqyq4hMP57zrtIxwIrrlf
cUxq33bQdIzoHIYr5wJqSlETevTU4XCcEFs1mqWvu9LC6dd1Dm8ECDiPjW0xsUf4RwHHoyX39hhy
//RateA2bwW2oDhes1EzQnkCfuX4HJi5pLj0+gzhZlRJiFi135B6rLyGirQW+rKMIbsvkmqbi6Pw
7NiG+Dy/79XXr2SXZspEGtD58MNZpeWal+y3QA39TYDqa/vDlA46UjvevJN040/f3o3gs8rO3xuA
zPdDHe0dFHrKwHWkiAnquindfAKXPloKzOFCPUJnabelMbMbkHYu0rCFmIo8foHxhWOeyEhD+gH/
tCSw967gW8JJZRG7eL511frK6CL/9QjRD6r5MbzCl+SInAApDPyeAXs4Lppul11rfAdQ4itmxR+b
doY/CmDmkEmeIyDoXFKE8XnaPd/pKUa6YWiC0+FhjZ9/AvpGlDXLlaHiRpYOOC2M5/7fT782cbpN
TPXw75hCkK2SOWO3PVs2BWhOMDFr1FGLd4b9HAZrKuj7jgaZ/y/BSEVmRYykYZ+d2NDPEHlheIMv
m0yY7hSeA3q+6bpbxCqNBCq338AT2ORyvX6zly6DsSNZkZ1VxHGP6Qy0N1rT27M93Q05WJTZlgcn
5FkX/AzCgbsMIQx85v3Qa/bmSKrG+wX/CtAgeHWOjBHHmyftR0MHt5F4mq6bo/GSll8jJBraIp6n
7kgSVU59FACj5A0IYvIvOpH1KEoHtVPQf+czYS4Arx2kgTjmzSh4JgjV53i5pC+5pRCp8aJ4CLg1
Ld/PXM08BE9eri1pQaq70eTpJXyru8GnWnx5KHXv34y1nNWodNQOCSG+Ks+QpEUnQR30TRkrtymQ
pydFbY6JVCAD78ZuilJaLuca4AtCqZpvjU2u/RrDG7DgSIf112NjHY4Pg3xMT0d6BgJjhfZmM8Ax
AwfxQ4AEJOw0wbWc1FbBysitnftTNVjAKd62GcnKDDlalbWCEbJic5cK7iZ6WWXv3uqFfIVmFB13
yYJivTh0sCxjAsrwdd1L50fWTdoTs6lyeKuIBM32kW9YVkIDccasAamYIjb9EuyQ2g0On9lMBXYP
DNAq1YN2h7aAox9z/3NkiqKce0RB1jwPrm0CLWI/TWFtE3Wo49HbG+Whh6UcWv4M/bY3A366U2wC
aNm5dAzqMPr/dcXmls2sF5H+UdedNG+6Z8SeyQoWcZwmbIMrMeQmfEVpDo2EeTZAsp4hNyWAGTk9
qUoH1OgxZyyBeCPTeXOkClRf2MmfQ0H39VH0nPXK1oCD4l45irOkWmR94CXRz9dUhdC3OYKBlh6/
4IwLuJAaF59PaY6JVx5TLkAcUpG15eYw3re231CrOTPGow3MCuJ+H+9zMzAXi9VOv+z3ldF+k/4d
QqAXPjcUTGjsjFJ5ZVahOIhNm0WSs/ngQUYCGP0IwCc+japL/APKjhDkrENMbJ00cmP5LGiG1bwR
OZok9Exmyl2Zc4Cs/r2imNly8WMBBhGDhHONZ3xcyPWGE+IhfK7fMK2AckPdZnBhV6ZtlP811VTd
BQU/8Fxf3ahErxGK7qxXjVIg9uKxuiFIQVMDl0cjhdEItYWUa9+RYmBg1fP+cKGF2e8hYE6dMaY+
Ds/aVQIyfnKyPw+ekTGUSbjAP5nZeiNfVgGr31zT+3Co31LWG+HHq4Guf7T6TZY8A9lPCJ6P1KbY
gIA8+uRLqN/grVnhVnLeIhq2CUT6buj6at7VIu1ollBgwOK6umtDaxS7FKTJMFK4zP/+gmeCFybj
F9JA/XfeSBTOzrq/AdQzx2LkitZoPJUTxF4jy13DEQUrS259qh9Jf3aGkks6uMVBKTk3UqWU0pKK
fsy5hw6fLRKHmDpoCydvR6l1g62uSV6fqMBEEgQvs9W/rM8V1uYKw2jRj1ELYcQg7orlVbNtEdCR
uh0wAhRM9KWJKozuwXWJzeeZbpfqku9J5AvJFYdz9lRS/czp6/rJJhcbyEfZp2jRQXy7SmUj3egF
9R71p7uFjHhJnIqiECqKj/xjxNsULjxJpN3aMosWDEoDwKKfKIoh+eGV13UYdtipWUk1U/8ZlXBL
+d8A21Nqpw7hz8iOCkkMaklXswSvyuZ5s3eC5COwa5xbOJG8GeL/5rVPoTQd36dkZrE8awbvNTPT
nzh0zD9DlbVuy6ajjZXiGWsJxcnB2MMwZP1a9sLl8elKV3zcdtsZwomDNy6qrVCrURxxgp4JnGXQ
hSwX2qowT32EJ+MuemJbO+1NO3IBYn4ydhQpDuhJIFmYvtmcbr8bqZMoZdKgz4F4SaHxdhSLNa4J
UBOXZOUDnJbqjrSrFIvDw/ebU3Yb2llmPMT1voi/kAjH9seq/hF7Xu8cv+d/zje6DX3fu2bvfHpx
fJlNePeKZl8e5EL0TZJmbHRB206SNHaWPx1Dc9Z2cy3BNDmmVImV4/O3TWRvtppJwdXk9lIgCJ7c
peFgqQmPK8SjVonqnA82DLNxwsqkwdol7RyaXyOUKDJ7hYXzyXv/rIeqNxaYa2NoWedo+n6LVHot
uTyq9Qf0IjdMxcGs56yY8GTowl1r1dNr4cnIoQ3Y83eGvQjZ9iHRWF4NrmVBQyTvVZ32PCmVEu2g
LF7KB6wZjLjRjdiKRpMnrHRZvjZYUM3KWud0YhsFY2erMU6Q4SUY/STpWhwVFIJf+3VraSJektBy
pKnzzoXYVVMU/0iFiIx9KbW+OQrrXDd9xdwCzcK2l1+m82AXnhdESmDeMX1WaSFsKP1IUK63MlWs
Zt5B9ZD2RnOG5Gx5bLi+mTkGAW5H9CWlGYQP7pudeKspZr+vDF/w7zfO4X8J5867oKcd0GXrXVq4
VQ9UWB4lgQ8kq4KNmLr3Iy+mW8Ra+fFDae9/jz5+FsI2hrUtvj2A04lBhupXVdiyjvFWHCVSy7f4
okUIJmzA1+0udNuJHTx17ZkeqlHBwMH9XN25NsEC4Z3cJxTPdIPjj4byRd3yzTU3qakPNVAHpIS3
yl9jjYLE+aswemx2O2ISrM4chb3W/Bhb8yE6YoMGGZU9Da6zYbuf7czr92GB2S2CM4fDNkh+0j9b
qwuB6umugOhdpHBDrtGu7iAlPAO+ecNz9olu9gumZCN7jgiZNCJW6Sm9neC5yDgqZxuVYL/IlJkB
AtveLwaBZURsio2E0uAiXjsfKnHf0h1JuCAu+Swqcm1JB7+Bz/L6fp92iaK0hJXdwS3NOnyXeQaS
GGAet98oNkj7VJ3VngZw03JajY9AxATsUYU42KNeWA8olxDHhe6ukDPQvWbC2HxVzOY6FQ6yH46X
hW23oHIwvVFCfihBOiphp9tUuC0T59kjZF+01Xzz5oAjY0PKRIPQGTkv3F4cWnWjtQ1AAKfpBeyc
VzHU1EAhUcA7UeX6Z2WTFKMJXS1jPUspb4DLU84hsB0Ql8YOcHLCqfWdJhoWwTLxDXehY8Ho4vLE
6mssUiojX/QDLjdmYBBNPCbBnccjHlU3v6ML64uTn35lOaM3xlz5bfbBDoXx9cwedUxTtb27Erup
6SQA1ZKfLWJU9SK1p+b073jxZ9Br44YLVGByD0U7QUz9JYbFke51Gkja6Rqa2jw2cfNSuFhcpffh
tA7Kc69ivl5NpT1wPv12EuhZrBpqNoGiYOvsgWPfR0yKFTriAyaQeaKzT3Fc0xVEjQJFytxiUfXo
DzkXGB7CC1CTSok7JuTgJtiH6YOrSBzrFXEUy5Z19mrGnDFOSOB2ffQpPpIkzS37XQoJpTrKKL4I
aRBD1owuIPk8FjJIqVSuZzeQZXsSMVeGSxbguqhRSG0OVQ21TQKDbl91s0zszxZEdVIn5iA/fe/e
ZUs9Hp2R6sPJkrIQJmGSpooVnNP0qkp+9dbFqXhXFLwkcJ5kxLEBSOKw1Nst8+NQC9MnUtJV52x5
QpLdPSYXy+h6TVXBJcvx8wE8IyXBOydsKefRzU4GnPrgtYaoZWvLCFi8pULEvkR7AsTpanaBy0MA
AadKj8VJ12RP0PAPcuvSzT1I6TW+lR0JLhyV4ztCEfPqIUtR3iey6gaXLzw3OZnZ9E4LHiaRAanS
Xmk5hRGzVjwgbMn2HoDDPgL4RYmDFhCeqGvFDvorJd+4rzQYKQwrUAsjU0YydLuVAPDjQ73WjfsE
4FIUw3FLtoNZqffyy0E34B3Y4YPJdZ2jlxvT08Gvz7Z7aNufmEoCCMB4KxF13C7ZLNbWZ0o/GLqL
bM+PkuaMSBuAwkprLMtCE/N5M4Hb5S5hgXCnnPSsRfPsAsnp9Pbt28Kv7DhgiNe47H8zGO+CplmA
B09h0zoXSDwfwi6aWxxUf4upMKf0oqm/64OHDABooYxF4r32Q9YGFzBjoo0XM0y2Wus1A+4vNltt
ghWpWmxsNoq+RVDIbfz+nHx757vzo0R8zTakugAbBC75OQz+dLSQYMcfuDhmyVvTQbcQpipPwSV5
/QEPHnlTkswW+abtADFPBl9Mn2OwJBn8YKVcxW9e7OZkl02FuOLGqR5Jmg/rb/Doey1gh+2gphAA
1Ey2tWJChu8p0B2AClucS9cF9fNJiiBNCYv+gglS/7XzB1f30YGp5uTTKVNtcdNt9SsJKTKFt07f
G54xDRhRSLKlw+yPrQlhXJcsM+N95taaYZV0FnI/LfxOoK5YkbH72pY7XSt+0V5M/qtBcgMalrqE
N5PIgq/dE+H+iBO2HUZJAoY24SJ8emS8mFVtYoo8m8t/w++yLUDmhESyim8Bgnrd8NnXhLaOj9k0
iRwBUJiIXZjvJjmD8+1xALVEQGpAYUoVaaIEU+d2tuTycSk3KOlvAkdPQI+ocUxlMEIsVyL0CR5a
6rkGU/tQH4/bTal3i316ePCW2Kx5D3fMD+Avj0mm9OTCyTAXEsx93R6aJ0W3R7jV7Rw+FxK6Tv5Y
qd1I77k/BxVZxDAd8wboyDjo6OyTwHboL7ys+CFA6wc6sQEO41QX5lj7L9+mvfmgC7AjRzNveNAw
kucFGqHKBJ5TkksNKlajoXCb0L5D3ikauopjU1Xj++/eroLcM2JXscX4G1jXDic39OdeFyC/Ncxt
9fwf7KCBhTut7XF1UqVKGfTotGqtqnJ//Y1cE061rbGmNSGbwU2XQ8nBD4v4FOL+9+ntDLEzZq2f
44fYRhD0K5HAabZ5Y5F4um/7A57dJrzy/bnVS3HyhNp/G/FgkoYKgMrVCNmdmmz0rLkDHEFEaZdi
Wwtx1+6h3zKbGq5Zj7vefuhcrRlhnrLq/0weSqCoQiCMr9W1S0Xef2ulZvtXfM0eru4iHT4d1fH2
tBCgZKv3lE0FU21TgxFmqCX2qyL3ZF9V4KGKvKW1eVysyy7S9uffu6NODXX1UWuovS9QWG/HauoL
vPsIN2DZhMIikp0NePQqY9bvXYB06ijfO0GUHWy11Wu/5DCaPv63/KWKA2NjCqABQZ3J0AHlB06A
p1DaCW+0n8JRJfLae71ZDbLyejdEiv7uOYbQSf4jTGODskvtHl5yLLan47tXH82jaj7i1mQ9LhKM
M1fIKc09DgXri88uTPLU8U8eEAEDNApQEFYBcRNyLkXU2J8O6Axw8m0f1CFmyk01BgQ+hAkNdwvq
AA2wYBPLqJ3bX3C68O47av2baEcQ1V8i81G6VET9FcOrYiYJuE40nzOlQgZocmm8MiYrU1dmWvm0
sc1P5qVNUnLpcCHR8+WacE+d+17vkC49ph16/UMl+6sWu56qx6ZXawbD86rWPqH1+Zu3lZH6C6uT
wR7iUe6X9R/Ay9WNz+QxnaKzgnr0pFdevYXmU2KQL/GbeqOT/cz4vXwfsNg8xMpfiF3cNcP6K9sE
C7olzwyVYTHEDlScRhtBxNEYsAhD6Y8nOsavnMttNP5AlsLWt2KTWMkUbktpO8g3dNd0Jj+tGSEd
CFNDFkFUkg9nFBnQLzWrFF32xsUcn8t1LxBR9vnkqeuNPGpp/zpAjy/x6KR1plGHoOurpf5Hbm8T
CoazyQ+q7Nw8ILBxx5KSfXZzX9Rc7Iq/YmSpzdjM7S1Q+6CAmsB8hSPyjWPT6835FNNmBN6+jcBL
Mxo+U2+XRZt8RtPCNUazwFsmin4SdDxQlxEEViUW/oDSHaYMEYNWjiBdF0OrMVLer+UUAQtPIVRn
SBPo4vyaqQlI3aRcyQyiuf+c3Tua+QFLFrNiq+XYxeUWEBAOLVnz382PBRd5a6lTDEgxv08VHplB
38Mfrk6OeBs50kLyHZsVpTiJ00KFyOEbweKZoZFiOjqjm5K6QxIEtkJeyA+ElrLLWNlar6v8Kfgt
LR6alSGWVltXKUt7ctgDS6Jxs8tqxGkWssnyPNVp9scD1a5mP/hLTj+0LkcFsYQu+65ZJnBdsMYT
Fm+I1bgUSjAuu2KvXc60Ka6DIQuDhMf/9mALO8xk7YadXqNwURMYQcAVtZ3fEnr62IpigQocPUWs
KDHgek6Y2xeAg/wnzXjHsYOhzbuUlnKkejwBJmnZsm5Sh01yGQrI/HhmdEeb45VWA7KRqHIhGdDw
shfcO3HmZkseZrId3GJB9kD6AtX5notBFeoqUU/E1mr19IfEwlVmTQsKs5brD2rUm5gD8XJFjt4j
OvJMbTFnYwsF3GAHCaP7E+OW9IbYfpD2DLdkE8imOhgszylCNwCkqKjEyPEvKYNmM0s3CmTbmjiy
WQrEHIuBgGx62frkH/3yxDQ4RhmRFwlPwcDHSV5JtX5MqA6yGyQ5Nl9ppOmf222ESxWaDWRrJJ9m
JOUUhutPebzxcJRbU5PQxzKuwmAvrFWd3VYDu8wWnszdmQE7zZy57/qZW3I7EYArUpk7T9USge83
btd0Km7arqJWbPhm8MPIs62WYzd0Hr9cWVrTUfXLv9/P0PnWuA6FxtfR29EOShU/5vYlmykKZcfG
XrpVkEXbhNM3Pf6lx6Nbay7B1NusxjtBP7Zo6Ww+eiElcy2SS6nMUGedY9Af2Kyn9wtCCNPr172I
EACClIHbCmW/UEUe00P+UvqA6zicH01edvwKDGz3hWE50wu1JnTJkDx/mQ226r9edtFT7rFmYu63
Q0dpqu+tY6JhtQQqBmkeGBcZAtYja62wcnmw3hOTMN8D2d4yRM3W4O34nNOO/5bHLDnBiBrzdopX
WmZ4uBHGgU/8f8bBY3EiiCuOCIet2FThT/hgzRqlsuDeolTAGYOO7iyAFn6pLDggdChik3uFD0LP
6ptEaHLURtPfgRkojO21vcc0lBb9+1esBzunmQcRJGCOMjuaYdY35moWZ2+2OYqmehxjB6SKkyww
kZzff7Pg/qSpdmyCiF/GVlTdpF330+uhnocWp8hKYUYu07RUpLU7FWrC9sbvD/rVSCB7rBbfvbYG
9tGpHifYZXFyOf/W6dbGRkZwznuAG42hdr7oWwmYUgazQkIyVgsYHGYBYvBdfma2LgCJPh4zYwWx
Yxx+sma/bDu7Lr+CKpcVlEopZ7p9umL9bsZSo7jVluiwWXxMzmA2E7/coU/RXyTm2qQ5U/etGs8p
ZE9/M16VL7VM68j7vRgDJ1DcOnUVyg7LblZLNJJN7eAHkAkxddJ9DZ+eZcQppApFs0OuYFt/sofr
1DGPKi7CPhORjnIxmTN+rfyhzkN0oOGFb38ClxlOka75c0vu0bc248cCYYeQA677E/0V8V+lAOV0
YSlOj6NVu1nzbCqu99m03+8yO7VfepxPbIGe+2dL3dYZFILkzakJT4PKYSAoNB07bqswFRQqfFnY
Vxh9AtFWP/OSdbmFIfVIBEhgnms+NGgI74raV9hV1TfkBXrQ+j8ViNW5AIJmMecuCPLDEPBmG03j
94ualaPEF+b+VldA1lpoK4lmy+l6T5DzvhtjQp/JiLyUDFfvAKyTwIgbTRnDO9ReWE3vOhmIY8GR
cVHuoMrcorcDK7za1wTLbnIja8V5MXAX/SIXu/9O6KY6OiwsbJXuLg2z98N4suwm7aywv4Fos0hT
L0WChYacnU2T7ygPp6GXvOKJMhITC95RX2bMuSHUGzYRvBIcfytE3EZaWD1GLJkGwJWzMEQPWkq4
kg/qhP+6FTKo6qUshh1SBWdoFlmbH6OJeW+jv99yX57cikhaEHpfCimYbSYsrdrp8uoHNrY/cyFw
NLHjJ+bFxAHFXofI5QUB1aT8rx1t+emcWRHxj5JDawleigTWhGAVAi5JJjcVBJhz4yTFHt3UH8Wl
3276+uetfHyiFUmhZ31CFT+hchHyQHFdamnr1DY5lLy4T7zxpVyk8GpNfKTR5mB0KLJ3Ta85RiWl
LDPCw6Roq1uj7k0X9aCN0yG8wds28fedoCrzNlxLN+vqSsrt0elpI1GL9zQOH7m5SnB49uMy5eYE
iSp9Kk5/T+VHKhZUI0Zpn5U5Q8E/cBtAWds5UNiDdDTErNbxQ5VRv8s9HADNclc0TW4q/aKABGop
3dOIIkrATR0uKqjYEvV9FkYxnITmT62y+Y5w4qMo/egJvWiw5ybNTV9aSROe0iP95pVFH7WlwrR8
AKa1696ZEaPRhnwSUk6veeqFIvQmx4JhlY862C3aauJwbI3f0lVZe9ThV54bpYkiIjmN+7SstzZs
NOIZIyEqbK0aLLyNz4/x2jnFv3S5Agcfm6+1NxmN8H8pEhUqP9XypgX6LCNpm2a3pcmWTrsH7s3x
+ww+P4c5HXR6O7SYjkybiFg5HHCTAhcUeQu4ZXpOyBKFJ8WMy3JjR3vkVSQh0zwObHOc0Ssk4pw9
RSWi2+HK9mT0u0ryu5MRvwr+5HavL/iWmHPtJJ+1+ComOptgG9QaAzlJERuN0BOY9b+7BHNNtsLC
y6M5wDYwWQpWUNnHKxWYgKyEJG3aUDeG9YxbwYITYr/1ye7mr9Gh+rYA9MUGE7MEGRnPdrkfOuOZ
ZWJXY0EtW/9ZZ9mcIHi2TRKc7El9kFwSYw3pwrqG17FcxflbNWFhomwN/plRdIkiiSBme/mWkk08
LKx1lwSvmskPP54Wvv6NrnhMOhTE36DMHfkXyrSVOL7DdvAXPapcnhWFB+j8JgjWuOUhnM+ESGkA
+J0cKUqRbF0au2EufRySY05PGu7hRgLxUJDDCys3Xn4F7rawkvLYgDVI1fUJwJS+vNfADPdHcjdj
TstPLjdAxB/7Bg3vN9wAns7dIqONvxtraHHzwXsl3FKpieOxXtjS89P9kt3RaeW8OtCNp2GvzYjK
XKaBV06OoJEyHJ2NC59JFoVUXLg2aYJUmlqmY7c6vamV5+3JE1veWnD8YBZCcqgMs5bkgp1+keoD
q6WjmcP7D2drbbaB+Z5YBISUfCLOe2X/65Yks+Q6B5gbRjMFyKsvvCQalSeY0Z93gmYRFBrrlGVK
M4lnH9oZjm5QLJOYCzDCFwlAHL/j10g+V4B8N/8uoUd49k/j42vMk8kwW7S5CfLCUhfMmvrfNVfA
akyGsGdr+J93Tt5Gv4o+JszIhHNZXwh1jN/VBlO5uUXyNW3VoaRKCZ3OW7mRZAY/YPqOe5y0QOzv
k3NMx3hYhquOK5CJ/tS649SpSOEnheWUKJzc1vq91YkYnKjRsHTJwnGa8wbahI1oQEh0No0zUvA5
5ligN8uvFinSPtGuB3ncA3galVkqfRrVT1hyokrGW3x2x11UXq4SbxcOuQBVOzDkY4Xs/8078XkJ
sls4Lr617KwecxzuiMb2h+RzxR/zlw+9X/j3ezbxen3blPhpInSFnXZsYlmuBjgZNG5A11yNte3u
v7SWfpHDCealhdju89MX5IiqRuKOv24vHNuMyEWDQU42F+epkvOgtoQZ00mZ+bkKfjNNg5mHQT+T
RPM8gCp/03uxiPWEC1VLpAjuUgwm6rJfHBRRX8KbTas9C0LjajHmh/x0Osbta+Vs/Pq6weDM3P14
5xeWKCc+Y+OJrSrODmAVJ5LfXAiOTKRGoeZUxFxi63mVGvXhy08hjTD0hwou9Rlmz26NbrrsWVpB
3FgqLIP/gODvjHRMgjL98VsFLSQvwfr4BXGpw4depj34VCSQVvlw1yP1ZB1pFGtoW0bdy6Q/NP4Q
5hh0vqkmUQgufovIIAugMcNmwnRjfQnhdn5NE8kK3Rvu/682XOeF+Xs5xte4xtF10+Hc1m4LeJKL
MgQ0rcAVswc1/5mGozW/CuQ8kYoKBKySxbXLPt8wPQvXUFNn5XBczFQNA9MH2CVaPciLq390f4E5
HpAGBIo2bMosOyUOIissZK4YAM+UhfceOVoeFtFi57uivrA4t3N8un2JWBlKJlMUuBqravC8Ddmu
9QvtW6frjaBJarcf513+tfnLOU9XoVytZiW9bSiDIdJnFrWfsJ7SFlAj42hWQDDAtpChMiDo7HIH
KeV6GlubSVvgDumLYXxhn2GwTT9yYq7HtZf2OUix4UwtaL+uKKEdXAfaf3PBR0PhLWGodGov9n8j
kXLeed9Cfr71sqU9mOnO1zwt6+sjkNoxquGRWqejBqa1fjdpbQHodrfR0eBshPNHfXKeShO+TfiO
5P5OQqWOozopXXe85DRijgGJvemgqHdXb+qLESxmrf9nlTaNcUQpT8WMa0nN+E3RUsm+NMImcakU
M2F4BA7g8xWyMYdF/Etryb5PoVeSXT2Qhs15JhAkeAFcaTcnL/Y2Of7lG+uEgJ92PVVi1/AHvucL
cAPryCkGmBWI5ZtaXkiYieyYnOvenRL1KVBUULEav32H2vuzq436NEL7lEVBBAgL2xQiF1LnpAzz
38gACkNzC18awFV/c9iK6LCXB//WHDqP0+bO7T2tE7ckI3kI84ajYcce5gNlGCdrXWQBNAuep7fL
etRqnGrQ/E7IFbTG8mknUduY/65magPCRNUEX/8e9kYgxJYhmxsSdmfonkY9/wdVQdNb2XioBwu+
mkve4Rw3c42Ve58BasVuPUnPyizCaiVeatXD8IOuAAAnFBuqh7wZfQJYVwpfmIkh8xKE8Eb39Sja
rBRGUApCbzT5SC3zrdYD2E5kvT3uNxQLutM/l/KIyPtd7ZQLVn7LhFSKSieE0eCyajFUFGogyb43
nFuRsCrehI0orDBL9OV6+0jLWzcmPE5kI/kzT9IprTvrud7J6wkBR4cZ+QlVZNvZWOgluBZFqZid
MZbdTmSNL73iAfeCC1+k3IQuVlFKrPrFkDnvq0eVvEvZ4fb8QuZmB2XA/7n+bneSPyO8LKbj3I29
lAQ8L9zte9xKChalvvnkER9rSk3BTOxoTbgBa5C6FGRTHpjLI35gkAk0ndPN5tli8IJLH9rdWnan
Eb8ABBeoW4DBuP0D1VJl5j5085GvczAlGIybKL6GS8VfgSQXHWD4I0FlgOa8VfyR1WKWkuF0rhvr
3X5q2Ih+fEMMo38idpacG/U3OqGvWOrB9uktFo+5zigfdY6Hk26nhWf//LCuYB7YCv99syJV0BW/
/rQozOodtJ7x5qZScNgkLWwzsslJggoilxYh17b5jVnL4F4LkoR4JifZ/byvu233CY44rtotj9wC
yBf1VChx53MQezK3HjGFnCcPggXK74JL4C3vnjgoLCgNL9Zo+0dTmK0FUyZvKTmvqNEyb3aB7E84
1VsokklXx5xhQ6DyW7kyPdrpsrMUOxLVgPCrvorzgAhM23B0w/JExm1Vv0KhTHXD4KmpPeFoTavk
g8UDFxn4/alJWwkrABN9rPciG0OJkYa86XVK4J7JrqSteEKTfAW4z8hL861X9IeFMcSjIOJ7vGm1
JmLvzlMICyfYNWeGxpcMiyLpwNwv0L2Ff1m0AazO52GLW5EDp7gfInydNGavzqtjOsnCQ+rGeIav
MAbFTxmLgLaAtFs1OTg+slVHGrkngKSIZwvc05JNVP2wLBTvTHJap9Z3RrxXTXq/1Cizxfr8QW37
sd5AS+F5kG/b2ecv+4Xiv3MitIc9V86RRIvwXpWbzpe5IjOlrafqXkhL9Eht7WMD8aSYQ8sO5107
hKiooTbRTJZcFTcWKMAxGyGyGNJ9pzhE/pP8iqJ20RsBhAx606/Zo0753dikCtm0cD3a0Ed2n9Cm
pgL+v8n/Aozsw8/7YQc04H6d3c7JGi3vvx1m96/MrdNxARbWbA0eCMQb4BI2QVXYU3ynrREdBUyN
xw5vH9MhswR+dfvtFs9tDD+VhBeM/Jr44mODA/1s3nGG4EaAexbGSmI1L3qHxwr/yWgs/mI+IGvK
eAqVMo0dwQ3I7hqcotoKwHfWqIir1MnfSH/FuNSEZ+bK3hKRCbCbwdt5dvMBlha7CGA7YzO+0V5Y
AhG2UYnN3yFlvd5uQe2GEp/JdJMovPEUGwNvxNT/jKCEguOL39wPJwORSOC7/U2lgiqSzLJrk0nR
KLPuynPE2WZNGEAcLiQIGeXuJ1GvOyYJJ1qLdsvU87YFlShFEXhO/0/MEN00KdnEi2c0M8uWFvJR
BPZINnBfq4eOXZbJsEEUXgrP5ziYpy1EzuLZ3qO3y77/nEWvmygQsbB5vW+GufVlKhi0v25W9/ZB
mvvyBPAq48Wm6iDLOzdsu271TxQE3fNOCayRFs8wg5Zps7gOTJGuLf9XOM5gUirM2OdBFv1LIQ2F
uBSXb1/soFfbXfMSoXTY++JIoUgGgkr7HQMDeoORr54ATwYkuR5BUMBFku4Ja4pK9m+b7dDP2NB4
t/e1Gf1ZuiVnXhl2NuR0zfzY+Sl7SnA4rhCiQJyaZfPPZxpJpa5G/WoljalNHVDoPN/ZwR/A7Mmt
RU2EwjU+JjiIoqN6exxltO/5ro7smd9hJP6tdNkiLNIPOXFkzxkKwzAX+ZRc6zIGdskPx9mPwU2f
ml3h2V803e6bQEhCYzc3mcfRc7Xl84+kBMNmcJRpUbDE+EA1k1HQK+4PaY4zEVRbrPi52+65nPwV
EN6S5SIE88rI2PDJwJ9H9w0apWPwGNYq5Pn1C9PrU5AkW5Ej4sQXj3WBbaBE/exQNTGLVFw+HFoc
ww+V5OqWi4g+ZT2FSenpRZJFaMbctwjQLzWaib+VCzJPWVTz4WjivbGosekUNDwr2XjPzDZ7GEJU
VyuZhGWABnZSoCb3qLcoyns4KL5E4Gs/OnTeSocKualdbep5xYKCGpyoRuiWdb2X2r3QcT5VYJhP
YlW6X58z4rCbQnia0fiH4YQxsLrJQn56ECQ0D/OwcFPfR1OF1CxynY7Cvgki6iq/+MgdLb9zBEQ0
Z2+iFkgyLMvvJ7wdtQu8pX12PesGihB7uhqxdtgigrJTjYU8lWAmhNtjo8W//zsmx8I4+l1WA4se
QVP6MuSzOmVsm4jyiyGAZmIzR0dweDTVTE8bHn6KCw1n3ahlvmYSB7m4sfMCrVsVrGCm8TribyNP
kqnx3ylL5DPiB6WbScFBaYa1CzmAkcEbc4sBx8L9xUJ6y+hQn/PuKYh7gYOzTYS5XmVVxXWZm+9s
vDVwVfjc3bvSNDpArO4xLvkY1sKPQQe2JUrBlEuGGbOd0jyTMuMUEQ7CPJV7Sogw43rNZz6TMUy4
/YXKmkhms8cUcYCKc0tRiSYaP73//XF4ehCpMLpFGygA35nTssH1kC9cEw9GMSwHtvx+8P7j94Pp
ByGG89bazGEgt5ojNsZTe46+mUsiZXI8h6GKxH54sbLkYe3tTzALCoxJL0Aszo/5l2DxixD5tTLm
SIh6bSEavcdpklZ/cguFn29Lstht8J7GM8oWQCHCb3PVfbGBoX8mSUpE9GTnha/L/xosj/8H9R4q
eQyKSfNXfDvy+hoKC26R6sAS45DmpbuyLtHy8ub4Ukwipp82hYgfAAd+zndWLkieC3c8VtufpSPL
CJhn3I6WZLwqTt/L1WSzuV1/FoyVlbvEHfwLQbS5Bq1Y7//2CfGUvFmoQtgARQMO8ZtlkILy4fcO
8nf+oKCOFAsJiVGMODx2fJQ7idMPU+R7goeDXf1/fQFwOAxO2YPhnZ+LNYHjUu3Qs75L3RwMj2mM
1xWfuNk++4jxthqPUxOv9tNZTz1WP7EZpELrqfzkV5RZeeMUJH5PdKjfuuDYws5mZZ5Z/dW0heVH
PTKv6xOuSnZGAIssEB4HsrApMmhTRo3YHU+CXDTjREkqrZz8TdgV272wcS6S/Jyapbn2vij8zeEm
61TYeg78PxHLq/fDd2r5lShZrGYwn/LfmbUuNXYwEbAqFGm7QyTMq3ma+tfkXl6hTQ9r1jyijhEo
nsd0GGc4TGsh6R3s2AYzMDGK2dg2omZ7pjnlSzEdGRXTkOcBS9Wb99MP13A4+71eWgxCC5+64I0V
0nb8BrxWglYNC+/jF7R2R30Y4NFTR+dxq5BS8necsDRRxRw/5Cey2E3e/wgE7Q+mWmymQY1eX5eL
RCQtTFJUKr5mUtAojdvBkGNU+XBDUe6y/otvzB+fP+xXcM2BzROpII5YLu0tLm1HyARzfnhQjn16
vInBCOV5Q1OhJFjoJ2wWkNHwPJcx+mwHhahKznFaNuveBuL/thVlmEep7MFCUe2+by9BHo0EWZwS
RLmcvWXmF6Y6VhYnGkvzDKYauA0IkQvNGWWsAydOvOUWhZIDfDnqZdipUdGpIenIARvVJtDDysor
cbSgBp3ThWR9sdRS5YgqPL03fyfvzuJvjZFVZEpxw2ugecWaV5qPXhWxjiIZxX9aPsczDdeqMXC+
RnGR6ErjVIXq5pAi/KiuJhKZm8+wfICxfalhbFN4Gdi/HumSzqgzJ6kwHTF2KpgHlczXQHM0i2Rc
AJE6M1Tke45qKBn9nGMuqPxsJS1gu1UX0aoJlPzUyLE5BvYkzO5Exl1GcsWy5FJ79RSHXGnnBKbc
0ODAhSyn2PyVsP+MeS/WX/P+ZAz6X/Q4DAI/6n1Qh8vUcOP2cLxWUp3UfM2Ep3mGu+9Eq38nv7vG
gk0XNn48ScXeJAyr4UkzDlDadUxRTekxSTdIwoMLZaur/AhO+MIOXE4o8P0C0SoXkfMSJ/dk0oNi
Fyqmy5+xkcBfxffCRLkCAhjukftXXlT2ZZCGRoSj8Q5mKPaSRs7LDvkTpw2dfmCalOiyN7j0xHHm
S6nT+9uTVELH1Og+WT93Y72i3zGea8mEInW8ofarnShxQL0hOTJ0+Xw1dEXK0sV2BWbVsS95bW4b
rzRlytnvAbJdyeG9JT/IL06f0aHa85Pi84VzqPaaeEWqLn+uvxgGXNTF1tiUS98tb7gMlZHgSlMR
WQ4TP5iXd+UH+oF6aKN/FKBUx1BXFQj4WXvYxj2mx3ozHPFIkEPy2r2qIGIY3nqsgct8ou3dfy8x
x0meWDedsfIDAsEPcf5zVbEyn5dJiZS9ZLNewPvBIiIDoHLm5MfTpxWQ6oYIYzrBThTISVUebeOy
sc7SkHqTmWbchWZa5Zh/ZsWnxsWTDyaXozFYmKQTY8z5XDdwg4vD8gdgb245gqydUH3AcV1pSIi1
D/YEBlwlE5+7oIZ/LoEnUR7qFuqXHRgi5ZAAgjSOOl+lfo5hyAutujAbCUGyrN3tjF9Y/IdW3a+c
nkC1qiO1VDa3brr6Fnx6hT8qA9vBaUBDV95haU+vpOLLBU/SPMjA5EKdyHTKUtzp9X5WF/3DTFns
dblXIBByIlLbY0cetDRogZvJC7Q13oO1EDMwKJc4sVvXScDudbcNUoBk3Ueh+zTvxZxWQSA9/H+3
2UM1jL4nSkYI8Mz287siiiz7WpO4Vib22Rl4JSaT5wJ7SV1AGnV8mJ7VVXYOMZFA+0VyK4Ckzhiz
1xhbUY6gaCKdz4K4Echhyx9rrumulxN+XILcxmsZ79t9RaEcSUpofySDCjURWTb1nUK6GCC13IyK
1D/kysKViwzEFC8ORu2TdVmZhK1npSWwjiAON+ROovLZKsEXlis4tIC9bbYrt0ds/MmEZVM5BpMo
RZKq3lFI6I9GyhxKiiiBHi5ppu6ycXzRw90C2za4PjVi5V4EohQ1R2nmlo/h4tJ7y3eFjewOYl/6
CrAeespvXvmgzW4sIJbCjYqFHkMstSCIGOLgvZh6kvXvC9x/SPbh5pVtshjRlHLeHi3kp5Ak16GN
JR3lfi6UQlMOGz6cM6nESCNujHsm8AyJcz+qg5xz2ttPz6Yn6KNdw3pTdKldLFQT5PUcWUH/mc/z
Q0joWwztLAnBXtC+rdMeupg1NtXgpxrcHGkp13wEUqiQOXMDss0Xv6GTmBeoEFlcDYgkjA2HM2XC
OwbMuMTH+qvYsL0ZddTTeQd77XBWVNKPkuKi2ZpC2tnkzcCZSllhPf66bUKlxV1JVN8yFxRzCrYU
62fkdKafbUVGTXVA/85gy96q2BeV9/uToujG0TsOpnKKO5SmJBXfLVgSC7VZ2AwgAJr8QV754m+G
+iMtAA36csj7dN4tyJ7fKm/ul+B9Bv4Lgf9icKmU/vLyunhX7LPyr739cTL/ji7HkeUREbeFmwMm
1vE5XhVUAxqM53zZVCjwUCFQdUmsNZ8S/0ukt61XAkI0O7BuPOjrl3PdWC+TbBuOK7iJMnNO4xcN
7gyq/nbOkq5riMgTq79KS0BHAaBAmYWLsvUXXeIzUBzHKacRPuFiRF3CaziihilHDxlqEn+LPzAG
HaLK2klUKA8L7AjHexa/iLAyEXYBqZsJrx61cHfAkCILogcpvJwJi2IC3DYfuzRBgRjygge45Glh
sI7pbvWJy4KCsxDQZsI1T2tGBeBynXNdvhWgsRBxW/IEqXdeP0ME8J1FOSKTj2BpWdQYtpnI+s4y
fAj84oxxgKUB1l9ELLlbS/ZSms/P7HJiTj8UOgb5Q65dizc5Z1tlxtbah87qGx/tIYH3XMeuhaG1
kEFqkJWN0SxMAIsbJ7A7Wt9QG/FF3puFBI2sq9kmrv24NjwkevTfd9uYB1Xy3E3ZAg5RQR/cuj6z
IVnzvO8GLhUrLswX7MvkjcNI/us+OBz7DSsne4/5Y0fzhVY57HVwi6nZQeEQ1VdKzT5rzGwk6LLq
aaiMoIhLv1t2YKv9iEkJGfX4Mhg5ib6SAVNRj77sAbtedFVMerOap41yIGSDW5C7xwdidwJE3Iwd
Pj8pw11jhFrT6m1pAxXs+gyIG0CYLG6ui8GpTWz9autXo/1dVtsfbjQbguUKby8gZblS+bYalsUW
v5ttfUkN/RAWQJIcxxqdH5oWg3vniQKCnFRrbxpk83IFazw0DCcTTtKD+vc2n7KploQqiAir9GMd
jEyVrxBlVe4zXUEisSm/7JC/4+ubNct1x0BKpDHt7xV/PecE0UdDSl30rTVoz/XOtRtCh89ddclO
Bfyoi6nQP1RUZTncXIjy1Eqzy9QOjnYET9ZB5A5JbGiUY7fdT2XhblbNsmv90fAwFRAg86dZtIkY
EgZoeTqK/W3ivhZBhAPf04D4GDdOukoGRAsuPA15ejBjn9LfafnbyLal5D/AptnzSZ6J/83bDw7V
5/4/wF7jCEgXvvnvDNPKuhH1KOlhuCg+uGQtgM6O+YTjprsuI86ppptSx71Mz9qnRnn/o+Jl7K4C
RNA/j6m0n5aj+hZac0C1vI9K06BDJrB74NlAYZJQIj9VS5Y/DYnI3+Gfht6sRZQahQmQaqDUBS5B
C7ds7LKpHjFY3S32SkhgVa0n7KtIoujSu1QRnZD7bExd1MtaZgeigEIn+vQOVEeLzr/um2FRELeQ
qUW5NNxA60FEgw8U+pRXo7feCRDAJjadpUL3CPrwDhsbCVCmP+wkgdJuQo8ORnR4mNWEum8FzNYi
TdTOanqBFPoS9xhGBXCslfs9Bve+pIqaDJDue8DlF9rItJ2f8r29kkx5gj9upbfY6RDsRFvwkWx/
6urtP0tVBZ3ghAz9vrTTx/zek23g8azhwuwVImHAHMjAA3eNTnp3QQ2x4PrRmn+TyTB7VyKmUyg6
mA7lW3avigtDTll3ZaesGBIqAB2/A+YG780nbraj05xEP4II0woteD3/Z/QQr9O/MjHM8lWg7+ai
dThQkm6gtqjOn8A/47SoF7kaeOjoIojiiDcRSgGOrNEHKLpypa+bwzI9LyWpirnSdhi5E7qkC7/A
H8cgmiVr3/5QppxHUvvIPBImcxUNMZznYgeE747S4lMfhUHaoXUnvGQL9yUnuYZI1Dw4URuij8gJ
KUg3Q7lvzuzEEoTzrrnAXhsZyZEr53mcgAqKGC6fb9/EmLD5HeIXx+Rgg+zHNmVqU2crR+Ccd9BS
1hgEreHCIZl0hsuKoygVTvY7LVq2fthm0B/h8HtNu5JuUdfKRr6FcLzR2jQOj3EinxRv0nck2rUY
u5XkAVZwwAQEap0NdvANGTkfL8sF6Me8gv4CuvdCcvH5lpa/ruVkD6ZtHnhVIC0bJy1NguwpK5pQ
NOpm9vhbuDd6jWhpmSAT1WlEU0P+BLjIa/ECHGEc+ND3hIezckGshb5OTP+Qd/QJwvLpXvpXdVge
gcE0lgdjpTKJMMxCDFkgcxSJ0Q4G3JlKH8/r0vlmrX8mjeofEs6Gjq8shtITwf55sLF2STuTZhOL
V2VBKzlpp/Ec9nm5yW8vZdskdROC6RPnzcqXU/Ue51IHAzzxvN87eJtdq3PlqOSF7ao2ZV9VhYZV
UiZRiwEyPqpQdc7W4V76G+XadNw/dOr7ACtfcrqz77+CMNAY11vWDxJm97MIDbwZ4IFEE0dqNbAw
TsJcTMLrzZFND7z8KYggiTylsxbBsguDuK41wLZoZOc23fgzZzBqXNvlpU+9fsYETzvidY7LbkLD
tWc4ToLOrD3arT8HkXPlgJizivuQ39Y2l9NsQD4cJpLwvFugzMy684mRXLgINx3uHlPcgPh4I632
cNc//4U6sQTAf68Bi463jSbBuwJcDRaSQQhXqzC3AAj6ZE5j4qC091aenUyKMXX7/LsegabY4wfq
oZmdVSuPC3SouAbYdD9Z5oUxTSKXQs+EDCbFiCCHD3+KuX3e+CCIlGF6KeikhvtTpFzqjBReT/2i
K7wACDw1+uFYGeIVWudfgSZpLvl2y1tkaqjCRDDLjnfQ8YeK6sNfZegqycq9nOKu3JrcV9x2ji9L
z5GxdfkTG6/C6NqDZfYTQjkwiKiEN62vPvupICqz6ejmh3NO67BzjI8qkUpsAlv5GF3y6xS/Z8tH
Q24WZMRYiM8c5V5e0ESnIwjwtvF+twH+J4HhOf96IagQcb84TK68ZQ6VIDrzmNoKPjJ8NZtgQH4L
GX6xwb0/9o7TSEcJO+InGItblCn566+NU8bVaNfuPCUFWXlor2Al8xZLEL5hEcvsaMG/BVOmvzr+
ux19vnxoJiflrHfh6m0KhKDDaYnKX8fhGwFXutEYjYeRv5rz/Mj3oA67NgYgHPeNUWl6cLlCD87Y
mMlF1xUexAPG2HGZnAnGNHoZSlJdyvQnGkmN0R27cm0vKWn8BPKWX564eF6d3h8wNBXUGjGIcZr1
RQ8YSykUCq5RpNsEUPry+JAy0DhbH9wLnU6INsT+RqhyyNe7iaAMuUUdPZL0tg7AHUDObqERhOPe
2WoeBcJNJwKbhpMPo5tY45ZlTSPbT0cAYZgIpMh/ZgSzY8tJZMZzWZD1pzUETD5WyNvly84Je1fz
s8GatI9inKw4+ZYOjYLuK50Ljc3/6S+QHMkDPXoU+UJ7JJvSrXFJhx+L07VXlhHoAB+5pzBcRUQe
k/w2MdWNiSKN9GvmmaCnU7NL0qd48TFcIyE52b/r29+ZUfHwlGd5QdosjMqywda/XtV3nHMojzWL
XBqCjeGh33NmM1bB9SsM3xhoTzNP63+QABesIlKQAMXI5sykd5/Jt5xVrnQ9Eb4OcQlomsyK64C+
E3CpupgZyOr9t1SSwI0zIjc+1aBsMV39He3ZGgtNTGrpzCydZrfHBEEObLcB1vCPowJDgrR9jUx2
dfdRk3cIew1bT0o96W7pgaZPQo7s73/yl5sj8F643LoKxNeNGVJlGcFgixN3i4Llyd731GsEjWTO
LB4bEaaA0SyOliNgbUytDnK/PSt5ajK7VC0CX6owF0f9VE8d0mR49i0VDARdEOqnhX/Y6MMwPah+
vOejQpSgq2ysRCeUC35qlT6oR2bfrCwWVF50VgzxxjcdIQSDRdj/M64xvmDklxe/bm16xms8Od4y
YrkEQgyt8bWvyy0SCx/OBSdmenz61jRV/sTebi2f1Is7aOr9ZonimQLhQ7rRAhNg5Py0GaLmPsuV
fit0StTGD8U8piAa9btDRHme8/eDP4yRqKQ6iz5gsppbknTY9LxhIQnk8VoYKonaCB5Jskc+VQWt
h9GUxYz1vEgPtlch7BhLLu6fllFHEOH40a0GD+8iy3plReMNhXYN7QNaiUhVdDEFCY/Sp5fpNn/Z
HCZ0W/2jgOBWnEZWKtXTmd9tm3gtT7SrJSqMH6GfTYVk+ADe1a/gYakY6snm7WPfpPRbx5BJzEXK
pMXVSy2OvBRstVkXSu2d1VvgoqVKZK4joTM7Z82S+1dXb969ljq4nxbjuCV7rW8sd1hWxK+XpavG
iIzHHsNrkj1IA4Zo64fg0R24zirGhq+pMdRHE5J/WTXcwXRLdlD4yJhZicXRzGq18H3Ros9RUq8i
0wG4rOyyc1irgSw75ZZCKpwiu+hviVheutx/sQ0F0zDI9Ut+zqkKjOA2uM8ym8YJuBeIjb7rDRdX
N1eCPePWNXam4UIMHKBEy2FNTJrns7e8QgqiDZktuHihL6GbduYhrWH+mP9iJWIrD0zdkD8x0+kN
JgbVX74rhSVSvnpGQiqmEXIWRvDR9kMyN1fotdu+jSYeQPh5haFTH3lQWFu8GPk7fBsrrrZlf/sH
vbJZSC7O2s4JFa1J9wFYlDKvXcup+iLq+k2pBgRPjEh7T3TnMpT2itsPCjImLA/uXtmE5kdaT+91
Zc5jmooOqdQf41s4D1Bzx2pNkX8WJdxa0aQleY8b1DxD24tzy5xdOtnjWfYUtQu/Jc8X+Xi+ikCk
4PLhcIZpRTuuvqHM7eX32Klp6dHNRQhMf5KkWr3gwz0lPCjRFTaYgN1vlnhgnzicIQbPCmojFgy8
lH8phbZIBUmgpjwEsH0NDZKlsmRyBAwK+NXzwwb4TSi22/3d4rE0si+yNL+Hk9ME97C7XZWVzRrw
oS8UzQDCHYwwpMZh9c4WhoFg91ZMWxY4wdbsnvTtKNqvrIENB2mvXZapGrMkqRV2VCQ31JEXOHw+
b3SLSjRqHkG7xlUHOlSqtuwTNXxEUPneUsmfiqLzLzFA
`protect end_protected

