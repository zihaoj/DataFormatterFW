

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HgA2IYn7DDAg50ZQXIF+3uF9LGQQ7iRnh9rRjI9Qf5gANpcevgVL1MizfVT7NKiRIjR25gpd/frh
i5ioFrwX9g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jGWna+ri4Ln5Ol4O2XYl54WWXvApiw4AQvHKyG5WPA/wG5gdYxJB5TsVgAEnuuZW8XaNRVTjEJ1g
xQEQ0pfMwvMIi5U6dbR13ZZNcJ6K5RD352bkLqoevz9cM6sx0mdobkv90Db/JxIGmA4NxmsNFJU5
OprkhndD6iP9cSc6xF8=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dE09sW8rfEVKAE8tJxbijIBoKg5aImi/bwGIqMNMo00RGPg+oZMfI/MapbgagkM8cCe8OcVtZRES
JNvPFDz9zirNP3oDs2Tt5klGXNXOmV0H9wo8twnF8t+v2V0VOksCnwflqXn3kNmZ7gktK4yiZrUo
GVG9bpriTIEerq9osaZ9zFU4gNqRGXMTqOCkqnVKc+guoVUqmu68nXogrnzzpdA9iZQhEHM4eRqL
2cZbraX6UijVKuKZ98sS+y0q40tEseAiD9qQj5m/TTizJ8N+QVgEEUTB7YndGZ2+7nWBRj5upize
jwxV2AwuUJL/ohewELTaCEAH54sauhn3IsA9mQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vJFMkpaFUDrnI4gxuqkHmRkcal6RLTHDB5pKdGHAIKJW9lwXqRph65+R46SI7MCZBwm9XXsphpzY
tUBz6PT7VpCSG2rrI2JAPI4Gi8YMyRIIIhcBRcUACFKwtU5BGWGL1kQl2dGkVReJoHz5rMC08XIr
8lHI7RXdVL0RJLoKln4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jz3Mt6krjLr0CAySESYUYpmpNSb2dzpouEL8gBb7U15BOyU5048hkAwGgdP61H9LcXSnDSLG06Eb
YLCo2Mq+Be79txxWDS5LuqgwrpUmspI0vd0x/0SPc2pTWWU4sSPsuw3OSHlXP83bjxUgZLwrFEE+
CZ9S5e26tFirr7RDMOQrjTM9ngvsabDng0ByxKwSSG6141sLFDk3/PcDxlJX63JCw4W+o6cTzXn3
/EfJownOkIBmT3+tYE1QHW4CylG4rnSmq5s9IIoayec7Lhih22HyCiw0LXNg8055ZFcHBfuVlvHm
nNiN81PGoBCrXSWTmw5QGIQtLWxsuW4jfy/Ibg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4016)
`protect data_block
BTd565oPHB1PFgXcRGdKttBF9UBUKxdvu6si4RF01VsLCYNeO+bxRGmq/sTsog5+iEise46iL8pa
bG+iT5iN7jyWolE0Os6FVHlR7W3I28ynPbfZAYVa2OXP2kkjxdzfqmgV686P0vs8NAah4sUtkdmL
tkRburpT/GdYPynJJuPIgv+yUHHK+ILmfYV3s031gIC7etuAu5fETeOIaYweWy8n2HdTvetCwOMF
UEVJTgHyyyTqurNbuF6ViNqzEdLsuLF0JnZY1AuwQF/GY1LnhD2SAwNTvGXPDyy4KmZpyODblPlG
YCP3d/8/nn6HG2M0CH64FEDAo95NW/Pr/+PyRvuEqtZBvEvXoYd/AfEb0EbLboAob/sVGkFNHwnU
6B3y5HbCXCs5awYWT71kv4OYuRsAKAdG/OGHB24QsgjOypo1/WZP6cMm8voa3s+1i51FBoTlilKQ
Dnds9fzD9FFFRlQqusuZQs+bwwDdFOe3YejWIK63pIvGDcSMP8CYoYXgTlJ2puwRM3OhhlkEWOwN
QByFSSjcbdM7f1zqno1v65pnC11QWRwLrMxhAGzEwRyEHbaDWhsT+elBelOPIlT+79f2DWQxa39O
rskhSPOTS885DXg5bRqMhvi5dEQrrpLIxtH8uhqqM6bvXHofcZe37NfQreCGvcYNl0tT4GY4ldyW
dHvWkLDbapzApe/rirsC5q/GoV2RnMmygpbW86nzm5Dm+Lvzb5UAcf/gUGvIN3K20jnU6Q0jysh5
daV4oN3+POomK/tTffm8NNrvPVUcOlhL0rsoiocNbDK2hAS5KuqHPJvzD1qnyAq0wJamX2+chRcv
s1Becfrkm5e2LKDTGqkrfYS05uU30SAy1P4WoWkA4kLNQwZd0kJ2ui5wa0alliR88qMK/S1YB0A3
Z7m7jjF3mGHFAzuh+Ev8aiOrkVXN8w0Zmi6oivj3ibzDGsA5Mw1MxDqbO4YpRE+2CvoZElOkSiot
tLKWieFECuhjYSkluouhEdYnwSfgCeSOzelcgu2GiLcmH9Tm9PqGeUCnJ/xiH1AWqYTE5G3lnAFQ
vcFc4rAFkewtlDtdDmPcH0p2WQU4In9jXj7wsLySfqKCvTQJ5ofOaj5l+ePQmGhQ2adG1hJo7qQh
aUEfqbqpKI9iyIFPqXFH69389c5JrGKFr4NkGjrL9l+7Z1A2Op+2+aoDc0qSzWIm8QPzJD3lkytb
tXjB8n3BjICIFtiocJdO2IOAXDNIpyBC59c6IVY7g9bqHsILjARPAvcGef2ILWScIktGGEsYrEj8
dzz7OYhwMJE4F5pNp5VvuklU1qST7/XmgKBLmob8r79aLibCXhK+lqENRu2T1sFJaUJi6h/Cf8RF
v4sr76RhjKOXuvALc193tjV/X30aQZQCQBhgDMgtuSj4KK3tKZxTWyRgVy3VwNV2V68hWhQ8yi4+
q6T8/0nVG0le5ZQpFWCzgQZE3rr6RRurZmxrFIPybPcKU3gE3HigfOFRB4TuC7W6xLSSf+UnNgtP
rPyL0Tii2e3dR2Dv6vmqjZ+AibGuO/VgtO/9E1NSrxzk0esUj/snjptbrQqfmr/BH302PEGlqLFx
ZcwYlUPY4TE7+ihvURsil1jcGI46MUgUBaesMJENLOmKTrgkB6AOlBdn70q7vwVy9lhrk+8+Jx62
pZklT3XTmfr7omg40SL/v6CZmMylabMV+Sv5LCLnudIlA/IG7qXHp4rpR0uY6PD/p5G1LK7T6e4X
AaNf3XqcFBk0e0uCtIOMpcuxdCOUqmgsGDojglmSLmpu60lTfOg5Z5vZDOootIeYbeQSx93lpTRj
xf3EKmpaocDo6Bebay0vGXMgu/Xic2Jv8lE+imrdL7eAcFJm316zy1Ja7NpWHpWBe7P1zymETcpI
IwdGHwUuPKLihm38yenN8RtonAI3oOJT+UAMWLLQ5cKcJ4AuvK59j5qJjTRkn/EFJ0KCoT3AfXra
8oPuX6qeT9aHmqbjtnh6GS7t04Dz+Rtgs2IlSSELAcQHTO4CGvhO0dLg1oq0sbs5pKKOKdSSIG4H
eMTNo5ahNNWPX7gF0svAKNMtc9hy+U7C8Ckxm7d+qNfG3grIXpitKuPPkXRASWwKpIKEzImHHyAB
7U5EmiZbb9I3AgkRpATZvDSmmW8H0/TfY9649zlFw5B/atWGezOJNkfwmsqFZIc1lIJsB6oqO6BC
6PsMtcMfjADfNzQLtYdIGiNsvGsPZ7APiWELEzbmlJ/aXt22GE45hAvXKF3EyRdcWS+ThfSGEYQV
PSG2BCTeeEDVYHlRuM1sJICZ8z9+3LtZI23hTUwFxJ7O6EEMT7yTQ+8k6dhRJIn7T4z1roEDYjsp
hF2b22m9+IFOb8/mDP14JQU5goJQlP1xyMntVnifoHRlHQ0E/d4meh9kdMHfrFWXuQYynfymsv9Y
25wCvzOIaDX1Yn7F48iiGvJ3h7+NPjERtH2HXOflBXGCV1o7xbHL7Rs++owrLHHBTu24vyEfj3P7
+gkDOJMW6q2JbENj4HWclp2Ntq7D7J2hxDM2muGSdj8XIVL7ngdMaOSsrGSFa66GIrtJHd6VBEvD
kZtFB8JFPuoFWLnQWfljVhU4si0ze75rPI8ZjIZFGA5RxaKhNIm+wQr8uE9k/EoPRUmiVAk5Cxi3
z1bg1qLMgnpDw1W2QLZnGIeIfR6Mv/zdCPKF0aRA59VvokshguYdDHyTrMyUmabWykKIYr7i8OpH
DE1BJxgf3Nox0JYauS6v+j01Q9ANRCjQ4wxOWvbHfda6R9e/bQBoK04KDi6m5bQKlUSDLAKatTmz
tw2TFatTm/Zqi8QewTmV2VC0aQT0ufsQlqwICXJTv06qCSZYHoqqT8ubq2D/i8aNOW3h9bIU77Ix
+1yHR19gA3XsA2ppCfg9/FpeEX4QeYoLXDkCwVVAmsAZJ01kVa9AEneiHUsAKNC1InmrxW9gfC8V
nAcC0gvfnYGpnE5QMwEyf5bF86xBUwdVKa+RUrP/KA8k65sJwHBwgcgYUYn/5JWTiyG+wr1AycKH
E/DC2JO2qVgGXRDPAi75+CdsUCw8VE5w75gK3hNdeITvZXKhiaeldynFT0V3KW0smfDK/2ibxObC
fmkkGcQbiIIDYgOO6eqmzFsEwosuG0MtAV4I7h7j0cENjFcA7PZcdAxuDDZJV8eewm6CuLMMrjbz
CA9zbifMeLrHvCcUPFL84oAf5rSFemSQTYakDpN//VmirEryA/luaXQFET5vXcj8JBnoLAfIz5/g
wYF+LL7xMUKOANkpiFGqh+RmTa/d8CeAbJz22cblc7J+lndnwONAvuuLxHdxdWNRYApPqklQqRGv
rKECG8cdACwsfv5rLVQeDb04Kod1d7veQtQh2UiYQi7Z0oH1apcjtDpnoLmk606wHE9Q0kKbiGJI
71sZLj47u1SslYws+MkT+xPpsywpSm7NFVsnUxbGt3oy/5DTjSi3HDBEL89HhLMHlfZFiR4iYQYy
2RA0bSFYOweflR4rnx8GvXfC/+ywveCwqxW7PD8ZysTKbsWyQoQatEEj5zl9YBIf1IjVJD2FSkmu
uhrSO8hFdDNtb+0CDqzV9pUdZlPwhw5qjwk8vxKG2oHf3IkX+RAG1lAgnutODwmb6amPdj4IlkWl
0mBSDsbFFeuATYslWXuktrR4N7uNDHlTB6/c/jXF+LxWfPmYCuFSrdwYFtEkFYaGcJFkS6tJJpck
sVBS5CFWXwddcMScxBLb3ffGThID/Q1rTzzTg6EIYr5v5mxMtAgnZW3RZ0VNAaggYTlqUQhImLUK
SIA73e3xhumbybnkyw95BECvBXyvYV+G5m1nr1KQukR6dPfOhT7sNJoBwFuS20YM1h08v8pZpHgu
NqDGjnJ9aRRPhUasA8k4VQdgFOTHtwdSsaUC+DiWEeENm90lcrKy7gNiKp+zIxDeIVyF3UDcLpzz
TqnTw8f/1RIHtI4kCZGPJtsms64qPtJV29fJZSvq1KoncqG/w2aYyouYd2E31p8aohbS1+YkE8QU
N+N0HhRK607sHz+I5mIQqJlMgDXW3XGN/z/cOixejfypNyncFflknOtxOFD/VQNDFGJ9pFP4MDxM
MwNu6yiThNnjBY3KB6BuOkbUdsjNYokXVrcMQfk0XI8ZAPV8yHNg1r6SU2k1LmlDwH/E9sUYrVN/
NZgo6/77E/C8JY333LvNvbcTZBS8dhT4g1bAp04dxx+tirZdX8HbU+6O5OAdOPz98tz3K/FjClup
87hW7DSZ+c5XohdoKIVy8MnilwHTzfJsA7m22B0jxgABR5KvH5s2bIrJT0xp7pxfqHsQeXZSBB/M
c9aUmlp0ilhEtWETAlSLEJeImgcUws8hC/YK9WhD0gnNnqTBVRqOPZOJI+VHSrqmPFVhDJZ4I99T
yRyYjVaTDx4/46rywWQAe2s8EuUTZl0IR4uWnCneCl5r1dZsjumefk9wMfVMzp/l6416DRDrrJmM
V0WUrWpkpcKt4fJ03QA9FFEOuhlLq3PIfwNbk84niEOG4r7D62wM2VNCA+AME5/HdPzS2HvL9OiG
GGtZ8YkSEO302puJjRUZJsLfI9NtvDCmAxuN6vOuKD28+PSmjICC3daWR96hazjEE/kO57Hcjgbi
wnOJr0ovu3Dua3bkrCgXetTn5ysCtPH44cud+zMTHvdTbB0Nppj2MXfUXF2NWLlCpd4pD3KDzhWF
qHRyCAqGUWUTGAoyczbh73NRdn8aXw7nZ/QHLm47lL5GAgIERVdqqwjnCAwRILF0lnwz0S0/VNf9
W4mw53+Z2k+m7zn046at4DgEqvhhLLC/qJm0ML7bmNrqpBFRDY/sygP11MLzmXsSJJhIz4GUB2AU
qbsKUBEhM5DzqSW1GZ+tMc/rILch5CQVTheKlc7+NP/BZWoI77hC0xuZrfZDmWuG1TN5SVA9sXg3
PXgXT/hsWwgTvzuHOfLMHtNKJGvfkE9weUkJJnhrPE+VoXBT/svr1SDGtmdklAlRrrF+IxMudS74
2P4PO2iS4wFiniAMnmKOpc0hXdWqkkniGpsJ4Mv4ubX59oXkF+LoHtDIxYEOYYUtAgyPrgTCmGr+
WwFLUDIErKziSHYY2wKqPLq2FOl8EmYZiGKzh0/Gi855wQWkV+JTTl22ULO2utVl+YhDiVhgzmd4
8n6NTVQgz0Ixn1EjDFmFjIwTPzLfMDxMotT021grs9jkpoobtPojPM0vB2mtFG8ctGTxvrdCfuWh
EjzYWdvQjAfexEuqjz9lM4GOIfZvH94tso9mGrGE6xK2jwud23vyN3EA2PGLehz2yyXOCByXYf83
TItVmL26ZWL3RoFSouLDYd4S4q9tnQKtmJk=
`protect end_protected

