

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qjH6h/L69lfQ/fpshTcu3+eBzk3cjtA5SGJK5TEt8SAe8gYC7kvOUZTDwj0umHRtud94iDtRK66c
0Gk3WI/a5g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kq4sklT4PBRNzE4t8+rEfcVjcFPywHeJHvgBXGRvFFp0ZvAVumaP5P4eiQHh9Yh/Foro5/WLPHrz
IJRbLfvT3dAyYaVmDqy8cesBT3aTlyQezB6dwBix7yE8xaYxIcjz9VKwg1pck1CSaly/Vbistl8i
qdWEqUipqYpNG3BG2No=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jNDEemmWm7BL1YD96qwSLXre9pt3z5EVHZqFRG6rrifKydzdejWeAP/El/DiEq2n6eTuFX2KJ1qE
la9I2PwfNpU6VFXpsYra0Pa5vCqOXWzufh8m3khRrty1eN3OVA49uGESs28fYO4NDevhz+kdHyX2
AqEe4YdAKibBc3d9WsrM0Sj1OUHvlRQrUzT4yBBZsbtUK96zZjqcCvuaBnR65ysCTAOgQ+UOAccQ
e3Fds4uXzxiWY3fHJPU3dwOLMIvT0hLuX0hfuaKNl5rwQ52uPubmfdmksmxtGbLtI5JL05VxTwF2
6UA+UF7TlMq/zoDHp1M5P4r8W+PhQ9m9bjDivQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SRouKG/C2Uh4IWSu9unaodx39OW8OGa3RdcgPSIqQtUL0oFvPlGZ/IoUcZDQxw/zLDzTmux55Wag
UYZbKCVu+WweMZzw8QS5Hx85TX0x1aAxsuFtNceA6L2Wt9KH7O+naD8SyTCVO/O6l6ZdoHQDkI9d
fGz7TOavt6CDLAOYo7U=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O3E414Dqw/uxwCMSYp8Bp/7AsE1RloCh067sSwv5pC8nwKuyopFMPJUq6wuGF1vVVbO1W2yYTayV
XZIZ6gUmNlj9wohPF5lv+HXxr19jtj9Wy79wm1ggvGAYG5minOp7BEMwkvP3Ca9iVVVnlw5Cpmyc
NGXw+9XYOTMSsIJoxKXhjucmlj4AuqGRTAwvTZJpe101GPt7r8PnS4z/S3oNnIbsCnieeyN3iWW/
9KTbZ289N/9K5uFlHShJMqDp88sCX+eTSh1dczD4vO5RnpkfI22iM7LCqqtgvQjH8q2OZHl6HePQ
uQrfik1yQac/oTIaJIJLR2cllMzIlAtSkpQFsw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24704)
`protect data_block
5mTcZYZWbOBQCmzhVsFqUAkOze+3dYo8xVUYNrzZODVn5EFbWq3dyLyA2mWPjjbNXSlU+eM/sjkJ
x2ykuodT7EO3aZvgXP4/nYPp94BD3YOLdBDXzyK0HGM6x+8LO8slCGZAXNdSduWS+FycQf1tZL36
DzwOiHFq2cXZk35sUvncLa2tcCMKyoYiR6C1OA4BmOUom8abHqf3duTmyrdryg7Xnd4IgEXD5QqS
ArVa42uIAUp32kwriEzvjgZ+Y6Aq+MfK/pXPOR7ON08TILXFPha1XBA+iQITL60tupuxLe0ZdEWw
K9K71vWhIL1+/ScBCpSGaO/UJg8GqfEZOV/Cdkvu6+ONr1YihCT2UD2bVdtzrBfb+2PLJZB0Z2di
VYxwMimbUedcOd2ezQPgdKHCmrIU1Mwu1c70p3502op6MRjxHWMdkGiiS3rqiCkdFeu/CsxvSCh1
0bS1YxO/m00HRqTjrkN/yT5FSgHRPOVGxR7dgtomkUd+ufX/7F+O6P5Ym9vuVrZQhJaq9ofumf4w
kd5lXG2WTlrckYj/KqhLNFKXk/KdxOfAUrB7wIxXfPmSoqP0r6adRf7TPjijBZMWl+6x1enrJP2g
QJvVq0/MFq+TCcf9z8gl+bAwcX5vBZStp4JjqXPpSjGs3fy3MtujiKme0lz6EnMmbk2WXzV5RO4H
UYPV3h6hJNYZGNnbn3TEV2KGFV2lA/TwBw+AoLqA/PfnmnZYR7P5qdldCxXTHJlAq6oqo7TxbVqt
pwRnFDo0yrKFZ9c7RrDvTLXqAX1DMFibP8rcv150oOSxVVFPCWPk/z/WyE+m7fRnwDGiEUi3fUjP
WvQnEQTBVGWYkhVhwMPRC1tG279VlOa83BgMveMOeALaahNoWxLwDbSzvLTvz/QiL5XI015Qc4oI
1akE6JLBXiOz0R1i9RWnUlXT1rSXok6q5hZEu3sG5obnlpHwdAIO3UlSotYcs6nyMy7YOs3NYqdV
oNGZ2XmpMjJBBMd+TKia/g14OSrGRA0JK4Yj6SyHcXEc/UuvVrTCWa/doi9np2OG6O+Q1wqapgOl
p4pfpP8W741CWgZFjrO9+C3L19/3nnYOgj+qnsKXfBganmf36nnIxAep/2mWemuz6X0o8QD4+heA
bGVWXuHgbq2Tl591arvPr2ez2LrXm+0C80E/iu6sFTpa5GpcBBep7MW+0wJzEBvlntqv2wjHQoWi
r1y9+IgWbOf1p/LKbQnS22U9b+8DTdJ29hln/d+wdewPVkooZ7/kodyJnCNe4QtZBoIDrmxlqRLi
XiE82MwdnQfCAB1uzTuTXPHrPYclhJCGQt/KHcO9etlhyNBIPB69yrv/3q+/EDhWgQctDkTsL6/J
tuxoa4WxqCUdMrfVLpW5cXXL6tHYuZlscxHy36g+U5Nj3XHJSyslkx6ITzcV1zV4h8cRy3Z6qit2
G+22BFdxgMui0BVY/Um/dasuPvEpxHsk4yACfbFp4v8F+yulQMw/64d2Mtz3AtAUBTeztuJ+v6PO
/3fm+7BdWJuDm0wYXl75rH9F71nysLsmDBbtM5rjTwxKaklr1WJIIwTcqhx2fmOU0I4wnYqXiEgd
kqy/ZJMOOq8qNOwEWYjoF4OUep2OvU/odZYcqL81FBzxG2+6rY6PkJEOFAds8DpLWq033dUI6YeF
/20LHdr82lOEDqlNrLNJPvQJk1prVMohNCCvSHH3O+jQn0TO+9h6j76BYvppJMA7xO4ahk8smmAa
y6+KDtwMMmOiPksxHQZlKkz15+vh/PxQzQ/6Uic0MWMRjkJULC8GzNY6NhtAybH8xlpvlGwRZWp3
KDz+u1bj3+ESvlKveHIm8HASOFdz8OTZLXNYWMtX9xsPPjSLzgkD6RHI42JaZl6GA0ppiBBqZCD5
PCOFbFzcadtgfC8c1jVwHDu04sBMTog7ZqWrQQxMetk5MahBETRFNIJ6GYI+A7p4PFqrPks0ivy2
SVM8x67uzyQKNxris2dyNZHY/XGRRigtH97xDzBGYyuKmaaCRS3CoRlXDzN5/6GIZW0XAKRTrWYX
bQd/CnYbSOgENl7p7PPzYaak2ejpdubrOjitL0YGaThzBS8ABZxBkM3gmS+aFsIfODGSrnuav4kJ
hE+3kuFQEdvv6K23aVfzyfcixH2up4QgLP5oOQHpF31faNDsd166MvuM2+4af9YwbNQCfyr34zY4
207b4e0TG0wUZwJTIwdTKVIMixUGTSiR4dgbCIRE0G4DjS61ycDCcgQnJBhxW5sQU5K2c8kgVIYz
EFAyeLGlU8U9oLPQGMXoYS9mp4PaUMO1IhTWiYlZg1bYN+OI5zt51/yGkM/VgsPHG7rxcHySPNmt
YmL/PZniZ0BYujSZV+MvY6mYYvHNsW8X7TVDplaoyJ8K29CNeEjDkR3SMVrH46HtmVaV+dsq2YxP
jLi93pGki4xxxuf1HT2BkUqiThAj1C6wTWW2BbgthrMho/LcKNxd4pEYobbw7m4uJa3XcUfTwZzw
KVPn4/hbSu6yQO6ymZg+LAO3+lm2lzmSd3g50Nq77kJOYZqvn7GsP8qXD15zeOGFQS68M7MJ9OeY
DQaIhbHv06WESAGVj+50kYDL7jmZRrrvbY04w7CktO9BA67ZUEpndSXmXFo6Xf2/C/EdBD5KUoFe
ZiWriN4Fl6CrGFbKqxjUeUBrhJrdaSac9qOUDWoG2DrK18LaDSgFNBjU1pO4g6qxtdusUdPMC+V1
+BUAq1y+PEs6OHm7G8wTJ6VpEqcl9UzcAUlnnO45TCQn0tz5GItxPs5A1+6VPuxulpObqbl/nBBh
eb2JQtN/oXbSRqjpjkgT+jixc76qWO4dOIyNEadz+QP+CoMw00uEh4WTUsDR2MaHvPWE6btWc8Uv
h2i57uoFWDzfYFW09U2V4y1VyFnRryJCbsec8KhzTgyhdJaD9oGzJKqVkHWrGEXB1+EI+NdjV+OC
JROcYSlhdGkQve5KeQFoXkW3Dw2zXttcUiAGMmhsWxnAy3Fu9r3NsdC4z74CT+2f9GpB1Bcgwfer
IIilNTFYhgE10YHrH5CyDheHQQLQ0NRvH0/B3o13LjMtfC8MTbPRuloz5/MiJVy+7vnvD55lz9Og
ZExqerMWA8JkpWDkR4PyGJH6p5BiXV93HgQlbUPk3LqifMnEugyOiFItwDwPUwlzlSjzw7jUJqBh
qUKkEnAqXyWPYrPQnCCw389zIl6A0mf3fJ3GWzmD8uOppI8NCiY9a2ACGZX6Sem7Mf8L3glVPIq2
Pe++VqH+8QS8jGEr1HU4ZcGU2NSEQxY2XoONmRHOzJ6WFLXffMhWmdxaQNRsaU3WaaiYWUPVEJB9
eN0pqoKz96Ev+3L+q4orKH8sm19fwBXg3aoMb9EKgfX2BPtHSq9UK54i21Iq8H8t0/gLaaigLU1k
qpFw4Ljqh2nj6APhIcKEDHgKX/ASWGoJ9PGSSUt7CX9104MeGebxG8RMdQAdoto6XQA9M1Hjjg3g
rFU4kZzdNT0lgmB6gVVGXk/WZxBB/eKNvTnE+eRFNQhVTeXNmSdZeM4i9+wfQy5vC3uZ8n+b3Thn
OLH4fQjaeyAEZiaZUlSpCTKvMzxqc3NaQFI/tSALBeUdajWuYdwpSFJxSO6qvt8eb6cJW2Hu2RZX
Hgh82T7Q8p2ngu6KlYT+bTL6tlAbBgKkymtaJV3UXvxVK4Zzk8nUpIf0fhvIoPNK8g354wp105uH
HZB/ZVpTMi+MOeo0vol/EmFMs6pmy9RWjDZfJb5PosX1F5ur7A6nnxaO+nI0UQ/S2847MCf66nHc
d2B1JWcz9YEz751kBPBOONNoRU9JYDfLvt8q1fIQR8uE7BUehn2ZNAI92xqI2UQk0yY/L73hl6m2
V5vfcc6gL7V2Hp/d/qtEhf+OHcC6iLtBE17MKGiygH4PuzKMFV/0NC2EjA+sRdY1cHwX/kmUuQ/T
xAMkSbkHjNWC82cnLqkoonfIGsr2OdWl1BtnFF93ebxEbEtHUn93J1DadD8wF8dMqPw/ra7M0OWV
TujIMxazFEMON1eRoLFC4+iXKFNzX1gNPR2AxxaTw79A1uMdh9tzJOxskX0iqewxkAMLmhOigDMt
hFEXXJbtRKDXCTrTPBVuw3bcHMrH/sFLSVMFK59TvoCT9TJGlYJPYb5Qr0IXH5v+ec8MjO7ebItq
T2tjgy0yryDZaCaDbmV2LdpJhj2+VCPVw7JzAK0mdHCbfs1X/5Vtzuv1JFaYA3JhEZe2ohDcDsuX
bDJFr6NtIDx3GUVfh7ARzlWvBtDEGzHnf5L5dWTM0drPaTMOJUF2JvslbOtW2V00LvEFwlwf9shC
P9lZasPv1b7Y67iKcZ3nCBhrN7bFHsBLXo5kdVlttAlxI7op6x37at+UphuRuhm4MQbi1kp+TDhq
KALSLGd4gYvMeVfu4OkScQWhmc5ra6PjeBjWMDAn80mX+JZPb7LJYZ+DKSHA/G1h6p5c0BoWjWoU
R1zZr94inZimV1rl6PpNs6lNTM9L7PrYigKnnsQoNL9Ym1Z56QJ6a3x9P3g7bz6Xfp57J60beB3Z
K7vWwn7fvJ57PhZtaoBzNqAVyi+wIobvIKk3q0LwcfndZCsyJU4CBin+9E4VW3iChAmpg4rRoekq
Ddq6+9a4EUQ7sA/QejqmfOfGvEETYHJbyTufbrBbCxUVQJXJb+y/arn8KeXP2sChnHkkdBTFzWyf
FN7OXxWKZo0hRtgR9GX1p1f30IdEE0h+GzJaH3apFswvdt2upXqb7/jae4Ku8YmW+YPaGF8nVGZz
bX+wYsgb4Ebr61tX5b2IJ5aytHCjngJIQB/kYlmRO18w1iWDNwJiP0lbwhMI4hp26N10wzcidFLt
uufETNML/A0XMCEdfDLgL9FnBxBBG1YngDCGzQlvtFecVRcGCUNv9NZjAb08oc3g9BpS254SIsyN
CGHNvG9a0lMrvIItj3y/YcicZBDYiVMJ+muAujnf4IJV8qngyYpYR5Ayiydt9EnxRhXoXFLuAeny
V+6WG5qBCibp/0ZrmCNUYdeWPyUJxLZH2+QcedEuGMyb5dbKLP9Zgq8uYEbb48SIkumJDM2h+Tr0
UngublYStYGwtE45+Pr+O5eKXoQ4rBLOMEYILT9eaFVvCd21eVwSBFzWhcjKB9zR2u+uaKqU21sQ
EijXzHPNOMxEJbW93/R6QfPhvQwlV+5sBryfeIK2/LWa+Nk62UyN9MkyFB+FkXq3MfrQMAuSBoop
nhN93YoYhneZNb/iisGXUqD7GHwZ92BS+9t7DJcjKafHUhqiroNEehWMZLk8gJuoBNPCZ5OYrEQb
+MBypqPo0S4IFVCCTfMFAzTK3pMGw6d8bBegTK+Sk8DVuv2a6tw/s1iaUkRFMumOQzLRSqqIkiLT
zcONAl2F/rjzGW+RNMfMnHyg9V9Xy+/BreX3pg2v3NKeA/kJUuk0xpQLEy/iIxXzx1pE4bVTfy7B
DKsgiC0T/aE9Zpp721lmCaos2veH0VxV9bAyz5ulQlWU1i60yQpebH66IvkLltjOfVgUuycUP4w/
kMNjZQTJeILuyCOowTVMBoftsW4mXHe/0LBBSRtA9kBVaQz4kk2IU2VtHoSMEZLFxPbqvyHlE3mF
fSp96cubKIijV7WSpByOnjz1TIoD8ZqHTV0gjgtrf8Qrhf42usV54stCub5MWGe8RNXmC9fWjK8d
2udpokcgcMyYCfFfOAKxDpoZf87p6E/Hl+y8dIHhIpwOI0qX+yFQ30naIzufrWgLMTCVr3kKRhhD
faFKAjSrakXn8rLbvJF7WDYHfbb77O3XbIXSlOvtRhVmqZT3FfM3WMiSGP8KdY1Q6RFCXUs3TLVG
V2zKoWOxLx1n0fv7uAK0+1DZ54TEFQ3UvIhOv8a3qrA7z46dWSoeH/1WUxR/QnsojUhT9WnzWo+q
hqQVwW7MEmR5quRnn6sSOjdKxBnS4YikRPZXYTcfAr4zc2DIk0v6yLWYsW3JsqkTGWRVyxCIxdt1
IPuK8lSU2jxTzUJJ2WZlaVb4VjkJ4AX2asxLbG+lm2ys+roTS4UHtRVwYwXsBKQmar8RjyRGsIUb
/VLv3gGHR8X9cRAuHyl06V/YCP8yglGSWYVC5NdZoHSFgbWFDJEEGAI4OjuiPTOwyB6PS6Va4GZT
5pHzpaG+CtWuBehAsaIVvJvMldCnPyWN9ZEyc+Yr4fa8aAgufodLPck27sKUJVCxXPdH3UN+hmP5
RcVeq1SuA0HojQ/AsrB+RuFKmW2yz0/nbAMtTxturXzbjeVLZzUmkQEUuL5Q7fHeIQPVHv0uhzrB
mGGKvp+G5TGwjr9cyiAOVbJRGeqPwl3rLq2zZW9xGqwzu4SN0I30u8DjryEtJnPN3U/0nO6ADRtc
GaMEe5gjHXoLZQXKaWLlpykvT7iBSi/OhpVCCtbfXGRmho5Yiw7HbWVy8JIEtGhEGnMGfYDyAB56
7LwL7uSyeMrWAjAd/xmwmZvo+mSFwol/wwjp5q2zVQbdkD9xRb5ICSwRP5OycgtBADmIFKXhWEql
XQuYL1qh99OV5674KJzLkZS0CsZDVdyg5iobmyYI1AE4wX80v7P++PcwOELywpCHJua3DXn3MhJ2
bkBmP5SRHG5o5cWUw+U8Gx+9c3J6DkC1iim4ZU6bnCVOeAe9q5wE2Qw+dwAECVXOSkqL8/zBiazm
+NOh0UcbugEYnnaVsqi6HP0oRNezGtOL30dkrvbedwDOObs+ZvN5Fhm1NNMVYx6BYzVY7ZQvbcTg
Hv8fVJGypfhZO0lpE4JFEF/RwDAwcHM8nNLxBQRr4/Pmg5VShlO48NGmc1ldWUnWEtfYGJ4ZtQ0m
XIpwOyVToEOx+xzGgB1GTQEsI+rwcTfEY9b2ngUDg/2r+a94sJQ6KuX4KxzplkAXDIoJAx4i9IFe
e3yeR8PVIYaVkM7fn7upld9L0fxgGPQlpwEe53zak8jnOtV1D0JLFDfsU6tk5l4DW+I17w1r4FZi
TafqitchnJCdl3V/yHOaC2US28ELbO7PsAAy2CSZz/s82gywpp4G5vt9AxRtcanB23VXJ4uu6A5f
AbCNUUvt81WnIajTRmW14mAx+pDt+/mo7DlXqTo3gviRnaWPv3QxMUemFkCPCN49RII007W8+GlX
zfynRiOUk3w5YIBEvOCZGkDi+y83U70yJfbuQPCy2NBjXI9D6ZWmTaRThWsQ19VvqL0WDXrtlSQ0
FbVnG/Y5mtlSq5G7xDVEJUhU2pgXsFpgdj4XdpFARBRF63SGMY0j/5hnZ6Jd+Q1Pq34hf/9K3jJU
oVDNtFyHrJGycpVpvfaUP+fH7eVw1/2xqGRXZ0nTzrynULfnEtjMvmrXZscSbN8RO7//IGCW//OU
C4mUwYhA5BlhbuQmHpIInO5YdIHQ9RQvcRd2fyK20c3IONslzpJgmeycETB2SRCQ0aPNxci75vPU
EK7M6ogBF5a01Uy8j02uUqmWARL+uzMn8YpgOyplUWNwLwakbenaBUl6ygVqqFhTxewks7eUtYEq
KLFMQciMvgRHPznjvsWl89zgYktg1qWhG7qoIIu5FSDwFqdBVVfyCh+Z2yeXb7zCu+a5dNWS0oB0
BoLVBPLIrlR1q6Y+G1X4UXTlkmiyOsIrN/9gp57O8jbmSU1vWkSaTyZhMOB5pjMoZ2UA5ShEwMpW
L1fygQIfFqDizxH+B3vE4hB3Im8lbH9SZR0qbIu5ooGffSy2mXC16X8jkHCEvd9/C2sP7d0qBL6y
nBjblOvqFLVsWZI55Nje6lZa7uapj4yPMWqD/bhYIB7UFuSX8m+y+htK4Mjka1JgneoExFuB4sQl
TUoAkC/zLwFJgpTvOUnCDbFEnooc09czAae64zdsbrjS4pBL7WI5TR+WqDB3QlflIyfe3ulgqDK7
XNwsvSwivzI+E+M0I+NuKC2RO7FUqEOM6G6cpm8RQbB9uuHSs8QvWlT8+86yYWSsA+GKYO1Fa5Rm
q+E3Pitq4/5XH7Tpd3S6W2HdupCp2RtArsoPkKir0zbBme3tRW/yfpa0VbbgxnL11Vyf28U/OXtx
rvOLQxNgQKI20Dj9Sj7Ppnzj7yieFrH30rn0qAfPfavXy6W2RENi158M1PyIB2V1B8TB9DjdB8O9
TdRWPzlz1tXXOOvrf+oqcWy6A2PmxEU2R2q+IA3pD7ZbKY7x84Vt5SvKnkU5TCrlbhcLhAH+uNvm
3cUQtU/9AiiRPGxhXlWZ2eyGOddw7lAW9i4PRKYhE9eya0JRgeyJYRm1MiQ4+JmLaZCpDfUl409l
YV6LiBcZuMG/+AaC9nEmBc41xSI7sXyvoYH4Fc8t2eyonIjRvimD1zKG3U9hl8I/ljJjpxEEmEqo
TkgaebCR9k0+LswmQlj2txphVtjFoURjL3zWHHjLWr3xwRgDkIO4HPwtXn/+XrFpJFR7TGqRvWZv
T80hEM2/n4Q7Lw5mrXaBBQLzsljTDMydkRUY+pDMWraes+APPSyqnMRmmUb2vMus3dMuDs350ZeN
Hm3PWwSMQZWmeTK+fCrhV+ZFViYHPPNZW+Zb0UwR4Oti9f7T6M2I3JeH/hpgPAvgE3yb2xN70ub0
8nCV4b9BYl9dNUT+0AbRLuZatlShyS8JdiMs0yuL1zkVi5UoFGW8g3CQQawr29V/yihHA6o6sJSg
VnlW+ZcVualbDSeOdHoiwxi+JLlGTbz/yMUFiJvXt+w27fDBOo9jBE+WQl7ndiehzV2N5yVLvvW7
MXKjm9xUsMXS2Vx41kGWoA8pEKvGFPvjvvyxkyNKjNf+ggLwUro8gbFe9kmZqnwVXETAKK9WDohk
TMXpGh7TufRYgGaKoZsvYLYvbThi94aLqnNLr+jKStK7cA38iw/D2opB4px/1zzWWw+yY48a/PoT
QZVRtSypn9iHpGBDyu1mP8/dhV/MQR9rJlJACxAn0O3YWF+y30zvKLbH5feWJEiACcVAlAjVVd5i
fJsH56QVGK9+cLxPUPKW9NtXMuClBME4OABNsxjGBUQzvh/7TcG5+pKs/3kO20QyE+yYXof/I2HJ
4dU3qTiesQqTzAyTPuSmbeUcCsc8l9l7bjq0Y9t7UAL0zlIEkO88bsRyrw4YhvW0A//OUPHy037w
THaTUIgOTXojVnEGLzrNT8w1wEB1xafnzWnWJevhieV8v5X3MIgAAiR3FH/3GG/kq/9dGUsJPt6r
nOsGYwWBoFiWQRXRao8IH1s6oI4zGAM0Q1VCp2hr5tNSg8OX7Mq/IstsvA/CbRwSAjNL8dNCVc3P
4MNucQ9P5lEYuaIIxCtOAlQlU2MJFlEGQIXeMqRKhKdZwlPbjmvuzCcAXWUBTuGo/8Crvs6vji9t
UNCDbyTCPqXRYlFJjg0m/MSSMkAqQnXeBedNTUt8m1GWZWEWkqhdXHNYYFGRsYLlDmvEA84BUUNV
T3JDCkd3t+ehFYdM6bTVZL3Izb65IRUhlIQEPUxC9qHBzqbek4W5Pnmwe65ontatsK+pN8PxRCYa
ton6qkjkYwofQtYRQeDx35305InwrGdHXWOd754lAnejo0IYkF90zsQPe5nR4S4HjFqdjV3yIilb
Tr3EYv/Yn+ysHnvfSYMqxl+pYXKDe1MVrFMTdULjVk0+FTpMwYN/sopxn7KgreaKyqy87nTQ0rCE
zf0XUR1fc+dxhrh0cQRH7zMk2SeIkKL9qSeuvTyu/M7cVkcjbMgJBxBizyTw91kFYzoBe4FEJ11G
QTOVLyjluh89zW/y/MzYcOrWTNPQd+onALASTp29W35pI3jQgXq5E5GpZQHeLqHLTaroxgO9ndq6
tf40cwAxXPqQ0VhGn/8QCz8wDVfsp908/5agh+Sob4/YAlAvbmwATECPYHWs6OfjhuiaCMpiVtB3
NWFh6HLfVl7ARL6AvLKSlmp3cfrYO8kyZ6uCSZoCbPb8Y5bjD63/UAGTR0Jf0HD/c1ar4YnhPibC
bffPYnoFW1/P+hppsdo+pc0ppmcmGP2wwtYbZH8BJ7p3x9QKRBgeQMdUQ3+trUtpaEajwvQPYDsy
/tGbpDBLwfqqM9KA3PFriG4QWAa/w0g4SkFYuNzpV27ZYVCfhUrRVwshJZyvKq9QKvu8uaDgQrUM
WiNgglj1W8b9t2DBKUxIDtNSI4yPq7733YzbDo6k8jLZpa3PQxTFLs0kwN04ldiVEXC+JCPEZJo+
N/sQFt9iy/pMSyKUey2eVBzDaO+hrNDoPzy8fRldmQs51/x0/nt+HgZWg2CFKJJB6m+Q6wL95VhF
+owdTGck4mARW/yJ35ANZoVZhcSt3BEf31eJteCgro4rEOH675Stumv4GhO0dKO7nD6uxwH1cJsD
OldXa/XfWTXz4sk2TsN2wA4FdwjnvaVNKERATWqMlPsGWRMIPIAO+TZEgLP4q0fVY58KPXo2gZvy
Ar9YOXa/1WuxbxMzwKpOzb/ThVAm5LW3xJG+Jdsrq9qfIsAlflGiowwoREz0MKqdjPsfKMXj1QcR
hfhcqTrWZkJgg96gf+7Sdry+rHofhAqoE3Ya0Sxaetqdx9+SoWexc6fRBk9rKSNWPdR3xqinvJ/+
w2rkGwWKL4VEn9h87sTOXICbUnjAr+dIaPCFr/wVVD4UM4f9HdjWbSCwehi5i46KZiQKhECRIFFJ
lqXwe8/mzQErZpnbD3qWLfT7i0dMdyLwkWsvHzijBDqOd5pu+e4KZGiFuhASHw5TxeqsaQRrhhmU
zyoSfejDLTwVWZOGuuxxcj0Mdu31e+97Ep9qOIxijUH+1ff0Bv4SETSR3bv8KtZNTjJdnkN3uQRt
Ozapkf5J3I+SB0h3ex4fyI+7ucu77y3kUUqT2XsTMmHNpNVonVoIxvvEgQE1gfZe5n93O9kMSBhm
mr2blrkQgz/FaMtYf1o9zflN4Z1Wb27wLnnNI0fwxeLR3tx6Xe8T7lyJkv4Fbe5xm+gWuU4/4/az
wYOMRCoOblJgri4fOGok6KcVhN3kK0lj9ejbLUWH5qDRKshjvgkAa+D7zf02Xy0yLTzB5aV02s/a
b4jBbxhDusX0Ba3c07iiOxJtejMqHMUHfg1rkCksnxLwBOi+zFTuzrd69aeICHeZhVP56Sl8sEMl
71UeKicbBWmyFVa5HoA1yy8HobeJ2e9bhsM2j53p6NGq+JfU56y4jEEt5RT28FZRn7JG72u3adsj
hJTtTBTKLrUo4JGoBZwB8Zy0Fw3t+blMXnZ4RnmxUu+ggPkGWudPaquMjYfrz7+FwEdKq/S+NErH
wDp8nFDBJmUyxb7Kk00o4degghqAaIZj8FL/Hl5U8+TY+lpIs5ZGhzLIW/mh9eAuVVs6mew2tgq4
EW98NqT/kPBO6ayLBo0crbamPYGRhEAnj7njfUP1rcxR82CLhaofetCZ5myHs8z+wrvIxCPfVDSf
iC/nDlJtbIDrB4aUFxE5J671BNoNl7cxBvLAuqwyHE4af21oEMnuFD+1sYTWBAfFTI2BD8I0sptV
qCw/stgeqGP+/decDB/kGwHpQHVumIcc1KQ5UYKRnj65DY0R8duP5Q1Z0g0Gk9XuWrcJ+lvpzwkE
1DftWgUTVpasXdOEomehPMQV+Y2NqQpJaCQ+UZUKKQc3wqg7W5h88XHORNeinqTh3Ndg6FtJ3UoS
crxqTGncFBY5BkAo0IbEsNrX0LVhTs87zpZvIFmfCkfN/rmknmCba6wRRsA06Mxh1IXb4XIN3dLM
40SFXIx9Zt2ee+s1m4xysV712kdz7bwUjvfpY2a58Najimh7mjZsI9dgqqXcFnuhn6CSZC0wl1tm
jaXDo4XiC9RId41rCQiHQcYr/xoc3UNb49RRfusGHqiQnntX90PoH/Vg9lK/UDp+rv/cFQYPh5A+
eb/Phy1GPCZ1YuTZo2khq9aKnzWZIrjfiAQtQ5qbmXY18N6wBTLI2dFc3F8Bpa/GGy385yc1++6K
fhBLqL62MI+TUOOUYIkooWJRugIFiAQ4gxiXTeDoTWv9AePjU6ofptPUGVv9Dg6p3xdd2Uc2bYw1
n1fm6Cyab6IbZZw1Wzgol324RKE18j49vFUUQY8rVvXmBCmzaZ8FbPi4fhI1pbleyt/i/u6a/Sp1
0VkBNCARYtWe4TM3GxSf7kwrFRkRDxLDYsZmEJT43usr2XkzjCcgop5kEDXu5fYfBoxtrJ9wRJk3
f4hn387+bXYE0XmrjyxM/uXa+J1dDrFkp4euxjk/7bXjMATuRx+CdxtJY5I1mx5z2brRT1vwoWzz
4aS5Lp8X/YPrcFvnvO9yBsOn6dDUPiACFgffcggzLVBQYNkEuhHCjHPhiRu7kFXfnw21426gY/oi
lcSIW6KFLk3jSleRKY3Ja0RZSeWAWYVSAe1vKn3X4MZBE1W7J7m0sFiaRDKBDsP57Nzbx0WBa5Pf
cXPfzP154+dMpQa4CEGmfGf1GAnwE9RPn2WXtzG48X5CCXmOi+iyWWoSJqK53/ClrTh3fVXrIi6y
JOovnP2yo5XYvnPYlzvvR+O2u8tq88jFxZx3XJr1lhct/iRr8B53UBCWKH9dYKjmSSc0IPEfbg/3
+MF7mR4Gi3Zws/yaOyd3+Kdj3O63EESEHKCft0K9nfAuB5iJaI1yMX+jrm4v1ApkO7eO5E9NqvOh
GD5e7cxKwftsaZVMPZOKUN0kSpwzeUoMIrb8a809WitjvlrEfg60HnFk6YAzHaIOTEFNVeCiCzPI
X86nfnEmoQ+EGiLHu3bMrtrmh8KNS0Hp+KP4poSyJ1iCGZ8dymvZGpdswnFo/3HFUG5KQx61j4cI
AEpzJcfD3uffpx8wQ6CUTIGYEVXFIVd4QEkdAC1qrQGdOpzdxbQVVw8ZooDZ9gVd9S0+rMYsBZcw
c8XXnxy9bc75YL7G+pgKA+6yeQE5x5wmcxVoutjivlZMz+52fFldrwnfeCvaXCMuqdq3pFeEsk2d
cILOWkVEthy4K3PVCcfkJIB5i3SVSu8toyBWc6yd7gFkExwXleeUfGSzdlwD4UqzXCNp/IiX0/QG
i0vvoA4NYtc/H8yMJleBYBljNoEfmmOgTnqU7FnlPgMwsXJWobWMY5MQnFGtVlBlLMJoGfieBfO8
yw3wPoWmhHplTzYYVeLyx3vqGzMF5AJw/eDjegi1O5WVnUUWtYMf2qbokB25Lw05R5E++vwIVaB1
kNU3z3rTUU1l0wjI/6rhd+qG1ng4yvOYSdPwHIA9uoyGnZqaUgxjHSFmHTaia3d2AQGUfwoakTrL
G6ZEsTgBdUQ6QyZVm9fejcZo5OYfRZaskDhvesLJ6fi3ZTRY2qIyRgyoGmlhPS564tSXkUo1g4Az
1IM8/W6oC3Gj3bcFXJ3VM2PPKDCFeeGfRtVhy3o8eS6m7TAuJvHGV5vhE2drUw9QKQON6XGEirEO
4H4d9Sp7+L9+/20bwhWjwko8blolc+0LNKf5OgMVcRHDAOXVfKFN/H5jEvs1/LN1FWx0zxRTDJkZ
stDZZVIrAfo4GGrckpjt8YUq+CnABghnE4nrATwSUFjz4fZK3PAny9xHkDoYnmlbUku7/VFpBHxe
0QJf6o4VlqW9efn4dm32WHj3tbXZASnGJep5zKmYkWqtfMz3D13+IAOFW2woEHGPVEoiwz+GSwL0
MEogLWGSgjzcLpWHKp8/zWHpal3UN+UG+Fvh71fC7XHjftbXTAbo0NutmAFdC+rn4oy9CMGKaYdw
es2XF7GZwWeCIcuXhrBhHjnDBAlo/UMOSjLwZ1FI2HE8Y0bozjFjgiEWK+odu8Axpuurpuhjssq7
dfUWnPFv4Hw8S4E3/ZhmSu4k7mITi+jPyoBr8X4dOR/IlF620YvLetAN5qD8ce6w9ocyW7eBIgE3
mditfep+TZhnpvR4sMQJNdrzJCmyNXYsVnQDBJx14lp8aGhVApy2CgJAFW+6xdqk50gUTxsoSlgP
x+bFr49omr5/rze+fUtcK8yMHwxybfkmMQTpIDq0tsNfnerBHATSVC8Wkf5CQAoKVA8UHvKrys4c
tx+WXNhvG0rZK4xbeIMbD7PCnDfAMAJIRNZEf+3QXLkYTu1q2rUiRNxBayqd+7nmy164Hp7aY+AU
H/FbhY7QT6MRloCiwXHR7SIHH858w8lH/FN8VW0XPvbT30WpLHu/kG9Almd0XV569Co7shj3QJ8T
AANsLFbyN8kXrpQ2AjmwpHUgYBSEtDZX20jp08GR6S1xbwYrORk2MXIFQYZtkFYcSTdplhHrngmG
REuvxyJCv/jFGMenkcNP18F8TiuBUgnXbjBMi+Ao8uyuwrOLBIxE9rk/pYUHCtiY5r/hPir70MA8
Csndw0tKWG2HlXIXJ+EPGFXeKtNmr8bRoO62ptcaqid3NIMBtNfJFzSbxztLFRZLzkZPbSXgqKmh
MUUHRqFHDr7zJRXUW5S4J2tPyv42YiY/hL5vm+8O8OzIaDN9wBgXqlBAlrti4kmAb+KgVlbqzz8l
/qfli9EnaVLLFz9GLgSP/lv6yuKxNCHpuqQNDxH1iNm0Z/IeOW1Xlsbt0DNyHJ3pZM4EUJADyQ+t
1jWPBzARdUUO+wZrtSX+IQlHfcj381sQYuO70452G4e+swcGPxt0ih42SMHhjpyUvGnue0y3zDPz
i7Hxd0MOhasIQ7UZU7Y2bgzIfyA82oIaL5nCtv0kVx0l4Z/VpBnC7U5HBcfILkhLR55sYVXNo7XK
0YhW/lgrwSTwCb0bLeb7ECcsF3i9375VH+NyuqsARpdtMQwIjGwS5D73HgvMOPB5lb0POMZUeJI5
XBhta0Yv5gOTN1tSC4PQXDHlxfiJMfvqymOvUB9qUx+Aln5BHd84QdDrP+E4yEqGX3/qrXq9cjzg
xGJsuF1Jgy0R1ZRwztVnYDxnUILOBfUWVaqcZCFUWqOO1ST+KwVlF9DIgcSj988rjxRd0B9TNHJt
WNJQrwEEygr+0GvdPMbRFctZpwXAbkoKJlge0Gj2BgYw6xLsEQI893br7wVWHVVIIOIbeuBnbGk4
6QFUjdgvPKEy/dHe9sYAWtORs4y38rntWBV2HdWQGp7UdN5hEE+Ofh0xFWVxvNopMiEHMOjatbLW
cLrNukllI+3NFeK5sB8eJJLety7cgi/wbarKkVD7BYd5viTvrB4j+Q5ZzLtAV3cKGIMlIJcgFzFJ
8YpNgxUZnRNbiW41pu3hQG96zgEMB8Q1XFGfFFvYOJ03Shnrphxhg+Nku2jNfd2sJ0lMy9QxSfKw
QPqd0yBJGkIBCJML7akfd1GXrG5Wkfnfa7TA38WA2jiL8UpNhXx5QmlGdIJfzbrdmXQ3Gak/d9IU
sUjW1MvXxxILYSyfmiUsZfe3GjfXhnto1wXcRO8ZzqspWlIxCiV1LFoepsjJMRV7Cuqc/lO4f4UH
RHq7CJxsPAjXvoOTHcv9FvtU4Ul+bnZIQcbhnntp0k5UOQFH2x2UYKVJr7KaE1MKFXSIRdgJMwAv
unijuM/kISSbYH2wNtBBPs+cZDqGoa2Pu7i/TeRDT8ULV5ODNcMJ7SQabox3GDapbvcGKwYXPk/5
yfDdpEp8JNPe0FlOlrS3Ajz5YGXKlbAUgK6WuHkrJNLtz1Ll6MYUO+2qv0Vhgf8oS8+LmZD36ONs
KAxqflJ43qgJF2WIbSf+LsWb7c47//6AHEegHDcIw2vAp1XKhpS7KHc0LPMUXCxJ20dN7ZAwnvER
hQRw96phPQOn9eidUxxtywwkLvXpEUXFgvheBxDF20+eZtZWzcidWYjOyE8Rl1Ps5RIJZ3KkDceg
X3pjNwia4w0V9HhoCVuU5CZ6mNWeZEoAIa1B8dhHtPAnHlGXXOzld0/FEQfHJogsX73MkcbVxjuz
4/UAjwvbazuE7xW6Z9NUlBnmofN8QG2AlqJQGVqOnPHqGktq5yqUZqpvKOkSyurHz+hgptQ74wF5
WK4ls5nPzID6fdPuvLfOiwAwXPuaAZcp/4mEJi1ZYL24K3IHZWXWqPLjbNizTwcw4DIU5NIQ5v+T
EBneg0Y+Nqj2H3WkrvnXrRYghk0YMi20w9kYChPyI/dl5T8qZ9CZRSD6zfG4ExLe9S/UqREGG7qs
fjJS5P1E4k9PjkhHCHoBIEfwElbd74Qgnz8NiqZlTRoU3teIz+kq00qkU1JbP+lPF+FnK9cU1++t
El+pOD1yibaQtmdvBzuINGbGOV+37GubCdJDycudJcavbZZ0fJDZjspXsc/ZxRKB0rDgCSmCnpkA
iapYVdVYFN/sp3vbWR+bRulBLlFfq+QG8pME1bG5ZUbVldk1xyDn/FTiJThsgA12w1MNu9imeFIX
ZkrzfrCvcRDHGCSEo/q4sbt89R4ctG8krpxZBnNOP1f6p8jZ6eSF1VdwvumVNHjJtGqOayGwIG3B
eggn8B+uY/9Bh73wU1R3Xr8mN1bYMWMUK1QLnJF8hA8wv+H7L740Bjm+ESinTOXiONkmlBiapxYW
iyvpzg2nhXaPBfa1fvUrWlqgSUt0NYPgsgO8EpK7HBZYcQ8xA8rx67beYyoT6E0XkK6l4wXLuvKC
TOgY7LZtJt4onEm6gnEzqY9raRlhCeyjgW8ed/tmf3Zeymvd4FnZmpJIEsN1PtDJ05RbiF/ezfqp
LVKlQAfa0O9/hFkTxFvbpvx/yslU5PFKnpDkux9+YTBGRD5jxNrJQOtak9LTrjYKhF+6NBUO+us1
ByqgCAfJ71+EVvupwlEiRnPC9EalKjb/7N+q68wjcN3duXZbAMKpLaQUxDWzGa45g7xf5+RP70yA
09RFd4Cjopzo0og+KrVvnVmSp7tYy8GZpuhfSMLmjG44rsY5MAk/01xGkxEkKq6R5zboM5xy8o19
+QYm5XR3r3wwVlhOLZkNlz6p2xyCaLJLK7K51r46+kBQx93YzThsH81NAhZAOr7HGZi9ictgUz7l
iR+WPs2Ub26o94XpyXDcD8S8OSM23WZvKj9VwPpgVWsaw61F1xz1TzZ88ymDNZ2qYvHcqqxkhSfs
R4U88u9Fi9/9RXDu2PxPliH7xcYxxYRRSQsJ8BffLmMYHmugQgj0gnv76EvOfray0nLbTKk5nW6W
kEg25nFmGtYxAdopXg0TQCKCy5y3647DA8dtRJSXBhJF4UNJgC1RPPAs79k4hQjT+j1Q81sqZFqh
sHAwE8xsZgwg1IcDSHxiPx1LIVfUZrQor+hK7YUDEnDrhlwmyROfKvxfszpi88ftnS8oksVk9nG4
azRK7od7coOpCBGyc/8ejF4F7MiKSjnBZmEdA4+8Nh9kClxVw7mk3YJGgJ/tn0XUtMwA9OHBmXh9
siba40PmDuDiEtAqOHVwuv9wMFPL7CCZj5dfU6PIWxKHalncwXdT6ASgWQbg0/AWvuBdDQL1Ths1
Fs4wVOCQm3x4Wj5dLNoZ6gbzz96h6RtmfUvgonbxjBZBRXwueTT6fZ6duS8kOLSNnYwLEL+6iY8U
WKZ8lPtH032Syp+JS8mjZLiD4gYRVWSnSnkvZ5v3Z4mFCBqwCBAvNSq7UmuSDOnKKtLA//OofAxW
xHqUeGKiH7ncT4GbJ20VzJHBdhmlAT5wS8LPAK8eaDkBYNh8L1TkUDLKVRtY0U8D3NBhBUZ14f8p
fwcG1SrjcVYJ2GQdCay0MighdDvltmk1QvQqh3Gli13w15vFtld2Aov1DmsyilmwrPTF3N9gVyML
Va7DzIZrz0qDA4g4PzRaWTaFd/zgOEi+xIGUApqGYNGv8LuDWOXBQpxmVNyzUKivFOzfkH4FS5U2
6Cg8e5KcqDI9PS3j44Twm3VXAOcBWtV4unbxstp2PF4601mMuKJFMpxfKRqh7u61XUYJW/bCe+b2
30iHtUx2nSgX9Ul0rBa+XSWhltVSca+5W0qyORHkqaPptpMwgRlvisq3Q5nB892jqkxVnYV+eVlr
DPawAUxZddZushBe1k2G8RnoRtip7/7/q73qHWQgVoOAnZjuENvtu1LH06uBEbh4ks+VWvrPgXea
OQxdwEV9NhVv7JecGhsG3YGMeUCLHb+0ct7CIJPlaFC8DNZcmLuYcnDE6pLPoBPjKJtX9Wm69iU5
FsHeN5TjZNmc6RZ5CZ+piC4YMZbwn7ihAIlZeSVP11r9XM5BrYmpUuJw2CLr3R8zK08wdxoErnJ1
wRkpZsQyCkD9c9hZiHIAzzhxO3Evr1btdHN3pGg/65GS/67jgfc7zBRUFwuJJSVRGkQcS5lXqz8i
sjaB3rUj8pc/CBQgeXAO0anVe8YQcVN1vFdQGG84GcSYuMKi2OmUG+6ArmMp+/l7VUhZ+oO8817L
I3+Af8rLlDQH2m2h9rL2eVt4kEYR68y5kr9PEKlLQC3eubxx5jl4Wb2/SnNqGwK6cNXJtb3AGefI
cgYP6uxcGqbt0r0aRs1jlJwWLRzzM40JPq8McjNNIYrsbCikBtmzRyCrZIx3Pu9Q0dy3H5EMUsAk
T/U1/hxTQAB0nDYcD/NheOMz2sGC47F2NIm8ZUZSEbIKCZs1E4zVhs01dqmCMcZChb5beWy3Hb65
yxNFDhsLb6+aSmCYLaUZOZQQ9xAhNV691pmALe/geoAPa+1B+BDIR9c1K6VSejG3i8namG/ktmWV
yE8wU5c3PT8e3yU32iHtsXVvI9o3uCMS6nlmDFt90Qu7YTZWQIbGJZ0xC4eOZ0K92rdPknGq/2X0
I9i/NuWnJXfJxwr3A7hNPyIPZ+O3tFeJrXb5t33YyQFQv6FXW9L54WKyn7ub2ttb1d3fZSfBKqRE
+pugDU5nkJuSA6EO9EYQEaWBkRUO1mkoaPRYtgulaXe8VT+ZPwvmGURaNRyv72rF75Z1Qh9+QBKd
pmrm2NZ6Nl19jFXmYu1IWQE5cEizsWAY1NoxtjyqMTXndcdHbHdTF9hWcMAL+EFwUiOgZHfDGWqo
VvfGE98WRT0z5MQ1f3qPy2i1HS+HIYRo8pFt7Wwl2pQjNIrmEzI7gTHiBE8tboON4ZTicsUP0QwK
uNZF3MhwbMyV4LESMlvIERwpkBWYKbsvbs/bdqAFgVL2akCiA+krHjHilZMI2QMPIhlwf4JYStNI
eFgnUVlp7NAs8IcLGxTnKNR+0CTsE5+zT2EOEoAv6L5v4uveFt0e7ICPcOXz3j2/uCYWzlBnGDKn
dN8ma4z9Ku+yDlyNlfwUzs/ib6ai/OzZOVxP8nsX+rwwG1kRiilYNuPzUcBwfYRMg9W3oofyo9M1
QloQVSKWIdG8grTCwt0etTPxlv/STMdOJHZNuXLPWkfiMwOLpiAOMoni8tZ4ZCJo/Z7UPq5Froj5
jhT1lcv9YUpE9zOK/SlWJIIAzn5AeAeDSq3L0xIR0SzL4fznz7cGXmOCju9Z5pd+MRmPL4MVs+Do
jg6dgZxBDiagKbEx2Qv3AzEC1YAJajU+6kEdzcySBHobWs2NP5dtOng2G2wk1fMtChyQff7lPcip
megUquIi2KKj2eEy1wQAofwDc2/m0QDzv9bIqjMADyThFbQcZv3aZiHCFF7nw0ZfYiJgxZAaHBvP
SKc+ABfoQQiT+lPrjOgsAlA4h2ScgA2WEO0WDkkr4zdWxmw4Z9lFad5e3Q1oOzs67GSCeJh5m4jC
Cn7k4x3GnVDWzP3Sd29SUYC9vu5mV1I4Icj311eF6NQcaEF/oh8DLY7Zg3kp9DJwZCrgVWhnvgcl
i0d+Ospb1Z61Uv60K04iWBxsnUarU3aAAxJ/4IldlEtrUqI7fc/6X0h5nFJ9XZFe8wixaNk71ZNI
lglO4QsLoUQoxf5Apq7J+K9p28gwE2OqviDG8FViOW0IbCbrywMwoFl3lOwLhoxykKpcvsdyeL5L
yfPuRT2WuHL/oGrU7rPzKF/kas+BbNrfXgldWhBg6OJglQiCBxyANamKkMt0MZl1wrYJbxeCKALd
/fpKq72SbCmJ5Rh2XJXrh4cQNQdS+MUyjb9HQg0EOd0Cg+8DhK4P/XenugNrGH7WfhBNE6cOqBzf
ZAyxNMOcquPjbpZdCYrLa6+MhTRmKNFFKMOggEQ17ApSdFdgbv3FZy8AzmudjHGe5AqUOtCGQUcI
BXNWPQibAnM7DGZAsShv3f29vnDz3GEt5Fyu0iqwtI5Lat/1NaR3db9gl90BDlxAM4lcq4uiYgLV
c+KPVpuXKvumfjJjz8arsYE1ymW4abTstKnkIpXlYWd/M/Lv2HNnjviJ1Ucj5av4hmsisaQV8flX
lWBjzz3vvoo3tmeZBlmN92fr4xtcY1qXSAmQ8B3PUZvZa45XN1mo18OiKX6cCYDKSf09GLwo1QqA
m86+aDlRR6fKMpzbSAiSPkG0bi7tzcxWAv146Kx+W2UomdMPsMXKKpaefknMhXwRDYA60JvoTsAr
e7ah+W3gQ+HaLqm9wqr0c6cqau9/lHvZKeYbnPfvnl95tzI9HS6wX5AveYLxxtOOS7yIszAZYdI6
yov1QICvfWPc8MWKXvRQi+cllsoyj+E07ESufA8UMwnOtd6sLX/+b1NeZmiLLgnacJOR6ejli1P9
50I/kaBALHw+F8DdmWB2O0jUkIWsdiB/LYqefweHeij7RsUtqehql247F8Gld4l5sK345aXYj8zP
XHXTef/MtoV8yy8UdxZLK3kpI8yRGtcSMOhLrzm25tRXunkvuUui3t/KDu7G0hPEAFevIZImtVrA
Vq7S3emkDxs6YEVi3zLj7n51A7ifsHbAZsG5cRDTt3WyqzYUkOkzE9L50rvvPV5HMq/I4M1NNlYE
tiB17BhmbcvA+sGz55LvggjROve0wARidp7AN7JNgDiUN3rwzpIz4eXaulVmMJq1EC1XSB8O7rcE
TAmNZhj+nm0Z2QlPDSncRh6VSFANUbngmaH5jadwKgh+2XUh3/TbktR1YLze9HTJvtyYwWA3gETs
vB+gL24QpY3+M+pxdQgm57RVC1wCc7UUMX29EnSqrjGZHHIKa7FWQv8D/3y+O7CfkDj71KrTkWw0
F9HqmZCOWWm/z3JkXWFLZjiR4wZvigtJlmWuSxdE3yyyVKKvn615DQ3GL/yHwpFEtTb1qvcM+w6x
Y6JOxGzojad+vccxNWmL0+v4ivck7Ptr5LliAogcAJHtef/7iOzCgxecaFmb2M4eqtsjh/xMDVhR
ufA6xhsfrWUYHBMds8hrQJ6c9ZKd7jnqp/x6kkBqR2f7/tH1JmKULapLVHHMIHgQnyxypNK+0z5F
G10cJT0iZ+V+BAJMnuHKiPSiOwI/VQR99LtvHOLBoAkESMpI9cQTsciUoy/APXef9kXFVKojBc4D
E3TElRc7T+n8fHoPzm3bL/XhBCiCaydIRyjQnuzdLEHN1OiLze9EcqZVjKa+Lcf7J+X0vaOIls8l
RMhPdFrpZkr5LiROiXH9QB9u0lcDuV1W2Z3OEtvKFqut/2F2vHBlgzgLjIvWJfhdLmv+t/xaWL/J
y1YxE6ra6MdbG+mbqCqAtCPBRXhgVLpuaM60KfBPDjCCSgAr4X+ZTg4/hwHX0toXF5SJal+V4Mrx
QdcgKvVAJmbo9deMxUv/Onww1eVwse/kpGv6xP4i6xHpWhYhfq68nIP9tKckQsjlia4KtmV8o7K3
2thidTrY9WNpIc/Fs3y9WGulSmH7SBw0uC1SgJ7bOXolnfivoC4LEvIIueO0JoODxuZTgp+USB8M
hnVmiu43mSJxetRZ3fvXL6kgSph3OAoJ8QACspA9mPS0mLx+ionFUpcpu9qkNa/MD4bM6RLmQfu1
AuLY0wxnm/Rok9/OS3G/mH8q3UO1GFKFGtc/jibp/b11zhAYVha7+hT3tewvQnIBO0xKbBU1gh/o
9T21x4ECfvD6X3ssY968M+0LVdeQzWSTznDwA6btN5f2Sj0lflvDyFxeHSaYBaQG2SO0dX7mj1bk
n7ihTXYOI8LSwGWTD2mFtfDrEo9giCRb+TcOea4Oji3OYklPZ0TP2hS/dEFAb7h7smjlDJtuuiw9
M3LF3GrKifRmdJtbYyQKdfYvWXCsYLrvWgdfoZfCN58D6PazKJYxBbtn/rDmBqcZB9UkJHYM+QyD
yc0RQC1YIGyXJNQQCrQqNB7cc3ozOoWWGypLxOnesKOE3Bir8JtxNo5iv8MLNXcf/dwisJPmIQvH
1wkX4zjNEt3r+Jeh5qd21lWcjnSu0a8I5lz1V2HNU3wap6iPUfbPdc0NWRbDHqA9ExlOrkkcRvrS
5DxUN6dPB/bGi1Qp/91T8Voged+Gsee2TNOnRKnY4h0rN0lST6Y540Fi3D05EHF3j7UgoyFZBv0w
GqQCzLpHFOwmcrZbp9IqAMidVrleixqHhjySCo1yRPXwH+Ez9nuVhmK9smn5ibANagJeF8WZU4ru
EPFBR0kF+C1uVsGbyPFSRtd4Q+uA7n5q7lQ9Ky0eP7xqUHFV2WQYcWEuoC7g3nVVGQgXwFvPAw6u
MUyPAoZmoxSjGmUnPNO5esjvOocGXv/MTxllBDteSiONQO9nVquuy5aUkWn/Y4yUDJJZdpnlarAb
gb8UC9SuzHixtsd5hnuYcT9lIXFoDT9fC7g3nhebZG3u6tsWDsfNYvd7+lBmfZUBh/iqV/DP1f5C
PmBcG0vQ+9jJIdTUWu44/Z+kPKGym39pedWmQlZP/fA80jJLQyu1Zk7j83Bk+6o1CItbw2lKo2Nz
zrPE7pw0LRcIRxwZPXUmaR+AFnZ5BXtAzGaZPqokD92MMHFF4UUuonPF2KqbW6VaIZy/5WszMCcb
bpQE7ozh2dIJd5hXcnP/z6XyAb08canycDKwiAyZ2fJTLfcSLTYIBAG4AfN64GVKBl5Uo7hFDVnq
vorsa90+6cqahJiPldNE6jpKvFiYY4Mn823uGC8B/yd55cD79hijkOdv5sQMqeK8K0zfrOeq8DDX
y0UeFt6tr6L1Ka5if7w2WP1YfWF7hwrZfglqUS6axVVwl7CI7deeAj23APjgwKYkyVHwo50Kpk/0
d/2mEmOAIE/PHMo3qU4fdJNHvRk80yBiwSpU6JyMo3GdDmV1LDdVWINSSb9xQ4lgJ5D/0Cu4rxRw
V4Fc+ivGo/I/v9ntagoSpEQ7k+YaPzjlmvH+FT/AcOkcC5/l8kBYScepG0+b7hGyIS3qou4/aOgq
s/7Gr2s7E2YyM1f/XGfMmdSzHXw6v7Vd7N8w+4ugefGIVPHyX5iRB+ip+uDwZpjlCkuq6j3JWhWU
ZENaLIuUiduKHS0E+VF2JFojqq3tdB4H7L0jHYyjINkFHP2i942Fk9cyd/Pw+UioyIQFbKN93vlL
UiaqnN0ZVMS0kC8xaz41znTIa0CoIW3KVFYISHKm2X0rJcdkwrt4BSmgVuZ2ydr90V3X9dsVM6Lm
5cHjOyJk3NaIRadwDVPBJ7lYAK1eMjiXyIXUhUU/aviMr6pwzHO+ubI+ywrj08XU4UHewssQDu22
pyVl6pj/A3m+D5r1dEzzakRlBqPHq0WOBxlWrgyLgvG/PAylMY5mfyPShadHbWci745mmJ5FxRVx
v0j+aosPu4SdiPgAwX8UbM4y7DoYDHmATmrrjlMfDUfOjh3m8g0zt9r0Ikq/QXosgs44doDTD7Ek
+DyD1Eqbh48eKx9mF5qETlg2evRvSDfWaMdrjqsK3EcluOIf+bSi1qy3bM4tlA65FUsLvefdhI4i
J7mYAuSNDXBoYutJAnWIjWlQRNt5baOPy8r8ln3hoBq5jnD+6EW1+A6rj4y3hbrT0f0r7S3gNf6h
NCeohDtOFah/nxEnE3MgBM5rEFWew1kgQGQXUD118XOEV6Qxqn/jg9Yf4ygXU0WXhAVHdwo6PciO
1pFflW+6MLhvDzNOJgkdw1zStUY1GpkQCJcTV/CHxw2B+bx/Jn+h36c45O4qtOUnCfWdg89H0xdW
LMMab7blL5Bbrd/7ZhgYAzm44TsLiaPWf3cjkg62kMYCCcXIpIoJrW+ITE+zoioMlNxYZzmxArzN
IFvh3aE7SE3fiB0fbUEwvul4nqUcaOAJObM7djcdmXQJrYtgy3f7eUs+WvEWIg6EROwkMnLCq6gL
kbmTpIdCou/onDSRnILXGPM+AABTkI+k2mQO5+mFBpwKihhlKZVBXEBRCv6iKMY04tzdA1NYFYy/
ABzbY66HYBxwB9rHt/PCCFsFkCCJ2SX8YgIlybBRDPzO3bV9b5nhqp+eNPrzc95vFZO0c2VqNa43
Vm8B7Tji4zv6PQydlusREn21X87Fsda4A8marUrJWePgKMynpRhWp7rA3q2pDTmERiTFpZw1Qt+F
r9YneSQ9ON2Yfx9Ew7KXzpO4mNXibFGWfzNB9oOFDf43i7xqLVQ1eXNuGeIRi1XimJnG0QXfHcLt
lHasAag2Ll5c0WX9zQ6qr7B9y83ecKSt6s5/FYUctt5SdmuQy41RVEhJZLh1cuOnUo2Qp91TmwU3
zFhD5/RtFBhlOiKbbZGGGS11jk3SXrvn07+ApquBq0pyLvlRylz0FvaKjrQAjvzhv3Di3YteU7W0
wTqyKgSpuC1cCJVWnmlkRrU7iLb/gWKkJz+PSP/SmHmgy1QjKjmlzhN+UKm9kI8Hrk4ax1psVqiL
SAkiDbT0w3D13SSIeFhGSfX00J6XWcEnafe+6b+2HR3yv0JiVkiZy5UEKiVsWkYWaSCbBP5/59mP
MRVjmAniCm/uZFOjNpGuomd4a0KJjnUDVMug0Ps0wuVdixHcYt2aXe9XelwqLICEbucA+ZvMaxSC
BTX0j5rwCZPPzfTJFH46QfeR/6thxZpfVDIXfHi6E8+pwkAtjJDf4CKD9lzo6KfSUunq3vHwjeqT
c31hf5gN1fa8dLwWX7OCjzI7OtSRZmgGNhmWo2lGuQL48pEmkpOk0SHwXoWEm9tH+xyVYFjG3woa
26PdNx4OlKOnPoLMdGHh9m9ScYF9eC22hvpxNtgSomNCo/1ihUqN/geJdEnYHcSVuwCmnBM9im0E
TxPR5iSxEhOPUokIPBpIh6VHLbn3oGPnf5Q5jspQkDKtzHWjefpkUqn5JCqIXqLw3S3Zfvsqg4Ps
/SvvTxLtvcePxaOoMuB0XWe6pTUFDHSKBxAsaiPkjNINQhbhNRRGE+sVzp5yheQ2VIsgNUP1ZmL9
4P8KoL4Rm2Zo3ceIzPA3v91S75Gr09RNny31a7W79WaobPQqMJ7CvHUtxMvkuaklfaF7BkgqWJnF
2DroKJPa6QV5azNYA5bVRAvJnQek8q5EbGtYe5uvldVcLUBWWE229ONv52/8Wx9FPPmFjD7ht3UN
rgBMhXWZoamr9YUZLISBK9LiT+lenQJp2mLP4spgMsLhyT6mVbkGbgu5ddV4b3Zz0isk0cJFIPK0
UMt/NzL3aiHhkv2TIH5bRooiNo7/ou9BmBv4hxarRd+Slnn37392MGmAAkjI9kLSSs93GVhcWxMI
AmFnl7/2n0clVOy6G8dqUZ5AxQyjRo51tf6rXy0wy5ER/dUmaOOmY3LkIvXbJ6ga7xaKHhQU5o8k
vIHnmqCZyXC2/GZ9TjI1UAzqTD6DnV9NWLboa9o9K5RUPHY8qAZKFcD3mhlBqHhiI0gz7fObzoTf
Op3N25nXDBk/YLBkf3wWk02m1WuWdyfiwurl2Au1+kuvfMTXiAHyDe341ZSnjH+zT/BOCPaMTrur
nRNkdBkllk+dDmd8WewwGZ4KDD2HvKUE9tBqPc2wp2Qzy00VgZKPwqAwfMSZ7nWfWb/nvkS25Bff
peBQE6+2jiQpghkYOuHbKJK0X/g3fHrexFXaucTJZ6Rz6XNcvk3FM1g9aWMdSRfceUQBczuiSpbA
VY17/niSx6t1q4S2mn50cbQ9GHDwPsJzt+VBWpXXdTyCyGym6sVPJ/EhehIPa1TkfxNvcvmLW6Ea
RmWWRTrUlYeZz9j8fIw5/Zpom8jHxitxGV9O2kdBvPLpmuAAymWLU/RtJ+HgLiloHqPdrrBkOpbp
Y44NdzqcVOS7xZIP2l/pwVT93Oz79SEH10Mzy549b1zbEdiWl0INew3kbeTJtRfgtdk6v0SIHjhO
4lPOz+V780JiZ1vCeKkc5POCt8j7zyPmn2g12EXvW2Oa8LtjQ53WkjIzKr2WGQ3lkfWAU2AfZBA4
gHNkLhm5rjvh3Vfda9fmdDZdANjpb1lHS+TnJSq4W5/VQz/lZghMHImH1bd12bk8A62bHno+V2dT
URtHcdIGSxYsC6/EAUZty+aiyUDc154T89vURnV1JUeUXuVm+htPvwwXNlH1hwa+C1sgxyWYCi5G
IX9YpGByMihzJoieYe8+135NQODnEempALfEEp4e26vvUMEX1Qgn4mxGhb2n7JKDErjIRXvRVYQA
K8y3tyS+AFDCUMutcpVx8XaOt5jKex6fQ8GPZU3T5Nh1jBe09SrxQPbNzewQ8M4SS4x6YXyg+s01
0QqqOXiYT0hvQm+F7QTndcFlEe7n9hkPYoStc1Ce5TFs7oLCn/w1Fg3kMQ1poBPFer5b3DYvoEuc
W+5Nqt4gE3IjDnFlJ0YCXIWJNzsGSnXlw1RwixYAWfm34xj9lQHVow5N/M7zWmhtNQYiGp/+Jb6u
H9FOGq+oU8LL5YO1gq6SMumAEj/ufR7eU0UVbuAvpfeITd5iCFizl0NHPD3cgyP7Ne4g7RXDeeg+
pk6RrFVNN/DkRg3Mq+MqCDYoOkLGyT3U20EY91L5olcAHqbwxKWhRybfBmopVUbFrrkaj76Ef5rE
hN9KSw6MZG0kMWDehJ/VCw6DG8aSTUwu30IJ1TWlpP90UQQV+6cS5+2RObkQqs926QvkbOSmi8oT
gcFExVHEaiibXpb231Y70Uz1vZEZ+rVW1QNRMOVvojfU+LKG+dRW6LrxpwKRjvrv2fAsQ0GsvduQ
Ds3L7Ic1D2VebbyDwehR474gQd6/xmvLYB/aR8bHth61L6TxIm26UTf1VIJE4KMGr2i1EOeEqTAV
gAw+3RZ7GdQzhvUZ7AzCSZ8FUlqiRmZAZhISrcKE1rrPsHpn0itYF8FiXFhxLEzn8DCtTN6+6plh
Qo5fp1sk3R72/PnJ5eLGfSJi0l9riWw5xgUb0r43A+M9IIPEM1KqKI6x1h1lEOw/qNGe2U8PBEcq
Jljb8zhJN3VT1G8gKS2zFvhzpILr9ZD8tmCdl3oNPs7tzt3/c3DFcW9NbPYMSyHj6OcEkc69j7DQ
ZfELmbQ1ESfnEPm45gKRrk1mQeVo+sPlOmlOfKDHUFPyDNn+78vnn7oNn+DwVNykbZd0s/bGChI0
7vrBFB7nrkmRV7REJOTjvFH8jA+hrxpr9IvH4FXLHxZsqxBlwk9200lsYbZFHCRSZlqdzX1tKDGk
VUl3i2pj7HvMveRkzxLhFwvg3pixRm2GRVySPOq9IK5oFgKpFpT0rUyOEJksixGukWB/yIF4Vh0p
RtnEtIbfyxFwylLTKYyTtg2x8TUwI37WqmtSpGTWHOBEG0B3aCNPCGNPXYwasikNSTVkaX8V20mb
htElZZc0vh3qL/cUJLWdg2gB3Nrjk4JZnvvKbJyiz64yLUoO1RQ+P2NFPW/AEC9jUilWF6sF+0eG
O6w/RQilI5Uad0zaRF9IhZkMMWsSCa9TiaZoQcnnJBpoDyGFezYShu3EoaVZGm7Y0eIQ844Tjjgr
BNffoKX4xj0HCcH3Hg1sZALRz6JuU+X3hynWDdWfyMFMlId9uagpo+UqpSU3bZq8fl5CcuUx09hm
rLsdyliIUCK8AYG0nAmQwVcFQVGFX5idI7/iwxamEjTr7uFVDADN5ZOCIApMr7Bsuyl+8/WV2OBh
TfTcha5EF2CQlcJ4xuMQuz5uGdHaAwD0H2IQi1LWK8f6FadpNAIJt8ekQulAtD0pUKvp8gZ+OaBp
dhVyMoF8/oRz7Y2zCZxafXYAhuXeNhfaO+WXW2pxu3s+lVGRHLcryoOydpLGdYLVUEN0XYYV3SCP
QXKbwESJZwGwkyU/V/8TNpRtPiA9YbSwP+MkVpulMR8EfuS4fGXPoHWTE6DXICqXJAqRp4p4YboC
dUjaMx+/Etj1t18jWH8qoveTipJXghFlmcUp81B1BPoWCw+Zr3jRk1XXyvKTxYlkp0P96VlwxsBQ
9lMt1eiRE9UhLZ7yWJTvsnmT6+iWT/H/IrBEFj67GJm+g9+NWsSn+P3ek6zQZ1YLaMMit9fAePTI
GUZI6taYIpMk45sqfAx1gIOfSo9Pt0Oupgy/I8DoIulRqZUu+LsleP6rrs0unQudiM34GziX6Ats
IVviKbgnpSafJREdv2hfcvq9FGhR0BRY0NWEWpM634zYWiROA7E6ICOj2e81+x3YXbPCKBb5EdEL
vCU5mwHT2xNg6jlicM0oib7u0T7irfCofKMzfVpYCeTdVF6vM5n/PumeQt/tC37jC87l/2i72ttW
bDdSCWsc2ZyVMMTxHQsTGTV4u9tVkw4Sz+sa3q9KCZhgOU9coF1zu7NroPErTMBvD508Ls5d3QF+
uXr4hl79OS8IEE5axC53xKaHM/kj3AHSgFieFwDZsIFvMUl3uneLuhpMPHqBfdPtJ3fnPw1RW43k
siCm9N9JEBKEfLu1J0wIl8KBG7cikV1WgHWIvkqbncyg8ueAYKcq+NqHnP6v2uZfvJJq0CBVbP3K
TSu+0y3YhCJ5bmpf7sYviV887p9aNbCeGtp234SzEwKM9QZ9YuVj8bsjeyqGXmFjgK8V+CJRaXD2
JIEFpQu2QGzZfKvvjYKSWEPUgbWulpZIbO9cl9fA3XEhMhgk2QxIPmlW1gPa4c2rsy2gAy0GXLi3
fC26KuctAg3UoEx/VUTdc0YMzDbmQo5LlxjIlcNyT6KHOY4Xl2WsMlfW7GGuC0DL0qB4F8bacP/g
rzAib64tXilTXPO1lezMREpq4DxO9+1SYIB/koozUzQzRV2b9sWAld5YFtOYT47evGq75uGAHPKv
fYaQY47fQLY5ps06F2WlH6YUDojUe0ggRxplcFb4au4EG543Hf69rw5ntRi9d/Tz0IYHKZLhoX3D
wmqc/fOmBKJNT/hmW0RkI5S5gGdhV0JpdQJOsHLI3tCNjXLfJPOr4m0bRFHnvh+ex5KxiBwa0xMm
uGY3d+GdiY6VyIhH+DJllk7YG19O0b5mTnP6Hd8DSjxC7YDJBFKbt2KFrrfNXBWkmKDS7DgpjgD7
FIVUHuAxeEMLN4XXq85IMcn56J1RmBXOJ5zch6TT4HrFeTnom7OTdURPou05HjE4CMh2yvekLA5a
X9SCcAk2bbA8+FP+A73EzfDqJlQXSyRBWi+0s1I+VSmO17o4pv2gmTIw0aWN8odZsIOInhEdsSEq
V+i+yhIvNxELHSdjSwb1MTwIOOti4aUafgBcDevCEeN+y9txi4iaK/IJzhMGzT/cjvPu1nV1EipC
aIYkxEM8rpiYjFI29S0uKroABXXM0r3k1VdczTrbyPSNcGHGccrV38H5DguSXffs1ncp0xijzTlD
5pmrXbn/8uopozeTSKp1x7riVWaYZmFgW0QOdMPo8QR6HRccsg3cE9AQsAWBS0C/G2rS78Wnmgvk
b/dMogyKELQI1apRpN3s4oi/10A7f0WEfzisotzKMjzWzuRGvljabnvhCRZ6jaaV1/8dfHm2j+aA
GN8Pf6JhO0CN0WSF1lfZJxvfeY4YViIYsYwb6hJsuS64sG1j0x8+XLDW6VjczlrnchYtUu2J4ohu
spipniCS/1Hn5iBVG2x7iPTT36bBc8AbkIMSYlSM/KWmCdVI0t3k5WThxbjBW9asxz9qPwyynucT
60xLMWdSH+i67xWU46KnmaLLXg7jwe4iRMZma2U6BKo1k33lLa3J0z1jZ+HXrcIrDQfIfTRW7crN
LkkMzGrvaay1ce2OxX6Oo+H+2JOwc2qHKMWkoqB7Gppc0jgK/8D3yrx4H6jdrWN6CoRuKK0NaeUV
q5sPeoTNk7PReyr3dLV1yMrAQZ3mFNZwxc+C0caAV48h2LWm+d3DpmIYalKomYdbPQyuyQQPC863
JhyNDltKDVAG6YFDxXHMlmUuHg4Bm0apNUGdxAYu/PjEYPQTarX3fCFK6c2xRpRyr8EEGH1Zg74D
GlHHTAeepe76VtR+i7W/jwgMh67R9Pm9OzmZfc+lullJiw9Rq2Q5j4fdmYCuvJkPVAblzcsBmTpx
r/ECehvfRAx8BIVPqIex5ev+92yFEYzn0dRBz+tukpBCxq4JxBnEjWQ93sXRwjPOW5e+lfBo929W
QhYnwuU5xaVDyhEGs4/L81W7O8r0qmQHnUk3txawITJgsPapuhLLG7k2tLk14GHOoeTUO2Xays5O
gURNy+NKpViPGiCGXfJFctQFpQK8GXous4+oL+fTStTL2OVBTaK0jy0UKiRXv/QfF977Xmy62wXI
RyxQsW9sRGIg1zWdNbD+tXYLS//XfKBCmTgjAEXC+RD7rS6EAgxotJv+eeYrudctZrEM8JS2lCGc
AA53xRS90G+os9yydxw5qGD0qg5STx888uJ4rcCaxbAeVmCb8Mq3siPwbaBzpGWrn7vqBiYG1/Cp
1yuDOA5nbiOZtqC67ILHa3imzpMIn1tuBltj2kjbPimxzZNs7cGAti3nWkxsK0gY5A5l+EI/a6sy
5Fd+7OSfz4OP3+T50+rtvk0jBHLROUKMh+EHSBpghv32sXOl7KI7IvX16ARIAAYbp10vyUKmUWa9
UcllWeRPybNhS6iZbpAe/ZGz71P+QNwB8Xc2hNbyz4VlBgCbEVMr4kjApRAxgZS59h5FIV3P0SnK
wmTU1S7w16jTyXc+EnlYP5ryzZfa7jx3UQKqtQQTKJ98zz08TqTTePeGIvKLrZ52DOoIGi4aUdwx
E+tuEDgR9t57BMec0RIntYVShvyb7qC9iH1q7g6GkQsiVtr63d5cb0VLawHSTzCRP0CCdqHzfvww
lb5+bneyJpuLvCGaEC/QPQj87n4gfBPjMs18L7R5NpRqTodID46wJni85a8EL9WOMriLVVyk3B+r
tzUB5f+kuIju5TlMTp5k1mSbZs1emzhUK21zVL2Ghb9AEWjtTNXaJkCXJZtowuxHzHsz1r4/4bNe
SOL3f6Hdv7DTqud0etoxr+sKS0ZQhQ2lqlphIyT1sppzwnzX7MpBZVuzcul7h2UB0+vrKlgL1n8w
LX4Mv+yhpq8Ied1eaeGCcApo0fJdim9Y68C6sXyOUXEaBPx6tynyqRHHwEqGvwne5zTu1DRbkq0P
pEdC3ZQKH+wnX8Qs+hl3PLeU4H7Ebco1s77ua56hNXN+csWebHZNdz/ZSjTy0E1FplNiT2+xeuwl
9yXWv9BjrcuZkEMoD+gb7t4weGMYQhFwHlhg2/HrQE85qkbZzTrT2bKH5acXagXp+51U6kbouOAq
6jeOGNURF1yDi15Uunm3wntW3cZxFgOi9PH8xLQ01u5eVQYtjc/KlLOdCQcvuO9t9FtADF2HpDcr
qR7ovKelB0RXabU7uW8wlCPPHeaEdbh/dmcgh2vIfnIlsLCn2u5bLFFqsTEi3KX8ryMBn32v8cPr
fX9nRkFtAwm5tlkvaEZdYh/O5g5YTMxe/xgbtjzKz7MP1HVnhDgsy2nWWrmtCDh364lvLG4dortb
bgvwcVI5yIhLBUN7q0R7DyDyf+l7ngV7e6ShO3mX8lIPOjmRSy4GKjbfPpaBfeneUbKtkDIB5JnW
ByaFbS9qYXqVtpZaVUVgKczOZeeMSwpUsbtdf5rk4Szy2Leejc/SpSnuGjyc1r0bY8wyjK7N5xiu
vHrRhENFjOMDuWGxiXHujL4dHLeeej7wUo48dz//aCloXYmT+DGvMYUEXEnbpjm+blR36Xe05gu4
OBRufFW1kjCwMxOQvcEAvCi2sT8FAUl/FLtxSOsp8gHwkCKQUeB5WfgUypu6J8OZZ2O3hvW2wA/g
Sp72GsoXrnolgSVJ+4DiqQgw2I3IgrXdVfuOuczFtyXYngV36NK6RitHerbauZzgASY3RRjXoRQl
Jo/Q4b0Azky7xMNyI9Rf/YlxJwjL0jjlTpRTs0JP110Wt/GiGRoSwgMVN2BZgt9B6vMWYRrahtEn
8zhzpwTmBkW6HzYvDSkjuXd58u/VHTpz8o83Rq0OTtjbcntKQsYH4QBzl5MorDRxc782tZHzthUE
OqSt5pE/ZTwKLbrUqmmC1r+L0WIasnfPFXjgZ6b+OX06gJAMX/6uOxzGEPZTjplVe14oPgrIW8ue
F+VUJ2MrwXyJquSzMqhQtepqqsC7SPnAYPZ3MOuEGf/9Xdwciz7hvqd1l666vV67I0pxBTICYrgv
StybOUogOOUB16XmeixoRgQ5nSrPHpa7d3xAU3Rwwed6txFJIkfdlYd3KFBxzG48ZRzD5VLJWhFD
buLJZh8UjsY2M2Xoj06wzyY/RuMbuqearwhXSYvCjpv+VMjkAHNnNxO0np5qiMm1bCXokoev4sJH
SYUIMvTU/76rnGs6B2PJsshaWKccsjNuT08CbmVA6p3eGCycn3MSapUULtagLof/IbNsJQVvc9Gc
CrzvFXuS14HtjPwyv4iTnlQpFxwxlqe4TIyWWMuVBMA47AQdmkUEvVVN8LpAOimRlqu8PFfvjF+l
pxQlPV4zovZt1355hZ1whUyKxguEfpHMUMuWsYb69x2dlfw4ia9ASH4ALcw27nQq9PMycaKhWW8N
F4Tj3eFus0HZ55xJMZZfH/sRlM15djokw68X5sSHO3h9U6ocfCICfHYxyk1v4flxcG1X4IhdNB8P
JCBiRl4h1VxT1M91iFRhC0a6Ophu2y/6LLSUL/vZxCRcCEchPSUn/SvxZDCFlvMy0RkLPALpBmeg
iRpv1SqDu+Eh9eDdWXcEUOiHiNcJr/YGteKzUcI+0+1vqK8qoKI2vbvhymzCV1SJiFqfhZKGZ+cb
6gfoOVEVqKxqgi0QeyIUckaZMKnX1oBL5LoMJ6XPVRIoPMpZQ72RnUxAMN/HtEtQSq3glwVo4fyc
MK75wyFuUFBEw9J6ylfuQe6WJSZE+6P4mlpkXI2YpiG7TYblQ3bMl13Qneg4hNthV1TP35MsETaZ
TUrsJM8jufMrzlUrvstugztxRQBYTIo=
`protect end_protected

