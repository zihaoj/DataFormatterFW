

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
adET+ekeJxXhc2rpmfsg4JpDe4j4r/h3qaXK6bbjnnJCR3NbN8WIg6DBXLdjLNCpJrXNn78rYe+e
iChiFer+Lw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EpPptnOuZr7qIWcAEuYBvzKzA7u5xTXGn47Gj95aP8z6BvdKdbYnb0fCC+OEbDdgzfB9ZvqVnGF9
NMOM3fwphT2Jql+yRVsPQ4Zx0mTl+kyA54gISGPygeH+aCjxF4alLsuk/vXq2e5xzafcGsYMn2+A
o6LJPevzzSgK8D6moJs=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oB9M8cJCuGIeW7xleRmg7VDEqeLaRXwHlLK+VjCPJDDQAxTgk7137Hm+8lEMHbl9cIi8e5wc3wCf
qYgaUTWAEjqi7LxqAWUAnwtPsdKk6AZXxJa7sER6jExfouI/CfiMASx17XtQYSdD3HmGA1EWJuoT
SSiSEn+FnJmxgoKCEbGavuIlxp7lBn2m4Pw3Zwj9DUgnjZ7O7c2BocGHlWFXl4XxBSR6yzh0GKKB
e7zDkq5DnRa/tdChxDpIZfIi66zAHCuqSjTZy+ohEE8zu9oE2LjapQxY/Y1L0hAaZsZMaIaYrrAY
kCnl3I1N/9xxIfcBj2FuPKX0Iehqi5pmaZvzfg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KQeYm2dM7TbDPDfDu/5jHPAYWHKekaI6XImwxJa92M4BxUCESsR1003VS+8j+gFawZEIl+w5yFs+
bLwXoZ+d1MrdSnJuR5CN5yyFuPP9o83pgCyu29mBrvxvtU9M+1BTzsfbmTxR8+uNneE2hDIObcGe
BQKZoLqui5wEXeT9uO0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iDjxlA/jX5Zgo2m9+lGcV/fDMmaSNvYoIcpF2bRzDAGcmANVdBRMlU4uzmG55ynUETIX/UKWhk2J
+j/xAO0bBSvQzp51csEIaTZ+bYKNZlRhEL+QkcU9RVOThMJK/ZAN03/r08V8X4asbe5wdeNfrxQg
6RC4ZH5U47nYrztjLmYVWYvroct0WcyW1sAqyWVych+3VPPhQngVLB52egaNrRO5m+7hNvPUlpp0
R1tMtB7gxgGksEyn3Ord3AgQlskmciNW6wqxRThWfTUeKAA9KCwZPo5qP9rFKfVJjL6zBWpDawnK
JQAeRCkSl+1nAvdh4rKqn3sXc0AL7dHuzHQYzQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 43328)
`protect data_block
LBvt0vd7va00aYSeJiW5JQdRLEv12UfsA1x8fbLn/B6vcJD/AvCGQUTEjHuHf5aJxjCQuLfiR7Ks
lqmS9/uPSzOEpa3M7uoB7HdTL/nDp2zJIFaNDCnT0eT/swvrm8VJvtVYk6LDjQ0FRJzajV2/dwXh
x3PbHm0UU3D8bQ1j7VmM8t9ujV/pRhobhZvtJLsihoJCe+Vigw2Yni0zkYDLQoGx0PSFWYgIWUV9
ZTnorR0bmWiN6Y/mdcAWz+kiYxDiWrC9HpdLK0rtxDrLal+Vg1c6E5WhPD7xdM4I2dsCLAndG1X/
jgmVGbAy1qbfO8IZlfQbkugdgMkz0Pz3sydHnsg38+zzk1lddMV7//BIkM8im+tCX9+HqJYWu/un
5nm3rfWUubr1ddhHYPkolOjofoozmhjthlwm0ctQ3up5MHOGV3xfMwB1GauitafzEdE9+rhKUChs
QVs1AYw4DPHloGs6AxP9XBut4GYaWFcKh/3ekwrOuI5XvC1ZPvUL5Q60V7y5qcAKQ2C6UNkUyZ2J
ex9NcvXGmAGuItZ6CXjQC7P7MZxVBcbsef/w/N4qCScAuUAvWbgPTDGeDg30VTKCDo6v78UQH8GK
Iv8jK37UuiykQbsBRHmhwUysNSTvX1POlfLFeraChG/hNu3pbWfHCAGvWkYyIM2czZYj5aZXLV7E
jlR2wCjFTzaqc+T+px5ndmWBulm0UZZzEpLhKn27AcqRbUlexxdTMvP0aJwzWcwihl8rWAjoQybL
7hygW2N9ZVlzZL99gD2mthGTldA83/6axuPjOftmzpIYsDyeRzXEwQig2QRtKJKRUdtX92++1jxJ
2gWqFGn5w5rIPHdkCBrp5yEL7uVECFen4RTupNjXDZ7r0Av0DaadphDk1soSngJnct2XIm6rgc4q
Ew0lHozjwjcA6QxnywdakTy+7wad6UQ3a4mT5mioSDy2qr3ojJERWnjTVfm8GLbgnt/avBH+Ywxp
XShkAV+c6iHCK/ve6Bhg1+b3WYkEu8ry5L6QOY/l8doNd/Q3og8Zozt9sqmSz2UAilBOCajbpxW9
PL231qdmivE/GUkYNN8YthVlPcuUwo5KMXMuWF5EyMboNyu+8aIPwyN+1pS1aVL+br+R5QiFCEXP
kalA/OIaG1QWZ4ONSB922OA9DM1kz+rz28SO2NE38D8WdmG1x9xxopbOeQTZEcqUrVM7X5F/twj1
S5EWbzagfJRDj4uYcPmop17wx2jLRUH550CPxsgjCGZWA7xl1haBNSfn/AMDgubjnl5iMjxNups9
phUHKgNlS2SafdbrDmfl+2HatLT+hmKk2PEVg5awNDYCoAarU9RP1lqZcxouxib3levRPaHpeY/2
xLglJbTby6cJRMHJ0gnloG/l2VRiOqlXguHobx+y+RE95wZkerP7IZJPnYjo64ctEOM/UF6842WH
2wHWjxGl8K8ELG99pVFeGY78oMayJwZL61EmdYW0yai9DV/wz46r2HBU3mRU2UIDw/dBD6bFXrID
yCYxpITcNwal42V9MqM+zu90cMVRrN6AlYNaEU7FPbI+ysY3t/zDSh4EKly6e6EevNN0hMbEHpe7
zgbFfX8XolKiLrk8hGZFM9TUpY6V/D9YCLvwfvQ+HMoue/ntGHAV8VCfqVN9iIo8bQ8/dqiYqDx1
G6qW37AgqqRBJOBiF8zoEY2+TbLYPxUttu0nugZiJJC1FpacsQCKomnRu3IBl9KLmYmkPdGtH/Oq
DRkg5x6Ua99yUOplu29xuBT3Y95ycIhUS6ngSBWx8v6YJN/vQhbBTFwNSivzoXMvjUo8oGeMcFxJ
F9vMO3I5tM42vcOB/zn9Xlq4JWxnDiO9Fi1iDSoLUIdbXaQ0D5hIhiwBE3jESzSYJn7zI36tbtnt
CfNQTxiSooSyCaNmln8s+Ag18NAJY2hUualTgkHYk5jW1FwMXj07FvvYORAWxLGPhhtfS1Yd/xTB
4ANqW3hemIt9b4JPC5u2SoJ3yudAZWuaJegId90Os0nJQw42pWITVTmxruDovhEtxl1GeYJyOstU
OwjhNPNRcQdBrVU2nxAIWQKPu7jVIjp5Oj3APvSiQyM9DCIZveL1IjNL7yWoYUpUYNpdCP2OVGbQ
6+f/C48I4HA3+Wc5BGvynEC7PysEYzb3ipCehzoJc3EUcIAiFEht47ZCvmgYnjx34B1G/UqyztEQ
jwqHX/aCtfN1AvTcSh+WPpPDEDQbVQVHktrwMrsezCZLeqCm5v19oVULe3UUjFiicqv3QYa3klmo
63rM4XCCcWt4Lk1PYOXKfK2rPl0RVxsbfBqLHn7JlwMxXkRopJ/uDum8S5j88Cftf+ZP5irXfVok
6n9blAxmc3DHHe7VqRCvaDDuWi66uVwdJeUWnY4jyf+wkDeuC0Tu0iM9gZLkkd8+eb8VKDcu+vKo
YSRrhBWTS+9eoHXvJVRwAg38W1ujStUH5ClUKfTqhEZeYinPO7xoncDPDZthOm216xp2I+J5eztw
ie0GWH71sXrYSU/iDqCPOEVphqnkFFOlSH76+loWkYwG3tj5yxM3ODhmgFD1RdJYIkfByucfACef
91Mh0dn1stzzon4GIhIeJhz4x/ClvSxDOEoWVHtJoVHf9v+zYzaPjysDjZsFO6QXW2Lf2cW+F+KN
NxKVLXsQn4KCMNUQGBEOjQQZRuB3t2D7jVX2tH1BKRHrpRdm6f5eHfPCsj1LooHXjzB8WJSOnEkI
DaO9Ww8JHsjri/6o7VaBGnf4Wtb1Zyhjj2l75TJOoTXoPJ2lBaR2GdimRTBpTzYBLBFUto6HSKua
znyUuV5ulBBfNDilyq4Za26xjp6w+qp2ovlIFNBXUuKmPkmK5q76H6vQHizBJCpEAr7/Gx5Ss5yP
hZnQsMEZmDVpe9+EK5JNrTDYaObayqYpANfPauKXJTLx7W37guirAj40hAfdISDN80Enq6UGot/k
JMoHzohD3wbqJr27KGZzH7ayMWt5MM4qanYLtDXR55Il920Yd1Rybt/XoP8JB83eLpxIAPS0RsLF
QvNvQG+XbBASY+nJiuOIPqCFNpx3P2u5MMX5gSLdmPBlYHk9YBhGqd0fL8b93YGRlXAto/qTAsRK
W2Om8hPQSIFVQDgpbGsNLQGAXRVkdNUDihQ8NFO14bqgf9VEgTZ4cmCUe191GmzDEwzohYNBS1Wm
Xafp2jTTzNn/bWi0iS1xEndQfo127sO1xQKI35cLVhb0iOmRKFC43KsOPpFLJjl/FlU6AFueAGMF
aqDmRwCNTLg7aZa2ErikkXdoOzwQ3DQ/A0/uWjK7LN7VdwEukVGgVVCxDk/uHHdg3tdU1eWJqlBH
5J9WuXgs8mNrWZAagBCcPP6MD4hU/3Ol4QHvnqSLV49WZnFmJmCoLKXSyvSzqWIDfhRWUcAw1fCO
gK8uBt9BHfSfeRmMFWErVCVLdnLESrRia3E6VTh5ljKvX2tOm+wEwuVcOp+8IY159UZ4ASN1P7tp
p3D/exEuiAuXD3Zbrax2VJ+Pic9EghhNR3Nq/geIizzaeH0xxLvo9+qoQajFRgpAXFHjgHCSX3zC
tTQ66XVobgGDAqhqIcL5tEiJJsqEoUpeSLEO751ibUOTfZaTNeyVE8tARy5LuBobm1PRyVn58ocZ
GB9t/ko1BK0HtEh86fWtrKpRGb/PpbCZd3Gm17KCIcCJUskYDVrVzzwm93PASt1tFKUmmnR5QPX6
eNTM606BesIpaxD+jgEAvvT1y1Ufik17q76O58fM0R0iOjAI+4d3kjd/8g5tD6LCxyXJFqFSvL8B
M1/AOk0ix2buam49rkSkqobb3D3mWPPyvvtC7RkHxrx83i4jjzDnOQBc4DJpB832/HjNzg2sHDpo
h3LptnNsrO3Ul8c3fJOF9wXISU85F2M3StpxMaCTk/bxudGTXuX9ga7y++AKNxyAttm/K8i7cUzR
vBpPoZ15998/o2a8ln+o3uq633rXw5qmwnjaZUjRriAexcI1BemUKaMQlVuBpkSHMYM4wY/vS+aR
eCFC11GbpJuBioCrXjHKjlB6GC8GDbD8F08qOmRLgw/lrLZaJ5OZxm8y8mVERENo8hguWioqfvQN
YGv3Be/6S3VIqIQyKTfKzPpLWOzpaaxXDkm1HvE2EtdgiIAqUHVNmtOA44IN28bKa7hDcpDfJKGD
ZTc2HDbt6oORySfYCjnuoxo8LNAM2E7cSzyhe12kL4ZggvLrURujpFTxmLn+oknNQaP3iSwr2BhT
gqUDwu5JJk/wusI2uDChGYW+cUyz1QLZlR0zpWW5dXGRDM844eQ/20iY5xgh5dxbXHD3ZoYfO972
kJIHwOR5T32Zl3YGrccIOIQx+uAmolvN4az4WCZ35rvjd6ln6hHpQvG5e+Nyk9nBRDvoOZWAsDv5
ZxcHZ48WNlvfo+SQCsgIJgKuNKf6WEhbnI5y4juScm3ksjb6wAsgbk/Pbq8EYN48j0vyOA2RWTCr
MwB/IYHahHWFkXaowu/E46qE0OFWdc7V4EC+sDAoNbFpoDc7+GnDdq/Q8uMstuRCrLS4ncfmrjJb
nsnVqrvdOb0taNiXrWAI3T4sZmJyUlozEMjPpyv26UuxVFHgMHgzTLvT04MoTp8TCkfy/BPbzs5d
mMguJgaD82kDEcVzHlaKZAZ2dKuz4FqQGuj2H3DdbNbMUQqvRT1A7125r3aBHZB36+pAs/eCE9N0
TLO1DBpGEEagAGP83naFWxq22SXpa5FX354uYpkB7Zvxzo12fugY0NSOsAMX7i4Pes4T9iDsNcOJ
PVtQFNJlqd4pi6sPa149eBg4D68PWns9MSSy6ws1dSJv32X1JakjKcy4KFKa4CkZt4YXRCNt9wFi
vuJf9wHJ3fVjWS/yPvwh0cNOtvJj9VRqWVTHw0co71iLNF3oOrjGMlWufAXPunhr1Yxzk/VHvLAn
8npY0l2N5M+8c/GtjplXA68Dh3lcaa5W+6rKc0myhEUECfuYD3S75NGz6smzgUsPuUGiV0MJIwyc
oNGxVPg7YQMyAq2NsSlgwgnywdqTXfL845ufkg3XtlUQxiXeKuRKNFtduFb+4nNYYdfI69kBetxv
6j0OK5aZEpxpOHSAniqycXQTBv934YiaOKOdmlRkItdc3n08q4tKQH6hEdqV8YHZqu1kfxzDb1qW
hrFtUOUp4IjKM0wAzJwOIsBWoweXFRyVX8XpqANEXoOTBn4r8+Oh64ebtvYEJYjoXaH0Zv88NDrP
pjPktfSk6JL4anacesSwDdnmiG5lAPUdOWmdmeiIBs0ryJPDP6cKj9RXC1a8giSLWfQHpajJsj/m
Hj9WozlIn9kHe+d5kfkF57d6D4fo+wLORyhR6HIBf7Rm2VzJSzJytgsIMcauWZVcjlDiXHu9MV6V
Te8nGKowdSNLdxkqNTcBPFqFMdw8EBTV+BKFeanJiAYIv0yqZTCP5HZZuh/89e5SvhvZ/LkOe4n5
I5UilEfeuWltDLUblngjlhxtWdJJeWdfQKdY4ASXPbV8ko2tBS7qjEAlZ+/HKE5NwWWknOIbw5HB
RbACMEAgZpmJd16sPAi16n2Qy4Fm9G0ixFpGtqp3EunT9019ozeo1qVKv2dku5WNDRlR7Oi0s2GH
BpBxDI7jQyg6fF4U9BTitQmcpkL2i/6vjBA8ZLlmsU7IBUTSKjPgkfk0cL8a3ycNlysL+Bz82KSK
fvTF22YAZMMLxhpPFYQScokZKPGSoI2MiAB17I0aELXkN3ntjPgsvkA4tJ+BW917Qw2mGCsIvy8U
1Dhd1BTd4plk7ZFgvcpjWbPNpjvQkEaFB/w/TEUkqOu2huHv3TWw6jhGRbZHFFvHxFTvg15VrDSw
hFLIj8kbaC9SPKeHOm7R9XNWhjncyZKAs6LRElRAwuQkuNcBAHMzzw1euhmLJVsEpOWXjIMOe3tx
3fNOSVxaQVr0qXsT+uf8DfHWz/rb2S/+kk/h9OgcUi4T4IiaRWg0157cyqWZGQTRMyPti52KjiM3
5aiUSrZVG5dZMmARv9SNoHubbWh3bz+hncu+oQvwpZ+YFLqybeLQVmtTV6D/tFKqJHapKoRD6DNp
20QJm+uQtwA5KPkqIDumyfs6UNz2WVydV/OsfwEPlLVgfES3ZraK7q0a914y2LDxbi/1kaJ9+wOx
EE3Tkl9ETcR2bj3QdxgfWQiqZMQ3VQ9FzFus4/hKwvBP6YDnT8B6iM3APNINb+3qbpyaTTT1BUrU
g8Nmcz9OgfJUyqmTb1JCOyKZ0tQQZdGsIV2XBg3uUIv4+Hq75HqktdM3T2uLRYZpZ9IRww++CyNv
O/VtWOqDtpznWdWlf587uL/0U7l4R7n993tQ9mWTp2CNQwoccCuVSLV4f44j7GMFOaAdyz/V+iWv
QanUkCSBrJsodevAvfQlMztegczENbUGfxIMyuf41hnKnpaXzrVQgKDvbixGXAEtBEERWLrmZFs5
hKe+IPXIL3UaMdpNCcYZS8GOT5j31tU3M5WGVJai05onAwJn5r9bHTJyecrozcsPDop+gNdPUtuS
Eqfu6p/dO8nZ0vWMiTzWASL1vN90dPKi6jGNG6JZrDPuyqBu+VdkRUq4fVAZactFmz4Hm9vxkqoh
AqEwk6i43/pkulOKy4DnsDM5IsVU98RdAst5vyChp3qM/soaXpkzFXUidQLRgC4jLKfb1hDxtzg7
lRlaTouVw4Aw3MY6W/Cqpm26NkKu92+PJi6jicAWZQPbPu1wKPVpbdkd//8OVyRr53TNnf1mSpWJ
5HdnmKAVfYCXFtGlvW7DmsL/Xfspo+5jimvVYT1vINEpvRU91YwR7fuNFBUJFIHijollfIP0FQFn
42bHKmBXuI5L21qJXAbd61juNXuWioPUduINTWbGYIDtn2gnXezbag9P47oKOIU3SgMZJbyBPGH4
PFDy34oQ+tyAkHW1F1YYPgw6kjAsefJSzGNV+5yZ0yPqM0aPx4pjIOQFI4sBqo+hpfPtGqao4W5A
4g3YTo8pSXm6YDO+cia265hccofkiRyEz6gJiiUhya6D7MznelmBNhCkdxpxqU2+NNorv2BzxY4D
lpuElO6sBrxWT5+zdTy8IT2h8FIrSfu4Zu9aiL4bPiHxHu9z4kGz2ZsOFXdfg+oHTZxXCqP71Sqj
CNjPYw0agaND6vSbXmHtS1fKlbpWeUyBF7panC1X5BiKy89W74iCPIexlK5GqWENgzE7aBVIu+2J
cxNHE8y4DP9y3dNLcZ8eMgreyPP+miTPDqAJtbVj2QTdGTBhiz0XrGOZgSC8IHt16Sr2+gnX4EsI
S7ew4Vn8L5A/sapJjnNY2Er9vbVCoqgY7NURuHKjRtaTIfStIPZrwUJTN57v7sn2i0Yp3cmxRJNX
9HrKV+HBodHmPsLwjKRISN+dXVx5PXiCOTsLAgsiwqbFTHfbaQaDbDz6lZs+vKAfKLXX9JvnsN+G
EBJiZpZSkH5JiApTCRQMv4uq4dfnmhLiW1im0DHdDlQ1rhIjeDzZlVaUik2AIUV8caEa6DOYTTYw
vXhe03PDEJ+/+EvZe/AOmM57JpgBlMQtoBfpmRfF3LIvj4mer1bwp7FEEsrnJaFWzzxrLnGz9ORk
JUprZ/0+hvwlYKEVQ21YCoWsnEw16VGne1pAO/D4A0EHBEJ9SzbYSE4xt4rveQJh9EunSRdUOdeB
hMyHEq1nsQKpIgdBpfxmpk2880bP5Q0F/TfzmBz75K2meOgIODUUrkf9kKyAGpp7bBD4LHQhxlEl
uPRBiYwJQl9lgHp/t1s4Gdjeb/bcmd5QyBUmTozRRAF1l2e9Ni6xaOX3oErLS8czUtXaI4c0QtYl
vPP/Zo7LS6zVI/Wvxn44EO3h2hTL+gfKirHx6mAqQAMQ4uZy+kMdATpt3LlsxV2gA/uSuay+f5If
bLM0W8/dO7R7ATZscFwUIyohT6CSqrs4O+UM6uWK3135l3Bpz76j+E+u/Mvgr7U2qxTmDgm37Tv7
j3RUy8TUhYAIQJDyqoM6X5rxqE+VkMtjOByser2iuq68d5pl2aSdQlwc84DUflnqdazWvOlasp5/
CvOu6y3V/IvMe1GPyvCrjHTQdAg3KXD15xvi0ax0f0E8U+SGa+4eGz49/c/sEpFOzwBO3zp8pEDF
hrKZvrZ2CnTkxVKRHs9gWiWubir8xuH6zqrMvfoY6BzN4EsAEsBqUuz68VjibtbKSPkT1SinkfiI
Jfp50uxzewJyxHpCBRLnXkzUjylKcVOhI6uv44UVIyhAkEScejUPcKkHJFVXphv3/F3kHO3aW9WG
68V14PCDryyXtEnFhUnAzO+O9Vg3ikoTGwFAqc3nrLV4IWWOV/3wCpcZp/T/N0HF+bqY4h/zbD30
k4w2jm6ZVfjIP6y5wLBqrZymOopuDwuoclt9XyPYBsEvCOtc04cc8T8Uo8upp5xADSchXek/fZo+
nbaOsm81Ga9lKLmOcI7BHcsrUthnALt6cEswaphqb7S7xmWTA064pMA8D7qKrisucSbQV5fIQhK3
sGtgJeA46SBjnVxxBCuvtR2gA9O47eIBNA1YDZfjSMcomUAvVjXGV6fpjdbILt0ISiuBg6bZQJ8R
rFJi9GkvRP9E2ZxGgpOPoPTkNURpz3qTs2M5+gzyPQjeDkXcUKQCVINqYXIqqqLRtfwjvfglX7MN
fQv+7srpL9ZFdMQKxi21j/PPFYyZTr1iqhxahLpUvP8tHp2qQMSJmWX85D5KqynwP+5vD71e1tRP
3ePTK6mtFaV4V9uEmc4xU0jIxkcAw707n+YEokn86eW1lh1B4DPt1FzmgzdANTifFQeIOLVgMIe5
qHXPThTKuxXpf0u9HWFRHoRTVkTf2OAmChquV8W9WdTrUeTnIjsyH4TBQeKv3uDafTtgbFA/5eHM
cQhIY4dYVdOYRELnHirjqZlRto2xcFOmC85HtST3w+87w/a95GIBtm4U4jouxsCXzz9BFZX6fK7K
i/uyTY5AWHPgrfXmyB1LwKRyuIHFGL/rV8DJwg2T1HoPy7r5QQgT0HCKirmorYenOPdU18CsH08T
5uKonWgM+saT14v/5UDgvoq6eZvORwvYwZTZTNs34kVp5pNEpOdm3dxg8ddyXUYyPAb7/glNIiYP
4oYfmN86Cirrt2eQOSlktf6NLj81AeAgz8m2cRdQ8yJUDs1GCcQ6/Esa0fgqLKJlskR5022BlFH4
X9qjn78RaBUcsfhtI0+Rsm1+RXu09nsmZYEVFEfQFNKEcvpYiDqBncmBPYFbBDOhM4MCE/YguGfu
y5h226kGBLPqQHe10mI7VtaMaAXVzOgiRs6Tyvr42JaEfM/MCFk9JTQPeMuxIq/JwoLUtSEn46+O
HJE3fDkb+uLJE+/udBhRN9V+rqq4vGzs6exRcynUJDjHkS8lBINmtlF2hABF+CsXMJpkQy6dwi+U
di0oCMwOadH4NsEZiaO9oisfbMrqq9XyyhE6fBkZlmE+oNVUzNLWPeZ/t6wvnldz9WrvidhIy0Ve
hVdUfT+BegtUn/dlHEyg23TP33vkhmAHfMyX9zSdAnW9d2vVFI7rk0jbtQ28mQFTNfpRh6QtCwIC
RdOuAGPjP+NjR1I0AN1QDxbbbUNB8zavy65A/elz8o4yoC7xK32d5t/rtiUBelwvLxtY2TmyzoRH
iWVmR0XJs/4VzUDMoHNUo7DiPd/gbXAV3UjecYWyEDfIYLn4D/K07ujzC3iO+ccWhWjgwkCErQP4
c7Cp9KBPpx4UKwUFD2S/RW6GGoG/fnJLiBILW4RkRgAwrzP5bHStRc0bmfxQy+Mt6JrwtenbH1+y
AOPqvwbzCD6hVytTNjBkNiCxFXk8iz832l0TRJEK+gQaIFre64twtx0iOUGXa3IYsZ5uoOjepMS1
ZRSKldEZkPG16B0f68YO9Gdtu3c43zXDNBnz8Me2CKTjg/uro1OkWkmm4bL8KOrux9NOC2Dc2+Yg
XoraPHRSEK4TqdvmTCqm+CmfqPJEZ+YS6JTLQ+K6qmbXkK8yJO7EZVglviqjDh8SomBosJrdaD6/
9FZ7k7TD0e5SdK3owide87x2L/Mj5LAM/cZJf1pa7m094mhvSUm7m0CqZ1qAa85okRRxpRyk4HIP
uxPhcAXwWJqqzhj7n+kOXRJhkoo+lFRoP4OI6dCpD16/GIoqLQm3ZZebmRZpMQtlKtNTgisIotvX
oRgb12IVysR1/GxOsI/8SlWDZAUUjrv+zNqdaCDd04V6GO2S72Bg1Xu1PdHZS+WAmZC0BqEmu/F9
dAWI7tQl6Jx2OwX/dZtgsH04Kot+e/J3V8AQWDxv0bjkv7Wmq+5I1REO6vgea4K/sMbATr30lD5T
SGY2/eyQ27PxHLMrNpFaOYyyQong36A47N6it5J/mEMwON2JGd4NqDj5jsjPs2/fcnqCgyeEryJt
IOuwoKWzInNateo66weost2hWCLideNp56WBXze9pWLN/3T0glYJT2ZaAs0vRxJdhc02rUJZrq7/
DVmg8tZZrS+kG1pM9PXzg0S4AwTztgBiTSLM/dj2ZaTVSkAIO8/BAEAMa3GNP7o6LysmFXCeyXUQ
zK4hG+0CtHkEkJvGiVlxBgzhrLj0+Sud2RKP7lOnBkFBvwpw/YUCJ1k3jTuCZzK8QgR7UphW30Hg
aOkgeiVL0tM7KzwCPIPijVwwrQuwbf7WZeR6wsxvhEEtSG1nrlO38xYf4msLruN0asmpvikO72CP
t42n7L9OwCMbeBxL8daVXstSX1cpGnJ6SBoYruvq+9TJxz0UJPj2jwBOlp8kobpYnIzB1SSA6rHv
YcpQnwb1vGC6LfHU7NMxn2YIiMnnpEaGwlN0FiM/K7TiGpLCt9ie4TPHAqkCPwu9XRIYtXL5zCor
xykoSerkmEesOLRakwdraX7hy3p2ke4Xw7zSrFsd2BckMZ9OZpKBaJ3qIU1H06Fm+14TlOZ+ZpLP
ikegW78bF53gbH+SmzhaZGmZ5R/Mu1d/kqpjBfRlU8qAyR6L0aAc9y3A/7+brUXIRoPcCHAKKRb7
bLd8248Vl9vgdfzRrfz2nj40pBp1Faj2ZjsdHySrQVUcIUNgPps27Khg+qEmZPmhJxL7oXYc4meJ
5kcOud1chopr1j5f3+GJbk7VmTLkwSTQHPnSotE1WMqjbuvZnOc7yOdQJJDQRBaliaQGhOztJ3th
hmyjtNDY3wNJ5/35K3m4G9CyxZAdz6P1Kw2aenhjoEBxh7qdm8oCJRfI+9HMMr7ycfwiTq4XP5Zp
HRiGD2pNy/kIj6/kia5wEIT6QQSnhFsX+aLJ9xpj9osWQbh62zlz2nzrI8NfH4wjFPp4cGTV0GN9
04dq0E53Jh6zYW5m+uPkv74iNCh+CRHcNcCCYO8fKZQm8NBOinQxCVDrURF6kC6i24FXCwmHu//f
zGufeLWEkJ2m0Wim6YZvLMwyOR3CubgSnmmGTpihWLZTVHuLf3lThEipzui5SzhT1kMezMVAaQ4I
ewy7O8F54QGcG3WArIR9+5Ui66bk4m2BkVw5VyyugSrYfzi4NsRg8nYptsaNsVM+z0SVR2DMyqj/
IqYu5+KBn4GYxKGALA9MrYdMfWlzZ5LqQBIkyoz1PmYMnM/HqruKN2B0A5dLM7jM4Wul0dLvBBwZ
mgGt7+X7LbGBJKH2Hv/IMmWab3lrz+0CgBtKyL1A8czMMdwlUGLMa/XRmL7lGASVkngtPr4O+jhY
X1qmanq5gLlfhHj66n6+6vKcEOdWJm8n0BS8x/SSZiMf6AGF3Rb/M4O5XK1NvlZUHa/nNXZMTQuU
HOe8j3tluKppFmKjaxqyUNTpgHyYf1B8f1lOnyC5wHkSKYXBobE8+1DncZW/Ax1bX1MGWfTpW/tB
dxsp0pEDzY4uGolZQpXI+Vr/2YHQdOrihz71JryfZuIRKcedX4/3GZlUt+liAQzGMofKrJORrqVJ
X2UNTZVLFFbYW/yE2UJDqkNijoBKFLC5oCQZ0I/g5+dJDnNfJlvj64jd0VsEEUrOtzZwIBippUe6
L8itZnXvB4uq/ZiGnutihGWXEQI3XV06sE3iKI+i8mQ7BPUwlUSSYiEaz6PNxyBzmh9fa1Xtl4pZ
ZdhXEYfdJTckSXzTshuQfjr/9BulhttTl9ARE4Bjz7oc34uf2HRQkv78tu6vy5ioteBEREMjTbCa
qiQJEyw7BlwCu9O/2zpdzovyHfKo+g6Y7FjFvmewdIrjTfKl2L2BMNie5cwEFbujw3lzub3/BCte
IhJJcrYUOZTtzmkhHSRl5N0VNHuT3IUhhsZueggXKMONpRTmWACdA23/AQ2noMXASA8rT36LQcpV
zOZyGPMtq7oB/DTyCvzx3ZjgD8fRBdmt2EetNBzt2/W/1VxtzcpoCC7SWzZaw4y6QLh5YdpxJhq7
idGjUkX0ehY3hyPji8twgKLaZtW+Ok+Pi3pELTVDAWqJvZddDcMKuG2rPEQ4g7Ai7VqxWE+YcFIB
8qAutdA2RLzUVjZ6HtuhVIAS/ZoJ/C/wkg8XaeHy+7NQxh6jodswXfBw5H1nL33179o8iWfhOZRA
eTNeMJ2cBjKwhn4kFumxdGtHhtFNOFfDzITMhAw+aIjtJ14+QfH+f5qEQja9jje8HkGesVSBY/hw
9ZG1YU5FFLfirotnHFtaTMmbfjfpxEMKWCPYxfiD95sac1OFHN8ZsCprVBb6QIjCD6RsBtihKNI+
BZuTg4f1qPk3M/20Cz17O1A0/9lbQdWf+y2HGKZcbtguBhbYCQdxvzxZVrLink/6Zvn/srKSRvz9
GO5vGGO6T5abjJlhcNyX7ehHQEWuYFgMlU53savrX23yBUmxE2JO3jR0tbs44GmM7/yRkBPHNMSh
dbJq7jwuV3CQv18ZPZoxa6jJDMcU+Ubpt1zrHtuh/O1NYMKq7OjNu6lNirT9XAuhvPM+o/ckHHLR
cT45DZY9uZPbtnB2P4CVpH+UsnAiYUfAx8lxx/ByrG9CSXm6gzJYZVKEtUgnMJKh7tOcs82bYtxk
Df5460jsC9LvfO1P8q3xocsPOpRj6Kca1uY7VnQwZRrDBSULIRSQ8HSLfS7wjjsbr01KbZL3Q96c
iKUm7PkOeUGJiPoLR266Swny0wsSR5Mkj0j1xyOCfaUTS2BumAKlJGG4J2orcRs63iYooFPxi3Ln
lIEUGtVYAVKBlbWehL28WbH63jvxfQ+10F/LNdsitMacL2rscc4DCx0O6lBI1ekQ0Nn9eQj/JmuQ
DBfYpArrXWi6N0bbqy/9dUR8JHTP8NLvnafKbFF6odR4Ok0m3ACarlPTLLb03Se6Vz9IQjXv9t9P
OlVriTEtRt9ggArbRWJIAaKuS8/1kJdbi/Bcm+k7uJtF/8wYYnU8zQSLMpjxwK2YbZ8xW2A7xMNG
M60ZC3acTrcXfqEljEbDwP9uWnwP/DLQdTK0HTnQJzCMFlKWGVg/vICF/RGqRell0VoxKN3j3XCm
33G0ljRr0pvpipOfW4mxCagmJlTaDQCGAFTc2GRJ0V/K2eYr6ztpNgnv0vKtOVTEOaK4gi5ywx/G
TH6Mi+1UQIXf+DOVo/ZJRkDBErQX5OYzanz/KwBJTQiQt7k9O0scixP2O3tcXxGFkxsyCYxIIauS
+7cfTRS0D9b04nvC/3WDwtcIT29Xm7jUbEyxuYfN8eFCn13P5Q4Yk5DI0J3llK5/UDTUP6eF3Dhw
77H4E0VcNQCTtWy0jG3wKILPMTpPWZfA2kFYVNZNNcQP3fS8K+OBS8JdfrntMMeUZ6afo0iAPlf/
vNnKN9p6PEb8aR8IddE1bhES0C02KkiLcsnljl3TXdCZaSPKZMQL7hM13ErrXk0PKzrjm8Xrikzf
DcgtEhO2+nOygK+sTgI/i1TCYi6XBrxV2XQ4GTgwV3KA4Rshx5FywMEhfT3t10kZpwhOUVuF0vLx
bf4CgpqBF/U1gwUTcl87OReeb6CiHp4y7ObXZl/q1bbjRNhh1cwxcSQqkcS3cBRhQP8c7vYnsKFW
A5GclhoJ6BgrQdwuTb7ZoCNxCFgN8ui/i4MXzTV9LzoY28MOwZqvXjWu3AhNASL+pboN+pClmm+F
JeM9j+xPZCGjLqvN/au83fomGZr3zc5V+JWVaM1B1fl5Xa+FRvVvBGgBAE/lWCIy4ZvHQBHm5yKz
THFCEm/2Edy5HvY85EFq6JwVBpwMj6bHHcvu7srT1+AaYtszDf8Tf3n86iufN1qiqjdjql+N7SSG
eRjKq+tCMctDKlTqEoABBOQ9nm+pyb0QL7IlH5slRSqQdPa+Yy/ZbiVG643FvQnwqx4FC7WCJMy9
RMKVW5fuBxoCoyMjFZxoQ4SEaouQPi/XVhttEw+VLBcg7TWNA/35+xVbgQvF/ouls9g/NXHQIQiD
k+IWxmZBFbWnSLPFgZrA57Q2inXCU54/6DeKNygW4rvTEH4h4gUV7ORI8MmwDPBA+RMoQe+DEJty
tjk1ABKeDCBGER5PeoCG1z14nEC9cDbRNxwoa7ZABGPDfAlT4tHhoX4pb2T2tVIwL1FtzoBVB0X2
yu4hJhC+KJelm3HKobQY4wyRqj+UummKedM/q1r2y4iqXtf4ckw382TvMW182ZBLOKNqk6aliYt+
4rn14HRcJKW3X3Dou+KdDezmLEPChY6zcHZZ7vbf1wkBgIlhWgHiBhDfkEyhjSvTiV4lDFypq283
Or6AZB6HfJx1RhHJi3UQmBZt2J3PB4WNzAzEEboRszRyTQZs6oeKHePf+9xZl8WojIHjQrsA/bkO
e2llxppd+/ydja4d2LC+7sPdBkleLGyH4GT6RApRQH2s6+SqfFdqC4KNgEfcmKsXspf1bNlBzLFz
x3hlBrqLnCR15D5LNsFrnbV93fsp4JOV6SQMXtYFsSAIAJxe6rycWUgoD0b3F1bQI7iyXaLWZnYW
WJ11ma5U0lIH0bC5lCz0eIKPMWpennw17l3N+ZvkSGmoFVuJotIO5wAoo8GaxmWxgnxQVtFJ4kkL
agtUU7VyNlbw4rpZKUw3QTSegMyidwTpQ7DgqUD3y045o1JKNZItsZnl1pXknKX4qvNLdvdbK5MJ
W3ryqu9dklG5PT4Q9gIIStabM7r571DNzDNG0lO3X3m9Bn+h35jFGYKk7qxQJ54TeFn2LK+zATqR
2D7wNkRR4jgI6Ma03nHKs5G9082+vcQuuWU8omFQUhzo6lDViopXKYuW4qjs317Gn6c94kH76p30
gzQ6cilMu0b5vaw9ek851IMtGclUNw84IcZJhabA1/bq+4vDGt/ZD+ohTN0j4xfqU4I6sr3nErp/
h6lOghEy4OSu/G1suQVU+cjmCqYjUbdBHgVUbj88BIJpl9ZHedKuTD2ZTwAkjE+jjxRKdqfoE+zZ
cNoYSVDORWD6FbdWhuClZnkLZKHq9rvgTORnv26mEVH91v8+1qdfv6pxdY/ZaT+1PVyL5hKCPyQh
OXK0M5H3o5qj8EU6RxmPuf3fSI4gM/W0ZrvRbIvkQy+fcwkYA21BwcHZ93Cw9gL8dr5yv9POcWz7
Bh9YVAokmSNbKIzYWB7HTBKhFXdEKmcqLjbpjsv9HDutY9m4ZFAg2RBcxuXNflz3z0YOWxAmZd2I
YunWpiEmBswdHKbuDqPApB+TVuqSNb3r61QD56OU2CFDpsWQilwn/2qUisi7sxGDOTSlZKQs47BM
pG3+M99nIUbfPUnyACoUkxMrxAjP7d8sTzJ2z7ow5TPPw2iYgfxEOTXh7dxPJa7lqqHIVce1Lv0m
oy+aUKZT6xoaPE9QZHLakJPx4ORHsr4Vf0Ce8ozA1H0Y4NRc7Ck1XdPHMzQEHT/WBM3oJ7nAQ4q8
KsZs3ugEWMQZRoRRU/6vc7YKDf1NxE5trbtDw1VsS0lM7vBur4vM9VmTxbL1LLA1iVPhpY+z6vUk
4ZM+7Mu9WuSQGNiVklBlkhXsQR3cDJEmzbxhh2qGfRn8rtPQbvrLSpx0NqMx3hGWouD0GGS5puY5
Ohfp0yYQro/aEXeOhS2QVtH6Ji5IhvPk0bWyNDS9QKqOq3qMAg7oyVd+KnAmvBzp7SF15irlJKrp
G3p0NZKe/tQl7EKIlxv0I9+zeLrULlDX2Bt7W09db58glAFPkaRLntIHGPuaGfypf7eEhv13S4ji
Bdb6lvTmZTeksN5kvE64xFche1+cCJpAafFC6Lh2fTtVw7xe5QCnft4qjbJxzztu8+nkikDOHnb7
fPY1sbkM+X5AsfcmRCcB7kTJqSppGOd2BNbbCIHJal1L7S/gwAXemb0G3p7Xdb6k6A17SN+UC7g5
MDbauv9JQuvn8eDz9Skw1xtMGoPNkdpowgH4b+ZI/B+1Rx+sjmTqUoM5sEdaysyOecy+QROJlft1
KaKE+xd7goyb6xIcCl/MDVMwjvGrZKjmgHxaiIdT2zufJPbfvN40ADmLCXHV3BBlvtnM3zcyYUyY
KGGKbOpKiPdsWB1t8VdXv9kKsxTq0t9Lpm4dt8amWhfSHZCjFwhlR1Si0Nyo+pmMv8c145NiEMTl
jx9G6rvt/4X+3FjJTLZxsw/W2x15fe73ESPRVvcrSmx9csrr9JSYW1nMlwz+YFMGF61LEuAtm62u
3uwkfkYDRDdXBFUULwUEFgMH2XzQ3apJOGXEit5u8nFITWtqwHvjxWhJR5C78vVvaZpme6y9XfMU
bAgSBNx8lwlZ5s0M71fU7lHMTLVsvjsSnBAvx5L8qCaWInaDDidRAyYunnjJiqPiPq215q5mRJvy
jcn/NKhnGwynVaatpc+s2/uqrbd36jpWzBqZ0c2JNqKWC0tD6w3FnN6Lq47GG3knB4OQSKkhJw6a
ZXlPeNy4ykxnCdScYD7eOt/CJ0Ki9L1bNdR5OZlKFsUFDeSd5rc8mZ9L9+J6ShcMA4iXEr7s3arZ
ffa+kPlXmkKwsZ4nSVlzzqDQTCgK6RAS5srlMtQbyhLsTJWo5hLorTC3P04WR2WH3hQQ7rm+7BBO
iBwVMP0eBO2mQvZyvT8oiOKbF1cHpcCYeiJhpuX000iyERuIdpbMUJWlcnI1aHPsHomXVVSPiDHp
mEu11VkeGz9/PwV6bXFX+YSNBNhq0oRnngsR9/1mXfl65UtlEfl5DQBj4zkQNfrjFGWvxfp9mwlS
upQyT+m7zUd4HVGtO94nzk0uLBUSMDC0C2j1nlpc4Qsd/0ARwjNV2/KrQbWbsZAvjKs/y7XxM3en
4KcIqWo1szD2Mj4CofN2llGDpYqBYKdYoGOZ58jvXLzZ3/okQSjJYqZIYr8gEhVjguQYhhz5wjRs
m5wWKTSLU6+GOYo2kdqJFVXw9K8o9Q1wvo+iEihCRB3e6q6cPFmPe3fIUcEZjTmmsVQv1+j4Civv
s40XQfJLdUZjTLcrQAkKtf0/BrlKa28K7DacM/a0sd97ceik32JDOIGRH1RP9iV+UNDfH4Qogm9/
7EaoD9XtXacyARWGo/yFSoptTLhZRoUV5vi6Z/NQMZvKes9rorGaCmi2gccC1DeF8UAIooqKlN5x
vkKUTd9F4I7c50tKNAVGPv3PRatc/1AquwKFr0AnHBahbvVlU7ab06PwT5ju+NYrbPq+nJt1vrPk
vX7hGWfsTAMncnmjf5idU3NFpsz2cXQx3Fo+c79Mkj7uJCs8ELtLq6+goAXYpOS+Wx1wma8WiINZ
JYdQhdcpsgxcZCHFyemyYNQk+KtBtaf742XdCQk8atqO+8uvPjToRv58jg4/wB6eTAUqChUMCmwR
SNdggGu6Ow3ywP5sEFfjoSUP0dUZ4JzkflBtt2lknxwWzV5TAqO8AVn08On7/xquRe530l/fsOyL
kNBVjkgNCsv4dCprgitm1WczeJXAHEq/DP9Qjy0IsEA9P4fbz+GwoM9p1Jb96Aw5lUsV2v6FqkWo
95hNRBp+Dqr/uex51aI25aYcCwfkZG2Kew7UwshPOtvv+7cksQ4xUSs4H8FtDGhphcuRtPh0jEwY
cRuM7Pr34GMO7iCq+9TAYi7JQ4gJCC/xctLDe4Z6io+XVlmFNMSJpe0FNzApzkg7Gw4OYyEv9UPq
KIZCSygKGu7RxJVEALUMeNQFoYHZBfFUcdR10UILwlwpc3A3uoCqNaGAtMIWIYouYXUCbkpFnPOW
nBN6owjBmV9OdaefVHOWgsFV2rxttvG7TyjBpZwcyvzcVNVP94YWw9w+eYbeX08GRpVr0QpdAUOO
vapdzVzoNExBWJQC6Hsr+YJAFmiw9ycpGnC0Q/oDz42DQVJfGAaLRJBa06Y9lnf774alBqLwwceC
KefjPutPYeV/zM3NdMxc+pKZJhy0u405w3JbzjGGVtmJLPU9tyaZm7TSgmUFEWC2SzBjeg/3mPw+
qhgSPdR50HWq1lUlHRxuQ1oghFvBVWszxl12qEpqibqb355HtNrRBk+LI8yMmL0dNIY5UhEfaijS
XRT187aG11wF2CFmLpv0VIvKy5HNAPdyuHwBAhOP4/+8ri68SXkJFWRJRIV1OXpAfd504p310jwV
ZTN4H1KNuOimydgGElLO0pXU6ea4ddDN04DqO49qXBlxnOyxPe9RthsS7UinWo1xloytOGptL6Z0
8RZ7jHSGyiRFr0QfRH7NqIvepa3pqaZPT9VYBLIohAsjTgnwcnfR6wmPdzqneq65IALFAqUN1y6K
OhjMxDJCdYKA9HsSbDBu32qZ/rYibP+sGmTqNhhNW2UZtP3fWjzIQilHw+dw+0ThX/kxgc1No19s
4++acUmtIUIwvYdbL6E10vyT2R17gpoRc1RHT9OnsX1f5lyv2TqHTQ6f+SugYO4HScq/R9xkHu8k
nV4mJ6KZEW9V3j5fEEXnwxOmpnGv1gyGop8Vlvy/osHIvw+9JIGQbnTBgRKsWG3kgkQwZkFrtSa0
E4VIKFY1WzmOemNpYnqYUTmpi+dAoBMN5lgC48z5Ugk92Gw77vlldK7UUkAKbyVB4MNAv/t4UP+t
PHRed3LUuzvlChIjCxYa+/1zOuAHXlJ134ivwDu66yQlXtu2mT0sm5zT9muiIuEiSQVyWCV4k4vj
CaPW18tfvRXJma00/paSZPNDr193pbje2dXFZ//5xC1m7qisltjZDQsfA+aUXbzdYApvsprLAuF2
e+rqS6iGKPJ+BWaZwPxQ5+ZFWfEeOrZYbGdQh8DGN557De70PY/vQtIkdtilP+4w4k1oLAyOD0XF
qeFLfRprrLOX2AIHjo9u1+9HGKhwARCaPORGC+GW494h9QdhIyb7l+d7gBeT4JKN15ZE+NfaxDke
xw5iR9APYbl/4v9ZaOMHhifTMpcClpg7GOi6s6D/F8w/8T0ru3hxgTCFYhPS7bg31NylTYVdf5YQ
9B/23OZwiPFdKHIEeXuiTf4Nn3NGwedFnlOVYwcBZ9xCu43RohG5pG1GnOXZcNvg5Iom5kG9vQdG
Ncr+3L0UsflR9IDWuLv1a+pecQltlRSTTQu2MPMZukS3MxZAhbo6KvW7ZyhL2rMhwSsCy2xWt6a2
n1jBvfmcU8JcALgCo6txzG6y0VHh+RCp3XH3IKOkhTDWD9zxhPuhlmheAFz1xmoqB6pkpS6NEYo+
SaJjGy+6WOlnjxTItAmZJRAePX5B8PdrepQVqchLN4IOZY8fCqxsomV/av5ez25Ohoq5cJE/jsG/
XwKs+JmnYu/H3g6BQCMH7al8wGNl2vmG+qGsdXHspTEcn5iSWqz89F/yH8cb6ltukj6Svq8S8pkT
4vVNhe2QCrAiBFwgSmELqoO2MDA+JSZYMwP3Q08PIxzukxBMSTpaPjAZi3/GnX1/RXxWrACe4++B
J/2BTZoWAZCq0HDKK8GYWd+oRQoHEsm3JHZKP4Xz+I3/Tt5dvuYx1AXBH6TZmgN7sBGa39ZgsRTU
1KPcMlYxXTg4EN9i2pVi/MHQrE09YOnwbwSrmu0rIkMAGLRaV8MOAW6wW4Z/pAs9kBsn072I+BYI
EyEBuHUNjKK6Z9JyzJMHxeb41meTz5aevf/Zx8BF+Q3qGKuJs/JK0dwwQusqZu8fn0LX2tz6t511
FucTxeL1+r/MPr4hzjFLwQyDNpygNqhr473+gruO9ko+IU57VTAz87w5VFHsR8XFUSJYNfeOE+TX
vcrOMC3+1/0qbTi9T3YKy8xF8b2/ISYCAwKo6KfiNeK6qjtDDsd/E/XcrVODeYA5GX4jqCtDzJR3
MaUAYT44/4c8C1QFo2yqS42+0ENJre5q/Eubw3aimH8rjsGNXgnKvqZQ20ke9GtZfQuTVLiS+frg
TjWIKQ+vV56XQEq5pJ4NRAEIAc4C0VxZurdoTl1jHgLYtnPgqkvhH3+rSlgYhAd8SGFlYXoHm4qT
pLc+BZjPwX/fJY095wIBvjC0IKVETsV3hYdu/+DQduUz+CyDPADDoi7CuUuzIneghhpfVD8OF9e5
O0Lv9jU8ALYiDy7VOGKhEzkkthmOY3SE1Eto7lQs0MlWjbcT16rTlLKgxk42vIiOQeNk1G9+G0CI
9nvnZAFFhoPEgdbwWomI1w/KavQUuAg3ZQmZEkDYSId/LpDK1VT9GDm5c/13GX3b5xgvavJaAqLi
qhOqX4Fo4ZwAbBf/Srq3d1KCJm4KgFz+txhaOnoYJ/xegLGtQJl7vC5VxbFdpLoHCrXIutKpJHYm
MLqiad2S0S5rPIdAjaWy5k1+CUWFMsTWUWbExYvitZS8/nAvb2wXrRmp78f93t0l1rA8O4Kia6nh
rRug3NR8AyNI9CDT7FSWNsme7fSBqXmJoi2aJba+n0f0zt1WAow/tK/y51nK87BFHck5U/lGiY94
lbiUegTuXbrJUiE5hHZA9wG3b/gpOnoaeQEYlY0XxIk2bXP0n8dFeWTmEWLP4fXwg5RI+sqUJLDg
R2UdA/dxUswdMAxiYelV6QDaZRRzdtz4YBX+CHlVNI/rY/fJK+5fTk4wsQNHStey2NKKiy0RIU+X
ONrMUBYKEgGwfXMiA36N2W08z1Z0D/NoHXm837eXCKC20onENWdTE7txR3jAFXufONotzMzPrJj5
2KkCRn5V50P1ooWXC2p4ECUpe0sA9Ol6lId+B4h1xUvKxI6+3i4FRnQ7eVc747HJLToH3wVKz46O
kGPAQ1atUoba3hRSQfLNKOfejCdseVjXmMZ1MqTOLc52TXdNTAjoXqZ7WP5bk6w3aEG1L3skAKjq
Evf8R9pR2h2Ot2OdKzecoxykPa7z8As+qpEs0edMc8+rWonesehe4Ijol3FZoA/EqQKqgGgPQgaL
FuYaniP1i7SN6UPaJPUGBumGwOF6Jt08QRy1V8qlhPVA9yG6XZXbOPooo37jQy6SlTS5c56g/qcV
vJBpAo2US4z9VOf9qNGacFcP8b6ssDFGqcQqFNeR2tYl8c7SJIXMyqzPpnENvKyeOJaAR6DuFSOR
2RdCfMXfTLqgaKa7tVX67U8L8XSXqLhpXtRFvRRokk7W3R04WIe5fimN0RN/bzYTLh1OJ6yIW++l
ItpGPCLHpS5xCwOOuBMC8byo/ex0n/ocpPLrW6zaUBZfNPxGlILDIALYdffwrLXqhFmRXrApmu7B
q3821VKw3/MG64hj8hbxrgVLbaF1tMy/ODUokG3Hw2y43TmOKazeFioB8dHf+R/KDYSKbXQ7UewQ
XklAtB2SIR3pK0VU7r1u1pV1Ry45m5ZU1clgCLrQeZaFyWC5kXaW5dTSvNcakU0uJh+XN+vg96Q1
kFne8szO8SsY2+p5k+4ViE2qVdd65KGOGKJUE1ukKXnDSBul8I5sdqGS1mDpJ+ixxJ7TkcLHQo+4
+KBtulGo3V66CQAVVg7PCyX/hvaIwaHxdRQTo4yKr5FP1Dwex/pnsVrnL4GCIUCMDlpljraUITkI
GctDDzvvYwdvc0o2dfoRJds5hpOIE5VprxRD0cflYv4uQE5OTepJ0XYFu09hkllVcMOCGE6cvMNu
4AFHUi1lo3ARigLb8dUI5FH4Btt6Y92UZe2l+4qMMlkNtUV/+JJ3FoJdTFyS7UBFGu6QU7fzy1IS
QcQmBl/ypkgvZzPA/1bmwqr2ZWf9hgLBp+LLbqCan/7QYNEK5VaK+cjou/qcLXa9swJfuHXuOKSm
5MDIfYOj0UUEeZdHgfcoj87t9NCE6qh0vL7jIIr0HJE8faimltOieeSk0zhEYeMShWoZwWObKXMD
dHfZODgtwan783zGCgFla1POEsA/KneEzqdAinmNlfwqsrXMtzeKfoENJTHsRXdqbAOGdHIOW45N
d5e+ONBBXuoQyj3HY12sbSZj1IRPVcbiJc6OBpAR6ybQQeEMabB6TwoJhUfiSbXYW4S3denmqhaL
LgRtXEl0Sk9A6vXGEIsQd93Q50wOzL5gV9Buf8r5nLbSoEhY3zt5GkI/huRu9/7CV3QccklcM/lW
VeYtmPql0a+ZYAQ1Yq7v4/sQc7hxDUB1bukx0EqUkP6WQunSe+ZjD8YTlBvzea2Vxa9rJDZaVSx/
fvM6GpmblIKzeoHpOd/Ylil7iT0hksQxt3CZaM3nIz/JWndzqngsjcBplk48Q1YCLpG93QFKoeQW
iC3fP8v73Z2aY/yg267carCKZpfSLBXK+iPQSA6pnfVF7yVEtqpvBbP7iPn5ksD069vF4GuurHAC
Hyt3Fm6EDvKwH4ppDZ5rR03GXygMn9bfTSY/X+A8zZsjXLqrulV/2kLdmsj/rpXwEQ51O2RyhkV2
GT6Q7XVEH+sIfjE4sw6uKXDHNHqMj2P7L7u9hswPF2n0tMS4kRWyxo5mebDSVMhT3VJ9fBvjIdGK
XJPame/9oFUpGZUO4CDSWPPxMLBQ7fXFOhQd+a/opFByvXwNJjBppdLER4Z/KPALdD+lTUgbEj/z
BYuR+egjvd1hv4wZacagP4IUVw6ADyllkmJoN7PFq7okptwvk0xYmh/cGfzOW2bgxZuG/uHRuZ2n
0wCFKH2FYXerIhlY77AjKyCkUi98Atw9ibfWu3uCoJ5S5FVUWadG6rjQKZTXTJjUSLGMzAoKhh43
5Spq6r5fUpBhAwE0bZ26MhJvod2ju67r8rX+BucEQ56Eay1HEAW8zjpmAQITwr7iA85LgpYnRb6W
h+op+Kg89pjZhVAMVcHIMQezL9L5cxiwSnyVMru+OoArDOosl/cfsmNCXbuajarhtTkEa6ovIZhu
sLw2xKdmOApDXyX7A1v9u8d4lo15gF4hfzywc0khRp+S7folypRyhTgzBHSyqa938eDK6pGoH/Dp
73uN2L+qcOWEyB/EPd3SnIImVMmxdY1oqBf99W0XPXlSnF1aekbb/JX/iunoSlsAOap1BLAJq7vA
9hbyx9+LuPAtugtMYTUls5wdqz4ZqSEIULaGuk/hk+dgxkC6TuUVatJ0Sg/pGGUNooIz8xMOoAue
fk4x15w7fOV9JrZ5OwxI4/0KeV/hcPmcIOiKEJCl68VSKENX3KWtQr1WXUoLGfMubeEhdjDnltEn
uoidKF02RhroRmvJ0QZVKwn9dS54voOYq4hWkii9j1OZSzl7QybSzjplAixpF/ViWwe6Z2uaLspT
DYy/5KMP4zXDC/Bp59DBaVVQFz4KFghmVWJV/sU4Ca9963CdcGKDxdoRMf9hv0dElNeJJjwVcIVV
k6c0J1K+/pryzDgrgdQTleScSheDR/dzVtLr1BglqXNcQjhYJ1IbfxqrdoclChI2HyFO0D61UFcH
qXJlTG/uDKnqAu8OC2K69Id1Axu1AZukf/fmVM3opKZTapuTg1/HwORc1ZGYuyqVLPteQK1/UgYg
GKnSsn8SCDRKRPnbHYGSfUDhx9iISf48HzTmo4n7pnpB1dsOpj71tl1DNU7gqlv37JBeJbJ3HLaX
GyjANVSp48GbU4UH0iNdXo7ELQjb16AP+CCJ3OcmoWwNYk9ubOrB6mKRUZV/893qhEm9mX5SJj+4
X73WzzOc0DzOQbYw3dT/UpSZyPm0qCOirjw5gurWbp5TBY8/cU3hWMHGCBzXDlfr3VKPHj/7Xtr0
pFoW/QMU1EAUyc+21f0yjBeyJGm7M4pdpjReMfNqshJa18IzIYrLzfUJZfabhLkIDSGQw13pequ4
dBhcEKWQuwfcfqXCInxUBHmOPSCixLgKzrUnBtt/65pgwcBJlRUYVIIZe3CN4TBq7N/6jeFJxQ26
jPSSuBcSFqAQNtZHaaXjwaK6rm4t9bfOI8FkuBB+xXpiYgQTkzgPGMW0F22kPeQzxAnrNIeLhAZi
7TwDRTcpmtGMiPIrjJNCus7n+FKM0tPmCQqxPU/OvEzKPIlePNVpqhv6hqWAlXUAYsJLzqSTeSLY
uZWR1j4z6cdnK6ifTmtLd04tCidV42n8Dq5KM1fDlZsr7R0ZAwQlEZ0NP+GrKM457nOHXRBLX759
cT2QS68w7HJz83d2EEUKw8moGe5TQk9aXfj/42+CJ4dpLdU9hzgjszZK9JFJEi+eTfmGZMEmPeQY
ruD+SowGqgULDKwIh20Plv8YqsFSfPhKG0Vz/L9GxLHuogTC3vGyZaF4OuujBefDaAwHGa+ip9tV
zmaX0UStxmicywKVD4ajmLohm1Fk0wD7x8Q1nY9yoDOdX5xX1oGrI2a1Z1VNHSBUHSLcDGMFeEDu
mNtzHMfF7kr+YR7Q/qVJx0M0K6VMtkACxwKcCNBOQipJmVfFmB07jEAaMeolyF2NVy1N0RYz4GAM
TOiN5jMjb2YCR1mOISGb8Qr0beIFMBPo2hHisxR1tHC1209rc6WVSbhXbPVHFydWYLQVMs5ImIcu
WduihrH4lsrZUZ+LB5RXIoZJLJW0XgpuiIz4C2DUET3FgXaK5mb46H+L3nZHPF8TbnkLoSOkK8go
H0pDXPltJEM9IRvMiF6aptPJ3rfEivtlqTf18+8ofRqyuw7Z8s+atlpNwxcoj8QS7GZrmLjmmsUi
7zHfdtFqkoMRPIinSqqX+ghudSbYc2bu9iRZ6dBNtP6rJWt0RbbaYFxIblQJcMYDCqST/DEaIHqN
75W9jFFLYfjzebdkYrBZm2QhyUoZ8Y9ZTOknMugcO0dswTlLQ+3B4jckzOIG9pGLJPrcFnu3ZUqr
pcs+nGZGvtWAwswBAkuuKajr9DbfZWrPPiGNDX+XsbGQg+DvuzPuj47qfudnqAIdezB+nuyAO95q
P0MJn9BdWK1zJ8Qz8m1L3VeJ6kIDFEgEa2siyL57LhXpzg3ukX7AqK0jLqIVxWhasFvesZw1ApJ8
HSJ1xDvsJXhCVhFix3J/sDJ/WM+I7WIS7YiGc5/ksf6HLHjbpwfn1KFBkNEIjc7sLZqmj+nGpp86
n9Ptj+kpGCs/GiLWmjLmO9OGsl+/AliAHrwsOSCFGRhQlu0AVgJEQw48UF+pGT4r5VLTi6nIpe8W
WvXdAAawdBSg1CaA31S4vea1lY/fgOMv+OFyQhRLTdKXHz+4lTQ06gY/JdSHQluW03/fp3CcNH35
WXQa75bnSbF1SJjTgyS0p8bz8ZQ7P3ijjHXZy9OOzOqfMc385n0CuCMOr0LLzKaUjW3DKTqDKH3s
wsAcI20QrK7Z6FR3INpYB8v6z5RGxiXotCHGkZ9e0M19ra2ZegPWtwopQLMfQsKTjHovUMsCoYA6
pot75/HyjZ1hWNOEBll8cwCKVYwOboBi0t/c1jAN2QKwjp6fDv09RhjScLEKTaJQ20SHzYenYpX/
WdVtuHg0HOtBmd8O0AXBI8hnh02rrPv/SxrTf7ldcAyX3sSQmERlPaxI4NQcBdTwo5WduxsDTVzK
wjhtLnC88qA/yIz5AYm8BLeWkJe5z6PmHjWCitK7ROhCxbmOeso1qG2EgFrvcOP+72KbTf3dyJ3T
Vd7VVXa8QOKutiuLP7zr533/dkNAq8Uf60thsDLMS6ki67CB4uQlq0c5sOFbDGxX6CCWFUFHcWy2
dHQ3oOGXYv+GH4SDRPK5RrICivi4SrrKy9CfVpNUnWmgx6mJf9IkQT7PymZRbm9kTgjLVkk/D2jj
5ZIV31pJiw5gDm1SVQwfefU4sYsqFeiYPMFZVSth1CRERCgOSRR/GNHOv3HEnDmMn8G6OVkZvKU2
GoX0MAewXFPehQjuTi8d5mezQweZdvmBZAVG+PkvNrGeSoR1ADSdLPKkJAWhCuIUayfyQAyclOlD
qd01oVjUHLjx+OYpH3ZJZqdASK6X2igUNaYfXQHBM0isHTEm6/9J3r2FqlbbPbCanWLbXNVJlLsp
IwRUhVjTX5hHaVday5dZyPpRu0zAQCmAus83D4GO7/EnhMmcW58NG8GWCkD/7Uyphh0fmeA4D0Wp
kw9bogcCtTPR7FA783QQPf7rivOCIysDpxEMtp92ckxkchNvSqgBJOuRI6evL/S1raevzx6SkKFE
71y1QL/M1BGPOU/fH+KNzjvgWi69q9OzfWmzxiop+34rF/b+kXmBNj+78pBRoRJBrveIdodYnrUW
xRyZrwwq/8eTG4Gp8imX+PWs/Xl47yxF70HhF07WfljZAwHca5hiBu+WhzlPGZtahBJ8LuEZlsmm
I62al95Z6N5ivhfC7GnunTnVVVFy7D2xBIhNmowxDU6o8wI32y9PsQfKqZRdIzTYMQk+UXT9DILD
3YfYdOqGfQQOXZjN5csM7y/5WtYBqXErWQoq4p9TWyoLLkqarekubH+HXV+oD1LZY2BdJksl4W2G
Qc50ou5BrPm6tP0IWiGPSR64oOE/wxTyUgX0wHdZAH+irgtaZic3tOHixZE779SwxOqoxQLy8nWV
KXTS+poGKOs3fl5mlqwSnpwIA78IeIE5rOh4X1KnsRWCplPVgOdKmt2XrpiAjTipdracio/Ie60T
pt1prZQstMWsu45+FIr2tv9Pxyswz/3u/f14p7DXW4K686yoGzIJoVRnmCdMaaKLy+dkP84e73Kg
z4NsRyJ57FxzsVd9GOYaXMXgZc87xXYvmyq5VIgzEpptRmy2YrHi7t99qFIU8eXWGD14nfU7HLk9
uczFFi9hUSgWVomCu8llsd7KBowjjN7rk9yFdBc/XD8WE+DKOA6Inr+XA8vB9H5qSzu21HO8beT4
nZGqh8saSnyhioR9gjHVyKVah8JZS+xnKqg8tVymC3mpBjJ4MXqaLwQgmeGHFRZ4TLfrLL3QRtzv
llGsKqcWPy8KooQARKsT/arssW3kSbuBF2iX4+XvozItXhMtx8cO4KwR0T2bDtb+BaUVmx6DYV2D
rT6ezAyBegUPayUig18PcW4RoEGSThWsk5W4s+aOPUxyNBag9l8Pnu0b52KjsxDiMFawn/Y7sUng
4v2kb7pe77Pf8FhuBPioIRDtsl2IKOEjBgnrJ/CPRb3KSujyOnQ2zGbxIlD7hBUorbOFRC8J4Up/
Rm6Qyc1c1UId9rUypKkYSEd3K99339kKTE7G/D/15sdSLqO/y3yNGA99eLv68DSBAjfqBMVgx/fD
C0nKVaKn97yUjorM1085IDRi+G9dTmUkunSxLEqE9pXv8aNU3kOkDvv80bAWx0RWGGlu7iosnCMF
i9SLtSaN/7F/JEF4PWe/5vR8mvXUk86T2eSHVZIsrMS7cYhRgda+r0RPeqKe+dtR3cYvDpKtQQSB
3iZFE+3VCwjlNbrDaKeV6orMxCj8g4mmMlvYWlbhDnAWls9gcmCrmCXV06cpoz3f1M+Wzdbt+K94
oD5mUkLB8z2aXzMOX5Tpw9idmFhkNE25/1D1003ZbVMD3rcTF4Jv+cEB1IOu+GLL86IgG6s0s7iJ
BTlwXoHQ9uioo+cBRZFrp2OTZsvUxwvgr5jwcYUGSUbsZ1kvoJsWygHai/PUOYI83DhLfu9oSZbA
b3k17u9mANemb/BNtySi7mZT80sraZFrnaQu1VEAkqOXdwR2IZtbQx3H/EaTcDuAD8KTOwszGsYz
MFpy7llqZrCINu/wi/7aPFnOnWESi+L0gFzcxZCkbQSIBEghr+3PN7R0uM1KoqyVPOlobOoaMcpR
SKk8wMzKwrG29ehAsnLPXFrr6JrudqYi1LSAMmiPFCtfN2UtJbqFoJOf+wtqV5NYoUAVmUsahFxz
ix5NYjXhsUrRnq86DcaPzeIpfgJpiFZ6Ny3o1QNydUAFLLuHg9Q7bT3JW9wwK0xnf6qfD1wO6RYZ
ilkL/XkE5U2xrOcDLqNd5t/hwtaI+BrLLAUfeIidywDG/hDD6YWvx7HCCQMiR4eDqJ6W1gqhRDBe
UeGLwQ0wymVk2FIB7Xdtj5K76B+/e41rd+28eDH4Z5K8DLZcOjhzGkIiTa/ldpifFHK74/OFVzas
e3jczuT+v+38qKBFL2mtwO7RgbMNWI0tyqCaV5x3YUcC4UaxQ0SAny/qINO/gztA/1bptV+cPcut
tBWpkFn7BA/DrXEG0Qy4ehq8m4bnTZEB2LzVNoGlj/Vfb3Kree04WY77HijzgabZ4HZ7wneVFvPB
EklFHOqdhux3iku8bJexEt7erMZCua1RjTTRxiadr2PQ/qL+mTTfxcBiUhdVkZd8sHGGmS6gPZmD
7+8PQgfl73mv5pAued/n6Ep5nqMXorr0DVPbzYfjljoytzVuH2guWzXT50s5CCgorKGXdCEcBB32
lEXxnEeBVHL/73Wbv9dgsy2qVqBsynfpvXZgbkqutgTsImyG/nAtBt+d+i7cAy5a8T6uDnyQ418C
BiW+Km1tGUAb9if10mDO3E74bRTfP9b7IQ2iGawTGwiaBlWYr8N2jsLvp++sKDsT213VXLJM3VVP
Waw3h0IRTmxKP0zCaKmb98+b37iDwAODkzD9oCwpK5qEsU6aSqfoXOhlCs9AjAFXM2xr7rzOFP/W
UqoGoPOE87vCLeG4UHd+VHtpo5188RBbNcAQBr2Z6XyqfGEzczvC92ZqKTL7lF9i8/Us5v4KGi7W
Nz5rLr0GGWeye11jvqRMqQCnTdiEbxPCxDEroaGX+JDpMEhT/CeHGBOKJASu5TqwNWLWeSeEZtyA
L+78LvYc1VwfGf4PJnBBxEZ/PU95jpS/N5ro64mOYVPAwpC5LMi5ZgNg9M/sfXEop1Rg/4AEf4cM
flIL+VICWljfGT1ii8/jzjcpQ4vH1TpiwIOrstWNKbxkvRq+DnQqIYnMncOr4KP4eCF74BQWbaiD
Q4H0+WDF8lv8XinVxUg6bbZzfwZuQ8bhYyZ8gB4hR+BVZ+iqdSm/e8Cfd+5QL2gA0OBPmd50FVe7
O9ArvdRI67svCR/7RSy05O4raUfaWSNQvEnxBHeIqefqKWNjlf3tcT4md1EcST9PZr5vfHPQz4SP
FxGaw5xFeZKb6KNl0f9/aQt5DukkejD7JkLct5pvqL618qfsWNYJ3z3hVmB2mlgT9L4JkzMT87s7
q3o+pIVoJrR1pz80BRvrDrYciDBtyZJukwofjMZQijJYO5Q9O6EcPq8c5nImvYurHBHE0dOxZ/ck
1wO2+LQnbWXi7+khZg/jhcmM0C02M6FAeNQvK6igBJ73Uinb1bk84wrI4i4l0YlQDjaRdifuynTi
g8UnJLBO5bqUYWN6QLH3gwDx/hBlEc2kBROHu9KxEc2Qz5SBLWUmuXKMj5QyBLx3PwPwIG1+rLVt
AKt0RXh2LBbR6I6hvZP5Gj/mD7U7sxbct7SmIQ/ROac0rXsDZM2uqlZI1TYZdnzitmw/kVZWg699
jrKhM04CGiAzc99q7TAXReTebU8Hsp3/cKGAbHHsQPi9xM9tPkpPWn0WyzjyMwWvqZD3pILntWb6
cSpJZyp1DyLtLDdMHI7zV1jfPzwdalfezOtMTCNmvnJjGHaKBXmWWxHmdhqdsM53AOpTNnH1WmGm
YXxJnhmCT+i7/K3XP7AnosgjkBR40WamrW6tPHvIelQMoB2sRvwazs2ToJk2LGaMgOPcUOnmzOdl
gNpY1Qbb6jgUz1ffeFWZ3HX5c34W3WMTBocLE3alF1ypP5clXK2EryGlvUgmP8HTSO1jkeYCAVPk
0dpmNavkbBKAW5QrierbIXpJ6qCxXypvRR/jE0r6SDVrzndZylEAXkhbwRPsLxsd8YMuvW4ckFpb
JDyjxOPPm6X6c1LkZOSNLq1Yx7nhB6cCDOqr0y8/TBNLD2Zg2eJSBmoUBA9faLBn9S9biTtAFCSF
yyCuVwUgZSCGPEcdIYW0i4pRXp7hJewCym+yAKfHMgfT/AyHSmNmHpbGtYIINqm82zl73VtCH4Mf
IOsAKGW5eUG2sIA6Atve8vOigb7++WxwaNziJ0CkBACUncilK71Nux18T0ckO3QydImJRyZeuXe+
RmvfDh59Y00GUDHuKgWByIOeWsb6KHwe/CHxws1axXi/sBimXtS/VRi7KEBMp7f6A8YrUZSRgLYR
iS817qIuOTe4Z6JVzSJ35XvpqBcTPhytGBNX8GE5mMvd/0NoA688GdBurcUP7T8X0RwtjomF2qFJ
rswSozb4zS3SCmVdmlaIIF/ZLTSIer3sADclIjlKHRK17QDivYT4moW6qQmwpALQeYDu4oP19iRl
iU1hzbFhDehoxyWpdewz/JyWYwIxOW5HUJWdhPn3udCs119icFOyIsinr2D+KIpOC/VUGIwxpBV8
siwT4p0Lihmid0NGyyRbhwbbjFjTRXETaOZvJ1iUamz+BSog2kuKoihLjCAMXRZsjvZc09pwDZI9
jQTz1E947U8cPsus8xNVPiVtEbw6l7aDBzY1piCgM92LkKs16phhEX95vmR6IlT0M7zGSg88O43h
GAMN9HaBw0AQyxdCNaiAhKZVe1zfIePEaoyDSKCDN53omt31iTEqKj5XYewbRs30ppAyLCjZkcIp
tNVcoAwV7v+21RjWpqagpyfBDi6KnzjBkBEXsKFmH9ll3Eb3rlxSmdhsARg4u5I8zkQu66WoSDXW
3MYSUR/NQQgPGNXiSVe3Nsk1iL+tKuN1gIwU5kKEwymmB47rdRODdGsDotivCF8m1Z7MExXbvw79
dQhvxhqBnLtT6+sj4Ut/2wvGKtZ2bEQmZWRBEsXz2ddBWQrUV4ziATflYLgQMKn8y88DYmusFz2s
pa5FpzMbqlsC/HATsTWvZeBqbDiBM+/GomGCnBQjOllzqAoVfSwS4yw+eShmI0auhZ34c7QWz8Y5
PJtrftYMVQjtjfkoqruz6EnsTG2c4XiBn/0SZIPBD3wufEFOHZJ0lKaGzQDA+AALqB9qsbkaPJm1
+SqG3+x9qVT7/zx72VKcBPmW/VKyqBeqGElqsU7lchgkIGokIdGR+FJ06kigge7twjsztpey5iYE
nr3Oxoyv6FoJQxS6zk7rg8DeQ4n5ynIfz5xzC9RIxqrbgIBxMsj7vat2Ri/6T692B3MMZ3MgBlc5
daaAAlfFATxF+URi0f+k9YzVY4AsF9/BeigMix179jjR6Mt1i0ETMy7XgAIGALs2hGPED1jLb1xr
VyJK4mBPC+Q47Q4fRtYYCMc7w5B+bYPK6F+ZWEjbA2bDiYD04B+DmTY4DZhQwXZQj73hloHjBm0T
KEckx8NOuziV+OZDGrgTGgV3e+43NY0q5LvemputJzMe37q8oT9dAPqUfePnRKOKDXU+Z47pyoni
tc6ba2PSNO/f7ojtCDM/fuVH6K60JQkf6CbkX2ttxRgs5BX1r96qse/08ZYr5Ko5q45HE4XtIJqu
hf/V0+luWuWpogbRocacKT72hdXFLbZ5hO0M5+2XxCsB8QaWCCV0lsALSlakbpzBA8ViDAGg/UJi
24XRXAld1aucGJCtr8mD0B2MHGd5+GEJEgASVpq5TrkQPWAZr0KkmtLQHIDFWIr0DlEc4BvCrN6+
MoNhCRrXP3FzswZUQFpfXiGDJtULvoYO54VMQB/0Yp9LEeofnhzu3/NV98zdDTS/RzcwCgXjZzQR
3pO+myzTBq/SQXgFpHM8Yqit45aH+CLiXarPt4hzRv9Z5cMYscloQ6mGpAih2JZasA9bif+OaqM4
Urn5PpUTtzZaCU+d9aTyPxP7B/IY8eWdf7+nvS/Y6XhxeujtmzggsyqdF1HmGgnFno3NswXcEbSR
9ronv0ynS0J6CB5Y03YtrfOPl6/zoaAIzJBpYOo/ZKOf41GX7RILGoflCjSIpr9XLmAcFcSFu3Zx
6NGA812+l4U/omXDEVBe+qr2qaMWzntUhtOLfO9lobBA8IfKTCKKQJoSyJsyhjQtYcdAG+ArSN1e
zvZb1UfS4K9jra8blj//c8we3Y6Zir565kwTdnRmQPDra7m9qyKH6IC+r4ARLjZ32ZO6ZTG79d/9
3rTRUfjvOLV0WsyaVfgMP2lLRcywnMrNzoxzKvqoqXEQbhk0Qd69mp0pZOw7DXM1/gFj6FOSiVxq
iNwUMlAZasVhrSNeRNUpos7Gbn6lXfM2FAlFYXk62UpSSoo5X3VcZgI0AC/E0VZc7SZmrZHcTyg5
kP2EEpF/zw7RtZR+za+j2SU3IqqiJWDVidTQg5+UM949qfEFlsqOseAHb4jY3G2FN0UrKYGMa2Dj
5Sc/QX3kSO9S0xob1cIPeeHMkGNSsytkiXZ6D3DbvDi48e4m/4seheWgV6u6n/huozGT7E+VI59s
v6gEj3NCaFyEMxavqpEpw+AfNk1U6hSIs3qikVYI300E6KgIkQP9czISl39qhEaifLbf8USnxUEB
HwLCX8HpQ05g88B6L/XmJ4TVb4LGL9QoM3OdLa0tZ2uUreMaX0tEY6myZ4mw3bd7IOVMYALNtvGA
l2u/JnuH9SEDnC2DBMW4rSgCdnQPMT0MgC84LA8qzd04srmJfjjF47VHuW8M6kfKvc2WtiPGwJpI
V8XmpJIlUx8RofFcIpeHYA+MdFrzDIxt4nuxFMo8wvxwPIr1oOmKDuV/rQGFe1ygTV9GGrryYzBk
QXeiUj1oXdxQNpg2YqsbRTB4hVrvPDsNk1dJf4MlEfZHxUmBDTkHPhBZp120Q2mq4t6nuV2YN7+a
cTw6Y9L8lwXS1bQjiBlayrbdVdDqcHRs4Jg7UaLbtCxbDBHAosqhlgZNYK1CycgTJc2jC/UUG+8z
nZplZstR/tFGquKwXWRuOQu2Q4ApJ3shmzihpV6OvTePtFuEZYbZmJlZBXxPaRQ81oxffHTu/2Uu
1x6U9DQKdpo2jZDVlryuNy4/1MnSAuS2uWJ5kRX0dY/bfmkYQOAs6H7yHNDmkwAlWqi319ktGc2e
307eQthHp1MT8kJCivtP0rCnyJsb5c958FjZFdhGJVtUir4UliRiraO8zo3Rk65sh5cmE6tq1tWS
/1zbHSEF4X8qbyPiXWAXlHklvwCKcen3WeBL09o1occxflvtb4AvPDswUpMJhytkmhfpVX1bxRbJ
8wrwwpQOooK8GGCtLwGeUilKNvsc44YScoFQwiDXTOWh62F/yVyK8SDkBVxlCW8QvOsV5Itnuduc
Sgf8UeAVeTN7dChcbXaAwxTEQPNmA8erFBqZSFYTxMVWFZloP5DrahssbMT1iRw9dTn/t/4v9Ct+
nim+dMjqiq/wVgwVVVHsL6YCvIIiGpoZZNY4cVL7lcWT27DOOdWd9gijBTW8AKLDDzudN+sWxAKv
gl6orxp5REEJn6IQ3R3i0U6Avml5c7Zdfnps1aU7xy1L6RBjqq8Y0HmuhwtfDZi4BWEeQxM0hyvC
dYEftglqF6iN+K6T9sMStvK/32yXFWz4VlaknXeA4GtjgfYot3oo3VBuPQyGRC7Dcrd+AN5FQuz3
tTb81DiNT5ZHklakoxPHlWqP9pOAqzn1Jxx8cp2t1NcUbyb5vPOlOZpPXpOq4J6os7FqIvAW0Whd
NfKz3tUVXQi5F/2Hj3gFF9kyMDxoi4Uq3AWAWqa4cDE/rLOYHyUrmaTH0wmoGDpn64YkwkF55opz
7DY+7s1BcFTOmVcxJrJ7FlpYk8qytkFh/1IYFPwfg8oPFB859Kz/LFEss2KXmn+eGI7qr0zJGBXu
+jlHGMGZ/0RDVZtHwaCfv5GkkCJp77NiQ/Uh9MyVl82VPZrnKpFRXzf8uMqBSOx+N687MBwao9LT
ZRE8ysr2+qVG1oVmkAKtEcRL8JY7qy3V1m9dqGtaeY+1w5VMJ39TMJYkaq70/Lzao0eTTglHgUuO
9sB3AXEs5mUfer5awsBUBTTC1qCEGwnVrStNz5miscJuH4Ttu6piW/yep+9zfMXjG6UcKcGOVrGI
7oR+CbCfQak1QGKbeW+nO25MZeUbUon6RLurUK3O2Hu0ry0LjG1/9BeMvejk5zoS9JA10HBAyM5c
+S9xXoyIZB+NHvKtOGJjfvMDe3QlU1SHh463Mg6M2/68Q5917gEtXJzt50VECtgE5CnQ4vVa6jtx
YO79B9P4ypR/iyEvrORl9IpS0Q8ahC8U2H9R3huwPElSsFOT4JqwlrvCW32se2msMT+TjUK3Z2X4
2VVkDezSW+WUpVfxoW0u09OHVKsZUjLKsK3Pjv2TcYvsA5zOMZj5VTEk3FwEiYqfhP9ZTHJbJbLf
nc/W1hBuhTvTr9bNTSAc4FGIaPYFg9cZEY0WjNLjhJxS3e8ue+kwp6eeY75kCC2X7WviWLvIkqxl
VvQh44Pq1d/jEEJvgAbfPod53+j+ky26M7tg+jMzxszNTeHXeT0rIew9aUmzQ6naXJCQA4vqkvia
h59SQEE2yIM74l5ErvqT8K8j2S+4HickWPBv3R8YzlI6qHtwIg3ps/DSy8id8mbV9dXdUvN9ZfrD
/xwMFe07doXfi5HltNJ8UJf55zJ71VKPH58TXNj2deyTTU4x6tOYUjP0b3T6pDdDhhQJX93GjKh9
H2m6impPfhY60TpCutGIfvXpytvW4PfJtpLN9vvlysg41rbwIULqdMNHAYLMwbpPF2LJ1O/4nQTJ
jUOwV8OCfEanEG2I6XR1yTYkGdx8ks/yDLuDm7BY2cbi7+NLSWvjpRVFuviC/ujzxSdIHBI983A4
lEZKYHRZGPS4kJBwachUCPUIsYFIEpb2mnIoIkTdlY8CEiNP8MWX2ZAxYXaBimoVxtpxD4HYV4iz
U2cJH6xK0ApxCaduYJ1eyjiG+I6rSaPX1zyrPtZ3V5Ynxhx8P9dIpQSz/5nnQBjtPZW/XCrhSPim
yOF3xYyyd3LYeDwXFCMqVK757Az2leGWGf0sDQvrDKYHYd98MvIX2t/YJgJDdwaz3iiVtoPapRjg
9mD/mKG+1bXs24jO2d50m5edPYQdfrwlpTePx3B7DzVbPixtQKcUJBK/rsLvqZE1c15M884Nc4aC
lSFWMrhesswyfKi/6F3B1jCKe27SoeIqjfBaDsqpgUiz9pcscp2H7SSmhBlmvk+QcqdqQYYb7pqm
jJuNmPXhbz+WslnctWm/b2riaxlYkawkOA15RwoSwFQzA55BHRhtkvl564Nx1QfHxAfWCQyWzDkN
vGKkhwZjXEXFlA7eoWx2j+yyz5lrK4UVtX7yR0ZSjYkvLOAN8sucsz6HsA7MC8G9KgGoOySdq2uz
54ZVbnAJsCMk4AEG+tCv+aQ8O2UzHvPc3jRYu6439wrCvT70Ug5Y1GD6AxlIcKIMvv5JxNrNKiXa
ogJNFoM7B0oqVCe4RGWtcM1u6fr5Y74eLziycz0VV4ybkPwvqjHBSu/iPV4jzDTQ4idafrCCm9qb
UYPzlC6oEj1+yj1pcnz/f8xoIsAQNGDwMqmlYFO0RIAdj8QZjxtwmUQuEneSeBM+hHOhbcn7Iu/v
X31EfNFE6tBpcUw9jPXl7qTbFpHegcuoyUqmmM/CD6Gbl2eCPgd7Psj6WkmWCb/lyxaEqnm9pGfJ
I7+toQ1d9XtwmO5hhdk4F8pThHvLWnxk0vAq4uMqv0+H1yhHTxdki7mTqYqw6K/3FC9ggYtjxqNO
nujSwQF2/EYZNs8foAKUtuV2tPKunVmx4bo/nNuWx1HBGcMB5mC7ImNzzppmYBPuhBVLjA2eja6u
VIf8HQck+QrevUHN4Lu5qG1g1A2qwR8msHRBGBgFfoDOM9C8mDCMkJEICKoIPDf9HuykO9xRiIPW
Y866va7mIWgjDZX21gaViH1Jf/r/fdiX5/0W5tgAQkN7mEmqvt9J8Tgu/pZVI8n+mVnFFpmaKzPn
kSjpJOL9pPj7+VHX9tlcVH9QvnIsvcp44xLyBzYsohu6OjdkBzXoIgK2OCZOCM/jhv78gR26yhbr
lJ69pVH47tdSn1NiMngMvYgw3OHxc64c66+eiWBzAzRb1r3hDfeid2XN/rnl+Dy7DLnY/TRK+TY8
UlTlcAHIPo6Rm30kEai33560PHwKljqv1G9plgU1ajFzEWu1xKkni+sAu1/5i9TqX7qkfje8jA0W
einpozX1GLMshFl89GXZWG8Y3ix5LDVn8fs9KF/gEOY6cxZOlGk3LpK53asLKFj0XEtGnd5R/Bg4
vAEAQ99nrR/p/L8faTjUZDGMV3ovhS/7br5cZ9Dx6jXcJknf05AkaP9bAs61fHbEo8PhAZCcbO1X
Y3omvB3vg4bNS3Ko4mRcrj9WL6B58O1tAEvFBam4VoAa4CG1nR0GTjRlod/C+xdW0ebEnxuLS1dm
vF2F3gyMc2g62pK8JVYrZ9eQ10r8cjhvoOFO16OYpR3jgoj7ZNcWh+B1+79XqiLq03gx6zsFsAQB
+H6Olg4kEXoShXDJPeT1ieIXkOqPOdgxK7BFJqHQBwEEA9NKAH0ccj4ZEslgjXOlozaP+MFLPR5+
sFPz21MhONamjsX5olKYJuPmzJkiefTLIi0Z3vL7eav55VAoLRXLCGZcnOvae0IOevU4yFDTmj0T
QNjwE8R6kY/eCAHU5FOhK2h2HYqWgB2TRCP/Op3z8sNEbxaBeSp4yokUV38+YFesc2M51s9nQNwq
1Xn1W7nkrQkTiMGXD6FFfpGo1rClY6GxoHQsjSknuj/zAKVXkBEUlSzcJl0EGc5Lv4C0yxFNlxkQ
gxKTiP8tcaQ0dlCryvwUOkAaZTemHXMYXM47l7wrnyV7QA8HhCZu++gvIJ1EZfU7EN62iais8mxf
izmYukfCVcvshij4I6JNdK1CxGKNcnrqLMigjKxWwMmwFlaAZrLSmg+Fp/7Yuv5BPIG1E/noNxgu
XiVwA83uRLdhcEKzTdTDcImAMkdqQpEI4O44vJNvLOZ+e00fe9l2uAiYueqRP3NcJqkIRZqLMIwO
xi03CHghW/Z3OeZ2selFLPnwQjL6bfD1UnWPQphulahcPk6M4JqpBdagNazylbM5wSOb3F9JjWdC
9RGbYG1eESxs8uZmAjR7CvaszIbE0CpQ6OYL9Y6HWgH5hk1nkMc+hVm41cLPX0swWhQdwRo8Achw
qiqwpYmCY+Xa7M7QKzOsdHLM7m/tHJv8fbu9CvQtGiIWcEoyZprblwdmh7N2R+gmc4hrnq0y8qEB
+evQ2LBuneYNaQZ29Nw/wfgQicAs4kyuJ1xNfASuVPEtUd2jcP5oTptQklJrfEgiisLVWhXnrXMd
RswBTE/dQeHXTBby28Hjy/zmcGmkSapuXUkn/f4ttcjkNwOLSmKQVFGpkefCqLNaduxTEcsgMaX9
4DeHQJOX9i1IOUQS96aQWGjjXI/vM3ILNPMzf4DCbzWO3n4zFTTnOph0AtkAlIPt4RzjLFKaAid3
9hw2ixVe7+ot9RFGaTNWX3+CfO3bZT7AHz6bNVxY8rbsjo5cQzcQcqCYj5YK2xLW2SaPPJfqDW9r
cTe887DnkQtgxHDBsUdVUIXjZK+EIz0t67tzfEnmi4sWYIczYVY3kTi8A7+8Skg7pYvjecJaVeLD
nUgfXfgS/bybPG6ml6CukIRUuY5fwl/rGA9w4jRMPYn8Y8yQTgkOoL6p0n2Gqat9zyVkDP1Mz2+a
8lPhJSBbSzlHMfwWdj/nPhFpFKr5XnwZpPhTWr9MdqXDDKjpIzkPxxT455T39mGONnliL3iQQRTF
1PbJQSlCrCLOSreInd2PxaIazBZJcShEl4MxIxNlz69KMrmSqKXe1uGBNX6+sgVz5CyQtEnxBQd+
2LtOnNECqQDL0K0ze0bivQ0um/HhOOhhIHMF26zkKwrfyeWHX27xetk9ZykbpONUvd5eQ6SixAy5
CKcUIwTk6O5/BfTXIKnZZKbAN1eoeHJnzGGdG6iTDdMZfmpIUl461nLj81i+EN19LB9kMtTqBhEt
MHW8mrHo2lBHpdbz6xv2AQv+71TTcKHspWDjV51OcAr1tFFCtD200XqtHDupRgBZCuiJeXduisZ6
ZnPDoVghljRdoCU71YOU2wont3gmzuJk237Xl3msTpeoMVvrThiv9gUnM1gN9wJexrNAtoYX7pM9
Q9BFu0xoQkRIcAMqd07SatyuzVTPp1a81iR7caV5Nmd2j7sBRpN9LglZVBsIUkjN4SQ+Un0XUTkK
tGk0MG2lGfRt0mH4DzxLBJBRWGWQB/Q5UZclWOqzF/ZuXryfXKZIR2JQxsOes2UOmdmJ4kHRuu4a
M0A1OlhJtSkLHkyYHLt2thCGjK92XbAECLHyoBGpl3gnp9Jf9ZEyLitdFmxdZOjDj6qkRqMmwRYy
S2QhgTOG+FNPjlZrqwN/2GFLhfeWOmzClPa+7aWBH55+3lO7qOz9XB6kwGwXEnrORdJj30DdUs0/
PYcETL+1ZdpQV7qjXOoVbNxNOhUXbP4OiJetIRFuQelDUmkYOn/8V7jAP/PaepBW9zRTUu8moZsd
zdShPR/m72y88bFkhnXNrtMz8u52q+potxMPwhd8+XJfgf8WTLMEtAZcIW5Dmiu/TLTU6dlJM2MX
za0zeBcAG8kv/E7JW5+CCZLhbaC9u3nBsYrEcae2cWWwPeKST1Lkt9AdjCV7GaqXDuljJ2B6VdeZ
7YvI9ZTwU8b/qH9FXiTQ9B5okVj3cEMXHV0WUc9ubc5db89Am+r/F+wuiPVbmIBf9ursrTjlFAu+
F91jNWgKm18QVkBySHxfUmnVmNlzMiOlz7IhKZOVkYYbw2C8V1uWtDB7TQ8EgzvUjeLfE2XpotmB
PIZgiO+4Xj4bOuSkLvpE0WjCYCKr59IqHlsMFZc/4Har2yCp71PyBF9JRlCa0RbkXB+S/VbwGBcF
PqXsbP9cWXtx+Ppfvpciff2yh3I9oKO/3emV9MGUV/kxFT/38a9TdLnCQSVWTT2ENKx0NTqO7tRS
zOG0MVgR7iWNE9G+UWRnTKdMagm0FsFCErgUFABalOVVES0ARP6Jd7RSpSFb+AqKz3btIT3eiR4E
8uuuN3xQMmYbqJFlI24UUaFBE4Bqfl1OSpjuWt0Ob5mEl919yclNklFhcTVfLxH8J20Su7Bal1Wy
IR4hFJaVDGPMlP5DJCE5kkr+WqqTjpo4sFogmcLjuoouqM0xhx2BwPx1YAHGOm4JSAvuU6VFkDKb
/gRTOn/Ahco+oQtuY+BKFbMwEMGL7Gv8f43rMU7M6PA4XzDt14nL+dGaXxdeDgpJ7Sq3bxMTiENg
YrddDH++osAdZBK20VuaWDlfgLlAOkbdWRD8ECVyQbIzxNxgerXxeq+PupAZoAdbO6x4glcurOCK
o+2/vvi58xxo8gCCPy0LJFKX2myiBksSlMhLYGVw82VPZY4wMa+5LxIZ3PNvW/KIXQ44XmufTjqT
/ugS5Ehcuhb9MQwnlmjsJG5u2yDnqGzW7HZDDdphd5YLgr4wdrpIwCrULpJct4HRrPOoMsuXflwl
do2vityxhWY/kRuHWUcms6RQsawLAKfYRtyKt9eRQVfPR2sR3p7DlNpvbg/U3eYBhUbEVcU53XdI
EMOrew907riGuHoETegGCpjvnAsK5YSGO8sJ2jMfASXMimiHmkKMxcZU/HK3sFf498ajYScWadmV
Ek5GHr4U/sudr2WbFgBH1fknCiCze1TGteRitB1uhQmUfv2ZwMi/DawucvhMvEUaphF84pVv1Xz/
77YYinvA7Q++BERN1LKCcQUjAY9xPLx5Y/U15xjg6rO3VKWkXjZWFbBpOdvJX94HJplPTRcWhmWa
CSAT0/qyZ/thp3ukscKjiCyWjHDAXRdII/6dFuJmrmww3NxB7FlzBa7ZzSTNhi0B7XaCcXpBOQ2l
Fr2CP1Bzjf+9cvkTrgEW/yBZ1/n5IiJx6pMaw1Op16RqWVe5pT0DeJ6CN6G/dV+sIW92V7Bil9TW
Qp5pRE5rSmbm4jrKo2WQqOQyUejTSGzOVpRtbRZjhRim1KcbVOizqSCZKSIMb2Nogwnlw0pzIPav
9qfK2ANU9ONs1U32XYgu+tME4C/LFMYFaWaHFM3DcxsYpdKYH7FAC5jiWRYQll74ParoVDZdp0E6
L29Y8H+2PH24W+E5MuRScb9UkYTZG0xsqMhzLj7wD9/PfzYk9ffo6d5xlY4ZfovercHZbWeSo8g6
Jqjheu4l1RxB/CvM04iMaOVtYld3W28EQCMMX3Qvc/P2i1+o6Qes8afbvOgn2Jj/zJ1eMWWF4rhE
1GbycNYHmw3YvphJHxSrDvEAnUd+joU3iAGlB1oW/T7T9BDzSST4nrEV+2XAaBJmaJtQXSV1DE4b
GJNgMY1V0wfCSqPlv5cK+RxPj6YXdqrDflNWCNWGPVuxj2yrWrq5me9xCGAj2uwqurnHNO77w8kw
MYZ3WgXwA51/798f127sSx6PfuGnFvL+p1ytKKDHIMbB8fDEcTjAL0iC+TB4A6bkh4X0ZVzXqdEn
mAkjZ44Hq+LPYBPSDD+JTmA29PS9UkbsMBqhBtEGqhpXu0oG5BddDGwWR+Mlj5EHjDJ9r5IYZja2
V0u7RYXbMjtOcE3n/WUp0pntgXkz1+r6SOLCf9Rm+DeQ2051mtQROaVPkJh22pntjUjfs4T1WjKR
GsSgyeqoT7iPDPZ8a2/noUDkSpTK7u304h2aOYMvGkQB84944VdNwlUe0Uwx/LO5Y5+tGR49dyYg
zmS+hU/qSeslrvrl347L7+h/BTMw1fYZ1QdZVGPCgN5Prek3Q+UbPLszyFXgMw+b7k5jiLjrTOcN
BYMm9E66MjNlYnwKVn9RvU6aQ3syhYMi1YVnQSi3al40RdyzXnJ1I+JYc8fK5KS6MvNjV3nRmYB+
zUYZLxYZ1f79kBkAbzOpvrz/qVDpTF2VUtAp1fH8CMHCyxOHq+Ezas1N/HB6Xm4jrgpIlgX34uxF
UAKyOc6foesQwMrXxxZaOcOKDd89btYLiRGhixrdyTd5mroypxtS5rDC2sdgeow2zslec0cKCbnU
TCbi4ylA3cGWpWJzwQxvVUodPMdI3e8ntnnOWXDii/Pw2zsl6DNDGZ4jLWEhPcauE5wJupy1IZYl
Nt+XbNeVfBhZxHuT6orDAuI8A/pJNsUtbabsNKekb8CCCiPCV+ljogaiXOtY+8zeb5Md90mNho/Z
wurTdKVaXimx4+KunmuBbuG8KJ2EQ7BJvG3Lmeur4Vjvs13Wrj0RXvNnMStstZn4z2Qzi5vhfi64
u5tGc8fB4EgITH00qYn1zs5Db7r9ck7utnWx11kgECMR1afI7+GqSnXQwl++nes+x5ZSyrVZlVCg
OoneNMgaRSh393k1hB3Zy1Bdi2mimE8cNZubWWQjqUaRkyx8JFAWMZN5p/5RVDUDXw+dXM3qosUl
3TabFLOvKQTmQxQAEWbiJNK6PBlTlO4sMNZpkuAQ9FYJDh2jJwdGqp2m65QF61kcbdvk2rJrZ8n5
wyWpkYQLAZSsV6BZDLhbhevuRxEi22A3vfzctgZXlqcjTr3F8fAdOTcWL6sYZEZQBPeLKjDPGLsU
WV+cl++WqpLwPYRF4WPZVdpxD+S2EJkkUmCkZhJWibxT5rtQBga1yc5HgsBBz5mTS2Ie6e8ubufd
ZeBVAWusLYBAOzkxBVvPMNuUL/vNoqZ5Eu7eAcQF8FyXCBqTOLsURzI9/4OWAiQnRpwR5vA3lquO
ikmjRUTUl79Ep6YfkGytKFaV2ItycOiV/okE7yyQHeJKLSRSeA44zsLqcBVmUYoPIhzDTCQXMG5E
eBe7yuT7i/7hEEkRaxhR2AzIDR877Jy9x3th9ekrbZDgINjasVXfrzEWbpCrTL9JhxNrofDQWX20
BdliTKNfEh58myMDJkgncaZ26vHs9nbAS3rKSdZKT0faC42hqeAXP0AAtmIXJYXYrPal+ntuFQN5
32sQhU2lzoMAkmkLNhwV2CW5fK9YsBuLn/YH6zh4YgEWRNkTc9qsBDopJGx97oYnFjXdW3R9QUXj
SvD1U5GmXDP618kQ1QtACb5SPtbdur7mcJjjrEYg2K9fcCr7i+LqpGo+Gw9q8sfxPJhXV3yi6b/v
BGFunRQV4B2lCKdsVUyNkCgUzaM2B1iXh+7KJenF+MVp9a+SQ4U9IulZ7Y1MqX4NdYHcaIdBkq6x
8+v7v/Aa9yOQSoCXHoXHQBxi9LIupcda+9Y7PMKBSRpvr+WwdSX2LGzD1VDG/019WqP27/X+oBjj
muNbiXZOhDjjtR6cQ0oWlI/w14/GvpmyCdjZMMkMCXgs8R7itnPASexldkaqBziNKV0n8ascPKBp
FDvJz4BQIMEiasR1kONtHUGaqLMb8AdCrxuuQR1XtW4CT2WzFJKP3Cbz0ZzIa5cJQLKhFjNw8ic3
QQgDBIR5eGuMjRHNUrESgzJ4Lj5PJW/AIWWfDdBsDMrBGeo5NqkisXlsAJzCBzWi0W1++MRVdDHj
TElriwMdrG9ezIZQTV1TsJIEu2u/NUstE2FZC1+s6klWul99wMlilLB+RESK+aOr/6JPP3bA6YiX
/9JWV4hp50ePVoQgpchYDF9Kl9EpfvpjNNNMhnv3CHVITd4e+99NJnaa2l5u9Q9MN5mFRnSTTV8Z
3krjBegBDbjq/TtzDArYpCG+uiq2KHGicLMwwcYDHSqMKG0bO0ZxVgFriCJS38zWJexssTJLpeG2
p09WuPzdnxaCf0e1Yr8SBcbxAtYqwfrpI/Cfq+m2/kMU3eGqO/WV6BcISkVSIsmj3XGSBPLXnqxD
4VGZdIrZS8KGtxPhS3roHwS6anpi7praS9BL0dXeX5nmB6f7/kND9d4IjhWuU11F00uvCEjIsS5h
td8GuDNBwcNAugJ47dhsPuI7Go14HANWmtUByO8j/EFb9kfmMbvzvsIlDXgRord31bmJ8HbsyNeD
7ROngqeA+NRz0EmxG1UE4CmK7siyK0d2MWI4BCmjn44jl3WF/SChAitIOIkr3Z5lGIykjwGR12QX
3oIjEgPMu7mXPkC73ZBuXeiMPPq951z4E7LLfBdQqjgQo4JrNqBwkw706UIxZEwF7h2WmZzf2Pvx
RfkFe5NmRgrA/WGMhZpT9kdqyXw+ppsXTVhWyxuu2rcVHFo9q7cOMwZUePy0mlroS8aFj1PEbEnV
T4G8kt6enoDnSd8TFbmUQTaFcooFbPvTYHJqrC5tqPnzHnKWb61JHP6O4q1D+V5LoOJcMl2iF7Zo
GWBhmB6m8CniDH7QjVcKUGGjWO5H/xe490fejduaSuGAIf6rrn8RZB0ewhHiy9b7zEV7sY9YTE7v
ROZecZJj2N0QU/f8StZzPnmGrpi4oik0I75jpUJvjoJthng50r+oRVFg/R5fNjbsU2kqkRxNGoYQ
lkGwntgnlHhuyj/c2RJ5P9LlcG26+/fbFgk8flUKVQJQDLHahOJaN7VvNJs81l1F6I2mJ/ahYw0C
tJjaefhOm/SJWCYD0eBY5lAGOR8pf0zwbe7VXx5el7St5bdLpVm6Ukww3KH6BLSgiAk3gxCbUJ49
8J3K+ozJgC/Ubm3SjTLCT6SCnbz2V5tSl68IbWRRA56NAokVMdrdhghDJhTpBcfabOfl5cG1bt6G
l6vjcMZ4gCm1pBhSvvYzVytGXS+xg3Q1HdNue4CiTRZFVUGPQWZ2WziU39UUVpc++ly2bClM5iiM
G7CnwDBu/e+KNSHT+mv7WL3dabdVvvHyPULrc16USUAJc+mVE9wZ36XauaOx5vTvpOGr+IKUjnFh
SCBNa2hRk8SzOPnFJTeIQxHTDzTzmBjn+8Eiolgm/k6v+CzBQTpxku2z193zCnmM7HRn4X5mWeOX
lqkdlRe6tkheo2a5WuEbQAUHIALSPQzJjy4CPx8MmBIhc+Q4NB7NW1U8sKbb8HrJn2/sj4uGhcTG
X7FhYHvV21Vo9PFhBoHPNkZlrs/HEerK9RKpyk+yAf4xbOyXnh4u1JzsoZAyXdRqaatZmiiguC7z
c7dwP/ulK2YwSQZhQuUnU3IM+9Cu08AYKLyOH9gBMC4XoD0zAn4in+0X5DYAkGKhJml1qa94hx++
rNRTwRsG6u2y58nEKPhrMmB4NBczb8mNb+2Dmo2FWWcQAqel6mQBO3cpHA4Ya5gawJD4fM1y3d1b
aD1y/C/IuYeGlQKjh+2vvLDrzlZTomLEmMk44e7QGQQA0oeuCY25u7joplpghe4lYY6ePCpJ6r0q
4SrQaY/r5Di+bimlz7KXbgAQ7YJwv2sTkvf2ZntdYjA8UGVnZP/tUxrcW49Rg9Z9dIkpNbvVD1ny
hEdSfRzHpJpwNK8SZnepST5XGz/M/SdtgrY8zLBx75bcttEedRRq7RBIkbhrT6zc9nRgMoX9rGnx
bnqAyvVS/GQJ2JLW6/0bxWRyOXMTjYINvZhbKetV3AeERZwNyHHDxPWNAAQiA5lY27+rFVwk+plb
JwDfL45HBjY3ntcjrjmkDKSwaBu5QKEaM/U33A7aruB5y8SdLaB5Ueq+GMzlDbK9telDq8rj7BCV
2KnZ0AfT89oKw2E1hMopNi4CuTxudCB8rAOoFf7nQUyojYSjmQv5VE5HQCv/bMQdC0XJSoAxBfbk
sZPqmyHy7I1u2iFWqQ3n9qeUPnwsXoRmoA7xlQt11zusDdhe15xEJtflzwogBOeqmNXGnZfCdfSP
c336Ss00hfme1Df3iFloiia3VFhxtl9wRVU3m33Cg1FDEq4qFwWEwGqri4n3HmXwYC0TopkNNMag
Qa73W/FQ0EOT7Oazt4BSSPbDzA/0K4Y5S1Uj2mDtpxizZYjTOOkkZ0r6IrihUxpW9QBi07WalxIP
ZRPkmevCo5IY6atbSRrwOV+2F43c8tUTyduldX8YM87ODfQp2vrn8527WPaeUsqb1Iv/8rZRJTzB
DmqNe3MF5FbhqZo5M0cHHPw4crdB0iiMyf/YOgurk8Jmi2yi3wIxJG+vQ5URCPazMctapS2cUe2w
1K8mCuvzj/X9SNFYoEl+BLnjy0nkjAJDmAtPtUaB+59RxFpa0Ig4X6lyur6hMAOu11ZUeWFN9P5y
BW28b7JyMj8d1+69VYavSOBGlM5SbCg5rsgI92hqhq779GeZA5TpxfglNRTpTKYBPv9Zkr209CEl
t6T9qB+GEjuBh8P+EgOQJAIjJsBqwFU4w0UA02ypaK2OURma9aSHb5O5KLaJCc95DZ/9cwI2qaYL
+mkAbNS7qzqOrU8UKtcxQQsfoR4OP08+8iySSbeswdsOlIBz8mCG7HM9pxQ8uxviqSjiP9Ldd9/D
dItIyacEv4b4+vnDKhaZAOaqKWX/5MOp5VvrBHQp1udr97Ci7sNMx7uRB8/rn+VBFeeCiZ0G2bdW
nm/ZDHD2ok8mC8B+zlp8Kp4uQrmNxhSY2/vKVPA1U5Om9aaJpP//IHDNd9e0Wn+MVA5oKsmQfGrH
XYxN+BtO1sxGEplkh/RvOwrOZjOBTqOi9KvIxXh0i9TpyYpbfCtw05N61U5MZ+2x1qGWEEJYr/rv
MzmjrC47EmzllsW9S/7Q2e1FGip4NdHEPqnlHq2wo2UMdNqF9sZktAmLDM4jDxwE9XfvgWL/INLa
QqFwKlAg91nNRUSfad+pZEyIf7L/UNu/NyXLgwcf/FPnjCuFrSz6HpuSfUqCwZmysCvapAmX3WWW
CmMRd8Qmcbvh55LCPfJ0PjRP53QMaVn5f8oMXSpqpkSfJYisKyNzdz4gc8gAH4+IzAX8dIqaj6Jb
qA5rctL0b4nevHYGc6bCGFTQzLLbgzxPUcYjPO16gYrKCJyrbUncTxRAcYkRyCgxInhtzc7qq9NZ
JGIzoaEYccjPvAJCEqU6XJp59PrSVAlCByymnLXc3C6ES0tvUn/y28zBCr9B2E/GU/VLLqFmI2IO
B0SWQ5ZtLt04XSjbq5SVqB2ZX2b+pDJdHHIMb1USogcrAnWz95Lofj56eA7Nh3P4BfstmpQESX3h
vvufz3c99Ir9SI567s2GEMH/ONskE3daHZsRLA32e6ZpXx9JKjJnTsD4fHDpzsAxnIon5Hpmbtlh
ulDBesOLIlQIokv/GvnYpb9tUiqKQkhnIj2gJrDMZykvlrxHx1Afa7B6VHm38FAXsXuXNwAmTxNn
q5sqxHmkjOT9AVOzfef6QP6z+yv9vz0sTA6JYvVe7LvNTbYjFSmCUmxM4IA3cYvW4ynmjmACyDOV
KJgOPmRW5Y8S5ug+xhNTfAFK+x6iQIvsA/MnFuutSG75kkWZVPR4wGJxbBZNk5i7l1YOCp5KqTLv
MVXDgOzZfoNigltz186WeBiQB9Gedr+r+zXOh+EGKw/9OpBBNz3hTxTlGe6Syf+jPREbOLR6zrcO
Az+rWL0Mwe2Z11Nzzqu+R1KgNU7xhXOytEikSzs01cGqLglGDa1Jfew7cqAc4KMskEWbfcPt3nsN
R4dGHg6xXNThXEqnWyzudMVCHXyFt4ZPJ8UkbnRSOdcdOp21pQaXIvKbXoX17DjobhW5NYSaxcjU
cyLVww9ZFZynx7zYZ13Y0C9RSRypcg4KHu1T9bOXKo3BQGTV4PuhlpxrE6nYrLi4ax9SonRzfIzG
xfdYlJPWpnhyiTByLqINTJHkRI5lNdKh5N/BgyeDy5Xr1413RbYPKCZgfbrSu2FmIMeizr3g/LHU
yw4bC+VKyCeIguxPlSqZB2vEmn2LS2GDsssgCc3hwuF1X/BoYmy/wpSx2XzpXXuP06arUqEzXED2
Hfo3om2c5v+PCG5bWw/0m8lvZeTVY21gnbnWFSQA3rFQcXYqvODzRyQztMtL/Rs/w7pBIb/Q/yhH
uGYhKfjZTCURTibbzs7uaSCpCD5cTTm1IjigSUPmhPNUvFopmgImsFmKJn77RzWd6JCLbsJig0PE
Ndk3zqjNeof5QGzT1SrdH24RMWSBKVKskNkSuJAVjTqIhX5svaYDOZJjE8J38mlwsdP+prST/Y8e
otaEwbJWT7Dm3mT9fZOvY58g7tFoor+RuN4xPXQI1kSWEVfk/0EuIygFPPZA5dd6b+sf85As6yd1
wljnVhEHMeCiMIuSHCjViGfqBqqtF3izCzNXyxyLN0O2WM8S/xMaeOu9nN0aahmB1MDJCZzOPgXS
54KBGwNJzFespRXpUXmaEmCN4tVbSqKjavaPXJcUOpU0qTexu/bpKR13OvjdSqPRzkRUklDqU0D/
D9+6obAMmYMRvohYpG0AX8zPkqjBof03lMCcP6F2U7Ca5gBckFL/8YvTSgNgsqhKWHklNLcCXuSj
SiXtfM7AXkR7dueFuO6tpBrIzMPQ/DK2QS7gsM9EoHfyZ6GE3tL+l2yKmLZH+ZLhNtrsUnYVXtuG
ww/VLgN2Ml4bVT9M623igbX4XYcZort9cW/swBj34XV8Sfi1pWmRuOsjfvyaNczcB3sySxfVvzCy
EU5gut+mDOWbRTO9T2Kz3PNYf9S7eCbVFkzP+GufiVLGklZ+fvaq2ZpVtdhjaiUyzS+yYaLzvtA2
AC5lMP3KIhRAqjd7Oo9hmz1BiuwVrWQk/en0UF/dctydu2z9cRrGKgnkjL3/KcO8hhUAS6bun3tZ
9QoPQp9aEnKR3AtbbBj0XY7QsCkfiA5TC3nFvAlIgtYhzugvg4SoOhrRkN3y66xtbs489PK1sSAA
DzJA3P7+zOsBBgE6gkt7AkWJ0Kcrogxi3tjolo1QqfZ3xyoeCaenx8rFbtYhocYlR1j/gNAAKV0G
zHJloSHhuQhk8rHW9k33RmmH0ynLk3SV6Qkj61KRK5aBadeA9DuoffHBbhMVVGUNbS9XBXQ0NKCw
GpO9ZtTwAt3p158jXKQCwiQsTXUN5eLnofzW/EC1oaybCsZQO5hvmLQiyqzXAFexEXSe8vpEh0ZG
vfVD61y+ZQAFtMPNAOjN7TZ1aW2cD186WbvhUzvDxPhP7+MX9zO6j2oRiAyNumfE22qxbu0auEXp
wsb/EsFPiHQj3XJ7Osqo6krpPxhkhNptqweyMxYqH9YkfyB4v3np8jTVEfdzYFJGHVpNe6tjpBR/
wD+Q2wRkmHRVtcs9QfpezKXrwt8AtYpQcCdIvGKIFqBhsAZQlFatQi46StXoZ+/5XpfprBNcIiaD
roa5sGjUfbx8kt/kAuaPATGnQauuB1ieeaVZI//td4tbBLVhrH9oMXdeWbmfTj3bM1M2BrOowNwy
Qz+KO/eAn2PYLQmQ8UBVaWAS91TN0J0dYhW6zpas0LWyvZo1gdn5K1XMxhQJOvqya17+wz4gUmBe
k0Gfi3vJyfuscRXE2JnXU+5b6T0x88YUJSFrgHiKH9Suewh75gb0sPMysiOWLgmg7/glJcgRUsj8
sbhnB/FzSlpsx+pCL/Fcm+LapiCfqM7vMcigjFsoMd5u3km4/qiRKngwqEWWwbBT8CVptdxJ+0ro
niVrZ66V9x0jom7HqJrVs7ZwB+P4hpO6QwRC5m7abJxKghYgG93jehyHKpJ60XVxvvKKBzykAOls
JBTg/SfJLBSINuQ4v0zRZbxel5DQqpcLRly7C9jVBO1TxlD1cIAVtioh/jgUfuaOIyCzfwOLCWdE
iXOAWIYbmtcYYriVxds3U8ywbMzeFw1Yx3BwkkoVa7HuX9OZXvuepnN0wZy0hyWqx+f2EiU7n9dv
tUxPu9+uQUETBLe+JVOHieoLCQz80cMunWvgl7DXmMzZAoL8Zjtg7R5liqqs99mde1UQFppocw1i
97C4jOCfsh5yF9+Pcsz8fMNjQ3wkliQEuRuzK8Ssdy+BGk6ko7+kLfd0s/hkVk/vZo4fKKj2Dugl
sMog02ERVnCrXOq5GQrLM0g2yC0rkE6mK9iZjMwwnjQw9ZJlqYGTYvSJH1WVmfxSt9FXMXuq33WQ
SrsasY+ve06bLMkt5zyzBsNRlhzRv7RBfRPeg4X7/8EM2CEEqrafeD0I7TQydewct3G6hug2Fh5x
+dirsP2XcOygPE0j6Uk/ce+PmLdEHPIfhFCLgxTRFYUUPJpmqufApBXNwZv6TNamIv1ky1h+5DzZ
lAASBa3ERIUwJsM+VSP+98G6EvWr7u62Y0mQQYJGSuSQSO9EwaxJaxo7mT2ErwIpRO+fUYfWnXNe
0+OndPFp+RSAESlBKUuS/LYDHtOuxcfj41enj3QqkxqfU09+6+rd10+TDMocZ5EkFZIopGrKCiIs
o9kcbFVgLQfmBohxgePFgniXe9mMo4JgTQru4HHwFrm1e1WQFshrbNiz7MXj8asUet9By1nFqe7S
+MjZW110deQIAj0vIPJUGUx8bFHPr2cr31KmzXrOftoKTGNJeOPkGdYdczLhz100xDicChKp9H5B
9cUJO/bTSEqHz1csxenWAozaGTDK9B5AUujoqvPv2MATllWytTbMM0dwLWSDhX+f+Z/8HriKnIS/
AON9iqEstIQFiDCELEptt1royq1dcn9rEkeKNeQkhcCMc/cTdh8b3GJIgVBSRcbtNwNUhSkWIH4M
74+vkAtrSz+DeLNz3oi0qIMspO0/DzVyfmIHsKQwfnpzZ/eS6neK5xt7rIVMVprP5ZB755lEF4rY
bqJoh72HhGVqo6FpKHmm7LZ/I+ZHRkHpVLVtJwu1xeDdrzW5bKCqZ2ea+E4AmyOKbpYssxm3JSQK
8Pfj8LBb/b08oTOVX1m79vN9NEa7vzpBkZSKxf2CoeU5/yTM54rurcZGnTHySvyujz2DPgcGNulP
/DEbqrmP9n/MxaAWbJ7kIoLur9U6YpDEXfsx0mjl/wcOaLIoyDwWF30/ixz2a+dyD28LZ7lqDRcB
IO4pYR98vDmnmwA4RNoc9ec414kUXSwxHnmhg2EmvhfHtrqLZ3cB0I1qesOq4JZfgj76gNYIAHv4
8NxrTftRQumAG0Ux7ZpSkBJJv+r0R2Rz3OmOlKfdzl7XTd3HlHa08SAQgOb6dztclj/T1geAF9Fz
mPpi+Eofvu2V4S6EDLmMQoRQgGlBiJpFbXw/EmgLj5YebdLnOiQVCyBF9VAO25+o/wj8NNEaIykR
Wpfj53k1Q6/7NpAcXjEOIHNx4AIlTPJOMyGppynindwHVC1ErlqXilf9IRB/FkztJQ1zKFhqjUkT
RcrRraozsusKK7hKK+60nsFHsVQxW4C4z89obnYxFMlTMAi4yju2/Nub1XLG463AsxN2/P60uTjm
91EeiI+NG2NmEdukgNXqfvpuqtGZFxgeH8a+Hp83zlD/H4efzz12Hx1CrG5nstFeMSd/L3dcffzw
lghVOcgoHT4NL8i+0pZtSk+JIUL/9DuxuIYAbe0sokzB8lrSt59AR2dbXy1BjcBpRTkcKpQi+0lT
9BkWysEIJwzM7apxsAdc4qm3EObchU4db0it+g1OJTnFBf96uA81OhE9hs5ubnYYqZqCiLurns9K
tapIFPL+eN8UA+UoYhN40D/ahv7vEoamdpBEBKy89aqK17k/v3uI16sMClbjl5WLcKG8JmZWzuxz
Vqo+u3bz31wzFIqUVp30e23kPzgdDouFnFHNRAWnjz6cWFOot1qhFzJz0oZjV78dau5g4FkCOU8H
ExVahkUNIAu0+eAUlgx9X9dAPnFK4jWy8E7lVyNylpU4G8uEiEaH92LztlgKkJFK0L33/3uogfbf
RiiwvOdLzoCeAVLskG3A6jVqgAgh3GmLxhir4V3cULWewrBDzFddRQapxMvm1sbB3xe6JFw1Um+2
6rcx0I/0v8yKQhf3Gua9oizUL3MCTAiuvCDFy555mxxq6tYRSG9ttMXSxxff6qDqt+3G6bfobLms
jSVYAJwUnARyWL6vzoc6ljGvXynpEs4aoQvKiN7FaxbCd5mv1Ot1fQ0hY/Gei8S0xq4VWm3/0lap
2sFEDgUdx+IvEOTfT6FVWyyR16El1AXTQIBSbxrz3OAHEF3ztJtyTX9pdKh38sPpEmbFohH+9HL5
6zl7p05NCe0vHn7oCQxOjQg7G3upbVllQShyjVzRMJXL3MGs8lL7Le2vSyfvj9XFktNOf7adosu5
nroaFqUxk5UxnLMmFd3iXwaU7rk/gQ0mnL+KRXNjFl5lHgLgldx2erKhmhGyevb5n3mGE9qm+aSY
Yka/QK2fGCJ/3atc0eS9hxVtQk1AegYL2IMHwM7/zvJbfzm0+avuDc7zy4nXGaovWTK0YW45i6q8
vFWPYaiA4RwSXDbm93rZouzU5VtCmOdBoVzcsvBFn/p4IE4XXlOTv2SgRwvzUkCWrTJF+JpEVOhw
75ON7ZbFz3EbRhY8x5c7PlsO9q2rc6T3StoF9tcZDWDtygAPVuMxgjyjhgVl2ke+9Jb9/8fjLupp
+zjrrhiR1qrgzXrIlFEVMSSvWdjQAwwwJeAJKYsrkTGYoVXhlo/qO5AHOCG3E41AaRyIGafEsmwH
c+HedJ3JOCA6tyriAO0sglcGNDw51VEj4gK05SvN0vzHqNpVKkrWnfIg+pJJ6JUY3Faf8vk2Ibb2
NpB6oEPxHde3IdCW8vj16ypNgmY0ceIPDzkZwTPaIwKMOqewmH0InDcEVCfxCWxU5R0mtge5BqR9
FrrP6VjClnJtxs4VPw/VWIgfOeHVzdv2pKbytitHuSiJY1FqXkpaGUSmvKQzkz08ZcsE0cY6Wj0K
FFTTQgOKSeujaT63MBjxQ/igzQuXNEJRmmgyj6M4bVUENoxLNXsf6jRNXhqEuuScTYOGGYobziAb
M4wt0S2+8qNgifP1s+2Oc6QlZYNbu5Lo4Vz7/04ksIvVBxkalZkDQigYdT3QTmvKezVpbXTAvN34
kTqwNLvscoE8ruieu+zKdcfiys7qzQbeV3qeE+pj72ZAN2pvbSqE9FCe1i0/puXnIf1Ri8IwYACS
+/FAW8KRZITM5ONb2OZcfauQnnnVn2PGbmIwVXdSKCRhlJnDSLLSfZfKOwKACuNiskPyRt++6Uce
OHeEnqdkS80mQFdY6QZSOZtVPOmu2FoLLU3K7htGKvwa6xaQto5jZI85suf9PS/+NNI4QC94NBvd
7wYUA4jflbJFWn0aEylhSt+oyrD5DYOLhSCPaP1wXo27o9cNjGjayiWXQXoA5LiDJy2rRIwYlaTw
d0rci8eLkRWpYe3NzMYncbXof4qBssgXg3DKtlbbwS4VOlJiYuS1DNBDSwO8JJrcIxRDSw9lWI2U
9mmONHIYqVjsDHRAeeKF39AXKCTt+gYMGgIqGy6+5cAWbw7OU367Apni4456c5lP1EqOeZYozBUz
ZrOca42hLOJaV9QDTNOHKmOO/Q8iuaME51jY43BS5GUJAOb6MEnyIE1RBCsYStCeCRrp3fXz/5Yh
7O63Dv/xiqIXw5gxLQwvnJXQeA4ed8BF5lYulswJqGcRXEbdPetmFMmSrY39dLK+qad/Ouka0Ou4
QxvjZqVq2ksDrSf9YRA2NqYjr+vGNFyY6vshPDgdmb49eBTibTV2cvxUIdhKU3R9biUe0U6z2a/r
Hyxo0GIhu22jPnHfYsV/0ZE3d0pNH4vWeiCRgYr0sCmMuNSRWxoYJwbOUeuAKf6qC/Oi1ssnQQ5t
7aR7U5i+8hwBrU08Ys8b4wtW2v3zGzLpfbW5pk5ZLEwUMJPa4jC3lMJPQh0CXNKrRMG2fbiugNKQ
kWs8qoGL8QQ/GPYfRNKYR2+Gv2l+GvuFXI9LyQNkP2dakeW5aaB3hAjXP8dmG0bAt8EN0YPE37Qp
4Hh6eEcuW3Q7YbSeLWKK+lfEBcs8SfFe0qfCwKGODpCZSzlQJj6MpFlFushhRhPo+dad1J7Zi9jB
8K/tHdiUH6INJd5U47IHGUWgIW6mYc7lqeq+Z7h+YzUMx06cKlPZtWfkXan2PrE/GuvaVvFrSyZy
eA3f2KxlsbAXns/G7Ucl3t668ho3bkmXXOncJiyzngPBOftexjWQDmAu2fwdjTcJewt+3O+A5VbF
odVvREAvDGZLk5jzq4VX0e7FxDU83OEdHysOpSgPJsLVkvQfSt+2SHZ7IlRc7yH6L7eTXOhPgHF8
Ef8XQQXIjtycIJA9dAljLB3rajYu7nLD4QL7QX4CCvDaJQe0hpEMPBHDIkwcRcOf/EoBE8D2EHQv
Bv6hGspT9mUWVBSzCtw0AyoByZuR/H2DqSiwwWVmoD2GJ8C1qGx0dUlT8MN4eXmjREIhC1MLL7vS
tC033ReHDBQZaBhKlYskxTuMZ/DWkzrtdt3lRyWfGPjRax/I3Rn/+TnKTtAh/z6uHLcU6QJpOBG3
EPjsk5VOiMXboOHnaMNGFrLPQxulDA2bRxy328HYf5T2nLKJjAGLoZYZewrQSekX4TdpiMNM7ddz
3sVNap+Uru+4UKng+VOePnt3Ll5ON5sRnpCzBFRZfGIZKsBdpLMGQGJeddPoJBQC5USAzrtFe1Ya
woiTR3kWLaMCQ1vnGNeCfUqU5X5wddq8WSI5eJwQdFIcDy7NptX/V8vEPypLPknQULeqI1Hg5aHp
ZpoSXdvlp5Q/bTTyZBL1s3CRwU2JPQkQFMZt1IwDfPj9P/FWKh68CIdKU6QEqCBO4xvb3ApDjYIO
H7ZBXpapUKf2WcHmwBCkUCLVaIpQV8P8fpqJDGS4Xk9CdskVIbqkSN8iQqizXL9vOEBv1COedRYZ
FIPiBb9J0OstHh/0oGHx1elw4TGFEuKQRs9LWk4La/UWiV9dwT9BNWW+/bkenV9qa5TzDj5Uwweh
jWb/QvcZaDxs25knqF7qcSSts3ZlZQoMS1wU+fHzrgnP0sKfW+OQo8OPMJb+bAGRhDtIyKr7APE2
X6hrt9VLZQvHfBs7m8xVWIyLbcj+cKtZxcH30OOgYVF9O6vPBKE9uMzL2t8y+G1AZzHcFeX+vQA8
40p3IE+RLUmiz0cxRChCzlDdCzjZL9Bp9YOlnjATbuRrd5BmqGxF9vom55Uy6hn3ZTj/fu7HdGcx
m9iYoLfW4zKjieIbEZuLfQ3lGs68t/+T1HmZ1v5bKARLkgRxWGXi6aRmvS4AeIlL5TQIOWtkBxBf
aOtGI6aSIelEK+oVuaEzVUyBkRPb/TsBVsI+QIFZtPEfp+Y1VxuULeCZ1D3d/OxKXPVhx0vUf9EJ
D44Z5laN/J2PbabFu/IEo2LbKGSLhbwTsC9z+OycA+lfvUME0WPS3XNvtGBgoz6e6qH443PihtKw
N8tlRKXoMj8z6cNAzyb4idzf4vhvn5Nu7sTcpdPmitvbGukYyAorLBUlT+mnO6ayILDz77RbqxgE
wIno4/X8PhAuUF3l1EdGZERZzMv+YU6lBa70zfiOfUio4rvJtAJRpr5BNp5y3hzkJSsn17Au+kb3
JY+uDd0ln8OTmmjux/kbTw6cGsy0wDIYRgPvUNGKxjzL3HW9P5e5ZQnN2vrNH+puyeIQifpExnil
0mMzF5GuJOTWeDWMaxh7gt1XRU8j/OaGcGauDzuxLSk6H58GkP51ZsI1Aux1lkxO0+dCQnWDieMF
MzaoyUnKAAWInEJR8hn3YrDaIdPzAogJHGMwG3JUyMfkP9D5AC2mhNT3KHl7qHa/xUKzscJdHCpu
2ezXTLCWS6ITkWcY0bdYYwnMk7jhh2mAxbAyZQyXFYnjvpl+gBCjxf7nBPXCGn0zXaFDA0t3u88Q
cDc/lCe5kjmVwrjwuWYuDpp6J7st9ziCwMBfyGoR0rFFyRiBblTz7AJOuPtFUS4I3SA2H2Xg32xs
DmLGIhkqWmUXmSEYO1qjFlX0f+c5P2Tmjb7z0NIsZLnFW4Q3Daa4wwl5C6jMBC0nLDSb+5exjUc2
xGrBRlWeG+9jSJoch21/0XiWPqGwevRCfx/vqaIRhXkNcOHve3w5z/I4TBpLCBh2njIVPeWmgON0
jWFi0qkch7H0no78wgyV9G5ICsFR7XBa8fV/gthWAqiOSKNjjCGi4rRsb9gPTjn8hte8ynpsJLoZ
5QBHE6De8rH6zlVknEP+1/zkkitdyeUxCIt0L05UpMdo4AS2lr5hMypRFFLuQARk/qXXJobbEnXS
zu/l5idheACwimd/iZUq0f7t/eQxjQTFv8/6vzOd4sGCN2Rjr/QCFhgsFrqCxYITioNoqLCMjSNV
Dz3evsxm+CCwN+dxBRuZjKv8nG7bQFY7y2Aide9I33+dbhimynKcQL+Ychw7Dm/OxYYCcTKA80mQ
bEAXITWzyLi/9k3rY6mTtOX7IUwgSb+AZ3vlVaCtZogbsUR4M7fv6cOEp/bSIa0Dr0F/hUCPQV3f
z7puc07gt4UtwQW7cQWknQaxQqWfXY/2MkXe8xecySGTmYmNhR6osXxRX2TLn5+C8T0z6+ING3WR
tHPG+SPUR5DffjaXCho1WKu2+dGF5TgJmFFSnu1x0vOoJVjWA4CoOTC50fDkWtMSt6bVGmzI/fTt
I42u5NiJvNi8GO01KY5raev3XVnuHKHQUM1cDFQFUeH0a7dxKf50aDjXlQftY+bwG3KTaq+z6YYj
0cp8YEwxbjPcBL42QLCSHODNU75PBwMCQCHlbFsXCyHpX61mPvViDb8BmLNecZcSKHbAUVy6OBIf
LoEz0q+iLdSMbDYcp55GH33j3HoK23eEXpV/N5kIa73fsbG5Tq9SeN3u8j7kpi5LEBmlG83xf6iY
WpaFX6Eik7PKRPk9JAsaIfZZYMPftGmBR8qmD+5vaUNUDWYrJeSpn2hv+Np6vJbaCYCCUzx7tWWQ
XOrfx1kwCAYmoQhySRM2aROighrlQRCT7gAfDYUvfstvyqeHanNC6TmCsNKp4D6Np2V4DVNEn+Hq
25gDgnT+hlNxvXnRFGEbkd567pqZatd85OTFFjWjdzAStkNjoga0CoGuzuhB2NnuTJtfnyOi4+Ts
+OZZxuEmPiKvOWv5ZaiDotbXpl+8qGJ1pEZ10QwuuQTscDlXVLCM+R76OKlZ2sa3Np+LWXVVoObQ
9R9HnUpQT+4JnYO1yeQEjYGDCFRZbwqNXJz50hxzZUYCgK/BOob7Ie211KtfDnicP/Gm8bL2q3t9
KMHE+KJ9qOu7qDwpc2fOdd0NM6VcRMaIb4YFdLzozV9ZJvi1P4Jh3DjQccxzhIVsVKSx+LfrNT6I
weojaqURLsa+YIODtEEh09RSKHyluZD5RSUNZo/hMYj9zLSMYxVaomFjlG0Igq23Rz43WjwnbIF7
HA1eyRrVSGebqiSBnpNkqmWteLZFDJpfcQNasrnLHoAGr0Urphlfu6bJPeao8kv/flcAf5WO78iF
afJD912P+gfvT7xRSFYo4Xma8dx4zUBRMllpeJ8lSqCufR18nLfA25lxRHSWtRhlKqWoJ41OAoib
X498l5Iu9cz/7nvyp921HkTTdlVuEm99s3t5MH0pLsK+RRepn+LjeIsBlXK/ScM7LfHOhQtY5GNL
70KlxotMC/ukINsPJow52KBjyP1OjNI94Q0bwuKf3GJ+SlACy/f5W9YiDPTixRbkbioqpI8ytGz3
Fb9AKXjnjrWi++4MwEaprt3odPEko+H06NMfFK6JsZ8D/fP7CwrEUQfKzv8JDxfR01ncJ5VE66VW
md6s4J4ABHnTdLRAloZZTg3bgdoes1KMtnsMKZz9uPyarW1ztFRWh/nLLAwOTGgExq3DOjZLCdRD
aaxi07XiuLff/XWgjxcDAYIStfFrdHrk3Uz/RXaxAbWlUL8AhTLKz3DBmy8Nm53goYzu67l99ePI
PvGkAgqojC9Nxgzaof1BgVoYskic/l5s0oKdD9OCVA3jYUd6ihUfamu2E6vyU80dm57v6/POMtdM
W/kAXEufAqJeuq7NcBTsVE1boqBEUD/AN9Y8cyxQ1RMT3yzMOxoWF8eiJe5+oqxIN90maMt+a5hr
a7sDRxzW9kG4tuvmkIY+tSjvTVhO6Jpuf3F4UIBIHP+zdXV2/WIyYWFb/JOMfuBQWV4vuWPefydr
OFgMP+GPbTpc3bwRTu7OSiJ+vdSjw67uEGSeNCNyAHky7g6WN5MFwlk0XXUeJFAK6JR+T6a50tRf
fM0EwyrfYAAIttdIITKGfdcQF0MiiQ4SbB6xUcXuci/bpE+pGOh6PtuNhtl/vTYRn7654h1pUzWa
X2f48J/4riLU0yX3Hxwjz6fIdYg9awrQ05VnSvazObfhNR4CfUx4Ms2AkedPQ1DLiGktyw0CeYkL
WL+I6o/HZeD17F5zjoZ8izV+BUZZlAPnTe3rlQ/cbxMtb0e+NlLqeq+HxJAQ/nmHlf9ejGKvWTEQ
rBPomw9CXDzzrhGY6fQWKX3B84yFkYOmvf4JjhoqRqQicOo08VtEQM/vj3YxgpH/3Ke4NhujVtSN
OeKm0NDPUOgdgcEtSgY/LWg+bcBQbcuD6xJ0aHuxz+JiL5atOVBJYvd1GWgWc7xqBeHIxIzdro81
G8Acua/x20+mkSmwu7jF8Cp2fR3JrlIeJna3nUeUNIKN5nmxor7JHhLjWa9I+59LWd5PSZh72oU/
gUhSGNQH92o24Kr0UjniukU25zwBYLfk2prj26KXOLYJjGo99pAAQp/g08zHPOtYu3FyXokc0Tq0
HNLaQaNEZpQE28coWAUlEypwuTPRsX8gn/WpJ99Z7mIBinGSOtbCqiWud/0SS868jqerC7fSxRct
pI3kBMytSw9UBrdvkfJDYSetUG6HLD/wXwHgqjUpMYjXc0jyk5Hk6QaQUUIRPWH2c33HSGgzzQMu
W06QuvHWjzvTHhDsv/up6jnrpq1pjUoIZGrCxSfLv8fRgxTT170wHWvNjc5hlxF56+XwV5nvVojk
YFtdvsMiK8gROn3WJcJdQAbHPhYdsjL/BtqcdiNewhWDSgT8HLrpaOMf6BhO3Rq7JDsTauLkY6Hq
6vvX9XMA9Qs=
`protect end_protected

