

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fXHYm5mkuLNhnUmnTjiknlB7ZL41SueP42RWxDXqGkneatmPVJHZrei4oGr/dQVV7lKVeR2tQEE3
egLhBxa0Kg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WoOJ65R4pBP+OOZOhxC1/Ed2735KvV3HrXGww3ZEiXLNp2gHGl04MW2ew+hy2RqiCQgxrLzZZtwz
pRdbh3jBqQFcdo7oWNnWEtGSqv5fArZ3t0Jf8qCZ1dnUi88dcI3R9vN29UApTTCS3+qubeOEf8QH
wIIqcHE2KDXp2gACDPw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oMJt+BSOIP4qEWsNLoRbgIL/ulCA7nN9AOXw2+CtDh3AIs2XqQnnlr4QOmZu7EqepQxNWNZnK1gA
sZopQXBz+KpGEwAIgVh9NWcUJXON17xr2aUlhvW4ARJXkr7vVzTMgEp3EXVKXLo0Oqs89+L42sK2
Yxqrvhuau0QAG4kh7sYiS9sFSis+4/sqXZtHCiZV36ZycZQUTJANcriGaZ1h97U6BUKkXdowBvAT
kJnWUXnPtV+v45JVBcDITIasVAi7QUZ4GfLa8t+uZ4N12UarS4ZxybzaRdKfSW2/73D9r+dc69Ca
na7ziQ/qyeNFneENHvetITzkz62uB96evWrBLA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QHGTs/vH4WE3f22R9lffOedA3zPCAjArDOyk+86PQMbaeYkRU7Dh0plpWTAiXHvLVQvws60EcJPg
TqYIV9KRTZ0cyFFu8twpDPoUGVIu3UpOMJY739rY3J7lZ2SYF2I98KoVVGBTkWC9olpnS5XAt8rv
a36oXIYTJKx/DJT9GeI=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZrFFaSR/NK1DnF0szuZH+rS1pjhf9DgJBZ6q66ykE1Fn1eTZtiuaAWnG8ujJz/i0y/B+gGVORtDG
RASaakokHdEMaBKHUknT3mAaCQh7quZMdnv8IGTjsB2Cm18dpJn+x1Q9Y/N0bI80jJ0FWALEJbBr
yzDsyXF/UstKihRI6mZNAvjtK3X4lkn6sOBy0LDsz+XUfvFu2RNNgF7yW8BLlrQw9Q/QzN8aMlIh
5fCSyeiwUUlVyEslh3jvVqDMjKPRFnGh1F2iDlx0FYPpzKKrQSRF2nmyhChcTJOY0l36wYkATZV0
yZkyaYwP3j+wP43g7NhEYQKF3aMQ3blkB3c9CQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4768)
`protect data_block
/3VIyXCMafcWWtmkBsZ1kMsCP1Gy20NUn9VEFl8HX0vo1pmgX/iJvU+14eXPcaLmGET3rM7pKGq8
e6C4ygiDSym2mRndc4WaGw17N9vV+0kPePyN1nIZowzw/LeF1QW6Hue+3DjKWNZ4x9Lwm0eQuQBC
2lnu3Ho7VWNyImypQDSgn4AK0Yx9llLhsXHVeKEg5PdIdkHBvTrlJQCK+LeRVBoUOrP5BIObQrKx
rnNImz0M5ddrnhRH29wCqMXGVq8kso11ZXfqR4gb5ByCufV9+imqsH+XZw0Cb/ALygKiZM/KXuKG
OrwnLkQOYhOv9gs+cmmLIlQNrm54wChQY+UAWm/xyFi3QuIjmTxi86cc0qVFyXuuyspmeXx9YvCy
S7j/tyYIe0PIFHtyHbt3HocckJpBiRMBGxzpIdTyh3/7ypyIq6UyrYs8KcrCV6+DTbJKlXUv0QUr
5niSZk3d28hB495fT2B0CGf9lQDIWG2fyiqcgpxQcRhcK3ucPoF5j3M7J+hYw50Dju//QBbSn4BP
7klAkbs8yxrBXOBsmcYgj3qTNmjQoiIX94aiiejiv3iHrJscSjEbRL9OtX4fEmbqtI2He70JjTw1
lkF4S5RsHnhaNtSNYEI9+pBmHX4/ySmet0bogNMwAFgVU1l8AQ9uWjv8f9hvwJp73Y35HqhWUKx1
FaAx15VOJCS9WFJpHkA2C/je+znzAvYFvCYXNWng8jfj9NDzyMCQjuHN+EzbWImiea7GPouMJsvA
MhaSlFTGpoBVucMH9IsZwhTaqMEe8AC+HfYWprUVqalxcatUXBcpFgsmkVkuQhXiEpEZMPxnTJp2
cNM029enQCdH+qWpvVVTfyNGmBmRIEvCyCZoJ+n4x3Q+5YsqPEZf5li9UDuozvquS5lmCLQUGK/D
vWJ/JrfhqhphMMRsIMEbL+sxGARPLuTy9B/ibGBq0UKxvUT2TXbdJjCubTNT2b2wT9+9iBqOtCXd
KXE+uQNELTGN87m7HVgQ3a1o4ydn6rlT8ROp1eQfASCa2zNugiwODUnGv7JHZ726tb6KKkBP/+RE
VcXwYPWubFdgvrO/GX0yRhpUc36nze9JYHgu+Xy7yYZusthIgjHV6lz2hcmIPFXAOrBRW5Pp7LKJ
69MKyA2dABEIzAarzo5hrf/gOufmwDIFgiJ9CvflsFcNFdq5rDAqHQAGSa/sTs9H2NGFpV5GgIXr
rRbSjutcu6Iiu5hKwHqJuxDCLIjNEoLDVmGrRCBag1pnrf6mGwxBL6USCyD7f91SCM3IrxLUGa+B
hkJ9n/w1od5kpm/Lh+qFf7UIbjEDNCiePIOxaTUdN3bXf1aFw+hw/oyzPfX2QW/zAlGYk8+BFxps
E5tET2TXdozL5vaERpD4Bkd+4caxcleZBOPiiUjxtlnJ1Kod51ACV+CbIoEm+gAssx60x6aAtQGq
J90DZRrjz7+R2A5F1rBa/c4smgIdOXQzOdDFmtoR1jTuztGWWNWpqhbzFxmsWLe5NrF6u/s+FY0w
GfQAV0V0c7uwWTWeLwm6DtXjd9p4+LTShAsJ1eJtZWkgEo33DzlDHv0ZyB8PbUbD4pjF/wxugAiw
kt+iA5lrtAQ2fX2S4JHJ9OiHGASRbDVvHWV//ZV/M7abT8EhQ+6vigi+YnGGA4o62vgobvpHtqhm
s4vd9HPCfw3eg67nsg+fsGrrNSY5EWpfb/gUKtRm01JLS+JQ2XnLHyjnbYGC4g4KMF10ruCwiYAb
7PMnqodYEFBRkZaA7d5Hw4amnoUAbsaJweCZGKZ4Fky9iYVy4v6TvoyxlNU481AdI/iBxftRzS0I
9wLYaNw/4v1fySAkNmRiwWe+DGUs6yiSjSX+Z8d5z0FO3ieWJbDE+dD2Z+QXDVhRzXRx94fDBCe/
3myJ7/oUETBUQjHbS1w28c2TNTUzzH5OkpddPtIUsmEXK0k7sVQhcQex5xPBCM28URuB3qu86LNa
ahuA+nNq26ecRg8ZEjwn1TrAJhLJnMI2VXCLS/80SWEGHdBNDi87ebqNrDehoqHwvHlXXDZYJY2P
6rgh7khZ4Kh0DzMcigJCyE1B3qbV5UrIYmneZL4ys5fSimrADq7nXwo5qMfb/zZFid4K+cgEJvo8
158BT3dfCbz9G+RO7gOuQSi8Ufj1/LcXJFM7Q1zBvMm//uMMpBM1l2ELtuywtRWLRxVE1ngV3fEY
mpYUy9G4qZE6TIAVKE9fNqBDyNCs1KM8gwXFt/IJbL+JDXNazZN+XR7bSV1rTg+KU/mJUN1lQekk
XUd7LQhmr+R5o2psC4S0/iasthFFxzxzKGZ1Bhk0JYTYrzMpu2ubQOIwJ5k46xKvv1vLqQvOMUCW
8ved9zxCkaInLEI71Bkr6wWpUsQoHMgxpmd/fsM1bkJjjLiRtzDoLNthY2xCnzU6QERWsz3HEDgH
ml7nIz9L1Kaknb5cq9PiJ4v+uUd0/f1+cEPTB5JmL5bHqZB7BWvrFOew2xvHHp4ouT5U6RBM3ZHA
QDY4tgQj4996hHhey9esPoaciuQC6NPCuwsfjKBYmlQd1FoLQsAzANCb2ildto8oOrRiruMjPqtG
b6+pPFIsb7U5yY5UoUi9GZHT8a+p5cZDXZ2gjVb8RPTAiadPzeS2iIGIdPJvEn5Oot9hwU1gRwlc
5fVQMQ1Bgdzt5iE5qvavZu3CpC/fbIR9Hk/puKBsPPLlLsCfxnFmgykkknYE3+fDBvLZPoSiw1xW
gHUDd6K7QGpD5nDD2N7yvQL31PA2TgVJozyTpI+MWJV9pZPSiC9AVf0BLbUSVB9gaeBVmBpOWyry
59ZecdGlHsnZ2vgYMqCCcao4dWxsD17u6sdiRx9VE8pegj6PyhM3mCKxCPTqHgkRmPbK8+/qnCdq
kB0d6gzQjhkybi3a3iWdAuo5Hi23HOgKMi5wWQ2nUecAMVJR+g9G4/xpD4fpk+1rE0P6xQkyVou/
5bjpXrdZMFWaaaKE/TBbnYCBm/HAzsjfwILO7dBgmEbWFXQuIwmyfTsvoWxSNDC/UenQXh1JqLot
RmNzR2q4rV8tnjaUmD7rZZbK/OU2oaNGXQz9g4G8Pb833ynH+gONzE87jcaJO5fQCSR9RlSYcgGb
NhkIRXZV3m3w6ShuFapolcSArH+TyTeCsl8jogv4yZBqQ13ILkhX4JwjfHvvKSJ6UjugDnoOcyj/
6tcR1NaO4USIPsVayCKV2sQaOmbzRa2kAuEtMjPTURuSZYz/vqTjIaJ7PBrRr/StWBAsFTEQUZ11
Cdb7J74kIG/NjflBM3wmCoLak4J7T/td49HpxaDDAEoq1fjhtEpTbnVz86uJCnnDJVMQQqzubEJL
tuLzDKXYj8cUkOWyaapgyZTfbEwqueBqX/Q3cjeaqmKqFqrgI38KThve3qoDfOreq+3kO37OlW4c
Z91m3mxOUhUfyXMhilsZQmpSyo0349fX1JK34yrherJI1uPxt5GOEurrXRKrA4+mGh85vAhxWj0B
bSeNCNkhYBYw9Sj0z99szJljMnY3hTvdPyKM5S4pPysxh4MYm7ZwlbqaWqDA/VgbjLfNDcWQiGET
G4Fidm64Oh7DJdO19YM6QqssGGn9jTkc9uEWLTM+gh01V9fuS44nCQHCAQOPwlbCz1d1Ma2BNd+s
jvZetiKLssEOi56aCNAtma0WY8/X5UiSadObEMUiz80oew8Vnj72v54m2RSDyu/ZMF7E9ezUq2UY
oYkmuuOfJkCNSyJt1hTNx9CtLyLXZ4nLw2CdC1E+bP8kgmVxvA4ImRM2kV0H/OtaFUaaHFVFwxrl
GIDRAPkMvxKt5IUQsTkVUQcVLf2PIOSg03ZVgu3q0lGqtQA5RZ9P0L/QpQpStWKD+l1SaHSnrHtT
KaAHKdHojcJ1A6CgGStzTzsZMZAlhK0881L3RjW3KY0sG3fZZaXx0ivjYCQWSih9M3Kqx0p/5kbr
rtsBT79PLfb7n/AXer3WRu4t8qu6CVgVRU6o1TUsCNQLHjMVCkUai1PHzDy+60ontF0T4ftiEtkv
xcVdvY2hBdz1pdvJ2ACCyz/yyigomqGlNRX1FBxgOeY2Y2tJZ9BIeCOc+twoA/q0PUS8dWGP8F53
/oCODsCTo7od8EBVM0/qpawKSpE95QiD/2C99Ztwab+isSyOFT8E6imAXY+kiW6owxTID2H0VEao
FeBBSHAiGAYM1lV7lZ02jaTX438Uq0tnE+RpMHTdXXh+kxkgb4STaXdzFNpNmUKA6FYEy0PznO0l
6kTiFhqTh7s2DHExaopdjlTinL2vFk+UZpSnGPKEfzpvKDUvY7Vwu3pJvxpmFQJ+Ur5jJetAG3fh
eJu/fzzKeRIch9Tte2mZHW3mMpfMFXNWz3P+vtrGuFkmKoMOAy00JAqrvWW+CnnP3ccgVOntQ6o5
Mth9TLt5FcYDJNrYhtEWlsCgaElb8w8R8lRmQ4MPrK2slWxfB5BLbYVEVN6TtLRulu8y1XAFWAby
DcSs6msDsxZk9u7+1GyhBpHlwttaIlfOTCUFhlXbyatIwLfxAacwZcgS+7wRfA+qqSTDk+CzJwGh
6U6b/Qb0NuFV2uzyMV9tnirD/o0WjxFXL6LeZ0d2VzWFh/2QWpSeH3ZlFgiWc0ntUv2keDOtWvT2
4nVLndwdGvHa7iq3dlrpYB8VskMXri6jAuceKyeK2E8q8i3chsEGI0ofQF8lyXvwAmJGpxDk+PNX
KIqt88yOlkqXFrt5v3cWJhZh8awbKCVpKHe2cesdmQu9Qa5E2fKjF6XFgraYuUa4arPLXgT3Dw8L
42wYQ49hAjuj8EUOnwCUMkgUI4k6A0xy5dpOOs2J7HgivsxQnvuhLBnzoCHuk9mWJk690uFkn61+
v89H6jwXjkwbSQ3up/sIqbGjviaRFxEwlwb0CSY0E6IbkARVfEQwBjgidWj9qvfQqe51Avxrq15U
MJ24EPeqwkxqvLkjvIQGgO7hVDehDZ6zT0hPxNesajwzeMNCHYCw7nPK6bMyXVAToPeNL1qWp7wT
KD5H6LmTkzREuvMv1QdrJJZAhScnbgeeYOs772V89M0BQspapbjGrXvKoLMvoYBiWL5ZrHDK+4IP
lhEaLXXa+49N9Iq0Lb/q8GwXEvoEBSa6QGslr1SLvQdNzrObLMlhtLWg23dGcV9+v3uww12MkHnA
H88e9QulW/Mql3JV4aiaNlSFjEYlgzWOQXRZ4LD8Z3OP9IU3AswLBPnoKs8/SsCENql3gHJVAWHV
1HdnfDzyMpKbd35dfOawqXkh32q6bZY6bRfrmDjiDu5O1Hps1ZaH6AdnHvxiqdAxBfXXqneFQmgz
/V6HbBxc5zkqPtw+3LmvjWJlnmSgrBWlP/nD/WZI5OdgR2eloQhOAvMPC1NOzGgwRT4U8yOGcr8N
V66NP5bSBYToTuNqpFYCmo89r50F+S0MwfddlDRedNIbWTODGdfHRXJ6FgT+nSePm7cw9AvigwT1
JKHL66DKGfl9JvJ3ck3kQCjBM2aOTTgm4DPih+LC6DwRi4wHcS1lAQxB43XSEBm4F43D8fPi4qex
kqFMpoULeQh8tOMsJwXlgOWJ0rpQCybj6FKZUHOmT9BIxYcuvDlYfvFGcry1wE2eUTdjIdy/HoI/
fYCGDCiDho5nGwA5dfSuum0GHY7On5cZcR3TFsieSMCvehxxD7r+BIE1ZNv/Hvq45gZyzZbtwAVI
oOwu0SkijEf5hmQypDb9lqvNzM1BtAVJTS2VXUz/S8IiqesiyHSAVxlPmlXVfSm/N3RK40izMoUu
qpfi8ATxvcFDBFme1k5Zv1PtDcQboFfS/U+lmcbLx1ZhWSt1BSsO3l3bVP2mJiu+9eIAw4kajlbg
x/fcGaMGAEH4znCVt9NRvL4ciR2vF3Ndwo9KZa3z6q2vVzpHh0/weJUcUe2yj+6noL276IX14aOz
0rt4Ik48al940C13Fb5caZMPYY9s6c2tr6kc5xjsVEu6x1MHKdEiNuBE7VEKH1XX1cV+Iu1Uqnh2
Cxbl+LZmJP/9VG0BlgBYHks6VBXyvmwkOvKeRWu8CGIXxV8ctfHhL8CIrRTjHx8Xl3cDsPnVSg4f
9/OW1hNCv+sv4S6D5jJZahvRTFdFlY9BVID5MfZgSkGZE3/N3pMGKIcPT4WHg87Btpir9Q91Zh5n
7DKHJVgySQRHXj1F4AFKwFM0DdvVcK6sL9bz/idogH7tq5d/pNxkH2rtzxedyZ18iSYElj/lmOJP
qWa9yV3yuY0Fl4VAHXf3zdBjJTG+thYSItgQECXuQ6xkj+X0ePmuvJkeWWiZUiZXC3R0dy33gKKg
pzc3hzPK3IYngAzIYVgFd+UWZokHZnRW5jag2Aeh9rFxomFGKg==
`protect end_protected

