

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
h9CI8NTfKexOjOkXat5TvvkDPaB4qdtM7uQe4GI6LIjh5E/J3tYhb2kO9frU8JGTAwiNSMc1aL6X
9YMss6mW5Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DIM9e/7RX7iZPW+feNFy7d034FqnU6WUQwV/XeCV+I/y2a9Zum4j4TuVfbdtM8Prw+LkBQP/O0c1
6opchv5jq3ZreAwlr4mo5R26DSPF0haFP03teVEzu6Sq6xtybxeaJRP45ONO4ftBcaqWTCwQ4V9f
StTc+sgWYd6/7TYSYck=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qxmjaeHokRJWMwO00VC0pq5TMV7QGzMS8aZV0rLm7SkhmVqv5qCpQi1aqc2tW+tvmSS7RLLD7Luu
AaH5VkBVHhYlvM2fGMaTMfNaveh0D4KfKF5Gij9WbWsNNwZo/TWDnbbi6bKgMKW7ZfYYuKpwEBiK
DZHY6rIp3DxfGmNgOyfvQ8F5jkErMgL9YDSsm02HD+tE54uJA5xjgnjAv1tkW9pBvOuGeLN9oEeQ
82abAlvnnBgYEF91byxypXRgTEJ51FHyqKi3eC6QHnr7Y9uvM/i85hSKa0OmHcP97uFYOr/sWe7f
VLqYI63YRmM6cE5fWLx72h6h86o3tZfVbMnYKQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EAIc8rA92GQk15pzWEx0k3MI5vFRsZjnBt7wTzxHXZpiKz7k23VHX2uo95ArAq5d00geZe3WYYW/
B8AaRJ0uAyBAeGF586TWIp04c4XWSgk9h9S4Ou22Y/+J2QoYTgtz10A0XUQCwcu+XgZ/WvvGUXR7
hbST0wuFFOPuWuYp3i8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Cp/COvKUkzuJkXNV4T2k1e1WQmur71ncA/lr1KxFRWAZmnMPU9/doc6oIo4o82/gRQdZaW4/9LJL
fmk/nYk3Ugv6nX8GAb7IExJt30Opwho0P6KO83o8uh6mNX/p8RIlQfTZ/8sOuQVMgj0htzkM5KkP
5BjA/wChjtokreXV9KMpJ55grx/NnjWUovk7zeaQemXUFSQzgAQUGHVsZRSzgOZvjnCB24b1u4rq
GCtwV8veCTju5Is1pf2k/pgzdFoLWPwV1jfzmqXYYV9XFlDCbIg3NDrGJqMbbNaPAfAskNUoC2O5
4PEwxUoMdLpkJ++vj+f5Cq30Fpx76m2FWi//rQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3584)
`protect data_block
gL/TZwPXraVqO8+RxMgWnwCgyrcjSkPrWrDBSAibF/rsk6R8GinIXJUI61qirZzca9gEvfdIpU6M
RqurwlyaQoMVss4igDY1ywTg2x4OyVNK7tICK6yV6IUHk+TwfwMokgSdYg+1CT/Z3MdaTmAmqdLh
wOh/3gWsxEeDPAd+dG5YDdy3B+l7GW4vx9vWUJf1+o2iGsZLUqDfNWHEoGJQr4v17EZg/pbtPP5E
ecTNUspFqvLpDtLkP74tDq9YPLdSOBtklitMbjbHQ38NyWNfISptpRBwWqEjefbHlg4PVDU41sT3
DuQU1ueBXpiez+uDRo/Kpg8hjMDY+Q04vm13wJI97dOxCKPs6cu88T1XfatgcTZo99H/rQEjhezA
p2+m7MG7uUgv6h2msSnTFSor/9OD+1CJ4OpGjeGxH5aifvGM4I+mrun0SCIKCcA/7W795WaDoIKW
UaIMW89Iku+h8s8LPtvDX90xyR/2Rlfrj3oftdwN0vs7oPzbz6C7XyuYrx8wZuIMUKQ41tt+qaW+
DNKdcACCJLONmu5U198mgZzdjSi+xqZk7BRfdvO7G0t9oFQPbTa635mYGOixCWQqwGAUUPFoAfM3
meVy+9YOWz0Do1AnOWF6ipEq4BQ9ZsG7PDi6F/6SwtIrJeyoGebXP5+jNouEagiQZMjBoRllP2c2
KAn+GqwYzCZThT76ULYqdjYOIvxHki1d4rWIfReYuzphxZbExlbJ6G2Y6YMJh9mvx//P1JYeLhkG
+oP+/l1MstDka2Ck38J96WF2kK0ld8f4jfYBD6NOsrLsjb1PFUqDSiGFbAKbZKJfFhxDwaaQ4S8I
wyowpkA3iwQRUMnUMLz1z/NhnDYHWyznQo2g6G8d+MpC7efFhqV9lJmysEHSh5HfZMU9Vasuf+Cf
KNkEDP6y9aHqzzz1Rf2QKmK6siNce6Ju5y2MC+cc5iPtfs6JHbbbpZ99i27M/hO6LzNYvORviSOd
8EL6wn6v/n/YRUIoP8H1DvjUH1h+wwsG6cynxqp8hn315J5lhpuyhcI2XDvzqYEBpt6AdKBBj7nR
B2Wio09fsS9XQTtpVMdu51QtRXQ5jx/PdneV4UHdSDPaAqEYoHXJMQvp82IbC7zelrss612U7zfD
82WfR7NoHYlMwJIFDlAb5yp+MnLFlFGuAG0DtoaLP4EBwZgQvkTrS/d8zTgje8pd6l/N4LOLESFc
zQSX4Q89sdRrRkZZM6q1qIA8yuQOpWHAdbtrfp7dpaRrZGK85HHut8MXSFs3k6CPZnGUP9Q+AbYN
GhPUjsqf3RqNDyhHh4p1W0IWDuvfAY7E6Q9dDV8UxN8s1cFEYFuuyH/quzBZW3Bj1VJ22L7+ZxJL
fSUQyUdb1scdEuc8F6RHr/1VBM0XxDJTGW3MfTQoWAYGYbPPAtDgXbUd0NOHmJF3zxVNpOs8338p
cPneAm8B6bCTMFnjkif8RD5o9ARV2c22SvueuseST96QdTPVB9XCpAHo4YRxsOphYoh7YX4iH52b
HZxzVEwAi0TmEGO/4EJ5dMFLCq8eyCKhjIQXRL+MiXviOTxPXiHlX5brwJiOPMDVffCe3wSfZTl8
hnVzcEAhcTGfRPzSn0ErnWxb4XnYt+yvDvSqnIDdqi5x8AydQqk12IuObnLoCOMj9miW6NeBoLmU
4S5TVi3TVu5Hh4ZnDS164vH8chzniy4QaMJuSH+S54bFYfERBUxz8cMtG2aJfADCsaaRwV+6LmtV
/l1fFkooFTY6gwD9FMhRYSOlVlkyZ2snJR3wBjPcYxRaJcCeEnoL3LtG4LkUU5cXn26wNnW8KX88
q7ON0BDegIC14wFHen/44WwrOqObYkS/5V/TNx6CdsmBq3D53OZrelARGEvZO/ylrLS5/SUZkq5r
UVRHoqxOnO3d/a/xp1FOd5+xRLBiYR4tslUkiGXgyHwjHOjgWE8gVtmitJiYJxZqldy20XaxWJ3h
HOzCFdP97mclo6T80rhQrIIWniOgTf7DbQLQgUj64GuR/udma5TAU5nIIwHJKKbYJt87OyxqcXzP
jHxCFn400la1mWWgTreijJlHNa+kYSvowQe2jtccPCufuxydxroK0+/E+TTdqyGH3/fw97AJ+KIe
1yOMaJ7YUjxGTORsZ7HkkdOfVmMAA7oedds5TG7AvR62d/6yf7k4IjqdMhUMkPR7gcxvGDatNFy/
YzABRWFi+63tnqMzqcvAmOHnmJ1GyuW+/zY9Vg5x73mJTAMeN5Tvafkr3jVi2COkBQYCSffBKjgA
Hs6TVTtDZAvPIxOUgHftHWTvoc0JlfZQOEd/D674v8qEN9n05JAqkI70MkHtFdN4LLpSzlORAKw1
dtx80Vw5+njQ2T2Q38GO1OZuzfMZwAdL9GmpwBw1rr8zTA3esDIDcVrL4XMQmFfryXBp+Oo4URgM
JylrzdrViKJ0US5jAs27DB5fHO67L4tGvI1an7w5vFtj+g2K0XenexVqOK72fojs5+jud9g1Wgzl
7L12p6tnaspkSuGBrhhjDW7oKtD3i56Yvalw5r38mOfWyUHQb201BQ93CvqRsGMGpbs8xLPzseM6
xInboan/JSY8ABC7Z5ooUFxWrh+XMXDpDRWjteguNvf3XyOsbP8d/+YGf7ON+fIoyBxyGmG+sTco
qbCbX7ohsOFewtlRGD8tDO47pagS2Vk9T+3kfoS1rizz9zRLwg/dCqtc0f5p8Cfj7oI4t8Q9nRGo
u9PRvQ0sLPkA0XZUkW3kUbj7BusyvFcStp0QqU/VkoAftNTBNMsVc1aDC9iho7Z+9LuashCZc6W3
YdrYs9VDfQ8vNlGMsxbDeoYX6MLwWDTfpkWAeChVLFqrJ25x0B5eNmr5CHjCm0p3GLg4EtJMYTXO
l7PPC2f5qtJYXve8ecBcZNsnmXQvbcxbzUxHFCq9Mcnm68o5Bu8REdo4OersnGPZGef8GQOnIBjS
mdO2rghmi86CpACz6J+xwlxv7XVM7s1pXF9gzx3wUU4h+Xep/TYUtl186fiVkyilpv2/ujPnhcQB
C4NDyr5P1n8WWLkNO/AFLjMW7Dab2rFjG9sj1TAUd0JNTtvdh3KKc5qUq+Fz01yjhjVGVmUr9QJV
vu1duT7/Tv3HPWMaNdWM35PbJri9gT0KvRj6+tHeUmZ8Af2psi4V8jpLpzMvW/3K6Izf+nm+LdT/
jBT8ns87tBcg2nBHLlCrewj6bQfNuX5ul1L6SI8K2sYDkMl6570z+n0630iadL2MlxOKxFd0XZTx
k0pfyn7SEmjrWTNCOAZFqwkVGHcOtNAf+fbUFXSUJSDKpd7Ex3If2Kh6NJkFlU1TKZXeX2/9UlSD
QmFJguLMKsxlQoRpnprmLgwRAFeffebQIQ+pIeVjxf6wV7qpnG0l3tjIQA1vuGzjxBmlr6DztJT1
nH2DTiUG+syabONnj+tH0tFuAUo9jEVNRUtV6jg4kAbEKgcVzjlir3nxZe47DuMUB3BYLD/nwXmC
qMNCP4sRuHhUf8wYoLqbW5LHNGmwSnOaLkf5pWxnbFq/nDK/jBRqapVUMVHngVNy8GVIqIPEllHc
BMK7AhNbtzbtkPUvz6Qv591Fg+h36yTdjlqQTIqAxcZnOFk5seMbZw5e2XtEaxm04lRhxzCGw0TI
SzNwvwu4OjfCLE22nTlGZcTobEeeKFxhEo7KVw+tdhvMRU1i2I+/gy+icTMIYu/eFYWoX774x5dn
Y1CLv5F8dmKem6bEI6z6qfhEJc6xTxbg6QXgRiidl8xEf/7qrRBV+w9hsju9gDUPfDw6LcxejSQX
yrbqkOFbnslogzOisNuK9l806k/HxDzeONG7P2pMI+Dqm998quBuL88AwLrNcW1snuJeD5klBveQ
fgVA8kMknmkmsYNCkWg9PXTjZ+CVPnOzwqCIGZ87JNCuea6e+hVIlEqq4Lm8MscNzeWsCnMpZfmE
/AtQKgHAP4hnQMZSE5PFNRMYZGBfgc4D0boJ+MXXupgl5sSV5ScTUhRK/2S0vinV+RYKQ7pHvUl6
RUvhjISuzdHzbQv8yzD4bOLkxUd6R2mVj0ohbjZT9854UGaN0pM6DV9v7x4S51L5+v87AzFAMQAI
a3fQa8TDRsb7efiONq2Y065Y6Pn8xmIljbLfbT38hY2W0LnUUiTKmBYfS10JK0txu+vaRKyBuHW1
8YpxVw90dJaZ+0OGGqjunLmm//eDSKorpTgevK4xtlz+LWkXShBKGJVcZUIAqHedVPVGFWclUb0b
sfPj8dspu04Qatuv5D2cPrUvoEQ8H/XFfozezDgEAb7rGe11r9wcCUNGMqFETj2/t30n64FfjRvL
6Xm16mh9o6w28qEYLEarAd/Tppr5BC7tILgttjQ7W1cr0So1eiipU7xNnGqd/x/EReKSD0X7diiw
njBQAOA1/7G7G052FqPFYM1DwFs/XZeDkJFnnQj7Ehv6N7ktDpGVz+hEs9N56kIjCxSo4wmrQR19
Of7f1rgMftJ+roh2A58uj2NlCd/4X3NrO5rFm8Oi2dEI6rkYEoxYH/rO6S1szsFd2536Dt8+o2Ia
zZDLq4eLZktEGH0lHlEmg6HVr71U19ewPrB3K6IhgoXGzWOQ/w29wID4wPf4bElsERLmXL3zO3z0
RVh/X/G0+mMywguXevKwhW0sdixgyNW+9qr8CcEbozVLSW4QFhcwDK2kmIsdAcLYTMXpJbKd4wjX
mf+vyl7qMY4JhRCaXEOzEp1xNwlQg6r6oBgFvQ5N8wX4W96+XPv4tdz6UdbYMvhQvT8=
`protect end_protected

