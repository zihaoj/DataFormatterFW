

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g+1wBrOUy4OCkeJr74G85/IZBWxnBFB9soJKvSOOvaRieICQpdUX0CTulhesB1dmYsJMYMCbnopp
tYN9YpIvWA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n84iT50N+szAZCQcYtLz0Z57clA01MSOggD+K8HZ2z6tTDaNLy/Dzn3v8SXkyYI5tc9CeycXlU3Y
iSnLFXq7NMIFsPnoKj0vLtsJAly5uHtdV5mtLOxSz523Q7tlTC8HTajM/mrrDoml0VqIYM7czbL9
ITUwu8cBnpxCbbguL1s=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dUnznpvBSSu0hZtUy44SZBfS6Faz3mUlhM5J71S2XkQ2yZVNSW5eONFgtr0vlY7rlFVvc69ypAZL
6fv1VmI1bL21H4mkIbL7ewQ2tGKVPw1BDIRM2ZuYkxiRy5+fpXyomRLMzECv3VuBbvy4jojM8Kyt
9HA2YN3AhyebtKbrPORp4NH1U5WLQpE3RmJIrjeD10TgE0V5l4yPaJdnNezQuRz7BYI3C7PQ5j/5
r0yhdbDkVOrD61rfUqJpHxjSAhFftZaQJ7UrsK5pyBsxi66irwRVDMW4uVGb3DVs+23HdfRqAOaC
51krPSclz0psOn1zZASNRTOdAcIFHcAigpFo5w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hmIUFIhMIZjZAaXc+XlsAjlpEBdir+X/TkvpxE7FiO6BOB+83nx5yh+7DxuL4DBiIEb4rKaKV4mN
Miuw8btHj9qvDS6iOiuDmTAHy9QWhIfWcPttdcAWHzyC7MMK+L1Bz53BJSs5rp7g/2gPkgO97WeF
qm0B1sVLEiXYCtaK0e8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CoO/0RUodC9gYA0RNACP/fTFl3zJec2+ezrD9qieYPfO4Es/cypdS9Q4wuLwhEZWZoN0B0AgwKWY
ple1VAggBofIuhP4i/jYfWPqHbSypU/Usl54LKobjJWR5+fOwQ6COvNSGy09XqyOALPP2lJgpBG7
a2fCLP3mVpJbCCX7IW5Dr/XAqR1rJxZc1SEnQa5dtsvaY2/NJAslQe6jG0ha7B1cYk9zvMwghOXD
Wu5XPV1lAy+1ao8jUqrZ8HHV4cWQvbFt4Iy7nzU6NeIdrlsmS7K2uFRkBjKwJAyIDXgvFASWl84s
pYSU5gi5GvjeCZHl6h7fOx4YUbEn3ihqgRicnQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16160)
`protect data_block
INFLBAPYYVxmgYn8byer0ifh0AOx55ebn9r1KeHEUTgEkIzpIYjeVpF5aUXjFr3x87iyllNKwWDT
LtNy6j5k0IcH2mNenq6sy5bQgY/2A37Upp6lWHbIUrO/gytGX1Ium7b/tO/Wo0F+czXL9kGPy6aw
eDckvgrBjAnZPXDt4IfhLu8iB2I8aQx85jJHjTtuKI9ArKWjj8+JSoPQEGzxIWm4EUONK2C1f/Qu
c77bwxtujERDsLzSc7RjHzzzcQ6BONTxzWpbn8hWmahIOaJSUAKQx/NHTiTIODRE0qG58ORGlGFg
ofPuBACjw+4vDjGK9rUzMdh28qQiVBvdMKo2XP0ey57TdHFpsz4sqRmOyZfwaQxNREIfjR59ANM4
4CCE6Xk/PNWgDOM+HdRxFNOpvi+7xQmOlCuY0yntsyEoWOMZv59fWARAc+mDFyHiEqfcQib4o34q
lGFasTga88tQQOJhhJfLs+RNbDD0+6lT+aNk3GhQLbgAQ6wjpMwHo75FFqRUBOaSwEpVKoFmVP0A
2YfNKgGGNZxqMTPXlsdGzrPhW0ZXVdWFqKboPAiqi+M8LE64QbhzrmOy/NDdLE/suZMFpFFiDjPA
iYF2viwYrCmSJuO4exTy8Mc4FfZ2C59VCsoXNYw1wSfVeOmPbCDL7aTdatdxmS+0mkw3DYiyh7x5
+0PFwLnoJeLSuLu9kiY/lBD/PxkHcngzKeobcMuXC4HjUFoSotxxIs8dDj+hScnDvOV0HYSK1Hbp
r11Ifm0n9Bhdj/iFAJhBts4izjfuydX6+yfJLGKj/axHPalF2/O4kIVoMFIlSSRRnrmJeYAEBiOB
o68itTFHa9AaWXWxMUfV5bmhTmWMKVhgPqq0V/WtrqLq5dPVf7SCiy4b9HfU8CjbbaustelAWrSu
NOO5+qvRp8HLVarm+8QT03AT8eMEzfPXcM6Pp3a2K9u7BQvwmn3w2KkFUAtT9F5WW0q9fzAAun+A
/6SNKk1CuR1+4jNBjIm3c30jxrmNycX5Kloxz1Kvf/89GoJT2Fp8PPWBYg9cf0sfJKjN8CdWvQOR
37ZhHASWyUQmpT6odeffMSZqIQ9CPOBoi/d46WUCwV3fF5tU4csnlXhWyB1p+C5V174Se7YA0gN0
I3YBrRq1eP8xCxtsSy657BDUWn/5evu4vZDq/YZsyC8Xw2j+JM55jMUhw61vGOLBYJ2wqxax0JeE
aWdGU0kxeIC5nb/O4uRT9BBs19IIONXDvvLfOGknF3jcAXSb0D0sWoYcbC49wsIYPyLXuSDaV89x
BJZcWURgezxEhpygVREx+5uN45Fl/ecyqh2BNf3K2HKx1g1I3YGWxAUJftzHW5r3zZgXf+rCp6G3
etncONcH1qYjOi0KKZKuEoeBCEjk8wXFfRVhELy3PMI6p9/aUsEvd4pXsSHbqJ5VJ7ttOks9ftAA
XH5rnJTf4Er+I0mEVeNqve0yMQmNVPvVcYIsLbNEAyjAg6KB1pXv9QDQdOSKjZtYGx3vaOjUcMQr
eRNSmWIYHViDmEwH8QQLbhzG9eeYvRcxMqOP5ZZyYCptc9BWwUUCLv7hhp0XBdgXTmXJzxkktUhT
oK/b7EuW8359IdnBzdsa9uIYd/krOyGHs/RD+OWq4woj7EdUl6xl1XGQ7504oquYK9HzWF8HjjhF
R1PrsdyF+UcAOqZAIdSY7WBjj9WO5tGd/nIBFH/OUH0KQy8kmSaj/qOdRGlJDstsf2QhPAPkcTl1
0VyPjdBxO/84EzJEOM5F686Msqxf1pA0bxFHKNwXywXvfYQZEVaoOapOk+I7D2+DuSlY5rzdZphU
H75KY7PoV8p7K4WpXGW5IpXpZa3mAZSf49kPW0/0DZsyKmh/5rE4SKmDaqeAAgJ5XTT++IWPszCw
It16cMUbhFDKzHyQpOWPdXTu7BfvZxMID1Sq2JrGLokirZJEvIJbgNkVC+W0iQ6gmMne7CI8oI1C
K9nv0Fr1H63VwiKOHM8j/9IabKx4pNE5vSDi1ZvQy0hUS7SBJf2fZykzGGkZfnJcZhvE4emGISqg
CiVpxC80wt1pXygtK06ZEDGzsbAEt+SzoXC934ZvdbiWk2cEoZ/rY9+1/RumCjfCzGvDxBGJU3CH
FeZd6PnZLzsN7XO2UIJYp7Sr9Pce0lvYLXkmrUuUovC6kGi4Casjvz+Fa8f6dRGJ/BS6D/9tbR8f
X/NmFgZexQcAPzBgXzp9aaxmNvHtEvscgltjBcd6g2PKQMNUAvXNzpnsaDDXxLQh3h71NPAf9YTu
i2y48rpRhGi9Zi0qvVKZ05A7yd9UTi7UlnfVY7LIO7V4KVvHAjd5ACvWOs1kONMkpvQ41YFSoM2/
cXWqh1NdvnCkzFjwYgnnVC6sAn803fx+t7DeRXBV3xyljYh9+EQRxJG3peS9dqps8lqMIyNxxeEY
17Hzll3oYcbopKjQTryiMTopWHkL8Cc4lEpr+GHAe0JeZ6Yu1v406KKD7P9S3ObCX+CqyXzX64zr
ov9hOeWa2E37WpBXz3veoT+OUS9Gzep1vdq36pEkxNbsR0Au9v5NDs50M5lLzkdX7KoNsJZdbvoe
Co8bWtMZrlXiRau5ftT/FWk/wlXyhuNCffy65siXXJDPCVswUkvfjeuZpra5vBh0BnzhvzFkf3GP
fyZ0RrS8RNlQmJ4SuoKTtu3EXsS8V+NEp73u6zvS8J7bwuqiYlIFiH+iHVe4ICkkyKv6LDsNnLuK
G3S6/eFXMlBY0wuedzqq1GBXxEZnmD+eFJAcCdzOMhSXQ1sVLk+Ly+61hKSqP3Dsvd5OXYRi2IKO
lR/USAu2YgxotHbdkBqgFbjtWp4jlN0RZz2U4VUuiNZKLl14ABjOLYav/pz82ar3wHnCtdRVFpLP
EHsALIP/9h1aBkCcCBSTV7ZfPv4RGojp+4ZXWMUEWxLs27+xCouH3w8tWlJtLNiD+M2YeWz8WMbY
BLE9zoJAxOtfDfqiPDaL4WME4oKazPch3FtNEuzgfqOC/caCB0gGorguB3Op0hfrUBrst6pEjqp5
VeZXtK3kZqWv9sm6PmPE2+j7DfGp6gN1XmMxqmBIMekbI+pEFtbKxSCV++17SM6RyjN6z8maV+MF
CgpEXHp2ckimhf1fYjzNBfYXeAW1Pur8X9cQwgpDmoiAWSFOnXVfLKb/Ncy2xgh0d5UYADPggQsB
qjfAytvxtN7fzvZqgDpHDayFxf+ZfmsxJMwdyUy13tOlbtaHyIZHG74lASkSQ2hHEhVDwMsQEUFX
3henypS83T5uAOs4cfHkZEZ22P7f4SPp4JeKYM/I5I7O3Tn29JVQFN41JKtRclQjQ4eiYmcqqtcf
R3t+rjq9VWmGmGupnKBe72W2+r1W5G2uCDTekJRGbT8iitmep9BG2txAxCG3zB5fKG8BrT+QpoLK
2p6tNhwJwLJ9qGkKmeHC3EQUuVc2yPNE2jcmBKfPmg3Fq8sQIWUymkd4KUSVvnaEhADQ+U7LJdv7
Cjf1yMTFzl3hVMyjf42cFptlSjwAqde5itG5BpcJBGb3rtoPJt5xKDWY7tuwT/l98CYqn16foUSQ
J0fGQV1dw95e6RvJLBvzEPRN72Ex+dOvduqF3o8L5iVr89aESEle7Nbc6m6yQB98zjpvYXP7tgAX
BiX97vwuT0GKjaoQXP46QyhvD07oxWORNbbAEPD7TauyKeVbWVqDlxin0pI4U+Mjc/JtxGQ3uaXs
0jPtgA4dVWw/BrqoUR0awB2YzB+Bt07WT3CIq1zxQlCK5rIkdEbG98liHPbHntjClmBT73MF64ow
lHoiVPL7VoqGxGBkJVa4ib1YSXenJy5SQXzliw2meOZ7IMcXtG2KGOq82eJTn8Hr8Gn+AE3tyx5h
xAxLO7o1bbyrsfiYLd+g6C80eZ6PjUQt3Hj72hscT1acBIWUB+l0fGi6HxPh9/YxNAXk8CE0eudR
Qqzbq8uXJYJOiuBXa3UDldWWYHOlpnH3LQV93OvDJzaMFAqwIJW85WY3D+qRoleQVcFAF3Xm2glV
pX4xMly02l6ISLrS0wZ4xrzTQAFejohaUGujFZHPY/A5NSylS5lsbjj39RkzVNqEOR1JREoOfPAq
mr8n2DLUYA7M5J6Y/cma4+kCq77ryTJ3oPaAURYHlBANYtNEGWVkMvdgcCit+rfCKQQ5AIaUZrTe
NhYKTgcgEa1+BcEtUWAMlwdbzVx0lo1grJMwzIr4SkufpFP4l1CCKVSf0EgO3/9W6YrXTfpAUr7U
pbBOI76s5xWRYpn/GSCkICWEgxxqKqVE7Nn4pyjfim3tmfJk1TemNfpW5LG/d6MZJg+Isa4X+mzf
2C9I8FRMRbv1xuy9YTcg6AE45nKzDReQZAyIx9lkBgOd7X94sPdJYcXAXPPvpGLlWcBnFkpyswYM
gE6+rIvUgozHyHmiATJYkf1+VNqQ3a8CjXeUo4VXES5GRNirhEmFBkftDfm5Tt5EPttB1Zp/syj3
IQd2kIlg+lT7hScwNKu1QQQxAfS9FzJQHveSIynUPyIDHuVAoFRDj4wR0vu5RgnHUGpc6pAzErYn
Ya4HtzYGYNn2NE79BWR2wls/ZUNpdPz04nYNi8XDSeg1GXo9Ew+bsDXnM5r7udCL7B6azYXP1lyg
P/Q0RFb7oifA/wLjybDF+KvJ3cOD95WnpD2Hz33l5MocY7V16m9coKDizbZp1kuyd/RTZINx9Rom
f4t+4S5tIWR5e/ZqPFWYRQaJ3ZV419DC1lUGuOBtHjUy5A6+6GsV/zO6SGHe7T3txv466owSLZWQ
rtdew17XtWzRdJBJas0IBGkHlQv+ZVBNo6tZoBtC/NloqCrA0qskGkU3Pd6sCd1+ASKbV846dGu0
8Qd5FEcBvP/N+N/bpBfNaQSg2FnfUG1UWQB2o7cxVAj7jiOYItPCbi/yPrphwi4kVL0qkDC4sG19
JNqbJ+kxmHQ2e6noTPpG2e8V8mpGzXXsUUR/GpxNDs5Rr3ojQTRAkkpzSNF/QJ59VYAWHJE3N0W/
mAikvngC03XfWtBDiK4294FPwt/XiSfJNm0Ppf3Ck7xb3NxEsZwpBEW1SenZFZtwjJFpCf5rM0ZH
Yd0glpUxr1yI/ag5+9IDojFlQI6rnpvASTHJCMCOl1ElsAh2w6WkLAcYhqq/AaAhKIY2e7tzo4/U
7o23i5CZ41VnO36scKLRoZkeJ9rZwwbMnCkJ3guNZZpSG7al6rYeeHHwqKZg/rABOQ6b+ynSVSY7
2D7Sgz2Grr70ybpsZmi4Y2+eEINT7ZnQDx/JoJc6awqK4DcdQpEZ8dgg5ykjQTzyUZayjSIisIfi
rqDfmlzwsLBiWTTeZkYTtlZC0Fq0ph8AfjhBn+8A6HpQ8fE2Z9a17kqd3GLjyoOEei62Bz8cXvj8
boi+jQVW8TU3dyOAIZ4DPWQzTJTdFy9NSm/EDHvE1j9GXbx9SbYEY/4P4UxvHHGj6NctaEd+9FM2
m7hGn3A/JdxCpXs8lksfkFF3x8nHoLc4jZ2ghDXRPnHIiIPleOvg7LCwmzDEQFfIQSriDpL+lzKt
tpiufOkWH75+yyRnezkmekt4FxTEHaJvNHx9gnaWD2TdakZacdBeJ2DdGmtSaqlkU6g200c4MKQd
4z2WcBFQn2Z9O2Su2IkaUOMs0jO0Ud4uFCfjCihlBjxP9qTdXuZYBSMpIG3uABRXdmwIeVG4YAqa
Ky7kPorh0jfY9fHqInrQLiAezKNH7rMcNfNwAjSxoAvG8hC9uljareY6+cDvlbZo2AIp+scgVWZY
X+OztXJlBgiin0Y3Zp3flemYyGT6kxf7PcEEMqE21/U0Vzx4n6hm8idYrFTyMYQ9jPhJ0nSGyUH6
X4DXnI7ngxNKBT+SP1TXMoEajRebfHaazKKfDUYqEc2Dg7FEeKrzyHrI1Hg2kueJE0u+Xb0JOJT7
V9GnOxMWRSPJNQqii7cUCD1dp9Ez0TtsusaMpK+VNtd2yUpcmp5sC/zIPMVwBCCDLrvHOplDBqlB
jzQQhmoVheWbqN6ykZYWi3hvCfAloqNOi9G5q9TV4HRCmTrGFAUGv16YFbrsKT7VeXmJusaaeak4
jnKL/RlmHh+DBbu2TxI0n7Hf8rDD6hJoYIbdwVYjNbfnA6Z3PQcL0pQDNMLuNAaWTEhKzvrVm13p
prTXM74ZHOrt/uDbvvxIJNM9wiavTi5OKlGXR+U6imRdZZfVf4gCQB3QvSqEosTZCpCJ8bqrSMWN
mJXbiYMkuX5uNDL+FLcZozQ0d+uoWQzRPXMEvYGKA6WkuTxj7m1dNJRM42ASyOo1nBc/UoQf9Co7
Qx98POo3YUfdAdvfjv7ppqoxWWncVYnb41Cb6cIy+jHZfJXaz9+WhmSGCNl6An2Kf2Pfgvxth92x
7R3bef7c6Su3XIGN/WAWCsJkGL6swU6hYiixyhxdz9t0aEquSxvGh5231tSHKFCkXE20jk+lRxIk
eQkDYRCSsF36WzJCGGiEnAIiwDivCKKBsMpNSkowIU8QDUpgiLpISGpTl09EX/z0RzaOh4+/vlaS
1UmDgmYNm3GA7j+Ts2LhpF97+SOQj3eN/MVBBmMiaecujIbjjtXBvkpC/G9D6i7aGFA3/remujna
s7/krbQvS5QpnrQCioW7CIgbkVb896W51h6gSbzX0UsiQDsSbKXNPltUowSQ88xVfXAgC9BvQLZg
m/MkccBEl+jVZCYynpeccu5bBs+knuklTAK9HTymdDCJw4YfxTLEvqvoCpeKsbR7yZHT6nlbi12y
n8eymGXMibkBltnom7Ce8TuCnbPvYTv5eKf4k7t2869naGrr1FhX9dXxQij2IUAr4+nJj/a2NsFY
QVId2hZqpWQERZ2AzHXmdrw5iZrpAg//ZUDaFhfqTwgjwhtZ/hVgbz85zxRZsqCmqVgXCecZbzHA
presGjceZ1edifgJ4fMveOgPEznHD+HmcK0JA+b1FaS1vbH2EgM3hOyaAj91NHpoOLw7l1hDdW2b
MkkrE1quil+pxv7mwFY9CeEadGr/VqSm1Qrw2xj7CszvadXbK5IU3DJet9hPRaT7WbIlwgnJ89JI
qxeFzoxEA7vH8F09GQ3w9tjRltAjnfmJJB0SzrvhGDUl1EQFBPilhMCd6hiRNRE9oTqop7L2431/
R4MMHJr2kXeQNRTunTC7hPPipQ0jQyiNgl54qK55HkmrNmHHNQrhlMXng4eFZg0fQ2z6d7gNeajv
rOH+bm+aULfGieT84UYI7uW37ikRyiobKyF2d7VfX9L+1vD0uN4a3lKB06XvjpEsEw5kBWT7NRyi
4GS3w0S3JnvNj42cc1uP8hOCjBwgaTvGDzbJPcuP6Ok/RVPQLyEUF3rZtizvPSmkzg2+bDScqgJ3
trvkLz16En7CMzwvxiHnL8DXcyj/dCF+Q8tDsPaqY60UjHolFhcYQWSj7PksOPaY6I1vSRKb3FNL
+4oehtNRJu1GxaEHq5EEQWGUZCss0cn4JBqclxRtCJUfjZgeJmYLl60yo0kIXSVOpu0vbHEnPPfB
xUHsiMxfo9jLC4a5mJ0ZHKFeEz4crUiCKm3dlUPCDnh4fNGt1PNXAsYiRl32BR5uwF3F6yk1PlV/
fRT/jtGX4636DQHfaPNPIY3/vqMa0dXGan6fkT/5E4BKalK5TMu7AibRLsMO88QNrKex4LLp7x32
0vjQ0OkCsZDuqQcBqweeP+GvMqFzlp/mm+l4mqDq1jJcOi3YAVwbHdGMzrl3WU9KFR4TZgsB0f/o
3ZKKHVq+PNsBKdbWAghwFnnRuy12duvgGixLGLNBFxGfx0D4AKeA9RbqwIsJd+Q9DjnFAPJVNt4E
FE7T45H6ada3B6UDbUXSVWqexpjv+su6FwFZLFYMCfoNXH/jsp5b09E6UJqRIIQajUR/ppup/nDW
D0NaUc1XtNRUVR0gSlsztaj3m5ncyKOvLOIX8o+D5sW9+CfkOp7YMH5hma8pYmsLmKLlXPZ15W/9
yk5sJ5+2wLYQLZgqRwGuLZnTZmaDErqqk2J7xw3I5CFQrfRt5TIva/BNKwVtzsAT1rraCk7BfHeJ
M9QVLyCvEdLkzLIA7fqHLVHuBe982soqLw7cvuh9XpakIGoncHR4Gq9/5ri+vWmFdwAq1y8C08TQ
bhwwSshE7n6v7R/xjHP1dlrXwRi2hSkW7fqVf5MgRbqTwRIADHsLqMc4RCgDG0q2+kEnHMqVL4to
DgY8bzuC1DVKYVC2pBFwB3ko96DjtA7eUKQZSj9q5Ep/OF4uT6owwjV/TMHF7OSHy90oDAthOKyy
kLJcwsdSQ5bjs8tZkCW72tuDrMXtRl1BXHviW5nGXhyLFKZs6XYjNC08O/LrtvPNTSiiDVIj6Tvc
XndJfisBP+emRZRA2UcAX3Hw9z296dfkxisGOYqGrsivSEKUuId5sCD4uqC+jWlNf0pWVfkLJcvJ
IR3JHO0IiFR9V8XINTRMOHj/7TfQTrk3tXj45vEyx6jqeWZqrZRo6naNt6T748lXGwjVOD3qfQt8
kRnvELEYCDWlkzAsy2egFh1jfW7NRGArJEjj77kf2kkknOUkDMs1oJdEmFhoFc+xLHrkoVWFcbT5
VbiqwmMCXWAmB/gioZXSl0s5MFcpkmu88nVMUqjhLIfnw0L1N00izjQBSScb0sKj8cMPtYFtng8v
IIwM2rHImLJYaK0JM9Iipaev0jG7CimTU2jmgPcNCsJQM9p2i9BwzJfTzMNhs+Hnm8pj6Em7+lF0
sFzfdc5i2ugPOlE89Rwicqf8GhxMdr/wPxWlWbjeK+V+aiDr9IwV+L805zy/uojTj/5kCkrbvJvR
oXEhC4XkCl/bIv8CWxcWx9AmTwOKWA8Dp/SA5jimGlJ8QroDby5i4/J1AlvCuPDfU7/MRe5Yv9LP
mWyI8VypJKcKkE7i4dXGkpwKcGaPReUvweZoHHU4aDYMYSRs5G6TE7q3ZqzmjDXfqvnomyH6qwTa
aNjImfyEVhO4Sj7By0Xkc5y1RQgoCem8kJxIHTuIZFJTNbT+1w9k+vp3FwiLcWoGF+agGF+BBzI5
413UY8PTVUz+cKwkNN89u+lgvLiVOVhAD5AMyevOEUSBUv0+EEzBpZCLIc1Kpt/XaWEL39v0t3rb
/Rd1v/GGDPt0FE9xKLEr6g2gC4u7Edpwqa/D4jxFGL2eGnWgUunvHJMmQ1bcGOWh9wwwkVUgvs66
/4eOvpDSBy28GnYG/83BFpsQ5qOd+t5a2dABGrUghX7z5IlMkrJEBC9Bp9av4rCXWHzNPrAYdQS9
++hRqOnXYXg7lpD9tvF80XmP/xh59mnY5Dv7HFg1+dJoSQ7Osda2mjYli0N9ro2Du9r9saFU3MVA
IHRkFQuQ+gI4Sq8ZpXC4ITSd8nsydpYOq+bfpqG3BCHUgp5cvqGl5GBmKue94GzcQyzl93N3/gov
TTKwF+tXt2JYBDkIZLfNo1BmWdL7AdtwqLKIhvsX/2X2kvnt7iMvutXkOoNH3yVNlghhgA1Z9bR4
zPiSzYkmtOGoAzoQNQfimWTeJNF0/QKQUFf1iDv/rUBPp2IBYlrOQLPqG3Hp98Hhc163BEfkU5Tz
WADs4TQ4DYl8HVT1+1+ng66thRbg+hBYje0HtjAehOTXC1o2O25Npz5tUF8v49tB33ivEmlHrZUm
S67pjemdeu/5YpW/anMw5Lbtx5j2h5FFmF71KV3nNODxeXf+yCH7O2/iK551/GytZvLogcFJFtAm
HuSXRdQj16eZ8nCU3rKxILIwauFJjllgTXkDh8eCn6eJSPWl9hDaAU+qByR+700fY8XEpkFikezj
rJ2yl7cnIkCL9gIlIUzrmuF4dIosSuKr5IWoxha4WMmS84p/vxNH/EGxdftuZtGu0uokMCWhhca7
HEs5wnU5IRfQ5V4buNy4l1bXwt61MHeod75OOye/VoA22usXsZlE8ddif+oOyhjZ7CcomPaYajRF
za/QXqd18tESzwtdhesvdTL6Pt/HUBqjY2vj85q9oJO72Y3lc1EOwzccDDGF8a8829T3yhcJDfPY
cMna09x/6vB6ZI6gZhv7lrBNzILW0eNHGIrIFBsYtnBHsTqhN6weUvGvQVvp+7I3y9ovxvdxZMuY
FTiDPP73WPup3N74Fop+SHQ8vI34M/+g5q2eOO+0ysR33vA8My3oclLIbza0Z9T43P5haJpos/2R
wdxa1pJf4cCN/x7VmgofbvpWpfnz8jnlYOpDQtxrCsfU3JM64xDxEm0Hx20aGAg7PTaCX3XCa4A6
hIiL3wjR50wN4dYN36OWpxftCyjxG0a5somcE5IUZ8GKN4f9ZcqZFSTLCuo86du3sbXszYP73uO+
IjnaQhjpMCy2mZv8Y/Aai33AKznjRjwG+uSCXJWpdq5CVgARXKHesrCMP4q9ukDJbiJQINXqn+J8
3JUUeZn1YHFJU2/I0WTYWOAMO29Dly9is9+mZx7jEgUAqDIZ7npB33N0+8n4FNZ81u/sClJuiGCc
xwe0ix1i5ZHs9oxQOu6kVqwRdnEj7kqR+XfJIw9AonN+aDEPyGWlSHq+bBRuA8nDJKaeyXi+une/
QsrSYnKRPaB57B+dWrMvdSNnzY0f35/lL1S5mObiWGyG+2UfZK6hues7VwiRM3tqvZTwt/hKMwjG
ISHwnmcUHqV/tbyFGrofNpOB77XH/Mf9jav0UklPiJoiUl0il4DyuOQeRXYMBwlbC/rbrfiHSRKk
3NDzKXbaXoSbrVx/xbY9KWhVkg8FxXpvK/tIPuR+dTom3xduTk1ccm2dDIXs5gNMtYvDnkNDNmRQ
rGFSs4RBUPYad1B6DbGN5oFDVlhqjZn8xfBDMlF64idCa2lamM3sa74ZThtbFDV2WyzFeY658lCO
CPqtWg5Lo4I6Zi9Ovo3YRcjKRbmbuMrLeljN1BzViVp1QE9Ce1ivneqlGxk8TGYTL0i+4Yrtgsup
sK3+Z4BAYlthu72keb5xLwlnUhXnCiIxFI3+z4ZjkUl/BdgmjzfUjQ/UAFT4TKX+yXlTozfmDvUY
/XakGEePYXV0bP/I9pecn+djw/HLlHcq95lzT+hW8KIIe16nl0qQAnKJjrDWOO8LDaacT/xi+pta
LQ3n74vM4kFdKYUHjTJ1jnIxZWEYY1eo59s3nNnZ5XMMJrVpx9q14RvPcPYHGuzQeRlGQE3hDlVk
VRYvVVhK0aG2aOKiNh7Wx7EI/Wt/DqdnwhxBElAnKB3EXiQ5OQjRWgnRygmwMnrA2DS0QG5YyPoZ
GTx8fB75t9ZBpfk+bbWoUCYBBclidNwqENO4ObmtjMDviZdn7Ci9YDt5I+SvYM45ujLKKGfGuJtd
jbmUXoUvg+sMlVw1YvRbKVkxq60cmwM/Hx9/Zpv69tjOVmFuMDJIM7p7plG8hWioeIEt8jFYoENZ
6HYDwQLrVSphcuSJcc0E+RjZxnhcsOONKzc40QmIccPP2/mmcc1SCS+a6P8V4vkQMLdbkVkRlYb5
3oFIs6qMyYK+uJoLqwuP3zhO9kb740empQXyoarMXPkS5nzRHlbBR2VoYit5AxDFtpOlOtMDxw/h
R3MXLRUnMOmckuo7O9Vs/yLS8KOyNTIaD49VWvhJDGMCbIoiqkkmaAtYArCoI373qWueHAKc1Fhd
ergRJt/wo2EmTiT4wPv9nnHrTfimK3ay8sQkc5+zYJNpxDttqEBZPbAwqpJVCtESRd59M4YNhY8a
o+ZdqBmXkt3mDPDW8cCJarykY00T47SOpMNEqnep34VkVfH9ZIzbA9EbK7CnGYM4nO79fnXDwkvZ
BD5ZXgo3vp7TSBup+Lc43K1nb7/1bcGmN8kHlwiN23DSy1YOowILQ+bEGn1u5zKQE/rtzL9TwN6l
1qhxk8WGbK0796M5mRHu4VG4x1cNKRiWXGT2csmdgBnmZrdLahEf1tfg8Ngtu/BYz7VAjaRJDP/1
SNLYy9iPHO0cMgXlKsdC6CvU0AsNSi5T5DmUKANp0xlxmRuTcJkG6OS90uZLJqpftr74zF4xPgLB
yQCM59B/k/f93cTTxlZEuvcu1i31CTlL+a1lDVEvwC27NMFnv5tWRbFxQI6V5QDWvdPbVCrzBYej
Py1RgxgLcDLzKneezt0rXlypF8SQyw9iQT9ri1NVfZHymwU/aR3piA6DbPSWIZdbVEEcXqkh0I5S
h0IfBMbpBqlkOrQpS1IIHlKlfRbP9Pij2QCGuyTuX9R3Pb8dOTHoUzgL1cN1+2JB16DYiF/eSIS9
Yqep405v4rpYKmKJUL1lPFv3MFCHvOxQXITWeAmyjaLBuQe+UyEXw2+Gj5G2iRCMrOJMZkeZjXLr
BYTfU87plJcIJB2aV9DGkSRGGkxzfOLwFs0C9Or41ZnMQ7ziz+sSy2ge3cBntbWVDxm8P9zZrgvs
/tAXo2WnqL3M5HuqBvTCPy9YGTtgLOxfW7lJNHSdNXPfmZtDjhtbu3L/6vGTNzBXZiQwjY0lRoV5
L8ZNp4daJj/OtobYWqibk6VG3j6Q7yt3D6HI9TDWmBYFT0Qp3vdaJmQv3DkZS2wRsEvy+ROtbDzm
+35//UVmoxw6H4yM7FEzbvOLxfKqCz1EEwmJKghta/QFWw1Whk9piDulyfmmeXEpuPaJ9YpEXUAc
vQzALlo78vnO2NdwYCTIKpx9vMJyPJxH6irKNGnQWOiiU/lzoNpWk1Y/WVYBIbTvRaL8o2F9x/vK
u8VvCliHoS6JusHkJP+RL+9iMXYxSvGzee0AtWTUrelArLe9wz74mzgJezgGvyuAaOqPFXObeTy+
G7Z11UpVq3OMIxJV1YdmD2Oz2Oz7Bnf3YqD3gpKu2Ef0qpzdr1Yd3q3P59eT4RwkSarvPNzcYiUg
gjI+O6GtEpDEobXokfrIwSleBchM8LM5YvJGir6m9USfqJOe0Z80t3idQWYFKAs6Ua5AG/fqrLH0
P00xe623xHCXE6RyAnlVZkxreBwHlI+iGQgfcWG/04Xb6B5SGVPOpmcA1oWcop9AIZq5MRF2gFga
/GkUST5l1SJVTlotXwFLssqBwdOWZAE+egc32B7hjIzqSDpK4EfV6uyw0NuFbWQ8t315H9BaJvja
nZ/LAjYBQYcTEK+fD0/YzQsmk9a9vRkrfOtux4AGI2QJ4jDfEVe9+Pap+skPIxrj3AgRwPxLRGmH
2utdafi2A6GSLpMV1HByiDbNstggWKK6ecPWeFr9nWAJ8V36W7S+/Jsy+qiE5E1voXC7Wi1bPgAQ
aC+IW/jtDB9TsxpZVzXWoguuAhJHSUV3OxazcFmygR6nhtcIhz0oPbH5OosVDqPHVUkicAH3rf8q
abfF1BFpmnrFE5wnLet5hYst/Aj8zYpZEIvwFX4aGcqHltMrzfXmxKVAUEtB2srfbtBtJU4LcpcL
oKohLxI6O3IEu+VP+zNEU/dZlXDPszGaYSPffAVpjbavAE0/Aj5Bb98bJZ4vJy15WMD20txsp2GQ
uHGxPTlcIfY2KRVtOX1PtLYVpZ1+AnrjwfSCWFvd2grT/Fl7aegTlC0/euaRZDHXNIxBqUqMhJ5O
QSFSfhCzCZ2qFBcfJxoE2SVP7y/0O03B92m2NSvzd84VeFiZjsZ2F/tz/+bPbjer6XyZhWzBhXHT
os1pArIwnvBJhh5sxfyXK+dXeIoqh1ls7hewOeZik66JSbMgIuevabdrGp65IXWyGFj2iZFiRS2u
et8Fksos5OywKt4MTzDu8RIl2x8k4+nNYwhmcAGx1vH9AMQe44IlQWFwQtoeSzFSy+5sDNP75Aq5
34gaPPbWtVlnOeRTzrJfZ8u0ZNO+AUU0ME9lvpugdWlv4h/pqRd3JlmCTzH+SEa2nxXTvfKl0Y2X
wsGff4VbGlnjrC9BSfpWuew9dXORp45Dt7+64aTgYuw2mPkwvv7ZtprcTDXaTLnYLUd/bc9BORAW
LLJfQUgUZi4gsvu2S7Cih3C4MdjTtHI1Mab49iXiQDGBuZixx7hzSJrDyDaGSBwRoco669UGOTP/
Vh9+pO2fd8socRWp2nLsZ4ghSSOTs+B7zMcZogLBltlnjfGPKSwt0UDO0OtDRPblOK6jmxOzv84E
35zjXtB3bbnKl6avcpMrSQT1jm72IMSBYyJumQr7Qt73Uy67V39+KB2blLICOu+sWR9xe60E2MkH
k6dUftl3A0RkvcGHC2sUsOZafY2Kl/FzNulNI5luIdLcekPyQ8/y6dstE65+JTA18/NXpGWmOvyv
NnGTA7zfmmk7l/kpRgIHrTzG/F7RIowrGt0rWvUPIuSzEa5mo3Lzb8hWq8YSIVZfhMQflPGV/myG
VBBobUf31ut53FsVFis2nh/gQawOekpxuYWIo7idvESyarSaMFirNu+vfPYav1iDVBwjPqScj2Cc
4Hvkt7Xl7gH9FFOrlOJgLfiFzo2QQ26jdV70WlDRrLEnr7MQ3BV393U1XilJMV1h3Jpo7kQ3MtVX
SPKBdccMe9dJJoQymiHgYwlp13nN4vp58k/ASMRgI3ndxR1T++J2+QlhDChU8XTSgFbbYs9+5iV+
lESOXq5ZZaTDeQLUCLhbrjdat/HWzbRbVYNH0zIodTOTpgyPceYxVSNjf9XHSXlNHrsXOgmb5B0U
+Z5S32NvkipCmqtz7uHMjkPQq5GodmnXTiWUydqByIdnz5icFDrIwmUISM9qqhpZizPZQU+DISiC
qplos6ykWY2BAidJ0HONRAmka6dQT1VPVuSGQYV91XN8V+Okqtzq+lRUR6VZqAZA0J/p39DDo2J+
bAQAMv2PAbHNMrPaSM8m0BZ3m6SgIp24DAzKS7DDE+EkaQt2TaYhs4c8dTswDqMPjolKqOfOrtJf
p3FFrUerjhNOQzoy1QZ+coeUt4xVH4mW9Tz89wyadszWNYJ2/nt/wQRaXj0TqQw5qCohpDRE9a/7
K4MktlC4bWto9dRXAtJf1sZ9ql4PBMwUnxOu7NaJNXTvkjQk6uh6yiimGUakG8ZltGavfJ/aRYPK
8vi5Iirj48LFHh7pO04COZFiZA4FhJ8yiMb7VXH79CVFzWov6tgV0oe4F82Sk8Q4KzfNLMeIukWV
zCVmyaiaHVr7uxGnZeBW8WneOCcqxthx0nQqVpaReeT8PQms6u1sAwvVarS6tb1/PNEv/8lv0Rh2
JZzBOnv1OBxaa8vr8I3YplJhaS7zJP54ipyV/eTIc3RH5FPO/kB1MN+dryz28IiTdK3lZ3+QHvif
5tEYIDQ/v/BJCS42YL4wM38DeZadBgqs/0OyaWkujKoyibQnG7468qFdaERRyrHtt1hCLSibgdex
mSB7qZy0pVGGUQnUUPdcFiPyL89+R7UV5XjwYm8Gw8fqtK0otmd4cUn6JRyQ6YIVxfuD7ocGG6iQ
T0Utvb1K8fJdjNyKeMdpE7G9/AnfbWEbAsx5jjIHMouVHNfLwvuzczRthvBPNvuJPsYo9f3ERq6O
hN598sQvZyM+A/iLP+A0rnPbd60kXebOD5uvya5GJFImQKrlvXxMztFIWE9I10Ax+ULBbg03A2Ax
I0/3E35UA7VKCwDsjqGVGzTWg0APX10lj+8NpOHrlgSB/f/X86PhEExTfvP2pLS0pQVvTNI9iGGf
+RbWNbDWIvCdIFdUu0MVif3a9Z6xkeftwPj2y7vq2iejUDFCJEKXT7hT9agzjpbV3d9iD3YEGoqD
5qvyavfyU8CpgfxPIsPDt6CC6zEm4VvYXzd+ozq67uvVZKBe/SWuZ/36w+hFUOhLDv4U8OaBhl8b
WgSclCRoDg8SxoZN2SD262fYmBDeiCIVozhXS6FU0YAwa5kjTY9NinYZr/8kuzVB+e4H/jUln/JK
U++Dj1LA8yyUy49/jy5MaXnuGeXIYm/BqauWWmMfUxSEjUz6y+xXqMidegjAfxthSWJllGXe4iqQ
BaZT2LNxUF9j7UShPFJEHkZCCKF74r0FNRca0UsBKJidPx+kl2BKzyG2XuQ74cUQoevrdju48F6y
ZwbOHikV1gqxwXaYEbC6qHx4u7vAQ7Vludu8cMeHO+0B5V7vNx5wQqFGg2fPcym9XGyPYBIDUVeS
anlcOJ3rTqN0NRa8BJMXVlEPWRWKjckR+cTL4BPtFITgGa7axsGyyDPaabHTEISHq46wUY9nojrb
OV2U4/aK85kAw9uBpQR7hanxWGZQ/ZCHLTKVkkGX6P4EZ28AfnEPGwV1MZdDuAhCY+XKflxDZjko
cvzdOjNM6lrerMrFOTLXr2/r1OYttyA0uUTse6u6EW0rZOaAJxN3EAuI50C35p2IGTRm5yWvp+6q
sjljfzTlvR0tQn8xoSouGFPdTjLxsG3BifInQ5ONvJks+uQ4Fc94u0uI+2S/EfHBUsoXipvvR67d
6ZcueL0IzlpIPH3s+EH+vnZvj5bPNO0QeGYXOPN1rCDPQDJpDP0wla4b6ED28ZQ0tCmx4wSvPfCq
jAibaERAnLxyxXR93MKNpl7yWB/tBIrPBiQapOqX1p7Qz7eE0zfxMFsHbIYDIMy7os8kwrLgYFar
Irpl7jit80Ux/Gw/n8pLOB1Q+a6N4d8idxK832S/lypI1iNKvB2r/772hWrzlY/W0vWoED1mZqHp
0v9/LCI7c/AAocUOwSrD4133W8rBAcE7sBVZDQ5yxqCrC0IsdzMbitBXQizd/caqwwYRaUBrqjgB
QRWEB4T3hviaKNnGYUqzYdtP4355DAM/yyNc8bXNn6f8sjuVpUal3hDJplyFYhO9NVA7BwcqmW+I
goYZC4ahWCh/4On5QgDgvzhO9EWO/Vxnn6H8lng+ywpZQHcO6HCqV0ok57RWHEsG1lyG/EZHzWO3
zTHLDUvSfNAvDvCO/mXbK5EFyPVp8xZ8M4nGCZHW/j5lqKT1UNtcg4RKD32WrI5ZV48E3tmmVMoZ
qm0MzI/UL9l9BG1OJxOhe13+eaIbVSYH6hqvap2sFGMpnAE8s9ngA/W4LESUzJJM+LE90Z5gdAUi
FvNZgBK6z0j9h7bSqdpoLsKNwDN4ZnMkcIuos0wJJ1iemY7T3S92wSuT2rWx31Gk41o9te1RfZWF
QO8PiJ+YWBJi8XiwF8Wlj/yB7HzOylutD4dlp7d33HN55p5QZfcMEuP9k/V9F55/4JnxE3t8SeeF
dwdHelMu9bJzxCR3zSl9dG4cLVjInkLQS+aIgHloydyBiUztHCsksyWuKqJmniZT8ILbCYPt0YpX
MLEKV8rUkG9X7JlRx/34E5lwha5j8+7l8UiahkgBNb/MaS6PZZmuDzoUNTF/wEFgAHlPxzEE5K02
i433aFMMOLlNtNuEUrBbsrIWl2Wx2wql5q9qGYzZ6WNRQOLeQxkOgLH5ZfZtpgztcAzWnYDsWzcz
6qzcxUI6zZHF7hZ5Zr40XJdcEnvUmpMAVli64KX6mopcMrLyDbdcrko62vxk5wM6LSzhvuUqZoUK
0hqeNyg5oXOQPh/z9Pwk66r9pgK2E32gukXplYbrOaYEOL++azIv8FXMHvAGrmqWDNwFgy/f8d/H
JOi9+xNrEw268UOPvQsxmvlgy0qB4mf3SijkPtN5VR95UjhEtaQh1KU7PHPML/csPslXDeErgBfR
U1uFWPN/5sffidarSFS0TipV6hOMU8arJQzopbKLT7V5FDGWX6USRcXYzsr2L5eLXn44fesSHw74
FdvLsS7TKKc69MU6UNYK59dJsbvD2ba0B3BTq7FjqZqsZuBE0KLiuLZ1OfgsN8xyoOqnYSriK9Pm
3TI/mK4RnvzdHEQPM6tgbWMX01qYLOfiR5iuLozfBu7tlQ4jFpZonbYEmTEdpm6rRnXzaeGEXLOP
xxS3aY1oPw+FNtMKFaSMCSqfdbmWmoAfRo/84TSmICwKOqfuPRyGrKHu4jK8GiG0WNpJ9yEOUeFs
IOBI0Hj58ODYNNG1ToYZYbQawdAKGv7MaTOGEVJyKLyl4YEzjE1KnRvJrBtc/PTCImaV8jQ18Bgy
AG+uiZww8kGnCjFMSlVaYSUNeVdmack2tVc9deaaUKNG/ttyoFltQZfixFET5v47qv0OwU21dug4
VSxjc4HqVsH9QO4NQm+BElnS3qVCSwYrPVyS590o75Q7MfWpMqbNh9EbCwIPtq2xbs6NSUCcY/iI
Rxe0JMWNGLe6cmHDtZUe69hSWAyZjHJ+QJ6RNewSEK1drLmuKR/cSWGIa334dqvcC2lg7O0jMXHY
lHKxsHnE7xWYIUYekVychdxZX/iCa4ef2oqI56p90wD537Y1QPbXzS5lBcnt8EJVF0Cu+SxaSTaL
0B7bw5X/KN8mExnTcfBQh3YDV5NXSq9zNNfyhjIGvHaKrIP4IOSJO6H6TyrMa6+20fcT4jgeichf
p1koodIWTdOqn+Rfp8Kpdqhp5WbwLceaemdMpJAIO5EyGCOcm77dA3r2kxejfeO4bMp2UInfALdv
hOu7LNhg18PTM3wVGdMy/SgjyBtklYkzCkz+UVUkUoWQ8Vu/yvspV/uDfT/ipXGOkHMxeLgTU8TR
eLu2/Qv8Oa1aniDiiSlZdXBMDXIEKIMQ2Rv1q0MUUsplz+LTvByvNeGVcFqtXyRjv3CseUlfSzLD
23rjo4xke5gEMa7BXnKK4+yzQ2zHyKoKY1Pa+bwzt1HwJidDPIn/19YEup/gObO/fQjdclsfxnro
Md9THOS/Kx81jS0dnsiT+FxOUETiefaHUt44H1lKBrRLuQFIp2rnXnty5p+cV7jqkUhxZmAq1Q8A
r+V/5ZNqUr8owNT0zYIuNmhnE/fTxAbrDVTqAjGSEy1T1KHkQwVWVEafbGM9rNbhwOgjnzl7MMA+
Yix2D7tTPlOUn2+OtRfHT/JHOKynNSQzTmpZcg5iy2y0ERYpgBAsRz0QWJCiHrahZNIUv8V3sGNK
hqimXni+wq6cNEBXpy5usDD2cHb9FFgd1vZ4H/arvutCL/opz+hr3rgOm8V0rvW23wkKMARp8Fk/
+IG6ZMmn1HcxCcA3GUIzMwQd0WyBzSd8BGjaXp0Qc+W6Ehjqdpd4fX2OaXgABfa+kd/XaXLnIKJz
XXQAtrULRmwTUZQ6JE73a9UE+/fhmUC1W3sCO5/cTr5rIXZnVGplfinvgyI/KXF1zKhol6z92urS
K2kRwYZqJju6m3F9k0xpX0xmm9HzLT4OfHBL1J1nSR/EtiL8tj/0ae9vxOhLej875vgNJQuQntIf
2KQ9OG3S3czhHlRcCpG6HEwYZm3SKUkVa2658GbrAZP5TYBJIR4h8D2EoWEbCHUyUbkt2j8w10++
cdrzJQSYkPcN6ty1BWnhW5p3hfGIMQMQe8aRn614Rbl4//pflecQB3mQNgseskTaOyogE0R8YGQ6
WNag7dDCv5imnvt3yr1pvIyfb9PkhMFu/pg5r2GOMAfEL025LLkh53Av19VCqJBZFgCe8KASfxvn
E3sfSbLthRSom26+wj6jpoP+4SLOhdvYv+/8RdyHBQ/PkUWyvAtnEvjiDFPWmGHUoXPVVELRBFok
STAcLSPM4/1HnNYwrX2DS4Pk5Pws5SK1+gMjdyH+6PqETmO35How6YRSf269tM7vOAsYOgJ10xwA
1IyLKxbJKUu+tBf3UG84VwPvqni0+hI/OL3NyxAZ5wn2D/7FwQLm/qBaxf8NNiuJEw5+mWIu+OJ8
noYO5+GoHHOCR7yaw4/KlpMHazs1ljHhcxnSA8pCSaHdXzQFVU4vLKaRwd8tELLdHciZ4osU+xYu
l8pkLDZepEECcQCGvouqymcEXMzKe+McT2UFT0XEJOY4TI2Xa83AHq5H9yDZlv7pZmSrIT0LJY8W
cF59d5fY+1DMQ5rbHwHwEz3eRyCs8n8YCKRPAUo/f09i/ar7RE4s5UOfjKp9DoUsNu5fX/EBRX26
pN/++Fkui6BThBni7PD/R3X/MvNj4LTkgXF+DLonWwHQaPym/juSR71MRJAHspCums5MbOyZvzUh
VgaLKFTGgSFNqP8SvHBmo2dP2dKHJGoV15cfqmu8wfJv4fulnijtv6y/OHKF60+Nvi4jh7AQ0cH0
IRB1BezxUG77aIrYj9Mgtb5l4G2c+sDNMWCpL6PDP2s4Y76Zjnx0dBlDcub1/uxJcIMmOokfuSSG
JJBTbx2tuEia2i6JLp0+2pY05ZpZumwtV4zj+sNQDbkTFL7rO2BdTx7m/sRHm44mkFIwM1x2CIXr
vNxga5xbrVhod4CEC3XWmKnwOyhpcUsa8Ge+3dwYE8WUwSN/POtLWkELoPDRM3q7+eSkhboUYP41
broCRDjgyVwr1RR3Zdl66uuZKbzkrX8HbJ5A1aAS28u0pmeqtNo96fZZWYshNItZP8UY3Fv/YdDf
THMYU7u37+aLVef29UaO2/WhG3uS71Dq/N4V/If5gdTeHiLxpPyJr0WP+GojGkRoRqvBZeFZB84z
Ti2j0DHl6OaaaPZE8BJaRWMKAcnZbf/UPgp/FYOtFqSFqLeMbDQUpVn/e1enPs5dM4nG92fxVpQ4
x6jXQMFVr6c49+0OvIv+JtV366vizuApBx+tm2n7KccgqJ5LnVmEo6NngkwJEjwyzBeMAij7P9rk
kNHw/Tf+V+4gciZMgV6zqZd58c/fUTGcwDQ/KsliQaobu4wOI7WGmiQCZV0vTpbex8zqJs/phQUR
ylXRVY9Dvia+ilIa7YskeNPf2d/kV7ZAqo4nA9/xwxC85Jb8k+qHeEHmDHiQn0cfXRGAWG2EeBWO
dUZdDfLL3DWDjv2/DhnZx5CnIvRwxDi4xZZU7jC7zqyPhUj09f+3gf7Gx/DSVt7nNADkPNm7Y3Wv
hKS1X8tx0QBY7GOQvpqGdWo1gYFmVN/2O08NzFZ1CLIadFLuG25tKSvZ9NNlHQT8XBva1beGPYhc
P89XBwlwQ2uBo+uKqUxcaiGrU3X8ORwCZKVed2ymJUMQt2Wm2dXzJNdgXgm7tk2MgXrxACD467OC
eRXZsU/MHv35U8XYiBP7mYUs+dJp2/px0FX6gyL3qf/12p7ki+wKmdNCXERNqgUZFeWUXPQbXdY+
Pbk+BDOJeJcslWAp8usj8iDSg8v6OowGdkOdRW0wPucuGMh+rdm0YVIoyOY2by2lqNH9PqGZAwlP
XNAdUGzWVWBTSu2eqVYgIp86DVwGUc53pNorw7OSlhveiDZV1ILWSHJDy+OqCrPjJysBlgll6NSR
ynVQUw0pMt0/8M+fSEG25vRShpXXkvseJcXuGsLvNCPXIECIk6WM4WNqQegJnhbqrarQWwL6+CuQ
7ySJ8ih5J2+3wPOo915Lx6Abbu6rRS/1ajQpCz85fKwFNh6unQDydk7+z/bokqsuN6RF8hwXInr6
obmfWhzXGbXmXHLb0Lia0MirkFvSsi/CkO/K1Wr93b5E+cb5Y2OKnmOAWaYMnkVfNt+0ePx5VatN
NDtl6zjstk5bzX1Vn6OKc66SPoBcrhNQr1DomgUjycfo5aul2B2W280ggcGzOhufhPD2HKYnYc4b
EbSCVpJ+IbvlulV5XjeL8sFw1p+3fmDRRT1JtM382uyzl8IQzQ2nDjOGfjwpTzms1Deu1zbwfRKe
dMBQCRUpeuolgncF5/WAlQ47X3OQg1WGjvW/5so=
`protect end_protected

