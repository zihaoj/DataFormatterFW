

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
W4ihmw0SHnxv/qHHP3XYWn5pGrBTr2Gt7T1nGzkJJ0fG0ZuPsJtJybNxJCVDjkEPLSVgdzCDp2gU
yg7BKAMBLQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JdVQn5lf4JOc5cLE9Wv8cqeyc7U6QeYKIT8u+5QRFGxMwMEJF+leRExvYVBT/b6sIPhUUwZG4/PV
6OnRdSEaVLEoSirhYpbF6JMTVrwI0HVRLHo4X+ViP0ROJGUQKiY8RuwDzd9rZnbvCXr86URbrPvk
A6KtSj0hSochpQuJRhE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Y/3GHfod0E9RgmwTa647zpY5r3YC3zG+53j7cbOPKgGh4vTmbneSK2AzD4JNKtdHM6/8hbdr5dF8
Cn1BaGa5lSzDAxLscVzn9IpfxLWMUugzQR9GEaCyX1vhgw/+XnRwJ/a0y4S4kHbcq2UxdqnHNQfD
W+FQmA+g+9ik4w3sk/mEOr3QCeH38vz0mZTdFTDzXzr/Z0d7bOf7t2FV8CsE+cfLBVngjRXOj8Ww
+1OrYsJZ/o08DvTPVCRZlTUv+IbXQFvCQtx66qZHWiKgiQ2eOLOw3cnKtNsXeHo38hYwd0jS0IW7
UqmjjNWSQXZC3uU4Brj/c4iU58WSdTq+R8hCDQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2Nu0IXsHL7gf9cvUYbq5riKYRQEVc3ar2+yZHz5VU3jkzPNl6VLkVsGTnELPU8FGlXAzTWjnKZaa
PNtFOJhSbdt+BHE6atiYqEcqbBgA0ihbGIq9SxmZpPhvTKQNT6G/S7JvlCJqHMl6Ky9VhO0bx5t/
etlqyXhu0WBbwfliCWw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Uq2lcX7kRmke+UnutEu5TR3MKKYCsYq4iVNl8UyJQX938u6lUTljAFAMc+K2EzSd+AyTFcVfyeI1
fCm45tj9phc1JsNaGj84/Tr6qSWsEKyX/6fRlRyGdQMkNNtJ7KhmYGiPUHEWkFTQdDEzLRJOnJyK
S37a5WCt/VoCJrYxJEiMg0QgB0MBBGwOnQfs460EdGoLvU3TCSFlx+JMpv8SGN8YjnlxFLsnsCFX
8nwyZDgwTrMbxGjxoFerog0Vt1UATQ+EB3lQ/kUr12fZqUOc/rNDlOfYbiZmb8zi/XQAPUAfIiq8
OLpBbmsqAYQflSIFfjUJ8uy1v3Ll0UM+4Ck5bg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10272)
`protect data_block
MzF4BOQto+EO6qWmbYEH7KWT/rxfKDcCT/pZr5Q9a+X/nKqisMnDD5JL7sHS4Fu1Ku9thRipeBqY
ayhTbSt1b1tGau54p0y4X0ojgOZAOztothAq4fskItOqOthEROX+fWGTLGoHlWdaW6DnEub6RuHo
uEkmG7nbE8k/HAUasfCIYWwDyaERjPRz2mMF/DDV9/R6mHKA1zTFEXI4kfniAfM6rv07y9WQHjjP
jBfVaXyB9hLYHjs0pCb8jNsJKaHqCVt0X+Rnh8FhDq4EFOMGsVJHBNJXiXTbxcT057qmzVuiJpF7
Ru6jLtybWuGuLvXcVMdkQv72HqboDr0FnDfs8GyP79ChuU+qNm4L/aZht+U8mTe4u13Uj13GpUNZ
uRDFa9RiGVwg9ra7f0hL3hdPgD2H5qKMKRL2RQb7G39jquOAj4/bsBf1DqSSjuRQOB/29dDNS9Sy
G0HCKjGjMasTTYFgN1DMGwrlaES7EL8gDf/hQjq5yaNsdZGH74+XNWFCGezt3i1Q4VXsdkvsPIks
8a1yEPM1/8Z2jIfOux5qVCPIMQbpL0jkPx78V9jVOc5PF/d/rQz7os2dSCmhvApmnsTn6vjsxnbJ
kYS1ExooTwWt2N/ZV4gq93Bmm9uvWW1z8BkDvorwpCyzNqZ2XwjiSj9ZYBXwU9AcQZviPbGDRFXn
ufmQqeIiyUoYDoZ2+MVTW64bFhZiUBidBokpeYc+crYnVTsuRCzOsfUYS0mawwxWWETJqbRds+OH
BD8t/cJ9/qHB+Avm1l+1hayvFajtFX0fPxKTMCu1W5nvQZsRnlGEDs31JzWScaeyVsah4OEGIuB2
z0Jl/0Z6KPYWBMO9fBzjHYISUZfhxa+Mzd2SsWGm0gSxfETEWfyQazhfleKuqFkTpf0vyV0gX0PT
iIV2LAeLXzo+ddbO2DKTI1Q7NQr8g3Z9XWBYurxwqdyIIwUO1wdjHhyhaLB8US36KjZcSBo4O8O7
pDgS5qed6dAOpd+iAFunw7E8L6TNKqkHNBnupA3GgRI9cyYOgsxSbpoKJlPfhcVYrnd/FSPJGrKz
PHo+WhcHFZhsGJSSbClbxzlDfNdksBae1utJSg5Qc3rUc7EG/OHRw7HK/XHh2xE62FQRdVkfb2Is
XF5LGVlYiSFEgc4luY8NPH+36PPZgFV8iPxhAfQ1PdpZlkcEULQnDMdax5mfNWPLkD8EwVHV3MTn
1AkKvC3zD0g9y6SoLJO7d/O/WK7FWzcj6Y+BIB3SeHjzJ0XUq4ZSt4iCee9l0EhxtYO71t7SRA+l
fqotjMRju/06lrEQi1rwk0whJVl9DHKiU4QWrX6zWAD/ilF69kUXmIPM/W6NX16sn5wlL6hiFPdE
C4qlpmCTcu5XSzNYV2+cs5olxLZXLY1GymS44yKpLVFu5ljX5qB16Vbj5wvp622lnPvzhECWoXXA
Xy+f0iBl5kuErXOUKu8EcbUQH2fma2o7fOyVWVxU33rCHkfIiypHSdzg/NRrFtWrLu79qFChFl97
fna147E6A4RZRl6np1j6R7o2/L7POFyiQZMTZFhkQk1+CJLXr6GH7ERggsvtlj2saXVn5QkdLa16
sDhCw9aM+1E99WTyfHTS3XWWoXLFOVYvUQfsBuOgM1eXXf6FetCkdAal18/Tghyzkz4jpRhu1onP
deSuRKQSYACP2XGYYYRAOWJaeSRNz+3cYdL2gmXi3ioNw6dI4RlB346hCXnYBdlgadcLgobXmUPa
cEIFqJA/mCq4OVJzB6wu4Mid+1B90jk//Yvpw1BfLWTo6hI2UR0MRHu+svaSp3C40Bp/LbmETH2Q
fp44SbgWZwF2C4pPMsKYEOKFnIbCLMIdwVlb71RS3xU02FuaIxq+cJ2/LRwFyKSLdntRbBES4CEl
kYDNclvtCL9Y061J4mfioXNij2mmAlQenVJeInZUfHsOByp0amV9Qty1KKdLwiIHHInrsGD2JHdN
AhZZgceic4U5KYbUVCBCzl2e3gR2l/ilM4vvsPaSX4u7rM8r6nYFPc9sFFaqEvbb++ohywiKr9+i
uxAMjXa6jYHHlg/ZsRcsny5+y6o96Z7yOPRhRgrgWbbvDG8M0gf2JpE1II41IB8BHUjDM8WMDgDo
Ltz31JjofRndEaFGIckU9deSqwYD1YrCvF/1O3rPK+ae+NIFT4glH9KrFjx1k5knctYo7ctqb7sm
JQyCPejejMme/v8ER9E8nTENqBe5PFTTNA41Jd5JGaIwUeFKG6ZYsKwh0PhvAhkoludl52eKO3e+
5bcitsdi74dPJM8xnSvqxHA7E54auUfH1P9CmMCFtMmi0mLDa4IkPgoKVJvbABfBAbOEqjOV2Ku0
+MJr0Lka+Sl51UZgz1tLT2Bwceeb5UNprgaVPSRrOqcZ8fW9zHD3gEbD4SjwnvuFDij3haqsL/B5
wMimQPGOr4gGlxxxhvuMsAKopVvHziymnjK6+tee6I5v+E1pNS5Ozoo/wQOXIUySLpyccJKYcqVw
hFAhOSmFaoy3wccqbJFe0rdVHJBn75HkVatTcfFP7gq3pRZugkkJ/RZmEYrnmqeYHuqQjBfawqwU
C/QMAXd9ZFnbKdU/zFLjdS2GheJkw6aUCU2pMGIyHqAF+A6T9eIjdF6rt50N0WPLCz0jN5JISFQz
JoJZ7aUkk31Kzlu1zYYq9oqoCdAj2w8yOeDGVEKW311ANBTkL3ZLs7UNVaJQby7F523VmoNkVBee
MtyHDNDBwBcAfhkfD5vHHe0TOPyGovQ5euHlT09mQl0jIWj+EorSk3gAShtat+qui7NEX1oovcCm
Id8JG/JKLdTPIuPUCL02WDqXlDKGnoAGpaEYixedl4K2+xjjBs8BbwIR0h+ioUsxOQuBL1mZwRrX
n6p1KC2OY8XVANTIY+KpfpxDhDxdfYc4+0I/lqGlHg4TVvg1YzNwr8nTqnkTxU8rm4v/2mycQLsP
MlUVkrGguhX4MYYcrtdGeznbbU0x+s8NocSjKf62jCeas4lwUlRhk60x3R2y6bhcFu8NfYBjVtu+
JacwrN+seJVzXoT6fBSGcHXvMpoT1Z008y2G1BwhaI2XhVjYKP93SPcMaIKtxA/rfauhVE6+SCoX
Gy/2X1F6LQJEghsOVygMgHhCo/thgjdApO7oVI/PRZLy8acKxUA+/y7NOfqSDnb4QzhmuZLJHmBP
WEIUUqi6B3XpOBzIG/3PJ4/17G3qYdrEuJc+XKoQOiNsBBBoG3C6kRSSOl39SAxRbbPVKBH1vD/y
PE0v5xIBH3bBafxWbIjsaF/KiAej16OlA4FRBY9nCtbS461Badzm6Gsf52fBpVy0Sa3l/pIXKExS
GTliNPwGU/Y7T9mZoRgpvzSl7M6yDnFTPCJ5fP/5XjmKZIUcMX6deSsLBQsUigAjX5kyaUR7HQX2
ROK5rvcwJdDL94XTfwUR0TdAOOF4VSp9FDxnGD2j/uYy0QJjAF/pziVt/YTt8UacMxhYIA5x9fUA
1762xQ66qzl+gvGe/8SUiBhFV2a57w69eXNBmL2eyAAaEJnfyCgIB42u+LNxRexLYJternQoM9K5
UCyNgk/cUFoR6iD1sswLM8a6CejQjRDTgTMnxx4NnXwegF44vwJykFO19k0slidj5F/bhaJ7u0DI
oK6qFLv438ZDuYXc+hqMKmayCviTJiRawBW16JZSMOngHmfwqS6FTkafIPX0SSi9HzsBxeOfJKLl
Dr/4NlHT01WON9GI7ZjZqIgViDDCnNNdQwDLlAESLrczARSMbT9F6Idl6VaDLoCXXrDlZ1WtRrg1
WdjJtvCdCA9oo9NHr1WOVfLa8T61IHhdOxDsXQEbmxJ4j0zmMDgR0OWTQpaOEicQIug52IyaSU8v
G9hKCR6b8xG1/bAi43eRid38762ZJVu699FwqgfsKAyftHbygl0jSXMP63PpIv6jMmxCn4uAr815
213sRAhfCYn57Phs8kB5A9Stx8Oi4Gz9KyXWcgBbUuYIUydMI/Dn0Lu7IwJEgXj6kRirWnUp6+8K
eB8O82/txzrm19GD2K30vjPTfF6kAv/4UWeza2qPnQaCEi73EwauLbz0ObUo2cHEdu1u9obgZvmd
xRj4ArVDVx62GlQv6DcJYdNwmcAun+A/06zRxXzKLbFuz8T6gZ3Mduor5LZFG3JOpdk2f+SgHTvE
Vz7hqHX3KO3Vbm94LfGmSLX6OX8ZBVt2UvrNeT7gVGSmGV6+HrwHGJNoJzn9CMNd4zmaycKI9gfI
oqjYwKuQ0H6ZVKj7HsENbyOSXDGn2vh3/5as9iN01TC4FswSuFEi06P5g3cnP3UXS8w57m1rz2K2
YZNxuwK7bWkxd6j0MHB2KqbRvwA8oACwVuQFiaIn5X7THqpBaHVIMAk6AnHHLk7h0C44azmzNZ/n
ZLyaqbwK8dS8X1mSd0N6PWGtjJEAkDnTUAuSXuHZ5C1mkHo1enZ1c5V93up0YV1m1HYwxLOgjTJP
3ZgKaxuLqbbznhUhe7P7cVg/6LthJ446noIMt+X9/tfevD1guwBS3COqQh/apajMuMblqckWT0m+
XMit5Lzik5slDJlBgVERUz4xTeprVM9pF/7G7v2azqNTGWS05GuZdXPeAYD0VFJlwzBMsBVp87FY
UR4xMoZBzuPbubn8AF5a7gM3MrzfuDUvITELnJ4QV7cx2Xxxp2vCj3imVfWeIoDA+qb+gqcHSTe5
Wq/uDDyulvh1iCXFGv+cCeWbYN/oidtuYyBNqR/nx7ZKN/R9nCWC9hw1GVSUeuIcvyEYxpDWCNsg
Dux5EISDPJWOnOFtmlz1hkDjUaaUpFtZFJt7pYdreZxRyL51U9MD8hzgHM/iLjZ169f4d1Xzgr17
AGP7eZtL0gBeolx8U+Ikg9UFB3zQkXzndgJ4xiiXeojHhn98x/qBSxqQ7IKe/wiCLawWXw280iiF
JWfTHNrYs3/MxIIWRwIJLiqquekW3wZl+unidpOmRpkTJvDh8KVdXEwsiqm1qQ0F60LU7Fw/t3Z/
7HpjpCd7EmbiWghwQ2XeQ1K//0VTr4B3elwdhAEW4Ewx0E0Rt/SxUj1D9Oa6se12gq3E0kOHgW90
TbdZ1mLRi1LPHgSk9iUZZnTupe9v7t4oHuE2+hisOI1fiZJ25hsK6obgTi0VHm7yMCDIXJwGN27q
c80hbipyrnafzZm1EQX7wmaGuzQKh4g6iiuv2LHfkCrDVizXPF98VkUTp5nHbwISvnLXG2zxDNag
PlEErDwbrElLFvFQg0J6fgbLwHS62ECMGjyjPceTBX7pghw9yL0AUkMlSMaTmQon7wEKAVlDLPtB
lT3Ff25FJP2roVnvhQk3s12kg+uiqIDWZnzQMDAPVPU4TiEEDLPPeLM3gA9Yo9R7O1qfwrrkexfK
bgU2DZqPmHAEQbgtstZdvO7s0F65gy3s/POElZpxN4svj/indlkykclUGQIDtwAAc8jrmgIpkM05
seldGdfNE9SAedmSGmhfXoC5vRWDDGKcW7pA9WUiU2OSYaE7vTHPHe877Zsp8lb/qSYW1XoTYYUZ
AawRQhCHQp1f4qXBhpAUNjQh0O1GEJdewu9FZcuPEThNHtYbfcv13plVW8EpdRQ5UkCKG3nUQEyl
cq8pF4mjUHbh+8oLp8xAs955mzs3INJbYCSoJdnKnwgbZo584e+nFNU25E6vWuuedbzVxxyuz3p3
HQ6x3W9H8uWlfqiLcKXIpTlB2oorO9oC4FjxjOx2DoOy3lHa5msxxD1RzbhNkX/KfyKtWsUgTyto
kbmdhaqC0K2FOsSanvbpkqTYROcAX/AanAkyNlzrD0XRrWBRyoXwHfidfH3Yu7DDuWoG46hPV6Ry
8VXgZJrGLjDOOTssYb00uvI5UX6FqOdbXl9wOwBghQYNRtK0r7H2xmWnaKop2uF4go8+me/fqn6t
LD7cF9UJ5/2zcfp0DKlFnHf/fBvDLbik9zcHks28DZN0UNxRfuL0hCaMf4PI1XWfumd5G3Pjg8b6
s1j8NOE53ygsHMBIMbjARNg/5dbfD1LIQe6hZH1/GMiUJRYrv00bkCCC2hQJxhQzpxzLzyHzXnkc
+NFZV3oIz0VrOUWOwaswObE/+oFxUIcvlv1NKQ/8GTvV3fNLOxKVuZBKzQNmeTbpXyLVF5heMgbK
jIGZpy7uzE9oM1MMYB9f+57ObVRxgS0tsA3illBXTd4mUjAR1pMjYzVhWEIuPdJzv7FzqRKXglpM
V3lJhq/QZNjp+H9Zwc0B2O67hCXsHNSzo54AsyvM8ZS0PS9yJy834TiNAcn6+5bhYVdm+E5yrtXv
7GB71kyJxD6AOgjUV2DjbP9N6BQl1EWlVULqEfF1n4HETFGTnpJOP/K2VD3LTN68fBndM6+3kBKT
ArdpanvLMmxNvtwex7MRjx1ko9e77iHMFGXG7xu1k5kSxvcEiYNJgmqxeJEjcCrGsGIAKHbjL8zU
bc/1VwOEw4FsPhlyd4fapYxRGGskuMOjYXorIa/UedHpd5qjjdpy1ddSrwB+1JR1/peJJjxVq5as
PGRXaclEQ392wqE0VnUUDTLdEJPrinHhzAMKMqZ2GUhiGIwIPLUVzmzCr9sKtK9N4md/9miSXDsU
l7twx0FNz8+v+8lU0+C4I9Th3o40aMeBLyuwu0O+Kc34MUmbrnACwbPZcZ7JhVBZUH/f2VrwUyDB
KDRfsRXQTB9yrBQTbRGIRp9sShkQHm/ebzv9+jxuwAJ90/rykhBh5mnpDUqqIdDedC3BTi4HqMiJ
4LlY7ojz46Egw2mM0FPJbxnmzNmR6AMnqnZhCZzrPxsHtKW0JX0K9DKE6WhrcFt8udZ299ycMOGz
vHNnOo2O3hAQR+CFVQChxV2TjZ/Q2byhZE/z1EP5weY8sSZ5Res8Aa172rRIbfxgw1WeVLzlsV02
AyBQ2ut3S0YEUR+PtgYP3OOqr7w3EN3x4IJNIw88wVa6swVH7Xpj0BECN1dTZ1Z39OWJ4P2kYyN2
PikD2aP+JBWbk8RCCUY6sc8RXp1l/WXXgIp999RFKv13H3q3SIPcd3qfs/A0f0GnqPMS1uZBKkFZ
QM4MRjfxUzVVGfHDQbOPT4pUNlQWe3x+1oQHjbOmrhIZkbbB5vgdUBdM1phEJ9mVHf5511okkhL8
d2v2hxy90fSosroR23XSv12tgsU100AxOud5pcMiyl7i/CPIVaxubBW4fp+Uaj2Rn9pkFcBnGOUU
2Xfjz2mHP+lLocbZCzxwWkZEQZiKF/XgMMpR9B2SYws11APf/fBqdvDpxK3ZkLXqZHXveZA69foW
n7If6H5D8JyqgAq4mm6ywlqLwJlUlIInTRhWw/AbQN+lvwnMvubVl2nqNFU8p7eF0XVIWh0ORlYp
Rt0GX3hwpBhIwrGvH4GZvIKgKTFZ/CbQIMcLVsuGM0lyN/mGgqasxyk2eOm+DyVmk3Tp9twvYQPA
5YNRLlwX16UHhZWJXJZQj6mrl7FSXwO/m1MPhxjBfapkW+pRyUe4bMZqW/D7O2wYjuVW4jslsh3J
vSLErBBwcadgdw0QTYOkEDkEUqvg7zrS9AKY+uPtpsccL+XtS5S95jFJQOs6Xdq98H2c6d5oatXD
8XxJ+AYSAoNPCFAY/5qI32BqgTqxl/Lrd5S93Fg2jY43e02Y6tV6JSmR5iwBZqod03wWmW3Oc4wf
kmk9Zlu0qZ1I0x+8EHKlWB1cS+Nxfo9nyVesi4XMbXESUGRg+5lB6325pXUMIKIBwLKgBa22CZX6
HxDms3IJOX5CaW1o/jFFcciHkAoJhhQEs3ccEEfVampgyxV4tLKd+gaYxkqkGJt5xG9ZGMyd5hE0
feGNBdm2fRYIiApk891q66CAC7Cy9IUbs3tlyd35MeCLNdVwYfOKRtTyHozYm+xj7W9jkVleaYbp
/DlysN+ZEAuH3U5hT4iB+KlPAi3ietmIt8lfVbip5NJmRGklm3vsWuML06Q9UHHpKezQdmye2XO7
uU+UeEeUgb2fA9o/DU0rv1XBbpuUMC8H1hkmq7tzE3h/RjQOwCZ+Fw0UQcabUNdJKOKwh02hdpLO
eoTKJqsimEf5iONDIIwH/CAFQlXEpn3AqQYSuLXe/XkaqMyxX28a3b69AmuyJDBDUEyAWEAx5OTx
kxMakAzo8n+yBAY67GjYdnPMSLb+BGc049NPR/UfZiEMz/9vzKm7IIJZTF6UoAM7vRhlKlLSDgIQ
A8q70H48DoBRv5wQcgd0dQrnREFs3KlwGkXJxDG/+UdfzTNmAMkwcr8XkxbIJyvoj28Klrn6GrES
2DovaxxEFUWOKcWdt78iqt9Y9Moj1XstOUkQFe7xCCdta8XCnILMDwl5Wukay4K7VN15xy0vgcA4
M97PVnQE2eQP7JLfLk0q/l2Bv5TJoVlN14IWKHmYbC73v8LwumJiNk1CwAagvPDRnTXI0+pLCk1T
iWp+l30Ym5DodH048PEbz4gciMWs1JxjsJKMqJvNk1C3OeV1SENubIRVlQQ7mspxCLFA2MYmYEid
CyKXx71tRx9YPCrHt69B0wwNAIVIPCDyFLTIQrPQEXv8zfSRr5ChHReatBPbWNpgckcbXgccPOAF
6VPszSCI3mWQ6gQm7wXyjG9fX3bSCg072lJU9eA+L/P0aVr/2Q76AdMog2/FNTS8NG4vRtpi6N5/
rLjl8322WNZKWMZdvg3u1PnfnTEz3+LkYqHvb5fWijSiU39Yn6hLrWj3GNRZiVaZP6S/zwP/nzKQ
+XxMvxCOP3b0kzEBQJVk+/WmUX0RjLG8NE2BmI5LU+snvSRq0K0K/ldZHWVfV6Ux6pD6JHiyh8d2
f7pIYyKrr+hv+E9hdEWG42CoLbXAfvLmKgNgP2Xrw8cex+WwT38ZMCtKr0J6V/jz5k3sYvr6kyoj
qbDFYCBys4+R/QFZngBPODKCMJiB+fXOkQtuTKuUT78cQg/PhT+oA4+ttIRG5TmNjU0J4DUponQv
hfu+u68p2365f1zZzBJM6ezcU/6qmMbL1aB8lLao4Ehd6cqinESyIkOuDMoVPW/jkxNU+HU/Iyjy
ZZe7J0XBj/0fLXaEEvTReY6M7LqLMLP7+6IFNIC5cIeDE9066C60QGyVlQzbMdFbc5V5cxIdcJZI
xcJ4EConiWP7taWKUDFE/mUQM6vDGij9FvbGJOLDVS+rJN714sZB7CWqy2xhVUgGVQAkpFGX/NtG
ElWYaSW3Sts0Rm8lCRoOsJu1qMkntERjccef8qluV54DjtsZUrj9ZGmPpcm3eeWh60jYi2VvbmTW
SgC+qdas+vWiHA2wvTLWkZdQ3FNL04lfq3+YKct4QsIV8eJ9/UGHtK8IcF4fAZQZ5cLCp3pi7vRF
TUDYiAtPKK9YrNmHaAH0PWFmnUntEixvwD/kncsqyii3pIh6Z6XTkkbuNXcyRhD4f8D9ImKnkD2w
Dpz3xtPlfgbOK6Egpevs24U6DQDApPiC7xNaFhnyROSpU7VfySLm4sIOQBajPS5iluPkbnlaTcAE
ZW9kEw7/qecvp7QRrTJpEDDMUYGHJ7lJxOq61T3XTpSjb6dt3E/wU/ZuMXEovbDhdbyhhHKghOmn
s7lXZDqC+K2d8nj3fsSMTh/brgNoDaO9eWFWCWwtOa7/wwRQhFytH1V0taIsIeaJ1Uf/yZBzMKnX
gfau2PWtZ2DIyd877hNz/rYODKI39P5jns2Lfbf8GFvM4iCoP0vBjWFzPP3Qi8hhBuiYOz2NoB+l
v5CkhQ2lIltg3G9ic6w5IIgm+k2sJ+ZIFvmyNhaNkdvzfG9ILdkU49BgzQ2BiQX11PMm0Tm7Gecc
WNw7Z5eiMJqxmUKvxJVC8Y5y2tX3vVK+QLBpZp5hPAiEg6fJsx9fyv3IeksXcMDN9GpDSaJc7C6a
NPBsA4IyyrTa546bpjDoz9Sdi1bx76kEuWUyggkfl3neNumfw3XlqZ3SPFU4p9mcpnioslyEWUrF
nsj9rxPKA/oBd4G1fjLO5SxDmu5BgV7wPuXvVBpWSDQu0P5kBaBDbNuSUXg3F9XdFxmvFRA+Z+0a
QUvI8h+MGaBI78e3WpjMifIRt3K50PkE2DOUz65s5gAyJni6IXcSIgs8KneQHtAlI9MPELQz9wCx
FLv2n9INm6i4cci2suz7LBOk2gSnyCjr9ugYwK+rww+9rB0n0mwB5Bg1CZ8NwEth06LpfEvR5gBM
4/8FTcnn0RwWaah0BhFVGjCif5Zgh1sdJh6AD7zeCnXsXZbUjFsYtiL7kDeatgpzd3W8ygTUgp6E
r5t2e8puRGseFhNA8K08vDykVUQBggoCrCGjhoChkAez0zxu/Y5tx/vzPIqf7gqGERv0pdXCwgOd
T1gN5aA8gVHpVgrNd8olQzpErzvNPh0mTfJNcQ/KeJSCKG9eBpPk8f2JH8Xxc6CI6b9usb0DXzq/
wPe9HKTGgpX2oK+NGwTwa/B4ZAb0Xe5sW9x5veRbQLs5cCcrikJUxZ8u9e38SWQoBLUJ8sWpHFkt
R8j8tllyEWTGYwf4bjdYwTteHfUd7+yYCErclVqeAYQrCpsw8fapK/y7POT7jZUF5Zcq41wSUgfu
/5qMcqmz0caAxhGOstYZaORgWo9X76QUPPzoZ11s508ki4datdtnuKPBNdF3KQE5uQrc7twKoynd
OFgh4DSjERHrnHTYYRiaOdC91tlqff1nEMlWQV/aG+gPSzkKJSJiB8T2DwrHbJMLE6OeauoX67mk
WeLGE4gVMtwe9QLLUpzr/eAmW1oNz3jebjRwjXLCS2VoUAjBT9581p9I4wBah6XGv5teaZfiKb8n
xzXaw5sjMi96+o9DMaT295oAWEZUoZzZqaUWwb1i8avlCSKqBp3mgAQjvZFR/ydHaqHKJWoQbVsp
WMu2JYKj9XulQaTzDDszQeBwiX2BgFyfLtwWh5ou+TOFEbBLJ+Of955xSDPPU6BcbWEQXjxfKPyk
k23RqxJvYYcocuZOfcCVTDWf+HX7kHRQ9GYFfca7TW6axheOw5UjuRIObSiSjc46xOWtvVpTGxXe
pxYbwiMFy8IgEg9OgEGV5712r1MubpLsbagnDi+wGxtpqogDI1yCzPHlQFcPRSQDoKLT+vYRTnIl
K8a0yoRPz3v+6itackjVD67MDWr0EsSzhrALSgqtvceLXMtpj4jl0vgJOztwaUEa7QDlamO7qTw8
zcCb90WIj7eTGpsZ9WWrrq6VIZ8jkUDfE1GeK0lrhJ/BcZ+lJqA0UFmQkXdpASjJMwgta3jFwCfn
JNU9plWebvOxmVn8yFqp1sXcLHXHg6DFXJH9f8VIW++xYmZrYCYjumjQE+kpL3ecVUWbzl2wNF7c
0DDnUTgreegIqCOCcE3BDnBprOSJGv+8RPUWOdkLY1kT01lSEC1c/ovr41v4gDjmBdgjAMotVN8v
GFDB+TqE1zw721kLEmeil+JB1kpP6hp/3CkDItNya4bSJBjdabQ5aSzjqkBHlRQdbl97lkMHt77M
sBrTwqnYN6sHp/H4iqdtl/9OqQ2TCOVqnoSAm5Jq2/H7Md+d4NZMdgxc8SOIweygq2B0fPIb8Nuf
wHfEPx2fqbvpgmN7cJhpbr6CuBa8GBCMhCwwU+5DOmrrGxWd5xCkyq9FPnKd7LnvlOOQncXtwgqn
5Km0frxCr94OBxZvlK0mEONDrjTD8V3wf9E7vVU7dG3CHrA+XV6nnUksrfP4u8Xr88RpLrcIVETl
N1w4H5sKTMhwmiXeSPAUhp2r1HpLAhJQTmgMwPMkQmRJcm9mf9ZUKRjWYWZnArur2bYT+yEddjxi
/gF9Is8W2MPv1pob8/DoODdCr8x/O//PQmyLLYSBLoHpkQ3py70cUZTpS20sJUCNFp5DXsqYP9Kq
sVjaNE7V4CgWkTfvZgHJWuNV3LRlxXLoXvEXS8SYbCGjaX73LHoYarKlP3GDQ1YOs9DKAIYsvsjI
pz7PEiOQ2iWMXvAjsKgr4OTTahIZv9TMw6kAcbf2PZzGRlKukE48T3GIjcpj476+rR5opo6gijQO
HbXnot8zf12Mm9iQS5qJxflaQ3ELoKuSQIMmxxmnNwJqRY6RhYRBabyfBp+GsZEWSTjTv3kkBZZf
PlxqeCF307AoqWvlzMypEcvK16gyUd9G5TNvv0djmNej3xbSf/L3elU4youF4/oifjLlHNZ+0C9Y
bPDxmNEU+0R6AnTvN6IP4nsOT+q0TED0sva30THooFKQl0Mls3NCapeVxPnGTb8HnBEh200R0j8X
aqk9RPpmwGOBB4js8CoXCfOrSe1etQuwGDMorRt1bl46sMa5y5PKZ5RfE4vGaTL/QiuVtkw65+LJ
Y8SQcwR7yWQfbExWhB7k49VBmPtRxYUqcCOO6KJbJXiT74PWA+c6PU1Fa1ZhU5Eo2NytLqqOO7us
ThMpEMrXr6Y1bs8W3PJF7FBk/sOEo78yPuGPSo+opg30WcEX91dpvXzyusZJxvNs0XR3+NXptXaB
oNcJGjw3NIMm6EyGIOxKTFu/FHIJxF8B3385uKAOBbYe3uZjHj2bTzsHW0WDqCMKf/ih6SSB2LjB
BrdY0VXyzb1+tqzoj3zKM1zuQncd7i9Ge6OPmC9DUzMSKXAwmltr7FHgIdC+iWBj1B6wGiPAKwSI
gUx30R37JsGXNTstfAD1/VCbHTfMuWwQUfpIhep1M42AHd/iJTadV7R+PMyifRKLlbzVGElMYAzg
vaaf0JwfYYUexnlm4tPM2quOT33HCY9VG4hS6tsxble6vN1K6ffoq0SO9LqkYPwu5e9T79V+tJe/
UaPBcj9BlvVTmxjgEyRA21ROE4/5NWQgTPx/RYH7f+RCajV9ZbxA/zIO79ulD2RSTAi9+MW8RJY5
d6JswJDGFTb/EIkCXg8/m9fTx+1H+8qpnT6c8DnLEaHVowvSclYbY0pvcqrfJh9zITswFMAUk86B
CXNC2QoxXulMAh4qsR57SpDnBHowlkYzIdFKT/zzgfrkj8c3Hd1aCKqcVllpPS6DdxhpBm7gKtmk
fZlqWUg0G5zViR6qTSFIeqbnRXlkmFPyvD59SW0KjaTQ43uJmtw3JNRiIRhWyZQguHkU0wavmpeI
fYuLJuf1ceRMXjpBARrUxqd/nIR42LcSR8GKuOrILDVY3CsfbJreO18sMXV61qSZppeIR9/iGknr
MzARCrZkY7KfMP0n9BXGGwBGIkHljJE27PIuEzBI6tD+eM6kSGIkorUkjsCAlwRnCPaRv0sjrs2S
EM88u+4e/HaDt1gaBbFFU4Wg09UCXOe84xfewpI7PNWDyKZzHMbYoRZobEoWskQLxwMmDrX9dRP4
2DC5Dw4bh2bg5hsRg1ZBWp+Pz7wNH4HILB3Ey9MaSnYkgz6YJodlICZeXGYRGhB3NYUUaOec1Rkd
Fls9reL91grx9Pz011zpzAY9YvQ5S+oiZ1QwqvNMeCHw4FFALkKM3bFXuJDE9TFDpfr4NRkS8fOo
yZPph1ldKGYW0Mx15FOHypg+OyRGKBPDvtNq2Se8Z0sRcR/K0ayzXdyYlyaQjucXWzHwa1pylyeJ
nCgsevzKi74juGVlSOUFzO5KCM8sCNNwiiJQKJJeN/5bYUNGA4M4u7tnVzxZry/er+JsoVLgKOJH
iHK3n6MxMLd0XL3Nwu3tD3lLPjNx4PccFKpSlaIg3GU5Nw7p82/voFdTCHFF9SVhz+wyhl51gg8E
PXpXI+8tvRJO8xBG
`protect end_protected

