

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g8r/7sde1iyR0STftzcYOcdH/3R+q3JXUCZQpPRz/VObMWWqrxZsHW7lLAXgWiq4LPjiaWHF+vPi
AECUpOzjEg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WO7DgZGyzsVW5LpO/Eo3jPkPwTvvisAARwFpj2ThVqKHqWqYz+cfigwxmDVkJRua0WFfWGJfALzZ
wH9inJ1f2CNVtaotQX0lZ5c362qhx1ui46ZI+45doxR7KHnJYjtJt0bjBJRxWiG1ibF5Ibq1Vypq
pWOz4nlaE+qETERLz8k=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l/QRLOPuCKHCQg9QTQMR7jaNBVIni483AUdnDJbuUz9G/TnesoE+ckhte/F0j4T0BnQXltD2Tnpx
iVDzBTduCY+rrKSf4BDtqZQWJixR7872ZqBGdzwwbc3lZRFia4ykuBaMAKWhpB3egOY8nll78wm0
IlvLFfiXsSWw6JaF5MsY2IumW7cs9XxYvVrO4NCsL96xF17E8iSUPKLB2HRiNN0435RV6oaVGuFP
6dDpS/axWCBwmIlrR1/AJYmARBBTb/HJMKmuWtKGLARg5e4GekIKL5niXM5CaBOaK1N2RkA9p8cv
1ZaBmtz4Yz5BlqinZppN0hM7m21yUJeY3vk0LA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SIPc+Pr9P1+9JsBFlLDSyhr56wAGsokSTHVRjBnYtNQRv2Cm5GaMw9a4/GZLBPH4gUodqp7zeOyV
CWSlDOlDpo/32Shb9Z69I9aAKcLsfexMWcoMotgY/7e+Q0QLV7cYrd/z/ObLMAAUU5jChSdYnzlS
+7VMeKlMLT2qVS51Zgk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Pasliv+gc6ueSrwDi8CYMLQuGH7X/hw+ACS+RP+c7r6sIaXZM3oFjtvI/1vDkQwJt1DRpzLcGPpf
nX1SRapBAYpWFD/ImY3wBJ8C2f4pksIHaMrjA1wpWFNCX9VFKYl/zBBBB3CLfQ/oAH+HyUHSfuky
Q11Q+PE56TbXHxVkPRT3n1MMU6Dz1GmFhKhauQh4dtuk68rUVbIj1iVkOAV/24pJz11QsRqZTsaY
omz9cQKbLN2TrFSoAkUJgbRAynTACbr8zvFgBQybG7Ha8oZ9TmwUMCoCzJ51TocJML5Wa3hez2Gv
PJVH7QQFGyJyKD2iA/1Cm51lM15588DZ6VeZ5w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fitjjbF+Uadig+MOn0ROwIXMOGmAsKF+ai2aPPzK1LuoHEybEUjV3Ow+S4tCN3XQ0vXQwlJ9qrkh
XjAxKmcndINrHSnUQUnxaTr0eUO3vd2WqvZ7Ju0XJDR4+PjdZ4oM1DsnXl/hmdtnOjsCyplOs60m
9W9MbYlqrIN0NheOVo+Zaea/RQAZCCYgUcu9j2btQONsOmorBJXqpSvBA2MTjrhGQONrMBGpIptc
e9X97HPIpJ+DVROxngOntMcwYa41rY0znA1gjAtxPvzggRWl9qqUkQqmAlth9BjTr5K+UBTT1aTi
YdQaO4qgUwRsHEtK35jViPEl7DIlbfQ25Evt2A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16112)
`protect data_block
Gn3q1/b6Uzor+Ot9pFP8ZWE+/6WatgM/LOmlVtVol7d194t7Sg85QRbsaMB6M5iXbPNM6MA/JGic
uYyv7ujpKQwH4Ch4uFollr74QYUJbH+0GdcOihuxDmhM14m8n8PYiLBBbov6swhTw1C5stjWCGrN
BO/UezUs9tUilTB8dOd04LOuG3e6McyL7+tk3czOPVQ5bTtYbbGpakrUVWoMo/O0KqkqtnlAbWRA
ormqTiLE8puB6nVT8REf+Aa/HUMCYmluYINewMo7DbrNdVeWzBV4kJiEgpwWYHuewefhZnvP6qY/
Ruyn702hI3CqCu6VlofOAMoEzOGbq1tU18RoZ/4MYnQonL0NIAmGmhiSvOp82Zk0U7BNSKwhWoTX
dy3eD8fe1lK0Do9GlUfMWiscWr2sQl/l4FCf/WNkhmomca4z+UddBtfb14XoSR1V54XRMnfl4gjo
CbP+OukP/Pe/N5+b5IKMkMj4g/e6fdnj+fK1Cp36Qb9vDzWTWOC/i9GQ06/VtRxwSYsNimvPAzXm
7nQXB+Gv4nvgjZ3Rm1PcDUwLNraqjAdevpRBt0h2oQGYliPRtb79N8QvAp41JXGyxB7u4uhRkY5V
ikpSWS/nXC5ATkFfCoXna8fddvimDFz2RIOM9SWeVXcRDVIP4GLRVZj80bucGCB2ojYgtNpxemk7
V0NC/EpgFTt1TnVMH2ecmnbR4LZqCtGmkToixqezi2PCSrAJyHjxdEyRJpmnISbXFEpbr7Pdim71
MZ3N9W5+wZkz3henQ3H5ylDWxKR9TWuDT5cbonXzCmIPPWPPqyDOWJfOVEIUIKzBhKejKNN/71RR
loivbE/99QTlNgMTfSUrxF8qC0jxYQgJAhS1DRHkhk11xuyppruTz6mKwurqe8LlHBqEG+jh2e9n
WATZPbAf8MK0cPrWRFVADpOw3lixEXiAmJ0Svvuj1SQOFAL0jpTAdAqdd0el1iAVSYcGgrVFO8/r
iTs7+hvYLK9tMdjMoh+VYPdy1fRiWQmqYKpb4ywnXgiSEgbMQ7JQlfbXrqRdCouKZ0qVn5R19+rQ
7nbbGEs8e+JYPs1lD1y/jFGJwl9n0DYucaNGkl781L08YN/tMGrrwizzs6yIYDcb4GwMDvk2Ufou
d/0SLqRrvpMFi0s4snp14pqGpo1tDqFU+OhZcTwUDDFVNrcRtEvMn1hf/Jv5GQb1kYSNmfxhwG5J
Z9IN99i9ZqBfjzMC4lDL7X0SNxHQTkY7yxDdwUa5J4t4aITqvDMmhejk9eXi1A7HhXcTqcVrUIRE
sm2mjsiPlk6JiWcDX9D8FCbbuwre0JC8fbRyNUPYe2GUmNyQ9LWgmqeaBrLF3WvSx7vxM9v6AOIJ
iZBGwi7hvm4X87TYuABa64wQMlHehGa1coborYlhnJGdXkUH4GvhhN9LN1vSEmEHvm5GvFI7+3H3
5FtCLwuJXZD9j65c8tIPSnRCuvKAE+wPtxMW8eT8FuhaKOrV7pi9Me7idXTi86yc9X9hWWfmmME+
Es40H2cyzMIt5c2vHPCS2J3ULlz0cr9OA5vWsWFNVpGEbUQT1RgZk+TDTzzh9l08vhepCbAI8LVv
3xJx7k71w9VldTaVL85YjtykOFNdBmv+e1WsMPz2hextHL5mpzKK3sDGMn4soTC4w5OtSEWoArOS
jFQK4kvDo1yuZspp+iSuglBLql8A0FoYBHG4lS2BncWjEhrAr4tjvdjr6ZVmQPA1JXlFGh/sXrtQ
eksHNf1VKTfhKBl1Xi84Keeei6AK67ucADmwW4FSCSJZqlqTPbjbWlsCBma/BMsamC7HwKOxrLd0
51YGgTjTqu++1KE+acAHOPY95e6U8jN6fQCLDiq0kwO8Skwrs3dSwihySb/HKQMTNMGm8tcaTj2j
EWp8wtqrKkfMD4IOEkF3yr4MbKh4tdx6H1EZ0sQaesdAhz40zpCHpmOafV7dcEzvTSuBK8fQYeyM
z7fFjvX5ghBZ9dYwtfwfNhjV3h5TCbFo3r6/Zv94JzovrxNDWwyXJUUt9u3O1hTdVHWqUK8r4im5
0BxzmhtkXL6ap5lLqsuvX7e5rhHAvW8OxGxe0CKXti1vQeMyJ2axM17mGqnVV7A1YbNNBQA4qqHW
Ad81k2R8sVIfHxcK3l4Onn66SVgTZUp4LtkO8LnIaSviWjoit9jeFeURmeQ1u0cm5fczCsQPc49X
l30cz7eoPcrXbrAK/xtWPd/79lQKvEjnVrXjucd23M39tFRxR/neSnequMnHyE4VswJ5dIv2ZF0P
1MdDmKndHjH49Zapps9XeQJn7SQ+8JYom3iaXx5gV0iZEPLRpWhidQmug+rY89oS3jnTGLtdQDhy
Ve/OrzqKWZ044UvxgcpqGggL4m5+uXf/0K4NIhbQ/QGVsBIJ2+GTSwVCsT9DYtXt2KtS+bnKr14T
fUgfnLG2TfUC/9oKuS4nqTnHijhM71oeE1nBJWnpaj1tvgxXixtolbLwu2m2xS3nToRX+nI5j/E8
3L/B4iSCwiJHNYKetffCqDIU9dEjpxRjqLOYAk9+9yrF3vAwDWaV3GC6ybjKABsD9nJAzG1uEgSn
6GWYk2t56J4CPElZR/xFbk4YOf6jUwF/OwCwVoUrnCqE8Ap/S7DChz0b2TnRkTRU9GbzD9mB+Ve0
efNU3Z2jTmMrO1aTes2W1x4EiRD6yNR57jPFnFSJWS6lwo51EaZLs43Ht7y6eH8e8bsUJEmvqNPO
j5l94+6q84XR+ZtM6GSUt0xVzba98K+m4eKf38Dwfq3zT8B16Iazo/7SxLiroVQzXAUInZem+BRP
DmYy8Hhfz9H4KwdhXD/+qto4zeKnVTROmCTLPhXDfVBnnWM2J3tNcpPp904eusNyINOGDbq0RWPa
g3cGvz2l8QayMZRpz14gFqqkx1ioJ/H17+oiYp0lN8CueIQ1JmFns7hNgKLHZ5Zl2Jp6xSiV5xmf
TWtRVVlIF0Jdm2wtrGeP8QDxVbloWIdjhvSut2iJ6izmjuraFwiCRe4E65y2iBYQNMjAd0Qd4foY
fajkDAvsarJPDyvEMPe/z618c+xWt+w4lFMMz+qc4XbfQ7UngzeirDPgy/J5PXqTqNzgm4RYDN8h
/kSA1PQhE2EKa7LafqUjjJukipSAYnYFBX2wPYw38QSqpKkeVERtQqmP6sFnB0U1anjGKkz0MHX1
9tYuRO7wYFfAiC0o3JPq7Mu5rfl/pRw22WjyajJd/p5RCE/B5AcY3LV2wzzK0UPcq60DGZ1HYWpM
edqknXZO/YmDMS8ulJ7wyojYr299qON4OogG69gdIn4NtpUMwdSpkKrgaXgf2qSUBcQcfPbu/6Jj
KAnx7uBwyyEJ53MwXzi+C8FG1uOifnShwvv+VEuRrDRBzGBbnhLsWngVd93j+JCQBxfcgy/cJiMx
0mYp/KPrOQ+xe3YApU0DKWV+LxXe+yA64HGwxJP45CzHUwYI8NgdVXdFNbl5rqXEIjUuIBDDHvv0
bgO0c+qXdL9nz7ETPoanZfWbTA9/1W+TAsmA118DAV8eXYL9PVyjUNV5LAMP7QoLNF5CDXgLEC1Z
oP0rjG+n/nXJzr1Y/MubEJyYItOns4JgNTbhNI7fPCzqv/81NB9iUnVNEGw2DMHq6qD2hcZtqo9w
FnSmUyxLAn9ynFxiwfk+ISMHmHIMJ5f8KCcGYG5l3U2NN3WjKYKxu8oAKo4SsjKNN2vHY0n4NiOo
YpKW4Ada6J6FbXOLhGqemyvhlBOkFoAZV9oZz3uEzyi6ThpQtT1Ku/lvb77dHfBX2CHR1MO3bmLp
YCh8nACWYcLhKPpdyRloXjCZGAxXW86U59Ai20fmozBM1f0vQBPuqAB/pt67C5zNCHp4g4yoZkQa
OgGaUsU/3oSQOgRDK+hSYGF6yoipBr9bL+H1ClL1M/rEKTD/EEP6KV8+sG+0lkCbvpXWU4tlsTIG
I3bVZsr45Wix2x6eIwKafURTuPTMTlSfSccslS+mR07ARYfXivg7WO+DOPo50Mh133mXwOHBv+NZ
9t0UUHoMR6It3bFILW2m7OKpW1r3bfsSXz4ZRZA+k+53HMTdQJRnhMudUUrxsMkyAJs4jX6/mpkF
W2ujlwJsInrCWIdf+0I1ciHPW3exhm2ImYMVDKJOUfMZZnycfzKVocKMjBWGwrUYD6WJvN3Tz60i
ZXpspoO1hNehg8VwBMmvAK1QGCSnnrf2AWpE/zE3UTFInjLsyOqKqiL+E8MsUWPY7p1kigXCrNNI
x1PbUk8EROf8IMU1J0eF+nkqbuz7nSKj8buaYIVtjru78Zq1dQk9Sety6hWh79qVk1JXBNETbK1q
zAApyMMc6iDmSKzU+aemCS5BHKzojj+RKO8Pf0bTLu86K4F62LOLonWsV3liJvskENFn+OYksuRt
IW82RhPHS+TdNkctEkb5HHA11CloMoIUUj4o1jdpoOh2cL2cChAPn1/oByS+j2a6RYTE0sXqkMrP
2wcIqhPHrR4yN4S5PzghhlfVXB87TAn66ycp6kvCVknXIvaUr+GwOSywOCPmj7zWmvn7OlaReWw+
Htq/nJlZPR/Odo0yTrjSg2dmkDlHksSSsajNGfvaBe2vJ2fy5dkoBT6Gfc1w9vsDseBCrnX1S9/w
1Cemly16Z4q7dCBkOp7aeF0vyZjvGM24gI0D9XAQKqQHZBObG9ckQzWhaXMDHlbGMfK/gkv3i/EQ
qHZxyTp4mDmESpUWYxO+b53FwPzU4Z3yInq1KIW2k2F7nyehP9gVR1ZxkykQhMc8jcWSzScxVPcn
kNDv3AMB8YMZKBn+zuhFTPCEOxLHsZBBXfgZm9eQ0NTlgVyQT2T7qfypR+Mp3xYjOTn5/v/lSBb1
0Y10BYbKn+c5JMbUzIvkQpV4vX+PGay8ejBXygyMV9diQX1ybymj6FttJlxAj5nvXKEWeOh/dIHF
8mcoNpbAl4n3zSNHtVVPeo7++X5/DaiP+B7FKHJDWAm8Lz4tKWAEbfirzOnA5Cbpp/Gyy0WSjqlc
Ys2i03sA5I8BYQyh1vfvhcKcTX/+7GaE92yVMn7Db36J69dnLgtsoXGcwZZeskKm36QQFvo79ddm
p80tSZsGTLHNd2NfpmqzLOOKd3/uOzp0oKkO59ybmzpM19YP9jU620e1ij6ComMxH0O9+Tett0+t
4f/NPlcE7NjtJFENmztTPWE4rlkAHifZ1f0qnl1yuOf3ryUGxwxv/V9V3P/4tRU5gMn2olHJ+45c
qAaMsEVkcGSnrPuT0hpWvWKWcW05uOs/rEm137NCX5VS3Q/gtXLthxM4nFNV1r+ySFXE8SnU2XxU
1yKEXbfO8LbEpqdXHSbTxnTTcQouRYazWfl8Qi8XVymMGWn1lPBub84KcNr/q1RRd+rg5idYjHOF
cyCWJlOwLgtEiuNJFuHRlDQRBBgPCRAvCEcETI6IHlhLhWTWkIShLXRCeXZvYmc/MDUEvmu9o2Ry
t03lnOFHLiuVmf6gsniEv4kPeTj78p6XrbiUWvz9tZnP21SRjUBYg5a9740sRRvPCc3HzYjMCYnR
j02V68WpeTOKHArCv5YQvPXd44F6pIGkNnJLfL++uyNKDSellNE0Zq+DZLRi6oPg3hfsmmAfLayX
a0BS+YfgxG5k4gR1/Ew8EbsuNo1ecIa108RDIUa+1lhwGq60ZpB3YjnSEUf1DrtnNGSqr8qfXvuC
oSp8L9wYrkgrJD+9ccRC0+G265mowiJr1TmqX823JEwX7ICrtpmG7nCKYbz0eACFkfMr+bbQTbEQ
rdm9cnfz56mtPM/EgvfadJzhhqA8Aby2OVcyQ6krppfP/0u2pV0Zrw+jyd9QgONjt3txNsNw21pS
yUKt9Cdt7FR10rLf6nNVd+7+BYa/vGNpyikwH6H3itFyabG8BkIiacgMrDFui4YyeoQNlV0U4VL0
FufUUFZ4izQRsxndyBYfeXKUHx4qe/OeBHnq5ILhBLHs6OWXVPboUGIMw3PXsdh2KdEYP9vOMPSJ
coETG7KhfhPdLrceFAyzynk39xIRHhLRdTs8tRwo8laFO7Sm3JPjMEZ+YPsasXAd1M8YsrbDDbPL
Ul/ORieKPw54OqB3TP0DnvQRv3kWzVB1TgaxFqt1xoroT/n91+wsdWS1DLHY4Gz8lI7F/tHCvGg0
RFyHksU4tpTAwunAbcH1Xi751/qEng4WHQBNPIqDO/t+0RbZqygmJVZ8B4Yvv5sTRsJXc3REvnVw
wd1z+/UiVAmKdrIhQgRsLADQAHjAdcRRvLhEw/GsOhF4Xal5VzPpE6IU3GGSXvkVv9hRCvd2uevm
3EENf/CWdI1lI0ormZPkmyFu0bu2SarXZ0xlhEJ/Jnycxwu8a3tZrogC7IZYBUNtELpaGjm60IDZ
tHaXmuAOy8c7oStij3R0P1E7bihE5Klk9yqZwRPOvSMTIFJqi3qbLJG8AVGfcfPqNPVKj82BGGLy
EY+spnQIClD4lL+3kG11AJJcGFN25CtGmbpmPgui0g6gEVLRMnehSVUJETp4fSPX6ylClzVB/CSv
LbnEyykbizzwAuvJhS6QxywpcANbRrw2cNw8KxgCjI5VObgNvuHkPlcjAVEsEgtrfYX0aBvfVQKO
S3TY58C9d3gBv3jmKQoOjpIhgURoSstQ7XV/SFohOoPn9ltbfLD16sOTvZz1Eg8SD/Y896saTSRy
H3hOfZ6Vqg3dxFtn0ztQG7lJSMGa3akxNV+FKoksIxS5QJwElIUXp/q5X+28AYrfYHhS/9wEJUhH
suz2iARdQHrx00TXf1ypROsE7Du4rlQA66uKm9tYoSmzymKJ9r2P9y2/o0DtqpwwJLGoLL5K1pPN
ScM4y4R3R6Y3CUSfZ9LkPIZ+Z54FtAuYgcFEkinVbHfsNjWuokS+bXVsDpZZudgbEPYlIdrlOpPs
iEsqvTzUf9/b2M06m76TG6MRb2nwMEVS5P/xRTT7O5jlq8GNs/AjQby991le26eyKWs+DTNmCxU3
nLe4z+AuNs5vhtiR8cPenUHqMwgCViILoSF2nh0syCZnljgDFHdy+bJd9rAZ39qkt4DUwgrgkUA2
Wxpqf/Q89vuRiCMzBVCB2xrxjBlr6F98LBU/DCP/yT0lpoztvhr4gPbUiypRgDlb0MFDm21X+953
y5z7Emd0kaTd4TeHx+Yd5ViPERwGvyLQcaQK7CDyw7ViDdOYogbAk941RhtwszvhcrEZf+UNcR3S
joOrKXNwQhp2xyWG/JCnd8r0R76ofKadIuA38+OHeBRElzdACkzYadxVqb9sG3KDg8BPmjsqG3/c
NC55Jm3F0y0xqDFmE+MbdpLGd1VWEzNJrkTMRQUdRaxO03wgSLP7DTWz4kXLAzBckxEImNr7xOSq
CopytFqpzWQgVpuwoQsK+Bzyk251cuDruZfkMoRU406OjPs59fprkCRbPGmSV+7c9Iz/oPL4anok
WzkxhFXtghY66siSf8ti4WGHb7B6osKW9+K+K0WNtwFIXB0U28E3qOiTGJqmyOs7FhYlEnlvnTSP
ZwUAX5jZ05o4creB0DMYCZBNzNRYM18Xtq1tt1e05j5fkmFyJjRBw1Q2PpeGiVSRbOv2cexV9zHb
SnKTb98zlP5EILh/z/mchUiqSj6s/RRtiggbDO/xwkngg1rTgsDEswkXmisKmbuRLtXEjVXcZGpo
3uu8AD+tlLL5Dtw3A8/z4VoDsl5H4K5eYxVmCq/avcAzOkw14HtfTgo42EgTIW/o24do16LEQ3gn
DpcMWACrbOp3SxZ5waQSFbZYbIlqrmT+ErAAgYJbpGt6AlT+q9teTIsHU0EWcTXGV0jeEtakTteH
kI89ZSnmGYpHovIGNKiTFfR8RzPC/sJaabxMDo2tyiwksw5fCS8MY4AUESDKIELJwzDcwaOd+6z3
RDffpSqUyw04GUyi6J8FpUb/hCYn3ZT+LQAA06rxaIT/0OlGpF0NuGK2ife6kcbKUyoazcNuSHOv
bdB6rPHnZbSmk/N3prCRdxhbapDxwHe7VG5Rf+MtONMKGL3OuvArid0pmyxqkd0RZnB3zqM8z7Sj
lFhp/YmDqi8zWolJA4OfXazvETD0vi5Sr66N48NLom96K2pSFxSI3AHc3LCoZBpXwHs6Mr6BTu5m
ortQpP47xfwIGypazYTMjSp3ZLNq6COC2ubIRQWO1pMGlPOThgcDX6bJ4UuSZTkPSBsmfP5neeeI
zU1bPu/tcB4Cmx11/9oi9eY8+k5K8N2XwptbggKSOSvZ1lhmPaw7ebUcNhh6nYSonfNGsoLI4fil
RMOQZY400Hax5uqJm4GQdbD/oKUON+S/PgJwBruIPbu8gtvioqude48+aReB+M1wlwstCsgjouth
btfLUOKKu3pK250gNYJLVPpfsBdZ7ZFQpivWsT0XcSV6cd80xYmjZMQFDip3gbOw/ZQtmKTlTb4f
y7Awn0cwd5Jd0SXqi6l7LcNqUNIw9PH/wPPhm+MLKQw0FgoS3eVsk1feRArCqjom+6HLLkNaDTBo
m/LIWYOv7L6O7vrIh0lZnXR4PUwSWjrjKYZUOroKfCqdGW/tNC2yb8W5fhRPtR4WlrGmm48hOejM
RM0ZqUtrGqRic/dKRkNtUJBvRurjaz8nU6w0dvDDflqkx7Il9uZ0jZBKtRqhS/Y2gG06y7Rs9OMc
zwLsVvPdnxFF/uNcfu+KFPaxLsuiZDvizsH1yoLr/ix5IsbUXzXPkFM5S2sGsAaFFD7AWY2zKxoQ
/FXNgt4lQYxqb9e/BMz5U6lHad2t6ODu3ElCnCOZHxyIUPJIWr2X16PVYm3hh9qtfO1PssvOXhN4
x8XSa0bBFWJqYxncWb0hvUHPykyVwqmc1Rigy4v+9I4a8UQ2MspB+YyE6hcO2IecfLhHDLAuJhyF
tmLP4LsNOZqzEwdiRCx5v35mlHKW5dKaTPmBi81usqymsEioVhMtdaV/XCI7LXvwNrWQVvDWuqST
r4Kwe3la48JSUxowgmdygo8p+Wd/dQboDu1X7oq3zCmgr7S2G5XEIBDEMDGPkzFif0E2M7mbqc4V
tcAOCPC1pOOPjP6OpcmejddXgE9lyQQN2BVRWLV7M49L8e+o0DtzgNUDIYH1ZsmhstAMmfydluBC
/l4EdZE3jU5wViFAXei2Bc/T4HhIczwvlvkjydQ+fkCKNNvHzTFVumoWK8bR65v9oQxbBzTxcGRq
cr1bJUuSRyNE/DRAm2e7vSGJZh5uRwZGC5CdtNnQ206EaQz+BxFTBRKUcWwdVikBXyaALc/wQZ4J
pnftco93olGwIK7t0Hmd+/rLoMn3WM354BrFS1kbZYUIcX+/15YrGI3dVQZrKIqegP4AhnmIDKpQ
kubyMnNrSpdmBpfSsntcpUZenXJbAetpvYkhkAnlXKB41+hCPfODozeYwHA3VazXxBbVcCVTe4FE
GIoyBSjGMdMJ8gcA/FkJHmdy1BrTIpPwderrks4WSIdRu3vAgduj+UBlekGRBlUlk6VXhqd78CE8
rP2VasubJsEJsDIc0+LmlZBL+yZornMGwOL2lgn66bQruHSEYj4t2jidFESpCAiGwYjuQNqC57l8
nkaWWia4mx+kray3rEJBrAuTgcxFHF0ZFc+vba35Nvp0byhTphr6+Qfy6iwaNFotnoXWJLhQ1oNS
LOeJdsdyVFi6vtVgHgLj8qWtS/oTNxayWN21nqvp6kLDBb7JIT/jGjlAZ9MXgK/gRaG3qQYp4WCl
JxjWBAuyiYIgYeELGU8083aBwdKdd7wsaCbG0hyWyXedTVULbxLqM8IzBdm/pYnVOwvowK1hEQDC
L1epZTb0FOyNFzoybmR3X3T8G4UoptehgCI+7/LQLvrlr2zroipAeRS4bv1ywN7cGHNkfVEHiTIW
Ci2gGOlrU2vdHufWJIvxdcMHRrGIFfb3LXv5kHSLSdZObqA0eA+uYRZBxOAZ7/mPKJf0ahGp6i9h
XkY/OiXDQLYQH40gQDfPwATctlg49/k4nEeIvPJBuFbMqFXnMRyPgn7IOZ4ZBnpKROxlAg2Cdg2t
j8ahwtRVk3lkwBYR2NcXKF7ThPAkSCYzfvwR0Tl+PISpIskRbTdXZB1khvtlS6/Q9aFlo0a+EMtx
tisNTBVTZQQ04uTAoBPzyRGYA+j7dmPWLVPJYRS/quKGHHscufqMw1VyorYEJ4MbosNy52AA/ttj
aLznA9JTJO5ruSJ63aiw0g6rjSvZqvw8Pv2gDeT/Qf0SIw/nVoynpOHl2Qox5Zpk9T18ic7QKzA1
Rckau20sNhnThoEuDx52AW1iO6PSLH2AjAawdjUt4TAk+CAv8EYzY6hX8n6BUF2/3iOmKdkG/VFc
Xs3GvxT3PGdmujyt28XzQMhY1O5J01LAFxjDURcSSrEf0fDaqMbQNe00YcoP8aw4aGKuh7Pj7LsB
IODn4bAmfGe1WclYk01IzLbQae7T07PZE+B+TESVAIUzEDZjSCj22rm/9LQwd7zTQVWC+xw9Y/Yl
y1tUye7HsJMWJupxVtMOfvbaST6ubgfGzhvuisUxeiz0jnW0z8URCb9EU/0gOuGqOZFFbWDuDTs1
vN+vGJ2dOfKIZpFtLXEPJLEejlu8ZJhLA91F1fGVQXC2PU1ZCOiJvq+bZfdcWtbhwIFfdbPwA5dX
oStoqpumhnHPbdKH8/a93fviz/ciAXGbyOLDcYUjb03/OYD65SicOGa7itz+LzJtBsFg2Pg50Hgo
MbqccEZsicvJtKaJLBuykZMKZvZ73L6ByZj6Rkgg1Jf4z9AuN3pkLDPtPQHTCsxlkIVwFKxV/G89
/Z0IMyNAHsjzR405b9KwtTU+2GLU4QRgUZlFFeWF3M2mKI1QcyC2GyHTeQ8NTyAC+XanUiI/W2OS
D4Ho7NMSdeArLkSdoK32lEIIhqKf/ru+cP7E92VUR5ryE1ws3FM6XOPwyo7X93IEiQH2zYaJT7ow
5gljhlny+HC4PrCzXcg/w5gMdp46mF2vK7PY6fKGZT8NAhqlNT1z7K4OoHl+lP6WJWdJhHQEPoSA
KpOQMW2xGoOMhXcVyVE3RSRwc5X3YhsBWIa2OcAQLC93f1d9j5uYK6ooNKVLLg35icHsqV6I7Uv0
tJhG7rih9Lhv+bhjpudXp+irSgUNR0YfUKV+ih1BoMrZwkldgpb2M7385dJS8/8z4m+8yhi4fcXe
sqjhCvzo2yFrsy+qBc/MhCRRUVnwhPoOXMoNdbqTuB1yfjV4Cigl9KfUOi8dW7TYgJQ++vdgU3+O
5X0qG1w3PtyXyZ3rN8ecpQNpJz/UHk2Jig0JbQ2BK2ShmT2bNBMhE1aX87B8mOGW9OJxGD0mZwra
58F0Kmauh1ZV0BBosdUmMJ2rXev/XKX0OAcnv6lOTT07z4k3Wvp2Py9QA8y5JpbobXorKtgxojUj
5njX2XahZkcmIAyqKStueWIc9RSC4HtRs/AVstJwSFWd33SjbVoMzTXtTMLEuhcFortxgRitibz6
UQ8mO9aVPAPis3OyUn1WAGbuln7hGEouoGW05gqjatVWVHz5lPqpyqIgL9vGeSTodmMKkNK8/fb6
bMbGroXb70Bm4k4rsh2oG5rr8SB4viMQNwOHIHKT+hn/HDk/1w2mVyY7BnVZIawIHrAArVvjO+FB
CJhFjb/4A64fCpN1PkELl9p/pDPsrX/GPupQiA8CBi2qXO2vt4iK1FOL21eqW6CuFTVklKOvTAbV
K7jsVXBDfqUwRDOdkz3QtdbFc3Ma2inNW1NdeEwq8EAm87S+hN8LrgUk0nWIfsKC/qV8SOa764y2
SUcAMIXHY8wd2t5TM94bbDxISX+I7FwflA1V/16le5NPGgN1DX0hYElC0eeKZuk34txiXcwo4YR2
ebXX27fdFLRbSzx3MM+fgC6rzTmrGJmNuEPPrD6QGvBaMi+a6gfPPJA4XYS2HpCyaK1gYCDHTMvl
vG5SjLlDk+ywqU88GK2KFOBcSwmVdVnJ7ZEVA9d8sf5Xq3yWLbcJjWVx/+gqVGAw0oXXU7ysKAGh
TFHn5npoF3rzKYtq7smcWE9EKZWoW2jEyVrUjCMDPlMldxYnFMHIRbjUB6A9dKynkeVcFi8JBChT
6G4ri5eyOw1BBt8ExYpyvfit4B9uYx9RXZNOHb19AvXvF7xALgCP9f7qnpZTbHfsrWZLFQmewGvi
oiNVcNX9iASPJAfX3ohUuYmxjdetLv/G2dTkD0c39yMeXX5ze5jgj/D6QeeGcwMOAMctwj42Efyq
96h8yUN0X5z5YIgApFNOU1SZaOm0rbMyqqavOecT2aAgUh7pK551M/3Q7s6OeDI2fZlzMcwKTrA0
js0La0pmZH0dBqd+7trJvMPB2bUlseOevMTtIcVoV1HgnczCb9VvKZGv160j+Ir2pLEy/qzdEpib
ClJOM0jP7G/NNw3O6t5Q/QyTjac9qJeEzS67gffyZtlsRc/tHBq5goyKWNp5Wwqx1Jm0J4JLnWYC
h6DLKUo9HoaB4Rzg6KJWhFCUAVv0NWIXsA56d5EcYrxreSXsbRmCkp8qAxD/E5sG0R75GlD2JwDU
pkhXyl52OIzSnOBMCznWorg+QgbElvbNvcrrP7n1SD/wqJFMkgeW2LAPXPr4TfL8UuieqEm4DhOY
iwd2Z5Ri5EM8oDfVRZG0cX602lMuirK1yTvbvax2LiF/x3m48XNC4O1xxs0rkwxZfW5eTlD7itZJ
OQDFWsIoyJ4NBFI43wJC9d80l+r5dM+gCmf+eDBOQpyw4Lh5UBDDldJWH5CAGAy4oLElgt6eP1Pf
rJpedNCrZ+7fC/Y3WaeoE7epb//K3ehtdg6RnMSicTkK1NYmiVdALwkYGVEHPM0oz+aKnypvGbHP
GRjn+R+pVn2JCR3bzW0vrdu4MpwZsXSXXUZI1P/5iYjFb8+qMonha+MwronrVkyGJWO19h4ckQFl
PSpsGNkglrzbTfEoXtSC57/T4pn64LDb4qozYCB5GpO4gtCPW8kTQq1W6kXE5kdtbtslnlJwlENZ
2FWagEJ2OPSlHttr/22FyVyC9oh4GmF1oUpV1ZyqSkwBHrjgWGxdiMyjygHonMllJfNuiBMQMuVL
t4NMXF1mlj//vFC1qdULMFs4PSrSFvmH2070FWexNdDy5G0s++LrQAIm0Px/4rmi1mEInnOoLJFu
iLmlMpnV22ZMFPkpYy0gBBGFnNvFYhtjKI2P/SS9hFzZvWh1EjS93lo6YxIrRH2ArwpwhDXesCA6
Z4PYMUsa4r5EMHmbC/16rjM0/9ZeV0Hxzl3DlxSJOU9bv98ANNpaj8UK2t8VxrDIqqseF4onhjlT
Q/XfSCdTzz04wjqUgT9eXTsDQ3hldn4behNH0R4XmlPaSW648YaCJw7N4hwMlIIFpUvspJy8SC10
mfOhmQ4Bcejew+L5p4o6f+eMhs0lvMRCGKJsmXPWIl9c8A+PPYpHYjhRPRjCU1AFlBZbmT3Q2htL
aU+xKnpE3+3v5ReFs6wvMnildQVwWhfRVCmVPt7XKBHk6jQFxD1Uk0aO1gPdKEUdorJ8deiL9kD3
2PtUNAKfNG8VCPU0m8TDOzSW6YVivh/Hrn2R6Ole1r2yxrPgo3AYZQi4HCIFDd3HjHeJJfSyxLPe
9KMEKBzif49RZyxHoa75FMsG0hbJ0hVpwZZaLpdkha+toodq4FTdvL3fbFPY/7qK/Du/lOTKVHua
L7t+iNflYU9OoXxamET33v13dmlFBYTB44Z5oEqS9DnMghrYRPYuBzEEhwJJJ9snlFOtdqeOOHid
JsPsnfZX2z2o/Nh6Xvk94puvKDcd0xoSw3/eUipvxAYBLeUMnfEih7Cz3chQiweE3JYPfOIysxG9
c+2P63/B+E9nQ8/LxbF5KFWSZx5u/FhPbQGiChUwnksKRXFnc8wEFgEsZ8DPKrbcBgXPEt2I00Uw
TpLfrOsvb55fpL7CgLsEBs6zyAwQlKf7v8NLiV9t5mtUeQiFjExAp629mM1UwcNlhYfDJRyf+5qf
ovYZaMOkDSOGya/DXuk0CG1XpSNBGebOTxKmfstKs/MhRIcGFvaFe2p/x7eZ6xEvcIs03NBgTPqa
ol/+o5lCfMlDZWpvruSSOlFBTJi2mg7L+PLHsife+gqSvjBJI2bkaAwyWA0dQgTDVkpKyCRXYa3u
afZapxdCv3ZJ1Flp/rg3ShXo+FFtAQ7PQ4lWg7byY8yGkoGOvoGNDU01AYhF2ZxXqPl71T3W+Bqx
89U/OjZeMlfGkHzwyfc/JXZr88dbzxvfhykXvLcEzbWGC5gVf1dErmipwjBlPLXEmwLWR0HSGIIe
7ChnKww4EXzZnb3z5bsETM0yIU4IzjUt9F6NlDAu+5Z+eXMV5SdOsEcNjEAIhKQbV8WfbIAVoRd+
ZZ9JqMEuXqM+v2DCVxkCLEIOWHs3Ynbgl5hP9JA9bbTfPSsmO/CSann1M0lO7crXNdgQWJE5sEsn
T2+JFHJvjUJVX81TBey58P0txUTTrl5eACfsbC2zL/Z3UldKD4XpXVXsJILTbGJ008dqMTJ1mV6h
J+JxxR8xBHbI8UiGfYE5ZJIsEYadCWUs9+22j6eWMmUK5HIL6SjpCrmeYnKfuZXuEqp872lkEtA3
7hmzJZc5xDUzFN8lif064dC2DeUVwv6KVKJv8mCnx+IBlZdHkcNaJO8r3aGTUrnCuxepHbT9E9UN
KnHbPPYsILIDXePyXS34RDKiPitAzNMVF175HFclQkMK5nTafSSi3S/NsoW5fR9e1Wmcci86Rx98
EW5ALSuYb+N53UgMB1q5bLkI30vrRFUrRBRMG174b9mbxDZR8isZhR//hgS/Tt78OIm/AIbGxI7p
KB8jT5SA02fsk9OfwyIdDQlTa3nsxWIon98a4bbY1sFXleA0mr+kAbzLptsxnsUNAsiSWruSGfHR
GyyqmGFmBdQcY+9d8OSLi9yF3h6EX7h+sRqocmzpQgvQhu0F1DxjTQ0Lfld3QEotPK012OqA4fZN
iyiUsq3cSb9ewsjL7IORRvxitO0Ff5b0ECWy/om93GJSiYXFxbA7HePacbkCS4Z+j7FdypAFPTnD
+Uo+0e9h+Lhqa9RzXQQGRIdgNXoS900leRHc0vkzhs46wW9u/INzkPUX5uPs5QlWb3pUKVRYRZtj
nUtG8Zd7jP2zduESPxRCJlXyfDVys3VKNanDxXXyc9BlVHNqFWAMSMWTHZdPoFKVuBvh9+2IMwL1
Vl/8pR+yFMtvclvFmdISaNb6PAWfWeGtZUH2lgcVb80mqGGFrA7ncTyo0GQn2ShOewNfZ8HXK5Fr
Wu0YeQrj0KmiNznb3yzh9spcnYm36dpKW8DJj6aiuiDRKVQny7LF5v2vbTdEaj/UwTTx12SeXFCx
Ci3BtZ8a5xyozY5oWvE5vtK9k2jkl7YgcvdqYLcVlyCfFAijMqPlFV11mUTCkSJ3uR6+5RhfPkTa
me8V3dftApeMEV59/z2uU/7Fzas1mwu003mp3rZGaujHl2/nOWK1uAGhvUkYFKUlu2dBqFjXquxx
6etxxJ7WP/yXpLbup5SjNUrZs5r3ij6V3ujF81oEjxWaYHF9fIQSl5U2r4siBjL3orU3eKYTADKu
JuqkxrIsxzTUFsI6Df41p201Cp2MkRV6kkQzgVtUdip3OWE8Dntlq5f5rjMPtY/NuHLaALkTrmY0
m2S++k21IebHv3yZ/iqp0eZbwMEUkVZV0eBBfCWgNaHn1vkdQvss6VDIiggNGJAn0pXWyI+1K2o3
xDQbN4oxj4GG+GqDx4ebRoFbrfI2aert3sJgtyPXCnK/7dfVDYRSVrldyl0ge2pYmpcdEhVciFkp
zmVXzMJ1iKqxgdnn1pVxEFaqw5X1bgHG5RPl4vlU6sr1ZXaAcMZ8ONooyOelzsufWeUTBYeYHb+Z
BJD2rXNmfGBrMAhjDAEsqNXCr1MqjqTfcEwDBBKqtZ5BJmmbnipdOMXgFMYiR6QWFd7sK1d/LNrk
W5NeP1nxmegyF6Vruro9QZUstMqRt2kaO5AfcEZrOQIpStbKXC6Ej9FptO/+W2Vxa+Oh6pVlj+/V
TE8zuEZdEPOEzbs57UUKCokzRaKUTC9LbQlzuBinwuxvmGZJSZf8B9LOqHxo+hMVPBEBU7Kb7M2s
ncShgQN0QwuiruLpa6rsPFgX4dAS8C6qS+Qo4ZmjagpZe2rTW9MhYP4ceLCkYoaWfMTfWVXdkcV0
Vp0J/5K13dKb6YAYzLr/0uZbRD2Kj/aTj4o0dvEUpmwNCzH++TQO+J1XM3gaQ+po5HIswxhLyM/i
OrdBqL3wlfExzN5O604oZXUqqcsbJCkjfiryejTF52lq/UrxP2C/xfyeH28AtiYHoHi1jL1iLe94
bwKmTLTvNcoDDinuUjQZFeIClG/7wMI6W+LIqPszSIXfw3BdBIz6JDlWc2YoVhdn+vvPVsp5TeRS
MVO7sCdneBp2uVyJwChTvM6l61aHgRcehgZ5/nEz33hxxQL7HCh/tg9gr/24Z+Pdkq+Z92ZaVCkd
yE3uYxvIiOEyb55ncks5qLOtspbRUGMna7yt5mEiEX2GWn9Qprx2hcraQENrqVnMj7xraGQnWDBZ
c8JjORHRLUwBVMvjH8djQLPB1GeZbjt4GhUs3l/ra+jEDgTwdLht82dOklezY56NiLeDoF7moNFC
FIsqV+1FgEJcJbtvTTHAvE391aEc+J1d3gk3g+rstB5TjdnTQ7Kq7Ipo6C0jkZySk/pD0xCZDlw1
cxRtLjh7zYyDzsmRn6eUG7m1eJz6kvprtMqzs7wi0oHONeTz8o1guQ8YpJv0lyTNn9WzPwkFWwCV
8cU7xLG0scsUbU3EIQNCnALdJE4c0dqd8CdUDGCw0PgSVtyLUxRheCzG8WKEFdaK3wejq4r2Oozl
YEaLxYRnHc9lUHaA70OJanl636AAijS9kusZtI3DnPffpnOOUdd/0Y2W/XvyZAg24fp5u2ZuPT62
QFeZcYXSNs23Q3shdE2m6BYoovP66Hfo9vQV5yC6qXxNMLZQwEfoITpKNDgoG00t6+K9Rb59Npmv
zmiQdbUtlKnAcybVd7riBisOWtUOiNBNE7hR1lRAD/YvBoHtREBK1JNg/OeLAf1m5Kfsfl0SKd+e
oFBZ9btdJQLdYM3T8VaxA2kwxej79QlvWpYDIndiCL2QnQl7gCx+HzDKMNaZSAC0brVfA9i6GTvj
hfArs+IDlxwNCuJpjGIMoOiY7sk+hytfXFAmxrZTtviAWdNG5OZ9pIj2Td4FWFr+vJYrdGSy2oG0
rz+TboGYSGSg80uZbdgbuKP4apr+QvRWBWObQ1DPR0U2glU9m7/asqtTN0JFmrUwISMIGg4fkgo6
E8pHOfMkzf5se46VXPncH5oseWOZN4Xy1HkFCOp/+915C/baQw+IQVDEt60qCNpwBj/O5wV5EBSv
Jo1eL6VtxOi8FiUwjEMkT+1kXGEHzryLLKv/Mx4PoXLHcd4dnQQrsiXN46E8ZuE9FsVch0NzDygw
RDRLnOFNdVFB9+TuzW8ECMuIgOBfeTVHYn6JFBhu1NE37+r2wtOmOwMG4tqsVzUnuXfUDkABOUtf
Fb2MLdPdun+dWrRIxAijv95sGfaQmXNflueAAvrzNmOjB2tRpSFyPJLr8lTMsgPFTv3qnAJOGUlL
R6u4PdNncbhf6u+K65TSsgjyYxO63WZhJdg4ZZ+LL6+BgUW0Bs9pJcMrWP3Oqv5yjj2fLhuUdBxQ
WibxK+I65sYk/hXesEw0BbY62NFQkLjvoPJuz9drGRJ1GKwZSy+A8wBsvpD7EhxnD1rA1hIkzpBQ
OZafjaUoMNaifkI2K2DTLqm/ZXL0kTFJd8gaxAFryvTCsa112DF1DwMHyg84cVDrw9a+ESwq+cEO
vFHVlqKLMCVUpNbk84Q9aPH1FqnZIpOuqJtUT8bt//1rPA2VwYQcght3fe8BV0DImTpOnxNi75f4
wO0fiGzoQXHNw1NWKJdMsvhWPRB//OsGL7wyRGUoLRuxTNrTOcSvpdZLE8ptyvCf20K328xfqL4i
okRQwiml9Ur6PD8xtRSn+ID/fm8o9Ygg5Wzq1LJQCPmBfz18qS+5T0dzxvRb3CWpA2dGYTDKtbMJ
2V0XJ5I1xxST1vFtnDxLZfHbBcXAsWG7oqYrG5F1NIMENKl0a6FvPpr+xZUkBazOj1Prj8dvLA2P
FGr6Ra6VaWM3Fiio8EftenBVNhyQpJBOzqRuthh+yEjt5sE2rsjqyWgxxFAL+j4N2/WmHkV6RCgR
BhxO1vFCymcdYCfGNFaS7fbXr8gBTEAnjvUxBMMsh+SL038zkhatY9nnt75qbgw2ixgQs/PfKaGN
xm8XEt1Noo+gvzSH2eetX5Q+Ho0afFF4yor4eBS8Mrcx1lc8qmty5qbVamBLe1vfL9lD9ZXrQOYt
/gogXSZTrS/LXHUQ3y7Wpru+rY+K/MVgwvKHEGS5pLo0fGG7DzhlBiUY7OsbEfHUS3Qq4FL8EPAb
gCKXqadLl54qUrNXl/JCDdhOxv2VufWIp+SAy3ZhqWmBIin42V+yOoUcKwUc8n/O10Lq5MQLbdw2
ZJdobLdQSljBYRuAv96+TflD/z8hrmlEOCkSe2NQvdhtQrf9moK2er7vR1F9uTgigfdsLKb2VWpK
ItVywDy0cTZPjrqdKOaM2Jn5sFkmwDFOjpy28fgHIqMOS0vPydKdPfGie6fevqB1xallCaWN7XZe
Mksg3S8LhiRER+AO4fEeKFp96YIoLEevBXTS2dhF200I0PhgTFEmk2bHU9lxjdqkHBJ7csgv3p4A
uX+ThZ+6NjPMqftNuQcAuUGqpfczlPsAvQI9IFRi6IcuD2Q9MkW1d84atgrzuD3WuK8Fb5IsbeVa
JsdzB/cyOhKpLT4nrmrSljOD0/pY9pT8Q6Wqo9qkfoN0B6v+tLczhPv36fzMnYeOK5BzxMjwTJMc
txp9sOIqT83Y7oqoKUIMwfj//FkSuUqjfU40K0Da/+Zotf4mWpddLAGJspVnKjsTw/Y4GTkiq0we
cqf1zMByy4rR5AW00+I/1vZyXNCK4yeXGUTaNZUoWMkJDT8P377mSQ9bOioHlieE30H0e//PPTpd
loJpxx4iGsWQeC3F32fqyXVQRk7RmXTB9LVpdIpk47ORFXOhV+6rvUKT2pw/4139jW+U9v7NzLoe
zMPwXTUcbj7c3ZVrwJA62EiFL74sXEvLoA2xpsTqv64nw3gmnfFRz1bDqh2jomZNQxdusXWuEadh
+RxlEzMmAVbzUuEuru9L1SnvYtCSgEntRcjM/5PWjK22k98gnl/0tqVZlnvulBf0W3h9qG6lyetZ
vaaK5kHWAkNmr2M4qmsvZis3dMcntvvvkeFByyvpKjM3wmtcwwwiDG1H3YSYrY2iWqIfMVsH6N/N
b4IXcdBTzxrN+Fq6VskL57rPMm7AZs+d9oVWV9ScEzRUay/62vp2sQYVPWGflR0yCy+yCcZ7nWP6
4Dq/5SoEr3nzjmuTDxWcNVPDoMKINWyEgLV3IHCAuapk1FJRKGqz9ev5R1k+MM07cNavdW0PAIep
ZHnfAEYebGP4EbEXbjdwx3OWkjlZrBcnq3+4kLYfWGRJ0ZRKCS1lqQ0wwBO2axofLomVQPmeAQmV
idvor8Yi+OBNRkejbBuU4lMf0+eTm9UrXpRcJcz0WIJ/nXTG5VXl23vTemjYZRjj/eVjT5ixqyBJ
4CpE5Rg+CNdvc3mvOVqUyQZ4W3AYFjAa1EW8AsMKXTqMsLVhoNOjUyeqM2pQ1uIUsHzPqnh6ClSQ
zZaJmCFGIjM7FhdOLkZHNgv+Gey5l+rlNMsZRDR0/eBrC4oWtE6bY2uHa9AS3rUhmZJLldnJiYiY
MjKog6oVY94TMNJWWumole6nuLyHZmzuxE6nqR35YSfvqXtohtH5DuuCk5L6XFdEEV42LrnJuXoJ
5rmqCSyIDeTj/2raXBbb6VdZcYK3o1oJ79q+0Ac6vT/YK6HfI/cdWES4YJdis6T5VSAU/LeE7Xgj
sHdJwGq/JmPcOBBy9k/ykuatyorPIePpGQIF7+3NA5KgHUd8ug7Vn0PK6zv1aCdEFHNoD/6huoCZ
K6HtkwBBRf/dns8e2D58qg6JaDED7lhW0fe+CZ3sQjgfT+RhFjqYj4t8RIA1jQlNzwHzJw/u2CKZ
7MfMpMtBu4AuBb+YyaNsu2tweByftjPpvS5W7up9UQT3I/PaYao2qFwORp7BrAWJHFJfMLV+RxOY
r/B5FPX+lZ2Hfi+beb6ttw+2EztmvGB1YqPt57ccE+pdKmD+4JmwG3OFLiFWxJM9IFoE/olCbE+z
cweL0V7wUVXGzocozCxrkyB069EmIEC+v6W+uMksmWOQIlHUSjJfyTsOfrbfQ4E01kG6omfsyz/H
9jIa4MhdpqpAdYjW1wsT8H9gNqEBWk9YYGbkzFeYv9Kv8QKj3opfp65PGjeZEz1IDTL0VvcrRTXs
p/B8yyKXBDfbaNXPYA++Jo09VVwz1yLo67aXVk74uxV7xW92mib3nGLDeAILQkSEjqCH7IzZr/yB
sRsO4nyxxIWnnwIFHNWVB9YO9gIuHNrx20dCZsN/I6pukvNPhja60yCrh7UMtUQadfhzprabm1L9
oea+pDBskvc1PZVnq2QI6OladtDgLVNKDjfw4Uv32IlUcNrEAskxj3jSQSD/VqdhOD4wt56osOz8
7/0PbYksHfREZ6acgamjkFV0koIV9B4Jxk2ToF/6oNB6toKQyB/u1bgCxHqgyarxJ7umUEKJ6fLn
2EokhMun0x1OsFIamw9RfBZkw9Bh6/0G4ZHqODQDWA7p+GiAhr04WSVQ65nvhoRPEyQivYAYeCB4
I02tOF5JOB7g9v2JZj5KrkNHFQdFtd9s6nh3spMfg+T7OAfDYshsFJPVxDpbsB7P5IsYUc7zKLQC
gOc7nd5kzIrT3UY1UtFvbs8p0sG6QpDPRFWDGO+tApwm2+4qtxsqdMW9OdVfIUMnsPMxp5huTOv7
UCVpmKnVai+0vkl8dAq1CrdxFIv4/1tpPtVjO01gtFQiOnRVS5qjgLAZtkBQT6EiQ16W0O9YZ38E
tWQWzSKpVt73IfYRl3XTbG1JPY0AH3SJQDGcltnc8kCZIyoIf4xhWOfOZQW0QDEoAQ8DcsOrhqLL
a9yfQzjX3tnTIdzhEoxRvUjEtwyeHoSdr8eJZ2GqGYGMvkuQKcyt/2pP+JWo/3Y65t2UjdmgVewg
dnYbV0qiy2j6q9BDHlhGcKiaBOy4sAjU8qkF7vDw2qk4Cl3Ab7CGl4VHF64dMbWQbc/tv3kPFz2Y
q7m8MK0Z1i0MF4XMKI9AiRT3TdjrpJ1kuluA/lPBRKFne2sQQq1pj0YbUfL4v+8WQFbAPUtT1TMs
6SBsftVvYhd2m26D3iT3U5DMo9YNoJqOrSL/jHZJoGwxcQsmqbo5aZMxUBrq9x78yAglXRxu1AbR
Zhvcg9OkljvuT5XlhalIUXLjO+K4YafGU+sgTN+dSrCNeaAyElI=
`protect end_protected

