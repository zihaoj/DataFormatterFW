

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KfHEbzufW5/np0Nq2185GfeO14Hv8fxr1TpOeiVTIxQc8/SA6asj9xEItMxF9eDI6z1E0Zt3my0c
Bq+X3hVMxw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aBpqAz7oWD3l4qfNWJ08PjD00GJgqni2dOD5/3ioPe3LmI4VPwSolvefT6ETYKe7V94NCyacXxOW
f7uofbPqup80Z0H78GX3AgfwMKYeiU1LTOovCbZaHfNoaZdryYUGJp8K/PgWPm4GGJTbBCxUfmiz
+1LeJiOadOMBaQu+Zu0=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O3SFa0MMR/qoHufDh4hPxq7lcm15rhym3L3b3azosCWJTv6sSaZEQgJUCmfSd0PDqru+2qXuswoR
CokYnUVHEDufDsGYZFL6dvuCmFwoq5nTxxGdwJfYEgpDq2h23mRAMdu/q+zc+4XauCq5MZ7x6iIf
2Xu6wbZHwpIq0/upWS6auXfGnVM8TJvHAwfskBEC/6EQQm8AVwhH4rySQEHYasrK0X+qkJtpmEbM
MuRcUjolcAQnpeJZEnpNpg/FbX2dexLKfxMMr/iukYQeo6dt8EiZcS5gXzLBIpXVHRh8HczVZSuL
APFoZP0XWRqOrhjMLlVGv7R+Rh98ZvtvKhIvFA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GdLafu8nof1y8qFMZ3bUE3/pmLxtqJkWwjMujEriRCEjVHEM37RlkTLEu0zpaoB3nLmNzJ/nPndQ
enllEIh1KXiDCsv0gIrQrNY6f94eHJDX2ESlUZN+2dfdlcjFBZSl/G1nKX3lmci7nGl18wBrO373
osWpw1v5fzyKEYtCEVw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DSEh5EmapiPqeNY0fW26gkfqG1L7JQiUGHKeBSEbiGF6Ulm/EB/K7ePgd0V+sutDnIv+dg3PZV9t
uaPS1kfu7ghAjIOKVpzNQQn7LfUw7izohcL0MLTgj+49hsu/ytcZrMX2AWvJjwszyS2SykZKPJ9t
oRAmU616JZCWLVs4+CZwo8AHP7lu396ZJLFh474FXnFp20YU5LYZUqV/WLkhcVUGBJrzWFGlXQRs
771M5nv5X8TmBP52Hl6rvoDa8nqerL191eQosoDYkFPK9VcCYjSeccAewAKqJ4tpcDAP7+NKQrO9
d5CM/sd+TZhG2xnBsz8pBaE2U+eNqT2LVeERvg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9904)
`protect data_block
ymist39KasajaSh+yy4xobjBiFZoMFbp1o/iGpJ2OgYYupp4l6fb/O2HsAgIotjFowhOMkMqMFWv
OB6wWGAouk6XsnBF24YC7dP2FXYoGXTVRHYh4L+s5SGuurka1sB02w20gi4U8fAsUp1VI4DL80xP
4K0UNWgIyLMavGleDsovHXId5MqEFX4t2dUOziHgtOsdar5/FaiQM1eeoZRrkG65yY8SNZk88qRH
QxKWgEs1qtqOWHWaNGjIa3kZMEjBQIcUJ3U0SXQzXuzXbzijTI0QSenHfkjoNhCpezmabupNI8ds
nD9jDm3+e0+RdvN9IuBz2+HnrxMdEUapdUxZ47jy3tYZ1+2M1HilGqYU7nv5WpNjcKLY0HzNgne2
fCBLNUvUI6Wgl6I0Xzfl6Em9hVQH5iTlaw4XgDwLM/05jxyVwB3a9EGnmGxtPCTIN3EsgS6XRGMs
7MBMzZrGXFYzXr8rL8cODB0uEt3nNyqtgBZlZKFL7S9c/sbku7iVK/xQexksJi/pEHKWRgGUpkow
NGii2SxVMTqh18B6TnyZi3OwZ+X6Uwx2Re3RStRVmGQLWitFhbpIIg2bSA/0/sCianoj9v/sKhSr
b9+fyQyD3NjZCl7e5ZNyxhkD9H5hqjk1JIy8Oi5fz3FdHP1vepCGuUcFLweUA/K5UK5nAHLBORrn
yiVJMI/naIgap+Z9feHITUBFKStze581ngPaXp2OpcZwhCa1toSZbg7qWxItOs9UNEtLLsc4+ccm
XQD3w5VM9SdUAsNJ4lnqCePU3zbl7ut/bOX7+BJehOqZ2f+9n2FE0Eb2sGRwP19pAb5tog9oXzsJ
s9U0ptXjT4IffYWkAiisobmE7dm/+EOY5dp9JhP34YLEFL8yVNWK0Fq0zEz8a2oswGsdvaORc0bR
tnQdMQoCefeMxzjccamIYAGDNigwkbRqsS29XXvHZCdoAiSit+dWyaFh2dDvs/brExLVci0N9h85
ykVKMJzlrrljGYci9dBEUE0I+Zbzm49q7vFbGmzwqt1p60dNcYZwkGdrlGVYCleqd+zOi/4AAF4s
f8+itPldHHPEBv/pckhrhEPeL6VDswZV5h2qvbZZRvdy/Lv+dU8BKL6lburtIRZMTS59OAxsPKqk
QMxdufnAHAEV1QrEXMI5f3z3RIy27CfHwmvOtIjF8CFNI9+suPJ2bYhXJOZwXCzJWo9UyleF9zvF
iKHrTyb0oXxijiKwsJxVsTZHNOqeim5bYvMSnQIEof4JGbDqh7zuiRX6uXIdlYeSx54XDUbmkfRj
qXDhhgdaZKkxkFvPLKa+Rp7lAkud+mpMREgheWL46IDh4ouzNWOPDKvvU3DLDlH6lt38CWE5TVIT
ghnRLhhfkJPSGCuPPtHAP08RCmWSa5zTPHq1dnmnIVBywam3zOxP0Pb53cRWFi+jkOayBXEMLCfp
rOm5P81C6yzsPsa5MLywr/XuwQAxfU1dOFisHP+MOe4YuAbsJ1O7vKtPneWFr6Z3uO01EC/l8aiY
iA1GBE74sDCtvHltkpJ8p12d0QGeyXr5xKo3PeIaJYO1in8swjjau3HtWxwz1K3d6If5OR6Arc5/
l6b9Oplz3OTpFzURuJcoN+JwmZbI8PicPua4WquBf6AElv+JkxVNkgfQXG+oiWT1fB29asBvY+Zh
wj8MzYGbhbZRUQaSD1uSoQGyEG3YSxBvRg5Is2AVYLk9J9PYXBQsuNWBMm3twvKjhDat5MrD/O5c
u3jJHVdDANZWyZo+DWGYOlZbkjRrs4qH0fxlUQStJEBXJBvoV1hQE+v1TzxW/kof6araKFGK2Hbf
q8Vof2vVJyC6k6mypmTaP8EKwHxvU2ek8cwzQn+Fly8FENoSnx2aegU4Jo9uo8/OgoFtD4tlDYNd
ZnI3Ld0vIZfZ7wAqrBl88o7UhG3wy1Oe8+0er0cuhp9UqU2iJVw8sSvQVWECdoa8OedFg8D0P92G
OblAkGwKHzxBCmeJlC/1+384azw8vjbDUsmnBI68gAG6A5BWBWsYTcsbG5PSelMLDpB2qS4tmah7
iMkNgunmmxH+qiquiVVm09A7PDIqn//oUML2Q57ijhZ/a/mWjSd8TxiVw+40sSgqb9WWXtlneRu+
wtA9EbtBBmn4rT5GGeTURaOW7Gn5cw8GjWupA1MNYdwvff7T2HgOFTiIquMD5/ECoy00t6+8ugci
yfn/N7wfv6N/U/wGaEIZLHCy+PsaAcH+IRdUw4qeOixeKc02yFo82Yw++QjE4fVX+Nk51BpIs0f4
pCCNz0Vv+Q9NUXmhJIRNmgbUy/Pow+hrmZbweWIXD0NC0YY2RlZ8a9ssI6+mT1FjAka4/4WkAf++
JnzE80eSXN4KNvj8LqMpUFZzOC0qTpX6ga2B72PEhSZ7I7y9ElOFT14ue5+JJ8SUhJIYKNUUm+m0
2vRxr8j6IAIhAcxrdm5ybcGI7LXY96rmpkyBDoCZanvcJqjpCSWAM5O627/b4PA+LUbshSoF5AWm
s2C0deYNeEbhk9v9UjtjDRJehL66eqwC5jecxdmnrw/oOQP2J/F6+b5QOWBYgL7F9nf0+suaSMrO
/jeotzhuktJMjXmeiwbNu8GKq+/yecBvLOkoHnG3AJJ73PDb8pMbloHKXosIT1iafKbhFxlwtmwK
dFKsbkHbp9z37AoKUhExHEg48wSrLZDutk2Wb0fbui2f23S7gGYFxbeRn9WFtyn2keOfObYVMOOd
BWDDm9vdpnHO56DTfatyl9TvsNlfy/rBFUmiIAlEOB7w9moI6qtuMCdCC+5BIzGfpa5zaYtt8pMX
/baom5Ma25hrbhosaU13tqgy94qhE2q7NPK8VVSvuH160ivijFi5zWAtju2LHnL65fjfzgaJygoi
UnRRZdWeAiIKhwfZUepirpDyjwHFss6tr0lQHYCujbY6h6aWyjS/ZfFc+8qcbQCuMJoMBtwzFD9a
V7AGkSA6bHNGLiqSuGVjjwIZ+1mHZYfZkLo4SFwSZcCdB9kq5XbB1D8eA7iS+wMLtOi6efuaMLJl
Rbg67O0t0jRrUcjXP6or6XQNmH/WVV7Dj+j8t1v5a066a5CxULRkEN3WryrhegePnl4/BpuK2X4g
pBFOvs6XZp73muxqJ4M1q3cjUAnFngU17zkg5kz/aWOF7G23W6B9Arf62zktlTgKwzN4/wogp6bS
1YATBNGbgmOPHnoQxIM9QfwUmhPvTZcrIyN2lGzzbJBMZzjtgWUElEiUOR6wRYHuwewOiTlM3zzB
SLrNRDc3+6g7xCNMYODSDnst+PzXwlqOXmye20l+HMYhYpWPDbJ3EyAj9hBBIl+cXO8Tfgems0/I
4MU1ByVk4UyIZGcslKWkFsmp5dFPb6ClCl9RjgusGsqax+VEHjGtxaydLFbshCUDMc+t0VMA4Xtm
cznKKlAovLMn8kRLu+dYihkvQ9NRiaaxzPhUdtk+D2Y74T/4Lc4iNRFQxEztzGDiCnW6uEhEhagc
HpeJ2K1uhuww1vemhvID1In60w02dOAKJCd7urfS/kLy1CCV51W0PUezQCTd+5rcRWYV1x8zflXf
CfZ9sREIaCQtywOLCmlMmQivXyryqGC6kuH1AEIa2Dj7AbbysvtS8dp4SaFb3foPtXNPD1R5tZ5w
MYAkVtZ/cUzvw+VWZsrjz30qqyrLp0NABPEpCavYbzVolO1tsTSD58WElbGPaS1PQbBL7hSKw3ZL
pBg13kmik7NYVp+scmyz4ijW8e8dlzzADl6ISqDlSjsE7vrTJ01XhlxeGm1VlhVciQHL4BdwVDum
TTwLK6RoUyktJHBlCUD2iT04Rk/2u+4i6wY2ulOAiYSaekXTKIuka748KXJyRani1rDs/Dw/eVif
gZZcZMAD14HF6xheP/midzUagR8l+rPEjQKSqfomDDgW8CHXuCE9V9csqa3HAv4QMROkqc4MgDvx
7nGNoRXoDlmXgexU9corSpahAivyk1bOfGnJRp5yhM01Dqoq9ViXU2mMoCBKA/XTyTLdsHzgMz6P
gDQLX51FmzagKh9le7OlMOkzagnVg/RRKsDVf57BnblDw9DSsSbQYcVpOQMfNom/fLnhQrFWKTs9
Fx29N5//8ssdHPgf/kHadFXPzrG3GGEivS2KqPpbOJrphX9FmDseEoqgdIvZu+u3e6wxlubEs/qu
4nwmXB+ryvN0XsToAkU6cPu9UdnKlrPb04kxilJkygm7+cbToEgyc8VKzAWwG4aIri+MttbAH/dO
98DZ0VB9pZTU+AZGQT4QW985CNuEOvOcTGYbPeOc4AQZVBY+lJbgpaX2OBBt36HELTldOKIcV6YB
SocqDXhlZXIvB+85/aZIVOk+d6dr/5902DL8KtCB+AYg5RhKPtNroufnPuH3Kq5UNcDHAs4K578l
N1lBz9ljSd/KkWBwnvVBp/1dksYL5uW7h8JQKrumxChkAcpv8E4ctRtptAsBpaE3HhYUPre3ValK
4LS3IyX+C/Obsg9YkS4Drd6W3Hf7Y4TJawE6MwVLAULVDVTn9+/hpE7kbuAvWw/r46DKRmvoxP5g
RrXBbFr6puAkDNiVIL+iCHoi2i5baKW0Wps7TqBVrlWarOwgn2X3m3kpt4xN1rNDKOVDmPhGyfxo
UTvyUIitaHnQALJgVclI2QV5N9D0lsBX9HyB5RG8VJ2srA6gov+zWa7CV4iJ7zuZravPgZqioiTk
iUEJSoq+HKBCoPKcggOH/Q5i/U4MfJCHwO+xujohJZNY0MKeJ09KH8+3tu0ud/4btMRGqM553RVX
TSMY421YjY3zmAi82XGJKw5e5EM/l/v3FOgWGMp/JdeFjgY1te0VAiiAC7ReLsWltySOHul1HTxJ
Uga1ShPwJ/zpeYZgv26dEY4glvh1GTuaFWDoDSW1Wfy74SDL8F7F5487fRtM6bbLM2pCjN5xZCSi
fikK99LNJz4wB/Zlm8MokwS8eD2/9+go6raJBYzp/IDFT8XOwRddzty77fgaFObowgBLgBGA4O+s
tu2LRxWtEMoYD/aVCFWCvsMTI9xh1RytWUScGijbEYLJmdg4iuhufU6goRo8Jsq59FNVGD7J6K5Q
OhP013wbjFAaR/b7ljPhjUMkCafO4r2wJsRHZd3K76Vqx4farSVZo/buiIJ6KD8pBmXfCkgjpbJ+
RS0CeoHNIZVoR74HAy5fbdfUfB1ppsT3+KdEmI3daj1hTswPettrFiucUOtJmEXNLYyRo44q52eY
bAmXq+9lCu7whjFVQfs9Glewa/lOVIVGiV9le2RLeFfh9XuDCPmAQIshYIiwwyEK4piiLMew3wld
ojyUs4V/SIIC8ksBiijmcCVVwBEyCoKtZbYKmNWQXDXXKJRrtjlj9293ELY0c2Wci5X1pnhdezf/
rxMOl4uOMC5aQqU8fk6wgAaA7ESerONVkAn7HS6/tLWWBq8NURXsEw0lO8IVQbheED4pVnTd8BWf
VcCH+bCi4lIFML5kYo+u/bW8XP1l3wTc9FNBunFVXvAdLZWidj6DBnjMJJWDiVLj7nVwPyt0dQtO
7WGZ+j1YBbGIAPaOGTrJpwmgcm2bxeXOHF1l0Xv5StmoIfoGdnZU04pAJ7XL80U+ToKMmzx5XnKP
tWn2ChK0tjfqxoVkmzWnByCJM6hOgN+r54wHDqYGpo7cRkgb96P+7mDKiYNkF2I18a+tDTMeBMOQ
V9/j4N7x4aBz7C0q2aP9zUXejyvF97hbRbxRNdylp7XMBciuD7//R494r0/VamjhikoccTKU9Emt
dHI/H8FuYgiMuF2IjXlWoq1EeQkbT8YfwcuHWLa4P716Bcdzp+v9R8l10ABOOXa+cPtmY20dY/Y/
5kQB305KJfwHVlYLh5Xd3aaO2McBIC90EIEsBbUtx5Co5Sa8XRvLKqPze3hnYM+whvixYU7tBIdD
A/8DaIFuruLjPWQ/mHvL1ExXUGco5ZP/yN6oXznu7AQB8gOHUOmqJpjcznkdyTQusHGAPOz7Ilrb
AOlMYFKC+UxGfJS20fTrP6SXv37vQL7WThR4IbQTpIx2b6TsKiqn8T4lQVOdqpxPrHNnQmndV8Q0
B8cgyvxIik/x7X8HZSb5+wXCT2J4QvE8s5stZXF+C8+6KKtr2p7b62No3l4Mf59rEIjXFmUKUVvk
+G96dYnz6Gw1JklWK36etXbZLch9es5UaxymLJEFsDtix5ouPTMvV267KLwWogvuaOYYPoFWC0ef
X2qGZvJ60QTpAv5528ipwl7RSkLAenhpHaMsf/5AU+wTLAjB11Si8iDZ6YhZyf9ll9y/rndgBb1y
uu90V+C0z/xzy5Qx2lQcnKW6Sspd72dcIgq4Enx0/NdS8rZSb8+muUzzlxRgW7a9c2PiBH3YNDbo
HH0WfSTwBs9HRwPzwuSFpPuAdQCl78r+UgxT422JZdjZ9GhSXnrV37q7SuegdUdpCr8C5Wn3MFg6
tp4vL+CphOkE5W9+n4X4ykTcG+WzjHoBcfQUJKJQrVp3IfLgbwOLV0rePfl5jF2dc8UKtFSDTIAy
lTMjvfZLlCTqldd+w4+Xz6cl6UHqx/ht733nxHR6ad1+BwogAzTWQXrkVEyD98qjEH2j5+tzrCaT
3FlHjOAhY0Z/38DLMeFlzwrNGYx8NVqp7LXjQjLypD3tV97y6shVtOXMlgGn1dUO7E0/Kzq971A7
ROkkiGCsvrNxyLhkytlVZrEUa6nYTkJFHop+8iFZ16+lyFvgNP06/cvncp/l4qUi3GFdCZniD2Qv
m/eyotC7gXZkPfZ9CHh36kY3Y54XyKy30VQ7mueBqxOaTMJymVwmBFT9tmZbLTeovfwZHJfucMGB
6bNOUCEBb69stFxq3Y14cyIPypHQn921o+hisY4ZDvRcGaUnxq4AA1cXcerQLGLyLo+F6T2Dw8WJ
39lPBDliXT5nyUiZwEefc82RnPh9v5zK2EjZiT/kLv926gvDMmmS0xlD2zEIB+HsuXEYbRZk3kq3
7rCD2dHhHE62vaPrc3PJz6qTCvILb3pdD1np53uxxCh7p3pe99zXe4W7Wji6OBGD0mNVPmUENJe0
9kB9VOywaT/G7XbAiVg3sib0HmGtJ4DguoTa3EvGh2aHoi8M9IsNLhiQ7eWyN9YiR0rLXuK5qTgI
3aamuV5ECv/WvvbO+j51qUlsiuPF1exj7EWF47JjWwqGhVZUmk32fA8/9DeXQyKwlIt6bjkRhXDE
LFCd4eb+uezAMLOMlCO7pSmrY0lN0+c1Kxtvd4Yg+LBIHjpM4Zknx/1dcAQ6yRiau8DN9gb97Qa9
l2ShF7KQMrXiOWwisrvnPIgmY+jCQLhULQ6mwgAX7mm4aomKirACK/Mo47tCJGJ3yb3Y7HuIlQjq
olnGUUi7M2YTwqFCDF4PeOtErwk+olzn1Gob2WaXJ4ZboJUu+3o5MDnYgg0kun8AwnOpu1N4r+lz
qhKi9qoZXuVmWVVlPUypVA8LkoWiY+EybglPHZu9Rm2cbkEdTTSyWfQVoLacVyJ0K7bH4O+jzaAq
fvoaQye/Mk4LFWW33hxYDgTL+4uq5T445u2REX+HF4FChlaTq5olPAh7HofrOHOJzhrcM5c1ce+D
bpz/PAdzXuAG/SIA9N52nu9V/YCGq5C8COj5R+r8TPK91HylvmEOe5qtm5gBoWgSK0tKJIs/OpN4
9CN6WD6auMxOk/flq2ZSgKuXJM5zwE941WJ95iZIDIcwpI4VdnWhgEIRmPLH2rf5ZcfGK6d6baIU
cxJkzWsZ/dVRtJByc3mOnX5XSGRyzEpCwPXUaTjdWNot7PqCJ0bfVy6ERs5/d/sy9pwaqaag94kK
ak++MDH/GbRng9NX7+2K5LoaNT+VJ0ZeSCXtU+8Yblcd1/hquigpngKWW2mWMvu91/qqrdntbj1B
irVt9xQQ2umNUA+KOjLcAdMoyFkMHNnuIAFxzHJvBLeIdYx/q4lwUuymiadB9wzr/OCwwigup82C
bJuatoErobx2TxhUOH6ivNYoWKUKhxByEu6guZ0HjhygAt3VR3nbzshASn/C0oqDWZ+VIf0AtVav
gPrU14usZnYBxkmq2YVA8ZX29bqtS5cvUpQhc0nhXDhg6Cg+UwVgjGzBfYinUunJNn3yQDSKWt+I
O+pSgbPN6v1jAHJYPRomJop5cLXZcGwL5kXPBK9zxuYT8yAmA8wKajAPu5uUDiGOIOsOvZn5yIz/
bLhg4zCzGE9HRx8MZPEY2aG2cOxM2bmvrULUuV4I47+i26EGcHejhxsgrYixiRgA+5BtGow5BnPx
ncsqtaZfPkPQ+63SN7R5X4lPiVNW+Btie/qOzC5XytfE+kdBEttKvTJxDWwa7BsAHypoAFh6DBKa
6BH4gK9qyuluzMHsYCR/dNAkeyngGtQZzx1u3e6zbkZ+81yyfXvWJn9N777Mdb30zlrFwJ1tX5pt
T9eG9XwRJSSG63ho3fqft35CSYcmq/91GJKO6n9jg0LtgsQK7PusGGEWN8UysHKPR5h93c/Kl3rL
DtK2V/cKU8wx94tkiulkKrlIuA3R13+ZDXCxAuR//UY/M8Pa1AnKnfjwyo5oyxyKSPvQtqVwMvUa
IMM5vI/Bz38Fw2iDpoVyPEA1PxjvX8U/Va4I3tnmfoZUGWfhErZK/aaUFwkN1tKFDCIyX48WK9hQ
IeeHP3eBM9VoJ65+t0Wtz13Ms/8jq1c5nsFGuSynUcf3pUsqFt11UeROgj9JBIAE3aQGjF9wzRkS
DmX8iQCSLz8CkFTNnmZjkqVx74GlakTZtzqxevZsgLH120xRXgWq3k08QNT9JYJPyxMxKTu/xuTL
q3ubsjmIjerLgpAjY6EcjZemR9DPYOSEyiqlPQjJrNbe2aQeox9qefmOKraBI3nSXapVbYKFvSU0
C2s2/f373d+Fe+K3kVgyIxfw/h+osvBnDnN661uiANLq+giWtAa8nnyRSU+suQ/ePZ6Ja5nxFG5K
UF4CpauYURDQR4vI70zMwKGqmsSeRy7XGzqyMf73Q0ngWEYMnfvWgY9Fb0Z78Ah1uQCct6fTLth2
pJAg/Of/TYH6ktG+OvR66f0rVqRcS9acOPbVoh6TF2aePXHfSCj4uPJc5gGOgCAVW+Cob6T3VvJy
x/yWEo2d7qJt3Pno6dwE1OcDi0x4hET8a536hPTfzYR9PpYX/TH8bBwbykEhyCkH3g/Xs/uJjyYU
cObcx5faxiNU2VSW0Rss4f8DplF1ZtHJou0TCWmrzYS5XUjrHONbWtUUVnWbxy0NQWftgPh/QOmj
Rsv9M+PHf8HAgjMrs3qN2AAVMXd9UBC+lfChNo99lGY7XmymtNUoABvAKUqieQBAgs10w1Io4huI
0XgHhaAcdLDXUFTG8ESQUA00wqdvzFOVMcIqRlnqqCSela8eBlWb7O8imfHOVIw0LFP+J2pwiL+e
LhKQMMJQKwIz4Az9sjxBtdqmuvmfOxawxZ/cdE0AskwZr/77dEJBv59UU6vmu0axVZ5hR4Vxc1mx
iF6TtIj+KjbPfKASUkAm7Tlzxh3gP3yADn7Yu6Uyh8F/KAuZfpYAdeIDvHB/GaDMjAdEgBcixDrG
vCr7rWXksKhlZzR3GNk5EwcE4Pdhs3Q6K8NqB+L44SBvGPi3pnRCoHcSfcckF80fy3r9RT1lsp0S
zmvmXfvg48fCwJZrsIKHGhY+1lb3r684Rei3B+5R+FocRvYbmU0X68qy8ATUqy4aD0d4sP+LGKds
wUTyxW9Mno2KFRU25FDknUXBGSVSkYFrcVAJLxZriW4qL2tjRJoAvFxLszz2y7yKTpB/2u3MxTsC
jxReyu+8Sv8an8o2H2HN40yriexCs67eI0hV3jiJjXISMoVZ2nFBhFCOjx88sK+kXkbf11zsvxhd
duZca//BSwBkIzX5kBRN9rNABqHPalhgo80n0uFdeZra+lHT0cr6GoKwnudgaDOHIV97DcoAsoJv
wtMPWxqhVP3AR36olTCoEwo6r1CumNUEGFqViaOayx6gkRdd1+/9Oqx4JWMODJybTAqN9tF1guZ7
jckmPRhXU6pR7SU3dg+iUa5f4gR7XeilYAfCDxE7ztBZuVi2HfOV0r1m2NAUA5Fc8i6NjPpvCFec
BNByIEa/ZiGw/dJa5lV7DxPXxCkXpSyuKr//shOYjzSfGZ0gQdJAD9/iLFwbbZV+kiaWMQXyeYbe
JUPp6GjvJdcNdky/p7/GXMLYEPCczyHsyVux2pTM1ssemIIWfKxQTeAzTnIoRwla1bFJoEArtoIZ
PefcZ65rDKMUX/pk5I1+Xtmsr9L1sksFWQ59MhvRCzHJ8VNi0gw3Gf8fQmT3gYtejBMdVNlmRQaH
P2AUIh3mh0zkJa3K6KZ68uiU+mqDO39V2ztJxR5AV0pHoexe4VQX1fcZD4U87csEzYKldYvj0w3k
gjv9VJHwBLr+E0eqaB6d0PV/NGXvw2M4Mz9XQZjKj5LwqSkPagfA+oz8Ldq3ahSF1bToJgEBHia4
LAyBvS6MQxGbJYqdmiPovbdz3auqOWA0SFIghU46J2NK43eCOBn2rWvl34eFE7fi94K1hGnn8aHu
MIXqoVFDkIpCRhm5EetML32V9Inhq3EOIw9lLKXw/C0X37Z4dm8uCVbJljgCGjwelTF6fgEv1hSo
iUAn0PPXqmnbqVrx14rwpa3Zc6ILhaK86V3YSFHyQgiHJGBtaBGJuxle+PYcrZQudMt3YeiO1zdZ
uC/IVqw5NHgzXblyJVsZH+by3GtMKrBUjyGZDwzUTBftrX7enxeF0Nwc07sHnLRQ5vEqlvpKKujH
NHuQ2BcHQy85EZNkC6ELs7yqoD+N86k4wKtImBC8Y+lfFooqEorz4BimbE6sat5RfJkfdE14PcUO
qH4leXH3Nq8CEY0l8R+XnHy+Pn2D21X5d2zwCjAmjp/ufN/eFPPFCUiHYKlow0cu1r5Jc73T8ivt
4Iw9Og1TAGF3cK+CaOVL3Iw4w9upOp0DTNk3Nv+ls/p1zYrUcvQL6Is1sPq9Ap54eGDOLGJ2Sfsb
OORb2d6hu6ldS/fzITWgFl31Wwp6YTTQ2k++ClGjpOhDZJFf9M6mKJwbxl7Hz8LJpeAf0hMU8ms2
VctGQNX4u6yx03vinGu8HQWNyQ5/WwXgvQ6io9QiH6VUrKpuOPZbB6uyt3D3kHbqkSOolD4Q4Cgo
+5FUXltJIshTP+bgI8XK8eYF2U9RFHeGvElJo93p/TiiPAI4PMBuQvmJlR2+CG8Qdmj24scEmO+F
i0RAzAbXIJigX2CghP7Hi09Pgj8Mkotmwl9miSDLGWABTdjgwzbSU4nbNRiJ2N8J74H7BqEhlvX/
+MbDRAiEeDzJOn0s4euMd1nMePm5EKnINfeGAIUhshkjcijvSD0fLSygK4Xj+j532Is8o7E+9nHn
UpkRDtWmxZUfoGuEDONUun2zUrv6sYwrq7FKARmU7Kdl8MVni5ay6fuqrzYji0WPR4ZWEBzQ98TI
kiawny4AOCq51rBZfgQCXgGH/7nAhoukoKJNI3AehTVymBX0DOfd+zMd2MvrFNIIxjhAp4TbKk1E
YOnpFE32IDZVXbBpdOA9SFlp9HMauEoTUydMTSdf9EvDtc4LMBK3yWe06xYRGhxW8jZVYxwx/b/9
FS1yo8s6Ph1Xcia9AHNxMqQjEBQK7YnA/L1zR9+hfJugepUiIicRG1+7F1mVZoQLWk4qzwlzSQVo
5pRiQ8FJ+mA9inqY7mn5XQUCr/jB0IOV0Y6bFUg/TafKG0LbQkM+py2Sq9n+p9ZAUDfcccoT99qz
iatVUT60rKAKCjEwpt+2nrUtatrotR7B4V1vQSWKwNPivr1Er81v6RwnvqvnT/JDZUE8NCmBk30H
BDSr5Wref941a05311TiWUubFDSgWZaSwN4bKZc2l0uz8urJzaZZ9wu3eggQRXEjo0JvzpeQ/rIm
bGYqHyURLZGrhyolyYbSkmehoPQpp+HPiFccbXbxUs/k/ypViBfFwrWgPLwrjnTrVnu47+WVjd1z
6y3vId026ZvQ1lR4Ip+XVV+GuhdCyJB8VIqK0+yMK5hihCJsG/jYDOdgLvR4aiXFh63g7gp8T+xc
D/kQfe2WK8Ao7O9UOyhC69NZf2eWEBOb+5rRZiotv9a59M3Fj2e+EuCUsU5x0L/GrZP2ZF1eyhlq
O0Q4UHDZQlXQE81FWVeI5jzCT80Be634wTwpTo40Hu91TjYe8hpEQT7/SdujrCHU97jXZWH9Ksla
2gjNavs93PeUiKyEdoievNgNZWto5eFREBsQNbco+YDLghUPoEFtl5NsasCXyeSHwiduA5k6Tx/J
WHakqnN7oQm8CEp7uHA/4pAbATcmqhONcfzM3P95x3GcTT0CbwtrV5QrSsQlSS2VWvqeZBU9SpSZ
dC2674eJ74j0chCP/YUZrKDwb+g7UVUgaqH1g+L6V/kAU1pIXvYcCvZjzRwa+OwAOU+A6TOI1WNA
6AjCeNKv0PsSeGdlO7OCgDgvOgvW6V8qHAqQfNKYgkyy2Q6eRjv5cfamtiUTn4hnCfOtCPbBw7gm
BKjoHYuSjyCClgUo4IxsjnGiDUpAqd2CbHLryeu5Pwx0P+514mKWAB7gjpZrY4axeL5e7xXPfXWw
nt4Vg49rzEa/IAYGh9mdBjixtRCGkrc6ZLHRvou7g1/nLmlUt66qpolKwvyG36T+U4SgooqA1ejj
52VRwT3maAt6KcdlWVloRTNmLDfk6qMyQmY5XKPCjKNK/ZVwmstUbZbAIACcMd0jCp4Ba23ph4r4
fR7NPhINsCk/WbukTtkbQ9crOgu469Chd9O21qViTnOhTTJXJbh/d8cwQ0QMW9kGD616btADIZx2
GOSSOuBESIbQG8OVzD4OEnGsNrE5jQs9x3PMag6z4+cCtol4hneT/HQ925sNYZp/SsFRtVsIW6wq
Ulp7yU8o42CW3CscWofIH9oTpvbxxBuwgE8TKt1TeZGU7oO6mcy6yJrd2MYDbjhYX0rcmBv6luin
gJH0kWmXyomT3T2B0IaGiRk90ywbfdSDfD0kDMrfT0osvVAArC3/3YhKjyUOVAvJ+FRFDjXXZ7+N
YMrVADa7Mdp8/XVB5JlTIwLPxL25/GRVAcw0OVb4UKw6Quovkjpelz+NJLmQAzOeA8Fh9d+DfUdj
w/W+Hf1K2x8fUR5UkEi+8tk3pCeC8pGUXimw8+SMUG3aKOGSIj1IPcPdvQ==
`protect end_protected

