

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nvOgv7ZCjWXhLig0DqIYarjRIYNMgvBL4t+RjnW9dPwbE+2Dmh32daQC+cRejtTj4d/pTHalxJ1U
DXmEK3skRQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
e0ToDGmlBj6NVat0a3pVKyDwHKrzEA+UGHgXhK7OQgn7UuBvEGNAv8O1095qSG6Z7Ap4nUxIQGWO
HN8W9LyttSuXrYZwxN94RSwh8LTpJbvnyIYi7UKCvxXR5Oy5cXr7TEPpgeaKovipUGiYLgfC2CNR
3uJz/3+qMM7torm2K8Y=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Fv7qg58PT8m+ynJ9+MpU/vfVq9t6OiKELULZ8eRfbgNQi0mKRfhO0U6zpHfAktl8i6biNbgdxqUE
lewPF3GZGKzH2NZ5CAy46Ey6BU2Uu1o6ZRPZPAz5O1c4YAafngpK9GxjijwiWyDRgJqYlLhfos+1
TthFnUdpgqsAoQ9NtD2kMZTv4trJ39rcXB5r8eqdA3/HjWFo55/0e1t7me6QYGbO9o4j02WCJ/2Y
CqdYVsXDTWfDKKuct8YE/4EnDinZv5ViFX2jT2xSj6HRofzKZ8wBHZo1qFMDOMZPAHxGBF4o16OB
G6fknQ749sUZkcDpaNI6KqkBUxthfVzLwlR7JQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vFoT66pkN2So8U11U09GK3GCMg3zGvtB6aww0ejFwkp+kCApkz1FUtfoW+7OurvLGha1nuizzFy6
JHqpRCC//bR/aAL59rW5bZvtLumUP/OfHLcpog4o2Jkknfgi/m4keolMa5f8rve6bl1KHM+P7zCq
lswSgclYJiDaxrvBzjQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WmbUOreOtpRj/pbzJmDDVseOMTkM2iF7LTkKx4RCEXFMloMUOexcSsWaJjsuaCTUV4RlVxayjIKC
1Eu+tpQLZ3yTZLmqyMw3/94wD5Zc3P/Wung6Wut7iaMBcAD30CTI2i9yGrWoZvfm50+oD0lVDIey
yaJ7Rys9XXn3JxgaPWzVNJcXcFQajItPukj+WhvVOIdv39b3EBSWI9tNjZPLBLn8ije+c8Wgd8cu
KSmWLEix0GbbgKyTg3tTJ/hLjsymY8YrqsGzog9pkhMkWi5q+ZzJ0CzxzWzOn+s4HOFte+NKmRdv
yRVnpdnX0oQ28bUB6dG/ePjWYdVfyAokL+Hm1w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62128)
`protect data_block
D7Mool5YcSgEzQSh0BBfhAB+7Q6MIcB8ZQ4QEvxFvuyTQ9cVgFvKStTG8hSUaItSQ78jydBBh031
j/tnBQ3b9DWHnAosEP9mqW6V3XnfqgImqODDRGuR+3tPXpTaGX8Qd+UZAHqtimjSASGdLOsi2PQ1
F6JiacCCNCVKDS/viaL/GuccSICvgg97e3N6H3juGlKKM6qtnFCGHIWjohWIc+R0pEBG3nbXlmAp
NSfK7XPRqGw9veLrz3EeI4bwbp5P3kLgUtouHvX35KwPuFApK7f8LsRyWEU1McZnPelU+TcFlZf/
Tp93LF9kHi+blu6pDJkoaZu80evV+EnV4s48NYJtNdbdB0rBN40+IenIEq6W+kdI9OxJp5vaEkBp
p7NLyGXHZfO1nS8psGNstO0D4UL5OqanXdpN5Y4xJ1o5XdIg/38jyWHjWfiZe6Sv+t6f95tcJh4F
Il/0tqXKhmRneh3PJGHKurHBRbUGUu7JKIhFjr65OKN2Co87Qq+EhwyBP/OsMUdmBhL6fN9AOzpx
8CHE8VlcuHT9GtiZDqWftg1oC1d9j0XOAMzskarCXRf5h5S2sCgKIJTNo0EbIix8fsVDKr9Y6sPn
nKQqPBVH0olNckBYAEfKOKtJRDhKt1hzjmdGZnNNrzYRC0vavQO6uQ8FYneZciwSwocGiRf0lQA0
LTCmJjYQonFtAPa5noj2e5pSMSfyVsJyEfbm+/AzSj6NKVSw8h9+KiwNfxIkO+BDdrATwXPMbAAg
ffI9wWDqUFgQWOcF70NhnE1gQ6Jm655t840JQ71/5Bym4aThrn5NXfAQxwr8MB5Ah5fGz1NoXhAN
CL76FWzSMsywrI0T4iczqWiLVOcjtFYk8/bDBmhHrULLmt4EWwfALym9WwGO8ops5FrIqG0/APs8
rpm7HI3Ur5snKuKkFDhVe63UKApAMwT1dCyRgRN6h6eW8HZ9fjhlcB+twyFv+mmu9xGL1siRKti3
qLFEaOfh8E3RPxZZ0kEujOBgdp7ETeqQFUnq7qZp50hmg1nuLaAI9l3tTlyUoB5kLM9oy3EuGM3M
J/gZNUjV/KZlb1ru1xYQbXrscu/5RgqsCMN3hPj4qleYD07oUFP6HqjzTnacsAc/L3x3LXYjt8RS
TD8pOeJ0JnL4xfhStqnL2Fh0TFJRFc2D5VLj7lvhCrB5SGH+o2/LSTHcreByYzWx9RQX2STIbv65
xkb/B747JT5ZWo0I7TsMh4Am/Y3p4FOdXnYadwIp0t9sVFmN/QJNNskQ6FYLWeRFIisv4dWCQBN3
kcFW4yyABrHtvodmAuZtudkqDd1raU689YYGU6OP0K0tGj/9yGAzcQFnb66pPZcn0ChHNJE6mTn6
EjR8flIIfdu2J7iCToMX8SZcfB5oMQCQEPp48LoftItXWRoLnU48iklzh66X3ZBv/1PHLig2Y8mj
3p+RipH+X5IdowkT+DGVR46wroA8N8a7Oq663fAtncMIzkH1FKSWWVCTdyKvL9i/O/wrkYXDoeNw
rOgXWM9Ox+oEZjokUWBFysW9B1IIWpoT7rOx1/Cduj3e9pOIewVGiv8icro4+X4V7dnLpYYeDUMS
Q4O0Rkn8PI5c1HUkmyS7yGZZCAoUbj/i0OY3hLDIgzr6w+sutSwqkDuqQT7+tggBjJQ94u/rUe2E
ib537ZcbRyqNWk/xmQz1UKZzdeOLYLgl+YdK241wNoheYsOmA7SBkR63o4v2u8t9c5EpX+6Bv75y
Z+Vyn/b9ddyT8hxDaWY4OAa0BFhTHwvYdWL03iXa0SOITVF0ICz3nwH/6D6vKIXE1DE7TD+wsuBd
89AMXakDsA+O+3/oeqo8Jnd3foIP+NH9+7DpjbGINCX/HJxZRnKGmank5peImiJUH1fFsWWdlJSg
BZVT7rb5Mc0EF+SfnGPV6k/bRoLxGJobfwOY5Mp6ZQLWiuNrvgqfZEYiguYyD+4nY8LPOISYu1Ha
WNXLxwGkma0bvH2QhyauZnDB/C2WP109wMgJaZy/Z7pYstRrbdxwUcVglkTMjmyR6FL64j23+Riz
u2fOVMlPkjYJtlE13axSPVNMPLM43yDTg1Rdb+0wybBfUrABl5RR/MnkYRAFIsfZ2StQ/doAvqNO
10wyAuq8hfHsPgD1HzNiTBVUvzHFNx0CXRYfDZ499vA2OSPwvCtx8SAj1cdkDwdY6aXflPwcPZ1c
onoR20hWupQBglZAkYKT+jDDJOKfKs5yVfD2h8KkD3G5g61ASaZbX+BOmz3R/D9aqFmhE1xvlBMa
eC4+Cw+v8bPtP88cYh4L94r5E/+K7zFYem20p1dOklJvrWfWtoMrdUEvN8PTmBMW41EJ2Ov57ZM6
At97EEeS61cAH3rh1mndgfmFgz73GXE8SVr9iDUudoiyVNJCWO/P+t/9HdPCFvly1QGRhtTsp1ZQ
MV3y/vKfggeyaFYp4/hhnsnK6DrGVVUiLPKrTaXcXYCMy4aLQBvAn6knJQnJjiiXCE0XJztW13tM
2VOUtF0BNKB2G0xTuT6hTY4hgFu6vW0E2I0gyh0dBLDeu5uJ/inT1cw/gzTu9ZNVSNIBLPqW1i+w
Dp8ofrssS1ztbFuAGeF+rZOF5IIilojwyUPZawnSUzHJFK1fa7/DYGnsbMcFGlfyTsr+69+fo9Vo
PI2E4AynWqY2bIKL6ozXkpyBLU3WKxjUe7IHX5/LwtnYZCt5U8Wr0pX8LLk322pW+WJ1FsgnYCRM
wTVpd3nT1goR12WJEXS88kLsg66wDek2BoJcwvqUvHmtTg6xbCNEHSzgzbC4lu0oHI7pKG7XcEwI
5ROtlSoGRl5RFBYdQeJ9an2fo2IEd0tDdJIvJzqNdiWQQuMo4iokkKSXByqgtbwFnFkwxJJ/AUpE
PkufHXSetEqUCVxcpYv3pJJE3/fBdWPg3VpL8ePgxRf74cGF1js8IJD+eWdZU9oNlELmO36xwCrG
oa9Plxv1OdX8IQWu4UxYDpkqqpMSlKASPJlL1/XyT6aI/BDelmvrEUI8ZK5FT0FRhT+9s/JL8M0P
cLBPk7jzw0J8O076V12FZ9Wr+EI/ELnOlYEBumSVUNKWd1t+7LwllTwIggKcfgFBtJqivFecMg19
pr3Tj/fT23QuWh5zXimxaRa/Krk5NOOY4nE2PTTTx7RgKvI435jiM7ligtaR+CHHqb2RTzVyk+hs
O6xXfLOvZMrKwG5ePDRFFNuu+3mv4gd5D3cXz9tBYVn5pOP6Y/Wh2RWOj/sP5gkiaAhMDGU5jp/8
SgvfV1zDs8weB0majLJlSrPsVC8kNk2aNpj8gs9lO66cVojMsZ+TNMTdiFiUHclNCot7uu4L31Z9
G1XCbRMeboFRq/ESOWOjbJJWNgApZZNc8oQg6mY285ZNr7b0Ag0R7eP0THvLNCyOm7ZnMOUiJXX0
Qh1r0CIyt4Qi2gA7ouhG7xMlK/0GV2KA0ZRw1UuwwVi2RutyjhKyZlhc34aw4KRGqMTrRZs59KBw
3uOQHK1WCOOJfGhJLzwwbvvKuH60S1Zzr6uVnlZ3XPs93OY4HVCVBRCGfP6gvuW0RKxeEYjvGun6
9vcb+XpaC3/WuESD4NqL9rsS9gCy/5LTkqKmcT783DUbsWtpIHbc3V1m9F+J7XArnELWJSarYhZx
Peg9+X6blvaL0vYZ6YAxyjEIhK1aTo8TZEjGzHmkYg/BsLt1TXBrPcOGXClFyhdAepMWVceRigP1
qcOiPojld2IHqyvlK8ixlGUSQmOXiSTk7oNcVO9IuDGkI+/JdmN5IWLdZuEUJ3pWG1HGZb2EMDOG
hs9HDBUDIdN4b5mvdlqHHXGeWRUw4NaA3/g8abiTmzDOWils50hQ+eaQCRHud+huXqfUyjip00B2
eOUruVYBtIfiaQf6DdIcL2QHHp1IRI+eP9/WmSvNg/uXXu1vbBFxewjSFc5nXIP/W7fJprfYr7gQ
LBq0Jl7LvSJ1aWM4hAQF8cuYB6pZFkVyG79++E8LOL6Ez7auWvIAYc4V0lCJoJYt4oRY993+LnLc
v+qV/Ln52j5wC7OqQPGvkXxa/6yf9PAQMQoTxBhk60BPU5pOE/HJ00HPNxcMJ+Bfy9w0zIA4B4Aj
TxUzjKpuFuQ4ZlLE5HUWXF4BkJGaeMXVdAXAqCl5AsMXv0HLhZCAUi+kba1Kp0zLyPDSa1C3Nkfh
8Syk5zW8VHch+BThH4TcV57ARWIewHeracRrVBfVE2SEn8U6BMIVsgiSkYSY6Xf68PtMl+PL3xW5
PrzOhmm+raR7uqDiZGhvKm9hClh95bQqrr46XvjcxLL7H7qhbCMLXD06MpmcdIWUtEN6m+t5egps
M3v/OKzKiCgomPG5SHjw+/k/1HnIuMaVN06a2bICKM8QvxWKsQ2UkfIDHNrgeCxCX9Y/1RSeMNw+
RFcIk+vbTpgD6wR3QzyfPSTc9VXzxS82veK4atez78gWpUvbbpo00eINNgD1PrkyeFnyD8hCfVdc
3YDzMq14+05bW7iEEfg/QZR0VcGlamI8vVTg2NrZqRD6LR/j4mAmvdevWhMXel8TitlfSq2XrgEW
S4+S0oOcvYGhkaF6u9gPr/xj86+aaYQ4l485t7xCg8kGwbBxpNo31ljkM1n55VDcIdoQUjf0vUke
LvVBFmtr7qsZWPq+NGbwfe2uYi60B4DEI2mWwmibdC9cD316balhtoexTCjkzg7uL/9ZEo0K2Jpu
AYcP7TSdRC7FpjOGcfFnTsmfnDnSbGs/KEYHLRClpRjNbSnTvRGQv1w8MXoDL8cov/XW8gZ+GUAH
c0Z6uf0/rIVEsglkOagoKB27KlcO3hgbddOgrfiNP5eyBnK8V2O3OoMVC5vH97/Dj7Xy53vFjEhP
RYVX38NsPpAJp/5d/prZagzh9Kkr3+Srb7iWsQ8sLFkzjFWo+K0haTz98kBIWguXxn3xdEgeeVPy
6sxljRpFZEMobHLROe+mKy8gKDyUIGUvM6m//xVZpeQifhBOhuoDll1+9iXEkUUKOrd3P8sYnEH6
pjNA14kM5w+Gp61SrUmz0dj3mkn+9/qEJWlEgEhTsca9zHqFFtv+5/OfPmWXNRZcefToBC8d5s92
hIIYlEKaSUz1dX3CbbzHSm9/7hrpqbw1mP5KOLOwQsy2AcMPMO+NrBYHJAAP6lqFQNeE/M+tfV8N
9hVsLt0Xg+jZxpoMn0dYVBLc/ux349Y6FcqMNdO7TkfzOeEV2AIA1wly/AiJUawqjiFPOmPRvX5N
yf8OcfWSm9lmCimkGUNb/2azU08yzSMlLqySR/7ISbj2gKXsMpS+cdvWZjjKm8fv8yRZaOZPWZY1
y+WnEJvgurN+ujhpYs85iVt77oEJfiEYolnhDW0R85sfPcJeV8urb3leI2WRZgZPo0mUfJaptRie
TDlwMzdr1juy2gem25+3gON8Jf1sZ8NP532wFJ3MG3u+m5g4dsrDUmHKf2hkbxpgHYz/sf9A0NaI
EzGTax3/Fu4/EGhpWD+vN0MD3advDQYU1E7+UuOHmC+YDGACvILKMoX04Yy/7dJFwnFQNEzLZadq
xzyJo2iRfIGYd5LmrauID1lHLRHiTYLfXe12txvTEjy/ca+QYU1Mp3abX4in8cJ/wx8LMKchMiyt
bdd5XzEWFDx3Fhel8Gi94MGIENEaZj5MKkQ9ttKR9VqojrGZYywylCG/0qtAeZuzxRTbfd7AH848
UwipsH9wTsJKbcnMkGPszK21tOKeZsZfJjKnzMpUqjIgp1y4NI4sdXhArTu0K2jEiC994OKBkA4i
g7yOkcFKkbubtlp8Qf9IKPOAG+grdNCjhNxaMLyTfnqxogWbws1FW+/5BzH7Wkzl+jNvQSDKjGnv
DBXyL9JgKNHdfsbJ817Sj41UYR9W7GV+CxIIAvpIyDkKe8+GFfuMJJXtNV0SoSC/vMyUhpzw+FDl
zBzvea3AY6u7qaPSchuO1j7YdbuvNGf/EPaGG2ZUT+9mA1rhGeorAjnYe7m0o2Df5OomevvjTeLL
+LL16oR5vu0y1tLsEwQTZfBPeEDq5MhchHRuvegg1f/6t+B4J4x1Fgg7DjGutRXh26EF77dvOp5V
RtHy6h3seJF9ASUQ7tpEWWa4U1OqfEW3kwBuu/mO4TOfNw8+8OOx5KWJGTCLCdNmbkNpwEXVVsDL
3ThELUIMSNivyauQRKXvbKWUU5XjgRgRQORFJ1DfosviAXa3j7iDw+mlSha4duYoSVj+WtiNA+yL
TLAWXkrVFlxCY1fxtJa33rBEsJ0Iwh4RVkca6PU0/Vm57Pu4xeez0GRmeZ9i8sEfY4aA2l/U184a
VQNGEIuUigMZz1Ll0OZYjjxaQf3yVKH2pMf9oUrrQAB8ujP/AYhHNvoQe/oivxkWVfn8I4Im941R
Jch+YJNKBz/yyFEeYMNeGl9SdDvdhapu8HgHdKQd2+XteOL1YjSFOCn7ZDRgiNx3huH25vdAU4wz
JdWNEOlzIU2Fh8G+7ayvUXkCicxnBdwb7IbCTO+NGVf/+TpTcm7hjLzm6LktmAwmQunuhCor3gwn
cyIsNlAase/uCDsvkwa/CxbAWNj1vq54IbqmrQjeMAn+rrbupBySTDSV0OTQHV44zElJJv0qkrws
3dQM+zgXgVWRLFfHfmC7OQ4x/0QLlHQjwykU0gghW6pBuIuQcnQkLMNLidMLiPo1QNsHbxCBcQxp
1wGFUle1WwGvzRxgAwhRjL88/caPVi421Ld50Q+QFwd/hwMtZBexRhegnMGiAUUTdForgIOG/W7q
gf1kP2lPiQok4Km6kyncJJm1ZihwyNeEyNMKfg3IIg3li13OR1+DcZJJp99B9H8abh08wmqyCb3w
XWYJNRyKkHfgf17WuRXQ33+m1+rV4Fuqws8W/5uLOSypEB+UfV90XUBIVAtR0w8eW/mEO01B1wRi
+jzrgNeP/3CBuoTLc+gxnnYQEjEea0UL+Zx3GZFgX3/m2nZK/HO/kNJ2G7Qn6JxcdgQeoJS3hpiy
Q/Dhe4iuFIcn1hWkdeSR5pEyoTh/TF+k0AqH2i3ewdQgNxm2zusL5lMfPuBWViDBivIUxHCvv3Cu
xBUybc04j+BbQFXeP44Dppfy6qg2z/JDIOiPX+5FTYhgAzZHa/6o2ZetjNp307tbh1pVVbGQUQDv
KKQI3MOOXxjcP8G2qPGLIUO/NhVfXHW2YGCBwsw327vMcj3zY88zvBD2CvyEX4PaBYTzIbXXMvTu
rBsfOod5zDyw4RWY/P4FItE5xxXKM6dxEaa2UjxVjRpLf1FsgERLDNpxdgWikhVM+EKm48+sx4gI
0JrOBTkNRUPcFjXnWFnyoc3K6NjtSYsjfffaocv3RdIAZpkSIvH/xp2U3hg2Y+towrw4jFa3Vt4Q
I5X9zusVip2S9dSqiTCZKPfOmW00/Pua3niRe5IeVsjhYwAfhSdDPQjsrtDuWw87pUrcfU4RjSyh
V9QsRY4b3pLCApkIkgK4nJimpXjYHwGLbrHBntbyWA+oIbRcUAJakDKX1Gny3Fg988CVJKFJYs/F
ULjgFzMWcEApWOxgtu47TPQQ8HNwdofkbSqIz7HZOBiCzRWhOqQ43hHPLdPXwsrGbDt+K4U6sGe+
IPyt8katBzEGBGFSaGrMvoZBrrbRF7+f6K52rtkmyq3Tfb7VSsMlc/UREHTblWY5z2G9Jkvh8i8F
skeES+I0cY/LSFFfDTgR/QMLFr/GU0L6E113/wPuGDtHNjorxqpzt7YgoZELOdeOUJGhY5pfLAAi
wlD5TgU9wTc0lTq0SCtpAek3hItwFlrfEcj417ukg4dTGBPoHe57x8iYW/lSEeuD1mf71zDbB2W+
l1h0H7DDNWLkgws60pYYwB1ZdsT2Aq8bSRIRDb9/gjhufMaflIWfDGewUtgfb1b6VnMcrWLbxwGk
lfUOf7YMeyxzwOCrKBNYqdWNQPeu2FCaRZ42PI7X05Rlweh68cDqkPRmo2+TzlqmCFVDSy3yWSS0
Rg4ermZ8feQWXLvtoFCsJ3qKcMXa+HPMQs+TDIF1qX+3wFvjEz7P8BAiILey+B8gqcAyMmvx3F8G
5y4sCof0ExFlBe2l8wF7M6JfpzIZQVFdITALNeh9TVdeTC/L/dJzuIrAXF8I7VDPz/ggYjwhBMeR
hRvWgcaEYpRpkwvJQNyQtQhos0BQBuCwZafgcXZYCABP3Dl9bAJQAkdQrLQgDbGPZzXV0MXhZXp0
U02Fw96Su1xFhJEK9zV/jg4J90tWb84Hc0wfBLhKtJ+Pjouge+HJUpk7GEtUQCUShmTA70hSW5Mg
T+auAykWDOX0ixUrb77glyX1YLws4gNF0p4BWlTNO/0dINb7FXCD9xaoec4vBXdzx1vwHF0PpcNk
qXJO1sfIIVE7HuTVJiV1WnKb5PZ63rRkuu67arGTGdrC0xR5n+c1R7HD+HeFLWaXtfVo0NeyT0BL
WMtDKo5ziBYAg5AfUUl+YFcWkDNGIvHetMNVJj0uysjmk3n0M/IKaN/1H8QkEWrIvJUMosc3dRRf
SsfCejR0Vr77ueW54iQ6ypJsjn1gpdchb3Q5UlZAU4e+5g5z5bZy9o3iTPduYxZuxKC7xsrPeTcF
bpKxFmU/dxocKnXWWQSRW6Z7J/ZxcdpiJ+wcNZ551wPfEEpsBMZevmUdeFmsEL6QdB4+DTYjVHas
jERKJn2yvEf9g20Wcvp9DL2JdIPJsKKTtNNVPoTdE22niTBADHRZscjp1p1EjazmvIY1h4Gub4cS
/OAOVLcUrxByn2mkO6HujLQIutWEdf92DXiBX0b1ZhCjx8w7tlgFQjYLj4UUWF4osbcloLkL2zyA
WqA1ft9D9VYg8gpMn9Gj6FnreTo8si3Pdh7u+m2JTnGcy/nS4pQIm6Tcjrtcmg1Y8oQkxwI5jEVE
Zt+otwDqNaOJMHYPpBEOiWGxIoaHQN7SvMMDiT88tJCczGJab/agTPZyq3zaRpUvcp15wZ8D3CjH
kbZfXRzswTs7jlURHMyrthOxJQVU1kU6b4T3rFftORIZR2M2iU72q0XhvT0hfs8u9biGmvf1hCKa
oj6sBciIQ3ppGBT/8+1vo4kFilJKVSwMFnEj+uy5JyxQgT5vdcTGLbHVw+LDrPgrXdCH4SpWId1F
2watb5xsv1YVFXeFSmILV9cmzEulpTHgSWRxsfqVFK5d5pakTgmptjNpCtJiNsuO6c+d2KBw+zq9
XvEw/quWtT2evpIxTSNWkrTHyA+PXPmqF5BxIizgbpcokFKArU5qj5ELTn9v0CeWpznit+ANgW9T
4/uogGr5dMM6LXQI0AKSMScdhr+RVF6MxIiV+GyEtRF0Y9G0wymU4jD1Ktet2vK7bzuoCRqnG4l6
2cvyAt9cVFRYfgc7QNNysVBZ++WNbUlixr3nAVKUaGv4i1kfG2SgfWfi85n7uh+O1kCqdu1HeXsx
1jwamJodg8Cj61ibn4z/xbdUDqqvmql+hkh7OkOPwXf6xb7zmZA+xxj415Y53YBkfpl/iwW2E32K
Rbh+TjXbVrzxMqZISVVZsFttz0OCJ29GomqKd9zSfIvsy50siYdSD0eCGJ2sUmgTQOZDZWksHw5R
gAHeC6F+H4RWg/AvDCuoF/Mlc4xEIzmGaNCLVw3vwKJttwyZbJmEhkRBMdikNrJPzXvhrVaAfqJt
u6gEP8OOT/5aWn5KlZXBJJQKJbHIAsOfX7OY0Yi8qkSylgz0js299Gqq3CuLUhsGjR4HWUAFEKXw
tCOhVPlOHFKUnA/ikd9opyRc+1GnQ7RfQqS4kttPDSp5NDT1ZkTOwpYlo5ngKvAWUcTv6DA6HEpy
dgEhHoJMsSD3Rd6qN2v+tva+kBv5o1vyhCcevM6X6kg4Nj7n1dKVVOLnm24Qwku6aAsgtIHq+wPi
t4RkEClhHsbVzl1WYb1r9YVo6hPTQoKPJZVtnPz9Vh/t0KS3kvJ3wzcij1Hc6Z+hgVTTXFIEvGl2
59dSFZOpPcjwOUVeMOHoM4S5Dld3mRMQ2wG2OmcQ9YZzLLtsvhuW62sGa1rtjD+XZ7VCt0vLBYD6
d/pRKySw0sgJv88kWlwLQFF6JmwLN1EDjYl48gRkZUZXvoCIw3i9mWffYskM0i9UPmBvb6ANIoTx
eBzvzcvlqZ6YqaepS3jcOqAXpjlOySOsYUwmyTX+y2pBktGyWvzPzhIQCw3ArZ0DkOUXE1lmcWOD
KpISolDy4o6Q7DwQdtsSnkdhXagYQztVolDKpgYroun86doIOvbx/T1kZPZptg3cjyPhB7WlbYkL
193Hgr3tCOxDKPxVBivirsXYIqhUT6XWTSzaltxzBNiH2YcnmP7Ikq6xLaTd3Ac0ogG0l490Joai
jpOUUM9MHD6YzSlukmpORfYute1suz9gpUYO0O1ZbYC5vHtVDatt5gE9kc63wtqWvlrmJj0xtp0Q
onXweHBpMYtuKnkk3HLux/YpqXfTUk7pl9H/7MGWMb3zWEUplFQ12fcaGDU0UMwE4F3Gh0QZkexr
KzJWFSfkRrgn/mFEuBjfqF6xVw/f4aQkTs/cY78C2kDJMgEUvIgIjgUh266INKnu20oq5qOTd6R6
h4FubZrgEW+jGamtjOR41Z/UXZJIwbsIiVxkFz5LrL8A1+IcyQpH2qgv5x35JUfbhhq/6RWyVNCK
ZsPGdKqm7Zl+5yqxru1rIcD5xhONUf1/JAvQrkYLn8mVzKTsg9jqNJzq6QllOwEG35SObbVXRu/V
isYNMPzvDbklTNb7TAUPy/FwIzwaKCxHircK02puF0M4cE05VqEoUlwTOi4yT7tSrjtS3yleAExY
3n4+1e8XrJaG1k6xxgwhceWVSVPN+Yknxg5z8Tww7bOm8SE/I/FyRi1R2vdZu8Qg9GwjeNfOtLY3
OxW374EkWz3TJhZ3EUebMOwINajpEMOHE1WiQSEsmeXlSJsg50q8GAKdWxvGGrWhxamdGUJy4qC4
FMsV1P0spF72GT/zJHSeAMTL/4xZ1HDmKq7oTi0JpQunk3LLYSwLhX/bToaHGK+G2Tp/aDAWMGEV
kr4KC3c7AVTduTygRQL+NGL/dsUQOgd8r1lmFrGmuIVXhR1nROETzM/Z5R6dbnjSQCFYkTdzbIKm
WcaUzq9BMXo0hZiYhKrMENWCN3hY/JkFxbBOl5vEyfZq2TV/oxDrdTxeAxnvVbCCr0VQLN8JkeIj
h1Qp8TXTgM7qvv/+3GbZL7OnK8tAnqPkeiDwr40/DO4j0GWDYIrbEUdN6+jTeiJ/1HTaiQvBZU9l
3c45isBVJijDzprVQ4sbOIJKh+ZhnK7qlwiQx7kBFn8L9xWq2C2v03S3OlBXNDxuRIgBcBOgTo9B
oVKaKeDgxH3z+PQj/1wxXol475G4z2Jrdhtnd8XtzguybsL+dGsXolFD1k5YdCimeg47K56oZXfc
NXNgr4qRKnpW4tIlKs1cVawYmaq+rsumKg2Ev+0CTS4LUJ1Yi3FYgnCKUFYHi4A7qPDxap/T+/Uz
auDdZxE6cmDAapJXKn6CPGgBZ+qdRyJVbqF0gZFHXTd0BEwQ/vaI65uzbCC2/bwz2xF5akxhuCd3
OXoYfPL0Lqj6D0UaBOsD9Ppd+96G77S8smNhDJWrIgGDL+EIlsn/wgtDUBu+eXhj6kQiuRXpvlfV
Pmzzafsvj5Se6nJeC85bk/82212g3oXaqyL23uXxVGZvCudRpVO4NWd4hFTULJGwXw/TPgoR8WJj
xkIh9hL3TXAPIGroEq5RENslr5GTH5cEbpVsvSktaIka68Gqm9HUhGkGpP4tnZTsG0M8Uga2Ha9Q
DmiCyCgx43z5nLxqkzbDhKJbMQDaOEeg4iueLMpUypdNSJ/4sCPwWST9J+P6Gdf8H0ruCbgeslWq
UzD6J9vx2DuFIQ3AFJlBUa6RfMqzADRrXBAHTQIE0bM7vAFTVQNI9CzjKtRjMkX6cHyDyWFqaqj1
2nhoRO8aqIS4ZJmIW1NRVjRAHzOSN3+FXGnhUGj+50xs78wMGMLfIDI89SfuKH7y2+FPs4HLMF13
pPVOst8HxWsL9WEl8T9y4g1OuIZmY8cPXAnIuOhMfB1WsTW8+Q350PqTdcEMBdSE/K1rndCFikOp
39P6FFI1xSM+P0iyEByD0xXoXmYKF/aCmv0u13ZRe7YwRk7ahBuHXqNyEfpvBvcbxrDUAlIYGRin
HJfSLLIbjcvJrPZiWo1wwi/RbT/cIg6HmSn9MdTIjJyjCNHkpye+FOdYabymZoPtjnmGIZCdc7eL
sHc99lLO6igqBVGlQNJDj8j5fMH+SQ4brfKGT0vTlW9hOA0jav4xhW4YQmk9uR/iIcjbeqyYuhbD
CfQr7cyHxfpbZgYCdCSDxalLuCSkvsMDZ2NurzSh+pou+yMw3LrWKMd19BaXl0Zf6b44QIT3Ac6t
OpFdjoKNvRRb33rbhZyxkXnayE1RKWi2h6IwZiRPOdUdmbxHUrnbCPs9nTtgQwSYM5a3iQszEjZ6
i3ijQtbLRIijcnYqsai/c6swEzanmxy2JZ3s+djklHVVzm1OgmqwDTLf0xJCF5uaEzPSqVyMKtLl
5JgI2kz/hj/vf5euBcCsHug85MOcexwCooz3Bz1P2BGz7TOGVrXMBsWEvjOEAmjynEEG3JaieXFe
LV17n/ZWDZyjOb+bb3wvMkgKb5uAHURdX14lFA+nO6g046z2JmK8gLV8sXdVRKcCbIzDyS4qA82a
6QrcDMNta/4jelUk3Ro6aRSMD3VViFgdUYclizw+px4U9Djm1qAmbQXPym0HGBaIGeOLPIHKVog4
cb5BK4T/WLrzGIWT4+i1InZGSSrt6BKIAVkHGQ3kDs2laf+RpaHqgyavPd4EMBPYFNiBoTqo0sKP
33Mxjul9ialGNx9HRUaAU5atwx2B2JVxUXHhl5mqwZRTBwNwtM7IB64E6TtLYfZnYD/GUl4HzMYZ
KClaC5HnHRqlMGu0uHBeJP6Te09eiEs36GFi6h73OD+AszgrDchybZjihD2rmQssWvFqnE/GW6xH
Bkim7rXuYOQawUw9yAqFYdOj4qbpksYHPEOm85n+xkZ9MGcGaPghjvlrvuqsn5NMaUwTPmmhRweJ
RONxHgFpKetkTDziuMFyj5jgAUGDD0MA+2P34gtlctLmsMdOYC2CsIH5l/4TvYH1ADc3kkpqns/s
70yNVQmFbKufH18ydaZ6HNOSu9cZf1xGajwpgMMX+zeu2W6OXARKVughNiJ3GSP238HCYuQHe6n2
tsye5ZiTLWKiyE1SnXoBLu94t+TLvegI7+CGrQo5AZvoPRRuNiTpMiEV3YLil7ocpgdC00FOqA9V
6JqOrBpAlMg/HAV5oZRCKHOgCMoH/fj+dnVzwFcZqVVBnUArJnzHsJVr5FjXipML8a9bEsGi7YaH
T5plz7AchDLfLIDvCjuEFSCqpN6fGa8Rmp2BfAgc4PJOF/wdgrX6txX7x9i63Vqgl7xB56bOBzt1
BIXi8c1JiZicUJvRsEto2iKuHdvC75uM122NHEs3YYNqGwE+050ngK1og5xR25IuXUrXEaEBFAAk
/5FhnKr+fsZTZcvBqSFxNH66a/stxP0DViNkzReopYD7SHkGV5e8nBB5CKTTJC4Ecjf4pELfSDKC
zbt2dOG6DVYaKPuDMHri2IQ+eY2YxFKo+A3foApKdigdbFBLMxJthUA29V99KZIGPkuXYf513Xg4
PuR/zrA2+qH3/olPFHrLX5sauGODnfsL5mVjic5gzz9XmFHisqc9uIfl3nglNKdRqiA3R6/LhFYw
9gDX5Ts5iLOAkxtJ8RIyoltMpf0LnKwCjVhYTPrZcgLGhS9DQKk4E4UhKMS5uovGiEORFqLTdJ2a
n2EuqvEiD2XEAhfv8ORGnEHEfq3Mc5Cj9+kyNRJpeP+3Z0Whyh6vDyRHDJ14YkbE2xyg4MwH98dn
dFT6tswRgdOYfcGDt13uIDn3I5hVNfvgsuhC02t25RLsU0j08ZtUx8OQbJRn6zaEblXmfs4rxLbA
7NXQU22W6if2i1WSp3885XddKXVwB6eFMmLpiuKfTk96GTp0+8MOVOKpl93GkHq+hLdcS43u/zME
BYqG2i0PJWiGydgebR3SgTMMrbKIjADLGhO/pBhF/A0Ghv77PUOLlFeSa//SAcvkNntgYFsgqPAv
NOBhA8vBMyi8G1SqTT+uRu0WdQmxzaPEkfOcxefcPTaFrYLHz90jTQLD9AEaiEG7SgpaTlwOWyEp
Ds22dOP0NHxD3qTTCChVu0cL64ck10nWTS8IS7zb+9EsEm6oEtWtpxy9x/QkWk91mFx2drbVroVH
ZDmi9YvOFI6jkN2Hjx/sZloTws1WrxO5ZFiseCeOrrjHiLhg3jTjMF+PCvZbcyAmhedyuna5uISv
viQCTubn9Z8CfLktLnJ7HatD7yXBt9yYnjZQw1/R016Am/q3MjxknMIUEbMEmK+eyhvWtah+qwWC
lyX7U5jcGN+er4TkiyYVClPdtaIpt8ya6bOPW3SdO3qVB5mNQnoMttOaXv0/AcNTVvWFma9wFlLX
NGCcfqryWeaN3oXlciLFrp+fbb4zeJLrxytBl1Qk32JrXDIJdl0hs5LI7CEilbf3/55SNsxJYMry
Y+dUGKQv0M/+xEB5dhyXJEzJGrMXuR5PbvdNvpeooQM/mrT8RoPZF2TaFaPD5/xPdDT/OqTEIEet
2gXVIml7DWpkjtx20THUEBL8aRA4jpjgqnUzv0sqXUTsfuRuyzM9rTidUmBgytDrDU8RTo5eJWch
pX4d5+Oe8y5CkgqW/yU2UDpRSuPk57salou/GbOZl+tDd289lzhgrVFSA5KB2TJJa7vScU13HCug
3savjJZ9Cqb3BArXDFpSkwTTMmpKODOlC5/wvAJWmw4lQUF5CTG3HZSfEnyd/UsovLlmt+SmYqXE
1X6pBJKbKA4UkEngLErYnrMocbKHdGhY2aoaGBGBmKZrCWKwUxC7N+3hzGHacWEbKeY90z6BlxB3
4SW9NA0P15NZHJf3hGNr8HoDwLCU2SAyH1gLwwuUd5+PZAs+FTAbfZmFZRm+NqjBRWLWJ8XcoP2d
ee3jb7VJo73JIJiGJ1nn8X1yzEjM4IFAH5uTfzVRO+509zMQv5i8bNho62dR4G19QiEPsfO7swTE
hF8ab3MopbcmdyQXtm3TkarBsMKHjK1qhlBGQZBQMduJDOA4j5aRvjLLKXN+9k+/1xtlRr1wyKaO
pWzmkExhKHs/lxeQ3KKBslU2ckfzaWHz4LZCaBRC3dWOyjuDDyb7P3xgJRCM2NmTj/frTACAwsuQ
45E4W56zUH18OKETKu/h+ICsXeM6/ZkLsja+sfz52kYDvVF5VIfCxEddr2NiwPqMEVr3OlVSgp2d
pSleRxNb86sm+kn3Vij/rD21JQlJT12hZw9W3ZoQOMbMrezvvreVv4S1pAQWunhwr/wGiDE9+NY3
dNWh4ZvMVXmwl4iGb68vpz8PVc771xw0pFoejWzhK0tLMN1m0SPqkvbtqkWer67LkpRWk21V9zDm
K6B09x0IeAdQBQEk/CckujLHoXP6Z6koG13PK0tcd7sHJV72z29bFSXVcA0NXz2LvFJ3OGMOkuOH
mPTtXQXAHbV5utBdNHAb3p4yIAipwC9ETXTxCLs225KQzCOD8hB4Z4dbzbTopbJ2i5KBUz+EeTfT
eMItHxLEMB57DtM9SAETKGTLI/lUEyoOAF8GwxC5BMWSXFnmT3CeRroHfKtqNGvWNtVq22731AZv
BRRDErJyAzIjyplF4VHJjwCUzysDJIO1NwpfhqmzJoCrFk0fagHXjKVpFJYHPqC1CWzv2j1Bn+8B
PrXLOpvZKryeQst6/BxBizb7dDlUC+zbOwzTG1FJCprUUa51G57Lvmz1GmIkB+xPPrNdyekYyNWZ
7gHzJNLTSeHZzVbJB8gtesZsUZBHkjSVqIQ/4QgWUSHC/sVeAjWD+ZlE8Hjzb8cZN6Wvw8+MoDtQ
W6ffO9N2+8VETHG0UE6CTs2DzqlFc1JgF3BZPkkmYo32DgDO8NrFi/PRYtO0TRXB8/czFjtqjtJF
AP7tk3twbPZXr+2D53g3QZXlrh1C4t0rTEJnK3S+4ao0yPHZmFOYg6DwQB1GNiv1fJRgQ/R0EDgq
xDmPU/eBpboF/sK4x6v8LqlY6P49ZLhltKBBIC0qH4SxP6mrabArfcPXQ48zXs8SmcJfmAVgCASo
djY7EBq+2Cb0RXb6Qd8C+dhm/Poq3bAr6RF/u/eiRxNaun9JKyPOtX20Z6MLNyDn/FA6X6bFWuTb
JGwmZxCHYMrhjYodtf8qXrWlfsoarsWHrAkBVuIETUMow34aVe8xoZcNQXPItYPJkFUm3cUQlwPU
9lgSnAA7QUN25T3vFt7eiPr6CZU8qlEjM1MYvDt+LxOKrFs9mf9Y4YVoDyf+qEU8BULH0OLsbCM4
a+OZAgTKaicU2UAkVfvp7sEQ9xcQHQdDYhu7CE99EfslmJs7kfhpo7O9z1cswEto5sN1S+ypUMZR
lktgU0tXxTZ6N2QUrKYYRrqivGHo0nOrYCi89i/8VW8VABSm+wZw28KPlhaBVrHqcpJ3hBe9wHk0
ySvU0P6KDG8xD4NNo+QAxobnltXcAedK6ws7OmWfMfc/hebLRUXorhQ7ezu+IBpr9DyRPzOA7Y6c
YtKTVt+TROUh7gmTnj/d4R2hwCZOPludo/RKTCsDLynswfHq64xKXDzaXqudGmnenQv28iI4LAbm
nMxi+1yKC93S44wxHaeGsmyk6IBC+rnUtb77VuJypkUqHLEvHSZd+GVL3eBQYP9sbt1M3TkpMYX3
QuNm8HkHArx7th8h32kOK2/54ZECh3uYKAyRwst9Z72X6VfMHzpvA1pKzporw2Fm6Q+t4OuW4mPu
YnPfWZYpyf1WKgQQvpy6xDl4uoq7n+PpsDqPEDSmoGau65EfPDVxDtQAmCFw/CE+04VQRCRhWWrA
4DC1E9s0ZuCm2b8eDfkTS+oNRJWCM26ZueNth5JwDJRU09WX3+H01dsoOJVBAM3b8wnUb3OTsKvF
lYCtLj8NmcOneUTojDSwFyDwdgohTvb26ESE9EmIFQeLpU1yNw3OYbgvlnVHW9rNnwZRZCxMEZrW
OPZcmnvDlhn4JRJe6bealW61pXjwMFrQoYs8YNRrYcu6CX95nRxAl7/iHo6O3AJDo3xP2PIObBPg
5A/2ObScKKUz/W/pl4sLHdaadB0IAWZLyIbihxOeK4DilkV3rVSWrMzElZRKVHUprWbmIiGjs7Fc
ADR7U3ALM00jIh15aeJqUXkuDIG5qEcsbgBLcX7/s2uN3fzZ05CE9quaTJrw3r3IvTy4jmWpAWqx
mpTKuR5c8nlXCULb/yW8IlFvu8cgkR2LuYS3tBXQt4SKna0uEvWWIckLGEqp0NiZ859cFSVNP1w8
Z+SgKwf5IJkC+BKr5jqEAQEQaVYds4LvB3KWauDktF+4o6d5BTn4cITW+3LcNXmT1UWXxvhv7R+U
ACwDkG3bytSySnjv4om7EYU61fWTlbR/SvGcGwy/XuIld5yM8wn9grloWxo1D2TF5ljt7XSGL08o
tpLsypFzWUVutkfzcRnlwSVRFwQ3EeNzED1AZi827daRzQrz8pS8SsVlTlUMXHb785aIS6d+O6es
7F5riFK4JbLb1oEO2Pug6nKHkp7cfO6eLni9Azxq3XpDP8fMnXZ034h3Kc37COT5S7aoEXXxl1QG
aPWtoEpYttCY42W1s0wzll28IOPo9l8f2sJGpnN0XGzClR7cESx5Ddnh61YzPXCkOEKPCoiH5ZxG
d7ajpvaXJSAvaj8VlSTOfiJKa+WH+TbopmySH0fTIn0oA/rJGaK94LMLwdYzmqnCaVLrLC86mdIJ
6XtNyLZERL0MaoBiZfN74yZIF59h7OWmo5C0YUtKmerQtwFFtSLT8jhKP94oPgt7PtA7PjOx6itn
N7/GNDORRU3cNkhfK4NvYu+hPaAFccjzOIj562fToy2rCIWEGYd/XESJeNlOTBpR9Bmcyy04HVl4
EuQOCJ7MjZStQFVm9wgrQO1q4iT0A2Sf7P7kKSl84E8QByH+CVtD7mruqkVQ4lM5EdvJp7UHow3V
oN4gBOfuMYVBBNpceGNxjtz3uza0KWzP/jrAlRKDzfa1/hkO5359/W3k+egAjA62Zq9BxMd0xrOD
Y66NVEpUfSWkYaM227HP8+4CCSLbmuSaMzTgeJ43B56guxbTC3/bvZKbfDqqop23d8dfK7Xo5O18
sPgMB9oep749dwhqUOfx75OmtKIF4iOeAsvnowS7/pl3Vm9CWIBwKWW53L71wY1S/cXFU1xeVQlp
3aN08tao6fZQBCENVL4Qmh71kKWVtb5EUk+3JoPno0RxV4fNd+rKl0grMOm/yOM4+Xl87/4JxgGC
dGEPPaInbgjX/TSP9UUNdEdRq1a36SDvd52+Moza0ZK8dCbREc820ARbUxZ+gk2Wbr84pnYtbAC3
7qXFTzItX0B1cK+s5XYpzA3vFz47MoX5yeglCc9Gk2lnNe+6jN7cvrYz5JmZ3LSUJynNjM6Smhza
VX3Z49V9RdHtrq4M02i07s5CrwiGSPAym/RAhyn9RZdR94GCgeahfmkDcvL4EwmvQ4EprQj2vskG
7V0/tp6wU4/IrVdKqImvVMeRfrl3NGI7+4HZlEyZR55EApsOlwklTifeYBfz+rcJn6ajE+VUDW02
3VzOMCtXXOUFS5QNM3TWBZCZFBp3CcWYvkZg7aGFf5kOgvL3DZXMN+GDcudBDuqjznPb/gFsgwC4
o2Dy1HHmKyc5bu+pRGBVLQocCn43EIIW7L02jCMJyu2/6cDvC/SJLxcGL7yYrqZ1WCHbshRVL0wJ
OhvUD00tfnpGOYUzw/rH2E1Mz8teW5uVhqUCLy94czMsTyQNHShfsXqCJE8sEqF9q3qEdArjAEwj
g+O5nkWErFL7OwOY1+Boe4cE5rMQqyM//lHWyq2lJuWfkAoJpMUIRvQlMj4WkCAYgfG4dIb7eiRg
anql9npbeCp3JEoYgj4+FBIqy3YZHHDUZFUnCxCjQ8cVI63tcfUcKDFRX5QXBKrOoHoqzwt4vQq0
C7O0Ju29Po7Ig6Bnd7sDw5mOPRY2WMrlzP805RY7ueszxKOb/Hpr8OtHzYFUdeoUKPkJNRBM7OfG
Q6GKEZtzX42A18Ohgf15RI/J/LH2g32YKDRwGz1AqwNTIsJsSyTCC37yL96D0Rz9oOn+Jm2IxCrS
rTENq6oKuPePQgR3N+OT58B/v55syq4RH1sp0fcNKlgvaMtbuShG08bJV2u+IQV4OG5tA6TSrUir
TFpgYRCwDGKbmggKMaAJ2BMFuUr9ApE9DZvLsopQDSiSMsIDRrd453XIh73ioS4HmGGaUPeUrdAn
CnUb1Fetkv5wUysZnZ6jTK+dQPgxv5k9wSLFrDY123KPZNvDJ8iv848FJLXn3Fs/2FbuqtV3wN6Q
ZdD+VHhfmxwwEvXm7fyd5/T87WZpMnqmlawlwdG+XGuR15AnuuVf5jsvaW1tsPugvjdSfL6Iqfrx
T8EdwDDDzwnYEqBFUv4kQGYWQhBtWJ4KeWxyqjWgKqve9Tv+Db08CDzC0RqsGhteFnzL+4zkpaoa
SMMCbqC5caGCH+zd/J1Vff9P+rMZZn3ymHKCfyhPVZHlNN2fWjV1mFjPD6IYoZpEv5r/Wp+WxSlG
EYB5rm5VMrfIatGQz0AmsId4ToxG92nbCp055E4ahAdE/gs4SW5W3GnpKQnbVqBbmWfiAHmZB3Ck
zUpgdpwaEtCdx6/eG0tsCaT8j1pU9/4aQg/DhQxjbfqWzkgCtLPXHdpLMEaxy13YHMXXktAq26vK
agOnJugaF9Z+rXfnN0AlGUJhtR7sg57eruSszefbIAggN4UK7LocBYHF2MRjrLGsrfZY3398l9lR
3n1R46Kt3yyE1nd6RdPrNt0h9n0d+qRyzGllFTw5DN1R4X91b0eKeiIcOIuQiS1dsEDOW/t05r0R
m2yh6VCQJvZQINNBuVNSswZppOq4Xb9ws0VCEAT0I41a/1jQh10BPrmD3VoC+PXFfcb3YlLuX1fB
9cUctq61CCsxmTWvUnN59mJbYbjlfVbsES+sEm8+krIpc00YhcLimxj1jLiiRZTZ30ggihO/QY3H
EjBAMw8ZjO8oOSie6eh9S/hVvAJFDNj7AbByXYv/UXmyBdtzcln52zdqbIenqriKS9VZFyiX4FbK
+7DMON7nhGvTh8HQ7PWD6f/d02qmEIdR51a5USf7RxrGj8wWxDVook1jAHzwatAKqjv5JU0jWLIJ
A4KBX6erN9woM5PlTrxf1sAY7NkpMNSFxZnWNflFayJUSh1lSmGVZt9uUI/osq0uQOLIMP9RQrJg
2CT1OXIZcfdKyP9pUaWofZVhpI49iaSDPcOJWtD1dFMbE1AqsHxjXFGpUIvk2tzw4uWUiBgfC53x
Ygn5kLt7dHbysVyedrDA+qHuRwNSZowhhxI7cjbuMpJphMNQ5Fz3QkAVHBPx0nyFmcgKEQSYgnUN
JH3zchjO8HLD3C4JbJ6G96KVF5PrFMs0lDXpXOk2ZMzz05JloqhwV92jQLvHlHSg1eD9lkwBoWrb
Pjfl7K3bqoOlfcFqNDT9SV5+Fq8yKkVr1E1JwkCbP2tWWdxi4+GwVV2IEqAmyXCk296gg9osG93g
QALqHhKcuvw+hjl/mbgAoWY4X/dUIdbcdsMJyH+Jdyk/6bjxSdvdO44TLivi0+b0VIQCDJiWD6rP
IUDG3a8oyBlJPrCoqgONH4OfSGfoUp+CSDHuXPxn7tYFtXwIjEL8fCfLBkBG7LFf/FKb0h1efBop
7ZUMu/pwFnKMFxpqEAYNFB0B+jmu+IP8lRQFftgluWR5PT1TomNgFhjOMeMIjXStOp0Dv3ZwEuk6
o/QYgigP0JU8WeInoNkIO1vL5umPN3sJFNw7kb0BhEd83i1o6Bw1yd77Ll2joT+EW9ieYjV9OhvB
wD3pyb/c+GQWnOVbaetrpp0rmInaj3Iv2FCxKRHdmhrXnqxwkdNo3IOA/o1C/A3tLsvFIQMX6zQR
urzLW0zYVET1xjDb+Ok48tZvMUYZPSJ7ik6tFuNtsgTdX1o3xwXWm8UFJjGR75oX4EeTmMgsBdZ/
okmx7Rqk5wR3JlK21H+LvhpCNZRqjg5WTc7NupH3LpN91haZvG/pmEcD3Ilg5E4JJSqTFyfm6GB+
ql3XAPOChNyn0VJs6zpkiO8NaGNDu3Q+7jP1TmU3B+HzqMHofgn7+yQncAgiQBY/0rPoVesafI8J
uDp4or3l/dOhsVLAyvWUr06KuoEhlKzQAkYUtp3o4juvRrLx43FQ/oTZCN/CjbVnDGjHV5EAXHc8
6fFuonblSRq63kDj+7y9ozfhjKYusBJSjSrE6Hidb3L3ICara2gVWBnAICpSCU4MEAgo5jk9ptG8
EQP2fjeQhpKRlVU2AiMU6PDR59LiUVaabsUq0spCTsZsa6ySmAO25dSTiBjf2AWdgtk0F49vYAdx
/vAbyahKspTmQqfUJqgrTVZ6Ms+mhIO2PXB5AFXHWnM41OVlgT0o/7BVyWJ1t9dBYco0FX5xF4Fw
mgaEthvfCu/q3gvXni9aVGra67X7fhAi4tFHe0/FPOA4I0ZXeOBQveoqebkzNkYDRiMqJPl7/LdO
f6iEIPnkaxJNIKK2O4jn/BdUAqZ18dy89gmX7Nofdl4wO9duYs8qnT54sfmo3VLea3iMrQcbB6Tr
wuJzNAZTwYO5QppyZHfRi/w+CcHIFeEeRpHk7vMRUVBta+CPZBxOiwulJsskwq9l2WeKwccWaSFa
M0kl6heaROudYbL50hLLDQdmjeZ3I++mA/AWRVx10sYJXcIsKqMGaMLUUELQyGmVX21HaJTEmrzh
J+UtoWSMhSILTYJ5adJV0dX9mJwWdMYOFJxevTwdTMY6cB1PEO7GcIMO27idiFnwTOkecsp2Al7M
dp5IOnSMFuEqOh5U+yy5o6xSxerzweZTM5K1PFb6GJvAQnpEqmKBkg2UQL8E0TWjDw4GOiohP8EL
C5lwIB+JrndPpSwBxwdUxeC0HJrSfqNY0ddexFNqKxTvsJj7fVe9c1s1F4IxarCEebiECi5deQAG
KslOELg4XtDCBIuJERjCMWrd5qgFbEzmwqC9rEu8p2pgxQ7Dsn9blrO6Mli5wWhoySqbitoJuE9f
YGSqd2QRcM79q0qbsnOLOG0i9uLbUzRHIZsnkPNgf4CCziTaHVPOtXE4BzlMa7AdAdhLax89g5AG
hu0yRis0VGaHa1azwcoz6TWQATFZ1rd38n7k1uu62ypi90SNzsvDDA4V+WGzrrx8+5CzsrErC6Lt
jxWATqDGTa91wkbCEpYOSrHUifI9RA3nII6B3YoAfZ8bERBxWSQ+8bOI6yuuR6OJpx74+fiZ+eXM
jYv2mXoVmV+7ZIE+L6GakUr1+SWNSFzmHbglHxCGiGKSSBoRivaNPlOnrcdMKKKSeCp5he1uMpgx
D10sMa4VKqDWlBb0gX1si6AK4qJj0Aqa8faU2lJfaaVCcETIEFBkNfLSYysMDIJnygKJgc/QGvN3
LXehuTvhpLLlb6nL3ULK+xQ+VQ1l9Jv2zZki/7bsvmm7LP8Bsk+PukBnUkMAVKa/c+MmBVmaVIOd
sEGOuoGGtEZ0/yV8Jtg95xcnbsDz0oD+AIl3VoxHsIa9PFgF7y5Zvaps2kDdsUu27DjFHccf0BC3
2Aqi+yHfuwaN4BFRY1k3W465eIF5DIy7yqC28LpWKrDLdy6Re83DbRrZ/E6ZAFZ0fSPrbbZA5GxK
nottnWTMSG6CTxNDEJMoU+lfEIVdg4DvpBIWG+g+9ablpRDYvvzLPvwC4RL1V49beZ6sbiav+1+K
GFEagf+v1/Vt9zyj+jtkbjkc8ShZoGQyFAQM0Q7CDgFpYG+A6U2RaKn724eu3kNYK97nbUZ+ApBy
AFUEQinEJCaSvAM3nvflKSP3SE7Tj2F96Cnz0vdXdJoISMq2Vq9ELhk0b8AuqCBrGxne0OhuO0sw
zuudB0zZeeMT2v0/KRppzu90pZqsRuGDNYd8TKaagUsflQvz1f8kfazT9m0W5gcUXGjxPfsn97r9
Qj5IFSZ9sEq5NKlGqtprQkCY3zpOy+JmnRPldwySYBgvLScKXOjYQqW5ovwtLB725DCTOTUV/JJN
6OgrwG2THNF9EtRzxtaBrfVkZmv7xt5xuHbXW93ZnIzypj10UcBlNy/LaV216ckoEc8LKzKgiCm2
KxD3BOZ7msWywnXBC73SEv1IR/YRu4Xnptetog2BjlBv9OG36iaVZfffWNQ9dZqHI7b7udyHjn2R
Zca/jPutpv02WP1mK+PpwjUmeO3W0Jaosf92xAV7kBHynFwF/ufRkqgNzd+/tOp3xvThQ/VZj1mX
76/1AUfBml3RD0O9di5oy2DpLJnMpRZJQv8zxU/qA7FAK7VObg//cUGFvb8pRmY7FI0+yrVq0IgN
V+6Ur7pFZYIV+8uUC6z4FzhAdq5RadKgqnV/Xia+9gKZc3NRNe6BPnZFFFCsQx9Xe5wQ+0I2+3ZZ
pM7QMTSkIw5OYccC9cuUghKX2gYbZHVyD0TCP+GJXybz7ErGN9/GaII0NA8AdLPUlo23s2c7QVo9
zGiw6cThNJai/QlH3j0JPywuEY3WOp4Nsr2qMPvDokq2cp/fo0O01SNRWpZ4RUON/wbDI3aIVt+3
PFI7yWorNVZiGcrFWNecuMGiqH7WnqwZI1r/gikuY8CChVosVMOgXpOAq4VaiHor1ZQp1ffToWBl
NKDiw5tyhec1HsQdN4dFbQWo2EYSnhZpsb+eEAExrCGlcu97ZWIKNRLXZxRxhbtK9wmlZDW5mq4w
hpHl/OdVERWdyqjVdprAjT4kF9LQ2O3mLuA90Pxidu47dNZWqwqRmuy1+4lc4wKTR2y0aou2fEIm
fwGoP7mLgqZKdwvhLgAOcQs1PYIDCuF/O9Fz0y81aGayxCyJcUyu4wrTLE4j/kE9q5fXKpEmuLeD
7JpZqyl4bbgoXgklAKIPRTq7h55TARAieDIdaJ34GFjux4gLeItDSjAeiY/ClIloWZ4bJXbPGhN1
eQIvB1RLpI17SQXuMpFoxCW1UAhazs3URZkGmhVAmDtgeSVLWdJTqUMhMbOzn+ScIHE5aLuTwjG0
aJDM3Kk0frpnAstrLajc1fLjaw+f7BY82IO/6LXpXY9qCs9FRdvVStvQ2v3PHpM89uP8BrNcaVXH
Xs9bUtmc+zbCcjBPH1MziZC89PKxb1BnpZ24CY14urz9mI45cIqy4j3hlyi2bCFwNSR+6rj/YKXM
R12zPQVy68ysidsJ5rxAZuWlvRmLnoNX4JBnu7b59yV8G8dOusXcJF2+arxUGrzRRgO47wk61txF
xjGK1X6lVUBCcnNOkPGVZWnpdP9vIxUqmC2HPK3897rca5XDV7OGxzTiLDdCbc3gaSi5Wh6PrxHs
9YlZKKTR81hHTFS2VdS29MhopOT/f9kW7Xv1iw3yUecOlU7LSHNxSkcRYhT5Vi551j+JplDX785Q
hfhYwMAAr76QkPjt0IRR7PqFfrHLlJZGQ2ZASaeFcaG05cT3M2Wq0dC3IiPxEpZv/abwxqaZ0QI3
+ilzCOjVbc/lAZxq0rTeggGVfDWkBU2KTgBMqVXkVdR0Qi//RVY8rZOmk36Ewu/08/fEIgl4D0aY
3Rry2+NNLAx8wpkz0H7igTRVuZKf0XW1w03wWtOCUrEJP2ebH8/N3O9Spn770AR48oG5yD41jyw5
h2//BhHqBGZz3HnMroOJCOPgo74STEbOA8vScpu4uJnvDsc98Il/xZfp3ZxKyBpUejACrk21eb+N
ARWatLGCsUJO5w2FNZgERnJYzli/VNOgZVzsQhh7cL/ZA31hAwzYMnitMAEWmlN6PUr4p0jNEOWa
1DA1N7/Efx5NrKqmbzymCWITcRpV3z9uA+36swW9HdfYcq0/ncXYyFk8or0aMZvdiQCBA3N26mub
5si6aU6cYizoENneFtuCfAc4tUBWpeth7JspgIZHRyINSXY2Ck8ZfQAoodDDsQiReKgNlJvspS2Q
0fiXQM3eCDd9GnPvXAUp21A1CNCoZKXd4fU/o+lC5iwbMPsjtleKh1wR7yar8KO021JNngfRELGP
1McaOfGxS6HgxNH8LNXmMICD54yS26YsC6E+2zVjcOsrvubAwtELyaQ3gdBU9mYyyJyv0ActTpoj
xg5QY2uZc3L2BQizCln0mhuUZkC1/Kl2Vrf+Hba5QowX/JX529092kqTV8iSzy0oS//g/xnPNGvq
+avvVfbZ1xKaLgN+tIIfAI/YSVTdEEJEU+OFRlU/pgyon33MJv0UjANm93JdiKV3Zzv2ul3gRZPb
QqRgCzpw0qA463RBj7PxmfFUinJAR1qShC+8U5SLx1wFiKES8HYNQWCMErZUfoPRBDAJU+1c7P9o
m4CKcUkV8TAEpy77AALNVl6cINBTENaPuQkyAkqNycMTxTmR/cVPAokzianLzHa+1nbT+0nvsQ/y
lqzST95V6xn6WeygsV6vV5xsE8G+1BSONTFuaD+j4KifAKgSwrkw5Vo0oDDF9yv0TcDHG2CIoTZK
4fJcFPmoN8zKxODWyZc4QLb3opfIX+xSW4QD+OlMo62N7pKWdr+e5PQs3rb3GDjRKuHAc6QCK/9q
0FRoK6vY6p7zSCj9ZOxceIo5xfj2F0ABT3BwZvXs2IqhNPY0DgeeUowZUw5HHWedT1ik93fN4QKf
mqguSGDevHJ9hy5baYivx/YpvCftNMkOBK29QN17tH8MNrmMB3ojmJI/SufjRXjOmQeEMybR9PJ2
0+hF4Vvb+FiJZJeRmpI9brzZqX3Pz15GspNNS9I1HFAG+vi+YJQOwR7OLC4qCubbNWim/Cmy0AXa
d4ACs9LjqMCKFEUHrwE90cTiK85Mrya39bsqrYVMGT1lSsgMrgvNfCyxhfC8ud/oZP133fdmIR0f
LZ9m+Q54D9nqxiPOb7fsagxcMtBtVmSV7aZA0SW5HNJsUJUqZI7/IPcvKmo7qatKS70lAJglw1My
qsDrLvWlXiPvJ2cW/xemHqmeUHvoaNyo3XBg/mBoe+VOzKU3UVezMfc8BHq0Y9sJCKDEkgLsCixB
Ec9SJWar5YY9SNioe7WK6j0hlizjWJc/ipxtCamtGYeYG2LsXIeJwXhE+NO93tFt2VnNx1kGLZjV
H+tOZoSSrDFuqGugT65/e3xyj8PZG66hNZi1OXCG6IE+M2yj/VapM7+IT1ff6whd+TG7zbgtBBpy
NRNbIPSDzgUappBKeTk/yoRbMsLFKHW6zVtzH+jYkuHi231XNuPxnGhZOyvQeTt0J6AbypTLnOjw
Ika7+ZQ1jVSwq5NqLhO0Ulz5GLdPgzqxzC+GjFAxECwQ/uA2RjrnJfE4HE9dEG07QrhgHJX0Ngvh
82O2u/uQM3rbktPN+NmlXhCsnUIfqqzREFcJnn9B9y3A4FohKRUUnhVSfzafjfXnt8qYDEJSp6GY
C/iAWcN5niXyGbBZf7qYNCb0DXhc8Tiz8J80nmqTtQWCpkRomQNpGD/P6W2ixw0n9d+bb8jDZvzc
q8ViVwyRmT8rXOsu+P4KNCjFHtb5b92nHY3Cy49ez1WJYHSilw2ciqmmvzVxZcnz8vTupAg6YUq9
3IHfMHUFbo0Iq+wzHTmXx9LAg08SMkoql+/fhGq8m966p4VUdTqKUaUYm5im1o3i91n5EwEzX6l3
laabDp4OAooNq4Zat+FHWlwmjeEuvSRch2yY+IfT/JKuHidk5PtndSGfBwkG55zRTzCE2x+zkVX5
hllLFMPNOOm8r68OWrrb/g+y85/Qa6UF9eNc/jRJkwS4gC5wDoWfjHbWBp7Us/SV/ilbiGblKxaZ
sWI6gDvZDFrwatMdAdC+jlvbf6FNwpWOphTCJnUsdbUzBkHf7Pze5lYT9aSnKF/5rlBqIBM9Ul3d
uUNKqEuGXFDHYPMkQokFttPe1HWlGHxq/Nt02k7z5Gp/ChHh8rzyDJFS9dzTx2BQUnNCHz+V9I9V
/2XPn5x1UAZRLkeAS63Jl54DR21rNqxnzwvTbNuWYE2cftZX9Lxh4qVPZm7bJorphVI4jXWyRPye
4Ux0bHnAqMmbz3PgFBEo6u2hdn60rjYwqfgjENazZOPI4Mw+cGY/xgo9K9qDyHSrrl2kkn4VogKg
RwDHsSdtiteCPZEiaojovzxP45sRFoEWzS/lxxcS09Yf2Pma4JjUiQDu16sHyhfBx2XlWSnEMoio
DRvlSQaZVdqJ77zOlXn4KLBZx8zKtcmo6vjAUVsk9zXq2MC5CmvKerljFrz1eye8rV1IPxqQODJ8
/54eFgZUkL4piR1nd8pqUF2drtqJlHddn5eAH3dwvgzfFEtZ7bJ37gRt8BszS46TFxdgIjHRT6ml
pIITH0LnkIKhsoWoEBbQWR3VJVs8PuQhtExJsVxeuJ8Eriz+M5wrdyatdyv3YTKjf8R7dg3HIprN
lLvdJuZDVPJCRmwbr07nCseWmWKslr39StJZmCyyU68VQDllFE4c+noVz9L63QbKGlD0TITYhNbi
SEAPisH0TQ96hwt1Z9hSTrc7EY5KALj2/GkxqTTP4k0Sgh/TZN38qX6SCDj3MNMIS5n2kL7poeb/
QHPw4Z8VNsVqFXlL3sOQhTPuiSshKJLbytVgWklP2UuiyRHyEKqgs+MWsBhySOnvveqcYAUodQj9
2SwYbubfyGTj6Z/6B4EX4Pp/x0vgDL4IjZZCZMULyYOoaGUt81axvLUxgX9A5dc05GZiWrAeoLuH
vG5XfpXYJb106UApFRLpNzA9ec6ZNP3/K83RAS51l5sq2kkRIwxX03yde26zXZp/pKOuxLdtRV9T
aLbU6zfYCmliz0qEgSqKE8nRzInxkljD0b/ax0HEz5G2lQVxJ3yIbMb8MCvdU+2+s020Zcn61iAf
OQmzodyc8Kyc2NB+LzP693W7yi7I3WBdmVTd+gt1+/8rp8x8KWqNJ3D4F9JO3L0V07Y4atQL/uTj
/wG4F+qJJqlmuzGcmARSWzlvwozDHzkOcYJkRuCGq2+t02ggo/tCl/tdlg+8uN6mnOk3VvQgai4A
rFbXGmRsEYXY316xzDeSdo528lDKAggTcG9YON4bvnnJZo0Ph1AXsBSCPqBiXQtHmtiC/2uCY941
VdbtHZAY8mQRGC8k7C6ANYfMghYkQNazMTZ8gPivAdqhB3xcOUi39WKObQr3gtroI6QDqs1jRS8Q
PVxQo4jKrig2pE7f5FrrOo0vX/iDYhJYDd3x7HJHxydrPX3hDE8dgMY8TZPnDcPTUiopMI9hsNRF
yOTmRmO4G0xY9BYQfENM6eD4XlLs4oQgSOsrbIsDkZPrE8zBp2hYY4Wy0xt5TOoo9hloCadEG8Rn
lnDl3LjyTyHdfjQvkT3EUw61QSB6eekTCIM9bninTFHVreioYYwTnqO1PSZKRVQSRoPHJa36Cmci
rb62nP3+dyhst8GnJss5UcUxoU/BjyY7U4CCajeRlohczC4wGF0BgUF+B42mqwc39TrdXrO5unTI
8TumS7s6kke3L1aafnJ8lpy6aypbNZEvuZYyMcE3dXc3bah9kMknWWcxont0UUkNkPZ3bSrrv9QT
fbFN0X8Ox3WwUYwntvzXxZxz+lYnlxmB4frArZWYpIxiR9hSlfbCDTYkWbkVqJZFsEEPa1Nq8ps3
dGro7a9Y6+iiNdO13/olazPflcvRmWu5i8XA98Xb00ZgAkr6ixyWNEeSaCuvmmRzhXSCgv8Tf6u6
FDNVOt/kNMvnGwbx/IS+uMPpVchgw0xW/65UrCPV6+vaCjjP7+uSk8SdxPRdYxMdZheux1GzAHbZ
pjBUdGMYXltUFC0oBCOC3Zdm8tbnOblgubbW2EAkMHf2HEmLQ+Y0DAxP/hb625UL92soYRGe+4oq
FrZOC3XNcl7lS3UrvelJv7zVwLNi65N7DuwszB6HI4s8QF3GaM5uy/m8+fDGye56Ap0vAo0moYBp
j2rk3W+bL+amTLD/FtJqPUXYXtl8TjpQjS8Dz8xE3Lgmqv7hm2eBe6VZ9EW7mMbiz1zVmsD8Hnw0
DCFEtHbGfWWqFzACPTVXSef56J4CtXu0YkN3wjxe+gg1OlGSeOBi8uob6JfJg3ZSbhDOE9o4FHCa
10f/6+2pHJhoGAUMEOxc/WiLsqb1VtsE40oeOms0/a66WQs9pUlHbjr35GKkvFMCDP0HXZpqqui3
kwQzaCjVuZnVy6b3yIynBruEk07Z2iMzCMRUFrRJFH5Wx+6V8tJVYf1MytUu+i5e2WWS+bVBz693
FB4Kbz4oxsLsmqHQ/x2AeXvonauv42WfyV4E0/4chvxAlZma/pUZFFcz4wYJQFPX58wUdDondqzR
/rQTmJwh4TaN37Lynkket7yNRyr7BiT/nbSzf+aFkNhxI5X84gKDaF4Rdq7D4+Scraxvb4LyINJ3
yyEkiINwN7bOtzqyGR18VRftIJ244K2/2wH5saluzEj3Pl7D8+mUv+NI+E9EnyAGyBq1WKBk/iRh
PsqT/XR97BE1lULIAeD9isSZQvzdT0EVgOiwinpPzeSKCkBRe2oPGFyZziP/rR2Hv0Rpra+VjnmD
RNNWeFWRbQXoYUqvTzBRqVCu8wKiSE/5SC4SL1ynG+zGtlKltJnx1Pj2NRrvG9hUvXvTzFj2iW6J
ylN4bHQunWQF9+XwrIX8awp9OxoV2iRs6Krc31KsWmQF2gPofU0Mj008gZtjR5sfLfG5COFgqj4S
pTfou8uV7E4VGEqB/iNk3ajZJ9QBSQik1Lc/Evm7lH7Xm/gs9SNktko//kq9+91yF6QTrYPsMgrB
3keXAMcBBUGiSGg7mT7TtPEovp5DFxsUWhFC/VEmIAAP7n0cOgd2EwkHdHDTz02ZchAB4nzCwixm
y/ETl27KudFBI6ZmrNqNz8WsfnEZaX5TqKjsSfPwwJ/MNEKElhpDD0At6lKwfhpfzzaU7Ke/g7Gq
36NIsmpj9Ji4GF3TD6d7c+2Kap6Exj8gXEnz6gM2KRQsmwKbxDmIn6Z+d07RGyQr+ZXaBnnRSY7k
fwsRynFlL1x9IEWCgit/4L516g4ft/Cev1+euUXlIVB7BVLjQJROoGlChEAuKaCTkpuN/4RcHu96
BQ/m+zG5pRAczgq7l5dHfab410QZPZqXJHDrCm3K5TBufU8vbCgQQXn/6Qpxz2JaNMHDbCyajjwn
fqNtcfBgWiL9r+59cSO0nIEYfe0T+iMz2XhTXZPi3fz89pMka9kGVae/1P4mMWuSeVBiRdjdvZYk
HifkACEqUsgWBPV6jAlzZ20Nzjn83mbAEuhJIcTLV9Bou3cG8RQ48jANlbeYb9wd84x5SMZW2/NA
Dx55RsgxBc5+hqDAXElfSYY6xSo4rFnu34eWjz+5HbKV8O+tzsVaCvCpRgljc5odUApYy2LcqPnW
S2qjxx1k0y8eKYGawG225I67q8q5sYBbiclUVKeoRE3vyenYHFnzRrSpVGhMpZzCKAXZg2IqFkTv
0VAiNkdvYGGwwnGNZN4BXGW3I6SVJCaowFoRuZXvVKy9j0ACcbRgdyXjBbtPOp5yfvviuCtATLMG
wcIA4+bK0rrtXs5Rf1em14WHogIlBEZgENx08YDQfwnsBbEgu5IeGMhFz5wtvly7t3WG0Rk1rPj3
otVjtO51KwLqXP+FLp/v6jddMUlr29m6BIxYrn4XTxGQkQQxUAxCHzbPYO+tKOyuKbvuU4t6elEx
W9Kq1RNTcfMTvEJm+qCEMtGu8WsOdlqnSXDWyK6JXaqQAUHYSDFluqDIJvCRk2GKCJ3d8Vb2I6Gw
EXQvbqCCFo+YaGXh74aGl0COIPszitwUQDbEqy8bZjqXxj8x0uej+SMBNrZqHEk23N/zsw1c4IXL
zA6/lK1JJBu2mj5XlnqkU6IzZIiz81li3t8eekw7VGw5uI2YVp1rfAvKJO3Ik1V7zK2P3CFtTBQ1
m6bMcXrv3EnERmCUMyKTfiKarUucf4tGIS+ulalXE+n7WbBPpZ++n6Br39XVNbrKypCQ8A5t55bY
g5L4wFe801KBBS7+zbK1ZyY3iIQBf9RRzD3gxp0nZ07LwhJNoTg8R8+zk/M7x+yZuRAKScss3vhM
vsvVGfHkkibGv0I8/jFJCb4m+Fe3LnbiBi6lJtKJnyZ/JX70oTYJqkn9t2n76KYSYa95UXZ4sxhE
xLCKNhLCQPNaDuXhANVCJPbQPitlQyp8nFGc4OvnkUDd/H2AY2H3xjiR2qz7QYWrPuZPMGdEuaWe
yuGW1Jr7gSGkr4LJnsYhuPHsIcCJpBfJpbJFysTKCB9cpC9GptsZML3rNbTbA4THrzESjqb8l/nm
5TKrfSx0FRJ8g3r2mydcUmTFg+n+ZJOLXGb/Tk3uVkU6tskA5NALqIS6gTvQCBOkse77V0tYH9LW
XmSSgpOTF+b42t9q/AwKwSXaFNdT4JF81Mvu5NP5C/7bg1+Plus5D71U2ifmIA9hPWoNtyWYoCu8
yUX9f3h51S3pUTuDQWLGM/W8jy/dZ6iVhxCbpaPcAGAr5tQQi0cssM6ybYdMDEWgyM2MhaaouE0W
yJ1jzuzimTmCTcYInMFTGMn51H6JVZK7pxhhhw/T6u7wwEd7w4nWYQjfJGSIkUNgC3Cv0x61KFj1
eJOtua+7+Mjx/pGTRaGNdwo1lgCDnMCzLActtVm/sxoYMvkBVaeIjGrVAj6AcxV2jmF0fSlZ4hMR
Gr3PtMQAYMOpQHIuq+vRTCgXE4B5Lkw2cVqSGm9Xs+S/lvQHZ+tr3VvWl+lfeby7yH3PlV6Zokxw
avdk9ZbTlEmhHSqnSinyl158MFlsvn6frDIz7V0XIhRNgIEyWtFaq4LIUVLiZD74eVOxqKcjEgQz
9Bbuzis1Ls7V7jJ7sFi7cTg/zOjaqlfZx8zM668QUT1PatAx7vOPlWoBpiQXm4vpuVDLfOZ+6RZj
CFyV4iE+k11abAGZy50srHzd2z0C82n4MLdC/s7BhsD5AqrrZwGsoyTnWZi7v9i9H9IyEoCMmPmK
gtik8XwNhjT+G5YNaRyoh7dUr/Xk4VmqUVjGQ55Dn/ZwI0oh0/AdkecK5/BttTDMppIdgZ6NAyUZ
2vRIJxv6XurFF3XQ69ISGH8EVBaJcSRWuG4r6hAeKlpltatKiYlxOQi1dxIDbr5EUWF82hWZ+zvB
5g3LLORkjCosR0UAwbVMWj1H2UgjFe+7yuOMVSgYwbzPkzED6s5vgdh8M0UtLFhLynHMl81OIbZq
HYp1Q8lsJS3Cgh7/qR39BalCekEYw6XoqrvzHpVIVlG4ctpFG5iMoDoi8uaB5ZAA1myTeFgqGCHA
ejV82LWs1QdQV/xVkNPA4dJzYLzAZeLJGOiCS1N8SPrObGcqq/HJqq0+d9dLy9106RC38l+P/F8s
2lHvLxwzfgWkUcSOkW15fW5Rd+DvscQv5utx/b0QwEqgCyCMaPwfowrptle19MMrlzqZwbwqg9ly
7mSzDnx2yR3mRCRrqavwGnLyie1ac71SNQgCs/vpDmrUmdM5eGYtWuZIw3cUUtH/G10KrBHwRJsb
gNowsJI9dMVGGaq1FIHqYZ/zqY7XSJhfq62gYy1T0EU41ecmfRTcpHGB1F2avVRFYD1WHNNM/0F8
tsdlwmTo9ryMLuyPPUABnlGNMIW9HXDF8DcEUJIvmuZ1H35aH+rum33W8IFbSysYcfy30F6kC0Gd
gANzMxKO2f//0gFv0Sa7zMMvMglLqYYZF8/KTsZlF4sCUBP/wlsIsaUWVW8+DljxgVoGXaF6MY8c
gQOAVadhsJFlHEWNzPGjEQAomqolgheGLpmNfI62r7hTEYVAjxdpclXl0T1m4xVmpqMVLFFzVf16
RL4MNLQG3IY9hrMp+Z9ywNnTL+LxwIS6l+4Uf1XNsXek0kiZFH4WsbyiBMKIdEumXQkPlocWfs0N
L06g2AejL0YcpF7zxNFD/R45wHi6uMhIz1wQOTL02/5ViOvAAKckASzEisxACjWLGyLgxiLnpvmt
NfBVsZeWjdgHsZXuH5hFftsU7YMl3PhLMjTDEM+5wMd4HbPsQHGRoiEkhyERiWvVkXREnW6mPuxz
43XYw3nJf7zErBznV9/yIUbL+ZahXFZBDspb3DSLPo0krClM4GefUr/y4YYyoAr3Y5h/yJggl7uw
A5GnO0HNBqR6GZkxtARFcpjM/b5eWVrnqQieiJ0uQrUfzorA41L/oc/bllWzIn4tkqqkAeSgFyrr
8FnAvjCAw88Rh+YRp33hAXbBSWUwrOxKvvCf4yg7FInD3DdRkKgcUI2iVnI/cbF7DKKGfNQgmgNm
xwE3zC17KpYUS5cLLYvsLz49ZHsjvq0qvy0eOT64uYVxX4mEjT50RuZi6nx2XL8ma02fh3CQ4EBA
pRt8m6F8B2Wn6DqCjaCoKQBQfPkIcfQdeQBSkX8cpxOejUoSdZ+dwzB7XES0L6uOtuTU/RvU1r6J
ULJLW/0xmNZPIatPIhrBrcp05i/ukXPCZuNs6ZPavft0ngdlKOBpzMUq1HWkpnG05ZPD0B/HQZhJ
zCM2T2O5Vk21vBJh341wXhz+8tEDgP6aExFGPEgGltcRduRQVhG5SJ3Z+hAEXvcW1HJnMe/Um08l
2Lwwr+7P4slbYdkTxsESIzMOUUVKmN8Mc/wIpGGCjzSySiTiUiriMwe4PboTZm74Rs3R4waF1pJn
vpizxqLvsSBHf0QoDHC89KJk6PKdXyv/d3I2kPJLeAlWvUs96Pl4SUNk8FUztTtms7YdMHpUbgZL
4+IZMsvdKz53R9aMyIP868zLegKf3dopcpC0j09K5G4BtcSgmbd6pngaRotx2N8KEUMiEoEW2K3F
1+0b4QtdtWNmnzWAESkvhLhEMuWLzkfPF5HqOemCLjl+jYs5e3gRmpqQcQPz5gRRFsgJ8H2xF1oD
igFeBC3g6yH+B/CvWuHFJVWCDSYscZgtYxW4tAefXoMHmSbXawEHcmln8h+p5uCnPa2dMJ/w1r3A
zF0sgPpqVrqT4k+A2MX/t3Ltnwn5NuTeYPmTnmZpnDyOySPb+o5vg6toeVUfqjjnnmnXQZK/5G1r
XuKpdSxqw5qZvHNt20CUL0akzfrOKEpURaxMro9+UJX34VgM/UFG0WgxoejPT6eXhJ6ouuU4Syrf
aTV8rsEIbzI80p1WC/c9LFNOKwKwVYTxXowlu0WZfNHnJMNoEGi+5jM/VDoccXiuV5Vay6XF3Crd
eDcI5yWkaf8m2ntKBoFi1AzEEnPS7HRxr/PcWUXPV7B7yX0KCB2Epwa5d1MaWngqgVrqX2B9zdFN
hDdZhDgTJp2gW88p21BIK0HWfEW/ORLSaBHLoRRG6obSo40yjy0sm4UsXNZuuxRIiTqjBSpXEOmI
JdmzNA706toqq/wOwDVEER2GCuuk7dVXAqOaJJ4WKPeys6NekV5KlEIl4vjXAXAlTJV9utVpjT6U
DuoV++9Jr8dj3KcINUfkLG3Ceuk8M3s25P4WtcQncNQso+3Xw6spwxA5POl1w0YtVDvtOoCxJueg
tQip43Nu0Sw3h4iRBEvI1Dx+EVARujO6/5yMDXCfLyYh3ooAS2x6zMBKVL9FvVmQ2S0S9mTqK64J
F8DEws7Ld3hEeZBbNAX8AZ2USuxfez9WGyJijUFW0/U7gd9lMNshZhd64LKXqgVi0fu7fhUDJoH/
TiVqFCFQ8Su7/Sq76dzYwPIOInVYPMj4Ji8nqgqnIK40Q6lM/fL67Kbi5NN6cXnxpz9rkDvR4DR1
gfMwZ3s3H4jOuL9rrC4by/WgbW3X4JoOAt7YdqcvFan2RdMjpFB6CV0zNcjwI8NTot+7Vi3Tw8Aw
BtTirZCt6XNiEGOZuKRTVeuKP6+f264xBviuQFNT4LqiEWX/uyh5QiMhgJoJWrB0W2flB/RIBHqi
hJadYm4XC4Fyq1qYPvyqAIit8s5zPUbY9NXVBBEMXYGRDdwCRP3ww+ZS3OJnFDfjqJKbRx1SRz1b
u6fmBdMM6OAuuKVHHjotREBaYUij+R8oYAidGWXRMD8Skgtqo+hH2QO34n3Yo9R+r3XrtIIHfoVi
DYkwHLim6OP3jCYckcAexJJbbjwXaSmj+fwxFUwX9RFbtkARJib2COz760rLXRY6Y25QZ97iz6IB
jmjIf9i0qvhGR6x9Q47CYG18b8NHOWB+633g/19Dq45f7crQvyhFIfkWdmvYJ28LWI3N4TsRRMm6
Kx3+f7PYZLJnDEdwW4onC6XVsMYyWXC85x9CzAm79XAKjFCrhVbZOAz28TbWSf6kwbBHKH7aBxM3
Dd/aeRQ1ypXuE2OasaWnu3Hnh+o88w6+u4RUmcDk8xS9bnWmKHZEClaSGi3+ltptzRu4oz++m4Au
LwOg8ADLiQhN7CinBE2rouVwlKkITi03TvOQwqi9L/7BAiP2gYQiDHe/WRU/ALCO+zo55VCe0d6S
0jHpOIXXc9oAIxc/f0LTl3w07MuHfcDW3dlWRwzA0twW61PjwzD5GbUv0YqRho3x4CrNNp9IMKo6
MjG+PL/68oBi2vELECxniihMlgY88riY7F1O+SoOPs3Ix5Z/ocS76Jjlup3e7sjyHJNEB3NS/dZE
v80V0XPFrPFqsKb5vRIrCq8lha9Y+yOoVHr9eW0zme+ule6D+0KdjeTyKD5uCkiCwjNXb2rbzXoM
mOzYaxd7vgaf98SJn1EvafB/DWt/+lecN6Mk3+OxEejZsp8HjWRO6hUUfRFSAykcT+C+NjcKUutW
jlRkd3h5TXh3PdnPzeNmjR63thK0WmWLE7XI8PsreZhwzlHpzTF/zQ72Nq40nlx4NSlJJF4QmD+c
1wyI32bAJ7Q9SagPjqwjTfZuH+RSFjmvVIFki+qSk3EqQDmch+cgko5ym6pYF0wDpPN8Nl4wF0Iu
vqpXlq330cKiuO3mSGmDcK2SmBP/9mW1xIN0Wnty/suPLfePBaJqMk0rkthxx3eM1Xhe7wMi1FWQ
ZlHjwqmLIf/hB3i8kuZNwH9KG4fZ6wYh3+6M4tAV7WapM6YTVJs6n3pvUFUVxz1sbEvh0QPrtFOB
jN8BLiQYXn7nkj4tdXI3At5PAzd2TMsHRCKmmppdg83x1fHNzdLRnenaFQ/ZqYUnbKq8AgFqv9Ma
JXGhv/XqhMdSBfeDytBnpUdNft4zfHvb1FlWew2PSWtRIGAGQkkQCHpkNTBCSHvOIQToXSREt/lo
yf6dzkgf23RznJ6p4Cmvly49G/+YKbA187UjodFQKuS69aHHek2xGoeofN7jWCZiOxJISLt+eclA
5lvLQCkMUezs9CgFUfCX8P4aeza19HOfSGp0qizb/XJQvWwmxD6YB28bZ3OPBOu1g1ieDyp0mI1K
G2/BN8Pxh3Tw4m78s6oL0ecS1NjkW+wA8Uj+vpElmGJaSOvVteKRHMMoCOFqTT9N5flgGwXXIdRm
k689I3oyIOoXZrkpSD4D34pUyksvqb+go53rWYII+XLg5/WSiuU3AMijOPToWx1Cpl9g52lbrNFk
T+zsRmHD4eYrPNRHOhF7tq/MJZ6TH0Gh4oxKaRoNu2AVAG58GjB2YF1UTY21VPhRN6vh2OaL5A7z
qZ9Q0t3qNrVq+LZT6Ee7W2Zuql3IYotFDLNycB4Ijt9ptSYbWWiy4kG6WILib3kSUA4OVWej+qB7
328p8WNwNTxBcaHsC0mkMZh5FiACOKhE4Yd34I2VAeHOXM7cZxfJkwSiLdCljp5aRxMikrXsCqS7
Jh41wLQg97RH+iRs0GSfRXktj0HVqM3tU+GP+RTLYOn7uSJecQaRWzP5Jm8rpH8VY/OEsSsu2SEU
x3O8JWkcy8p3q9Ke6HV02x7ouPHbTl8G9KIwo0i3eQL50fjeDa1YcUX8Krnfpmu/Sf2d81dDbwCD
eeIvZ3rRJjJ/IaLzwgdlqRk5o7deXKVh6x9APAYSbbQ+6SwbJiroIInPTJ10rZjuRv21WjJSlzSF
7Zk+XTu5vmQ0vwOMPmdeSF8M76j1rEQJKdS9sjYQTRzcz0V7cxKEwnbYMNu5Hb2irAnGWDu4Op4t
x3fkYaD70CkEZjUY6vqW3IrsClo1VCGezuLhmM2unUGKN3mxuEUsvrvlTSoZh5BmIqscxUJwlZw4
7+H7WKmvEXhFzIvJ8txmL2Keufck8uG79iAO1fQ062EYaZEFehlZEMWUr1N8sCNLq/GKKFwfQrUJ
mI/UQSS7ZheRkN40/dvUArN5iuIlvRBoEpfIEX887vgz+2x2+uQCGgPnrhOnlip0DAwpkU+e2sNt
bMTCyHuMWaf5IxoWOG1qgyiQEcZcItPhNqdWDfV7cMD0JpXu3SrLSChjleiyTzFybu+Uk8IirWl+
QKo2WkGw/cJ+j50jrJQFbpDnB2WWFafDlJYjJXY2XdK7HafvfClOTpKKCYW9vKZf+E+vrhSHZcPC
IEa4OHHMrd8Xig/hJ6ubibelcafp6gzer9rJGDAiwf4RTgwxkdPhloZWYlJdPxS0WjpJ1IRy7K4z
NZ+ol2vY2feHajRcdXbn6I28feWies1gMoQcJxWpxwgrDXT+OWlTvYlIEB8Y/EBCTaV4hr4uICkg
owv6xMb3lWvqjtSbl2AX/a05mZdULnjm7rG5mrh4cBDqIhNR5XwEaIZr7tM6dY5DoRwP4adp7RwA
7lBHXU8npSbDoei55URk4wUX8VFwWcJa5kVssnsAb6o8Jbol74XipjNOYz4oHxH7hf9+LxhFImEh
+QnSYXoO+WNXfP/YnHRuz/W5fxEPjxJNSpwWmbjjyr+jCwymDpSxICp5qycMh5w9HHjwHRFp8WvB
Sh4N7Tt9OJRSWvvKK8nO5PbEpLhOspYWxNA2r9calux+lamv7gWUIpgayS7A2AWybCpFINmTrkMO
EpyDeDqb97ZlYGzqz7O3BlEHOdiUF0lnSiTGQDS5Peq6BKtkreXTCCPVIEJcubmGdZ0wKwtQoroY
S1Q5P0ldGSXdEqr7mfNmzSAoPXCSsxPemwJjrYc6zkKtXWGRFUQ+nFTFZa5qTmzpJiiHvWv8FCCU
2fKcmygKDma6SHGvlD/uMbCEhDOrx4bipDJIvFFNkbbnq7YhQcHKmjDFRVr16fJY74DZVoPYhTJc
CBCSLQp6h5lxd3Sz9NmxHGVQrT76aahbD/A5NiCrxyETCfuCwq4Bo2PvVZ+wu8zQ2hPsjQ7qS/z3
bk5P2GeT/33DkiWkONT/ZI2ltdayzBqgjfxFqzZAPFG1ZtcJIhrnQDSMaf7WSYGC6zg83dxx1Scy
X1OFsg/yGwmi+WH8tKeqtt3rcqtWsz3LBPxiFQMPa/yVyXhw6BiUXOhgZTSI9B85GQTowz90yQcZ
Rxq2WuFgY/QUmC4yuSpUXyTTQE6Z8VuU6q0mopy1xQC6wA9K1MLq21EIrf2aw0XooRq8oxDQrg4+
pI2uuzVRVs38TICheuYzbcTqp/SR2oT9aDia6li+70vHAaeejTz7X6z3E7fpf+AhKNomSL8o9DSz
BGijyfB/5UyhjCIY4DgTxSLHRQ6J7lc8So1sJluZcXjzJUCyErRbt2xHiaMR9tUP7DqyFotqPTbx
GLEucc3Mc1GS6+Fswaa4poDY9nKwp4WtR6jtS6saVGXMdj1q1XPNBsgnXEKG4f7TK/N8ISZ0NQvR
pFghIpA178lcuV3c7VGGLiEP22dBbNY8l3XE8Z+HSkSX46G9UjP2pC6x68aOZPszw1IvQ3DIgulB
zPLc1LObjprZwA4LbgNayf2F4Owk+C9MZxyyvbiqTaHvCH9qMtadOHiSz1/HDx+kKzn/YEyWufRR
FbPT+YJBJrFPrv66Lkl9KUaddykUXzUWl5wv3SFTgXIssjD6kPr2HS010DW5cLnFCNpl8oMMWL2m
T4LfPMuqX2tQI5+jDfYXAbkNBQ/59HZNQJ1oPcVY6h5lTnuChJE/CdhCGdvzVNt+JS1Yf1MSn1NE
ueWC8zWckpQk81fK2/oB03KpxMDU36G3E6uZOO0UI986kEt/Ertt3i6Y1pwwWBG3D3fWVloe2FFC
E86LmNw/t/Og4agC3nimnHSqZJ4FBObCA3W/XwW8oWXAV9wTrdmRhWVoDEBauoUYtU9HsP+1CS2a
LOxXHO6k22N9nJrswFdQlm+Bu9IGxqYexB9JbFUH5GjpxjlZc/VQdoStkeCsi8jQhrKn3+bJFWx2
8yfxa3kdfcVwfEH86ASFzFunr7n6fg02HqC0uDKEGqFrQBK+aBuPEyjt+peqxMXOhE6J/rKnkA0k
1evbLZ4p9Gs/52jd0JANmIVCmv761Cu9etJ1Wz6nKlKKXu2vvlDI9xNwyZsYanLOGUOrkb39z8Fn
r4yj20JHOShXm9y9l9ZULYZUusf/g2dKrZxzu99saVsrusVGRYgPcrFSWHqt358TTQop4hnJqWHl
nrIXaN/8ApyfRuDZJB1ZFJjWfM1vtiZHZT2xotwX5OkUI5pkTuwWAFSFKoKk8lBOdF4uVBLep1Nj
GXdJ/QqNrKNKy/8daj4BOfIyzhpHhQCsi3aiLMqI2YjP1lQtdb2UcgtTWBqm435Xx0rbqvxh5Ov7
Q0dgCzUZdjO1w6z2WKGPasQdSo7TLo9dhgIbwqCp8g/umWzpDZ4Z5HOxFBuTNwb7oYd+HfDMCoLj
E8/EZ1DHGnmbrdDUOcVuJYfq089mgHHpMwD2B6njq2xVY8ym1KRT9veAG9IEenAgFcnBp2QtUq08
N0EBa5bagYE7wuxTPV7BNP36kxO9cnvunQFCX+N4iw93Kgh1SydMXd04kFlf1yzgmg4HWQQXD9R3
JPKJhbVw4Hfnh06qACisqvzyRGqURoEGvX+rTBZZHQvMYs5N6Qs8TWkDXuhhHkIUKRM/0vsgR/Iy
3r65rmBJmrBUp6nXlJ8/iP8M8OrCK1DdfPKxXwtkqEBceAwEYwBUT8pB0KsFN3anHBKzGx4TaALl
Xcmww0PLbc4L9oNBtIVxrVdJnjb8uXuBMgP4TufX0T/ii8BE3FYOwTnDwvPUtM0BmhTZWffYFp6A
mUuVhibibTdiWvbPRHNWxRNmEcUTlNZrEI0uZdqL2HKVZCrZEKe4oBzOIHIamYG62KTl/nGEDvI7
E9iWnqolxmzOZfQdah8XWkZoXQKWdvOero/vhB15eXPFt3iYkdI+04m/iV/odSezkOXgqLJIBNf8
NN7PX5AHr/dXgZx+WwCsfaK99xB5g79DS88ui67xsFsPfsdJ7sYFEAXvmZ7gA7OItzMCkhaYzfgR
el40IZJhpBbl0gvQU6X+jMO41bnJ4qxCgXlIpa8ND8Uoefq5MJ5mgQSz5RoiuZp292ylJ3pF6qjB
XpSyn8+c/Qxyif9MlXjbbZE7p82YHaV7f/U9nMcJbXgWrl0mwT/lc2kGv3pTC1DGDO9my80eUSiS
x/2r1MYhAxE/J5EvhnWR4DiCHYKimz5NuiaDJ4LM3dXFHDPrLfsAft0bTe/+EeB3bvBkFfhwHlmE
jfJVp5aZS8J0fHcJWuqi4xorXPMr4VjUkjPxu7h51c/Yvte5ZztwxxTHIrBuGL39PH0/NPMR0Z4N
hBCqY+X1v9Eb4S1jqzLGzzL1h86wk9zzPNMSdqwMFAvCopoOy4xGf1GRaKm0Q8tTbqhwx/kzc4e2
3ApeTUKGLuGSz57s54y4Vnc93x9lnm6fJOhcZnlkgn7SYbJNoURy84MbUmE0eOJ8GTyYtXK4MBGY
RbliYcK30Kn/xp75/ZauK/SNpMtkkp6pGm7Z340e0VOEsn26iuZETjzwsrbaW0BOnJCYVncbioTL
nM0NgJ+eqmg9KLK5zoyH+/SYB/+XDq/jKB6277QEesqRypxbQRzUIGYDZe56QVUgU39Z8YFywdub
OCr1mm46P7uTZpJeut8OAZC7+1DrLzDEVvJbrBtKF8sKit9Trf6RWKI2kouZFkj3aU9B5rSb2gfj
tWN6rB8du23lwE5PkenETnnLwGjeMXw6eZW35TWBDLGQ379t7+rhn87pnzZ/ZgQbBUCsEJbIhnz4
2AH2OYvDi+ZIeLXnLJcazMg/4yxvl5Hyx++Wd28Ux4Db9PL2mLkR7NoAyFZtHb21RKw018YqqPnv
iZqqitZosnJP11N5W2JhgEv5IqHMZR3lqY2JeuC5MFnrw/JdJViGreSEVlz7qNHotN/FMG+WtZJQ
vof2g6x5pLj2X4T2gLjv+tkeH72QJlxNcfoMPd7VxB3359vm3e+jhLfIASyw3MY9z3OeG2AquHiE
liO3DM1iSgIRgT/rz222+miLtt+uC0F3460Yh2vutVtw7MvwXowlFVZhFoFfpmMXfmIlrwNaaWgt
Z+wJ3JKzg7iOCS6ui3bFN8BCm31W+8At5ZnSoPg294IALHvXC/bNB9ry8vD9xhAtVOZ9pkq5L4+X
Obyks9qmCXIn7T9SrpP9NJPSED3aYEKDJWjOSEAM0f5wl2IDCmcj0oNh8F673+rTvWqxHvxTrbID
+DSeNk8hmlP4wytwFna0iIEgAC6XmaQebs8mPU+G6SABV8MwFj4XsQ3U/ZPN307LdIjBqpL04US7
PfEb+yDYeTq1P0iHu2agheESDPBD5Lq883rxeDetpvHUeoXLLZ16TLxn664PA8oxOmxvjmEppc+o
93WeKyJYt+e2GJ5YMk+sdKKhm7PTEzvnAlwZDxhXKTzrv6YN5ma2bJoY6+td5DqU32rNKHY7sW2d
XCtiDiJkqZZB51hfVOqaRvpWnadnfY77zxTDhjbzWvfkpMwl+R+OZ1WH+6Rkc7YY/Vtnz51TjYJA
7wvuqiUuxw2sTv7S+QxPQ1RMLF86Nws5gOpM7gDN5eC5jGvuN9Z9UnbL12sK0hV+BANaG0l5CVd8
uIRG5inVQae4PKraVxplsIcK6U3iC8tNsWy4qV3HawN05ys9sPmBMDUEeyZR4uUOBG2dAT9+584F
8Bx/3TuMIoairZoJbAjFWEX3mV61KDvAH86k+sre3dNb2gXmcmaV9LtuAeb+GG+sQTg2unmqdFUY
LeoViWlxIrqOiWh0vQbEHxTOYHBD2MnDUZJS0TbqMuZspUYqqpEDS3LVG+MgejeswiaFSOIcGGHD
vqkdclH7+gk52IxrgdgD5CVp6gq9T6+9haIDuZksH+SdEsl3+EOCf1cqyo5sk1pvqFlLX4Gk4ybw
JG4bYFrwTq8JZM+v0aw0COBBAejnIPT/MPi07OXhRzwUgSTD4nFuxFXHT9Nsrz3T7b+C2IdVdLTS
zSVdFYZb1I73B2S44x8rt//yMQvZn6lSExgV7EUFLo680yaRzUkvao1DuYYgFk/2i3HOjQVeJWA4
R44JsSnpyEOhtXk4ii3OP1DYAt95kDfJR1x/eZIWlYvoRbkZBF0zvU26/TUjuTke4Gz1yNmoe3Zj
VVQGSDBi202W4qFlBewe4ZRCqT30r6FnpA3aVunAs5TdE7ht5IZMBiyNlw8RG9YTJxKZi/oEBx+2
etMvImmkEc8CmxCYgTXsmG48e++ZgBu6QgZ41ETCUnUBcbzZS+2dGXroaBEtuysJqb9v4I4kcrhc
0wulEMQAlbogANvokkDbDIBAiDxAutLpAxGGRBmPHDyhSgxUg+WXTjzH+24xI8Sh/bqqztKgY5QL
9pJ56O+RXjx5/9rIoh01AmUCVnidIW0FdRLLnR2M8rZnEPAlJG651AFNvMZvWU+PmCNInrEJe0Lc
mpGmA+KetTb1wF3yR/VuH+HYmdcNriIj5ktvWfQ3p4rNI0lRfH/HgEmLPGFw3hPfS80k5LtY+v2h
WT1yhSQbLx8SJqYvEj4vGjN4dmttSAh1TVPGQiqwLaTMPg+xDSkm/69tTVzX23r3S1ydz/hH5/Xd
yI9Q+qHfHTMkXs4q0vDErG165bh7Doo88XmKJz8Qocxm79BosLfb5j0MTjTBBlMyLZ67JoCIUybi
L8Zugf42WBSPKxJxA9v/I2T1DnPKON7KSoBuBjwE3yZeO0fC9rZv7QXiWe++RuiUMviI7LFhJt3b
fgegzP5WLQN9U59vzaE9tGCl8YCNmajA6oeyqt0F53KaY9osWW5MbCu0iKcHmdpeBtHSlQxQg4hl
WngOBDLD/OgPINObRDCXHXd+LagumIDxTG+IlSPYUtRTaIyaHM8x/Vq9RbZcUNrj9awA/SZ4CIQJ
rNtfhJMtldxL+mLU7djbuiJWrJSBBwNGa1fRUfXojnnm4COUOBv7ENFH47DQP0rY1k2SqzfQ0toj
yNcC1Qor45rnS2YNFwsIoePGIVTlVM6HPUZSUMB2k/1NT+Q2qOCoXs/vPJCUTxClzpkd60vnR3pf
jMDXj/nVug2LxYhursrLj2NdDj0+zQ+BpQXQAPhYQY1UH5zM1YE4Y6NN4O+jbSynotgI2dZ93w19
5rMIz/vdcfGmAKoEHWrE5rMtDBofzx/XsMWf/ba3M/c9tAGBUapAuBBw90OVRp6/7LF2waNtsQHU
odZd2BxdY8/K+LzxGguoQFJe50kzrIb8xRL3Wz0RugboOcChhu7FSbByeQqF8LO9otlPax8s5cBN
s3NmqWXx7VxDBNJFBCToSvgdE1RBuszJSHi1b2Uk7IE4yCbQUYcAjJu4uT6mveaS5Yt38PzFL1rC
FuDkgvNUNVJhD+rSore08rmDjCxKP7rhM5axXqftNWKUKdJdpp9PmxBnSNEEDjN3QmldZCW5vpgv
zAGGBydegZwtDYJHRt4Heex8WY+z9h86dPg/l4n+TCYVQhzlRI/KVBenxOHxdTwRR5qcLPlaXxHo
WvG1aAz9/PQViGe3kGJCeqd8syH0BRaDS31Mee/TUJjee6M3n3v2AhT/Y9p4OBcMjd8/mZomAyLu
bOTiC4dC5irMNPkOuW95bvbouWf6Nce/mLNp6vJoAQqP294naPKRoy37EqN23J2us8UnlmL8w9lX
jXz8kbhr55mRWh7/fCjjmvCykMCFzgS5/Ahk4Y3UEMtQCtLHfL4cDXAQIScA9/bNGsogk1AhiZRi
Vq9aH9XwSNGmWORgnByGFd8OR5xV5lkWodDh9z6FZmjIbPpF3lserOoMOPVPTWv0wjj0x0BX9J/O
/YOWvUbJkhlZg18wsdOqdtN2sCTCAA0Zk9Z8Sy0QNUIMrebR/DA3DCe72ebyM9PzSpNkTxkKkix+
8Z8X2K1XwKaDWcb4KqKBSORIGeI1B1arOyI3i4InCU+nBQivxBUu8y6wGgrw6ZZlSQO5uomm86k8
MFIHqexZOOC36pZ1PdCbEet7adhNXCdwQncfECCFFXkRvpv17eRWavEBbmf0YJ65oXXMQrTd63OB
1y+hwSdvb42eZehGZnNcSEb5E9wCI8b0ElH8rqI1eDs9qzeBvaJxwrpmPU1GKefonn3ePw54RFMA
Ud5cuOgKn/wrNyO3E9URllzOiIx7DXxv9TIjKqUjpGu7LdR7XqzHDV3UjcDppeHA4xRWionB+CkC
TKj5XnrwnJLjmhwqRgXGDANkBpWH+OqoKF7gMI3IWtfDFFE1kkfJ30m4I4/+tgRdeW6HQiaqRj/C
ThXlD8A9WgUqcx25ilODA4IOajctbnAki2n7do8PRlcOOqeb6ubpKOQ6wFjNRg2fX6ynQlBVGAxH
Gdwkt5hHt984+aKzO+dLkWC5gFkEdsj30Id8IxKlfkocO9W0f14tQSodoSdAZPriNoODrjnByE5u
yFBN4irvmCANmPuY9v/ZhZjaP48NUFdJ+00+gXj54mdEIF62hHZWl7uCutkMEWri2yEfQi350TFH
4Gs12S4du+6UaGE4t2YpMPxu4+E1q3kY7T5sYRS9Qa4tkr5U2ICKHw1vhyzycMok2u2zDOIfA9Ir
b3yFrEDCfmNrBX8tSyW0u5f16bILZt9NOWhaoNYiyZGMqPDp1A4Rb/lBlKV4AV0q20OYk4Xas5Qy
b32iHzly6/ch5LIukzs387ZR8YYYc4sWj/860/ANgOJrMlArvI83Vz+/DhP1kX0tZbyr9l4ZsRvf
Ot74GOmN8KbgBaewZ9ttjL9keoSo6X539iti8miBMitiYo45EXPC2rggUe3SiC9w9qEgDTTghpeZ
xWuwdFMkVlcq+gFDCsRTJAMWN1opaBiLC1OhsdJYN/KAFM6u3MEpvCyTaG1fwOZH+38k8TXabQsP
ZcGY4AcH4WJOKTDXnUnUhsFVR9/47TP3iSwtE9x7vECNmxnfO2Se/ZlpZWaP0lGVs188dROnRIHq
lgO9iELXNn4u3oIruuWALTJ+rVSZReM1LeNqKTLkoVLV3KnTYn/Act0nIHaBm7QSGQayo6bBHt/m
LjQ0qNy7JF1EqI/kMv1JlLuJ0FfZLnIgJtUYpSKoiSwmmWWqPSgwtOr14h4sN7s36GtxhDxF/aCL
IHAhElEH0E6hg/LvSuYVrhUfA6dlnKpi1wYaMFvrANPVyWcYKH2CzwHh6I3au+Brw4prqGWYlQXg
rRf9sdk3d9ybZYxShnZjXkybgeKnfSbikToEiHt2ZgAX2kdWQP06rVxLCOegRX0mA1skPsq5pDUy
s7w47L1xnWimtHmJM+kkOjGJJMeJKWDLan5QwSb2RFAreHlxoFV4PqYwLIzFb8lj4DzszpjMYS8v
Nc8H/sFZxldeHsHOZhTQY1/pukYemQt3wg3pLJaUJV6r/5LO4Re6RB4jB2wCg+NKCsVjC1h+lbwT
uOC9aAYh0BhLO9Za8Zf2Z+NQ1HDWceMGFPTthoEfW78z36q7Da0cmUO9ZfRZLeRAlNqwkdTBxTFt
y98HuPEKv5+JWNsFXBCtYGYKg/3ZYhjOq3UgQ+AFIFGezgTTFUvqGYoLCmgZ0HMo2lrbggBiXl6A
xjN9ecgtl2DVgcWBcKtlxAl8UfCUFXegcGqtIh9dgMJVmZwsAICxWgdMzML6W97LIGoPVdx8o8mK
+4FCfVri34226Ed1x6OztIviQ2xrfQNNs89YpEQ/oTh6Sgx9BmL16mY7ybGdId/LiR6fRhA0UQDi
JE5jSd66sdDCYBd8ZbZuBv3el31E0Ad5GDfWJC22/J78+fOFobOUVxpspNDXl6fg9PFjnRi/B0Tv
pG67st+rolXANwjXa4r7GXcH1hVbD07cMo1HsLQihlPPZldstOUlzOFbjAFau12FRpK0QdGbXP6K
KNovYksCp4RT+aQFeN//z4bakE+xGhYtVGWwF59u5Y8lthrgl8cLfaI5yI1SvjAS0cxnWAwu7kQ+
nuwPH+AkyQNKiMwR0Fb6h4dhRMlEzbeDaEx7MKE3TjmQKXhGNboZS2RrcBpzxO3ilOGdlm5chiR+
eHOMqJTSpJxeAm9z0sByuhcNvAVBnVLyRx4B42FdNs+ZrHIsck9ceeoh2AN78etl8a2AZ8K6arkY
RRgDR9VLGL+HN6s0fMfYLTfIjv1MVCH1HSuzUh/Qi6hpUT6iPGzvbTUjLV2JbIgbqB8oWACCgXnC
R84cGdCWIL/ndtAqG/bvBDUgrdw2wivI/aahfQUaYW3URkvx4SxN2U6XwGaEj7yaheBvDZW6mFNR
siOJWPuDzikZqljp/Pv8vYMaedGKh4nJS+KN778sDDmxr71y6sL7CcCSa0IesOh1jccOyoTIYJrL
Xp/LY6QKsomU6bF7Q8g5K7rKsmEirQOfTMMJc0UE7392GH/d3JShGQ204AjETt+639inr9z+imD9
gepYzymkZiO5JaakZ0KQaGXnfZ2NRoU4BykdNMvYg6IE7xWUloLkLOxaehUAtAxPN7e+7+nsEqd3
tml3+jqHnyNZ1kJ2pH0ciwf4TuTg7YubMMQJXhMQwMTZQSbqSTGp8BONWats5MrI6WhaHzla2Ngg
Npw0zF41F9z4U6vft8u9Ezzm4C6h12Mi55Zqd5IjhowEIb6v6aA0JB7mcZpWF4gKrdzKtOOG1phW
Lezei12m4JD1fSPjKYJqTjYpkc9Oak0paZFA433TGTfWqjaeGL43FEoZOWvkbNpUZaripeJjNr3X
RbvBdN7vMgT4BeVeXePV0jV2CL5JMjZwx/wrLVnC9+n6/gRu/C2+GeXeUBVyX+nOrliuJc1OkaGO
RGPkCwYBVNy6P+8NfyyerzQe9bHNJw4e/YLAsZTtfXKRIWYeoTFSs6KzfcAM4QZRGHRMQl4DHul1
sozp/oZGSw8IM7/hCZkhJGhOjHcM8hgIplgJfpF3tX5d/S+BdXiMz0exH60bFET4GCLcnYY+dYc+
TwchskJSEaqg4lwtc7TH9czWUrfwB9FbGaHpyjPi3pxIcU82PACCdhdfaaLoqbVyRGGIwLEoWlMX
W8A96n681062XVjfjm4OL2iyeScL7365EzvuzFSdkSqQ3Rd02RInGbJs+kWmMSkIuz9lCo47nG5H
Q1K0gAfSYSuB6/HlwvPSii43r1/NbbjrLVjww2WwAKVm+Wi8V0szj4T/55+XmmthhNu8+c/GfAjO
FgHaKgOvQ92YphwbwR6kN9vjESKlR0j+PlIPhFWtfUFOjPqpK0lWoacICkBxrNsCue42oBYvuHTR
UbubsqlvxRkd37eb+2kNM2jBb8SlBCS9mGX5Gxya2VoAis442eNnUsPUmsys3s53EZhyAWsEOHil
3/KNPXNvcOujxi15LNZ3y49yXVhQKRGydyT64HKF8eomybbj7KbqN6HT+2k+BSPzv90KZ3KBUxLD
P5BHrjEIqC8FLyZQmfcJw1g23Uxx2H1lQ28A95K7QwOpV1cfBufpwwButC9rH4RkxoPsUhwmBAPN
Al3G1tArg+/QWu6DaMvk0dx0HlR8oJN4mGfud4DTKciK/JHJGxAtli0+OPpGEb6iZSSqC6G5AIqQ
nAmqWW0klNm2WxOojOdYuX7W5oVkgfYL+1iXrAQ109iZWe3rLk7x5hwZVDYSkB48SHO6hZweOLte
dFB4mjeI6qgqBorvKgE55V5EZwva0HRiTPkwlsBYt4wxYZpy10bDe7mQOcJH+Wlgy4xp+uQVn66j
UnQdR3rObx/en+UYvgNJ0uM2mIqkf/154+5PZclxdZQYIlco4il9j4O524RMjZ5ovGkhqOHAuich
qz0Hj7EFrobf29AVw1sSwKcn3wtts+jTsrtqocztVulY9GpsJueEuSo35d2rjNCr7roogQTdKuzw
VsMdTKp1iTS5o/jzJO11+mbWuVEKFbXlUbESyUqHaOex1PaKZd+Ir66UKmw85ALeDQhik+K2tMcT
T1BHlv5gdjY2X39/8gyAg/7gi1fvY+hptIGXsXzbTonHDysnOlkfhIaP27sLzFk3+6lko4NI9R2i
Q4MVujCl9IGd3/60D30C951AkEp5K7EkHsOxEOycFSNXmdVvUKxH12NHDHGrPeIviT9IgQOuwDPQ
WfR2HW1bhWjj8xEhaXkJTyZ2Hj+aEo8x/TXHYu8OB+Ze0/bePYjJnVyQEpreKwHiZnd20674xaFX
GXOeiUn7HxOyejP4BLtxucrBd/jRijWtcS5EtVdg5ET5aIXqFflIouAIJMowGq+lD+POuGzm4830
6XtWxf7jW9QDbc4TvKiJqnQEjthZuDdVfBnI3ghIJv4R9D0U6owkxBKKm2PY7for8jcBPnLeazlD
wY9/R4AVenRG/UHxiaeGAcTGJmklpHgimxZqTbrydkn66nT6e7BvPFH8y69j7D8ZWLFHTJAEObQo
ZvEB+/Xd/CI3yDFxVajPC195eQZvfTUaIpR2QMULmj/V/IjNpul+ecxowIJYi4yF0tyzJ/6c6vnF
4b8wgezL7cI4rGBL6Rfv7z+jmNL2eoTxh9j2Z/VorzyYJsCpR6ROTMdci7Qvqt3G9CK1f2bwWeq0
0PwEIgjBiNZ9UHQYWgjh7H+EoQQRSH1Aie7xqj1gvwhmlAPa157VvYoYbdDerUINhM0ZaL68S4oB
aLsmjwFJOfcdk8O31PLr9CVIsVLghuuZQJEYP0hVttAdZwkUnZXDApxem2FblCt7zOUVjXlwu/kH
ULfk9fVLWr92O3jsnW40EY0qTOBBaG02vB8u9nt7g1/b0cTBVIqMF8i1qXAL/ThN0uuLxWtlXLiM
TWrdWNMx34z4TkawtHMwRNtT3h6B5I5AiKNj1MfELpkBtD3ZuRAUdghvsMeEnUAWrFh9IwzFsZv1
7cp/CQMgxSrDxb7+Rln/KSJyT/pVMMs3BBnvZt1tYRzbtfaTlcfuxDvaH8L6Shbxd4Y5jpx8WP2L
9Iy3kY1sMP8x7EYE7JArgVcVOiX5NdzeSM2BVd2JCiAwJuCQfQr6SfbN58RfVG22wuVnlKlsYPYd
r3sbd17fUVr7mZNqQ32bkmmDiZSsTBMOw8HQ3hIl1JrbduZp0vMmWu4T/8/EonrrZk6cMmE2q6po
XiHc6FJDBGCbse9DyLOE4i5kJSomlusaufoEkTMRU2C3u9vMo4S3WpA3Yr2zspFdKXhdnUvUZhai
nJE0lA+8YUtigmxYWx8fQTiGl0ns3ES1olPIxZI8XHvrkLBMS6ysM+5PqMVhgmOzQFDZNrnoh+Kc
3eU8b1krnZmYXK+O/Wvx3mfMiTk3usBxzH09Oz9GiCzvTPrOm+fdIXUaPdbxyUZH9cWrahBQCdNr
oxRjQapkmFpaSz5p/5pXM1RvUvSUqzADT7gD8m5jBif+ML2doYJ5NPVNpH9RmjwmaEzKsLTWys5w
I9mfs+jyawjn3Q1nSguZfKRFHfH3eIz7txmQ/oyHW9qEYmAL+B7Ur+nyO4fwT0PJpccj+VdLVLZz
57aGAxkx76yvZoZQSgejNw9w4muwRIXjTMKQvVMvrASwGRsw51OC8mjsvz3XSpuyQaE/2DRajxr3
/njwcdSwMQbITZXZdZc8PeAfMzzg7hcj+ii4x8ymJzNrjjWcQlWWH+1LTOMrJGKkatEfT60Nl/fN
iIoXQ8agG8NG1e5tRtC5jerh3IzojwEBH7d3WO03n6pH63bTttaUARdTDoezUtBXPCNnbzNodsOy
uvAijORRPzKKXK8nIBz0FCy8kfsyddVoBFUhQ0A29gSAWgxXZaN28bBV6VnFG2HvWYDk0TCbEIDc
7wZ68dE67CdybU0fweblQ8oDSmHFUbFkb6U26VgOSzqa7ij9en3KS6n2xD6G0z8705tTkVYGNe1w
xgwtSv41nL80vBAOn5T57LE8y9cQt9op0WsuS0ZtdLMccRVTazqn/hSc37qJSTf1O68EWbDKQ2Eu
oWbHSgSrmRu+7JZPJfM03gCzfIbGqOVO9/pay9BeGAEVxgYWWe6Ghn0CyaHvYPHEOd6DuBKRsIa7
Vhr8yx0rVp1fGtnAf6eUuPKBhJY5Ss+P3JNVFQ1qKJr2w9V/uV1J4X3ut0j9vN1WM2mi3uOzsACc
yM8lkahLSbHlZ4S9qlyxEEcAhEV2We9swsZVpGi5YHWq0on3MC6SC03xgAg8mXaj5uvA7+TovfSt
JK2Rs4EQ6fPr3YCcncDH6GBOXZudFqzpkBMsCKXhzFVy8E+3wLReDxSwwvGfn0TvKdbV6qUhl8XF
4ffaqzT+RfuHmQN6CpwP5wCMAKhkmjyEvIDHadEA/vw/DjDPvYisxR/v1t/ifM+AicLrNd6CHpY3
NZnR+ZVGo8NPQd6A2FNamEi76/DwHxNEMMlHyHCFSvKu/8B4qsCDKOE8rZUL/hNND1vKqE2blA30
oKKP6p52/lJO30uUM9W7jLq0lewk9abfPEtYAAfj/V8LPNgvmJGq/K6EzqaJSkTwKDImwiJy6tI6
tNvPHrZicHmEcMbeHgET+W/P6nQtYOVgIZBHeResof7l0IwIM9ZPYTqlQqat4kWgjGhwVyDkZS3K
VLh6H6t1uu/Zi1Ed3gHvsWUcNjPkDav3I+bEa49mJPQoIy7It0MpC+LMovsjnT5VNn8lO+TlMR6I
Sc0aWANxwsuRqCIahOFCOOR1kUXp1zmsz4hCqVFEDC47nZVfYKCEFVT5oZ6vdoBnIrw86aQSYrZe
XcqpKtBo5f4uzBWi/BUDZfrDCHba58dguZ+W6NRr44tLxQONLNL5QUBGlDAAeH5Duikx72cwxM97
UWVB8l/fECNsvkCwzuvZ48oZ38zSs3yKlFgFyNazLuyvuE5k5wCJ2qO5qQpi06typ3uh/7816Bfa
5MWKMKBS3MzfyucxV3E6CV/e4z8GthBY6t8ClzrFPPKT5NlT7gEPTXC4jkrjS8m5FlFEtlHCSeUO
4RG9Muf+HJyRU5fF0ZTVowFKmkwLyqNmNYNWUyfLF3XTt7UeH7GJkcLV4zqQJzU7phqGfxykYTp1
whvMY6TfL3kd+0qwEEynEiiqnZ1tL8WzH9Qxj02lrLEIWk+P5B6Uk7dEYafyd2ymIgVzF3iIt+aB
sy85aDD2lIKupmzOvY4UgiUkNQTViB/9ERxoep6HddeWp1hUnLMc83dXwjCiZN9eUybSum3ab4en
5DSwsIfgyFPflMwLiKPBOObAD0SVAq95YAcwe88wq1p5AwgMyCPLQh1bTCCKCqFOXDpLWJgyUF0n
eZ3Oy0m03NXc3Y8TCw6eTyHBrjBmFylz/RRaQqq19qbuyMfrMMVnUmSg1yIngdCsNOOXMdPzSgBR
yCQMSFRoNwLMHWHv1J8xeoyob0CGfcCiM2qBOICoQYeYcsb8y5q7BHgvC+SXV+ixzIf2d2gP/Nhu
I6lQu2jsHFR5WyxeBQLB2NX0/KrK8IyiZ9COCQLgoKtVTO6bYEHyegFeDZr3kw/lpmt+uXzLps/I
IQHz6XY93OZbk0aJrkIl7ouAlpatW3YsFWQ6mPOoTi30X6HlL3nkCf+Dh844ugOIBHFGeDXby4eZ
6G49sWaPHGLOTN18xGxVObwYX0QjQufmqDZibwkaB5ClruPaB2Qk4Pw3hdXiNKGQmg3PGmuxcPPm
I+KU75E9I4fKXulrGzdHYvdHbbuT9ztHfVJTDNb0N9kUENZ7dwafmgZaM0RKHPvAs03gUEYdPT1v
P5wyzLHBvS0NaxgoYgIMzzLZ7zwoFlit7+Uw93qV2sHEp8MaTdG0I4DkDY59ZBI/fAKpByBMkLK2
CMX3/sKkIItsN5PSsiRd8dev2gAAKCb718Muqh0ZUAhafjre9vwnZmBQIi/wdNZoRJMVxEEvcRyV
3JiKOTBaoXyTzVO7l3y56AcWg76n3z8awSm2b4Q70Zp2ov6hbpmP/NP+/2G/4Y8ME+chwBxrAQTc
mKGZoSfBoa+rPURzpqCxfWyL6mzFkeir8oRpUVe3glP9weOr4lR2eLgGkjKVrtN3KVpilI+YrmBC
jKjIShX1pagiRY+KFfLykWJOAEPfOdKoymEaXUKzGgNQ4ymlKqqHd7SjXXmopuZWL5PjY7WzUh2G
TEexf1uYzqwG7+CvoR5Ke296xfLmyyntnu3n60oCE/IVYx6PsMR/vF79T2Lr9Q/rCvJkIgtP87if
CbhQYPJ+cShFw6Jrs80aGZAiePkD7z5vtMZJfufKpwu5++xQrCCjjRjtCZDeHMkNPxrAsNFixTbL
O2BR+AYmy8SFReJCW93sRQ8EleYRTYkAzh83hSabYc6kI137a+lv8m/605xUlx4ZPSFbz93TLSG4
7dIXyNujYrF8la+rgTRV9s9Hu9Auugc+EGOy79NWjovUoz++T2adxybWJKytD7AfWm3eNd13j+2K
Iv8G8Y3lJL0gFssPJpcGkSBYJ0DXzADf1dg/Uv/qh3QjBYMQNnlUeKPsPA3M3gZIGYSizTb8V53f
Z8JuHQq/5leGkNnPN8b7Cb3gl0tiX04rsSMMkEr17XSao/4uXeX5d/K9rtyhQvbE8c0NRTGVUwtU
Bc3fDiyqDdenj5mziYQH3Chz7wRkm9TG1JZG758JH0Qx5H5qKCLJwfiLKetXOS0/8MhokqjqEEVa
A8O4GoT7JbmhWqCGWA9E9SHX/UDOgrSdMRumYkZL38FLYyRtcydUaDtOjkBeJ5ei6CHLsabyx13a
/hj9MxT6JzpUtseVLJS3V+Hj6m1lcaEq+ahQ1RqL6VxDWYBzbYAYbaptRKHJDd9SsN+eoqOwwfdl
bgUk5KPsLesj6qP3XZDNNbsy37bHyYSaN+BJQi+mV58UyyWdU/O7bkWGCZzb/JzRuTT0r3xzd8Rm
pUpB/a2t6nMB5w8RKwPQHgB2v/B/sZgiZ3pRfBfRryzBQFQfkGqNQR5pIu99ce/uPF4OCQ7LLGmo
yZKba0kNDaND+DlBDl5xuE7VeOIpLboEZHm4sLill3XGAQTYWXzZOOmY2b0cN70r/vinkqFpZBQX
eG5d8O7oy6/lF1cPneP2/NQTedrSVh8caD+3RmKN7BJMFivClFA9orFB2jdSXlvfljuWjtVW1AyU
0g67quKo2ngIvSCgz76ZVsRlp6MoEU0tZ/Wt8fULzQea4yR8EXeZDuY4gVLO5wzDjlNYrs4hfiiN
XsHwisWPVKhgCqzSk2tgvadSnBMEogKRr0Aqb1kGVhYN/VWq+LfGV0G/Wf6yMr20eDLLo+8vYxZ7
ReAP4PD1NBgpQBr1Ngvny0FxmXuW2/fjGUyo5uLor6g91vpoijgB6u0BoJ9QfkV/dob+zmIZTr/u
DmdSTyWgtM3CMJl9EwR63wmyQv/T47+Kmdm8NrhQR+FBiX8n0A2iVDgEnG6v6iIdxSgrv3yJCVov
eb5rydV5RmjneillC/HvHUCEJZUjY6j893j7rj+Af7BtupYBlp3Yl38USbwSdF2wnBeHYpjn45Xd
lDY8+2pcKH/bXnGVEq/r/R7cfhLQgmsxskEzwxIeQlcI1QvnbtQsZ0IFTtCVhW2val/WgivyWBSx
97i1fo26/2tltSLvXoOtttd8A3fhTP4YtjmhNz4Tnj/M6KPGgN7rWzoZCbHGhuWnoRUZWm4BdlzH
V65Ouvl9qg7L89GNALNaqm5N7i27vpxbm8BGZbNo6gndVtxE0NV8u3470XTk1J6rH3c5kCBT4XO7
LsIro8lnX5HjhOPuQXl2lec9gvR10j8ZYxje54yXpcyq4uoslx5ANd4ZoCNxtAwd1qBVTDKddSFz
Mh9sqiGPgrevDRUHpp17T0n88zJ+aF/W5iZxtgpVg4q4vSXuhCyZVHWsOzAVJYp94buK4oDthWzJ
9cmqELCQlXe4mhFQ3yYG5hzQ78ACUGJZ1U+TENe98vSF7eIQIjePllKxctPjsqtAH9KRSzqSdy/1
drsjgLmF+LcxGUrY5gmFq7L05NvJzXS5gV8VNqWvYaDhKSY+n1w9E45ibzDOoWT61KRzoO5JahnI
cyvW1TVdirQmFoR/+IDCikPHHaMQXnIfeWH7zMcPj82dSrWc/6losbzoMAt68IXTte5jxFENNNg0
zuJVacdSsP/Oer4XiHnbJfzioJ1vKJ9IqYt0d6vrkPpeVSMy4woAvdRKjrFYThdNj2es/2OZLhOH
dSKDoFKXTxTD9VXZ0rmBjsy73iKuWvTmrFpgMkGkFUfIpPaysNYjgRHsEb7MO3ExOwi0O31ugNwL
klsE6bE6ShzLJ8k11068uy1f1YGJ3O/U3E/5uJd1rK9232/0F5V4A13+WsNIEKwyBTF0t4Oat69k
2rTE3qOp2d6wlPM/o7kL+Zd+EQZA9Dr0uVI+rKBwJ6bRDSbaInzrNaIfd283JhMA7Ac4OdaD3Ghf
CGJEPzfekePoTiLSJYnU6l9pMWVr8Yj1TRMNEXCwXg/TrQFMiE2uuK1WClQOy8IOOqyEkOGPcCc1
OgsvIIcwwHuWvJX/jtUffiaek+/Zq4Q7oqR16Bcz9A5rjZSaECu4tGsT0Jzrb6wrZP4ZAzQIhIvF
2KZlbdS7oBCD5rRjXenOY8cNwxsAiUpIgB+va2UzMIVgBE750TByYZMB0I9pxTtLUvmnFQ5SHlCZ
Vy26ofsbUQucthH+tooi0sUSavU9TUE9kdEVICfut3afNZBwaTBZID1jFklA/6boNKLrF8mkyrSb
Ay+O0MnL/bXM4e5xrddFnh8feZTOavzRVLvLX2WXMiMv0do7YnGQwd26YgzscBCI56ZKhrzQfORl
M4y+IdNkzxom8s+j8M9m/e4tMksCyMeNVjor5+AjvXGxlstJm2YmVLRkr71XtzBn+91CW0QGUfdV
i7rgs2goT0MuKlU8Z+aj4PEhtiJtzsLkdOl8zZ0Ej3CXpigG8MBWYj+vmkkg/RTXjA48fdn4EhCa
NllTyhEBAz9N6qWTpeXYLQ3C5n+70aDZye2le2DT6eqOw+xpYfl3pe1W4y8D5KXnmVsffXg285/w
qhh/QdsbUunXF2DmMaBgXXPSvAno2g7QOKwn2T+FtLHy1+XpnbeYufBN1LZBgfijjAgJZXVRUXQs
sBxDGOJTYfJW2uIvAsHF48tVZZiP9wMeFQNt3ClylMPEb2kNQupukzIIRnCQy3mXsIUo0Clsqp3T
u4ZJYFYTyctCfF4Pw7KJgt+R3g800wQCKNPEVkq96msKLrIW8GYZIlN24XsDGlE8E59vAJOFVPNv
inlj2oxpX6a6jR2CqpVYbyInKssl2r0+YQY8yB/44VNEc0/XVAewXsBWqmVaBWEBb/OKN+jCf9ul
amuSR2fyfbguXixBiZgbHk+3JFwchSF/oMjhAQbxIB7vMmncMbdgDwg19ct70teby055jeFQcEEm
SLVC943U2mZcYHnSnZY2pIjlNEzhP0A8XuHYAobsIh5Ie8obqDelNR4Y/PplauwhxhXMKHglaEiG
rGbu3GEWdTcOpKjtDXEffc4rTe1ItXgM52Ur1U9xHUXI6lOx2l+1gwmX1uoKjZotu/qRI8fawXZ5
nEKS6QhF+vIsv1caK0zz1DzrtS+ToqdTNnBMgfd3Ls/MnKc/EBxp2IDvyEu2DmMfRd2MoPZkvkVv
0rupYmM2SfLniibdPN415DowNmOzQubLIEOJrd4n9kudtJQ8OtFVB4A2BDSozhWpPN2Ha8J4CeW5
ZPCsGQTMlyvOInTkkQqQJHTFkBu/6e/Xa9XsmyM8nrOMUrBuq3DROX2ihoDLFCWDqM+YcRRzHQPD
s/VTIYL9koLuL0SJ/FHqBoCH9uXXuflL6vsPLAAkar0buQgvDcq3t/h+ognzVO6SvILthjRizJXG
bHCmh54XyipLaeXLg0SG11j6PmSfwYvWs4c9maRL9nmWkbCzTtlqqGw+V2b/GJoHpJ5lzuychBAH
olLW9IB5O+qclMA/89BAmZz7iYv3UvFVcFkrp4EHSe5+5sL9sLvwbYuNovu4ON3Ay2JI6tSaT9t7
bw4EiqKozjsdDpv2qG3K/rx4O2MLyHpv3ebxFFRA1Ff3ig/1fCwx3INS/lJx7VHW/z0OzjKU3AGb
fStubi36jvJdCNIlEWSdMwbgokr+KGT7RhZAoHGvPNJzob6cGhscHV1BL6lpgn3Zjr04runYuopU
8oVajfNHqRNai5Wpiz4KLupAjXIL8LIQyQZIibSEN4lLRx58NbtPPxBnSVaJTT0zteGHJ7EM1kFq
9gN+8mIJqvX//wTFcvkjU0rxkAfcwXSrIokheLwsoFQMuLBicmfMJNrzE/bZ68e+F2pd+nI1zT6m
wGVfG9gCBecahibpcbfcmupAJrLKKuliQM4IIvQmzMTFL4RY/enN2YLhhJ6Gf5FK1Yb4lh4cuEvW
QcsUWHz+elcB1+zczsASWz8ntGNIVqy4CDzexKtehPYO1hTpAl6rAtRyrzVzeDTD/VUeFRgUdzRV
Lm7VZ9tWh5ISnfAdjHuDcZYTACdx3lWiXmTiAz5F5//Q+ZFFHJ8v4o2bH7lApHtp1+ZIk16GaZkz
kWKaY3oBxb3unns6Fh9NOrS3UkbTSHu0oBp35VnZrlcIj5Ryaf+Jgoq+Lp8wOphVOwISB8lyHW9K
qFrn3MnDs8AH6BOhT6voUgytel3tYQuuaNfMv5gMo5XEzHqB0fbFHvsmIzJ2FCW4C/aGsY5WuqUY
2FIr9wa03oLWPHjwtpE553jq7tPBrWES6LFUGF7nnkspxBUYPsSUS13M37I0iKZgM+2BhD8HYvCK
N0lrsqD98xhp3e3SSlxmc1NjB7D1HbXrSlMqEmgyJiGW/AIdSnNRQhziRBKDIb44Y3+eXkxrwgeY
MqduhBBjPLNpMvAywhZ9FDL+sN9G7l0MQJzldSqLmgZje+e8XiBFDklM+TXOGaDLEDm6omd31RDx
IwwoW8+wxtnPk5A08cjusqRfpZERXmvNsyEuhCPbUvWiFQEurGTZKq8Z1oJdqeieJJBcxV/anXHG
jWFhFHbDq0/m3cLjn69MzXztuzUlPpujcTVQ+ifhEuEGR8jMD6FeN8Xvyc43TyVzL/hGVknE4U8p
UAOneMoKzGEZhD3rE8lwkkvC+6nBgrCET6ewTl5tLzsslC8ylmC3I+zK3t9L04JJudUNYNA3ChG/
WhiInA1jHZ0UWGQahpstzyNQLfLT1QKZYxlqf0RlpeEJTNH3/79Vwlo6DICb9gfXvsyRtZkQAzR2
h2s5HGQGnBhUkqJDQ+jNWlaiCgWkMudWQjAMDn5oRBnHph/vVU2U20OAvRYoLhK/0YxyFugXj0kC
GrJ2yr5BXfTcqJ/wi63yRPbRHs2f4rF9IOi5RXTvzif/RQe0RDWkL9cosEMs03848R27LH22FEPd
QYYwHt//BPnRw9WywOzXR3/Vxdh8pj2Wp8Yk8Kwo+RklhvJxZDzFttEyyFZe6/EY1nmxzuv3Rh9X
QWuh0fQCSe8baWs3Vtw6xmdrVHShFtWjRkusZm00wTBTFiBJFl2BG3wEYMwfoQWU0SgmjmXtRISK
vq9aunS2kf46C4tl1yHRDmZwX3RPOvMEtZoBcW1w7+AmCngaL57pVOLy8Evvtv+n1MjZAAAaL48K
z/rqaiTVOBWHKMoJoBSw+QTbZP3nd2P6q0MGv28weL+RsfUPSCNASkatCRTMtVMkAI2+jchM/Q4m
2mxwsTAnDQSqNaeSaCWZ+lbLMs8WKxKCLaFszCgK9Eayx+1+xwd64lN89xriPYwdyVVoNaPFQ1NE
rII6d2lViqpBGg7WFyh+7S68QMdFnLT2bDTACIH9G8qXEa5CNbPeWfKTXGensf1/IwuRWYHG7yBQ
FaB8G5dtm/lhi3+nkzrYpUxRngavNJPjXhSSngj6i9WV1qlm9ZKywjPTqSq2RhaOhCslnybhWJCw
Xt1NwAloyMCFecqrhDoTRwjdRhIpJ5o6W0NlQ3Ylc/ZbYJuFvKc4dk9taxcksZGx077fRVkK4co0
EUcyOWuBROOsQwLaYVfltvgf+veV3W48iu8qE/phj2m2/fxdvT6ZlJlJCMIyDpxwd7jAb29AI9Na
no1LCgPp+fZzvumBexLLe9C1G1Mwj/UHNh2/MnMEDJHdlp+ddE8smX53x7zgkRjOFoDvggGo0tvm
jpE+Rs61M0NtB08KCmVGQ8GHOwNyFiTcHXEdphXMIQaHBLtNMOrLXOGRX/GFO9o5hAXnCq6MZI9X
Mg82Hj6pf2PH37xHkBkbTcNXoNXWsWp/NVLelo9hKD7IFSYAmVyanWn6aWRhfQaS/RoL29OMDB45
Lwmtmor/0vhnoFx5rOP0MN5a7514ZzY3iGwPak6YYbnvMHic5RSs71u2jBAsKC3PYu8e4+r6RvVG
Q2Jg/HdKXYf4fgfaHzUaJj/+iNDR80QF6b4edigOjbxLmdVS5UdXUqoJqxUE3WDqWf7RalXoe9ze
zsUoEuXTMEPxZkP9kNgUhGdEqZM9qSXe4xpwe74Op9obAygLRZ4U51C2ONeMU9jvrmxUBUqRqISY
s/8pOhU+HFCXezdke72D4qxCPt/yApJ+vTDTIZPat8GBmq/O+x82TsbG5ZFBXD8pdi7UlbZ/fo9C
tEYYNCNts2nWc9R9w+kK/U12eL1172ZozYk3Abv/HzP1y2M5HW5gK/gnTL0nddYh6QUHCi3OcDSX
1XZoTqwlwMq5Ql3Gn8ws/9zGrPUNo8un7/qhF/oJ+tC733Ul+0xz9phSZrNBLJoKCnBhlo2LK63U
+RbUT30D4rAIKt42BIHxGzArnG5KTXXJETxHsqYPsYTQeZdYDiX4tP97QXr5kR1nBh8LxIqQ0Q6D
mvV1SUD8J8yam5iQrrR27lzxVDVzgwtymkFKTg0iYrjp4he9zE+59E74/Z31w9vb1L3P6xqYXbxh
mFIcYp5GdCp8HwIdMkW1rD5h6RFe+3qkuwBzqUphK9e8I+gZJS8MMROa8kENkE3nr8Flj83CYDf1
T1UGw+BMOx7d11b7t1B86KXpF+kxTbRIlDhZ3DXxy396wq07/8vT0kwjSm0kuq6yGMBswEXA0tkU
DT5iBwoVJ5LGFVLInFPzsqkSThR1hrgZFbmqIx1BZ3DFswFwY2dZPRuaiWS2He480buKpuGKC/4P
GIhHeYhNcXgqKuEdM2N7BXAW0Kkyj0R/32qlcU6vJpgQ6KPmq0//ictkgocz1ka+BWSLI4ofyMgd
xhLThhtZbKMNqcUZO2C50tLdJYeTXx0JieZQPMMMd75C+VGLL9UdXUwtuZovYmhv2+Eh/NFb3aYM
sis9gQOSzrM8IKyj/02YvNs0OJRyedflvgYdwZ5eeM6K3l1K85m96XoTTdkMRGfNaqLB4Yr/fjMM
u86c8VTY/VUFbdjdBHb8NfaaY6/z7bE+dH7hJgVDdiB7SwpF8kIbjdCvLRIibzcjzeVNpJ8Xzoy/
fJbkaWkAwhqPZv4vBqqTrDDngjxO/udxPb6q4uJwetgay17m50XYrYMaCY9zJnC4HAQ2vTch9xIm
VqkpNl7zlElttKYFeVndTECv3WojYQ8zPjtkbfYZNkqqRB7GGV3ey8FfLaqLOr0LlvOCA9GJFkr9
G7OJv03dmckWVL+xRD5GgdpkZe6usWqWQHHc6/ChLUTN0knpE6UQ2BBs9mkJ0xn/3gowqpfpTDly
7nS0G6HHHbYxfX5X5unIeLz3zgJklgKf5ZNcR4rhxbaHeSgKb5T7Vz7pBEYAVkDyP6ii+M8qu78a
4ReLa+HLbhzFTWHsTog3XMtVRRVdLTXe8kxIu9+EAd6smQJiaRda9v0fGzh+Zis196whDsdvo0z6
KPD6tuQD3BduParrdDAIm/Rlm3zjUaLT77t4Xkmdlp52VJfHME/TLFUPhF4LtrprZ8M/n24a5Nf6
JqRs1Xs/wAc+2pFL35PVG3A/Uj1zZ1bKkJwgjoSLKKvcwxIlDlwt3z263NiZGaru0yW2uS9R2e6n
CEJ+fD/NRUcWlt+bm/5xncB613Ofb9e4EvAkqTW9e23LPBF0op00eSivIRgt3kRriWrZ/3xZn1Fx
kwf+Y5yHtM3JzFya5LWmb+X6yXtOcbHoBEHxgrEuEOL5CRlmmH3p22KqUn7JgT8mZuwVt2NHsxBy
9ocuLMlg7AUJWCHUChD1ki4kmH3Z5QKHnH3d5HTf5rq4xsiJ1UYDGvCYFHSFse7motW76mWSms/9
T92vUmu+ltJ9VedM4CJ4Q9iDYh85NJCXYl6ntAxbVBzj4psqXcBJoCIc9x99bgsBNLbGoTPG8bNn
VlIb1BM6Z2F9H1ya+CGW8Z6QpmUrwg5CVo5WgN357pQreMHPJsExq1BaKWhDQv0xIXPmL3ZWpCX9
KI0+gGcSNNXh3vtiaCPMbjYPbF5pfeX5Ay94wVbpk4YsXWQc0MYhm0YY9M1tZyS8Ng+6yZ2ytm6K
bBO75FpJo/jfYBE072wHgCJinAAUTzFJwBCQ1GPG/do4ITFKryNm82qwFHTeNpbeDCDDawhNvPS7
085piNunpjDztkC6HATTEaYAfB+VgOg4YqxVHYjmjaLegB8UhQThgllgtfCFiGMVL47B58vgPPo2
+fRJIQNN8rPEFFRwgyu9AbWl2yzerACN/trY2LFj6F9B4hkybmOUKOyxs8+Z/G4H8Ny+qNcsJSLr
ZG+rdVUCDiYopmPSEorKx+tEchDHCyLZuP1D/6lmk2ydsIKWdEBVOWXdpg64LxkSIm0GW+kgrnbI
GSs92AifUkyO20+2kINUR9DWsKA4eBPfOmMNV/dYJghPhq6cJKSE+W1E3uSIWzlePxQpbBrRgmwi
gDaoeBU8m1iGz3MUW4vZdySxknWwgldvlg4VWf35QCSoyYewFQQN34r5dzEmAfxKbLuEMZHbsJZl
32uw3mEsm7B2Tv5tY2Qp++stUetro84nth2vlN5z/WIIpSEl5/FwRbsNvABOqMlzlfmtHwYO2YHt
+8uWoW1Kvn1i4+L1RyGEEiRYIAVWOVU/1/kToR8hti+lLMW4+4Vh+ybRWGXYAHA2xzSXa9LwRz0L
Q8Wjb9+dTfRhOUoN5I8B9TtJ2gZkksLoash1GGphO/zQl3hERpxqjGNRoCEJsMIeGFP2KoRYSRVQ
9zdJ8/IgjtkRNUzcjL49PshjNKdhxBudoI/dh52LEtew5s6/Yt1XvyYRdr7W3pvzoxeze5bZB/Dy
C5PeMGgZaBSFyUy1FfOwpzHuLJn2Zhpf3LYf9VPcqns+RC2mOyx1t4VfHR2nRf1/bcry6VZR+paQ
QunFmkOV2Wj2XcTF+1YJFXad5wOAq+BGqV/BApQ9Yhmc06WgtY1A9VoREFK2dHszcLl/0A/DSNGN
Jfxa2dFJeQxYXm3Jiku7R3uD2L29wXqZotko5po0XrE3reEOnPUzi1AD2Xp8s/0VXvrZokPG1/si
zZjnih+ozRB+zTTsVgY5+iOI990lJYp4DGpCMFS7d5AR17cT2hj/08BbYoURROtaNHIn7MN3q0iM
7zwtLzc+cR5qm6BCzWM30g+W91zKLOrUwtVc35L1zqME3I6e/NN2jRB5/sgGY6Xsp0r8xuqH6DLF
RY8JB6IZ3NUpRlcfDw2tjykPI/p/yRFlLeGV/ZLEvdCEkRBKoVY3D8ees8+94msGOnwQv2tyXpoI
hklvwVqYGbUg//i8PAJm7bL1YolxPVh4q7ravc9yAj9vdsAaj2SoSEBuRCn4rH0o9zkHtGw+LGEG
boLPevwDTp5wfkc69S50YW6rWmGe5+qcmYPISx6dqS/sC14BN4rV5hZ4ZfQoWN9mmy7zLY83AfRY
pYW1j+MW8Ua34GnMv3OV2XnlQ4lzU7hAego14H14MV5UzqjkYugY7IMVuBDdcf8SXEnKes/EwOMS
rbFy7BYQtRTX3qMDUrwffhjcN3HKLa5BHCupENIqDBmoz0KlUrNqgGGmbMT8AD6tDuITZ9kEjpBx
REKf0XFFDPukCpBJd6RgnWdy5C0YOGaMTrEoBfD6/7ZxcWPcGGPSxmZ8SWCBHpSgUYF4hkBIq1i9
dJOKOkxyqNAgUTDREOyGSMRZw/HY/22Vybpnj60L2tRYhprusdc0cu9teZ3mfegKQpOGqsSt3y8K
aCrkRXQNZGbbFmHMfAm13AEQH3+2qM6coytM2YUSR0rkyh7nKWOCbKwEtFOeWuBPVfVf/cQUe0sV
CcUhrpGjMZYRM5id73X/WO5U8MrEaTZ3/wACyLyDRPoNq6voOPO9qsCReHis426lEHANrp50EnDB
0zHj7ALfW22f54oCU+i0UZ9ZWuH6knST8785wJ2YAT3HAwGo6NJPuYCqb57s6ge5H8oaeniBnDv5
3knhwZDd/zwr7xceNiCm/0nCyMbZK0QT9veqFmiy8qrERyx+YghbeB91p2fYJz2IcnohOM9/rDGS
3iGbUcV9ZZMb+lHWo21rTPto/LJDkIcpmxViXgOKf0q9AODmalkvCRzwlODniMgVInibUGfnzqWK
gRFk1KbBbX7FdQV5roVAZlldvB7fQ/6hqBkAoaxdPlUbzJDPx211LCME/MAaB+So9DARSMDTYp9O
q1zY5iwSuiAMBkTdFBEOqISf6i3IBDkO76sORnaaombEc02BK/R3PCtJE1j+eVfNnJj6w7U8JP04
DWRHbKc5NLlZqwvLuJwJdsCFl99UhDlTWuix3UpfZOdp6zF7pN6oe+0vpggBMG+PrWwl4CEDXn4N
KSmHfO1Bf4mGdPX6moBCqM8NVFOozd92n+enyZpU5fJ6nws0+1iQGheFccgfxje5HwcsOYeQLYvN
bttD0E81mWk5YCSMIUH1sQk2qS8m7ZROQX/tlBCrthxAbQcGIkVboDArnPxFnmF9yM3trbURjdte
CZFPfQZunKcB9eWtwmWf+LisPkDKbgE6ohuUweiLuBnVomU9/e735DMZ19dJhBNzXGjUoQfOMT45
/rtb4Za3fjVNpGRO6ALg1tXUbrmWLX+HWalrco7tOxmge9/uJcwGK+Lxm6XCVbg0DSIyPW8NNket
L66LXtZOAEyLPWwnGCQrBt/urWdg44w4hMeVaL3j9E+6w84rrUSTEaCd6shXWhCjQtd6SO0z7TwT
nnVT/T+Php6B421Dpv6oqiBIqIAm1Dqf1ehdKCu1v/K6k7BgwsDYRAZGTXEQ/YIvLftt3UV7gAIj
sRxT4wYnUB6gBHXDy1JJ+c39euXsgGl6KCWBS2+Bv/UfXCA6tRhtvIqS7akGtPTbN1FHztBEAz6b
mw5z+S2boao8208rgtymBYBH0mQGksblmW8yozrdmkDeQYsw1YUnf2iRfp7F4UJQsW0y4z8IkssV
mjpVwccGSj10xWHEeU3MCv/mQ0lKZCe2/lHggn/3g83fZjGOy9uE2GkOS8D7mffkiDqY96L8c/6T
KapxEMsvI2Bc421TMVPsR3dXSbB2tSo69DUjWgziWxzchKSOkZ4F5/S9qTlEL+goJt6K0Qqprzov
yZG40JunM6mUp1pxYhEvebnb9jsF6W039BQUHOefQLRaF95nmVbK47bYvFuwsFPzEf38VWuBeEiL
PmWqOVBucoZEF/tZvE6qZzabCUF3xNLhl3e0yzcSPAk8+kpbKE8OnUu/g+IT7JkeK97STPQXYv9O
AiU5kJ9trOGQGAWxBE54o+FlHkraouncio7eUyqXmIHvcwwGOy9wSMWK8v9qBjn/QDIJ0jUuvKSd
81+VRa4kDG3/P6oAi08raoWLvw7vL9n5gp7bRpt9dyq28l6yPDq5sM5cr/X4wmp4FSSU5EyY8Hiv
MZfVQwBA19V55xs2XJGMKYoO0hfiBliEOlrL2MKcgJuzxs02r95M60vIqz5O0iPxpFV6nQx321bt
UdcxdzOwjgtB+Gb18p/tUvK0ARZpFv4JqxWoQGQgzKbv8IW9hbLFVgigMUGTBHSYPEo69aMM+vw3
0RuUzutkKtG94yjKkGN+2C+d1VdW/0I4nNGlFndN8hFheauAG84xI1M2JvYAqvfGQxBGlFfHicRM
cjnBPIhlgrYS2Yg9NMtalblZkEHn3JJtxh+JeFCcte6csA7cnipw0oKP/WW3ZY/d0kUQUJNmv0N7
XaHx5u2SoQyGPp7JKMFMBfLoUzD9gaWizzKawvlwRb5LrGRw9ipQOzGfOKlbPCDBQ499kuEBL5RW
YJW82+AwFN2P1EcDbFooqZtZdOlDeham1/NJZ5ehAd+Ac/WRvLjRc6udEme0FOuQWsxFXBa8d6xf
5RqJj4YX8tZUCkqOJNiuUzwb9cU5Q4ixEvQrT3yFkhKFA6CD0SKaWWqukEDXtnsG6AX/uFi089cl
hlgJaL0fhcfMOMZVqWHEx8ZvpJ1GlZxj25vStLDFjBPZ1tM6BZoFhj2AeVboBDh6iUnprGK5eXJt
XhxyBswx6JOPJI0EwDsujpjB0205JmDgaS349WsGhsZFtQQTstY30BkCqQ2yTEA8B7pxPyS09MIJ
aR/0NoQdefqv1sTxo/3eVLcS7Z1py59QkOJQ70wPjcCeuuAQSqYntviB8USftCbYJ0mr8LQb3gw8
Xhn3D7qTe9TcV0UsPZcyozZk53cpm0YrWU0GF2P6du+ZHQBBxj4/t6nszD9nKvPDR7p+Ak4ue4si
C26Tiw9ub8icAlhiumlnYsHo6f8c/wG0X+Nscdm8kAh3btI1C8XlG1PJzx/dxLVll/gfYP0SfpWf
yRsuGkikQzjc3l4OthjD/OArAf+W1mooY8GATVWebEZ7yPO3hGZYv+hFt808Or3SjJobqoVEVpXF
h45klNG5bWC/s0ggwBniZvLs7OQOiStWLGKXXVfFj2vIrWq4UNSvE+U2VAklbySsSoaxpLvxAb/+
FPfV2usenBhCP3nuh3UgKdzq5L0v3Mze1Ts8dZLcPal3e8KKlQcmkl0sLWuH7kyhepSAjek1rB4H
iy4vwylGafumzy3HjzV/eObR1nqcGvbETFYjP/RLESnzYGkRGmiJqKzStrcuuRsliORUqSt6i5VN
SZW74M4Tqgn5zHrQ66/w/pwZTjz/TeuBR6SY/CEcVKqQbtzhaqoo3vUzGANCRNSRkHmnVlWuYUaj
/6E86jlCSGWXoWye78uS748L4EjsXiMG2yia3rKOKZXdmnprH/k73uWpeMAxL8w2zp0/Drzf+brT
UW2k7o2N1Kqb/Djs/UY7Ix54MZZ7Y4huixU+0FPAQDB/EFahPATc88fw6rRgQlhzS0JSTYzgGKer
R4MHVTPx6p+xnXH3DENUFJ7gY4u6gzvb6e3cP+KS/92fnsnyzuBVWYFnXI6AOx8V5AY1jR9kffuw
Ng4roore4oco9Bo71OvqcQRd4UUwGN3aD9gaJpKkB1PODHvZ7VcV3KorfhEw7ylrjsSWo2XJ2nco
E9p/xvoHNG6vZHK2inWZyvxsL2TZGFCv6SZb/J7UmHPmZiqPiaEkbptH8iNVwsHKZz92cs+U5BxO
JnML8YZwHHEGyrcF0E2XzjuJKsWRHsyrjC1jnHfNtmaPQozaHnTETqhRbHWnM8b13HnzSjKg1+ub
nmAwmkfCbv/Wd+mZmwe1ipD0rt7naUSfk9dX1Y0kqOsXy4WJ84ZwpJwnrmkHd10Bj6WlGxRkZ1lL
0EC90WSry2Vze1mNt76iSrSzjmj4zIRM7KM7LdjmoQKLQbvgNa1DH5kKDESpE2NKVhwDsVBlu8nw
wnd2UyqeiUk9veRUks9NJ2jMvRuQ0fr0ufLW5hskh3nPzofLcVqteA5Y+dsU/sshRDj5zoCFZmUY
DOzyU+qht4q1i9tqbBWQnAOuIkD5hsVhaFSbvN6vua+8mbHfeT3b/Qv60YTienFG/EoCVs5hdbMz
7P2YCoSIPD2RKIVxADOwZKzzEHpUeW3OTjDkMfAJnUFhwt2+J75pbkefW7b7DTwCnP3baCdiqJTc
mg3Uwd6BDCET/Y/zwRuWR+U28aiaOf9l1foXk3NfVOzyfwZ0H5cWy/0XsmbIKgDQuKxwqcIlzASs
+w/lqb+wEPDycO84o3XUm6LB/6osMImm3PC0FFhFX5TDAucN2vIqXQQKs1tXMui9DtPcmC0/4lUy
c03GrfPA1dfXtBh0hBjbrL1zbiI+jkRV+/+yJTiNbRAZcCAu1YVyOlzorWkZ49yZIG1er26ZTJ8V
Rb1N5pTZ2dY1c7LNagArWIg6DClRT1nsiced+QYzCN57yZLCfRuStS2WRK5nOZifkO2FsBMUivbj
1U7AkUZDVPPJbYbsVt2FdOoKQ9Hk9FNWc/Eyol5wPlG0IUFtItTr+daI4XocDVn34K2pK8WAk4au
h1qJhmBCVfwdwzcGsI70dtYZim+p3FsmPMaP/akNBCO319t12cVEMtlRHG2kOh56ggWkt5Tdmmve
Om9YhGmzRf+9JwLKb2L9GZ/Bks/9MTHHNZ0CX+jiqtL9Bx0kVcDoiZikCY0wZd3WKbJtcYrKC3Qu
ccDuUyFM84pNwAE5vGQ1m7DZtD5TzZoI7I7W5LhbhtgSJ5RwAfclphKe5Qa1SVHS/1oeN2oECPlt
QORW2IUHY8eCDZpL7WNlTkrLC8FZzoHISyMoIQ9yVmG3RF8MQPCGb8T32snaaYVT2NYbwzrQywsT
nPUiVm6WxJkRCL6OAx6dMHyYYWZtaqKBJIkL4nnjB6bbd4kW3Zj0MnM0NxIrhHpLuQk/PV+epw3k
GrOUEzrZhqpIRS6A2LojTvkyKlcLJCh7lnV5VW6F8sZ0QRF4fj/C9w1XA0pl5cGaMTosxmuLhbV5
jsM24FibJsPptG6nQLvHcrxWTX+JrHuoWFUcE4W3UQopzbHuMAufSMIq9TmS5/ztx6fS+OxNDijm
0l+LicBPjBgOqPIY8ySZ/wLSeOWZuFgcstj+UEU8yqXZmMevPdTRMqHCX9Jm2AVHR1uGqgaXUYg/
RKUhRRdSJhu/pau+O8z+237RXItTWE49ln4zWzTsn2z7djjgQZaH+0zdtra34q7z7uEC54rgtwdA
oMoPtol8vM1ZMB2m3Exc3dFvGD/7/FmiSzuzBMtlXRayw6Qbj7RIjsbIrjgqZ3NBOWHKCpoSjNBG
pQsOpMRy2Wb8e3EnX+0gyiI5RYvzqbsDWrqPuciaplE7aqRYNQZTLoWNyIGe1qiePoEAnQCAofdh
WjnZ6BH79/pVxPHvckBW1FplArMD/4KFKGmMdNRPbb7/EGTPbEMbNuG8puX7q3ZLPhJoebgKv4A1
TNXi7cB1UAmvdiVoFFH+AL6y+DQdz/EqfTr4zhHIuLUg/lxbK5yJp6AwtXfJNV9xukBU55R5SaLM
86C26u3a2sAsXCQi+rKUb/VRAlYOGxmFRTu7ZmJbRkeYvlnjlyR7aLdjp4WX5pg5BqRhKx4Fibja
xRHKyx5EWDgIXhCNWywoLa5z3rodSzASMdO1T+4+ANZMIzB7jwL5yW7qtaXV2h7x1+z/eRSijSRS
8LlKGj4iOCvPxENIlY5hT5H8cKUsGHcE80zf0MlqI5gFthfHYwHn6in/z4K47ZFdqZeafxyZpJPP
kUpbIJL3+rOLMKWvoTtjLY/NNtcDn7pMmwwGG/C3NZxQC4gc2+f+PjuefFF60seGP3i1RQz73DeZ
Fu72g2VNFeEmVB4vCRvgSSf0pWYNeHamqVtgikOH2wKBYj+c5cbB/8Ze/QuW6AV6vjzmlPCMn0Gs
0KbFGpDz+mjp5T3TgF5czgWxCMZWnYW9TxLqs+pJq0oAnOkdaDf0YNY/p4mL7cJ0DI4GnWDY8Xmu
8efWqb5bdyYlOzOPjW3Yz704dUX+heNg/1oEJjEsw+VuenS1BADgV0SpcP7LDr/9elegAYY2BKVW
jxOSU796LwyhEGhVtnN52GWm1QoxaP/AUalLn6qk2nnVN3JcdWa+mHqK7mM05jvvefpvnTpctLhS
Zevp0/mCTWd7iNrdRY0ZQRgvmadoI6lECQHcU2YrUhlQlgSliUH8Ig1AhDovEuK+xeFap/3/u6hF
nuwGY0N7fPkIsNST34dBLXhCbzaIq/mkT08dr0Qly20t+/LTM9KP8RmKvT4KB3/d3GLJyS9Y5Mw0
rzYuNjHLkbJYuFq8lXs5AX9nxzrAzjRo1HAfDmwl+mmAlwS0DZI7gt2G1OEV3NQNKutC/dwh+gX0
cz3m7zJrg2QOr5EpknT6U5903hF722zzgNtKX/koWdtr3XNfByoAisfBEwRPM3TcH8ZnN71vTuPs
d6UFT4onizSJrlbvVkyVXB2xIfeRXbrIp0CJf3xj766mViPva8CBpSGnk1qcrvl0cgsEH6k/adbA
e3bsAGCoH67H748CWepNPoeJFRFq3UyrZJ/IfEttjS9f+OAucnIuwxzpbkjCFM1TSnP2F/znpDM4
6hdW4By+d1NaFj62KYAkx//YJVwxC4Pf2q8fIOZ/xybnD09A9enuPpQE24EjF5vM48z48vqfgcBs
tghRT84AkVyBp9SjmApeGdNgW8Na5j062/7xAsqHdJ1/MXS73bsIeQ29Jj699Q0pzgKYAfMQVeBy
wm7myV1tIBAq6adhTb/tvSHq7bgIyS46ujF5mipvKFHZWuOzG7fd3e/GCGtwfJEOG6uQvf8vFRvD
7FcnfYNbWMxy+6dWoJHnZG4vEZkVtoCijUlCJi0LFCtkhba6c0ENejU3EYzRjCtpAj2KXInC9CgW
vN4JtpmsWOzpBcmECzNqrt+GpCNsKL3IkaNU0ABFabMx08RTBwXNc7N/oiTGONiHvLlYjxdZXwDm
m1V/2ummSr1KuDsD/8tIohPw9aG+5zbPh9CNqmVM/7zdre4I6+H7vWLt95lPsiCeOJtuUXevX9Wv
xHqxruJMduWeTYCYVKZhqGFWBMgndBZIsnkBk62RlaesO10Cld6L47yJNWik0GbfqnSAgD8AWhtQ
NEIVYI67cNez9Vz4xWNRGw+L/dulSha6/yqzmIka/wVsBu341kQj5ICVUG8PdpKs/kwQJ3GAkJwp
gkoWsRLAhTcDn32xS3pjjTdcddYA2L5FTUbCiF4X4YRWU+zPEzL5wQ1SIAO/7I6R5baYCiDp2RoV
ZjMCk3mzjUMVNSmf+BKoUlUc4H7uaAGXzMarDWPMFW9XKLEDq/l8Dnq3ebasfyc1bcL/JihvdsJe
B52qOJgCLx8frCvkeooYDE1Bpp5+Tnky3917NvUK3H9CnuqLBN7Q8nOI3QGQr9KLSDYqeVJNc3UA
aoMBnqmJMZHdpdUvHUhAT7OVuBhsbG2NYABi0+p/nbfmUAz6vDnaM9WzXJun+3Z0wBi4avdwvE91
aDs9itTQbTMTnHGrmxsO8XvdwY1bMOyl7k4podYV5N5fJbYT0GU+Wrckg7SP9t67oxRPlXq5F6nR
hwA/dsTIpIYKzqI0pD1o/QjkXjxYqBs3nJSe0ndfcys6569eHnn0MKwSvzn55vZ8cQX52ZNUdm7B
utXDkY8ZtCTtC1mLwuQd4siAbD2baOeFOwcJpwcE7EPNKvTzeOx2u77IsEkkHC2jSPQRq7MdW+9J
WxvOxehZZrKvoSdHW3YD5j+nDvTAec5EUJJRcq3ICaiwyPhM+3KygH8mxuVu4dABVK4uYQ58vkMS
Sfm7KtZu1iB24mb/hYyZfqImKf1Je9IEua0Xf/upd6IRSMv4+JthcycAq4GlewytGhftfnjOOSd8
YeX+mgPatnq3rlblx1YA4/nb37FjHuDJYSkGPD1iIKhyFZvQoUr4oyFakR4SKcLOfTkuRgASX7jp
o/XFUoczZpD/ZFt0O2Vq6w2lBRg4ydpmjCTGJMEZRFbHfNhRCp5dLO7Rat/k67ScnrrSR6/L3VuY
58PSHnxDtpOiRrQYKdaKRRfoYRpeSjRonSzhrLefHofKmLbKB+ZJEZcGwvSjWbJOfJ/LSfY8gr8n
WwTFjImDE49wQwUjSQpWCs804y/OHGYLmjB5zZ8z8Y5L61IpryNuWe5htRo1TYTpsxFKof/s6WLz
0T3u++FlwOkYHk2d/BtJsqVwMHtVw6me08XaHfSTTCFUeFy7nLGvb4O4b1s0GM2RP0xNFus29nmv
3hULSRLJQUxIZwRudbdImaoZxRck0XnlKPzxdXwg8v2DtTSYVK2ZRDKwbQ8gCKQAlk0NryYVoF5i
VI1sc/VkoUm1ia/NG7fNk1Qj8PwsU000CKzUkw/snwPSPHRnTGe42VLfHW4eXpUXCWHsk9ah3CHk
jGOX4OJW6ohbzcQIAz/DENgUM2JTheWJCeBqA3NZqbSHH2iXDA7UmwgVV4bZ0RmzVFrutx5ZvmCu
MdGuSdwtQ2uA39Ow0e9cLGMpw5EkdEKIvDnx1P/njG25G/zdtNib3HKrJ8x7f4uZmyK6CoSls1Ln
2bk+zam6eUvQtSBT6lPjP5J7/25F8x/UHqUt3U8azZvjjMfr8tnDb+uCG2f/Qud4Id3G3Tf8KNMr
eTcjlZcfsqQGNvJjdf1fs6uueb0TbCnjn6P7L7+Fn7JCRfpzQ7I7UY7GVZEJA1jSvY2zZ4HEHwVj
h/S5BbxRuestxHKfKYxIV0bE0j+hm+WpBy0yVZb5NkWiBuTbDelAPvuO2smd0U7bayC4QLPDAbuJ
50hWAN+ek3lBsDNUSNnND95oZoUVYL75/WAXBCpTiut7UP5X4QoXFgu846RSHZWHwqkItnLJjW48
/WQii0op8VqDpf8NkkHlzdidy+fp4ko4Jy6OmGVfB5bPyLWGWEt9vB8z/7axX9zPaGS902FEpp8a
r8THydMrAGgJv58rGzZ3BgFWCTNGkmUUygNclc6zK/90ljfJkR8Miiqye/UPLtWt8P7rzA6YRLBI
1Eiaa+IJ20h12uLVEYpTF7IyROSfr2GbcVoO3I89Ih7zsuRS/RB/v7OfqcLqVO0hPlNljGrPLjVe
PUijeccgdEu2fsQd7nruonAbypq9JOb0H3DomnJkLxoDclMs4DRvghUGwV7ZDIrD0cFzCLZb3C4X
ecCa0/0cToUQzsh+FFq+4P0c9aIQ28uqrMEGjBHsJ9koqktf4hP3kfX0xUx1T3LvhxObhWhyafAD
+qierTLlAP+05ZqUyfLxkqJWzn7iQg1tBJwFesFccRenqUh7n6vb/JM7t0aYkuaDMp5dJ4zfHLXf
9fEc0lKaqQYJwSgxdGzwYCdgMNUEDy0W6M/Z6rjoS/DRjoLgHeUAEE59BPOIctZlSqGBSu/WZP65
LDyWgOK8JWr+Dg9yVLqV4B4Vb8qTidoWHn4u0vaGo8BTv8YOXJo0MzJyRfYTccmY2ckl8+e4FiJW
cqI7BN464aZeX03u+mzoUXb3Dy0KW+eBJLafHt2ffsLNp4cyRaD7N1pDwlLqHV3ypygCyPzRkeeZ
g/35uhbV9OGeDg17kuKAjWPB2Wlr/zjjAfJp00TPAagEX61oBdgoM+4l65M4j9/ZWgNhbcHdnGP2
+W80Gx1AKCFzQj7BjD0h+tukSn9NdVTSVLHfO5xY5oHvcGil3cSftOBaFhr9BlwjNYwWbiROwUax
ULQFwe5BMUwhMOSqGFNCb9lfReRIOzEW5+dFpf2tcbqcHXQrECc24ghA2wUGuaOuyP9/dgxBTM9G
i1M87ISrxLddUMmD8kabgNsnnOAVi7UIeD9iBM6jSGGc2L7Wem0vcDXu42JDutYcmzqSdshfkD9E
N0MskJwwXZbWxNW3JXNo4WwxT9JCrHApVZzwvX/2Dpu/qgkLmgCV3S6gwy8KTRgCm0rEEgC49Vnn
ahzHPASoTV9Euqnw86WtultjnehQTuNrJYDxIgbNcJZaNh3YUtlhcjQRDvsLHhIRsy/QmTNtMFKZ
NA4QqCoHOcp/DV5NVibwtzKSQb2lYegafQ1JYUAM7eXIX7r4T5W69sjTgz/511fGGhYwQpoX8dNt
zaa0OCr6iPi0lWYL3Lfbsq/SKcuMwFtlDq+YvuxqAHflKhcFv68EEt+mbyUrdVebNk4KuPHMtu3P
Lsxz6JofiOkA1iLrfiyNqpH2D92wpSeSULMIkKwIa4lns08kSRCfc2POGrBCe4vXuxfD7d/h85f7
daYbXb00H57Yi1klxUKLtPf9n4ZeL46fmEBDY6NouVT9GJ0vu582iE1PiVN1LZ+q0GoixwxqK35a
44zHsd1IrE1jUCCurZ84Tnu4veXc7VBig8LYbnEiMoIBBJzFwiKEUtE7Eup+KalI2AK8uLZFlaXc
Gu4ExifmmEQ49l35AV77d+IiuAyD/8WsdfzPLWmXjanl7KAPC/t4/6jbz1CD8Wb4I7jX+e4YY/dr
vBYk1oTA2aGGGfjtA7UT3SWt5kM8aJB4sXKgkh44HBfzN/vPzaN9agus9s+CcWH127fxdRR1ixCn
8exBQHEnseyDYu6TnO2TBO/BmRuWf/tabrsYn4hEXtPdqN8GqBPNwF7Mm9Tf7cYVIEXNKtwKL9gR
hB3G9aMe0D93W/0HS2Z/lcQNKGVmTtJk8RLr9pxzbvgAScKmdPOmtsa+Xc5ksKwixnZTOhJMjn25
/gFEOceFnHbnISzSjIUtW5pZE8/8FSi1D+4lqcHE3YVJ42pT7EHS+THxYtXaNPhtNbpvC+umHz4x
wpCgRAGiJB6weNwI4UJIDsessO0nJttOhA0RQ7qnklxmRCwPdguh+FI8ym5NKhhKThRm9ddz+5UY
tLexx4qtvNnrtj8dYF5/bWatNG3ItgXOgXSAIEvO5FWWlHNyQ+SKq4CuDtNNT+XYpq+p7fKcqslM
DuAfDazyDxz9WFWH/PFxFvvVpv8np7MeeaLh7JamXDEv6kJOx2V3ZKq7TSggKZeYFYQBQqtmwE6b
ceZswwiE7MI9APf79rOdxeiagMbM/0JYzUIMCV0GmWrBt3oXtfz/aBPgF/RcEpxQczZhFDw6s0We
mlXyHE398foVHfqOOE9ls3kzk4ZtjLru+lxwyseOcbvrFxE5k9ggGpymFEVvwcix/GzjT4lfY5D0
bkFzvbL1NpOJdZUfKNkqjJ95ETxQB4QdwCIfG/rDoNfefnohbdMPXQZcJJLvJ+cQndSykcD8MBAu
UqVSmluNt4yuT1H2xVQ8ZXziWhzlEtth7/05fLnwqx/HZ1aFssyzj3pE2doiPYhIXENQkzNfzwA2
k0JRdbmfcbQ4IZYo5b99IRInnK/caTxFKN0On73xe7eMluUXEbjGrlz/i1uXcAhGqpqfKc1VNU5R
A9Ye4PT/HQFac/2Pg0rEqql4UPvcnEaHl+vXCPj3gHcBcFj3sNwvSb3252ndDj7Et8uelqYMOJud
FauaCCmeTNY6LTMY/0UssC/TXfF5sVwretPrpsNjL6w+RCAhiV+FPfed/QfklakavczREpcIcxNc
Aj+U1XoWdZ0erimZwKXPguTbZKFcGx9uz5bkEp11P6shRgH5r4fOj8SOnhdseANStF0lpZgVr8U/
ey1lc212m4KAdu9XLxLCE/SHMFUT0+Y8j8kEKogEnwXUgjRYJ2Ye8COGRTXuf40OtyAh1gWCzrVu
yVlFRJRu6l7EwnptkrnZCth0zWKGRi0xMHCTLIrE8Q3qhs5Ug+axDev8wKFyznXosvf8GHmsD1m/
7wdMdAjzkVm++VVjq9el8CHLUIzIGME9TjdMBTyrMOiqC0Nin7ZpkfXyNt0201I/fuY5lHNWVHG9
qLblgrRrm3gIsW73P+5wATtTCisGhqhut4uYYgduJ8Mm2bvDWjK3PrLLzh5mnzYa9eX4V7QDTgz5
puCR9KsHAoBj3qoufRNFR35YaafzmUJuywwoJ4i9qvk3WXk6RK/E71VpDkRoQ8EGPjNfKhtAWD7v
lxXYx74Y4/iwpdpgn90E51atdI7wzIbZflYjByt2R9EXb2emMkRhZXh0fgX+tl0IWpiaNdwnSO/o
LXe7w1cpMXL4mGXoKxKIspa7WXEkVMV5NVU6TfGdyYsJFiYfHyuYWf1BXe0ELaZuRF9Ooha9sT3J
kHZb6z2FGmvP4QHy5vUifLfd+ly4ba1cSzq6baZyrBcKLtfzWiMV+XdHlQQR7hRFMkljgvI3skVh
uGUZG+UxQCQdQXMGn84u13DB+PjN8slz6qzOe6ZDeepusf3k1BllKWBNyh0I+caDuZlnhsMDs53r
j0bI8ZF+p4jlyb+ShdtQ/nCihpQuPCZ9BXJVWuQIN+bC65D95tZIY2tFZvirYdR6LbiO8mzxWUjo
5FbKvR8QU2e1C5esDR/FHhRynLsu8W6aHI9kYJqQWsHu1gYtiAx4EEBh6XvAY+tAjPtwAURk4Ju6
mLiuYou6kRicq7GxBnR7xlSIKK22wC2ZmBRl7R+h1rbAbFXYwqFso3vFyo1H7rkZ3AzirYCFjAi7
18nn/UgET2R1C/j7AZ3L75CYf/lezgJEiqRwx+wqLbSDUP7K/wCbKWpZZT6H66L4iWng6bZPzCoZ
lpsG/xuTfiQV3DzX9R39jrBGr08ibETAyFMCnVrLtvUtQnyX/Dka2kUCnodIQHexxuI5Wjp4xpAG
B0Am7MkAgSPMNyUakC1rvwUf+sAITbIn85fkZrmbF5yguujmLdOYBDePbVTw99IVPlW5/iiF+98k
yw5MThVHs2sa6Up9AoJ1f9/hZdivPT33En07oBh3d2GINd8KKuL2AMJfwP82ja6XjQrAu8MWf+EC
2qprWbaHNgvy8xnLKDzy0mQDfFeCKQ7B3VjNpufxc9VAsnx5JxG4ERBeTrAkw0ADOeCeQNjGb8FN
GA/OBPfvk7DAhDas4y7dxwNcGppUf5j7Fh6qhlkiWKLmmwj3t/6O1/qb8xiiRLJbjCbkOgBesikw
8BSh+/t95qXb1eqBzJek+PnbTk3V1Q42lUo+JZFf8lwSTryxb8Fkns4REAt3wJ0H7DmExAVTn+Fh
XXIMmYwzoY0z2E4SWzTEK+AvRttJfnGSlpdgs6lHrhoKfVkDytmohFT9xlLac2JvcSsi+Wamomkx
o2B0cYsG5BxBLie+ZvtxMWaut7096ijl6oB74YoWz0RiZFpJier+HBbNvL/l4lJNeraWWOerLb/X
8kBZeF+4UoOcUjICevsaP2MsFzqMqDkXyx7swuZZAGtLd0kI3WGUcizoiiVo+CwUJTltk1WqdB12
Ak2DWY1dVNUeGXR93NNFFIGexJ6lCmigSlk9Ji/TUyuj77A1Cw8gDsiEzIyoi7nMZyN1P0tuzBkt
tOJMGinkJ0l6jh8T7DGSVxoHHcJNr/F5dGc6Q6Waj2OHsTLOvpL/9mhCHJe8uZzIeGi6fyGwA1dm
Mh0WPGPmbo4XDMQ0Sz7RVtp0boB4e0Dm3B1NTieSHb5pQQG6z6YtxinbiXNtVJ2vd827lR9pETaV
n0e+cYPUX9ka0zjQyha+/gRHVVs7ilN3uIy53RZfd5MZRp/hNXYxt6XbB4z9DwzHX4/aXY6ucDQ0
q8mOFB/QxcgkZ9qkkgDTzkm1Dp2pyosSNIhA+spFN8R6OVbkOzeb74q1ISdfyfD1z7spYaVphheH
iAK4Cg9iODyZtx1q98KtZDFKqhNBiheMzlMGW6XO3H586TLnCK1NrZ5JGGXTZpeJyVEv+NurKMml
OGXQGr1FAWn/I/4oZl4gOVu+fzy3n65owE0DPCn65/84o/8CRdi29waJRG9W8czmc+a32FzKznZI
TsM8duVgjg02Zodq1uxrfPP/YEwR2dV2WWAA+hjTbUvRlpywfhnaTMkWfDSa7+CWN7+RdYwVEwKq
Q/iQuNxuBL0fXyOWGSeDjweNAP6Pdp6Q2rcWnFV0/K2DR2bsOSUmwEEVI0Gm2gCIb4AOWkjAKuvR
6olK3b+FN0wzNyfMExejel5dMRv8+W1EEV+prpAItUp8BFhLuD2RDUu56fpwzUjDLBjlWbZB5yF9
0sGQJSWHu2HlUg9a35Q3Egm0bxrA3jMrCv7BeFk6qdf4PxL+t/yDci/1gix2Kkfn5jyt3V1cw0dE
KR+Qug1nQpl1I4GrHsmxCjLWAqvdB+unxzEbJzRok8I6ikjnWReQDFc46og20ej2G4AnEyGwgwKU
9prtwOZkiK0Y5QuK4qkY7fFM/4RDT51taALhU89ITALoLvpVWV9FpUUkVMWdRZaz7vIYOqsknj+L
4Af9qnAM4ZLcjMLR2w+8Z/G5WDSt4NNfIje9HIpWpE8dp9ECxDFcb+H4VKvkb1gdokqlyhD1ZkPa
9LVDuqOuB0UwkPIf5Fp/ZeNgxcclf+sHZcfvunw7TNAib36XXBddcapi9Xu1irXATgPRn75O+TeM
emHQJh82MNUSGOgzPthNxXIehCz2PQHXqN2CF+HC5AxwRZCxonu8RPhZKdDyB5k/Om+TcPi/1PHc
dRVCVIl4Dm1YKn13qy2TnXALlxg88si/Ap7jL/HPdwd4hWRwPze3ljQzTiZaCOoWOmeOtL1E3faN
p9HeOwpMI1cH7QYqEIu+GQYNmNjsiPLzoIPNkS7Z3wCvkq+EqoWakSWJn4AsYv5h7zhOk3omGp3e
Jo9fr2YSOMtwLc2ZYjlApHWokpDIil9uKlhqFHjz+fiBL2MN50hTEwpvTteGBin7NDHUwSFmEQO/
9WxQCE0Qu6L30Edt+d9YbwLYE5wbpitZz5FvHMv00akDcEC54ICLt2eJNlv386E9qst64u2N/8nU
dQEiIqeVtpunqM85cOUllL6ktNI81yXZEOdlYhh7RaJeUJH5gf722l0YvwCJYLF8O+5IXLIKWvcZ
+Ma0i/m5nNzonGSUX+n5xpLJ5N+e9cub+a6rO9KsSjRCLj2awb/A7gOSvrcuouXBTj9HfJTQrLce
KkPiSF+xtkR7/Nx+93+W9Nrbh88vCJwP/8ElQbGmFwjnjvqgOl0oS5o0kCF3qY479VLyV7RCy0Ch
SV48P1dElKqPxHbAqQ4+ZbC5JJWmKokfPsFd1D4Nt/tXmgZY8l+eEaCMsfKldYwbS8lMR1x7mU7u
m5S3Y3fVT7OWqCEtEw+kQnZcWzUX14HQNPaMk++mZ5bI00+eeb2AB1sLw20ne7WHDYc905pUKy21
UmcPbHuna6uqQ+ZZVn8ABsID59Jz+y0vNmexHun2dswzg1fJr22RqQ6PNnyIoFZS7oKZ92N1+PWM
8sshjPyYp1QM7i1pTMv27+0VYbzJmqSVthFGTG5iVFx4woqDxXxEFvsFVNcbFLqNathF5WjE6K28
pf5J3lLWsKRJVPXxLGFq1AG5OWLccf/3zkoGHwgj0MDmyJeY4uUgpNyijbVsFT4OtjRsP7H2ewJn
xfgozQckFom2xYEZak26QJLUJL1g67phF0dLrhI9Iafu0YnYNsQsvQO1I6HOo7c1i0ZaXWOeFxDB
BDAL1gPj1c0eLe1qIFqzo7yHmoDVVe/9YmHQdlet6mCg9wlSNNn2zR53lMND2lFaXPqFupxJeeRP
guJuc4CW5TdieNa1MN7iNRS+4lG03xvMJydcyS19ka/et+BiMHMBkcEHc3bIWyHAqMIjngJt33xk
hvUyINHKZxFsofF6CgTEedW87pj06b3vJn7eRyDpXYykUNiKGYUPuceZYo6NJFMYHmTJHIvZHxCK
uVlA6rf7MWY8PYfuckrRdY8/Ccu9bgp1faKygCk88IdD5sYCMga3kLl2oPNYtP/Ehsv28eDJj0YJ
msfnZXa6XwGquhagBGDtUFgXkRFT4LYmLSIQrxBMsKfRi9UM94gDb9zJyUfH6veQT4fN7g7LDJS6
MgM69NVJq5TAzynQeoWx4T/9p0cG7lfNVlsnMviWH4/5lZD5pa2isTdPEa1iLgBBqacQ+4e35DR/
rVLD8VFwPgAxq41Yw2dzyeZ5deFXm3ih4M8X3FkxgGZgdGz8XyBPczyjwmd3myGGaUChynKzQaYV
dwoQEvYIX/4hO2M8SyET9Hcpk8/Za0ZlUq/4uD3HwY7BAto1LGzuPT1yeNhACn4INl3qEwscoKIw
nB/a8vmaC0ahhTlCVOtorZ5zPbIRJLvaCBy+GqhnzarKHt4pEf8YNTvKvI/yaWgUKgOgmxRcvcfB
NfyWtPXp8583+QbVN08PdRiN5tZrh6lcICoVcBVnDvgoyTWAmSpxCrEKa3lhnvvu591nw9jsPEMD
GbISg3XyPabFSkzfbDkNOvWBsrTJa7FT1xZqMFYBb5l8PZ9w0xKuuV+rSDaoxjuufY1IYQJF9MDX
Y/7eF69Bck3IXvmlwK4TYujQS0PODQEji0X0R6Q+LmH3APVKFnR9vuEuw5sZaFOPqmsmtqs8U9gq
CkcOZrUdonE0vilVJJnGB62n7eOoFJAj5TNVe8kC0/LnOscyEo5EElkfy4Jl5BqfD9NRqV1XXO2z
qZvmoItyKYgHHA6yMcUx/lTWL0n2mJsz+fniwxUXLPUwLqQ+prbo29okt+2fUtpAa6k1yqYvgfA5
Cp5JarWjEbUD+WEJLD9t7xi2HqOSyhRgysE1sLMKfsHcP6j1pjJQ3KcQDZzSoLeh8kW12UotocNR
ubxn2xEmHqEcdA0W/HcIYmmSrRYnirm5S9XL4f+rR7YCR/Q6gE9I+BHkPHROQjfDeT8Kz/J6aJ7k
Xr+amZ3H7nCQZJwJKQOMZChVTf/TVGsCds1ckXOwYByoXriQOHDmHb1Pz+TwP0W1fNf21wpkOlAB
vDQoXfEv3AmIFcSRYol+x6jwf+heYOd6yU4UAiiWxs9+5i1hIHDtWtgC/ZljsJMeD7+jruN5dItn
O+D/gIfzFNM1Zfpx5Hjec38HucchDx+LwhrxID/0RJi8gPQPratMZVh8mwDiT+Lp4/C1cIRBo/M2
/y1Y+WOInTIMxWHvPTE8qOri13eSB7TYAAeOQz8CSuWeHsZLirlk+WvAGTbMtfUndvKLyUHsjdAM
07K7Ic+1w8U7JLywOswPou1q8sxFg7dw9XQGoWz6BaLbAnnEL/hQnRY91c+q/oUhjqUa4mA3mFNT
9XGdfzevkvbfv/4lqXRmrDtgMpDUtKpcn3/xBoehRnMY94WUaMOnR7ESyRRn9OPDQywrQEm9spMB
O4sIzTLHJ0u34/FqPHHClCk+JcFD/cQtoRjUy11ZAVBRfC/9md9Lf6DyEjtDpnnZPg0tT9ZKldU4
qp8Nis5lmOf9kDdE2kcV5rDkM8ixatehDzwtTaNh90hn5F01JsBg4twTKgqZeHLRXKr/urxu0lHE
G74ID9fN692PIxqdzRlzBeypvRQRR/LHLIGY+nQhHomoDppnMhhPyU8YC6ihg/T2t8ZYtqY57osh
5uruhnmc/nQk+toNc/kR0vfVzMzoOg2gKv4eL36/kCEYkpUy1p9h2LiYcOb+PS2OQ1732LYaaPCn
eGIp68lQ+kGKtA07otdYjuqUZAqMNt2HtddK/lddHYtJaWbAU+eDye2P0xqsPqRlkppJj618KqTa
MHTJjuplRclk3pcVpcYulARe2OnSvT1IKDTmffijQBVcHo2eAkH0+EvmBztg2ia3EXT2vcn2890U
EnjYrhZScJmz+11JBDbwB+rmIw+Jx2Lvfp9LqJj/SsLjRxAaqb1iP541jtiPijCWwW5dPXe+rcHN
c+1HfirJ2v3ERE1lv8XBKdoqAIMzuUJ6pUxgwXmu4L2Fi33VdVkBwP4z0sBynfIz/EY4GLMXbAnV
pxIxNG4v8W9Ts6gxUE+IxNrPFYV/iAKUWeBnF9gjb2k4RWOzKiMHypDsuaWP+/rNqIMJXXYmOe08
8hU9v94ZVzSaYt0jJKweHs/4up7JLL2DyEzv3JtkNUttMzKY9bv4TDrGu6jn4AB3ANeGNPKp4oS6
6h5QwOx3wk7AetaiNGnXp/qkgb4liai2JQ7rjW3OzLmftKkYyRjd8SSVslZz7l43yBkvi9Z/8qRD
EZwNFwGG4cwOmF21BJX3UPWoIVPaNnFEaEj+mGbg3kdOBVk24fPS7fgFMXtmRdjG9byt+O8/pHEn
Ry+FAJ0pZL4P0vQ4jAWNLOD+soVX6XqnSgRaqesb49dx87Jrs7M01KrJBlTjkXEoSOLT0PW0p4Bv
Bi/bou6TxKcDw+4Ik+/wsyfxghQ1UPX49C/XLNY4qc3TI/nXE2huGyfyB4J1oYEJ9vP69E1xWqmF
3o29czkvf0auk1mQ4Cl7pwWI6m9iPuczNAjZjSml1XzHu4JL/5blsSwpGsULvmHTn7RzDXX6w+X4
Pff5LhF/H0RBSPVSBDBz9ubBIzK9+ZPvMgGCEMueF22jYWpJk0UmrCuNYXIKACVlojYdFF9tse8U
yJCOg+o6cAk8y7K2haZuFJqTraIG7n4UIQrvWVGs4YXx3TQAzKHk5zkYQU139hksDbJFU8i7Ijf8
T6y+SM2OEb1bi/PwME5kNvd5vNvb2rTdc/hYYgaUDAeCt8WMqpFmtjCnUhFQYjpeL0UYOjQ531z8
pjeV5Zzb+A9Flqo4kxJbLCRAcD/gQhBpdW6PbD4emDNMNWVeZkSHcdk0IWOFjG1LwoF/RoTdCRWn
OHi3QcbVlYFFpMmaoRf/bJHUO6YYtsosTTtdKD4t1+RuAvcljEIg3vaYilb1p7O2sQXWO0WLDCv2
DbQ8bcKENEphLQ+Ai7hFh6QqqnzAXu1EbeDBpy77I/fI1pkvm0v71n2Jd7oLL69Sq7vRmlIZYY5y
g4BroOGJlKS/aLui4zbqt9reRbJ4sM1XAj+BFjbvuukMpoWUzE5Gl/PcSfFmzOCujJGzndG5E1l1
Of7uiwYwGYWhoUB0eti+UB/tRjbVGAW/bEspqDOVSNUDkuieqXwyMnOmYY3HusGGfluFIZ9f3mbe
i4E6bBHiVFv1AtEcfUylyncPO/tzeKpt54dO20s7nNJxz2lFEYnFq0IOXlcLvDcAOHBCnNpkq54i
ziQXldzufycsmcxkEsnehUs0e/Y8Amh4EqtIG9azK8CO822iwPoBrylliOj1nmoxVBVdnzqjj48x
JOy3J0sKq6wgAqEZq+3IU9lyN6HDlvMdFXPadS4lH60o7Ko458wO5WxQUEyqfpOEKNMlPhH2piUq
Ib+1jCzm81af+QCXSc1d9mXKB6bA62ctI3pgBE+pzHTA2ilN8Ycf7G4AMZyQA0SHyUqOQ7wQOtVl
715UFeoU7mFUP3yWyxroBZqYW88/pKbBQt29Geb67RRSgdpaaMasFRsCzRsS10e6CA/ygZeRo6JP
FQfXYU/+JUOkDqJo9aM8RS77HbFMaHet65/IdDr//9yT2jCo++LB0Bvg4XqR5kfSwGGPLhTNmVd1
MNWByvViQwV84sOLVpkW0xc8zkdPyXQZcgA2NVg0sUlT3xvaQHiY5Lei89Rtq0JbXH/zP9DktSkZ
DLuPx5kpyd6MQ+P4LXTsRWFy6HXVUbAWNp8LkGuS8TqV7cCr1NxrLbVUhAh09c8gLD/6GH3R+a2l
qlG9EKqiFTsxy1t+V4VGrPQMHkA5DoYdE1BF6cuHm3NNwkoLthGjv3wzAYKdIAodxyXKf+10bmjg
9BzNcf3B2l39mhu4pr3F8JgT2/mJ1QN8fsiPRul5dKYjjIcOx0X5s4kyKQFkrF4u8iE9nKwICrn6
QZZQzE8UHP3ali8l3a/7EvQWlzHI9t0N5m8cj4CTKrioTkH1p3PvBuABVPgtPRfJmADMS5KHxxNF
+RN3VCLV/+p/xVC6BR5uwGs1UGlmUlVi7EqK+j0iry7RmS4fwx09yHAL2Vvh/v8EvWfFt0jFgigM
Ml8eGpMrPod4sFRTtbfgtCJ1IkBG9B4UO7bqH+llRTIfDBwOhNrCVjZ2OkIcbQ8DN3gAYadxtsBh
5rehvkzyyEbA0sUgsJQHbhRcHHapjAkh8jDlUn/DHgCc8fL8AUNnhs0KCVuGtcwezfSgskJTh2Yn
5MLXmBkyapCOntzA9Cn+p/ehpnXICQSAktmqAQjc6qioDlLC9U4pCulZy5GZbIXnt4NKNeOB8hmZ
Z/Dn08PIYHh1aff/9b83sMcQ9B3QN7eG1kT6bt4w8mq7pmEqKbyumhcD+8NuX97RI/UKUQKCuF1W
/CAenc/IveKKZIr9TDw2YdxBOGm5xvnn3aMjrvsCrE4+o3lfTjgB/htdpbwRuykwL7jm1bGiaeWF
loZ4sdtlfVHEmFK/63dLpW1+lQFx4iLJJa1v+bU+FRAgwuujWjWljQi/RQvxBq4QKXEY83DiTFHd
Ryx+rQazEvaS5JEBDqer+pxKuRMM4BYhxLY19XF5rFIzfMn4+gDPMzKn0r9sMgYTUj7bfQnKWSzj
/YKkWzY5GdHx+bHc1udh44pn4J2wbFI/4tJpscsN/N6wUHZEk6cc6dGHZQKWecU93+tBNw9teH/p
TOgor+RpJ0S7Mc0Q6cLq5t5w0Uq+5gsknbiS6BAyO8xsxlH258RR4S+pdYlyvBStZCMtuhzej5Mt
+UXGDuKZITAJP7rq2BmIjID5CLxHdAq8p137mhtWzKuZCNSaJxLAn2v7rq8MD/rsUmPw9jdrI++q
CeDiqdCDXjVi2FK7eg4nS9cDssh/2Udvnv0KmvJyzEOzKi+mLISmH1gV/PT09k5kWaTYaNuSjjp1
AzGliNpYik/Ct1ygX5f1KKBshq71E9KI5yhppRTewluiPN+LKS/XfiT1LAJ/lMwx3HiH4DysJYku
VWkib5GSs/lXpogdhOXmW0Ghrzqp1mux+22As9CBNxfsYMqVrKRxDjpCVeAoOU/9XOLve9WVSpK6
Mz5XB5HZAeq5Kk1GNi2KRov4iijv89pS9MyYT7p04GW56/SatO+Y9eyRlAtvq54H6UeBXBtGvv8p
kYbtUqmEkiYDjwE2XqN97YRoAup3rW4twoE5cZ4abvVqKyWWBje8NJES77vouDicAWCTTRKaIA==
`protect end_protected

