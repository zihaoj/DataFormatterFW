

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hMTrOc8dD18HaqgWvNmpZ4zEm8bBBYbUJD8q1/fmMBemus6deF/Rs3qv014OJsRXQqbxa2hesuab
yGLKKDfrwQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mSxgBrwgtLA2vAOXwyMHrrOann/C22f5E08+6DMf0LZ5hAU9geZ/0xmR5kvqfwU8TARik4RxiMPe
GoOXyLsOMN2W6UkShgCGCLgANK5tzZcuyHx6Pk44yHLUUpuKg164L+cH07mc8cp50IJTS2Cc8CtI
krKzpMgwe9M7J+GMH70=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XzknZSGCbgMYEa8u6l4dUyn/X4Z2Ja897ql7FP5SKS5fe3Yb+7ag8MRk2B3VKVA5Xoyj1B4W4sIv
+xA7HVkJ5qhFGnaIxXLQE9YDYjt7bN4aSnrrGVlnrTeF15jG6/33OpfAqBt5wFvtNlCAmFI6UBBx
g2e8hCldEiZakjnpEkpseVR8pjDgCSm6Ns4wvBhf2d1rxhnnEtxZ8gT8BwJdq3qbxox5IAs1/3kf
8FmllXrABHR6vNYYk5rBolu45OEDwNVpdUAmx7XYQ0k+W8iaDWMn5o/uh3S6WXr39B+2eCXFKqG+
CodlyF+RZCIldwTvMX2jtHDrcF4VoJKljv+wTA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o5iRsFqM3ce7b6T7svod/88zc9yVed0DgumWVLeL6+U0PCbfFWUs89gBXvk5fXcJ78wVSQZpoT9S
SMVqypRbuNsuNyeadNIPe8zTFMr+kqbvEhJWktgz8LOCYyNa8D1s6wjBMEvWOrBv9mYwWz+SfPeu
rDnf1CaEQUIGOn51rlw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I0y/MyCOFNO91xE5Xg0a1Z9Lm3XAa0vnInwPBlmj4SF7OXr3Z8er2IgnDAgtYLZRcJ4mY7izGvok
7oaOdrfmkgF09GXKIKaENYYEuxjKq3RDhaP2LPiYvfDSLbaZK05L5qDTnZrtUUdhXRKMlLQMJj9D
GsrzDvF6HP7lZrcyhXGF8/wqjq8e4mXVAV2f9wIMrK3WC/QjhRtlADM+kQmt/lq73Z+CLauXO1ba
qiyP8Kva34rNeczv3cj/jV6jMQiu0NrEDtr9UE6OwO88QpRGjMwvnozHvo7/+FaKbA5CxfncTyWV
8YdmEtExuakfJPBNLqE8l0vzx1GFI1YzLVkC8g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4864)
`protect data_block
gC4noZ54R1Qs9a3HFSI7dXKDyekcDdwM/HctN4A9vwu1QyN4uD2vBoMlU5MsVeOeem/MgrZ2Rayn
wUj7p0a1luaCtg72jC6fzj7Y6nDVK5MBk7ZKHCfTjNKUFaUlR3USjySkl40qTYWmYhvwVknJ4M3V
HdES3wBb+RkEZcQzwwQlcPZycXf5SqW+2SIWzY1IlqiHpQ7cG/Omu+7Pm1Iok+6RPpsF1oL5rFfb
EJI+Dxd2fVmKUkZvfTfUo2PqF9kkfZMl6wJQQKktOvGkV0h15DYl21pBR9LvTYWrQFYoL0S7TEo7
X8C2/9V01qLUbpA8k9CJVTgZRlmMegsmn4/4xVNNCMMzIXBn21B7Vo6EAmsv6Sh6qXvFMYWbcLzT
bk53GEE5yh3mbTpNY8SeCLmLEnV3jwAJlmG11u+XHHLZKuZ1jgN2k4zey82D0LcFKs/6gtbcJDCz
wA/TGmn4v9oeDfaiCXkCYuycGKOk94zJ6HYarA/O3Pcfl3e19v4t6rJAK2RI4dJUWVVlxxUCEMie
qxP3qfpjBVPb4BGra8DCKDJ2R2yr0WqJKwRH0NMYBcpzoNjL/mgYOdrwv8pvDd0j9Y4vovR+LseH
TTSKBIKeB3caSkrjKQfk5/KrwwLGa84t5yzTep7R4nTu/vez1TRUGWRJP6A+hPYLIA+q4jWlX68a
+BCBqauR0s9WJF20utBf3LnsSx3bxzOh6CB89FJVjPzABh+NzmTM47eJb0dg7LBT53IVd/eVwpKg
Yo7q+Irb6KjGYWlwCfRQJ4NS9O2my+C/w3Ie1bRx7SSrUdAwZINR+rlP3+M6cppBL664+/blOFKx
2tv6OJSwNX3dGS0ejyPQFWeLJWhLK7YQh+D3s/SNGqsdTqtw+C25le45gSVCMuk6H+cxI/UC7bGe
bRQs/jj/5JaITVYCk7mSEyl2jaQI//oJz2/f9lCjAiRQrcZbzLRyeAwcSvrMEc2F4+Gr5fygS0of
Tz+0uc9oFqVDfgIcZmIHP84xxb23vJNQvIq9DsJX28pQQitrbFvy+TspZTJfCVdxAAbPPgOdOyL6
YB/z8hT3KokFAXBqHO6Epe4Ta869JdDThwkkcfmd19FUtam54Nc3MwjT193O0xnEUl28Yxh9dPUs
Qflswf65AB/sNzX3IRBltrxx+9GiFB/9W8Zb8NDZq/35mJs/dl7EHu9cRhTO1tEGEoBP7ow/2pdO
PnHZHmWu62P4W60vz/jL4+eQS1wLSFwg3oLG8XAqmqlFqRAFg7Ni5BnkKxlVsbIuGuVwcdj2dOS3
fuFrugNtDvmojCFjvCuvy6JRHzoOuQzQuXIHjbeGBOCHplB9wr5syNi/acgEnXLW5wo+5IxV+6u1
TjB/nql7xnnt/30Y8Kdj+C3/yWST6ISBzVHj6MgF1g/KGUTYl36wQVerZFlJP6JEt6dcKy62803O
zBSu/o8ryWKPMDWC5ZomphFi55aI32g1nciz7WBldSo1uDCMit8hC/yOwJj5WycU44zju1kQ5Q6T
YHWNh7SHN+OZCTLxaPCfumGZKWyuOmvmNZrDscOHG7EJhIzVNRZVhG8BStz23NtqMfKVHAhnVNs+
hi+3p55pAbtmdQbnuigfk4Tg7b7YVXukT7/K+Xhi1+/C7UHWDppNKDzefq1+eBu1GAYks+5AGeOz
4mTYP3BY3zlYp/xFVRnZFgYHuuESe2jQFx/At6evepYBYxOmlNVFDaTweRm5KXVALx0+yhHiukjn
2DbpryojodEmkoOEyxwZcctTO4fPjrVqi7KVi7IiJiSDFdITNMQL7VjeYETk26JBcoCbgqpRDxvA
pNtOd2KZv5St7IptlSTyKO+NsFOB2Bj3bU/TrN0B9fahlkMxpIN1hpV70Pc7Q0YufJiS9e5eZIkb
8y8P9KxoZMAyIWPB0eDBkIYKvf5bmypMqLjxvHUIS5N1qFVINMRxQmbsKI02nw5XqsnQt0ebOJnW
XXhNASCUQRnixsLGBQ3aPSeEtp8OBtuPx/DD0NMZJnehHVMVZk23MHO9K0gpxQECb5DRHIoFodra
iw621c5+rVShS1g7yEFZplhv/kKYHY9yKzkyG5GZ2npVUkiV6Xhp8ItCN3B3Cepm7qliWOmjlljI
SB98aV3CeFPCTn+9gFF2EX30NiX0gkBAUP/7tfJOKXiNQaAV3CGwG4X9cjTZrLQ0I8Hg4T9Nl+ju
NHpKU1BFUsJyntAEPdmB0k44a7hOWw+DrB8XHY7dH0Ukn8/5aNZhC28A0Hg8j0Es0tNbproR0KqD
cHafFFzfEIvf5kftvOam3XojI39QwzAQ6SiQpvGihi0FQqF5PgzQb3AZEvupsD0Zim6ZpGchnWXu
k0g7prgYnDKllaOKUvtMyH676rB59F5JYs8/w4yQdZfFxcVChFgETFpCzXCV8zX2nEorQdmfT8qI
9o+C3GOr6KNt7HA92EF014/nId9E1TFqjkt44TXNiyX4IWTZdMNc2Sf+JQhwDZfnrFRKQrteFJUT
hyPL+IhvJXSKHT1Lt/zhMqGKulkppITzmBoNaRJoPWIxKFvq6QNaxkgY7AAYfpgKY3ci4jh8Pe3m
lz20YAsahiUs1WONrVh3dMPh2VwOf3AIWoolT30KulabeHq4TTCz+vWaNWHbFTLWBYvujQ8vX712
lkd3mU6h+uk2DrSkKyFcS4V2aLTYKcUjttO4ndo7LQZ8woW8uxWkugXi8xKRw/5JnT5la50lovy3
NNj3MLj4fjb5Iuprh2UVyflAI7OL0DKa050YZNsaOOlKVqBjRfCkQP9q6737g+5vghhMxbrlh974
haUN32NzHEqVDbpFHnDnFgq/fzphWzhI+Mi5svKMR9Q9Yvl0gxP33Kef71esER4wnBnuKdTlko9C
Vg9AacRDxFZS55pwECQbIG3vknqqktLJ/UXJGTBf7I3ui5KIvZKFdwecTuWVvq7mnGixc5+8L1y7
yVQEozdi0dnsUQNhVCs648iVGZCnDLQ2+TFswFTLD+jmzRY5F1nj1NWFFwAR1zNp/UoRI+ovjs4U
aMHhRq7gXJ2tdNiuUPs/eZqgRAMsRTuYmu7SsaSO51r9a2ugsDsOR3yATvuS7eyACu0edv+p8+b6
0oRernIcNfnZnVt5Jo6zk1b9dmlqa4PFF79HwnH6SGCsmskEmLxp7By9qIlImSIdS+JBjkWl21pC
hJfHg5H3hKT6PFQXScwdTLYLrJDJcA1fPH6vshh4P5pONXiE1gX9MtsoFK/RHyYVpEj0uVGIDmQF
7dSVaN64sClMsjmPZiSeJ9MNSkWUYWx7YYbwYHL7j2FXbCFl3LfZeUDH4aokgs8DpGOtft+oG/ms
bWknog6mUrw8ujxj8k+BFpF09zruOh7XJJCZ1XrqvWZs9b0/DGgOq2Zfm7JVDtp1E8E7Suf50bdg
4lpjtcxyv/fkYMWGCZ0h2eLs9bdbm3dlCLqCc/7iaN1cXzKVmZcpSmh0t/O/O5rKowFEE9Tp/8m1
oxrd8lq9OTdRTSZ5HXUwCJ3BDo0QyJA1tUlbGYO5Dlus5+SM3FYpaZm31nA5sDbCnvfys0ngwaMa
+9ZWJZKN4GG1k9A6j5KwDyJ97bP//Je09ekNLSu3JqKUEs7qVCmknTyj0j08HrjZGQgqW1rUBKAn
QmlHAobyjy4sJyc6NM7WLscFyWKzN+PDdIi4F36m9cwZ3m0DbL6tctjim4lWVwOcZYp9daID4D0K
2L5iYFNXjC1ZO6Ib5i6eKG8IY7cmWWZqMKYcoE66XcFzJcGnFNvEauCauigPO3dF1BiJ7vrBB0te
+8aE7XV21UYlm5gdCGKSGZCDF+tos1dGaqW8H4qkO1Uarz8+hXdCRAbPRCPJ+HC45h6w+yW+xR2p
xrDLXiAZUgDeez7pY22QKroX4E2aR2+7xHUM+/tP1KjQ5zZJ/TSVGQt0j9j4gTJp/1GG/UaG3Fwu
Q4UwSCKFQn2zvPxSLzBJN1fRXdhvkFjflhIzzqEzI3p8Qvb3vH+lSU6WRVO7ad0CZOCUbtlqevzv
i+18oU/Kd/9kufwoMNZhm14KXIaqrx+Mx+SoavPgCuVMD/zuxYUssanuUCsqnZyAgDecnQiTJFFr
0+dxuh6G3CbDQqQ76Zce/xVeCNeA+Rw1G1EctLjAnyER5PRNTRegu+esOE3YUfxXrJS/H3EIQS8H
r2PwGlLSAOC7ruoGfkKo7DvjHhKtDGdLQa3Mj4R4UcUuIP+OFgQK83Pj3tNEiLmYyh8NvnhmeZHw
v6qMEhkUC38fraKlr0pGLyZTANBOva7XrsweCMSZQZjnR/WDelQXpWTIqM1lT9/FdqROQZyYJV4B
F7KGcY2UFru8ECEQLop4Y5OspLNvbB9sxzhjIzvq+D4yw1IzO3RoI5HsSvStY3VBdyoew31UTvJ6
3+hRhKqymXOdBregFv92b85d/0d8YdFhEQxp4Tb5Z1tLGTJurlb0b2TQdxEhaL6zRCpMMuq4fg97
VbpkA0WJ6Ml+Q13WurG4f1RtqXFgSQf1qGGjYFBxSGP0OtCxNUQN3Snt/gemRMkFSPuBm4Hi8F6J
x3D4XHl5XI5CiT4De81za48Mak3ATFjUYen2jwjRi942+V6gEaKSs2vMF+ixU25odXEgXbUEP9AG
X+1on8gyBRbSc8piL/8QNF7mINNYY+exX7iROR+rtLKE5zMbReO4aicIkWW7LXlsQVIA5cCtp1Ie
Bap3YfeeqT5bjkWi3WRkruByYTyn3Q7K9qkZ+iIM13RX4GqYPRuEv7+PmIAM86wwLbxk7OUjb2FN
f0RWJj9QRbJdtWCqPgTgzEYAiKxZozK/64TjfU6vQFFZR/+WbrfrQFnIriuwpLlE37y+AvMWkSan
9JvR+MTDZE6eycJw+CzF/svLLJSKjTZbVe5ztKcsXLw/U2xcyk0KmXNk2lu8H4Y7sb01GycoGBwq
82MROEb1vlDadfyycPnH/mXf1uedPYMgIYfb9tutwB4GWp4tzOwF+ynBTwSvVwxTt2mQQEjCNk5l
1VIMaNWIKNf1BFvTMK7xdqevGlEAiozGz3SXeokbh/TG95YiQHjoj+IhvTeeEOeq6MOfsZ1GaoJk
Pm1T4WznUJPo7p01zueg3AaBujAhgrj7HDjv+Diw87mE0gVz3CSeRitUt4HKW2ExpBfcAbMMIq02
sG6NnI3zC41MDGzre7tcZOFAnh3Uf030GrNetG7fVDCliiGarAcvf3+WA3uxIswJUCZwJ1rrX8Mk
LuKyk32ATJo8EFg4WE8B32SNWkFpdnIERGXjbMGkSGosr/K2wwRSSzitO0k/lZOI05dXu6yAjzJ5
3e4dCdJyTOyNez7NE305++IP0zLMofpkbE24DATVEeJKR6OSrktjXuZQEJ8md7hDo+CKdC+Zyqbf
m7pv0RZfoERLxPRdpe5k5tC763mOYYzLb6CoiUE2hIarmS9jblwjE8JXMtBnTrel0nOO4WQ9SMZc
E2bNnDnOAPR6yMORtpIyu5mWsdWRYWvDuI7WdX8+Fy6u7/Bt7v7hHL48p13z5Meh5FCXvnPTxMId
6MNfcyDbuNfwWcg1SN8jSmMKMFVDhPdckuu6zDo7d4JQ2MxbrNmNDONHK8zoWXGpz6GofwdcWYKQ
HA03TykJ402cHLSkgXwPKMUnyHWGLLL7R7OYjeemHYiknJW5hm/b/QLkb3kwoxDzZjHm4aii2UbK
tDXe0LZms9IBVirGaHIeRy2hc+pdftT0yEpAQL1V+AgOnT1KGjLY6OTaC3W+YfaWeybkDJAMy01C
JZ/E+4dk6+ssBp8n83AjmWR5kn6d7kWRfyS1UFQT/MgN60iULi8QTN/TLNEJy2/8v/KJAvTs9MYg
JUiHFoVdGmCy6NGAl1MMrXkEE+d+pYN7DoAMyF1SS6f0T3CQaKB2mS7pW8Am9nYLzdmwXcVYKJfU
DMM+OxIMZBG9ZAP+5RSUqN3wv/ypanJTpJCyfC+EVp10EGiZ/Gnt1TJkEclzcPblEDjJIbZJk6Ar
rN4DtsWTWKgeVVTtOtpwzpV/WGhaaDkzvmVNA52sCw3pPeIUag7MvV8fQz8iE3ua+IOeJ0cADpUi
6wsIkSFelUp3EO4zvWS/ohxL4VXKrap2QqaquHC+I+nNY4mH/9o8SODEwk14hZ+6LGcllQenyH5S
wgTADs8aXkAADk/ynFtx1bUCmBQtn0joFrp2qeJCWqgP7ozWOVKsPB6DlzTkG4BSJfgh1KsgNP9N
nnTInPaqDEy0j6AxuSyycpLh51w2ggRvtiAkJGn0FRJXcDcmhqP0vcFqeqmljhC2TeL8A91fzUK7
r63aUa9VC53JFsFOCJdVCS0kHDwdgnFV+t6falS3rVlRxnDPt7EZVVZ2ZohFhc6PjiAfsj7jW7O7
OxwsHpRZ+R6/Jmlu4wdBVR3ZLAgj5f0VPaSHP7gKXa6NSYCBO+ZjmjGCBQUptATt8MZFtKwN8cbb
yvHxGyGflZhjMlcc8ma3xQLPOQ==
`protect end_protected

