

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NeaiTJLl2TdirJpB/LRMvm/ZOUDEf7GrOKVke62Uo9EY6Pcbn4p5xukWTILqeOPzhgX4A7PEyf2c
z0brjxQ5Mg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QljZFRkL5ZiWx+NL/HnRnJKoN10oKQwAcLDSiKlqgmAwOmVSjyfrHOxscv+NJS9cfUi9WZuH/0CX
OHbNw+3gPRhswJk7AzH11l8e1/o6sd19maLn/G1w8rn5Z2IpIMQm76LeaeWVENts4lMvQLlMCgVa
v7W1vKVUPMofOOkM2/s=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bVA08SnvqxGOwU+GHcL5D6Hp5TG4GMCcn9+QKdBpU86ZC32cUPgSY4Ut95ltN+wxxPf/81GaiEP/
18i4dkfbmHGs6F3OxglF/mmi9pplKDxUs87cW6cmELcydNwE1zGkxm6cG/s+Ze1IATKT8sW64GGO
0jUWyAjjMAJ4pPICB8GUgpVoLT8niBqCRmhTcdvIhhC2wq5TEivwl7Khm0594rBV3k7dRevjMWi3
jvQHZG+qMGYKHGmbs6wQrpHHwNDro8sDJxkDmBKeHi+DFSBIen/QRCcrgotmCt4h1pE75gZw2+06
xBWe+vPz4g3eOZydbGlPkFQXSB2SPDrcPm1cyg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
U5PBjgOvZ0lIcr4xuyxFjjyclYRt8CijGoTDEvdURx6zZimuPBKD/4XLtWuBL1n36IN2JjyiWo4T
ZY7CKk1XflCd9rB0FT8PKTqFxVgejnDzbWYLcaZYK5iXJ9dQU7vBLQU4FIjLjlZSY9XxeoiC1STS
bJfp5mHfD5dk0NYzuvk=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JlXYqYSf1CJZWXkzppx+sI4CefnseuGvf+ttxjMrEj/s59nNpcnxCNIBS9+faiAv6DpRb/Nb26/T
3uOY2mASn05Jlsv24BWKDEIhTTCepMO5ieMgaC60pe0dDjqdSMZ4GqktdQpMXQI3v3g16mw3Y46B
sYdOb3joDyf0PIGpIIEUZmzVlJX7OFZ2ZBNHw5oLqbQLiAFuunwoEfGFwpdKp/tzWkSCw8WMXMU3
PrQh91WUljmhEmHQfu/ARhWGgkDBFUi+ZyyR7tTBWzMEgjTOZEl4v/7fi0H6mjBdOS5tXxPXgaVx
YPrACOuzrdQmVNNh5eCYHysM3/cBroQ1Dw/VHw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10640)
`protect data_block
D83isUeKZ2CGvCzcKwysDKpLRGFf3S4pqm2m/quWdHc06FVuGatUfirjJvAiNs8iSwTjbRqhYBcU
kXaUEm6SkiL5fDQzKCvExXO2zadbm0ZUnqUigHaiI8NaxT81st+nS/C3plN5pEOYBn6YXt7rlQeD
fZQPSdF1YuIfvHk/s5UME+E9xgY+eTM0DorZLnFwJM6k8wUN19pu76xWD6Ndhebbn3DC5NtLt5oL
LA2SDd7wmhWQE/upDPEcZ/kgm4yOx/wq16bMxuVySLjY6hDbloutpG1eFUoH7z+uW88scDrpXDUd
v/80wTdBqoFYGaJRrprZ+CPazpCIXGY4KAQAmw4VJE2ymyPnjjezpGIBXBLBG4NJNz7MnqHdFIF/
kHf6BEl6TEvQM4canyxSC7sGu3R0gWJAQArB8iFuYR/9XBf/p+oOy5PhhknW8KOhKm4+dxOA5ws/
gz+Jo/ejG0aqUAgXorvx58rrD6rQ5iD/VPkVDjB69LLiO96vGu4aHJWE1UWY5Fa4u1jfVMjZkpEM
f/+3o2ZBIpHbUlG2H6VGRg/xy0fCgsaSuhA7+oxrmBJ6nezPrNhed4xZe+52aKUhCNSPD7tjob/j
DTwRz6A5SkLLCKfG06XnJyJGs8pbHVeWtqe1JntC6DEglwutg6+RtxD5+tAlhapqQNC2mHQSptqL
hSP3+oYwugfVjVLl3HAHKGgDPpkWJo4SYFiadi/PXSfJS7r5EyC5xZ+WOPLAa51ZeGpTuYSCHnJu
bRjZ0raNrNZRH1ZFmBNNAo0I1CgRMoCzTgmUo/PM9TtYUeOScb8pmnTcCHK0huu58wZzHA0l2uv/
6XIfu0wav/C2NSUQClyMfvwOFzKnzEgpoEBeUhwPkvGIk41E3FGLwn9hLxPz5BGx5ZDxHkGVcnoL
h5zGxLOVBkzkk+ua5YcUC4gkoGIQdca/gux3k5lCgCU30DNKe33P7npl//irMLrFDcjONoVSZr4w
DOluQzaevnKr1HhnO6yAzhHMpcniYMQ4Q9prNCekSkk9Ph8iX+mDqQiqQ2nLpNgAyhw3Uf9qgBvw
NEQXuSvv1tquKqGOoN3MAb0mx2RMp+zEfijRBke0lDsxeoqGBl7/LT6WSLZbA9mZKl2M3BFWauBN
zeIEQKFWL94fCTq8wykXH8NPe6UoIdsGfFNcEBPHTfPe/tLfX7+xS/7ucbrdM3osXWakE0a1FfeK
JGI+lXs51CTAivFoCKmIPVEe9QvXk7troufR9Dilb948qnCK25mA+/WmpeZcIhsPTKoZ8N2tXMhA
c83ajC9PrrrD01qSfl29goYyM0zq5fvWA4T68mBBRzH/yrNHcN0WlpCkyGVeuc7DEg5P4Y1hVWmw
2WeObSaI6iRgFyuJVL6jRr+woRvSsJxoo4JEx970oJXdvFpHF6Y0ufnATOcGAtfF7siKoEECw4yD
Uz69Kz2IXPyiunru9hd6O12ufLlKCxycjaIeH2+t4HIfhyGjROyWVilufYA1j1/pytSrflA8BgSm
nYbAs4g/a5my8rNy7Wa1V72pZ5U4NgikxifiFJtV64MROPfJ941qeIgC5LkOa3OaeHEVX4qS8wLB
Efig2s4ilDQ4du4y0t2bACDjM2GpJzYduYX1NU1oVpCCz07HwIINcyGISsAvZzz9wyP8FUpevpse
h4WhiCkrjUuf+b8WRfeDa6VdElDyXHkTSzbT1Ui3NVN5wCMlseC9SHv00xdvGXhna/UigzEZDFV6
UgZK925VdboePuPG/tIydSc0SoC9lvLawsC6EN2bviYBdZ61wFbqaZ/2Z7LXFEhJQjrzEjknkH6g
+Bwi6B2EfBX74G6UN4Mishl7SP/voM2bvwZp15p7ZJoejTT//lv1PUQFhOByhLlE7xZfAbZrMd1K
YZqXYTsExCUF2QqvLilsrVdvjd1lXQ9vh5Z+Oo45lqmIAgvpyZVtY8K23ZXXJWYlRPH46UIrMDdY
8IBjjXiHtuTvODVU4vSd2kzJF5wLy7OG/ELLMrq3gGVdINVL6E6kJQLaKWg7wsl8GQg/xazx3Ie/
h1cwNXDZx3UnfMgz2gW/59iV5AcUUbACZIehLzVyZ4aFscIXr+OLuWgcuG6PB0rjE2u97V3kZQz2
lqYMSEmZ8ucsr1eyh/LaH+4+JENurDqGKtninwnLSTuhlZ1c7T8j0pZ7YS4A6JIOph4sjLjlUWGp
PbOHMluDh0NI+wHmF8RrGy6CtXSX2GdkeYcNr9jIKJ8czqvKKbrdzZS7HlY7OzJ0bbjGhIZd2lKD
XGqY0TK2m7QO9mgv7xOPZCBiVpxZXJ2wmyQiBXBI70hw3ukIZG2mqmDIGEsQukpgBJr1Jt7XSWjv
OsEPhZV38qKYMNG43/N6O0BbM8zn9OoyFe6PcoErE5Q0gN38U+CUB3qALrO2AtxYNedcIGXqTCT8
Y08DOQvhqwd6nuk/1NT2QlFTOU8qaPSYrOzG5o/1KqthdxmCKNxkW91MWO1fR9AWm86/s1IrEC5p
xk0BmOMvwBjY0+1YKg6te2f1fBGD9Nl63qNJgRrXPu9SpEaeK6ZVybWP8h5iaP7h5TduUESZ0bS1
N8dplTRMqXDrM4C6lNen7lP/xPHEppMxFjWh56t0IxTbZLDPnXSzWWlpfiWEZ+3gJjW2vtwlr2Da
coxeujmTwUlm0wNZy7O4MJf5MXfQ/kwF/8Xk61oaubw1TxHdScxgouLsY8Sm4sUUNzfkUaiN6rXX
3YC1PMj4sUvbrnyXdPuaamuyTO7E197bU8usbJ6zpq2pN5AnVM2oDy06x3pccSoge6gjYcZbNIxR
DTBCerNRCrNl3hEyFD5wZ6YNmvedZdJIqLOtRKTUIxPEM5Nwrb6Qi/vOGSz2NHqddXWvNcTSyE0g
tTR5L/k/BI3tcKGcuRGt+aTTjaDixbnzIdmD1H3OTz6pEtGO7pZX7bFaqcIWIbGyXVlJm97Xbs0b
4C2fjjLbwJzwLqNbX8tQQy7vl0E67iAe0NevEwnjTfy3xEnJN18iV0kGYjxqUQAzdn/FJ/E6F6f9
XwK2s+vfFZSQX3y199muRLtxTJcaBwwPwOE5OYi9zQwjiTYOb0/QwONbqqz4eXSAGBu69jazsH+H
1sPqcOuBThALMFNYId/JmOHuoUW/ESA2KHCl4xaMN1qlqDyb6zIl8WLGqxbx60DvMFyN392VlrJH
u8LOYLQktG2mBISHoxtunUja38CWVBo1+GJ8DrsHVzLe05DTRq0Yth3V4N/gpC7O9I4kvETaLX6O
Ur5u97ptGXLgSE56xFauHK133stAD8kslY6dvM+EwgFBA/3x01S/A3JDNT3M83TMCgmLmdVq6GA8
ZM03bh5Gc/H8bT1XCxAJ4VyEevl6xknB3pY7lVPcLOqNK9hRYkDtnp0v3szFjGB2AAXCeSGBsdLe
8SxiCIKua1a81vOmBbIrLr1zQ6ddWN+XLhZmefLjrsPqeWcf4b6oBrXcLAp2mr28hL9EEgbyopvF
gekjcKfqMLggSTuVQhVG/FJWIYIpHzMvEmC+QZowyDr0YSxymHMPnHf3U+PXZMSvH+o5P3mb2dmq
7+TYJJycFoAIrhE5y6DqmNolNw6JJWZSqr1RAls74J2EuqC1tWQTZQ3oHulDZB0ow67iebpUiXLZ
FJc+XP0rqGIVaipAbgiPhrI45BHHZ9Bt8b5c5O2lAYYJxNdRneph6nVHjnehP1jowpcxZPMcTP4M
bFUbPRttbBosh4tCIkc7PndY8AstWn2k06nJBl5RGXCOSV4pEE0rlAdYI1/axC6Yuq8BBXme3sLo
UIVEBeSdswLwqoYeLLC0P1uaxmrUPVbwjSpBzHNvAdQqFoqZskinG6Pp/ykN3Ab9//O5MWXO0IO4
ktu4H1hAtyCP6Nd4JDOe9Y9mSuqkD7DMDoVGTS88P6XW178bJepCbAp067U3Zs+ObKSifUdJq2k6
gHDlX9gBwrD7lqZUKKNQdwPw3RAYijwlVHR8F+xQpMOxpX/Q2dcy0TPY8alSgAWAacBKK4DxHpP2
cSpzYbisrQ+xOyokb1jvSh+kMr4Xa+pKEuIPvxiWZi7ah7PQ+yplwznYkWN0sSJN4znf/vvF9mEC
mAXAOdnKtGNlqM3/KmaxGkdLGQ2lz6nPxcSBMUjOkcI5QumQzZGcfGqMZ6ocKJcYpxOVzJ4F3xb9
x4XGfFM50OSzzLnE98D77m0XGpXBO1KstpBUWiJ8va7GRUUIo4ICD4MpxXOEr9sTwg7FxUrxo5kV
VC08QxVY6UV6Lb9Y0FOetnbdonlcqZeN/C3YRtctTS9DBmu/IaFRBp48dDiZiLJZrRCuLgaaioXV
4sVptkL4b518OhcCQnmEAtAq+v4rgpS7ncYsDsN0TDing9yTHqoNT/G98nEM8duA6F+7XcEuDQm0
apUVOttvuz6ly8g0WlNPADfcg4Zz85GtLLKRzzbHyqdLKwOpc+RNpiNqoywE1ljTOt6iWf1L8oAa
rSy9TBqbFoNUUqBITTk+6eNCm6vkecbw51dVLBahdBZhCW96CwH3/Q5Q478Qm6eC7I+UNMpqFLT/
e2Iwy5vJPLe31rBVuL4ambEOrC35+5wEyAoBDw+/HRsbxZlQMGDzXOYRhegYBTutYM9vKTE2BB+s
GeVHf8Ke2NJCAywtYII+U9kT0OinJTCeXqrbx5AFIRk5p1rp7c2qptmFPZ7FSBU0yG97Z0vJ45Ow
9Kjouc4cuKNx2mruyegfCfMuPx4dqmXbh0ik43f5EcsaX1FLjYeydzKFnkDk+kgm9ff3SoxWyKRn
6s4MhUDFXNmFt8k1J5fWnwHryjgfxjlsuw2Cu/35hzXHxJ6f2ulEYm9YOtAaKTf7knfBjLzB0Qbf
nyIlEzijfCeM8plq4pSAp2vHugwDfS1Q9GH8Qkym+MiW+muQUR9IKEYOGsNIWbP+VEWelzTI/+b7
MReglwvuyWVC5pYxNKo8aRm/LeeOU/Ru7gC0gHv8B9D/KFKh+EJf9OQAu+dpiNaqpbWNQ0RA5kfQ
PZ6siFfvb7isFBDY56ucjB7J+GVnsBTKuNjuM5trDv+Spi7FuwEq5NVQ0caKtPH9D/BwO47HPAd6
qaVw2WPAyhGU/OFq7h+LK+lG22eWflj6ed35j3Mqhgzw68wE5yXdbyD83uPeB//lwBjUx2ipOXXw
jR0ADjyf51N2O6fnOSWiwmZIjgzKDtsaL1c/yn911QviRxCvv5RjWUJkmTOnYcrCsGYlJ1R61dNj
c8YL0ZDn8SRd1LNNyHT2DCCAC/qkfSVF/p5+Yg6XGz9JXM0f/4ikjlOawt8T+bunbOX5qrpjliqx
h0tM7tyAYYcBQ80ZEohL1h21XiI1HSdgHpcQlnx4ncs9OrgyUaYNHp8BTGRVXRrah5ku+LlZ0dZq
EF18JWpQWet38g/l1KwaGEyXTFFYE0tkQh5IUzQ3MfmU0HZgtFQ5uhlJIB58sMg/dtGgZWC2fwd7
ISHDDb9BHrCwnCHaro7i4mxiccz3g6Hj94NbDBnRzaiyaKp8ajCuCnfBgzrIU7GPC5Vk1wT7D+qC
BKNzv9l/Zk60wDvI4Zj/qhczkvvv0H+62YCyYL3RM5kknVm/Rf1yvuqY/sssJRtTAaAGw6Vx/Yp5
yoedjhOrIstBb4odCPpZKZdZCiRNMPlL8KkIkTmbFhBf0CioZKOHjdc83i1kG9t8xjVuI1AFPWA2
SKUfS468luBAzbdjlZ0abv6k9T41lWTOKOe/qkM5PHLBOHmmBOsjXbU9EDQoxqY1As0cokwtKoFi
nr7Fc7ddhGK2H3ZIp/08pbOC+YHYLbpvWzYo1tlydGJSXXqQjG42FY0hTvUBwsIW4qnPfvTHd9M2
pjHabIe6BGH8TvrrX66ADSPnhIcRrT0ttre00QYNJfqhZX14GvGNBEeGthE2T67xGpLXCBvTUJjp
PlZc2UT93At9wf64v0DGGaiLsgZde2uNe3AeLBpib2vjRNdh0f8lKeuSb1yl1oPMbhWolKAxy9lR
gtQGH/1nuG+62B0yuASuB6zqGKcXBk9psl8pzvU1rHTk9ILvy6iAzcjzZ2ruI6c4WKS8U6BrR3C6
M2hNbOao6kx0jWTYx3VUBaDlI4l0RplU84gA1jlZL4Out60EsM43/g5Dmj/j4PAxXyNqcff6T+XP
TWykMkvOq3FyyJpnxp/uPVLX2cvqd6C8EXTqKj/KuHWjX79aeIJ4rmnCfv9y8p9DSsUgQHbF1xWn
HPDxikrWk3momUbbDWrr5wO28qGOEAjxl5keRCEjlFlVIxo9HKTgGhSGitlGtt0hDBOPU1AFiSMz
9whxPZKbDuRfES772MVfqHGi2aXb2YJurk0Mnc2mG6oUworiGbpqrpdRvg7aeqr9oVC0DpoBpcQW
Fl61uLfN7VrrgOYI0+Ho4MDcmL+nVrvIztaZbv2bkwPZ8s4FPUV+QhJCmmo2xl/TyoGFQiM+cINi
iL+ea1VceD723ezEvsGpnhHWq1RcNsQaMVjqJNBlAquoLd9KUZ/hQefyZiwPatVy2nFmADQL7bZg
2Ox8BPW1Rn950uhf2BfWY0r/fCEh/fdgyLLHJ0Ez0wa8YRD+3X09yPXorZdAVAsKdjm1xNqw91am
xzo1xqN4D3CXHlwH7iXwQO2rC8nSCY0S/fwcvBThtIHun8bD2B3Tqkr5SXBypY4ETq/XXJV3/ZZt
NEo+tNDg0i2dt6rdPqzCs6IB6uP4GGp2eQBLBiL+fGpm9ST3Xnn+GzRMRLbIGtHEWdd7l4TDO09/
XOehuxTElJv3ZDx/N2f4Thur58roZgD2FJdqxs0+hraxypVNDWgK2Hwe+3VaACRfcMXTuAAcgibM
pE0m4TB0/MIg5yspFxP/L1MN4cegRsUTtb81WNYszCgAtpqnZyvliUIo8k7di+y3FlOKTxiJIJ5w
PpLZhhNj88aXejCWUfKP9Ox//ng6PWLbyUoCX9p2prZuiN8fBNsSk+xix4kEz6gMQkw9adjNrYQ/
hMdMu1QEKKxthaAxUpKTYj0HpS1c5pz8L7Sk+lMf68GVFYBw8LAi9YSfZqeECXoOMekfFjUNPsx2
tRzo87fGiuCUHFfRnK3NfkeMahPTK0FjiVwk8VlXk74R+x/+WNc0+qui6q5KzTMhKB6kacRaadbP
gVvxvObWlqBadrfskCoDzpxagK3hW9hhpH0riyi1bWjK6ntgvhnkwh91/RFIQaZBtvObxli9DcaV
jJLnSckLof/iaYijsvP2L2ttDDETKg2rx4WJOaxSnLNwkT4lnJbuh1ceblIRgTQmnUHtTJ5weG2O
WyCdjgNadSaNJmd4xXyHYQDp+5LvALrlW3kQ0ba1lpdMTet5in2eotByQ+FyrKhyWAfK7eZgcuRB
8281muot2kaiTsJlmG5oI3WsahMdLamhPkgKqqrT0kWENYzXQxHeadL9pklomUlZmw6GgwFqMxcX
GUs0ELE7EfLXQwTP+jaNEWr+85JzJm35x8I8kOACsU0EvlHvzTNo0zeCKIofe4xLVE+xXbPpKmyR
kLoxge18oGur7LSU60tJYVIDaufnzdgIWfv3i+gHbm+7VK2ebpcmWP4kndPNnmZvd1kCBWuTbn+n
9+143FV0MKh81OBCHBfDm73SCVvy31cAg4Aq7V2oVoicgGxKAXLIAk3ODMROCMlRTYn9Sfrnnheg
yIDlckiu1fwiP1evn0DPZy5YLS7hbTpg/eIVigfzcyCb5stW4/EB37MO/HL17Atu6weiFsKIeZjh
3l3Hy3ekZgyV8yNzddBYWTjlXVKuPoMziDqDCDUvKZXkfJyTE7eVVJ9ZhscQ1WWl3zhbblYerGwZ
rYjZqlHtcHyI3rjvZ52Y0NUZ0Lm1LtUa+xykgFDJXWdI2o5djMreUv5Ny/zUxSuKBR4xs5bJM8QG
H1tHK02fT92CyVoAqPW1jwRufZ3IsMJeSwR/cOH9kAxN0w4k/fO1IKBNLbZSBum9MidRHx2ca43F
pJJGztHJLw/dTD9LaQ3dOY9BKtORR5j2TUDmVdjTiBuJIxfX90dkPQTRlo7wQIr5vfpyBjLVmzxW
8pPl8ZigXpqb4lBmLY7PWfP2Q6CiE4F0jvR1A/8yD9bO2nmjKG3VqJpXQN4dRv4n5fkifz6wgLcR
6JP2eh5XPvRyymjxW+KtXiyh42Ut2rhMHTIEaao+UmdvInGn8ziuzjdZvBhuLgnix75CEfGZ9/Ha
yZTc8R95lbKrab8kbq1NNRAp3cFMSNiQe+lY8i0rLwvhYTJF6JfwpIBvUIeg/VvkhFXjJ1uWCey/
5qSkuxW58PgMf7eweA7+uKrNfKWuMgVk/diyjjG2kfytFFTZvcJW2bDAZ9+pZSoqQUEoczsumkSP
8X/JHkhQJmDk/507pPsibye1eCb3J1TOHFUhqjBW27aO7udqBEUF8qNoGCCnRbUh+6MsmyrM2coh
7wj45WskVbLjo7YesRVRYBYYlAPU7PzWNW4hfvU8ZAjazLlhPjhjoLtJBKBIKBV1dV17ptRYm75N
PTzF6aIvyIVOYPzoaPc5ODlgMl/Ec3fGsSU+6uPJ1wKO2lR5T6nmg7JBtkwD093gGFm+QCpG7HuW
H1W5Rqnozpna5sh2UMhLgMoaW0dkt4/Te/r0at19hqPMi15kZTLnb0gJM6YdlJa+dv2Bwx/qJrFm
KzFLBlQUEkuM0TYaykGDkw1uSeMwEVGp7wCj4N9EY7P9Q1qp95+ERqlino3E9FA53vPpwTd6fKwe
FG3g8xG3xOrGRN6nyGDSJPWtrBvNeuRl7wQoXd5c8R4HtDPyVgDiuxIzYAlfvRbPXC+0J3m2xe6V
/ddhT5beAqMJmGnzI1+2O5+i7bV45j8Wi0gpRvhpr1LRpFblrx8dSFf5Cn5z5UDy1LlocoDrbKAZ
k8L/ujoZIStJnlHTt2xg+tDhwIfeLy7AXtKQ1525nB47i/mWWZlhYhxSFZwhMPfXSMZMzPT0zxm9
w0IeBYnElr5JS/32I/Qh1iGyZnyg+3nxeZzVnnaex9xOdlULAwxMwXrfK3PVMHwHDL7aB2z4n/WI
aU/o9JJjKRrIdmslgPA0ZImrudAzW1wVTQ8efU8vmxFaUbp5YYYAf6vWcF15vhMlAb/BHYjidfrO
bYYQr9xWJgueocNMqlX4dbzhczwj1+4nn1hy2yKl/zpYG7yrQaoDBSfaj/DzXXRfwwsjN6lPftBL
KsdXUbkohn7j+C8EDWo3/1LdfIWLgQKppdsU4FgnE4hHC2TIWxhOsiYjXAzcU9nz9ewncmvrDFJE
mz+mcKrW3Yglld7Y2xYM7CnAvXavx+esd0f5UNAQ5MQd9M4e6zwRxqB/JToazM+A1ZG978KGpEYt
vVEgDSca6+vD/7fd3c6OsPWDEf9zmTV9+Da7r52ItCtOs2+BocUWADmeDAQugxtSn8TxfpqXNi/H
2WrN0WgcE0v1dlP0pt3Vh54dynnf7wzf0OJfUP8KASidypCGg9/waANuYU4+2puJZ2vP/T1W7zw1
u/yO8sJYsKDKCEKtVpFx6jmNmFVBbeEKkSKQz+oyKMupS1q1y4F4DlhoRZZ7/eSRrw87bbiNTXUf
BfEN8e5NAZAOdZ34ndGHNrQ2rYk9czkFTWl96ulwHeTW5SfVDkh90BsmPpEUnjJAJnsYgqA8NTZW
Jar9s0foZQLodzRWQEDIOCf4n00KkAnJSTNwZ3vR6lUCv/emtQQI0Z5ED8mzJrmGoMoYn5bZ/Y39
2hu35AEkY+dRSQzRjMMi/0+tfdhfwYptCaWxapuvOCp1uB986PW2QH0X3wE0FMZRrWc9V0Nk6cGk
GSl2MImfO4LH5altG7DJ2nn03yVRslUpH7tpFJy1Yac/geEuHxT4Oeqft+RIKYx63l/Dv4FUrjLL
dFDnPloR5cDuX2I+eOcxMYcjevGnahwjhmpFbqtazabwKtlUrtVLW3Lxn0/kOfxTfJK1iJWEDUhA
XfikC0eazcUnFySK8x4b9r8spIeYnUwE2cQ7xEhpgBVynxjM1P/z0ic1U1sTmEU6pKXMFktey6Na
62fZ6fT9Uo01VNnhArqAcyq5PmyoXuwgXSsfTVAQkRN4wgG/dOXhMpDa+4tnNlkPMKXL8jID58d0
K4kotWOfSMm4Vd3oRTPwvd+/8FpZwObhr8EFUO231vXkRJH9N6FODioTlE5zuxQXKTK5LHhsXEnn
A3pyBQDGbIV7kXkPzbGlFm0ksSD3uWbg9ZDM5Gvp9LXHCyiQ2FzhQ0UA+VA3rR6Hv1U0UQlOVTsD
syFvDh2tWC5Leb9CRh1GML/FrunUfVm+/4OMTpGkOfk3sBNZRyTcTAPuj+yJkcQC9m+sbM799kQU
Ay2iZVGdUW6nDZalzQ8F51YbTtLTAOQJmak3i113KSIyXbmHewYMANgM+BLzRjKi5enz7cXBHiA0
B8730u3C9Cu6tTX4YIGo+WLidnyIkiaH90ugtf9HEa0aiFGCcQ1RA5MsArdJo+YpuyVjLedld+UK
adgsot+AqTs1FPr191tuXU25IwI/+SY32dqYelR2j6k9vv3tPltCHKdO88Qp7toc+QlYed2dhd1t
AEqTDonDLoB/blbWBi3fDkXDKPio0bNKN7LZtH58XeEDOu+wl2CDxKJ8o18zpiDnqRDf0PtTN1Bq
j928fF2HpmICSpNQJE8xllHrs6uKXBeOoRMelQHXaThOVeLU36OhIG8jLP9huh34I7gKEVu+u3uQ
5viC7TubZud0qX1hzk7BMOk/gOkd/yhRG0+OsdkwLQcRxdDdKjbvLtV3/9VW37ARS6pSlnyS6mQc
TkssW1DpKnuw2YXZKZr1UwE4ul0SNQbZQ+hcKTR+zg0b1D95hPIQvJ/LbtrFwrTxIPUaenXa4fGN
62DT4lTdV9GPQnuY2bLZ8iq+AaQCGz9WQOPSwAxtEIq7tls3hg1OeOMesbbwZcipLK4dvb5/Zutm
Kjrlv+z8pAQRbXd4476XeKk3prlvUz5wSleizj/YdpPX1ebENauGKMwE0CG3+vO268+xBjQDmK44
flpCpEO0PRusvxm1dC1I/0itSDwBII9bzEGl58Hjt06361PmL+cFht+EAbxDLawpBBp3Y/pD3qLE
A90NgcjtXw9jNbypTqFMAvonIKrxeXN1d9DYsQpzgL+/9RTmHH/x9wwZ9zE7HMb80o3DCfNtqV42
Qwhh9pTJ01NTl8nbCsEvV/rlfynpyta/gS0c14mzF9U7VpYBPH8RcBhp0h07KrKN064jrflsMaFa
8qH/thjDPhwEMzk1DslWu1R27L9u4RdxNtN06Tyl33pMTh7CukA8In4sflXqdYQqNz6cNZeMPbg7
JBsLun12d469RIE3ZjsrBznPWa1V86LX/hslNd3uK4Z3crP0H82Nu6QASoZZwdlbPTunyUhukKcf
7AsBgvXPOIidbGMorsrBIWjUIl84DXJt0OxRwPc3mDdOfqcvpQkj69D+HhfedB8R5gs39a5nSTlz
+Uu5+vz4hFOWWGX8UqWzlq3B+Vs1AQdU670lY7sQu7USvmB74UfLrZkzZO7ne9GULzk+MnQwHWta
ex0cKhhnZEVaIFb6Fp9yyvZcPX4kMGeeLIo71siwlXJ5hgV3poEvR2uyeoQwbtA1HDwyryeDVewt
WtZVWmcDBpGalGBARAmJn6YydvEjTXmtLj6kRuJ4IGwcDEFLMvH9EsIvuH9ulHfbNaxtPoTDFh4e
Cj/v/6dlgTbHcOgLzSzrZUIN89TWa5/k6sM9L8jaDyWMNuM3K11NptCqaDZWGjaDKCTlbwGJQqC7
ZGDNRKrZEoyqy0fyLAmYF7KF0TwcmgFob6jWMeD4Mx7+6ZdED88lkM/+If2TlnZN0aK43FNSkC3h
LNnhhzfMo38gxQRN+wigrZbKEngPqvmUjRZReXmZGMyVK68WG7f9zVT3hls6kJ5/UhAhQE0s+Gx2
30jsoX0JbEpG79m2SyUKjtSYLx3kTX40oB+fIEIYIkpGO/jGbH+291Y1xhxDk7Vbn6OQE+6YHlQx
6yrVhgqnZboeDYNzCagB38/x658JtdoS//B1OdOZkNv4XDGcUGZXoYW29ONnAwAPPwkB9IlESLJM
V/VDy+pJ92HWbVsGIF2oe5yQWFWU6OqJF8O0tnOM8WDqJkjix/MujA3wQwywGURMXbsvAvl1Gszi
LxuXdMwXWWJCJoMCa9lXQMI7zkg9H8O8XwMLhjOpnH9u+7jvMrkyDdjwwDAbTYk9amwrocOsSpBW
QYLf+1e0RGYvCrRLkgJmP2JlU/wthuV0DZvlt29vShfDxvKc9iNl4iJ0OaheIovCwgg3I+55fdV7
hW/8V/guZIhv2iMaZaQsKI6vXEMYPJVwYPe648d+5UF3vTRTgh193KRmu/ToQ0ZlK4aKCIt9VGPb
yZ2Le4iUZu4Ux4ZNB2XZBCF8z/uouI0sikGO96F/J3/Dd4bCpKwelHUzE5MLSv09LTpsDtPcRnQW
pPl3E9gnT+NYss4+ckOPg2k5nRitrLfw7zpxM+EZlNRKO2OiMnYUhNMTxVARKBKALyO7jb+7jHX1
iqEjt8uQvO8Yom6bIptD9crGlNPEO8mW2MvOaD36Kordf6vxMKh2HqF8jMLVeYyN1AP719/akVn/
giAV0qvc7yO0EbVTZLprIJUsF/f6Bmc2clRz1PjYffLHCX+Dzm/avEiIvGs1Os38/uTRYF+0uDW9
2aiT4szqPEQOXqvTc8ftppN1hiRJfGBPpNqszTokfgv/JOjqcrliDN+WQN2ullBm+bafI6h49fYR
DttmzJwKVjYeXvWGhduo4CswSNgM5NyaZaYJj0Y9fKZ16s9fJkp219amRlyGsEjuDl/a6o/WG0/N
1l03nPJxbsOc/azdwRkkQl5XZhc1RuiqAUuoNH5QBj380hNs9OYYaFHzoA5/1r5kk53nYv44/9iK
9ry7AY0ro2CUTERqhpp46nB+kI7ZC2ikIpR6EOOGOksFWytAVWyVvO/MgH6UjvUneISVdL7ikgeV
RCiy2vTC5ZNvBp9408IGucazN4GvoAUUW2rnwuhej2CMW4X4ovzVPOooaN4G0eF93mdR0JfmW9kb
2gaO7Ub7nsmCBTZzlmyfBqqxgl+ryGFW2lmA38TVY4tOKBBqAW6yk2UruaRXXquNyS6u81c2xGZR
jimg2Xc219nteM1+3A/EwWLHF4rTP8EgAkV+00TcYsGRWU7XWRwOaPglgob98zMsiAK52wA5USps
Szm2zwO2p4Q3/ISyz1QVBC/weePZvrIs6dVFd2OGe4gFpJpW8mSKyWTrEt79r9mhybDNe8eU+kyz
qDozDpyShEQjqsd0GAHGK68KNiyIH5mRVsAtv8EdNpvqJP7Iw7HcC7nwTB7c6P0Z6ubcAtY7hDGv
y6pDoNwsQtZLWZhog70JePnW67ydlRO6X08ytTnm9e6IlGhuj9ckm4Z5pA79WUE2Z6UHhk4Df0OQ
qjDAGE13EXFsYVBO9sKcrFIsdgd/P5v3WRGQOGorXITC4p/DP9RS2txatH6EaPH6YoKNo3zRy4Xp
/0B7oV9GiPUtKR09ebrZHGXjCpzIeAFsIysAHPMyfYCNn80YmOvV7GLnrSDm5H7vgsCe6UbEEA0x
V6pQ9QsOobx0Ahud9yfZRczUeTWsdRsMUoO5AtnWlOy9Em55ykRLV681p/pdY2ww55dOuPLeQDfM
0ufuq6HTQ+4/xwRE7om6xtABNv0D45CFllqU4YwMHb4L1i0xfiaaoe/bzK5WmIDYvGHabXHmAcbg
e/++bm1lre/l9kE1svSiX8JE/KYWQggDkwtVOnvQ34mC4j1rmlZcNSG48mRYNlRna9EaNYyiU/l0
Ppe4hnI3n0/WqVImtw+QWMVda3hD3HqbCNrLSNB9Gi3ojPraOut/px9coFue7BpBCUpN+cGACvla
CjMh0I9NSM+7PzNDkNciOGIB5ZWcET5nRjg2WWbl5IXNdhW59lvKmGX2yaZFphycZa/uE/bvyKBf
Pxr3/lwQPsOPhseqU3wrlm/9HQ+VLn6BWQknaOoDd+j/99lvsPvRIPmbTB3zHIinooS77HlJyeVE
GWVIu2nDCHfE5pnnaj1cKR3fyML966Gwz0sBgxhj/XVVrIAzkc4xrG2A6q6Y+XQkVz4zUyYfiL4N
QoHi40nSMvzgTggU4a6qwDukec47jfvMGytkcfR6DOH5DdyTe6s=
`protect end_protected

