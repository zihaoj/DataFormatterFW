

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TCf5JGgj/7ugzS/sKy0pUT5UHsQVCij5kMFYoFTJ8tss1iq5w0ZsMUYUr3jpzKxBpD03WfXcwZSA
wetHjviYAQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UCJ06o+/kNN4HFRiq8296i5eutve9tCcrt5e2TfD/ql1IGfnmHwDww7XpwWxR95wLZ0hiU9nZmfj
Lw3s0XwfHU2NgrlFg0g32Kl0szP+Kdxx/k1o5CNONeIoyI9qzrNvwVUcai8HTb2d0mMFW5jqblFt
lCzqoWjM7rVPr35MTi4=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LEotkU+GtjlZNF3pNiQmTk7PYmxXham/0WU4S36F1R9sCsEeEKVZXi743WQ0P0GmzMoUulsv8krk
WVdt+58hcEp8TU+GzmWp16zuY+PSFGDJNbFXHyxv4RdjvUreDjvBn9I6ZxMoZOsZolEJUph5KMDL
YwB3DDF4fxPWGN1ZQtxP6hBRKtJK2HMCeA2jW1l4EizvArXE3WTMI8FtiFNufmRZrXapSnnzzTWr
AsaXt/ydEUJMd94wTb/lpbwR8o5vY+RIvoZWTULJo8bednl2A82O/igcAv+YQpt92NCRiLzvTCc0
mEBDSjEY6WrQM2ePDm5q2EQ0v4khEuZvQ4XvEg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AlLH/YgHj6mCBY3xSgnGDnQthI+brmGsURwYmiEQOK2t2bIUGrPEGqF4YLjOuzqMxH9wtbTXkH0t
4FrZS8vRJyL84tvltEegmAM1YWNuU2HKMUcl/r1E67WcEhZULYJkTt17CDGMnNnafpjmJNIgfvsP
RSUpXAbqimD9ZS1O+QM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mPhPeZbc7L4U7Cq2HPffhm6Uvs7gz7fvzp6+KTcIjExMeR13Iqd8726U0Y9I9t/WGlzGcfti6G7N
KJv7iiK42A5gaFMX4M739rF6FQIKnzLWNkRfLGyazDmpufyaw28bK5sLrHYb0zkKcZgIpFCNXDB2
+YObeA6WZXZbkxcQiYPYb+YfoGi6XgdCGTU8qh4v6JiRF+mshmKjRc8hvpIKi75csaLsU+/z1q/d
LWI0wg05IFu5WHOCd4B2g5MY4eFjpPywXsPr4H1echWFvqSHM+XniLfD3pwQFljHXjOK2EnMYbux
5cn+wIrk1WZF76IlHNa6fUvO/qFzgsHHk9im1g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3744)
`protect data_block
bwDarnSF9CXaqXj1LblbIFYSYGz7ZDZKVlnjtiMOG/wjKlTK7WDNuNcrSq7AxDZ4gXgd2XvwnXY+
u9YYIxtN1LjQ+lRn4vx1ad3RXyMzIoS+0ds2DSGyIwnwQ4J039uWENVlkxzIWHa7QRmh4oXYyjUe
xL3ywlB00Oley+s40G51ujtyrW36CR7sTtr8iSuet2YetzBNQXIutZrjWd+812tecgtCMizERie+
JRk0E+S8ahVgRZOEY3BvxQjw+cwza8Utuf+rsN+EwIg0UA/PLCKSF0cBdK3QqakmDkg8q4Gee9jO
fEAOEJTKNL2MUZumjavFocTcOwkGFkyH2/fKDT77Q8qRzvwGi7PJOIfISKZIX13lPXDoW0FLOao/
MF3wWSWZVihvF2bVh29OY9bTwSgMttDPfqSlUsrKSaX2oYiDHHE4P7UXC0C2caj2LyGjsqdq71gN
ABAVsEBoAYM9xeyLe9pevLs+zJKnfs8QvdaUAnDdOKnzfQAtLczmATBkckMX4TdgT/RLbMJ/LJvV
XgltTdUrtX0DjSbNJqKIo+jaPhOz26oqIFo023kheVVAejL8VllnLQu1ojt5qgq6CfG/TVr1W5eh
Gl5wMmF0/cLGf5IyeTaf+BZTOwxZRUE6Ys0ajmp4/ZdOdEJzJqxKonE7sJGUVYxgdK0hEDNDzuD1
vZ9dV+2J466QKgayZPR52kBpL/OR8Q9hipgYeqZIjtDwe9BcU9VYb0vTvKldltHS6f5I2oI/aW2f
XHKGUKvoAJDpMHU8jCd5Uc/L0Ib50K2O2N04AykcWPzz7J0WYKZebTPuLdiHJyZ0PdKkU4aLB5Lb
11JqeSzVtx1vAEPTi/yGXphTrkEjDky3OTWVKmgIgcjzwkGgl/gwiMJyKEAq4LpiPNgDsoPeVIh3
4bhbTpwmhM0TvHuKj+rdngAIcB7/iWmTdI3znsMFoIj2c94G+zcPYtWcY+ne7VX0R44AbI5iUVwW
yX9+9kqc0OmLwmKcVIsN7ZH4f/uHiTLTPUOhhPjy7GfYBP4CasFEdsxnlUzyXy5N0cRhHkrABI+s
Aro5Kj4rwEnfRNxctwAKfg6izWJUt7XRSaPnWsueXFhZhwZ/VN8KKYA2iUraiXCNS7rmjwVtDfIZ
kmJhPZMmaLw8w/P5JpVvDxjogbGClJgBS2qSXPZsjg3GURPoFb+Va8jex7mCydu+LUxsipnVj5Y4
7UwuhyLXY6MztUBH4h2AltcUO/YbrNaDiwiDw6eJHlVPyKtyEMkMdnH4pptnVY0kBXygrLFcRRNz
R0x+dKd1/3rL+oGH1afnkK6R9y5/0CbzsLwKGDhlIji2H9Wf1z10/nqEsgUmvTZP+9RoZ5TOuwzf
eYsZYoIdiXAsfcIfgJOziv6nzvXgePBGir4j79BRvTQ9o+abjvEqtrnxRkZJlnHc2Wcnjv5nmWCk
kDKgeGi7epE747QkJcuJrFpiqURmxEfBg+B583FJ51EcFEcLSv8CQXn2pknDsCXeinssa7cRD29o
KfzvClWZH423I2+VFcLlRm+iDJKQx8oa+iFjda5Vk8puVHyJ/oZKt0XZ8z1jRAs3IovsHDxuOMaS
99niXmcexS2Ro1XXURzKVJzxJY6RhgXb2JUw6wG8qIB/70QlLHWwUlB4uuNeyfLFlcMCNoCEmXLa
z3uR0CvkoRsGiOAdBZWUfiMKe4XEpMy+nYC2r3bHaeUvpQ442f0cN8PejCw1c++AiGZGF0aUpFo3
QkGqGZKxwW7tO3ODUIUTKTz9HVO3qMIOIQPiT/f0+a94rYqLrRyYvXQskkRX/9NOshRfqFy5XoVz
2v9S4mSNHtmN3NGwh+nz0yipl5IcdYAixfF81WbjfJ2DTYBMcGigyjUS10YvPhTxCVFt+1tQYvOu
Q5JYBYqEPbYA9SOq/ZIMh1kALMWlhhkoR3G+srpRAR8Sq3DcMSI3QK+FbDsOPtiMa3KJoE8FVn66
aeQia3DLIwJLXwJPJsjCCESjNsR7mANH1ngi6X3Cwi3aYoENxfR4z590WirQcgyfQz2AsyQb5Dnp
h+ejL1jMabBIRSGNOeWz0h/86hVE99HAtboZZizVsc9DOKl135y3a7DH10DbDru8Cdpwo4gQK9e1
LOGcubK5qhgUZ1LvuNK3NjD2MhfiYoJvkuxX4KuZpX3BiClSrraR6u2p3naW7j6VAq0FzlJX9JmJ
aSG/S1+MPBO5/MHUJniUhBKP/VvwRsKD0yF2K+dPYaM5dEM39B4xi73vjxxkBJp3KAN1xtrOH6mb
mBlnZM3uSp/E6aSkm4nqYEFQTwwOuZFOHhvm3X5ovpQ566rbWbMen1S23yreYbLLSbbohHd5R4hj
Bw4nNo1Ry5G9i3XaleY9sZxU2k5tnC9tgqEMFvHgY8v7+S5heO9B1CaAmlYpQNHtnmJZ0VoF1a2+
YaBOIQP4Ck6XfEFpaRIq+gt2NOBuFOjNK3+rpZCo46OEIfJsXR82uu5ZKuJLOYgD2tql9a9ekuMH
xk1QUab1ALmZVaie8A7YusX+OemKgFTQoQKN181dXRvopOY49Y7AKCHNGSORWzYNFO3DVxg6uR8W
SCk/6eoRAGGbV2y1ePgGdobofGpD4qNJezzXmR+/gYyDB8CwckAscaUA3HXvFQ3hCATLz10PbuIH
wGUmA+hca3AfzepYQc/FHiY01KhaOo7uxu/n9tHZg6MpJlb+Io2HolgN/B+C7/L4FH1l1WAPMh6F
YJf/Y5Z84KdAJbBN113epnrlIACzHWiA9XfEVkBaUPo+tEL7KV6M4VWyanPHapesGJdbBqkDUmDL
GO/sBGE2W83QUjMMO+6ZPz3Gug2EPWJuV+1DP69oQpVExRsFhvRIlUFSoHVpT1D+3OGvmEe4XAnJ
0GqEDGEQkLlzClF7qWUGZDo/FYxn+1ZtLWnFYgNFyEQf2pGj9LDM5GqGaA21OmAAIETcHaU2fU3f
xbgXUtQmwWBt5rTuQkfB+sdH3OvJCEKleGL76Vz4U5OX4bCP5CYm9bmB1rhrAbiMuUYZ3kC8t4V0
fzqIo0tdrmcP+OQRtvHCkaJr3K2VnCQCoYAATxdO/3wc2FdwmBggRge/HR+y2H263txqXJ+abat2
Yy7Nqzm7k4Le1Bq4dNtMkzYFJ9GhIDwh697vNcVUbTNR3tpKELSivuB6FW45YYEa4i3g/gpDLGV1
ii3DuJzwm/fDJ6WV0zpP9M1fTWQP9fsebGgtGeBMq2MCzmcIXSoAZ9KgqOYSIIUwghVjq5kxdT3H
1S6BOx0FRMZBh/v3NMo/su2rGH3zDQrqrCzuNCZYNgnNVefO21zLSlSVv0wrnstexTWiw3tvp35V
SvHqI3086AgkbVHCO1iXhruLIZd+6je5VhrX3F7/lQX/IaN2mPYst6udynYWkfCk5jY5zh9BKTi4
+UxaUC4/oyN28mjmmkZaftT1t+oqCTTgGZl7ZyZbNOnTkRqu20/Svb5G73ZbSqhS+hPBdXi+xXz8
Gf78UgyyGLz8XU3ER+gI36EIIHdjVb8lAqo7tIBFm14rjcfeZAKven5oZD5zV2FUXkYA5q4cAwyI
fpE5YUtpxMECujJOtr0kOlArfciNgC8R2FjT3AA8PIO1Vb21Pc9Cp3eIYVtfIvB0nL5ZfCiJzdIr
UXPsqKa3Zfj1JPtQxU0bQ2N7ZkvxaaNwQTi26cZy0yX71eUCt5E3iGCWFbfmSed43GX8V0iNFQ91
g5sx3a0hMYPnXdy1a31pJEJ5Y5J/tXkp9aiG3jJC7QO51jS4CGWppVmWzPhmZa1x+ZAHRjWS/bbs
jOMXP37Ta6W/1bUcWv4crmlpFA8PHZ7u/4x9Fk4MXeYXJAFBytWOME4Rnhmi45yptGhaT/BJ6Q/U
a/4m7PZyJNrQi0rqrTZmqsJjgBsNfZ/I4X+jqAGpRHZe1sh7Htf8UitMqbvNS/vAwP8KDSN5E8FT
W09J+vmh0L3XpdzwBswYsI9NA5WKCmHVPEM4nQtB3npWsErM7zfdaI2c+gZL+755dHpWbUCz6xRG
2uiJYvvBis3j1XOZK6WiIsRBDfrHIRJR9ObMblhe+MksvXxBFZMShA4F/3oDNu0YSXVrmLt2qyeR
a6yyAo+O+VQIhJ5CSv+Q/n96fZzduloAKFHsJDab/zOqBz8ZI5I6XdtbfjsqZF5KFfA95c1WPnVe
Esi1mpwJeBTQ79waqxeP52ZiswIlcQ4Yb1ltmpK+uK0Giuxt7Rrp9Mvm57JugmSizdeWrVlcumix
2TaSK11LfXFXE65F6uIF9LznizQDgn1aSlkTEUB65nFxRbqx4gslHXcf00aF+aUuEEpTa8KIOS4a
KfeDTYrAzVJdyaNvcpnx4zXVILU0GHEn06nTLCACR2om6067hPLYFx9j0zMPATsBeMHt18WIlA4E
yUawkMiXdSm4QXk00iJEFQBPk1zKWDEbbHeW/EmgukzK+B4+6Ac+mnMUv0mRXImS0GvCz4QD99ty
kl4OWjRluZx1Th9cRDYtyVJc4GyDUfJzCYdze54tOtWGpo3SqsELvVIRo/29rbBzxW6Mypj3v7kj
RvohC38m3QJhxHY5SNEwcqs/JWL3TdVvYnQjwcLOaIYe5E3m2uWNuuWb3D2XoizjXRxR3Gyp6JV3
kLCLhih1pFPISPNwz6l0RvMxS2NUGHn3drP5YFXg/ZLAb2H4DDIhT0NNFiwTTmUgEPq4bRx/uRs9
+ZUJVrR/IWNu0XcmFggxXYQw8g+c8pzGg67nT14F2EeLhCoQpB901MXxhAxI//nzrbokthfwJp6/
qox7w70ymADK1I8SJAyQPUpz08lFWc3fsjm1HekSJZWOZUmLYNTy6qGP02YTud8lhB5daFfC77Ez
GsxCL17vYTlkO7dfv1VUyoku5VL9181+3ph7T9eKAHBJwUBCbhSGrIpQtYydAJF6uhqWYDwUJLcu
JP8dF3UNKJEI68vZC19SJnvbV2TepnZ+jQ14TWiA7WNaIdjddWo6
`protect end_protected

