

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
O2XOryoxWHSJpVHdyGBaJQNdc8dOymHDuiuAfQsjyy00yg+Fygx/oSQcLoNz20CMTJ0oXsfO0N0b
OcuaV/bA7w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GVuiQASL5MnoVfjBYAuifaKQBYP5qpKi94ZTFg3hPhVSV5Z3K+xBNk7HSc26fljddtOPeyiQrh28
UfOI+r/9r3w7ch+EIVITv736T0H00tqEtDgqpJcf40ZaJFg7/DAJqa4bfrwQYMPPMtN/+LWpquNE
dRSjfIReTFFkjcqBuxk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kP3f3BnKcYzaKjuqBtrZmy5+UEIJ4O5AkfCZWz9sAHrlVU+4nM1IBXUAwmiC3k5d0krwcI3sEm4r
vt+G6kIqnFjoTn4NiQbiqvWYDmZzV+LJflhoMqNrJkRkcVVp61x4JZUlEr7e9p00rvVMbcTDW6Kw
nnCwqMLBkzM5UVDhuEC2tdG2CpSgECEGlLMMTk0DSKezGNtQXz+KtY6h+PnOfx+PFZwhFOBl/jB2
jTMtcKAeD4gg4WKoAn+7IIlgw2/HhJB3KvzLJpLw91PETbk4sabjQbQ8KStQpjvFK782EG+wfv9+
81MDogRQiFyFmN6oxg8ELCZnY8O9CQoxYornjA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
u1fw90y9ARra+4xSQeglVz70mgNc2urrAekaZxIT13N7fl3y5c7IkQ5+gaCLFemZ6U1NIJElw95Y
NB/VTj4qfRZU4t2hFTedbkAP9HTfBoQLkd5eok5logHyANc3ZiAYnVdPL08Ys63j5F1wjpsesyup
0l3zS8O13B+I+gzKcFc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tgz+QXmbbEHiuFJzeRhVhbQJi9JNitJrdU91eD4OUl255UhEJMjfDaR/UN2Kmj3daj1Y6N9XoIi4
93BpVsNATisoDDeAvL/Rji5I3h7VXyiH5+MTk/s7Sj/KtzXNgKZlWFjJ3fcXqt8NLD6Juh3fnX54
GPDGKSPlW9MCzzT1JtDTr124bXptK/drTliCAmE7pdznkO5CQgRoDuEMokxTyMyOhM68hW0orIve
hBJnTlVs0V8aXizs6E2X9cL1ipD/zg1cmKwssQsXb4Jo38wsiBwFRI72/29AenPb8DiuBit8capG
ogUYTJYZPuHqoOjMDVs+8SZ9yLvbdyM/mPqYbQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W9wfRxLjHUbwfTCjVdZcUlkVYIcSGOY5nHZELBaw1c/NDgsx5AflnXGqVw4ZcJVPhssJ8DFS/Hc0
BI96JG0oHrBsT0vEMRXoqAsIx9uiqFlhRbqlIF+e7F7IeBTdC6YXEXctyyXaAZNLmebzM3iZjvNh
ALtVke4lfkxz04zLYQv0C6ISqIwI+PlZWuqgIkOTgdWEtdxW+zW57JrC//OTuGggYGgTTtrpZN+D
56aBhSpOLY6ft3tCy/T96Rbxc23Ol2kCLBG7e8/nHNSSDpF2k+L4dRyTkMYFBNGDcszGyu7cghxU
TRsP90Nwu4h9+YZrBGgV81oXDRYKcIAKdTl2zQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69472)
`protect data_block
oJeKqDGNiBYjPNbC+BXEnyA7dDqbGH3X7DLuEWp/PoCB2/ghzWasrHqh9z3Elp3dUbxHL9J/BbsR
ks/qCJV7dUOKuwVeWt8OBbNoEFs9uuoDpwKSYyRYK81xl3NwBe8g7SVIVN0t5a0Fo+j4D9oKlZYd
mIdxQ1a96Z55aK7W45Y5wNVv9odKf3ml5ECoubtd0RrrU3hVGP5iKVgndmyZknkvfyt4WwgZTOr4
9/7OvmcJrP06VV+/spLgStiEgneIuIEb+NPX1ib5h35cgrdnNVCmUVirbzo9M7AWWYVCfYhZ8i+/
datcV33goeZnGN4vJZFMJLrOzg5bEngYhFt0jCTiMHKDQqxmJYKsAOYAxF/YAVRJfXQqmJ0eCYLp
+zYobAtUa1JylUztMeJQoBC8qQ0/YXgtoP05tKUHc981FK9f04kZSyVISpmJqVhZ0hbB28GMDPfU
/cY/GQNlFngfGHCMj9LbQQ3dv91f0XPnyzgrf4DV+78gzpLyrfEVJQ2C8Hyv0Y3/C6X4vjCV+qNu
Pz2yMnjw3SZsLgEHjl+5NKtHB2NiurFyWQ++Nsq5l5k7ifLfHIK0t/gwYz+CgSTn8CoHsKe/vXgc
Hn93ALbVEokYf4cd+V5xkhOKgBjhhyq7yOBJlZH99TXT+Ma/aIUJBFMC1bFfYAYfUZ9qSVBk5ru3
qNxiYK9Yp3RppDOoCMY2pYOWFE5ApALOdbfJvHYmt/5BG1o2OwXdp55Zxnf1yesqxf/MrikCL58y
/IxajH43Fo1kC4rqwXDPdxzR6y5Lph1A4vwAwu5D0ebdE4EbObtYs0s60LcIP+ldj9KxAXpqynOF
FT/qOK3eJH2bxMkazvQ5iI69eTtlFZ9XMnqTWEZ1aa4q7b92soL+eNYKMoEDreejVaYt6fcFXNk6
vGIt0V8ppsyuz/9nFADK4D8UA2h/QGh3bkp43OG097g32eaxDMdTDUatPhuU/8/6P8HsxSY7kwXW
F9Gy/vVOtktWzqC4pyoKymu2nT7uRd8mqvh3YaAbEDBbokQfMJbTJRFS74w7b31KFI//zVdFQ8fJ
bvFGQLc7aCd7QKasdBsc1qTmpfK+yBliaWgvueYdqZbelJ4UtnhQj8/wG77Mg2fVmbMbcxVT8hSH
TNl5JfCvcGoSZlE4a+uMpidc1TRYpZM971QX3cHjihKtDhsTpWNzu5aRJTtaZs+3kSzF0eCNM4PZ
1j/+J5tMdQq5MC/FvUZNNCSGHS4KTNNhANAlu5X7c19eS4FgiPKMpC72UodhIeQXsUFljertKGvc
cgQTgsA1koGBit7alAkso3ZdXGXKqrIhjFgSSWcv/37p5RKcc2TocqlY9oLp0sl0aJVm0KRDAURz
iSuV6tk8k9WNQyph1ZX/csEB/6FAOTDQE5xQ3Uo0iOzw9/mp9+KI5Hdsj53r/QZXUZ3W1PXFnVZA
Dq3AhSO6xXA1Joxlt/pOTzy3zexmDTa6pRkrVHLmIi1bnl+MKbCb4d4+lT6awp9pRI1AqjL5pcRw
PWBCKWNXM1EuIzzQuj2pPnXlir5s86Kom4U2rDT5QLB/Km/lvyW4FaQPMZbgc2F07iR1eU37jKw7
fGmfxC1T9o54i8lqRzs0+QaWaeWygwEjv50W7n5v5JQ/xF+Q3MoaW6Bl9EvDyNUTf59p0VQ9ELHg
gP7La0J5QPQU/WqVVLnIq43PXlgfxe5iHGoOJG0C2vA7mWcH7VYX8b8/7+194cJXXM8fuX2Cu9RL
kNgaU2lh4E5av+DWcE2G67Q/PSWPfMQfikVajkzWcp/QqKymdCoQ2IroLLq7R6ajlAeX8EZ5JJ4M
JgBkdrBbAMJDXJdDCvIWklAb1WD+MZsMkPj5fBdXwmXSRGYTsNFYd3wCjhwg0dzEZQlhHlD3DmfN
fThnDhWfuHDgGpbvAlHYOWT+IPX0qBlk/ABvQwZ3TaM0DYy4WqcApvXwY3cfUuamH9BaNMTv/D6k
hmpp6lt6Nv7nx/q/nCfcOUFxX5qgpRICVWrEy/OQt4AJjZDITZ2sHrMQ6PsMeANlOeaZj7rEbnSb
w+f57ixB9AHmePtJgvjvffysparY42u+Pkk7Dw1nf5nG9Qyeox+XRkF7hyu510MyfipbVTXc1/P7
mLPXngIisgx9LTRJRhbEezT4N+z6bstC1GyTWxTMVjTRW2Ae3285oRV2QEjlFEyfAWPi6qy2B5ji
+JmbisueWY2YKfn1htwCDrDbdDq8Zuk1wUysjG9KC3ConjuGYcvrer2NpY+Jr7ssKdJV4vxUx3OX
Q0L8xqbgMtP/i//TaDBjWD/l2O0JunZerfd1qFrygAWsLaV/Oy4Zf3NCOChZly44ahnTlQapOWzK
kFvBbMxxyJokOFYGNxnPlBlYbIC0VVkPUFKBOyppqiGkliHbe/PFCi6Z73JpT9OwaO/txFoRufs/
/nG0zp7NA1euQ4bA1+gPycpCoH4VbWLidOm2qe/lTrdoU2/Jyx5G857c2bxJR14WTH8/NJ9dDnPz
5C7KVIffzUI59eP8Aq84GSQ1Xg5hfKZHU3MqRvGPopDeHohXoFOaFrF4jc6P0BFzodA+wO7diKOd
iIzhikPZsMkRWFQ2r4jh1BJAhlTFQc5YZKvzW5dsFifIgJvf0PIy4rsr7kGqiOqKv7Qj7usPWmJP
G7p7eBIAAqwOI1t1U+Ix1BpJIoXYuSG5ylVo7LucRpUF1bFqkhpoaTyQ9imafyB5wvg1Ogunp9Lj
8pZuS7Zqrg3fOlTNG5jlrtc/aXJPP6tvOOVklLoMWkmT6ljxiWQT8FML8FiLygD0LANz+dHt0qbc
jpueYq/CHH8U/hcXj+MNUj7U05Y0iMwX/+kjAhncpVW6RVXvmn+aUKURzIYB5HrvSYcWiElE7ef3
1v0atnxLMPw40e52WllBVBv14bvMu68c2w4qBCwtrCTb9biDijf40OJ+Uu4VgWzr3TNSdVHCRMn6
PtdFFZEXQXZV+aS07AWo5+bOpT4roNoIxNNgP7EQHQiycqvdV+Pxq237DtBOsrb3Lq5VWkd67djA
nzupahS+a/r2Et14k3xXJFc91bC1r67oMUoS4GLbr7g+ltyNuy2fudzHQroqZ9vzZulUw/oOb3ib
c+0dAlSVb3+ZfgAOAPIjxCi3C0hkgPU4bkgeOpOitFYDfVuYVZaIRsPGOKGUMRJmcvzmjabzA2NH
9Wc09VHniQQAFpQ9lKkVUbWdzNuNyyKzLTvBnLiZZmb2nqwrx2UwAoaY1P253xl7rUpMfFe1FiEf
2/aFRqhbIY5XYp7dwYrM5gJPzoeLVraw9lAMWvhZytTRQBpfJu3x4WpCYcdQuMi5VRdMZCMgQ99M
RTqtcNBOX7uERHRiLaq/1U7nxJ6Ya6CfeUyE7h5fnDv+xqK9OoXf9+5gkAIb8AiFkT8LA95zLBlo
g271Yb2flhZWneoJKI47P7Nd9ACMSUYxKTiNeHG8TRxpMqmW+UT3zdc5uhJ29PWYlN8g6yQLK2yK
ICTlcq5qKBKIuNe2jc/cQzIaZ9UTCW/3MqDlwANTQkJpY+lYmFqqMAIk8huaqv0MxnVKaNs0Od2e
dx4ci79C0rNvvCyXyiBgsqnAy+mcXX6nTcvYB2hssRLgCFWhhKJR2MQdfLg0EKn3Hir9WhNNEoGe
bEyZPQlyKo+eogl90mWVHIYpeFDNkJUnbaqVhhxoKDC40kpy8Ib/dsSjsou9UzdvMAgbRWqLYnJ7
y+hzGGog2lAqgxJpn2qvLhYQh5n6N6IwnYLco/ZzczVIz18wRxXz/ORT2SZyCznJXHBQZZmRXEUi
4GRgdIhASsYxROlVSSSPwDDvvUHq1XCBY+jRN89+g81qXnQLmqsNpGiiJYX8nJDei2XvfIHXcT7A
8HJninb2GrI8M/QPHPa4uri9ogqRw6BviywFb2zYz47V5YhhqSLD/yFX8DOD4Ui5HyhbEqtxRQc0
UhBUOC7elL3gyoMSyTH6pK3Rl3IhniE9DQh4IfKexjrDsTkHj2Y+a1IzId7+tdJEZlk+WC1X6Ewx
QUZzjcrG0oh1c533+msayq9pqsrehchw6hSSRhzu6AbZQEObcyhi604k7Re8yASe3JhwL29MfBhf
T3FYNvftVjKNKbzLxh2/Fn/qGg3QdQAo0Hs544wiegUJFk5FppBFXacJN40nOpxOduXVHccAhMf/
cZOp82uU+MKjfZf/hLv2IBl98qU6eDFs81rzNlR0J7f+pJR5ypPF5zzn6jDPVdi33DSNElzVghEU
LAG4h6Mf0d1IriFF/BVUs4oMurNhWMMXTAVy8hc5LyTkrGr2rWsmvFDY2s/eDaC7Aa7d9IctlS/u
NdOey+sPpRMpeY+Rd2U9nJsmXCtjEdMVzN6jdGBJLFVZg5owDoiLe+JTmCF3pqeAviFjrrwotZLg
kIC3Yf+81ueOKJ6EGnRVTVRJyYAze+xaH9lmajAwV7OF+P3moKw9zQ4Wz/6rLTdSQnWnyK+XxCQb
EqTKJjU7EGc7JVdSc0174FLdKp2L17u5ddh/8rU0qTO6WdZqQcWtaKo4edQe0J9ZlIRq6CeEOCzN
ukU432HDOKhUrMtGQDSrRHO/Gxhp9UNc29rpN4lO7q6ThPv8ifr5HJ1vA3fryXuGKZ6ZJqeYwNmx
dVot6TGhKuGly58UZYJk0TEmwzBiqpN+J8IIbkzvmzL9v2Ybo9OuETOGJHTQqR6nNc0hU6l1zx/z
Na4ArbFq3eQbwHTPCK57+cdABNz38nlSNwXPdbZggap4iDMyKVbEhPA/OMsWk8g5w62FYk6uLU3z
AEEEU6YUx0JsnSHyDsgoU10NMoErJDKPMIsKvJ2QB3dMuIdtxDLt++iS+ozLkU4LUJARAek86L++
lOCJN9TvwRvJ81aBsLTqUeGDDp+lWss6i127Wrh+2JJShyDoH+jCY0BfIW8dCE/QJGLQ6oVWeYqH
JB0yRSOue6XAkdC/IPM4Ha+uG7JscrCTgqmgFtNobaCcvYXInYp2trm6eWM5CjsIJuekMtV+n6mk
gpC4Eq7Xq/FZBLggKOhfF8dCZcJ7dHWKAeOb9pvCqUmaNhnWUcbI8mTDEV1LEB0bgNLm6xLd/Tld
h7MIYxi9rp3xXs7FXoj/3TxtPzHhjOM37JG+pmg2bwZk72ZYYnSxAPY3C/WoFP2Nl8BXOfL45Nk4
cU3cW4jYfQQbZPgYJYCgQJ3PEKJG/nx5kdGYY/4NUk1fVc7Tw/CcKqHj1sliFEdkttSGc+VBCcFf
P28iMqpyVYU3ytNmsEIQzAklpYN4n1rqM2qPx3iq5nYk9kjJRUocIWoQUVjuWvo7uMSCzlUf1GSz
u+F47SbNOa5WLdwdk0m0UIV7+sAMnhMJG5EornmVnh+JVmfBzsIKk5zbYBDQmTCgymVAD90QTbkQ
6UkalJeiCIKYf+CmLTxOrCDXDLuU6zoN2pcIcxmUahGOtft5NMzcT51V30BLcw2PNWGxhrBpDtaZ
L852hksTXcYp0LUTlVF8W/ANgj/k4/3lBRZxWnrg8UI8xsg0TuTwR6Si3JurgFFgkFu9Zh663a5t
Afw+Knx0Cexo3Xqxflk3n2uE7NgCxz1rSWoYar79p4MnkH4vXcrZPbUsc0PhiEBKRf03wtCOtDJb
u3rVb/sBFSgZI2iBQnFFL4dGin0mfleoHzlopgQiTXrlgQ8MxasOmLe/S3A2ghkQROoiky/EV4ds
4y9prnXdiInPoqblpKtO/eTs69QdqofFp9iqajJX5KETTDcq+g7+wR0vCjpgS0La1JVHpNjpbMt8
u3u9hlrJ2Sw7XB3Nos5chTZiAtxVgsKeHJgzUHZUIXqVy5GrRKCm8tSDN4w0jVl52tKOem+VuQVL
6UQqv9gukNLM75RSzwkeVSD68hBBPlON4O8aK9JE1vk4tHwKPBvdWp0sei2K1VBMHzeju3l3qA2+
f4KLZ2KgazH41m9nz2p4HuMfJAdjY3BEp6vCs5/n0DCZ75eBnoTmIKoW0LSu6S8wof0mWmnPIxdj
ErYe87n44SA9wb3Gv7gMLxxEHZxH34SL310lpnjYqDe8jIFINzHEL5mLcvlx7+mU5v2a/8KnHovL
7PkxH45/fRfL6iWJGJOOZKBvSCYVmERF9WvaV0dHoV6yK8rlIu640s6zBokJ0INQBp/1hnHtr8hL
GewxNLK8xCN3vzN6iroaFapduhfgqJ+gIlJdC541zuzmnM5Y+E5AxppBOUn03JaQyZnLibetOjFf
W7WbwoN5cEd/S+RVFIolWDQSJ67NqEJVGwzdnAZYcHrzvOOafuJWmzPwFcrqILh/tbLOLu2zehBr
qeWD/YTuCNGgvFzxBTHa/kxWcodUNBC/BZNq1KnssfJX7c9hHxMr+EdxanaiF8h5Fwb5kMNO0GVs
Ktw+PAnvCP6caSDNH2nqbgpB2j+1ViyE+B33sGzmgmm2v8kNrRhBEEvlvEBbM+qVsI9XyJyENPBy
lssovHxVa+SXblIRRq5yyo6eGkKzH+olBrOd3X0hS6W8aRZC/ZYi5J5KRHgeSykNZdhi1h/uNHxH
7GQl+vS7LARLop36rKX//Gmmz299wZYQRJRy0528jGV99KRT5ON0HdNtcNW15SBdoemeGmxkIcHf
j7opgjr2QlYscrZbLA+T1dLmYNwra+MoMID2vWv2cMSsCyBtafB3mK5tpzGfy04l1LbYieqmZ0dR
X5kjTMPzszidiPT4ufcE0snbBdr9kBERcwxnDS8LTOfjIV064ffwZt3fv3sqLgzlVksphNEDTMXd
pOrUuD6bYY/dZBesQZsNlxFEWD6xV9HEJ2AmNygrvkSpKLoi3fXtpvLOrHyRJyIlrqu6+9XVBj4V
meQUn63osrvguLsXIfHX93w3qEv788/8nZYUvmEMs2No2TGzPapXxlGUeWf6OFNsBideKNQc7l35
KFfI4cFVacZjUK5nbC9yTI3KyZSKGcCr5drG164U72BjzQNwEnXEHwLi6mWjvlapE1/SqnEvA8Br
mF7K2vOgM6p+F5TghlDl9GQDzOjb33lLg/EUI/TztNtHbD1xq4VMllotlRhIBBiwTADGnjO+d2Uu
IDkxj06eWRG9LgXJxKsZqod0bQ73DFDNrBgFLDHlxy35frjoUT8amh8hvNgcNULQho5VPcGRKsJ/
oMBjuftjtF3c8MchcdhT8WHXb+sWq9GWcuv4pWxS6mywq3Kpmu+tFUZe1FflfbIC9Ml+lJVk0Ocj
JOx2a8x7SQzsXsMCj3nas6hTgmgJyRPeIGDZkEidg5lwfz+NxhurwF5a9dlU6UxnzjkrTdvo3/tH
rBT0kWuw1gI6jMJCOt6jC8FL2h+O9rcY9a10wTiC2S3kTFEHC3+lR+Gg1At7EUJgqjHw9HFWPVdP
9hB4ZkQFTDX3EehldbzGr+gpzOmpW/gIsbwCRUK840fXLG76n07A8Q/TTh4uqoB9u3Yl8PuUUNmu
Y4t++9+ZdD0KfT3d9zF7wTX94mBOIT5TaSl/oGbp+9V0y6Y4A0xFtrQceS/TUDLNW2okRjxZ7Wcc
v1H9BFq4QxB2cS8N8vGKzwIJd+iO4f2xlSW0m+cJJ1Fq6oyVYdOj+eJmvxc7cx2vbZf1Sx+byyVu
QOr3USUvCCODI3w0Utgi+35X+P/dtb5TudXjOtWqIrAiD4HNZpnVziK7pVZVX0vBJR3Gc/vRyccu
39bI3F+mYcPKGCkTZI3Z8wCoCuRY/5e7kb07PbAnOP5gz0D8WUirpQtuVs99gjKr0cxtvocjko7O
jxp5QGvcUjj930+RpxXUFM/xIjBxZ4BY8y/XjX6UCTunzswJYMPT20u/ow715QHUf5hIU0z+eeMC
il7js+XR/bbEbj1mgTlWbcz0UZ/qI127dfhSgC77h8Nrrb8W7Di7t/4kYm3WZdUg+9wwq/XlE37b
unzBHaMpre1PKdh5qf/qK2rUt8UWzcrJgXkX9mYzXhBU/o9qdX7JG/2ilJsDVsjrkHr5OYjHnnJu
5SvBj72oYYzmAFksR2akA/TfXo9gSN/BPtbTgTkeuG+BF0+FzOzcLe30j5n1aFnGrDWtlYlbq5yw
LzHPY8jF3wgN7UGziAgxMD10KGnw1TK7p72du4SMPAoUqwCkdURQInSxXK/HWLoulKhlNOiQChsI
5u6+8QISetwdPt7mhHe4mxE5hdsJBMg06gbxRpfHKbZyG6mOOifKExKU78TTpT35My9Hvwi+x/ad
h4m9CYq2wfp24T+nzsHvc8E8c8DeSRjefntZ7/FTDXLo5AeKnBc3P83d9Gh6x/9loMhKl5fzaEUY
erZMmgUkpmNFkspPsnSlk9dIrCW0pL9KTaUNDwqWN79Wr0LXyjzuVc+kfCTy7rZZBhDZsO0KDnGM
NoFrkGM1CYySH3SAxUgo0+8r04Z1YtKObYH8B5kuHWfkDroYP7/osqXNy0l1R5UFGIkJ+NYd9/EA
GcLZ/4/xMLF3/QazX9pnVy5WlszyM1M4PLD+vdnRZvqNGgCntTL9YdA7Xu4aNhWA1UsOfVqiRGxj
W7xXxHYGmTrlGxxIu0SIe8X55sPCe0lyiFZBf3Uin1lOL3XBYA2ohDHkRMW24NFDQV3KM4bGy+yq
iDcGlU6eT+ZCEU68T2LIgR0OlccH7je37gIXTHkyV9Hc383f33NLCOt37DtwpRP3gOgchq1xs4dJ
8NH9QRGZZNw8BM36/noaAty9b30/OH6Zt/AURrSuadUX9H4qqP5VfkQtpG4U8JIBKZHjhzluQ9nn
dR9JYRM0dh3pd9/+DDBkMPC+C//f9G0PDRkWVnDL83n2//xkx1xXN/C3GvPfjQoZCbzV4hKVx7uS
sdy8RZpy+PiO/vE0t8T58XWHtY7x7COMo+G2pTA2jMUkXOXldaOT97V9/P1TrE0jeg3zCKqFLQky
WCVKaSzMP9QWKyP/1xaXTKrczm0BdYYooeDQDQiCaZpN25yq2f+VwRTkMsjq73idRghltvf7GIIO
pDmX8S70pFTZpftmnN3m1OFtS6kLyW9kjoU8IIqerf8SWdmJirKxrkZzxcVeFD9C2wSoESsuYPab
PSpa7vWNr2exCKs9VXykN4Nw0WMb0K2OggvapmKCamHkWGhbIOVH3q1VXb7mnZG3W0+344QcgSAm
bNdxp/63LjAZqNN3Wlu8sbbuc/Z0/25k+cHp+/LaGjmPpUWWC3Mr0HeL1n1BBlu16MfcdT6VIQOG
48gLiJWMj+k2aw30+hKBWRFVrqRg80cvZ/Ei7Cd/FUIXxTWd3V+r+CzTi7nJRZV2EaUvfUYEuVv8
qjCtcYIxD4+CwiNs48WSxikXE/uGuAjsUGFVkTGwXg4Rj0huTrROo/rdWJF2tNxAv9j0ewXx1VA7
pkXRYAkqZrxlDwgb/N9GLU00nvPe4XXwaCp5OlVN/q96ItijxlGl0AC/CEK3JPTLcqktbe+rjdEm
W859aumU8Has0PhOM5EiC0KikdT1Cn0AWuth+hr1eLJXExiiM7Eo1rdsmYaXcbiO1mkxAvaCok0Y
ZiBRyyskJUFh1GmGx8Mq4y2l4LmBbqee+//NxsVbWkQtCe5AB6MV18uB+B+FeaqceApN2ALOF4Z7
A74DNqk+kjW8WTRiHr0w0KC7Igo+bQGOXTuxDDdVeI03ZM3l/AiBWtIRxq1DtJG4HlUCOfsqMzhl
av80n7aFBIEIFDnoA2ekWWXnwcvCd5+h5IqbQSWABx8ZJNAPu85/FIWuXTpXHkLmg9Mlq/+W2bxi
XnTBFs9qGc02ebwakKOhb4kOpUcp4YG5/1+LzKmZNijPtgeW06nliDrBKHlN+YJx7xndlassSPFP
HT0qhnqUnQBGEGPTa21AvzwZBbNTsXzJFSVSImm5LqkDykR+NI/ehMFL/Rshyquu+Nyi5evnwOsY
Zr8jtSgpMJvbM/rFBGI98hlCD3ADwOEE5pWvwe+sn3p6dqQMQutyOVHctA6KJ1Ku7Z4mKMi3jNL6
XWxSIkNj+F4Kuj6G2vxrurJtlhRgo9A/Ees64dTKIoAfmRtwcHbWXZg3ASPh1tqrz2ELp3NYWRrH
O2J2UET7YMdHMn3ds2KGavYPHvdHLujBVHKKGVLOYfmfJVyj4bVFFeQubEfJ1jHfRLvIjhScM8IN
TfHESALJOIeNc7qifFP3GtPb8S5ni2UvJK+1EpxLBzLWzHMaAMinPHnd5fp2T0q7n1hpYPo4aKmw
EfstmCVUdaU8Rw53gSXka9V1mznvu+eqXGHdtjjq7/TmTyuIwTJkD3dgCjDtiJTTGEAszGgol0j6
odgJ/N94p76q9/pizao+zxithni+fnsqVWbyW7U1/NHxtriHYvSZfOWBTzMD4GHOaRHiG2GL5ScY
CNKjXSBBqAfLonbHAfx+liYo3IzbuYtxpXOc4tZrS5aSK7mfzWCUvQ6S1LH+WpsIDr5S6FCvuvv+
DsHDWBqrs8uBjxn9H8IRgMTpc2zEiLewqsg4Qz7OgdlLAyd8GyXL4R5nXByEM8AnWxlFj6lCuV1m
F4FiNUbvNkPwb4Nu5QzBe/ITaICwnKByQx0U7OEr7Y6Jcz97cTmiom+K+5nmLdOGkN0vQTjFxawt
moDmhO6VlGFrEfHzHoUPTvP1cWtPH9sJbyZyFWYL7vYJsv9Hs02aop7FgNOe+jfx5FluJ9nuvMof
A5676ChdDs00AM0NUuAym5QdpGMu6KrRTnkqBo20p0oE6/HV9Fl/398+F/tdUNbHZk4wqAElbbZ0
5RHCfXQTzN+IAw4LxAeCo7S/Utrnhpdk/UIicY1lhYyd46S+9MfKoSJw6XTTGc1xVMK4Uu7mRute
Ntp1EFgZa95zFsNBQxykZMo/9w1XcHmpFK1vEAUJobPPjkJyUJnylyQ+pVVLnuaT/qiuDk+EBjLb
9BNzj65egsnr6GSN8iMuUEPkaGs82camvfPhqBbf7mcHclLd/RnGBmeNvvGYXRv1iqZLV6hmWXV7
jkIOrArgfrgATBt+16rF78iQbDAndD517kLIhZYQLL4VbLDCbPQW0PrFrLASFVufT5krInGRBtpU
P6mIG/oj/Ofw0G8jigbgOGUvK9qSe8Q7qhWODxR35VMlbpSfCDSSQAt4oHyJsD/Mr3iS1/OQxKgi
2awAEqww3+/QEnV4giP8b3hgMP3ZrqxUwolbYC5Hdx60OrbV0TJpVsY8yRrZf/mD9JlS0PrTa81D
oPejHUPVYT55/jpTNrTk9cp2dXfRUMnduik3YsPYnF89IJonY8XekuiohVSpgBKxRC3b9FdfZR75
hz/edp2QvpgMWzOUVEYkt7EsK63t6UO0inA4TUzYh2TI/oU+8O+X5WcxYQb/efICpZw/LQxGUhEC
ljA1q2O8tBefFVENWiWyfj3ZdfSD3JuCew4ZEbMVnhl5E10z5uvxnilYM3O6lQneYgAhrwsK+xTr
B7ZqLjNND1RRCeIIhd0j+hV3YdQsl+Pq44z5TbwASP7ZWCtphhrdKEDXh3G0q65KmzXXfiewUmhn
OGxzdhVOeWRqIYBQ3csrYRJOfC+H0+9jsgoELQ/IhiyT0KOux83mI+m5HxwU6Y6zLrUqFwE1KHt+
Q7u6ginYYzEio+uddj84TkvMz2OfuxcVtawAPnHaC/6D5U0zu/vyz7b9EAjQpG5JSwtN8v6VjXCb
nK4Yd+Xty5aAuf7wsGj5ZLhDfNt4NXanDLC7HT8PztYp5XYvYpBXq/0Tgda6FKbjJqdRJIglT/92
Z9a8WRfHxN4jZKex46n3Es2AeK6Hzjns03lCVXIgJh6RSSasawab3YlJ7t2qBG0ADm5pPoVSwdQN
Y3OTiuZGR7DsIlNa6ba/Wckmb6RZgRRxoMDblXVrSNbAVM6hPd2xeWVt3d/z7iGLLQynW+ENCqjJ
zW+OrNP2BFGWQ3XpcGPt8SBKzcvAaxc/7dZ25m5E+FBcDu4wu0/i368BXJb+/CZxZeSdm6zvSum0
80eVzWcLvvN3YSMhULybZHKC17XkleG/+2vNtVfg9MSwWd/TNlzJMw+CZtKFy4Z0Y4Qn11fd7PQ2
aTI/mZMjEuE1R0Y/DqEvnIq2sQh2An3/2YLdsplGQBMqawC9z/CMHtYyAlQz90GQaw5rXhS55aGq
j2iv6SgsfXo6skPC/eq3TdVaQGswFd85Li4bgkObm5o5PZMTwtQNIEo9cUkALo0TCsGcgL60Vev2
yCJkXvY8rp9G1EPq0Fx9cqfxwkJoFa/DDLUgdzEqsmfeHxWkCBhe4WvBZ0CO6Ac1cjesy8ciwumS
q5L7qZBP8OxgYq/q4BZ8ZPltnmh8k20Z/HdOGiIZUmyWigXYp1xLmRh1AhL957Zo+Lv9OsTxQSG/
7otJBMSMfcU1rMAkkLB7SbWGDRgMb6zj8yGub4yzoXzHjf/VJRkO7+FoAlLKNWeEge6jDIqCoFg7
xG4rTZ8gfs5kPIwxMBKdqcirtkkTiU0Csvm5kRtywuxf+sFV0xa4ocpvMQqEP0Sc9Kv2dxizRJVt
EEK+TJZQ1ndXZZe8t5einHg4hh0bfQM5sLZYoOk/fGD4t0UXb+s5IfhKLlMVrMfFMkT/vsmMeOk0
qfk+FZOUbRbALSeYvU9GoF3ZvTmNgAVNr/VFG6cHuLTGtS42jXZFX0it+KAGldi5KcF4MGtwhp9Y
qTfUiT+WK0VTjgABm6Ylkyeo5YByfKhXyL8A7MM8Gk9jDf5k+rl0JGQJOrIpzXySHeDCAAscpVGg
jMM7o8Nt++l2ftpvc9iSBDYHv/hvGIedJC6Toh5cSTgZk2keI4fYEMeZ8/bxF3pOYVMxLYg02HlP
vucqrQ93xDMMIEYtIb0IX5hZcBVPBPk4bWgKMviKz6Tvl574PghL85IPio3gR2ireUribYon087A
cEegsxNirM6MtOrFsE46t9741vlGQoijj4dT61Y647gOmpOo4+N2L8XW6dA31hrav18Sw3eLSyHq
I6Lt5hn4Dqm1aQyv+SsQpQbS7U26h4L+0PK49Sa6b+moTUzp0i5Sroy4GdXd+2+F2yvPImi3CRzr
yMyIUdYinVkdhC5fiOw0wB6brgBCtSIJfstqw1wVVwytdood9aNZgTuaYqAbNigNVB2ZGkrqpdOs
OQKVOPIh8r9CZzBJ/1Js0HjZpLpxCT9F//Yj2QVm3CPqXSVtwpDpsSO+ueG443qpC3vK78684FJe
swlecAQZ5YAPuI5eGTSkXuTVGtXWs8O5H7Jq4wSOJcKaAA6BzrYeBOD/8sPxsgYUYls4yIoW53CE
s0L1BSd3Rg1/kzlNNx8Vim0kTutYU77IzR9CuTCTb7a/ysFm/WE9wLkcr/kSCEMrPNgSh4/+zhvS
jRGOCK9HILC/tUgnzPK0tBebrjIWOGqgNROie/h1wALw9hxcIyeIBIHHtPYurO37TqV0OWhM1jw8
OwI8K4xBeyaIQp/M/ip3TzdvO/zUa5N4odKfHQ0LvCUrqZUKeakTUQxB4HvwGOrho9H6QHUboOw1
C+2sx5DpEbCh4vEFRZWVsfcrGnd5Fnmexl9U3vQIAdozwj81+hN6TkIPBnlYHkBBMsY5AxaEd4D3
nXOUTrtBi1Luhcm5PZuXVmwBfyPXUwh/o36+KZVQyuxp7CTPa9hq0Q+yEeiIFKuZpwYlaU+9fPFI
8/Afoyed49HC6EIwcamqmDXf8cWN7u+gQ7im4iDj5h1FoAokXXwq9nLs/1nkie9wnRFU/r/kVjOo
Rux1Y1gqR9HpI4wxr4T2bIKevp9d+5yrwseZzeH00cZvsmQOAg94Pzs8iUg9LeG3ngX5GJnLoln9
i72NYN5jT0JY85xBxoagg+CYs1iKbNw4eYE9ksSMmVd0043SFeerJbYb8/AhLc02BF6pbZa5QNZ7
pN2bmiyH8M77/QPrIi5E0JweT74bvd2yPhu2Bo5fEoDGuOtLjHlZZDGYva2bWUn9xLp4aiDbCUI3
rmy6SBehTkHv+vWOBRITHgTCimefZnLm5sLwKMYJ5zSin2EERdh6xHsv8dA/yoH69RLd2lvROMeT
WmOBGvnbxJm9PJV5NaaVrkJOZrZmtCvAVZmlclRXTLCMf8xqoWXoKlyLoCzgVJ4z05kUMe937wVX
Ll8IY9/P+lZocneEW6e4mNLwB2TP7fMKgwnMagMNBZ0kPMP4xU5R4m0UCJDXlkEUB8iCmbH7xkXn
8Z8Cy2dK08AiD7dlIIfXjuRfzJHFawyEsZGFLqIRQhs6TE7FLhWCLIlj1xnpNQZcHZZMoi5v2252
3UV6OP1JFcJlsDmQsW3GY75mZ7bwdLwJ8n9cdq2xafxPEIIzj4aAt3JBb2rb2M8417qwYaiYPQeV
w3KCx5t+NA/Lyzgy8UK/OO7fWnStm8mx465SUb5bpdowVMcYrYd6EgE0tNAtTRDP2LlZVoUIOOY/
Jx9PQNhfI8l+ISx+89AJoX+JgMQ76Y1U+v5nvh5ZjAx1Q3blKC8PWg+G7bU+BK/IHIZ6lRGKY07R
/RUN1A8xfy7aysr05QbAz5FEn2LsdXIooskVSCDsCti/X+2wrTvu3cmgfHWe9ne9pqOFQCu+IBfp
Dn/FFMEDBZRn9VFU6EuGjtXmSZUiLaLNo/thmtWC5UT4gdUFplYBlm9WhwVrk8ZmTMqqbTUarXoo
70LFnElGUMgvRSEysNc7qNuDxH9y2nvjA7hCPN0M91fAJETBWVVbTcJHjQfhyfPWzqVuCae9rs1X
eRbI+4CIiBi2urSCTJ62zMXZahXRkva3l8z34j9frL4KPw4+qv7TTgtO1DO55/chvO/4dfH98UZy
cKrcsbwZ2XVUOIbDIVAcFe2EXrhgOSO/UKgmQX5sJMlbWbCIj5gXcLKOVfklMg3gXQ6LlQE70yHX
s7p/dfrVjqtE6ucTYP3aeOFr3mVgeObQ1eATIX6p5lAeoJeS0B+vYxE+syAmSYa8uyM4iBBUjcGo
TxtqaeM97COz0s/4GiIcQaJRSlHNEFTaCc4Cb3MJzi8wYd6oWdO+uRkz590RVJvZ+J8H9ckCWaQ2
qYmGSKAnzzyJk28SDmeHQyF5C7fPVsxzmFiRUtwKNkkTRpDCkxPfy1xzlsoZSXFdElfz06qMye6T
Pw47rE2weBjJLRuykfAiJSxL23gi8+8CowgSBJYkBkWJ1WUw8C2pboGr9se0rBj2txWPoK/WNo8y
GxSKXZI39dPFfp6AxG3+lTcL4K10z/1bnL7G9vEKZ+y/Oow++eDXqKdFittiZ7Q5wNx0dTSmTyTs
q7//fJ6WIcepUanArX9PhgrKuvq8H3Mno0VLmEknmQuEQy1DDms4XFq3ZBd7+hf4JePUUe79XQ6j
yIfJoAuBIRrLFcvIrUNpyuskOwr50e4Y9e+WZE+pe8HUftZYGmXD7hy96bmn/qbinp0Urn/vbWxw
CeEn2BEOPN/V2MSbS1yrlV1GJiFNVlgbJFs8HCp4RWsEL4d0Y0iycdMIS546dI0PjDOsjGGfFKhN
Kyc2/6PmAAUUBtuhYLwo0/XEesIgMz7E2WjuV8EVtZOEyBygit8aIvm1zPVANaHkJVTXfI0R8bA2
Li52zH9pdSVkfA0jQ4QLmc0kXq1Njb2Dg1Rp4DbTS8kwUbir2a2ZpY8ll9bBqB83POBZ/1y2gpWK
NkcPlKOU3fXUQMcqaz60m7Ql0nX9tmgTsYMr4GGR+UttoGJTdCIuUV3bKPOcC4qNKzlushrwT37V
HZgwCX8L8ckRpNl6ngVqfO8NdQA/PA/bv0zzoxZgJHglPiwzgcV8ctJT4Xj/r4xuk7GxVmv8wOK3
fo7d+h00L3cT3ui51c7jZj6/l2fTuZ2IkBTJonlHe74YuyD95Px972uv71Lm41ysVqODqDoaaVZd
eQWlmmbWjrG/ZjVqzvytHEiQIlY49KeQlVKWxlpSNdzRNfBfsvSECMCKycCqAFt2HIS9iwS1SA45
C9hC2GepXwNiTc7ptUY+rQt2Igkuj1hMEkO/Z3xZnnCCZW/BI3ll+4OUpBitlI6XjKDnYuoUfbxh
1JHELSv0CadDrtzrsoKu2qK+5FQGIXHCuc9uB6B0mkmW4SCbvdpoU/W2p6HGSLORN5+SBcdG8scw
XprMsig+PUteTs9siVjZnWCeNAD9l3HA8UfFFvWkYljLxL/n/SR8/2Owoca0bo2zSluvep6dUu4D
nu1z1sRrpE4dISjuCQJMD9LR65Ez9d7Wl7op4Qs6etKBaTkp0GcW+7aI8t1rw04GH3BeFu8iPXOg
vroW6uH3LgrDD74v99/UziuVxlznCZ2XIrj6WE6eRid18t3Y7axb1AwJsMbfSjJVpnu0zECuit9j
Jf5u9CR4dtzTkdfWJqRaucgVyMfsagkIIysvFcHDWJo7RjvgCcTPlMlJjfyB5hAH38anJZEw8zfm
Nl9uvXrwSZj3Ca9fFVzdIP2k3MEMQWYWdIDx3gFH9aBVBiFu3yDuZhfTNAiu4VjH0QwYZDe1R8pL
C8/XgTLfR77dhFPIKQTyHjiOIRsZaAphLAng+djvTLel3q+fgwEn9SF8fIpXgFg5rmnepScrn02J
ABCwrzL6vmd+5egJc0Otc3gZDPGqp+EYAP4KhxO/uNtdKGJ2yukJm0svkOguyODfN4S3Mi2HESdA
Sdh9v3IxZbCrgVZaOs4KpN1te37Wjat0rH2bONP5JBPvWi4pQSEkO7S+c8RluacmgQVVlHP7pem/
PqhWPiHKcSVA+at7uH6sJuO+pwycz3OxzlWYUFYRFerwYG9DJRcngBAee2Amb0Su667IoYQGGq72
RftS66jb+x0ggkkOC1Dn+gOU/yO8uYyRlIR968Q09y4HTdvQ7iJixSRmQmMUaPz1Sg7lmTPrUzT0
LwHJmY09lVHlMmlunw/MhY13gOTciQ/181eaU9XW/YkOKgIbsvVRqFIMO/EB1AeVnxuLXoAFhleY
yoQCavu4xOWAhMcbYuatSSLRIuYiZqTciHhGClRi3EePN+vRckA7d3A9oey2U5zVdRkwhrT3dx1L
TCJVR6mAb7kdIkuu3w1d/ucrBwmhQTPEiawG2tuNlzSKQZBpNk+zAYl9m/YbXWVCcM6AeHWUlS57
ZPZpKZwXWre9OwiooHRNaT4PsUaJW7MTpduYMQFZnoAz9krpJ1IIvcZNE4m3xjbJFDOctJUHc2n6
nHimmkhwsKXZ8hxpfFnHZzi0ueFcFoyW1tcpDcks/mzhQKnfgu5rMKBcY66Bqf+4z8IRU3uu+sXD
/+fbPQksvxj3qZVQzKQjOKSyFv3RJZ83x3OcAVqoZ1hDSXXKVmCE2om+ZVWSM0nWhpDU93kzQQp2
h7BfINi7weVBCoyZtw8aiC4gBdUoMYxnD9DMtZBIxXZfEo/R5a4m8CkfUgPpAeHFlpftRlH0PgfT
FmITDJm1ji2WDVDVA5361FNQk470Tk9DF+R4Aupv3Guu4vOYdlKfcigEpHCexRsD984l4jbcgFUW
MMRpJ+Y9K5aoWGgIJLQbDq5XLQV11OTw6USzdyO/LM3ubsFPLbDwVGjYhufrd8mf7gTv7XhCfmd3
AU9dGshtApeewIVAQZXVQr/rVojrMiQaaWllYq62sh2AYjeo+OQ+tpTLHFpCKpNkfz/2mbEvJfYn
nhvmhVBs39StdJc5r19Ymg83c7ZnRgk8QmmK+CzorCS/Qmabm5kTjL9b73biRTVRIWUtGw6S5nfs
NDis//notBdbVAz+qvp8+6O3RYfaIMDmgi94RIVq7SqG6DYSM917ljiabq8EjBm005VzZ5lKSBz5
OCBXt7abzzvIS3gxAV5dJUHdQzBfag2sfvYPuR9HDkMQP7qwaWY7bCEHdBHVj2scq0tRB+xVepoD
4XgKvHGTB4AEa0g/Pl8wb8nfp/D4Levn/fmXgWyOGEsG5HXeMmKQbgxB/eCGFYoupOmYQE4kOOjk
/rlsySo1F2N407f/jEM4hXeZ0vIFz/+45ggpBgUun+7rXFkOBw46bL50yPoVgcTGS6wFuBYuDqiN
fFs0WlYrJVJph1amva7lMfivECBPgjQ95s/fYC2QCdiEiMv2Hxp0eWYCVnkSO9IcBktEpKcXyR6Z
cA5rl7v+dU7xCGYT77kHgAKfsZxf2emzEM3vfAt0CmRWscUVBiwqvuzaDq0DA0ooOiXczcgbNrZ5
2sEQnaTLH8A9sgpDEejk52qpC2u19pv1kKUfAAmpjR2D7aoceIrsEKhBR+C7jt9IHEz9bj/OSsJ9
HnYD4yTlLt6aM89ibHh9a/cy6RV3SRRV7eczMttFLuXKra6hL2ehj3XsDXjWFe1ko/YuOAOulGeB
Xh6Z16PIIZPUUOl5MFGzUoh3yBabpxJiKKN7X5dNcj56SXPQd3VSmGgNfz63zcEQ4JtVmO5q5Kg7
xsBfiL7WHj7b/k/ELFy5LpX/GXozDeOBh2YoqYHpa89dtKYh2o6JF+DuQipQBZXvRyWwtxE2WV4Y
MLAakxJBFMRrpV8YqFW+Fw6utFG0vOy/uFtvviw2+kD/6p+cGEVIKmvEQd7xb1PndSB2uXBhi/7r
asG34DNztWSx9dpWYog/Uyqxhd0bzYpSaMRK0XHWGoOHiWpEvFWGC/D24jRA9tnqoOQ3ctCDxxP/
a7qrfsOVuW00w7ptD0plowr9CTJprLwR70YVH9zNO66RDpF5cbv5nsLqnm/FfUXsfpIwMTCbVBQJ
nDtzeOPpIhL/w9A5dhO64c7WVBvKohv116mGORyS8I26F2TaBuKb0/IDSadDtyY4thGVAZ6Dn4UM
mFyXNriYRurMHgiStDlSrk9BHNj1iiNsy4tO2xK0CHxntTQ4+Gn9SEiJ81PIlZcZrei2BI/M5Jpp
T1Vz+iNvaRDEtBF/56Ybb1e5seQYALqcNKqhiLXv1NSdbjI/47sdDGBLWSZQ0F0clYQeOqMO26Xm
9ul1Jz1O8DYOe7AZKlTPTIfeJJ+Tdax0Q0ZdR24vrDxNfjq6FseSInyO/atb8NCUI1LWXH9e/Ukp
ODk7NqONNygB4F0wHBGkcH7MN9ZCa5vyMn99gLa+2DjtKSS6FLe5su5ea4iBpoPHP9gfa5T+zj3k
CD8vaTe+zaXG31z24tDG3sd0FjdYp1DSZ6R1Z/JKXCYipF4XuZIKEEmmQ2b/dD8Nb9PvkOzMq2Lb
Y733JodQxyHlowaa8g7DHRI2oAYtr2TM/0IkttYFHqO4ZzfmZmWo1IzWnitVUL++toR6a5oG2Vw0
WzXtapO3QfQUy6Ra/zTzeRbjNXM/nWrDrFMc6tRzzUA+sDkW8Jq7s8IDa49L4JdHDfK9FAJZhppp
LOMrJtmZ4KqTwT1+0sgI5PXF/j9otZPkMD94bQN45VN37IKFFiXcCk1OcNR5jwOPbwfvbcr4BScF
t8AKDNqU43E0YtO6lKpAOl/SKldVt/4d+TyqseNkgvNZsNZtKK6UW4hWiK/DX4FMgiEzpMH0Vmvh
gcz6p7XnCmoUeVg7yYiE0Y+xDAow0h2Wg+3xw0w/L/LIuY+xD3JrrP64h27xWiuKERyHTJoZsFAk
l8npAw7Ytv/FJoK0ev7E0FESp+kEguOOn6n538pnlvpTYQDlP6f3zu6hZosrvKG7g1Dh60u3TF8B
y2kL92P3xoFhAtbNLeWHAfrHv3mSkrjD6em2YihZ/8hqbUb6WqyD2lmz7Wo8c/GwjvgnbKRZwPck
5WbeIqQAPEV/cVq024Lx1yr1VlVpurPVYs91/XNSVnI9yx+lhRFcDNz6gUyygMHJXKvTBQotcugn
KLh7egMYR7E0wQttLjSrm22CHR2ZsIFYlndMcuLsfbovmb5dxorDnXABXqYC8VS72R9IxUVhizoA
kanyZEXXZW23VKEkxhnarsxsWgaaZgP0notsntVK3Vz28/4LzxczIRyzrnrE29bT9LGcRhvhOTSn
DfQY5ycz8P7NfrZOnM9ZhRmPHye9NuKL5U2zIudDBNIRkBpTwRygGO5/ACQW6FnDVazc6Ag5ZM/c
5DDJ7otiim4hCqZ1Anweoj26hCCUPBqgyCnAOr5OzS1ZsDXEhbWoAqPaGmMcLOCAXCNw71t+8Nvf
QXZaIi7Nx9aMLw5LGCKEJZKdf/4xEw6uo14Y0ZbafQl2Geu/vkgVaOlUDoZCzhQ1g4S4Udf5A3t8
JdKNCBihsuSSEMOXM4WWySCzwKKgP0PWnL6eiuRyeb/DavVkhdqfSHHscdsvMFsm8XoqHLjFkCfm
axY2dSAIKHwNg/6KOcg1fAgPT52zGM2+00yZVFfVyixa8ogx8rwg8Jfs3sAtzjcPk7gTG9TRduls
Rr/truKDeMmIVkXpkegju5ozt1V+wvpyrwoh+wB4DWmJUsjgLUX4MWiOpDKc8+heX8e/9tH+lJH9
uZcTM9PgfAnM+YLdq5LihlbDVdH6dGF9Z/LqpzbUwEL9nKnHjDgMaM5FNEv2vpr8RtrSiy3yTVab
EgyMk7v5KIFpGNBwr4YCjr/4t/K74eAe6OriL2nsOiEcIUIsScNoVlHcr06oaEV3TA3rrOQP4YVQ
AX+nDfYKAv+Rsc2YvAq/4L/WUMybbxQdvoXwkcFHjUXATrSvorerOVbSpTSW1zjK5Vq4HJHR7iYr
8AeWgL8KqpvuSRW8oHMVR8rMaQPs/Z3KLEaG4o9DznNqgdqvvc2OxwRHPGC8pXM9dkP5exgefbwB
4mVKVJ8Y+cTYoFzvSw09ssmnsn9HwXgo1OXRjFJb9Gqnj0M9MKQKD4Y2Bj3a+WwP54v28y5JSVar
rxF4kFmqg3Nm3pI62SKVVF45STaD8gWJiJCrjlfM2tWuXAX9xn9VSUSnevbaqmbSMhndCdOP133/
GB7vHLTRlcGS29t1KJCOgQ9jLLGPWRRNKxmE9qZndfO1fhxe3k58+hsy49VRE3H+AopIv4mQZrci
Z7jkDZoWRHIijkmHkPSCiJT1b0kXs4dVkDHxE2sBfxxFuynnvr/zioJVuKhkHJBLATP3JagWFEyv
qQ/STtsL5nQzpALD02Qk4h0hakntpmrVOc+niDfex55nPPOrC0Evx9PsgPjd64ZqJ3qnp6X91Ct2
yS1gInZchjR5QW1ieL+b+0JyhBBcDjsz1vhVfoxlmxpHWENuT0nGYGlk8bcTFBQWYVA/yXyME09/
ZYUuoJqsTHuKzlne46RzHL7v0fprP8vCZSJ5RiOSF2dmmQ7MT8HSoQzVW7qrJW7TnsOKJbjbonEF
nFRVJR1dl0+nDgWMEtTutAxAt8L9UdQOyseH4bnyqcJbBkAsD9c3LMq/L7C5umbdlirImiPcPevh
hcqnZM6PoIbfvS4MVJWNMGUcjdGkN9LYdqVAU83Wb/awZFWnKjn78cloo4F+WTy+1WirXeGoW9SG
mKNXv9zfs6qZ+it5GWo6co9w/Jy51vkZuDimvOQC+tJT1cQIgQssJ1tNhTQaHU7AYEJVf4h9hLcX
yZWd+h/HaKyr4g71xh/XSc8N2XenS5h1AYgXZeCzLM7JV5AxvCWY+B7prN5q6TUWc7vP61tySrxI
oXllk4PhJhzwptzvkVTW0Ot9mAZbZYXl2/9iErMyyFyP6CzFya/4jsUGHXVzuLYIplXK76TeNRSu
oWUC+RX5WnTLnxhwWqr05NfFC0FmVRHHdV4dRcIjLsqA5Tki9YTU1EHEezb9yrzYRbLqiGorYG/9
Hv2UOy9FBBEhhvRZ4J7HXcQD7sPMaryjfLjGpdp6QlBf2pxv/UrylU1qHsVUA/xM+UD9m3KaDzOS
Dq9iXs9AktAch5JAa+mewPCliwQCw9Zs8oMW7REL34LT2buusCJUgn9oSOTtJfrDti39X9crSdIX
wxu77dwChX/SjCRbzQGoPhgqhMqeSo/eSspE7/NFk3V0MP76no7wofyFF1mmCR/Jmok+JPp0eftn
7DnR4pFv7tJgyNd+tP3cZg1xn1VzYrjS2LXlVG89g4cq8fHTmsn+gvWw2XcCQSljOC6MoebxJYQK
anDfDZJJVxeuobmtABfZxyjKN7Kjf+8IeFQas5YxzXvZjHHCBseGfOT4x5XIyMSpFeipB2HzmHyC
8NmGU0xOkCnVvH35BMwYaZ4KZl3gqdlXs5X4huB63BDRvoCjZv+qyCiJuiXBx1Lp1t3J3qkduNU+
cHdFLnMZnEAVVoEwtqM55qYf9A36RecDXQqo7MPAoJK7dzgokbVjZPW7UORq4hnLDxLl/HjoehJX
Bj+V65RQ4n2jUH81BHURfXkjftcJSbx3X9gBD05CauBawTeD/0xtKL4Clj03yh6VPPYGEWZ+uWHn
wQa30vzHTM9SbnFhv8FEnj5DEsUglJzA9d9V6ouC8CoFaX9NQQhonOHU5J7rvbEvJc0rxCfGPRaS
n55VUdCDLt7XKLUNfZ8Uzo2PpFn8wUpSSEXKzh8WE/ROvl98aLnItjKaxQOYt+9iMMwEI8UQy5AE
FLbvTTTmAYx17HTAcmbtpLVYMd4JsqKs1MRvmkV0T50BLpBbEhJ38XCfdPxKqUXzSgE6wN+2purH
PwL4JbBGMCyVIDvAea2/SgxMwxCcwcmhat+FbDfg7kZWv4h+bOg+7A3WI6b6APtwoM2kU2XZpGpk
KOHq3LMs/HkGcEMYVPgDJ8ITUQHf4e7XogntM9lSu1CNCuCuJXjM9Td3htrKfX/moBioDD1ampme
awvS6a6o34WPO2c3RCDJ9a94XJ8T0gSwYsU+5oSO7NxcVI00DRT8XPb0aru2k0HFB7G6VqhBDDcM
TWTtOKpemxveCr/vLtIVjWU4ht7i0PoBJdTOqtLmWyk5lhOq/BQtfAyXFn9LODlGt8r0qgqB4g9u
JbukXuX2VeoWqMOqKYbrUJrN3/NeNYQp9T906L8bh7BeyklDObc16nbk+KwdaDKcakix67K46CJi
xpzdsydTmezE+wJitAJkiXd5oe6/YrzKuWXDGDH0Jqs1/XHqLCLphzW251IklK6jvnJmYMXj7MrW
n4jg/PPh5J9iQJVgFPeDqnBlXjR3Ugmm1gb52MA27CAH7h+GRo7Tem5qOVFEhtX4JR9JbECl1sbm
gusQFH+lPVCMnBHH58ZPzCc2ZgGuM/srOLox7Jpj9kR5qeTFnHG1Hj8lPJwcCA/L7wIeDTShbDF4
tBOOmu9LTj9TgN81mzZIkKCVhsxqKVYBfuU+7QWaa2uunbOa9ILID2lIcZSWiUVgEqmhwcp5tDUk
AcRmJnfPYnzQNHBD3YrO9+bUZvcc1fQuA5/siZozhmrFFJVhgJk14ujnXYU6FPX9RPd537HXygqc
YI9RYjfFOlttDK8sqrES6qyvYgbwh+pocg2JPgbHwACWsoYEwkA1fi1J8Tcmz9bpvzpATU89jGqt
Z1ELkIvAwD0ml6FM1bKgtQUHNZvCNVxOwjT+lEGvXHBA9Cnhk02y5zNYJT5dYMmab/IWT3JxHhN3
gKumu/egiDVm+mmyzMhilcw/FTeGShQ9jt84wn/oSoNeqns5hln6M/D0keq8NOLK+4eUyH/3ltxX
k44tWRiWcGEc0AW4jlFZByN6ijatsnWxkfzm6sn6+dxBxoEspZazmj7WnKIyX/EwJPfoNJ81J/EY
T9cBsxvVJUsVmnTWgaRC/znUJmJo8xyPxqsQHHOGOhAZSdITcCI/zZKjhdJl1ulhcAHVcHhO2pfC
nf3AHhEXJ9BVNZGTTkiD2lE1guWYRFjbAe65Cu8q4LevfEKNzsJwU2dDNlq2IWn78QUbdACLv9Bq
It96nizdo7waMHKYYFY+jaJlJPbKyGnQybTYAV5gAYa51ntoXWtb7p8eP4d2TLVPcahzkAiZkokX
z+cieYUFNmAqZ2igGKpYfxuPvKOgmxwTOKD76T8HmPZFRxrKQtyW9HE9IPtef2WSpzibSGKGqQAy
PnokdTuamQPKnO4L2vJa+8ohMqLogIRGmDZnWkZ89qQnDdQuiIRLzUhlrdZMjcw83UC5SDF1SkJX
N7fIXVi9Z0EWbSw2W6draWmHzLA7GhbVm95C7i0aAT6m3BjRBY23SAPM0HM7xZdSvOj4zeq0/ayj
1TmVxaXi6DGqJ7HBxO+G+EEdj8UQE09hRLlmMxLFR3R5S630lRUxOgVlWdoQdaiIHhfPyr8BndIF
kziEi5NV6wRAU4aPqt1O6gQCRJyG386uVlEN8K/ZztBu5jijCJorYNmYKKhkzkWAWjCDXhdGgyXe
sd8AArS2jlYgzlM1HrmTvETNe1JBe01CuuQNKIFb25Au9RaHCPG2+epRnkERHID9p9peFYT7eYxZ
2dqkeOiV8NDeeLv0E4aeY+fsEb6jv48y81iSJaJVMo/NAMNUOYRjZkawp7vgMubhvv7dG0laSWV2
biz4YhbFYJs4aAVy2N9nYlZXAZbIiEV8kxm9EjPXoBei0czZ4UzJlBxfh6zfV1U5Gm3YBYBtWLfl
kWP1Mf2NlsDt0LgAOSQP8AC7uL5xlk/xxGigEhJ8Q3wGz/v4TaRG6AbVhtU9XAz8bqy19cIsyjFf
eUdFUBLXMxRkVewTze2zM3m2fMFQT2XmRK0B7wgfmSjpZXzkBlTH1ln0fu+ALlbcr0bPdX1LHrpS
1awAh59DX+MaHJ8Tro0S8LDo7EZYpeMPS1Du+0Z4EDRWLV9qTw9qxbX9mtbKjPcBFTIYP5KdkdSj
+3HC7wc4OxHt1xfP03/vDRicCn2Kh5S7NDRU3KLQ4CEW/ekpujDJvtSLNLxdd9J7+PQNcxiLqrxq
PHP+RltzQ06wVdGN9kX+CV9Ccq7aB7pjtPns6Q4bTMuqc6/Vzr3/PUxoWU2/DAPov8YpeglWce2m
oWpGR/IG2s5fLhLWKKeQL+vtjREr3vtXrFF2RU0YYllpFY1YDftbvzc1y96MvFQaynzUzVfqk89q
hF6vRDvWk8Pgs/jBnRNVDll5Pyd8OU0p2h2yKubz55Meotgy74GYY0HcZNc11+i2rkgpcK8nJKuB
8Q7hzS4hWJvR2SjEhozbYqvNOxBvZnHDoIZm+il9B2So4rqTx2YIN6rRlSndJhPdhsvMzEVh4D6T
8H6fOtLC9xw8GzZGs5qu0anhEWeBmhjYUQYf4xjOX60fk0To44LyTrWVxI+r9JIcCKgf5tpmz279
3SRsKjOq4B3WMyGJOLx0YThfrd7f5UWzpYCuyFh6XClmvTTjkqT6xMVgzF0ZbmtxqKMyu9YReCa/
mFE2ya5BruTyVdG7Bd6A1hmpfQDzk/MOrETk0G/OMe4mCHEsANmAeOdjszEjcyAwWEWExmyL4/O9
kHkObBifD3fgXFhGEDL8anWgoFnysurDrwSsbKLAriPwkQRf4sjqQzkzl+buOonmNPtmDJTWD6Sj
DRUJkLTCz+Vcp1fIg0DCTYUYaR/V+qjw4X27SP8BUn3PMwTrb1P+lnJQX7Qu87DacjbpcpxMEi4p
1bCR6tHpN6L1clyry2yqO6qZZGzd7do074sCPpdZtubfPIal54z6RYrVY+4eXl+5BDvFZEKp8uD8
0VJ6X3w4iDWzd6kfMmFAq8H5EdyiToCGFeEcdV+9X6WILEOSJWBDuENr/YdQbspN8OhMjttZya/H
p8AD9k8JhgwYzZypw5qvGv3gJucVBnROZe3u18WQJH/vVHp57VJ5ZPtPuljonE8DAv2KF36hnDgh
yA3+tnrhPmqYVZUcIbTFM1KfQggecHvrDLf8nHa5yN7fLHGeR3fzACzijJ85Kw5CVFp88nsZUBOs
yU6hyCDDT5m7FmnVsZOxGOD/wj55Su90b69XvbDsttWW5QWKzNUNbgSPdEFBFX6fkZutNYFwohSW
3ZPLY/Jcu9grqfq9vKYhvtKm8SqWYUR3qmoz3PBNspoA/azNZq6FIoKVCclQ7y6xED2W0/yBLsVR
RtBLN08EdaxxRckADQV6rmCM5JN5z2np5n6VVs8AO1PL2bXCubSEE4l44WSrvXb+LxHkBZDY7CfU
WbX+6lZ/bhP7L+y1cy0qnZsZXVeJuWUJ33r71ku5yoICmmzdegL6zIghKyWLP8mIjAy0dd+YoYVE
8WL5ES8/R2mf5aIXRc4sIwWnmGhKqs7qHPaPZlAYvAjgEGZ+zfj+cRnPCrbpFfI4BvNAg3AE6lTI
SgbFMZWVmw105WSYzx9mh5GrcPe9yYK/pXoR124ArEFB3YyIU/R1KZgXzINUsGIepSB2vEPHyjlp
+vBHzvNt/FDzgUGk1A221Iry9HUGgJWDfeYLg9j0hHJd+zNe3z1vYFLOasedRPV8VuzZmQMo908I
Ps+q0u/57PHFNdItXb6XHa7oFt+knAg+qOw6eVyLiln6it9QqT2Qig9N0DlcNN+bH81tHNvpPR3f
6vjyn1hJLYEwwHvX7m594TlEdssZM0vNNXOOSdjk5YGwkhRXAnkuVPaErOhMP7wf9FlUdC8d3Oz/
xhgoiHhC5vPXDr+bPzV4Jfao1bvDrTUMFMZL/knYg71bZIwkDBCQ8cITtlGBQk0576jQiAalzRad
Ot/PJbnH8I1YqtzS1Mk5cXCxBB+dSRXx2SwXYSMeMCZrAQvZTx+NmR4f2YnjfHzHCVjDvlGO3pG5
y6FDx5aAA8THvToYvZ9V+XAXbLrqLq2wO25hoWJcOi48ApZoL8wZ9ZYmsc9/hEZJcgcnHuavROWv
LYrc29tcRPPcXjIir7+jNWaowUQzMUL6Sr3Ar/4YiuKLCXrCS4DVB7omVwe3q5B7oqSnWbo7PT7j
Chr72oLewcFC3i8a+S7/YWmw6cyEpPjbeCj5b7NwJrzlMiwuYMmCLMyTt5voj9hFFlwJLpegfITC
6oTeyxceH8tAXYvI/gEbuChqxPNO6q73YHWzYBj6eA5JtXU/vMjrOITA1fDBqHVo5BxCNLXQDiDq
qavBPQ4CKtpnQmuncLx60vnxdnmZncLtpQoeIhuh71ZV2mNTzrqo3cVG0/qiufh/zANVJ6qEfZjw
nT5jFlBBOhro7jPOOG3I/3/ZpD0L2Oz3GfIWaDVVfYw8DkCdzuRIjy+Cf4cOXY53q6XfxyiDxPBG
y9JnA2mApS22ajcpUt5yk117QEIkhKW1Rkzh8YROOxNKU5nR6gTxNjAhHCokg3gkGRPYDDBmoLnO
qmh5jZ2QWPcK7mE3MXQzhilHIFcdlbotQW3qnkFQwhCno9+dKTVh9cjZ7UUuKsl2Xv5aX/KJnVVs
x42Cg8NSvz+NnWCD+283xedbL+lFo9JkJBuwvfJHJhknxecaTsgfJFvvrS67pYDAmUtyTSwZ+iwT
kFTnxhxKZ5HLp06gzprh9qspo2PugkuX5yLdKMh7wyJ0GVOYSsGBgva/hwkCdQnN2A/U7lSiwRSt
fIGVpI50RbNB1DGqwtvioh8Pc87djKksLFF2QlB8FopCYDRHrYIxkZhIncnSKCYq8/DJ9QyXw3VB
JZtXXSpdVyfrrtzxFZCbJpcxm13EsP50bD1HPZOryN5Z9LGXPzMVojM6/JINkp0FT3eFtFxszBoI
gfStpM2WJmHPlAW/oU35LcbTSD3X7nVXtUhz8vkrsQLOkHEmdpfDs4PRg+33Bvc33d9JpG+lFvyT
Vvt50DxTiiKN6N9r8qKQISkS7PNUMnmFJV0Vqz4ZH3J0PVbYmpR48o5rKgKncEuXPUCPex6WfRTI
+s7Vmuo9hXkdauTAaMKAsg6DNYCOUPVcc411u85FZNKHV/Zlby++eAL9Pk7Hk9AL1unV/UL175wG
55tqvlGYJKC+t+FiL202tzo6X16dqaTvPB3jiUWTiZq/Sd1OwF0TnumKyAK3nzGT2CyFOn6h5/y5
EecTUZw6QmjmPNQ5nCq7iJGfqymjLMCRufCnHRSG/PGWKCmWdj7md6ospIXcP8pz4tqzTyocDFoS
hEd12UeTD2QVYfQJCbzdrVHAqFmdT98a1p/WBpDh26zw4KpfDVmoBqX7Mo8jhNg58vodQeuadoKu
SWYAdwsiccnAAIKT1sRK4hXDH7S8+vW8CDYQTDjqV5jUeA6U9F7lbolPeZH0fAO3HnD75jZidOvt
or8+f4WY152IFLF8CfuybzMGfmQ+594gHYVxZNgxUlIuDu8jCnSty1nEKtZinUQfUN70C1NdNt8D
SuPt43GCWAOSxuANWHhCDJW73LZUQWFd6Jecao178U8z0QCS495mbe3fOsEDQ3gIShClbSJtjWpJ
pXqGVuGInKRswTusDDm7rbOvvJBI2CcRFbJuYWF/Ag0N+x3/WR3qhAJXQDJUrL3XE0f0FvlDFYjg
/2rwnlZmnoVfZM1bjnCIkil4okiD0+nvFYYCm/aO4wn+KHdfCdkbM6CtHiVpFMdwLtrpcs6V1J5P
W4l+JWZ5fGUbmK0iHhTj5l4BDiEJYdKok2yYj8ESu4PWjgxxoVSvWImv8FwC2Z5x8xW0x2N/asAr
d1e+EqUkrY3uy2PvR+gCCVK6Nhu3GgJtiyyZec33wSHrnc6RBgR2iubClF/NgRejlz+l62tubiTg
JJtkTWSUYgMc3YBj+gUZEv/jxvtjdXDajjvva+4ugr4Gqo+NVOn4R/kuOMwwvxrKMSTmNVc/jfMb
S22nwSZpkKbxfb2HMmgVWdLZZhlUq3eZAqjLIbFo7XnzqqJFI9TDnfHyL79Z8C1UgHbvNtNu82vm
S8Z6FkLZMm+1vjihgFCEvImwIdnEeDWk1MPMA7lr+aGNNUjXnsBEECqFSRkYzT72nXTNR6fiCErh
8RNhso3M9RwR8DZAfdP1MPwmgNJ/QQ75m90lZfz+x1WBgvTklWlSmRwHuh2wSUY5g8Rvqkg6u6qr
tdQYTCuJ68WlhVI6FXONUQBFfScrOv6+n26/yvKx16f3kt6eaeB7ZqJwt+ysRryElLQzUoz0JTcE
pccKnulDSfEAiMdOBUIlV4rm5iwyCol34LOEtkzkm6o5b/8GaygE3an7p2MnZc9oqdy6PRr4uIZa
jtznv587Wjl96qC1xNgMkYYuAM0mDtWZzpcDVd6qK5NZkbOSo1ntyXj6pgn5g2gsf4O0CQ/CEB9s
vgbfevpOSC5nb77aJKdHAJYRtPBIacu15Inqf6sOrcGR7mM921qDDFR9A2z6x2Op3MTFxvN5wzqe
QmXZ0Bh/RyqCoY21qaTLdzJxbbDtjflX5MfswsyMuSpOTw17m+IfI5Zj4jEqmtKcbd0UT77cFHsG
Bdh7S3uBUappE/xhxF26HaZ4aHcCRNehpYlF0j/rHIMmAgT+shsOurQER9w8yhrNXfiOQtuocsKv
olLZRmUvOJEk49UrrCkx7upHvTS4fpeeHFfwqljKFue/R9Co7tlhRN0nGrbY8LeFJhigpOO/0skI
uWMkRMk6wuxlU+3bO+Anyz2tljM85FCO/MgnAyRbbt9wJ/ZUOuJzAdpGqV1jEo7YQ0CWrxMOIeF7
Krjd8uiRimvISGlI2jD2EpJv1q9+855MJ0WK0L1Ljdv7FpmuBuEaWJmAhvL/vZI+lT0XEbfwofQM
dxo/QnG0F4KHilx4AFezM/sogpLJZKtBAtmfgtpsZ/1Re1qF0PjYT6hK8OXufspwxEjjAeqLI5ZZ
ZF0UPZEC277UT1A7sHo+BmxVbDxkTvWBk4mQWkh6d8w2Gp7VnC61cSDDbHaWRqdckcTCETEJKvqf
7wBItvlbRxi2S6e3/Ak7+H4GmynUkg8zRj10uK82jvfs0D+PzlB8JV20WABgX4MWfaW5MEqXKoqV
jI0C/BMX8v+5JQcgGRXqIX6Hw+Js/GeWxddScImJoSL2YD7fbbYs6N/EdJ8V6Fp/k/jEcTsgtGXC
kovhnN6fAbi4xRTK56P6jDLi2XStmzql2H5hQckQBr43eHkPD3JvEMYDxHvztw9ZF5JVIe6Y680q
949HS/GZ+OnuxfhMpxA0YP0nviCUoWQH4XJVG2InsYm7XhRcRKmXw1NNBfOXs1wIV1IE1RzrNCFX
1omMQkGX5amuLXLVLF/TvxjkHmK6IrTDLMjkTdraOC/Bd/NT+rxXzBEf6GRDFiQW2susbQTjS9KH
M9XDMpkQ8USq2lGhozV5VHIIR2JRm0Z36lklQmbZHFdA8L6El680XjIHaYFMJAkfHbIPj/iYWOU1
onrK+jbgJzNo8Wd5Z0luJv3c9tqjqy9P7M35lQ9ZhlN9rVmFG1+QuTEAGJfyaz8G/ybrfhpoAUZk
OXgaw+lCvdNVxCYDe1IPajCVI5XJlkeKTv8NAvqPGueJmf+ppaov86CYYxORJD9HFmLgIxlzH8DB
vw+VbGzMDJloeUKtrkEtMM9krGPIf9M+c+UQSN4bBgbM4eW56z+bFITODmYxcqggHi1PgEy88ozi
aCLtTqKuvFSkLJJpUPHAqv12tIkaxKUof9x9hdEsRm6zmQvdKrcjNzuJ01jd911CFDOaxj3uqlZ5
tYiSbQ+J6b3mlZHrSRTKcifyjmvSO1Oz+qqQQmmz2tBqXQPnF1azi8uPFAuxvnptG3RJJI3v6vNe
w7p6Si0uZMcwkech4VLmM3gpXLzp7MvCr9A3bziY8oMrqmCyVqcOBQMltzgogpj6m4ZBPE/wXujp
LE/bzUXDNN5o16CLHOxSfbwNaMR9Ffg7ACVrhm67pZTmmlj7oer2kBGIPmJHnQIrhaVsllFCjtvO
8zQlUjx55DGyhHaSHm0sEQftlgmRosKtGIoPK6cqAPmTbsZRiNzHvKmFT+1o0wT4pOZqDp+FRidr
XfZZdIKRgr9g2gE8twA0sZmKPDQz9NZ/JTJGnk2FpXIae3B32pG0H/ppMYaHqKtAyDaXu8ZsWjBl
Sfw+lWxtbibsCFWkwdD8OYMXnUdQdenQpTBEUzD+6d5gs4xaFhPEp9bDMdJcGx1rElzGqes0B6aq
ttQiEZVjm8nY1mw6zdORPpXhIouPWMU1TmpRfVfWKkgvjt36NXhh40VdXaZRooD/Tx06Tsgechx7
EwIGwKkJVrOR0VpRJlW2wKpjU3Uny7zjk0bO3nsq1T0N7z81pp0bBWJOJzFPCU6riXDEr/xm5s5J
b7CD/lEZGLgp2k0wy0FKYsLTZsFNHVZG2j8hA/blaq79G0sT+CC/JGFSxv3iEphbS8TWhwiAGVZN
XLLf0FQbGMBPQ1rosB2dW0jgY2PrBwlbX8OsTBdTMNuUHZB1+yeUnurd1J/mxj9E8y7GZn+O5gEd
0YUvLWFCXrF4GLResGr5dZV7KMkKwHTyYc+KAqxZjDSB+Gv7P+LdaDmDSbmBZL227SifQAVLJyP2
aKS/yPOzEC+14GjrLn/M17popDul3RQkPaOrVucXH5b6+YabaNvjRs6NgT1dtQ6YpoISWFyj1z7t
p1aP1SQvOOP5SkDPiXcoq4KAV/sWz15iYOi6g/rmyHik5sx3AoiiVqgI4haMbfVm1AJ82MB0WWlr
SYZ6Vu/fiqMXwiWH4meGDRoEc73dc8rgH1WiD0V/7MMGC9YbbixNkKNa+5z7AKdk8EvXBcxphllX
K7A4rGWSr/1EJaK1wBoogeSobWiEk0VUvywMtrYxCq9Ub8TyFLajJ4dKez1Gz3nydI5Ze+0C5Y5m
4j0cmw21F4z4M2DZmz6j3jqh01SR1yO8MvcJbOBNxc2trUOq18RuAMQ4SoeFFGcgp+plMEDY/CM8
YE7LlnCMqDqgERBcmp4beLgbhMr9d+tchkSkmBdO5gnLMZF7DmUikl2erhczgNyJc3WcnaE2ePFg
7m5YBnpymEnXbTmcN/fCECB2BIHUq4MUE840apeYmcCnWkHnFg82AndWl7sbAVqyz9pd8fL6tWAd
iBTfyUY9R38UNd0UyoQtb84RYKy8sLY8F2wgqPm/lGxNUSXp6SVA1UszUnSL+U+3GZLGafXd58SZ
qGm4LAH9RO0MrHcB5ehlwwjkbCQhugT2xtsSCto06afipMEsggVZNBszPoovlgy7YYcfeqLNkwwJ
JdTbOmnpkgkqwtxpFyso8pkPyqh9KCwJDXnRzIuK2QJM3iwWn2wDQAaOEIJ5iV/nwAvDC3aL7MDj
TYVr9TlAtHVN+BqXjMmazze+jES8CRjzekG42fdIU6s/fMR+GcdJOsWQtldeaXJBVk/x8F5XRX8f
ZzkQeqke6bTW/WZlyzmqDIXmP2DrXcakLKiMk7GiwiAFuki42DSINO3k6kDau1In77NVpZhnu9NW
nw8cbm1noOw3daZncpYsZ7OX/rkA2o0HQAlnAcyqnUolBde1BmqA3LbfnO8VDkTL7IrhjJwL9umI
9Z2CxRLeJCqX3vz7FmPbTqXa/feKGB3mz7HR8N8hUw5+5uNungdCurlhnXTGK+pdkZux/XJVCOMv
ekIM1DWUplRZHxzUt0J7L7SO/Zg0VupDX5MYsfQyl79Iq/60Sja2Ru6N7cGRTUYIavXLsez7QjQm
9re60mSPFZXhNL4TXAJvUpEe414RyL4U1l/cpBmZvmrCVBxPzgeOGkTtWN1sqw9XhJCZ7o3r96VO
o+61oc3B5HVQp3SQxff0763jtWfUevBzwKd27nwtz2z6QAveib3bohQ9LllY+ToQtOe9gJUuzpKW
lWbAYDGUCzm4vK5DSivJyFiJBDtdokv9i3yDqR2prSHXq+JYpWrsMuWdCct2n3DA2D8zDGzNFXad
9v7gDsn51+YsNDYywfQCDBQK+rC2VbgQQOz/oN0r8eKGyxeqKgJKRsZjcrovNmgUIHVpfkG4Pt3b
Rae2iXheCR7/GkxFWb2xQm2Glhk4N4bU/0ahApptoKA6Ehf/r/r9VqYsJf12bpIUcQeI/9ArINN4
lXr2Lv9cd9+etFI0A2xhfueQs3KdrcPLVkYZTBu/70MAuJdGDIp0C1MkaRBlqDRykFcZausE7Hg4
pEqZdp4uuoKBJ3g6foUza2fkk6dJC1mLAskfeifW9wbaecL0tiUgwM2wgZWodsAgihw9gdy8h89p
jlOmsrLf3TfbHUJF3ghYYWLYb76/eAVhIuTM0uYv4fE1/s3HZVCzt6aCcXlTHe3EW9bvdfvvK2RJ
nGyg+yhX/m1zQm5z+pr2j5hoQfJ7mT+JXYup3WlwHP1Lxg7RqEx52jhVUQcPFqG/7vVcw7L/eJdY
rOFKYCF4V6SZkMAY3gmyPN+geqTZjGhgczw5KNswQ9UiXqdLCakRBHpNDAlZmc0Ut+fqDTEKwEuN
mxmCvbPdsu/rLehiSQwxw1luZ1qZf13xeie76RVwYN9T5o2cA9Xr25DLlyHoytJmRhmrf4ydQjpI
FN48txphP4p36wiaqFFXmqITvDi3DVfEOghDMinPIEL6Ff5L7kc66wDIy9D8p4JgC/mTE05Vc6g+
fMU+HU7VjoVu+RqS/bd0HkQAiBRz5UYp0WfqURG2XRM+qLOEhFjCmLgum+k23h/iPdUwdIqfOW32
EDSCmYQiLN9DU/XslO0BvFtkTMFFIuhL4ZVmSdh2ae24dPp/dTLT0jdhao0aKhZBVLGpTtnwWLEz
JRvy3Xh1YscHKhcKh2H46qm9m+emd15peKjFJXU5vMZsMl9LS/RZaKUueNs3ueZGxMaNoLuPi8J3
gCQnNsDBeS33yUyDHpuOyUbxKsleZ3e8FXtisLDjyP/Ny/ekL7a1q2pL5McpMSY3uL/pzX5QUose
KVjzqy8t15xBAuX/eaR4Ak76c6cHIVNdGqRV27z/2r2E9iemhXeOqW4tSzINut4zQe3SZSHzAbeh
V6AmpOZJclhn9+EiKH8X8O3ed6GrA3zoeRzkK+MQmC/Oedgmsb0wMdIe0ac/Ruen2XAu3RYIhM73
bV1gWgmFLorqSf2HlsnnfR0atcSQA5vez0afDDLADyCkqCKV5TbQZ572j6p7O/Khw+l97A3obKQX
yUzmHlGIMDo6A4G0S+uQaTADk3NdW1r3Vx5pf6UsGjUZQvDF3c+7QTyxwkBv7QyqNDV9oKxdiUIo
h9yIwuVOQlbPep+7zeh7Qt9yuSwQ5fJK5JDNldVWRpq/xKfxLppwn2oonb+7/cYEynJyRJgR/WOx
gDnUFpfl84FxjMkXI8dLMuNZGp8hcCA4byGAW43PmAXasIRp6wQcYHTtKKO0zfKyp33WLMuj+TR9
60z116gNiwIlJ2rDxCsZSlTGq/9usngjlnZCMrFvfWHYhieK83yfI/HIqMr7gxLpwFRQrPtwtITl
YmpWOP7I9U8FSb52DxtrvH9wyNzN4M7V5e3pyZid4NPa10gZjsKWuURBp7IScTnThf5KiRqBDklP
/5BI6DuPVCvn/iox8W8EBxGmdQFA1mTZLXcusRyfKPhkKN8XHUo+/5FsbKbMi4v83d+xAz5vw7W+
t2oL7WFN5kg8Gz0qHOfpKhYGaJz7TWq23yquH60bF1MZ5J0cxrKkBa2jBqTViLJRYtCT68mLR6YX
Q10zIs8FNVWNtVsHimG04cjAW8ZBKDWO0n617rGriscgTLjs6VanAqbmnHsQm0iI+o+SKka0SIw0
ZM5wrKPB35f/oV9W/GwvBICJ1Rg0P86VnylehUqHk/IfhrFLO0ueLhvNaQfOWgrajbiiVlxoTGiK
kYMKoiItf3ruhS9mvRv9ltHd/1ORqM9s2ZUmK/fJ7yiP5rRAMf7HRIaz6rAd1k9Vz0ELq85wZk9l
ca0CwSZxG+cpI12O3X0k7+OR26qeiOvC76Y2jqtkA/Em+xVNQnRdoDOw0s8IXpoeuo8WbUA2Bj6T
epVoR8TlP6Fn9LDiojmXuR75a6tj2wJlLa81pOoivQIO50CQQIS7Ksioj73mCITn9IEXYeIkybuG
8karRHpm9GNJ99V0Wfq7NqDAA0GsX2eqfdSrp0QIW1D0XkZiCQYN/xgRhPhFj1RgIwD4dqtIh7Gg
XeGR+aS02cjC5kvQ+QVykoJGUkfeh59xgUGDsdQYn6PaEei71NS1Hu2B55aayAIwS0NalWns6qSR
pe6kpEEm0gAwIASiD4x3LJwb4Z09Ri3zQshlK4tp6ijVnY76hSkgILCXZjsx99m0oziUCzTuSSz4
ivuYMirY6Z11pKOrplfpxFFlEqjmVX2nU1tzg4QSy0ljSlTRI5QweAsAcPFIW36LBcXDNCOyTNhT
WeGtPUBbJaIfCBMOBg4affEbtKQN8g3gRrfB5YwNBdc0QhTvpfil7wRHLAOw8bMJ4F/kYI/atWtq
Ymx0lC6WpDLLpIYucm5Bxd/OrEWmVeeyk+b8Cm3h43upMSy3eHMJW19NyFtCO2iHBjUB05ijaXe0
g+hWYfeDLbmwBJ0Gaq8N/LdA8UEbyddsqe6UZAer3S2WMHptrGOq+YSSUvOZqOI6rm9mSPvOphVh
Dv2n45JXitxudoyVKnZj2IpRx/AzQalvCe5Vt1JS8FYI1OaKVWNDoliIzUhgrMluAm8Q838LWjXS
RiAyfGlVSWyGrYefw2LcGm0LLWu/PV/HWRbV8+/+eoRllwIOuWhp6r4gcDPZ7DOboSbtbykfT1JK
YaH+fJvr+pnrPNWOIXlI8sKXJagI56yjmijQhlvV0dd1Yi0bJBpb2Q2InuiBunKRwc5rXVfqp2T2
ZrNet8mno90h891KN1oDp9Y1fgrdkUMqD7ZPcrqLG7y+9z7L1RAuHsbMnQ6+jryWk8gte0JEmgVb
k04auxPaoOWq48800CuN1mJ1ClTyT1O8xLAGP35ECf9MPlCzbFMT8A+9qI2jFoaXGyE8Hh+I9cw0
i3v8rb4hCiWzdhOGZ6a4gGts/a1EDRb4cKb6J2pPGgy5OZGzqnaOk7RqCchyc+fDS1XnbWXrJYzg
Ie9re9aC1Dcf+HHtDia6OZlvEkKnsXet5EWMHebWaXFRZYLUgCoJ+GviwhmFtkF7ENiteF1MQ1V4
ngraXj14+CSwuTDC3r7sMJ8LNRLLHRV6GKP/eXz/xVRIu7TwEpW00d0kQ1nGPbfVsfpqlJvtB16S
jDQMeJKiNOLvZ/bIfTVL0mBLGX58RyFRnYL5qskFsWMRfpqs+S4Q9iXM6cXgPeOArE2L2DD+BuOt
960mKcONok4juN1EMYqHvHMKhXNIcFJ96e6RFQo7P3Wlj70fqEOsm+1LtLuuIywRJOfFYkwoujJO
GwX6Echcw0Hr+AXYNOGyjKJ6yS9l7bpT+piuOaiY5k/kbaDWhOF9I1Ub/8kuaBcZzGArs68hYl5t
0VFUlQMgk0IR/wIqOb3bGMjkdXgU5t4SPSKEWeob4YBKWFNS8Sn4GjoaiJcRZi8WBqbJpmvankVR
rzfxXTYAcl5UsQtwJmi0PD/8lDjLA6w9U+ck1oatIX4iynwOUAAJ0wIXlOktoQOjUE2JK+k2WxW0
Un/m3EczF1LBBPszkndKa5Cr8RAMP0r5gi5SLoyyapc7c1nKZjKumhg4dtc2d+rDOrFy7VbtC3ws
DqgMr4ZeepZXGkVE3EX3FmO18Q7LcZwTDfAubxewUo6IkSFwN8I7J+77tpzW+DIenSgHHX4MZ1Nh
0inte3c4Qp3pWNOEx9WE78avgsT7PeRzEF1TkyH4Hy6Z5KhD4wASFRLstfdBxT96iQAfAZPQUUHc
a/ib5M8hs0jddLnLigdXl7VwjGS0tK55nATBUY6N7FbIiV89cU7lQbmT8rMvbAjEs5BMsilf8gzT
0TCBkK/DbRFuPmfMnwpEpuNUhJGrvHmk+FdXMvKc7fxEPuushu85vRMoQR/6lqIiw7CIoGFx1j0z
gTgRDTmIUsamxizcd4QjxizZbUx16pW3ACAIoPnuHBPZuunqOWADMUF6KRiHUkeFyb3IaTYXoZSZ
bKBsan0LHSFrDo/8LYMybXxOtw27OuMrXGiFrmz0Eu2oLVyMwO2Hf/1rHoDIT86ULDFrw9q7bgM6
e37PrlsHOZWXxqXeP0ZpH/mGoNzAyjCytb+VryYwCaVwf/VfetLn+Dkn2XB2Dt1YO7q8DF4D14Ab
HpWVmiIfZHV+Kqfc7SuH094Kggk/J4fHLLS3BYs0yKneJSCM77oMpGpP7fggTF6rLOqAHLiwhwTo
qdxhjmvwzZzNoOumyMr5T8Tg8oBHghvuc+dGQt5s6maCs0+qIrso5Ij8L/enr+qMpW/1moD2nW7Z
GdzIvo3BJ5g2tdE9apN/reZc3pKDgftN8LSFZ50dr7UnRpYgl4cpigumqSkKQx7KNHBLPxoB1PGi
QtWlwxANOAyRtneoHkKxu4b+9TfSSDim8ahKmzuLpxkP0Abl3P+cnqFPbTbbol1le3b+RCrOb4+V
PaBwQ1QbAbv9eObfpokdpkH1biS6UokVpJkYDhzOKUmfHGDKTqRTz//klRLnmQLQMJmug2NBsIv9
YIuAKJhLroap5Hc/fuW6P6qnpa8aPdqi+0xdhiXFu00WAI+ES3cUxoau4WgEx7XvIzXJkOZmUmwN
JNSlbx38CeevehtEIXfNg5ADHBmKn+P3iR4MqqsZbw8Sz9e8J9Ud/xirwx8wbuVG2GJClgyCQNyr
Cx3s/Sro5By9SpBX+Mrhly4ThWz8cnw3dpMPUwdk7eyLoVo70Fzh1liknlWWr2HoEj1VBJ/dgqkA
PR3PMd2B385U6TocqLTWeyS4RPgPumMOq3hyPHcVbS4tBKPPiLGQeXh/hurZptEPwDXbfu4edUsR
lMLxcdV0sXdtEu0yLNGO/9W2TZWI1PEL/1XCoPCzCIP2ivuaoRagZjH0Umj6+z2mqXM1PLbgu/dX
Uj8AatBX0oa50sUivxRMH46ZmIf1wEIVX8TDfOA7qatyS7URB9Sa31fAFSV5BznAB9yXArM7JoBu
V2QbOwQzPuzMpRf63IbljrUFxr3uFheXCvMTSmeyAPFIWJwh+bynUqy66j9lIgx7HuvmCLpl1mj2
H08C3XHS9pOr3v5K5NEmU6IXQCUMxisYQ1lbsLznD2Tfk166IgwAf48z+pkO+f4dW4yOAF+x08Uo
rJwA/ykekvkjvV+CBPWHVllDJPUn2IGS008Lc1h+zmlGaoIC5povpE2gvnC4xym5rHAQLpm3ZmSG
cyPE/rNdxqFnxAeia4BEvya+Ytywww5wdhtCbAuF6ZOhq7iCfB4emUex+UxKOpK4jiGjGEhG4Gfq
rSKe/djMZ7mUBYVlS0nYh3aA6wx2vooyB70smOoG6lXNer8K6NBL/bB4IEffX746yU7Y+lG6gddq
EABv5avxcGBSlgUcPa7PRMZpMvuu/JhA3jhMranVUcjZkjquhOAKqv8oCXWt8DAdhftToEZHGs3t
I2sSZhHBD5n27+igGwBfKvoH7xgW2sw33lHFBML87eY6jYBm9c8iZ7MARQTLz1tjgusk6O+09xcS
D9/XJtdmIf+AN5XbobAfRNOuBVZU+tqIAuWob5t8VggCKKSE53+ib21FMgQY+V6mOojOaQ0+c5i2
OTOvqr3Fwy+n/5bJGJYAtorpiRzB6FnAl3r7pjghZfhH1GSO1nH1l1qELInD4RfMnUY47jPIdrR5
mM4zW6d1UnPhxVBlw1gYtKM+7sJyDyCLioo846Ge7+veP/HNF9jRv9ez8Qql7quvnckrQqm/bJiZ
K3SquB8V4XrUEgJjRR18XWaz5A0YgiYBNpSD8sO6kVdqCRHRK6cDyTto8YrtF3Bx8HhBOS96Mc/0
OI6v2L+ZBntk1ztSM9K/Pudwnr85fGFAvnU7YNpsNKIOhNGNo6eimgaEqYQ6ATLI+m9Rb3b0BZjR
h4nJN9zBLD3fuzgaIA7CcmujozGp0lLl4rRJ+Er9tz419eGp8vM0xKjNZaCWUTg3tZT1P5bJTvzw
vxRDGPwaP+4RwJ5yNSvmzRuSTrvW0qmyGiphV6izosL5S8RQD5S4cx4HiFZGi+CAvHIMGob1b7nV
7SY211s/xJJjXZfK9VKVJBge4Gofm2sqBbdH1zrJMBllyC4kySD3WpIhkinWaaPQWihXA+fzp2Vm
vkfHGildP1csggsDWwVvYyGvm7xKy3dPx5SK9amcOfm5kW5ygXJ+iQRFWiM6tZPTG7qeiTrUXL2K
b2mRdlSMCWcOpno+q6rpjnGGXpWbAAOGyioY15me4p5xielTw9aQ1MUF6gI1WT34jNhA4+naLD53
PqPLRc2Yu/NrJH9JQvBdnha3R0GoAEzYa8EgDbYy+2Pv7ni+TNZjWfBSG+DTM6wyclghVeXL51vf
mDjmSpK5RdfY2Om+u3Q7CwtuAX3diC/iW7xzTzt74IP34cxsRmI3q8qMRrJZXoOb/kjAhpYeLtl/
ZMfqWjywN7ecgpzIajFSrgjpUKJRcgLscABVXk6KChToIpKpMtLcRKRRGeCMDAdjpEUgbzcmhLoG
PSkAdASOGeTEasBAfDnKpIGV/tENb8VIsg+WzeuyWfqO65WwPrNupF33vpcWq8TMEMGASW4GTFkV
2/1lo8qdg8S/GdEphP8iZYN1U7sIGJgdPrn2mIWxlvboLiVW6EHUA9z8x9Y09cEK+WLYdgtwgD2L
MUoS8/5C6FZeWuVILBG0Slo+TYBkatiaq4/jfES0Ugh9kX3xxH5nF0pHvBl+6I4EeJa3V2EvKkgv
zpS4tPUZe4PjlSXMjdm+1Fap8hXzpyEYYiTHoTe1ICSCtzaYUywnoa3miuEgTKzOQFb0GaQ2UA/o
MJEv38GY1O/tD0zOxpY1N4XEGtCb8YYbF8GIhxn0tl7TIWQgCI9LgdPBGL87Q+q4nYhuQZONns9J
IyJZ+j0zU122SNydNnrILuMUTvrsWhbIa/uRS1ZxJizU8bpc2rMInWdvaBrfAheSPV97V5YN8HAP
jbXiSgwhdLgu18gfitB6FeGNalsFVi4dx9OSNOcIAmdgjbWLSxApRBSdCTrxL0P6yDOAGcBLojYX
+rcexJD9Idw36sfCgzu+h+KyN3IhnWv1GnFFP0zoHBHHZQJpr7PnebqUjgFdmjYz+pu3Elm6VAX9
+OGQnKFehVwCE2cSbcTRyizzWxxqoJKB/25TQK67rlq9tIEuEOn/3wBk0rlaTPq/SgfZdZFA5RqL
YTYrWFy4ID/U1aJw5oBNaMOVWjqZs1unES6EI3pBI5pui3jjG1ga+z7EXhxmIpLuMMe6jiVqxn9S
9AFccOiXJ4uIsqW8R5J/3QSIuKjziPCVgcC/YXK28YCREnXxrM4IFmQzWTdqRyicanv4OhUF9o9g
qgVVUfBnbTHg/DrBgWvb360r8m5wtV4psOwS3CIxDL4RXDlqA7Ztqf56O8YUPvnjKrHhphJ7eQru
YLruOc9ff8wJdF1/e+Ue5A9RxRlP20MPCNX9ECmyzD6GfkICesqhO1u+lNnqj6dpjcfVPfpCl5K+
rtUHo8yHOl6r9LP5sjPnJiqUYp41CRIk8un414Y1ni7lAw//kjv1XvFxarZhCAmTvhuEiFIoNP8Q
LJrijkJP1Oq0wcxsQt+PUNIXd2YIz8OeG5yM2KWx2bWx/jLhk6NSxnExGEpNdxjbL52zf2xruMYf
fGoGdxPplWQRKLpT+z5ugBnAAFyOjwg7b8U12z9KJj464Bkw5O3YbreWu7iZ6ffRYIzVr+4ocQrQ
3px4kSDq6HC6RaJrQ3QHIERxOJuDDpY6ulZVRa3zqwF03gAgF63XrVTzWMdcv59vt9hyGe/q0SNl
cpy8bFXdmkHOcdCUgNOtdfzcANN0gBt4NHCRB3knSJtNctGOzEmtdEqL4wScE8PA9luAKuLvbio+
Sqh+IYrbmsEqgsxAdgR3mNekrV/QP0vAP7iJxiV5mEkcnHZYV2MqOD5gXBggkLHhGvHcRoWhSCwz
Mm/aszkbpAeucKoVyzDsCUzZXja9R6Bmv19rxLiu3EQEf3ffpPU0/JNAebhaisN0CUfYbuE8h1Iy
GoDH6KDmg0USpkZXNwbTg7JHZwZUZir5vUygvgoCLYFLLQMydakChW0PCtP8/p9ex9cHT186fBxR
8wXONoUonH+ceoM6YkmFwn5B0ONivCJskd5lgK0G0+IWFPoayAw1bivp36ya3m68IHa4AJiPQG3e
Et7ileFLTQuROixEHO6b1YoP/FRjC+l0TzG+BDQMXsmzeeIV2ya7wrDYMf7Duk3Y00kUvSSufO7l
8Awo1oMlGEp1uP5WisujMJjhxatJUW95RMStTlcTGDyrp15QH32YQSxVk1M32W5nwnDCLQ+WRdI/
gnHlzPMS36BZYzF7fazszJG5Q0TCOrRLcRzKAS0+bHzPib/h/tj7bjtzwLoZaEY5KCsJt4ocUj17
+Ea6yvpnC2hjp4ddpU/l/z8vRIMQmwohhjT96e0a1UbpLdupLwSVIS8LE4GytJPxvtX3OJCQBHmt
6tKHLrgSZx+jefG4o5dbKLeTZL+U1THubex8GdUDQclySe3LTe1BdB+GUjuKCWdblNdEFqmz3Yj/
cQgDWw4MquK9dJ9Cg9U+3FlSfofWRLp666j0y/S9hqi1U6H9/U4WGo56MGDISI9/FIqJYmUwX3wd
QT1p8TR5ICkeHTLAspZQ5FwfB1d2J9hae/3w1LjttqjSiDX9YYKbFhLYPp/+SCURPSYz2FeZ9T5Y
0c7C/g99JJDf9aovRdKF+bvjMXj0kDbwIope4AEcRx1oTrq5PDAa2lmrvyEgc65QbjIdX6O25xgJ
zQjMcMMffdGN+biBSUf92Ct3kAXo1yoB0ZiX9qyZc+Scj1ag3RkEuQq7kpRKzSC2/pDZxpSnLqFD
4So7lTtRcpGogo5WXBNVKDCfTDtpmghdfxs+ldBFutFF6nL4yOC6wbJCI7azE9tOqKIX5o7zcXwV
7J537kgpYQJJNEXzAPNHiH9YHui5LMrOUY5705AsP3DNBirv+s+Dc00KD5NqQEC0dhiFd6J/YAC/
HYgKigXcZiGpziXu0o03OQCVlhBcHacS8Tao6v3nCR8aZU/sr/3tiqhF0xGwCwA9IrvT2ut7dss5
geoxv+BKobLti3NlE9WJpOpkXBI8GoH5hT63Jbgp4IvzVRc5VFjgw2EnDOapRqkyoxOMfuIxzJD+
R9oVmHE/lHb8XUN/WkIOlVWgjEkmzSXvUALLD/FaYPN6DDY028PYjtBBd4e/bLww4qNcqv2wX3vv
Ll+DCbRrNzsix0sZIkoEPEaypUlvM9rlTcN9OK6p1oafuPSbnc4heKxO7DfVdTK/HS6WcTYg7jhm
u16pLJXqw1jyYWqrTXvKuYMnl+1HRl6RIMt8x8hJECNhn2k+QC6G6R/b54ncB/ztj/jn7DugP7cO
9099IYRaFGwgxODmW2JtVHYdvg6YI8t9U2lHjDYxekX4OZHlkXszM0lRVhDRPo4xi3A0PM94h3Yf
1b6WAS5GFr6OaOl8GlL7mszjUQZBacKdNTmhZuVU1ARbMohPqSPADjHgMLNSQmo3OuJsj2vSviea
Eu1/namrIxwT9Jv4zt+WG/19UrqRZ6RtESrbOPXVSDHYll/7c8E25hZCmBW5xuNa/dhXWLjO3E50
kZDYazGsLdzFnkA1p0e9URSUlXL0ehnyJ9FWnpV1op5bSkJzGKfZfEKguo7KyxCLDcsZVbBTx8qD
AOucCtD4QMttZFrYyYL5DEDoRQtOD950Tx5v76Dw2oA8Lu2R0y7ffmm+ptBu+Bm4gHNxO3Fh+9Q8
L57H+bKBIDxyq0GZzEocI0TVE/4bMVFZDLtfMrah0wB4awPbB7P9qsqzMccc1uz/2/nPby6g6oo1
HU6wkNAR6lZ/rWhmuOK1aG8vXMPc5hSPu6JQSUl2Hmt7JUd35xtVXUbzJkIQ+zAPszEx7jdCP4jz
O5su4Dgy3IC3yTtn7upb3J8kouNLtNcIIyGdZbLFaeWDcRJz95zjQvJDc5OYwGvHWVpf5z5j93Kq
QDYjEA5A2fj8hEETSUUxBQkcma65nYfL/uWbjvfmc5Bw25UHFynX5H6R49fS7OU3l/r/ZnoKcXvT
B3C7ti8Fpar83Gk4uJlrSOi8joeOXswYf+zOx4QGP3VVBivf+sfQ8OaqYA4qR/ySRgwq5MNXK7lz
OrTsiaqw94qfhYwTnhQQmrTGedNfV6VWCBb6A6rUOMvrXzTw0EstyF99ZHauZ4TXKZDAq2tOXQUx
9/pkUaZ0mE8xsIBkQUzFCznp0ZkmcIP53VaTlqv5orTtrDTjGB7DdQYmU5YQVcvSbZTXkUJ9PHh5
RzyHCfhiqOCCXukGEsU9y75zgno6EpAHjmVxoeTgsfcXMoblXgrY6L7dAglErTn59p5k2Qe4rUV7
a94VmyrDpz8KnPaDh+pY+Y/9O5E+Oc9VfHjIbVgA99Gi2Dx8d7jKXRNUhs6F7Nqvv7ufPGVz22vQ
QYyHrWP+9Vp+QZT5bvlVG29zHQVCJX6Vcjc75Lxq523kHRbngPT0MYxMdy87c3I2l8ePBWy43f/N
hSo29EC9nBeX+PZ3f8hJRO2YSvI5o1CUTozYtB7d4Stjcf0YwCgOyskKfpXLsOyolxxvDp5w611h
radQF2POi4xdEtAnBo9pvgN5CWIqNgxKSohRekGAxkKMObU/CtkoesgmNA9FU+dPOjiKat1+QTge
ExnIIC3en1b2Ddc4uhGZiQSQGKjMBTFFmq5kifRmlVOsGv3LdQQLm7gI6FWsWpoBLx/wS4NHXfLS
IFBlaaBVv75OI/BXBP3jruDgE2Scuym8haI2NXJmZYOoWXis9ge26ky1wt0o2wWy/7wLYTg/5vD6
VUkP3FAq3RlaDehsZcsx3beV+4o7T/wE91bmj4iFDT0byKb+3IUI9D/WL1dDjMELovlyIL2XqyxN
85d7ta9ODVGJ9cG0yp3Nu4aGeT1OoQwI+jIZAirJIQuoWG0uiOUDQBhbR9elWEjQOhaEwRbhbtda
GvRIwMCJOQpMwUTjOk+B0h51J/Wos3ehzwUY3ZjOzUErrxwH9qymwwEoUBxGJh7bCMc7ZN2ELme8
Rg0kLfEgQ7LTVUaH8e+PNpsaNkgzXc0VPuK0m7kINYWUMWj8l8+PqtQW7M5M/kAv9sx0NsjWGCVb
u4Lzp3YMCgfdu63y3tG5Pk7Q+0WeRji6MIEQUuVUARoV7lE9X/UgQKYCTyBO6DDfjS5NUNdsasUu
rUvHai+4i7vdOhOT5uO+7gJJUIgfPAjQTMkAhrc9LRZiHno+utebsUaKK0ppKMCtGGKPnxIICQJy
JUeoGXwpwnTVc7YFU6wQY01MqtoOZHhgUjwBNRWwgFYzj0qdyvw0GJO3vuFkOGWGKWRiGTI8JSC0
guTQ6IsFnRDJQW8X9xSe7Piqvbc6v197nJg7+d07CRL394QUaSCWKqYQokekhxROEiVHaWHYLtE2
GxV4qKRJvpEvlrencTyZ7cMF4FnoFZ+HZ5nut1LZ7wL9HgPalmUXouoYuciR/cuoKQbVZGOwPc9f
yx1I86ZMneUrYur3EIbaDeAAjeabjcFSfuhRahnbc91/BmfH0Zj1MLhWDDrx13k8ei9XzWL2mawI
Fbv/OZM7c1FtIScAxklw6KrXawtIIAzflOH+6LloLeNdSldFc/5AeZdsQk5yG7H5rmPFWkCti1tW
l70U+8+BiujBKXbY98aQLrUdnDTsdLOWnXC1pggiykpQKgBIm/dspl/1nuNAhFTAGmyOOcUNcgST
PZQU3u9Cc2fKVx/TXMTYyUOzNKOK/AVavhFTwG32dmebNJd57zsG9O7HyAAQz0YhIZ8kGlN0r9U2
+/iqrC5HR2Uo3rcUk8bPB4VBQV/rAo8QLZSxOEWEQtze29DO0ujNwlp62lV4RAypi7N17dkE8vC0
9U+zjwZWqs28d0nLFLpLdFDhe+r2q0XOPKixYPrM0rEp0Lv0Zp/jE01ANzimhvzxdPVBPqLjLia1
Q6sr8hbizryL3X0K+vV+LKJlGCG6eDR3t8Jh3h/pzSCSV/A4bM0XsfEkm2lBORbHnDOWaIjZCmgt
l/C4F6tdHAxS41sSLi6hSfPs7Y7xIbD1XC6ruB1ML82XKg4Pw2m8TyASpLJzBY91KYtgytZD6aan
Gpn8KH5XTQaPe6DByhBjmHAwzU5kJ9ZE5nkY+GKTaSGaNi72B02JOEypDLVqn8Zl5W+LaIIOKk2S
8w7Q/4pOF2VLXuKrflzHnEQxBtgoueolcG444z9jT7Tmqgmp5ej9XiW5npEDtBmVWIYpRYqJlD23
OHcHjcjkTCExp1Spu2l44rJ9l9eGhJ3nD1fWiodb9cUw0y5UCHIuEF+4BT/nsfukcdw3YTO5ax3C
muVdcdgD5raQaSGjhDOfWpHq6igTTpWJ19+092QQk9/U4TfqgtdvmzQADkGG/Ddd3GaMVS96wd9T
UzhgVR8axrzarXxUJPZBgNOqWuMEW8s6SbiPRxkeO7tBX5mxbWDdsPkBSMNpna1gDYqBAFZrrIPh
RyiNXk+sy+uwsQYtVjrhfvfvMsL+/sGOt2V/V7S+7W4bUetmWcVjxKRsMNyzilU/11w+sr3EKIJa
uFZQ2xQxT73Ik6+ZNh1Vm/wxWtRUY1dYOl3PN5XPRmwM/4VUPtzT2UU7ukRqvJIUUX13WeEWuwx2
HdKFLzGX0gN9X0hQwj6o72uEQ9t6nINrjmrV2b/6ztszb2EVuDZzHbP4wD5HSOeyxRVnAD0C54vo
tm548BGChh1IiZUNFEULM9ByOf03R2ADATVHarhft2tAYoZKczgc6NtOHrBVsuk/AgR0C9eRBmvT
b2Y+BfJFwpcWQF+zuX09gTub97ucX2vdQGZnxndZuZrIOb10I1nhAZ/+AFjvlHHvFW+8Yc8txssc
49gTc6Y86FQ2z52cmzN0WfqUKilEAUtUBFebFadty4ZtfI5PaFi69erTl6JLJKYZNl47CEAV/+VS
85I7cQbhAPtZcpH5chTdE6PgTIc/fBUVa7Z0a0GVdRIfBmnEGSUYOUtmhARj2nHpOzvaQ9ppQQuT
3vsxcKMXujLOv/XBX9umZoccWry2Vlqz8z72aXxPTdIyWmY7gcA6fDX1rMIm1J3DOc2spWqKVDuz
cWyqCq9JyTxRr7q1ZmytUZ9vykbOeny4JggdTEa0OH70Ge1iGkufPciiX2494tVfBftvV3KmVICX
G6zYyv73x2AvF2165xdM24DaPryAOv4hwceEtEC274RxCEEqUbztL5aAkRX4E9J7+PL5YECqQiGW
RvBy8WaqP2clWo8YSciPQ7eHI/adZWJm3DWGxJaggNaRzfJuPyFkhrGIGoYcD+GFIokDFsTDX5IK
Xt19vFv8evMCpR/dIN3y0mEOY70u8k9xs4HrSnIIqK5KX5EsXjVCiLfzPNBAVxppXw053K21tvjX
aqf+ocdKUZzLzEJBhnB6gwPJjX8jMlsMMmeevEtmY9rknd9db0ya9DW29OqfTTndZdVBxBz/5yvz
L/7gUHcSP8qH14jhM6jKS9XTEN/OEhngH4oCLPwlJXf+3Ki1HRAdJ8XZlkuo60DWuSPVXBVs4D+/
Okbtsd5A+Nf62YW2nJf8ATyT/7hChXZYlmz6Ej4qCCz7niOGNMOXnxjCpW5bGxIR431dpNPj24Kz
pqupuF6OqHFKw7SS/MHg5ibwja+mkrd//ylbxSJatDjXev5kME4UeS61TYpqmRR/aX6YMd2uXkxK
R+BJuE6Phr+srRF4LBBxQQ+isFbpJh6SnPlKsM1TJi+NQHHao+QiPzhjqIWtsIsdDfa8Kuqq7dHc
1b6qso8gzV41LeE8yCDwR4trmO/C0tgvbwQKTRXhfeZ3UAqPmjZ6uF3XsO1HlQaNsOM1CQ2kOnyD
wYIRiQVcoohSe1tg463RxbXKeS/c3TzkijVef96z0urLUN7tCA/ohn0rsMTAkFPOIJnT1EVuQJ25
typnGAqMX0MuZOfAjNIIASaLycueKbVw2Vh46Q+MlFEQKEVcOio5n+OOwlw+Z1tBs7J+gFL4PAQL
AJMcC7bkgwkCL9Psq9x71ToOgWxrXYEtZXLTnGonqUFdiXF3rNQQ2O/8Yt51T89A9kFnWpt68oB6
Vo8wsgh+LEtRbDmvKsEmnJ6o5gSCGRa0czajKyiOtOLgm7yTTJi07W8Pf5PN4Et7ubFzXEEOsySb
J/SbN3O+JtdWcxA+/hdwYjW8uv7W9r8OU6uLMZwAmEc/tLOZe7MpVd1UPZs2cmzndfTYjweeeoz1
Dy11/ekGb7wLQhjWWttuE2m3hxA/Z1vjQwvYr39rVoB47e5gu4tKZddrQBHTafwVDnt0jeZ924M3
tYkweLv9rAQVPsc+7YCvJzkhnMJ2GwyI8GvcESIVqW/zWBEDTZjymos0IQCbUgCitV0VGlOFq/T2
oj6z+no8yUVTisha5gYoPn+XdPMv4Lc6/yLWiWjwDltT/lTDZ68mufWXZxV7ogVbVPdKFVNsMzQF
JJagcOBl3sCOtQ0cBv/ZeCkWov3hstWJPI8GA9BymTDKz/yFYkrqxpvxebFTgDO22F/Ez7ciYdOm
VwK/GSEevyeYQt2Zec5kgKfM/ycTVs5kYBkDQXKaJrybAFGLd/re+hMqQuTkl6x5qgPXIzwGzhiq
5KHxzw6qNP3NAbg4Fdh3tCg9NUQZtr7WK1/iilpU+QeHqhaVl2swu5cIyXC/4nPkvilvVy1JlPiP
+BNRbmR3De/B/+f3ebaukKMSbMyKA/yy3JD6wPPiotOCxbXoGki6bktoiqIlPxbH+JN/aLBmB5UJ
GPGLTvPUQjOtzGlOrJpp8ovVDD5JfdHnfkP8BsrYMJSY582zeX05JYq1x0J0H9MpNuDMgW24TLaq
9F/aYCNfPfTQ0/v13SEeFP8598DEfHWvddbgJkbV7Oqwo7+xD7kTzX1MMmZzeM5n4CZhN+m/ts4H
77dIfFCPPzpWDy7vx3RNg/z9fBtFUYREeKMYPg0mPwBvbhubu7npnCIlbX3F4VWD1qqLg7DrqAb6
UlPdZY3BE4373bJLkEz9BDV3AFPN5Yn9AyZSW2OlFxY56EuCJR9A6kDjDIvuJhd6w0Shl/UaBICO
XAIO7AxX8sJf0Vd7aRIscEQZkhYtBkY6q9gcdhtbE9RS9DoyhV5E62VfVr2y4pSjcO4mtzrueUhY
v2ae3kuI1vIeWB7DfW8UcGDul/ZPvD7hijgjv9l0VLHx4mRsZ8nD9zEAzDseAxdbld4nh3DYvTfA
Gbxr2xqMMlpVx/Wx14JbSApf5U2ZfMZ63qWySG7qTxAIzLHRfebGQE+z5rw7XAO026Eu0xOGkW/k
F7qgJNSJYMTxUP4zTxWiB0q2GmUvpvAn6+F/HRuqkrXqHrZ/nPKMC635ERl6vMYW9pRMh3DHbjSm
4qSsU3m0SHBHQ1xdKzEIu6v6zPJmvErpULJ3+16uDz8Jn6amgOD0dB7dOuVOpqnA3vxvuVk/E/7Q
5SJ8vVlEgZeCs9CXpN1yQgIPa9j9Sn5eWkVT5uR3fuhlGwBwPHxp1bjgl6S6aNYeVCe3UTZw8Be0
teBJ3anqigmZ4dis26O/re5WSoUyH4Le6Y5k2Gol35a14TgY7cE3KnihlXFpzRUI9DhT67+ifoKO
rpTHl56iiBpn3cNbTozxa6YffuDeDjTkrCAvBk7p9NCEPcn5pqjPKYgEzaWdJirCzaqhYuLMjYMA
tGpGYWkfWlrINFMReELdQUIj/aATrh0gjK9cJBqyOugpJadTMYeJOSS9kKKYSMyg1+62LxSzkGDz
teJR4+j6Ilron3kmNA7my4DfPklxcno3gImV5gsV7rQ6BENAuwwu6LfHlfgvyUzdboJZ8xDczoHz
G5ex6HtY8aDiZzcBi5Sxqb8vSEt/nnclKqmMK69x1zS/f1VzV+VbRSIDF77NFcANVECWbzaCPeSf
fB1f7mLTCq6TSxPzJHk5hoL0FpMduvucBGYmrw2mFyFbdzBcfo1nDYC2GO1YfSUqHJbXZdu8S6Lc
9qB9uz4mF0v7Nxp5eCqpAM2UvYka2fITOMINCMC4HyyDowBxAM6TE1nPfIPLbRKgB3dpDEdATwMy
uZ0i9rSujaWnhbU5GOFpkUTU8nMZrcKy21PAz0rz+OJXKls6DeU4WpoEYp0ybsL/Ok4yFvDVQlQd
RdwkCmJpX+BbNPi3J/8RuZLjO/oIVGx0UCzrfm/GqwKcCkXEmlrFEX/Gy2t5SpGoum8V4wajuBqn
wVmysBT7aA30nRTi4F8vQyuPAYbZQyHYPMTcrHWlfpz0zcczhmJNB+ZUDAq4cdT4r/ZeEvfZJBNj
OnS9q3aNmHKi0QP6/lyiSzk7r5goHsiiNRjjk6fvUjmYIuesp+YjgQAtxx2rTH4RiGzIvlSH1Fmw
TWFzu14k+Pd9iP9lETu0lL5fAtfbwkwk86Yw8AVF3dn1yy5ZD4LGd0QJYEdBSDZlgHXRCEDRlRPE
M2keAoQ0nhPE4/RO3aGgqKfM8QlB8RXhvKxBj5I/gBs8/zU7l4fSFhxhYjj4D01vHjCINcuG36bQ
qrhebEkOx2tJbxrVt9V70zI4fQ73zAghb8okTov+QjaNOXgM2t9SmnVvwGXlzuvgAGxnBt0VWSQ3
NvBDbfFmcnPRRNIVFcXDBpkTs9ejuHslEjtYQxmPposbLoHOm76dVilFxWwZJ07VcVAitTmvAGLD
1G+JH1w4B+TjJ6VNN+caOmBemkBM52b8QzDby7mLKPL1is4zAgyfckB8jxzyF550lmd+amm50NJI
LAgTorYiDQ47NV/gq8VwqJ9KBkxE5l6J5fud5ybpzOj8VrGR6cA5n892Un8EEtcgeGm8AQ1r9ACZ
bk9DvxXabuvOr4m3fdgctmTZB24Fv+6M9U4zSV+LwjnbTg+gj0MJDBOyEuq8YjmbFt2M3xn+AlnZ
Yh8c4C8570Ru3fz88rPZ8+CkIu7+d04VOzqQkIVUFMdriWIb5gSAj5TZwkSguy8OiDFHyZYSek8c
/C3ECgkT5465OWwLUDGs+WvIOmBSgu43N766FAGZSxrg4Q4+8pC4SMuW4pBhLaYQhn19tqMoDeBI
52XGwi0ulPP9Wff+0jI4+VVSB4pOaevpoMrxOhtXhdPoHKfB2qhv3T9XGGjmb3uj++sFqsoCKEKN
obNFMs0oacssMiSLrUOq3IBd9NIeSMMK1/y8ut5NyLMuJZuHZHeFJExQv3E3icHMG6n/AdCBOLDj
akr0JP38xSIP99eZgShHsnnDORUrrtDce/f182j7k/PEpmGVJsWCmkTZNqIpBe6YtcoThED4fr4J
qYhKviGXd/JTsH9+YbtXfJTP8uzP7a2XrUOh7JzjdHDhSWd70Az572rdZ/DcaNNxJuZlI/l1xTqd
DCw+M5Z+yviCqL1c5One2mMOhz0sxMIAE1VxL9tEmeF0ivAWKCncxobyZlKZdYu57j3UEDyKj53z
hGCPZl9NLVhaeuT0Bj+EZV+W/wQImxWPEBvM5wOeEg0ObesRBtjTtOmbrEi2ePFAz0IX/hoK8qKQ
ZEcUQqumvdszRBN6sSdaNAOQzyvwVegIHT0LTa+SAFARYTgFZJEPPjdEJOHho3npE4Md/FboDIBB
a1CmKdPgMtxCs9LoDUnEvcVxtylPcLaN0qWf27xuEhjrpPQdVWf0q+6kaojF+pCWaZsp77Z7BdSc
8dcKAxJfuV8dxrWlmdIT0eLrrnlr50JYLHagAq0aPt3BH1Z2fc8Xi1o/so5B777N4o8XDesFhb5S
TEglmZyPV+T1tg8yaddvcLq10qWQqmLaiGQES5nWSTmekOdGcw9xY2p7Phc8Ua5Bd5AMU6HTMfKY
1uWIskx1bjXDJfYWtiIKx2k5f6RSCvhgxC03zCAxHU9VhFLlVPU9BmrB3n3ALayBtwx2xdtBFF7Y
7qnKvLJt0zP84cUJx0QNFfIRAUgwCFiz4pB7jIPL44rQne/AjoNLjyFnefmlPvZn/rZw7l7qSLao
f6qDwOIt/Pa8wZiJXZINxHeF4pnynJxmRfM4IODRMRaIcfArRAfecfgu+T/V2y8+inNJcHwn0Eqm
tUQ5rB4eFDJ9jdvTtp/GjqCHRtvaZZhMKqgA3nQdG5RofrJXTKYpH42p631cLiW2uDHWnaHYFU27
SvLsyvdb/N4lmOkgwB7GG1yTO2iASW30YDF2xREKAQYNNDmohBAKt30DN1Y5PPVumUVAab9k/kpn
k65Q9bDfFEkkzgpIf0mwNx5Ne0Y4xzNTAXLxHUYsug+YTulWpnY9PIPsEJwI1wAF31iX/8eSJ5Qq
HjjrDgFJ5J0WacrDOrXf837C1+MhjI4gF4aWtYDzBIt116yprjKiU+7sSMNdI9p5XXsaucjMxLuu
+u4nBHggZ682dr8dKYS7nhTSCM0bv3TUWHzeX/0XD4pDEcjUjZdecgro2MZPkz56ep87K4ycJBxn
HKlGMdvutF1sUyovZ5o3eo6KvSmQpYuHRfqGG+nkuncBSAIS+dO5GRrNlUJjkf0rvlglij6BAbSN
yyYNAllN11nI+QyMu+D66V5c0VE8JxZhOcLAC4oTUe5CIUqVwS3f79xvS5cGe2sXUhgKufbgkize
1HZG6JCvKX6RivZubMcR/ueKSEjGDv73Cel3ZrdaA5fLTMBT9tAg9fp6ja/7lxt2GDvlZGr64VuD
ckf+6ExU1PIx9b6aupFSASxlnrgyvRRfVA7384GVfKx4+AYdPe+cnnjugQ2ML39uvnal62l3ZDYr
Pwb+L1Qtb3hakR+Ct2BhCALKu51yMrzwI2JIrasTT4T0EXr/z4SdFgJoRbkCZDpqh8pzC4jlEq0H
N5rK23nX59QHL4Vf13wK5GuEfeaUo7aMzaTv7+3I2tip3CFeDPave+l8MdVEGUwSJPgZtKJOK091
cakwt54MXyN6MVFHdII/a0258WF8Z+9h7ZdpnC89bR/DUcO4U2FCxf+2A6o3/TjJMxGmRx0ExlGO
K5apLrO7gGdaGWcbuPd0bYwbQ4pWB/F1dZrM5gVl5zRk0jQHLT8wbGCMKb3AGrAcxvmNPqOBnsJA
tDR9vdP+BR7dJfYFW1CwsV2+Hx2CWmz6il4TPLoix0vkIlvohvJHu+NYKb4uUysEg+OLNldvOfln
qTPCRHrZ/UEvk3QrxLruw9icieA2Ly3T2MW+NpY8LYOrH9PVF9iO8c4dfaBziqzG1atkYSq0xlI7
zs/R+5/Nj0/Uk8T2+6/KkyNbwE4uBo81yueI+oGhXxcIEsqmJMO75loMfLlqkpQKfNCbnQqDqjz6
++NdzmOIOVzp6VE34O4Z5GCo1AHcqV09EQDsQMiIn8RyHV5p4dZbY4i+zgpekBVJ0U1DLjdvhNkh
cHPCAZ5/rwqrJHD3JrBDUdEUjeOKpHlb6svBWYItKu7cloPA/W3JAa/LDHgODuL2LsO3pezWak4j
yrquJ4tktRAcBQHskOoqSxRCXPE8ZObXUlAk1bVlKh6wQVTWeqLvbWiYuCgcN+CCIXasbqPC4/zA
1RM+eHjmp6jWaqG7fQGTaJXH8fvga6axxieCC7VQ86ho7A/0Zo9KviUVp0pkj6i+KQUNBs2X3N2A
9JTcAeHQ2UpVOzoHSYgJtOfqriDL7BJqpnePcVHqsnFuTZ7m64BS6/k/TVsSL+W2lS2SpL9BZAlb
lgE+Z6U2oaUzMQEMdPSybfflpfNVqwnzpC6hJm6xIFcj4go8GjIsmDkTl2jTHtBiUFr96WqRGvO4
ojPUURjln9lV0PcpxZIeGxIqKehz3avbgQKg6twTMgZhrE/TMkQjH9n3CiHhbNKPc/xpsRpor37I
R2XPaLspEJIz3moDZTAnaxEKLrglpCa3Z5BtQ+UJ2j93yVNS6irN0EJtSJukUxEdajJb9Z2MSQiT
DNb81oJ9yyaW30b6NEVuCn49TgJRA7Wb+Jx6dGdlku0/flcBz4cdjs8M+ZlS81KU2KxpwcKLCdaO
m+OHmu/9dYZVPj4xGK1jZpETqjSz+vyY1eOppPil4Er6vG8ChpnEqgG0bfcAD4qEBQsDXE7eez3d
dHURDe1shdlNAv6det6aosCCQ8Um+KbyNRkOF0c4YRPZ/THL3h/GFThjzOA57xXQrjZOXsCE2waY
Qtx4lIBdrLisMbKnbmdPyeTTvMLeHb27Tio1S82njA2NgHmQ694U91H5klFwKCwJNi/WQpwb3t5/
+3qnKWIxcQp0Q4rGk3CrSj60V+sfh58uq6LEArEsOoYCiU+5ZMxXuL4uITxSEx2HrsUkVYaiKPK/
m0u59flZtut7fpe9N1k8+BtbDbjaog8kIv9QmZ/bxDclugGp443AEPgkVE2cHLoVz0ISF3T/2XQ3
xlKWYpZyJSKc0vMIUmxILWvq9sCwry+w9oxCNpT8ZWCmElfZDWweE7b6yDXLsH9g6YahAC71vPK7
Si39Mg0UHegfZt81en67RSCG2M4jiLeKElSziePJgomkWWSVNPn5O4kUEfG0cn5rl4ug3C1+F1Iz
EoDxEKKOMOJFdtAvNsmn+7KpHeafNyULFS7Ee+sJgVbCtNurmJBrNyHS6QXRfUFjWWMHeuHclDUU
FL6SeOxIgjhwzuFD8uO8D69Q8xqVEUjYpF89vWYo4oQDONcCRPRd/XcyCQ34/Ja3S6buniCiGSKu
BLMDspRHnJO13nI3o1MtouhaPU+LWEMWcUtD3VTeKUC3PYqNF9UOzNUZ0jcDN1BW4m5IRCn4MR1W
6CO7nnMFyafGLi51uD+E8MTNZeB6rs1rG3ZcEyL5sYOLBrNp6YxOKlUeo7oAvdeUt85XBlnmDA8+
yeyfDr6w7+hQm6l2NoNISPOcu8V/vpxNWjkWjm4taQWV9XBuOs/o7/UH/jzrpVAMIEuyMTXPP75v
+L0v7NLSM/mDZP/ZTVkYtKCRxQGXUv9dPyaqtNvdD0FlOCFg7ggSmrNnT29ecO1gBo/+DWGmJmZ3
cgHDTi+cbwo3b1upqCKfLYu+TDE58POJWvdN4aeVujUyPXjV+4ZHgWoP94zJ2P2YkFzcdRQbgv1r
STXdnwT/rpm4dYxr0JMePtcxGa9G4/w5faGUocfLk3MdyTv8Jm1J9ZE7stQRLRebulQNEUnliU9i
JZU9iL6b0Jx2nJKwbML7HmmuxGOLtNP5YocXVCA72UYYhmwwvsuHwNaV/DrDHy606AeMgcOea/e0
z5/j6T4rT4UrowWNw42/qJzqeV7H5rOXeT9oJ3ftLcP3NfEyeopsxwmlTBOBqteZ/xd+mpznvJq4
vZ8MLvxcIY4YrfHlZ/cavhqr5QNiRYCZ/mbV2aVbz7cFWSx8hLtIp0xV1mNC27Abd0gHdXGWmrlc
iNmDhXyhvaNr2Rvj30j7iaNZvzDb/Pb6GVrcGMmzW1aE84e4qEVx83iLHknJBxGfxwkKjzJHFK1y
pwrqm6XyNrgVbe8X80d9fOMe+CKtXoqFAiKLKCcIwxyaB7rxJ1m59m1RTuEWSJYHQmusAKyMD7bM
HND4qWcJBmsXO9tKOIdqcmfiIYOuQ70F5PDv3fN8vjkNcrZ2RBv9Q3mk2GBACrPKw2sceE8aybH4
ArbIIVNt2pb3Z0NoxHi7NJItrBIWhZhPPYvGhHsk2SOU4b65CqO3IY+TBaL+j5KHEG057huB8tfq
FbpSVdT4F2s3IYteXSUfKtR+JKQONRtIKHUMi2aHdom/mj+J+2gnBwGOhS2Lymvi7gihpzcio3Be
3bQoW5sJhLBMmlnBoTYreEauIewYS9BsXuf8Eh/wApVTPv3ds6fEgMrsaurkVPdQMX/R1pckuTwb
sP7KZoT+55aaesnR6Ge2HLNjuLrtk4P0CwFBu41fAxBkIGLan3reU2N34cWOVcWFPWlXfc2gP3wP
JWkrjJ30kRvKSbCpBTmuNttRkEJ+nrcLvy2bOPrxW0jwcVIaDTKwS947N3rYm3Y0c7iTKCGWCLw+
Xs66oMb54hejbecbuMF4mYGqMpOAZQtStizUIzie9ZWQUeRu1xLqmlVMdGbgG+ekStX7Da4AyLjU
sk44NaUtjtGbBXywosWqR0iCBdUWY7+k2ZVPUbjRCv6kcr4WG0U0qAW8XtxIQGvSTpKYJ9Ww04DK
PJWmdY4AYBf169IRBEZFF0hx9RrrZPiH3lRsMjEbosnxXCplfesmHcmFYQKQh4yXjv8zyuKl6bu0
tP+h3znzcWhpZaw2p38zh0OrQmkc9d1fHYmUacrV2VlCYXUFJ1EXzxAxRViHhmmxFWA1ft1C0Rj2
Q6ZoxLyMBmsnnpYQftTqEKmCkOIxp8Uh/HRRlXbiHTirmE6og3VQCftK/+/iXep/VZj3W97nzwzY
fBAmIZZpaP6Liu/z2saDYbzdbtzXXFyW+ux6fP/tQKcj41kKeP+VM+jt7v6fLGJhwZa7OCama09+
zn73UUBUVmnNoNOodgE9zue9ubUyc1xlSy3N5Wq/Q1jJSkItB6GagPhIhPlYFz1EB+xMmSAy9Xwf
QV7Qqb2nnfmVXMTv6nS7zxSci+Wdm4lCsVAfyYbqYkNpBpl8lT5x7y8bAIvmR1Jz8uTIy/ZyIMIi
88iPPAcIrDIQlvEWHUtxaKl0B/718L+/+cVAWuQlwM7ce06INwRD+VxWfLIn6wuoCRkINkx3Gqrp
8Tu0V0yMG00Fn6cMab8h/MDLZod6FGR7Zk8PFK6wMVKkK54PDcUmD26cV9RkrUpSt1U3OK+XA3aR
rpcfqpL5XGR8nJXlEBFLKwn8Zzf5QQXjbLbUz3fbq9isfwPcVoqqb3efKbT4Sdn3ddxQXZobye62
fs9ynWj1ZlCRz7w30ruRy4IeBMgEpCvCQIjhLhiPd/Q8m6SjMykfKGU374Nhcmq/js3Vk2k6zJxn
WlOsJrM1s7he3/EnOll6XCI9HVRFHvheXXJz/SFWTn6NRls5kZCI0Bd3teSdK4gNb6IhRC2crj+a
RjXYmYB7dsZUoOx3kfkYGLQR2Px86OPXYB8gDBI2SbsNfj6xIQtPqmMBxyZ6b8EJTtMOrCj/K3td
cvC3PGte30HG5RvOnjSm6ImJrIS9/VmSOQGJSyW5VAGDzsPTGlWy9hDcNAACEM1Dm2zSG0FxIhOS
FHPwMl2s5LQtd04aOzdHTgfT+B8FBwFygTkMSDUiELohnXMvNXylB/UM9JC7v9OwYg0prkz6tWVu
R7Txc5qYICI9hH6RPsRGHmm3kd/ytfpnG5ut1pdZ16EP/KivTZ136F5rklp0ZQR+MsGWy9wvAFCh
0ZBOlk0hYL5oRp9vB+uonhg4GsE9ZjFPPi1O2a+IrXbYL6UtMBK4RRHaIlONUvzlpJScR0faNkcD
TRyB/ZtQlQUtGnmoLMpMPFex26ZSP4XsAYpkcWZF6GzlxrYhRHjw78Y4Xh6h+NT9yNfMiYB7Sj6b
kliRopzdyk0FjfVIdaZZQzL1xHjhUQpvDkK89ZDE5JwY/hTX83leIAdx8BThj0NyjDZNtJBIE7so
esQ5V9Obm6SzXiVZrrbTgn7EqbzIRLi9mKb92VVD+VPYjqt2N6MMJFjjcCLjRh1ixlBbI5i2FYYV
qVBe4Jjw9mB3Jdtxf34lQzMtFWVjd/nTc8PaofvQ6Fqzyq3amU41+J0BEg08u3gBT5caTesXo6+X
QVR353/Jgvpg9R7HltSb+IYDNoB/zk0yqfqaTIjRr9yEqu80pvOovCeHVCNoFlIk+U7xMZ1XC++m
LXWzzqkRI0Ue/9w8D/Ux964emVYGIqLSH01Ygq4tvbWsfsFRctNCpGG84N7vLKULkC7hFC1kZ+7Q
bodknIGW5hqwRedsHrXvdklrsjb8KRjl0DKt7U5RF4LUx/IKbXZfFw19kxoop37VWRJdaVAXCYrW
BwikJeet3rQViUTpAZQ+6HNeF1lHO2JxOhisInQSXtkvIuGlQwgnzgpeRUr/RCm9jp9bo4uqiYRz
WxKbaGpDtBaChAsS09gowfw7xqD+lOfYevtxO6id8TLwk3gUjve/EZ7oRFRKZ7ZbFYsc+I5PhyAh
QPK6cW14rVfDO8azEvu4QNRk8ONF2+BVbxhREzU+OJU+og5ssNHHPwYx4YJdc2yVKGRlw/n+wqRY
myeoOroaP+aMSlpZ+/06B9Hh47Pd6gORhj59tPD6/XEyRSjWvL+ZGUDSKJiE2GZwdNYbpMEFa71N
kZU+tvmfGYz72np/vWxl9fWLyr04huQ9LJC2orIyEdbxNqDUZV5L/380uSQ1dG0AuxjF88Uy77y2
6ZoIlFD3IQBM6WFBJ7GpLQUYkUx1jDwUrExB8rrGmXW7zeEntsgBKpwexzTk3KrrXrDXaWkdZ7OL
Csqod86mFBEff/axeLvN3v/kYdd0uiujZekEW5tc8CfPQKWR2yY4ODCSBtvUOSZXu3g2a0m9Lhlc
KKR4oWO8PxTprJ28K4lrEZVCNBUW3IIlKaUcNNfukAFokLO1I9tSDEotovPHU4yFHbKBaglwewX1
BB2h0QwbC+MdbfJOxDnCN5P9e3q6529AVw2WNI1GQlC47k60NRkTiwKAhTzcslwVMWPsXJBb4JV2
rrgHlYmLe+s2kckDKy4wSXvSw233VLyZ//93u1B8Kl+xOChE7nIL9qprZ1NcqptutDgvmgCEY7Pd
oY6u2KJpiEpmwGl/yd0XPSsS3gUVq9xNNrp3fJ9DBnl9wz12xkSzV2KFKN8XV+yk8GmdGusw5Tmq
YKBz5mmrF4PDaKMwJYhnhymlkea4CmtW5nitryRpw1UuAA0uZfxqwZnyk931aGWZ+vAnNaD5qsPk
ZCr/pszL7TgcEKixsVBA897YA0brKVhhvesVif1UVfNixfp0+640DOw+aCIPXsXziO7BHBUi20kU
7FGKCk86v73nGgSVN1XcWUezwf/P1Dr+kkl4f7cUQPJ5HSbAYFXK18owTgY5aYHSW+PC3MlGbQBi
mU9hsmj3BSIM2OVgX0t6EaoDOjvA4mW5w8xd3HlBpnlDjyVhG5IMbwEt69jYEqIVfVDELrBL6yOj
TGmR59Dl4ovTMHSUtH8tAAh35olhIrCjWA8ymwzee19RTylRkfwp2loMeESrTdAbWgoi/cKBuMWB
uZDkp9g1rN0wBXSdUi3YwuOGWSBiSbLX1kApw3+m0SXi3teEfP+1hbE+L3Ujxn/7E4DBFRHHqJ3n
nV8ELcVIUTdecCnJ8SM7GzFXyFK2GW5H/yL+tvu2O8180E5BttqZVK1YxJy9Yvuvgd256eBkSilj
bv+zReeTyyyQI7l/U0a8p1bx3/IYkjmlSyOagbBa76jZ8uplGOl/kEN2WZMsdj7+AvvPLfYirAIf
jY6miPlXhb2lO9J5V8Od4KBMM9rXWuXA++9IdfU77wb4T/HGZPQpZKXwXfjlaKbAJBVuz9aYH0cJ
b8mYc1rYVMnZUwcGqYpHg3Q68xFdQm8OM8SVHWqgHku8qzyfzIhPh6FnDwzMO0IwPUpn3wlsbgw0
AVpfU7Y27n3TbqxtI6ksAldPIMooR8Y42Jo4aX0MVlTn87YWUpeULpxklYYtMwz2tS3cOkunqWdR
LlgacTCNb3+mypm8N67JVKpiruImLeO8WjXcdEYeip7kC/1ZYiRhusF83vdSEyZG5MQLEkusjuGx
zDzhnNwgZhbtYztfu1QLu5NRdtUNOV37RHbc5dlV+vMphlRP7kTLltwYPWtFCKVr2gtY2stI4Fyn
R935QFBjANXLByapSpGS49WNTDZEDEuIPXHoFuJk4k3jReSZaDcOTUPl5luvXCP/tKYTVHscQMop
IOlbv88BxbXHiI4hLHy7GIlA0wpXOXdOnMUw1bNRUloq4wUG/7LQ5/dOTPoUz2kvkg1t42pjN4Yn
PMT6U3x79duSrGPRPgoqEhEVWwO2GgI/XuGhZDYRQEAx1i9N1Pz2ML56PecYGnvCYKcrycytaJxu
1+/VcU9/JIuuneyVaKk1qFnx4luxvPz/q+1Udu+DE8y/zfvBzeDZzWmulAZELvWf3j88bFatL65F
ZyoqZ4+XebKKrXg2bx6F2FMqJ1GV9Kb8TwDlytsFMvQoXT/ZjXc1epyItQuJjMK/4cRSFxQx8aaX
sqaStyEC96U1rZRSaMFPcPt35N28qSYZjckCDdA8et1+8gs8TcO+lIFkq4KXnww0jcHmEOKXkq4u
q5siHBXTvz3ebs948F4tT9qQlkw3ZtHTTYilHf3oDTLAPkaOM+h26AqZHG/oJZtwjVZFzB68BBIu
rJkVQt26jFGtFKhf/b/YFI39U8+o7eubVYzWLGG6+c7tK2VQfArWVlNjK2RIk/+h+2jYH3r7Pk7z
fI2aaJRUKcN1xzK1Ks/+6mtSWkoH6xTa/BFiqGmpni/LJsFq4RBLPsOTUYzSQQA6437KwShmujNj
3K8lmHAHw44L4X1y1gW+Xa8mYYtlheujJuX+r05T81kk86iZWIHysmIouVa1ajgptkX2sk5+rlWI
yTbfpnhqWXputBzDNKsTY0fl9xJ48hcpGgI8aCP5a3lpSIwYKvhsSYO4h9FvHO2LI/kovUJKRz+o
uw/22XpNyHSs61o2Sja2EQfY4FEHzUJAVwg9L4nm2bGjgivc89ks7CPZoQzdMrGjTK6kjPeoc5V1
QKNw8tVTkkB0yMMrsAtgSMyfFjOEbjHkS9zEybe5I/hoSIEkZUMgavRiGQcEu60Q7DfS+pk1h00G
cZEH6FaPra7A7FZQvSee8ouEzgZBjDIajAAkqur+teru4+CB4pAGhuDTEJ8JGRy8njQZcni3PP8N
T3GGTJJaqHeQrVlQKrwcrJdaR6k4TQ9W9YXRhOybBD0CCQ4yO2TyGGSlTcf63gnlfKCS7Hp1Hc1e
qqEvlAjmCvEsbrj87oDR88J5vuW4soRbyO4qnNaRG6dV2/pSC7i+rzRJrzv9jWkvI2W4L79m7vvt
GjEMdnFbGePGUwcHWUIvwJn9qBiIp4kBf/fg2HVh9JSPHdwRU+PpGyTXnw5g9+TPtcIWYs7Q7kwK
+BwmDMo8Ps2/4z6Su3McO4WPmuziAJzs4FGOzp84Rbj1z3/yq8tCgaCCrr8kkFn9J9W+DvhtZHFt
8wpUZtoAzHd4u8RWKoEBArtv4eNXysqyTJsgRMGU4NOHjZQ3mgtle+wXCEnJgUqmB/d6DfmkzZGu
x+lYEaRm+8Uo6EBWQkLDbCBXLBWekTJ6jcATUaHWSibEcS5i238B+oiSRWO7iiZBiDe1eNycfED9
QbiUeaFxzA0+MV6DlYrFkY92TM6YxtgJPsuzXpR1/l8VqwUxfJTKYSBJxUth+4i5u3YtgmUTz+Ii
ydQe1/Cl601hXYRJDVxKfhCvcpFdL3z02fs6XYiENxAoACfE8eoFVk7u6QgNyaBpRLmR1Mu53e5P
GU2OmsFam6ePzDPAqivZD6q0jvCkGNMmhILGpBrJj8aJSYFxBr8BLlrQ0opB2UQmopB1uSmSupwO
XLm/4LCAJxl0ZXYeIORHuTI0uOO/Hi5Uqtrp/0s4qyjYNPlf6LcQmbadsBvFWbSnmAM97R6z4TkJ
BB4RdECiBSqMPlxQDt9x/HCJbxYlKAz6cYCE5JjAofCjEq2pQd9TVOBmnHw86mfDIqh8qKq9IvGT
xIM7a2BN6h+fttgIbj06YUv0L/d1E0OXMD01F2LtRytFfbxLPa2Coax7+eADO/YEHPLVHWUrxR+4
9iemtGWEJjYMpPrtGXc3meVZJhiRW4vI6pWfHqmN8nqe2B8L49pWX1VUprxO6+tCiIjUR5MLcjfA
fHzHZ0y7ZxCURf6HezjoKSy9R5Newt6nlzIlTzeOMhrxZQgNdrqrN+Up9B44UCPtzCOmdkxiNhhj
VFLiC80xdOCylxqGzNDC1WIbip6dU9HDC/rH9z4LQrs58wcjHQhrFXaMMp8WsEezXn/0qUBjsxWZ
7H9xy7paL+g1pRediXVibTHf24Od/7n+0zYZ3HL2t65+TpIKGqq8bDobNmyhajhwa+riF/Qzxfa+
I//HqS1mWdVuMDecTZmMuWS/igUUZCYsJMFbS/hpf1DQAIzgKgubs00QyF1vCwle0jhD5K1PfnO1
iffnpu5QOQLJHmYZ3zXd3WXmqqjLwtM6pmkCO1Iho6+LSPBztwnCCMrmYjpzqVk5yVdbvltbtLvv
7LuPNxGWpGLdqAn0fZwXlSBDOPhqLdaNgY8aI0mUQi9TtmS6Fu8RkeZ7q0vkIsNJcHTsQJkfKk3Z
oTplPSngYCO5ThedBCCI3Xt6Z9sV/hg3ZkhU/UIoKgHM8qZUx0yiVajK62P3GN9ZIN4zgOxFQOEN
990LlQPv5kgY3EnFwjtXGQzE6Iu5KcZibegrXR4FyuErrgX0Mz+wFgo1DN8GMkLhEpCtErgOVStZ
PtF1zIQbyW2IfAmDDn0vA2o7QsUoTRR2fSKHlukxkwRF0939hKKVPYW+98JqhIGFCnDdmUoWHF3u
YfuZyFuCFrQTyfB7Lzo7FgVHGbaSkc+jTutQWfRK7tf0wtMdrH7xb8jW1tDtN5DCUadiO61T76Nn
RtUcwBQjiIOzZDzPBxpEnb+rsLBsDfGdx7HlmKxShE52ACxiR9HkJA6t1qofdjEF9ZmZrcnXeDvH
hECgAYQd2XJbU20zQAmTjyuyXqnvHwy4ZzPzuHfNfHMF5z96665JtHEn8FBB9aB/AJK4TTLJuKW5
k/O79bD+UuXsmJy9p6KeeiY5bGsmnrIQvaUqyczZaDWgr4QYEOHvi88tVGOn9Vi61xbUXGt4yQS/
AWP4RvXBpX1kcZFnzL+cML2mwE7X7lZjE6E6/ZmBJgNh2i3ecX3/lVQRCfOfn1VU2ofbIVg8Cofb
p6+YJAX7lwYCKAJGBN/VYHkafwZH2eHI65HhrhPAdxBxezrlSex2oZIGF8Ipkgs7PBuJ6RFCxPUv
/CN+PazyxmRFsGzP8c2z1dJPgsLCqQEXgUic5WrDTHAf/U4IqZ6ztREb4fBl0GApDhLbD0m8goef
WpazB/v1ArT6OWz5je4NtK8hTBWAgS9eqM5Tfs0VvO+IvYoO/dtXrWTtTmP0ZQOhCzrLNQTQcK+k
aQjb+GZTRVPeNuC7riQivKBHUEds3xEG33L4M4gUxvNYD+sccjmGl0IzQAejMd2Cm7czyuaL6qRD
eSwPmTBGYogXIut30KXdACGROSoNvLD8O50JiSzYxMxMpvAupCrku3wvFktEOLU7LZI/SPB6xjkO
6x61q4rGkfnPNLHU1WshIgoL/NugKnnwB6mpUGxsO5G6vfsZUOojQHhNibBpgCLuvXwDCiwtED1+
S5xLAOg7WhqT+YHa4Kl/1WnEZ/VooZEOvBQQ0KJbwRH89EvDooErW9So+RIk63henjlH9IbmA3zV
f6QYSs3CJU5TvZ5po1AhrS7K6k7ukcEAzjgjV1OZlyMU9Mwkz0LrSHyuQn3Mmp7zNU8HSDdxeJ4g
UOIu3r17tBuMshGS9STAUSyZT2l3E26zS1nT4MrHKNIAPw/xmweZ7+zpYoeBCKUY5FRHCVBr6dDn
W5ML1sTImDh23W6OyVzdGxGtqyxoJE1jYXMFV9bxyBxTQ6K7cc4uX0/2lRbkNmaZWrtrf8Yk5fOL
gXLohn4+I8URkA5ZaZUE35Z4sj+OIIZv00scruSjMnyH4Xx0nheV4IFjr+xupo8xeg6sO/TRrxVO
NHLJZdv0jsFIyu/OjtqV/I9Pfy+oLokOet6BHGr2vOzo80C2Y+ojvG521e16Zq+dU21qy3UNhSrv
iFUTwYi7YR7nmFmhpGM5AT6DIpMGigAuMq4Yp2XCXj0rDccUILfWhpYe8AxzLjYxvYJoCD3Yh6KU
gjUQEFReU92RgA2Q7sFi4ByAPaThHLQMCpWrPFK8NTXKXaUMlhD64rmTgc7N+4eCCMkUwMCgpsyK
wG2CtNRIpbpsKbtYHT7w1wT6PrT2hY3vIjbKz9S9qFwssYD0ySZdE+dOtWkCADYbFVK65uKrFpZJ
fwwsXiQvOelTCvIRJ84ujK48aSqH7izomIfLxxhjGU3alL89DP2OrTJwFAuQNI0oLXo9J/nfqcq/
SiYjPbm7vcEwjVYxXEzGeqi43xvLTSYoeJERlipbDJ7NVS80siVpj/jb3pX50NtODrPWzfTi1N6x
/+Yph6d0SOCP8qedcIStiLsk6Ibn/dgipVzxJuJLwIIUuKDkdj7dRhH0wD2Za1fYb9vhQ1FSKyBI
AgrZXzeXGVtP2YJbieLR5gzkqC1/F9+HIqkn7z2o15Nk1vGl35aqi5jyRShZD8MFAucJgQLMDopy
cyzQR6TpOM7g2OHW9PXxBcGBflubIHWBxRcCcNmgPj3MGZyvbUdMxVbqwEk3FpU9YT8rux7TihV1
jBalfMI13xx5yX27L+9XYsrNRRE6AYM2vZcg7elD2S8kP5fhsseL0d8K7q0KpCEvHrtxIyv0lgjS
fGB3FKw7/bcEYemOCx+VEvD4AAxuqV4E00392zbivhoHN08O9cHWTNQIOz6NgrZtbJUUMCz+Oq3D
nMVPXBULtPFg20oRQdtQvaS2P/NX+L06cKmiQNbxvdUaBP8r22u1IafrxRaMp6sMyZwPTQhQz3Zz
Rti56FvoE/iuRP8eEMyU0SQ/vNYdLTBx2R1G2lldZP8BOXcsDRpc9nXOB3UJ7fY3vgTxcUtCz9+7
CKad6jfOF3libHECvwMxYf9hCdq2M0c+1W4RYoDebW6L9aEKSVZjj/UNlgVWMxBwNHBZP9kzi4/S
GxqY+35yxln3gKA0R3MRldqjZkpxpePTKnLhMAAAUXd+Lueu2LUoClGhhWIu2PUVqHJSg5GgE/bP
Suug9hPcYwR/KuR3f1mXOPTBY5knC+gvQP3Pdh9IpEvc/SxUZN7zcJD3AjxEaSC0tnVOsrlByMoo
MLbiZKLvZFA/H1Qzpd4Cgu1Vd7rfyIgDbXFRMnkLJS+LTDg2A5/lyIIs9QMLHfyDUE2atIXcqS5m
J8mFdZ4FQMWBjoFeTBBShGGuKL7apfT4yXx2tjCDqMJjycryakWO/vYbyHbGRZbZBrlfK4SdihNi
PZem1SHL5346huoI7/otFlULlqRXO1dxlhNDxAsBjBpV9R67jSFKaeYxOIrDa7+lLsEn78Qk1g19
D1JVlr7gqav+Sgkt2IPr8lDJ+rHWTfElzyYqYIf0cBuccxfT/BzdQ6PGK6MOTLfCjg8fy6Omqx+v
pmkQiC+c4VP3vXSXFq/3rgfNjdV+qi6O/95G1f56TEoU7hKn6R9A+AYBXKNsDXP/qoBdvo6eukt+
FTLhJnzIMLPDAzdjRdxbyQe4asqmiXyZb+cDIV8PlS+oOCn2A+ArFPI0mahn5Xfa6hyAdNPJnEKK
Uegi3lralEv/xSe0ecTArg/A+A6yOE5Oc6KDxq/jhmDtEdzzGJJKK+JmPwq0sVjI36NsaVLx6dwK
/SAFQEHdu1IE65iDbO4EYI4E26k2p5QHoi6W/GP5A5ateWNc9zS6yvYnkaIz9YcIU8BOJrfSCMKP
4iSVPnKzKJZQjAL0VpPC0Jy1aAzl/PcU5PZDsK10EBMEFkvlxtEGhM8giuuZTOedwZfghfH62AmR
Ex64JaM+0PhN+HDQvRZCOupVOd7YRsXfg9NX7pz4HBpRyWp4v/TTMt2nPLboj0J6ORuUcYo0DAc8
JJmht9AISE+P8vlYh1+kff9JshP+rboOdqXy0zbWz9HEjAPa6SbKxLwXBzPqibw7tiK9pgyZ3RFT
irthC5XKexh8AjVvRkvNU/T9phG2WxwoWVLP3fbSjl23PjzWrQr8GxL4HL4YutGZn/JWg5M+pLza
UB76LTemINBUxcrtMwx60hYz5KAJ46L6yCYyrFGcjQm0uL3QLr80wZjD3ntxqhr6qmHbYGctDPdL
Rga1o3NFtJ1nFIOShMMIecz9AMtXVChUi6jzfBOCaiSR/SxysVUQEBfgV0GAFZVvCzNGX4LonhjX
RZFcTihziTzTraXHaHhFal8ImjeuhawUnQOtP3ycuSMlcpm8nQYFXNqtwpyoASKyAhkDngfXqNa/
V8JyF/eY/cyFyrPGIOBs2wyhYYaHw1QcvV+/HYCCc8pfJdwNmB6ZZApPMfRblnnU8nr4Mu6qSJqN
w/Zfvo/1M89dCXCKV7QgzPTOIc7JKBqMLACE5Cq6O4o5CCPOK2HeAJgQ4yuv0YiekrFe4DNjNjFA
+myZVZdq0xjY4KMQgMns7vGE2VjXXrupueY/dPqG47sjEbOXIomFY0YlhswBIlAz1uXFFkGFp4a/
znK+tpaUX4VzcD1zZSZ6W6e7vxmkspRcd9RbmYwNw9sCI81Dt68NdnqRe1JvLZ2RSpBpBx/5tpER
sJ8SAVN5iIBSNG17hgcX5Oofvtc1G7jfsiKYLfeDYf6xtzs4jXnJnPZu5U9BoLBwSO+O131jjzaU
A/+sTqY69zY1wB2E5hY4O32aS0SBP6YKrC03r4SZ4g1P/F153AHmn1/FKP7SqzlCrcOhUOh1903Z
lzuvrreMmpTlUG8KnoGmyPxrWodV0VHJJs0+t2iFbrieQXBd46vnJle8M22UzBObxwW+BOZUhLpQ
+hFX82ZXwOoCCYunj6PtNJpvTKcUsDrTgzbViT7sNBygZ2Ht5MwNaFOqv8wHo0JDGWczpUYkEctb
T5wyDCBnnRB6KluY99FobnwuRwVc/z3Op9f+Df1omhSMYbr8DqUG4eQrwiUHKifm++qB8VhPwQt0
+FUJI3ZCjXv0uLLspl03yShpreDMw3s/17ejmTy/DrvKUnfN2FcFigNjDA/R0qXLHlIrjnLERzlN
4SCexwKm6Dv4F+9QpSEmD8C63b772Ab7te6/0b/yItukQlpTtxRhPi7PBcdGCFcAT1255XkgB+Vg
6kc24KguK0wABoXyT4aod4PTbjC1lCI/SPRWrgmHN819x4Uro5ix307+2eNqIqYcRog6aSuouFCY
EnZ/rXcpC1j9J21RbkuKJCRY6zTfygnZJeUaWWrccnO5cL2SVVjZjcc6WHfdJqjdbzGHBkQ2fpzI
owsqNGhBHIWiVqoeV6unEYlUk1M5LWIWoOTN1iX4FOGP+beOJV+DVIh/9ukaRhDiT7puh9iSCko7
yjwz1Hq38CMSHLmlJlB0FsV/27caPjgdT0I5VI8FlYJwPnFwIuybLXhI4I+SmcyRVhH8MiDB+QO5
ljlkDLqXQgtYjLTBF8/jeFku1oWLovCo86g6u8ZO+n41VpBfHPLf3/JbLP6eGp93eRkF1OGn7chn
8w9Gvurk0RE7XiwlyVelyxjrRSr859CL7hJpPIKS6yXEbswCcTxBNw6IctED4FYSBuw4Ndpme+UR
aWYOU6rAglEW3sonBCXTtxqBILcgLmCm/lCfkgFf22yrVXiK/FFQsybEd4hdHRqRS0i911t/gK1V
5/EI0Xx+C8L9Jn1+rRe3Rh7Q96CaoKWgyyFRvgRcZ8P+CipDQbqdMqTQP8UVZbRoOZJkxV0DsWW7
ZPEy5Po+YNl9h2O8FwNjTlikuQkiMp4I9Ing04Hwb+s1YXy7wNaBifG7KIXy4kD0rQaCAZHi1KOO
N30mAjNWvv3of4USgiVWbiK5jwfGHAw9D/NZ9+gc8iuZ2+xLWobO23fwnwtVDKQEfq4g9/6vtAZK
VYsta05RD9OsFhMq+R7xmnMnABrfIA/RDIxgIcLQ+Kxl3n3AvqQsmil9svRebZB7kEdqoKfgkFNW
T0M87H26dyrU8IZifALS+qpYr/xEAhzxvdVIArhHrtCBlQj4HRyb9FRFFcIZI5a1tOvIhZFDxwPQ
lXhTQiH0sHV9uEzk2V5y+e5xqE4seDXpkVVqVOmSY+zISKbs5w5lc7onwpHlMM9039UpaIcuq82+
EXGaZRTjfpi+03rHvq8h+VCAfcwV1Cv8yAPwJ9bNIM0itJFqxbwRTR5Wc0lhzIYNjNWKAtRFmFXH
oNvB+3hi/j4uGqHAKHI9bPLLaN7yf8tzjbeGcBYtW+ZY8L0kH1F67kJGHOdBjoiOCUaEXTTCkRRY
eVhAtPYj07nQAnRKrxY028pK5TNl1UV1hAnIiKTObc3YtCu6DiZjQRMMCNcUuhpYWfyNBAwXr/wF
XtlcfT54B9TpJ8EXXqTsnlzuCKool4cdeG/Eon/MI8rp3YXvGALKDF9BifStUUQxbC35HRoY0FgO
bhz3JO0Up2GNjhdxFLIljPzoK70BTgMhRaXqFfV5BOwMpAYQbFxWa1DD4U8DD8Nt/q7EwLVLNS0C
Ixf2gDBtf0LLrnN8GJaJM1tp9HE0BOSA0xMk5QH8FBaQ1H9xz/XOWcokBbYot5FpIGn9/noX9jRc
hu3YH5uA27AOcfBHKTSr+xBLq3O7UNLiZL7cvnTbi9Q/YF3ch90ydpRdQQI2ATSr9ngMHBVYrhiY
ANrlLLqiKi22CxIh1K0qe5NZQfItNjJC8oJCT3c3kNXGYHv9LsC2E6FMqbNimhjnv0elHO7y6zeV
0lrn18pvv2VDq51JEwAqyZ8xrx4T/56/Z+hx0eVKBaaqgnafSLZz90plZz6rxJCEC6RqKLnBsae1
7CpPSFGyudMWQuRN+pBsY/RzuPANTqqWjobPQKWF61ppGOrFE2wl/g2rl+NJFRpJ+fdB8tTO4N/B
rCMNYg2GuIjgcSxkJqCvlcqNBkAASME4mhb8Q1FyNguV7ZxmvexTFp1e9E88UVOhCbPpKUgc0vtJ
GPJwFW/YPD8biT7kn4CM3enoYMv34MJRLYUGWzOsul4AduREbH5cDLFwRB6CxTY20/rhNapmwHd/
zr0JopOvLx1Wx9n4A6iYVC4mTB04/dwO3oDf/AmPo4OZtsnlnWFE6xOSznb6TYcmSon1JV1PC+QM
gVmI10DBlLp+pLsfLDBZJSMxIvQ3PLdMJg82Fx3miVOhzUFaSP+ekcNmtVGQBpLjsneioGgmZ/Do
9pUjK2CMiT5nj0ycqbFofAWzLegr7HKr4BRicYLdsjOaYs/ED1dGGc1EDAKii3tn5LZn2ccmv+Oh
6q807u+Ncq2/+Q9BuZ4AkPUEIhjSW4PbG2/1X5ouWC4ryft+iDPz/MZxuDy31z5R+00BsORBqJb1
bVweBMjPZ7PGKvtriUTO6VEWwXOjImIv1LtmqKxiwcZhWq+NezukVnK6/DwAfXvhRkK/ElYoLWbN
eV2p6mLL22K/TVskBJBDc5/GjcGuZ+KMDQhGTuiTOaUtJJOIf8K8MTbbLeqBbfjS0u+XipFedmay
wHFR4lID2DUZUMezxz5ELZyHX86o2iOXJo4AtYVmlS4faV1WMCxAgyIzv3ALqe3UlTnj0ymIJxiP
egijeqJMCa6L+4pl7IE5Ux4ogLTitTBS+2tx+KkTX4f5I9wt2ZWKMutGdy5K998Bwlq5j8ND7xc2
w/neeV38qlrmDfdgWFjyrfmfUi/YOAD/MCacZ5x8/NwA25a7Jhgs0/1mb/iFhTkcqjISYkSErDbw
6L9CCReTHepBoOzWoXDzSiIgz3ZsuBYhZAULMLwyVZJDD4PB1qraYVMJzEI7WFSmvsn9jrShdHNO
u9u/LO/9I9Fgp5JD2YR3+TtXQ9+q3gl4Nvj8LcZv20fhG8gl9//GUTW0UMIvI2QD7/YZ2zt16c0Y
wktqbnMH9LYRS1NIfpOkUwgpUSZCP4oFOYfXn1k8Lav+TWkhKOuE1doHaDc70WBZDPu5nRBirGzA
BYtwkkZv73iBmdoP4FcsB08Bs5yseaDgyOdhT5at/KoDdohzSlNFGuQklX3iwWhsxvEzZFwHi4jC
1TIdOY4YTXmxnstsx8XEeVdvVqsjK7kGX0z5dB+5qreE4kkgaweSL7KHJLUhgO3ys+vBw6BybgFp
6JxVsEl1zaLn5ddvUr3MwWzndvFvzsxrAh0YQvAnHXb+q28HrsGi/7V0P5FHYTzy6NRQcl7y3VAt
fIYcg85a1jkvOkkuHZ8dtEBeuN1Gwbnc1b/HQS9sE73eBjuFpYlDse+RkaiJjO6+IM3jjldp7cRW
n69D3UsC0BaD6OsosCh/iK7GPQVpHbJI1mzwLivxnNPio/yMgXZ0FPQhgEZaKwkh9nMJmDdOozjE
pP3jeGerVnZUEPy/zBjGoIuiBAN3LROoajMkBZkMcP+ofOg11Eck4/l3+Q/CjVV6jxeHYcWO9pza
+Zg+W1LvWCWGZi+zzzH9NUDVZ328qmsS5pDneQXu9XXIPlaSesIZfVouW7z6RJxiv9Ide1KYug/5
/YtofLAiiQEHRIKT9tesNuKWcxDwRarA1T7bRj06W2+mgHvm8eAfH3JUbyZAFh3gR2etnA1bMjW5
h4c7NOV+5Xfyb0fnWnjkZ6v35xLi8mHWspCWdcv67g9P6LfMmkjcj7jikmoxNZXmbfYPe7kgluJI
mcESIFJGTey4XW80R3x7wunvs+xm6Lzl7EBSJb/V+i0Ti7OrylUl0wZ8e7/2UWOJISqxLnLEhX7n
UrUsUAgW8pQLyQuIOLq5PL8OrIYk0GZ0qLU41UEclukZae7NGvz2umS5Y4+X3004Z2TipBvb3ORA
cK87yZ1/P7sr2Z6/lT+IKS5pkICJB2RIWyXksd+4Jyf+5k3hkexrpSr7Mr2f7JvSVdm302dBiUZ/
Op2dx6Q+0QXKT5UH30UIP9xFRidkhpRBMW1nzI2d/AhiFIuXcqiLG9s45drEuKhMF7BTB651cshq
rvcxuUBkKk4b+lywJUHO0DAZY7w5co+oXFGlTLw4t00SmKajYY9+4AK21aE6tkcqlr7atIl82oDe
w7b2bct0iyY52bF6+VIje8RE4D0Bf9yLgcEbqAn2UyQT98U8wkWYh+ksf4wPAehcssFZUFrtr3TD
AYy1DPUGgdJszX1LuB7UWrBsfn4E5gRSm/qbdfCNKJvtLbFmvvs6q5zIUSTRhlAYcAwKsQpf+D5Q
yjlJ6YiLadUEvu3RRkto7jt3KGYY/4WBOdDOj7HXRfXg2gqMLjRr7+iONoB4FSL2fsjQPdhmfXDY
gNcNJNOkFztuyUoOO+qg5QaDr1IFM27gf7fAQquB/hy2TP+0xFjHRTBP7rkwSUBuy4Jvh6AHQnJQ
tfju0RekvWSiK5v20twLMFXm1TOvi8jVpuVp9mK9WEAGSR0m0v5LHwta5FS/C+jk1NV063LA7RAQ
n9to5fMvbuZfULGO9AFYcNTx/r/L1yrmh7ujNqvWyfYlQiWl9RwRs+0Bqj3d8PB512JtCQ5ws0UZ
Ra7whUSgEBpwXWWaTKTTFq1jjRR0c/CL8C/32CFV185gXFOHroZGSBU7mPCD+6pGVMDVHFsfix7b
16aMc/0c94Hz9++g7MMNSFqDJLWBkZLF+2ldZKKoOl3xUUT8iTA1fshIlWbuo3MPZ4mUWZhMEQgp
LcfjbI9xAyygZ+soGahOK9sQE+cMN71lFtq5toQY6zdkHhqVd6Sv13Lsv1oR6FLyaIbk2xHXJn1r
EO88EJ7twETY00Kzy82yj/CS4AYgCtWKf+rM+q8WfDpk7kDnoNk38DK+gund/AR9qcqM46JuEMRb
hPB1L2M9Ks7tRorjI1ZWefQPzzqvNRvv/jkDEY4N/MGiZnRHqrJt0en8o9J+8WZnq2oedbZci4tA
HhQhoS+k6yH5Pqi6VCvBNxjSkWWtgieNbwWSoleCu5/IAZBmjVIFPDBq2QAufY4w6VZ3kegQ1ln3
yrvAQu9CNTn40ELIpeHtiQCGOkuQK06FJnYR88UfIIwLMn8E0vY3bU82VtSAYKRtZ/leMo/WmP0y
UnYNsMl0ViWFt1/tH5TABq4/Yqwwa5QPGWHvQDxwrCweuE4Uh9KktrjAOmZT1wcDgstGJVsSqK3t
Br/l85VYGfXH1dNkNU9BXhGFeEHHxhT3ugZF/s5+1mvGiG1950AExg4PNcg1L6tvCtmzVGhQVoQH
6XGZpf4zhIPWAp+Du35rrjP9rgIwc+k+DPUJj87H2O39vrd/ehzB31k5TZoUCOniE5kGLGJuwWPb
JcHxQfnqjqQP1R0OlSn2mE0Xj8GY7BGFv2o+Zhj1N2B+umRCAbzr4+jKzuArfA1j0yttPZ3ZC2Ba
H2Z91CnXGySATFH1/I1T7VXCWmh3zOYxXxU5q/iaE5gd7UWkVD9pcsuW9jsaY6gJRujPtrqLAil8
Yo43UK9jb6qT1CrpccHlDUIpX2WU5qwcVMUhLL2FxAjMNzxZEMzBK9D7Qs//qI4uA52ef3JL2+S6
CWuSDtIkNb5jKf4D9YOx4BBwdA14V0grAADnxDBccpXt72/MppwIHwZHnvhVGLR6BkMgbQDYvk30
cAGACqo6rjpDmr9vm51CbLwHkF0Dc55WldCLLVqDC5V1a31f/aIjqtjnpunCfbHj3KsfusHZpSRI
3tV5YR2ZP1FPaTEANEt0KXvpNK79UrHJgL/KkupRp0rkpgKlqK8wqGb//BiGFOX41zArV7Q0ecMw
HkzwxNRGdREpyMss6gpLRtQdoFZNcxfhYV7tzXZTQwt+RFczq5dVCf1twyOoCgiqeUXxKGHdR13h
5UQeO8Uii/rdgQs1xKXNjFHOSm8fNo06Y/v5V0759rzkCXtSGxZ+DRbeI1cPtwn+F00nexnnXze0
y6nK1vI8ZGDbtyBm19t5ZbJeDJzEZGDViF2bfFc/Bs7KYYBzjpaHsmryFs7X0gc0srmW78nhNMai
Rkkl+Vy/nkumaMNZRFfzIiqZoFMnXfc9qBKccJfsRz6ZtuQs6P4w6e3gV+Q2XpQdCCV78rQYEEeO
9qhhfgJMH1cnFxqwekH7vwTLNhfW80Njc/V/puE5Q3m12BYeTzf7qABhdK2ku/bChYYKuOgBniOJ
usks8J8/fl5ex2qLPZyuel/jiAhPiqkbDyV+USbCG05cQfuUwYm18TsKS3xmmErAqQ6LaKq9Sf4M
KGqC4tERyOwogtnzbbVHO/WVNgyXLHmtXw9HviOTe396THV5nX1/jbXP07og73AO6FAuf4A15lPT
wLbHekgyF+ThcaAu+VA8YOK14pz2fI7in3jguSsZRJtqLEy3azBLTRe2IrlAO4y/2zw9BBttscUg
JDm9KsR6uvH16kL4UbACuRYQbOq1qDJxfWTCEf0GgQBa5N2aauUbM+P6kpvvx76XySYStosePE8O
vVsqn37Qm5TktOcZLetA1FrAuGJJu7KwgvCyb4oBuZAPXaRQgPo8gzeQPQmiBh/gm2hVyR8LDMNa
Bvcj4SGTYlK3awTl2qYIZUp+VhzcuQn9Ar2uhBf6sjVqv92DednL8Ko8Y4YaF8AzVsKVryXyipEv
EH36gVGWMy0jWWExaaav/NAZbSpKuef9pwYeApAvz2A2wiFktxtOndgPE0vfhJH1n0dvJ2hQjClB
dnNvVsCtw9fH/tIKlwFnZAbfistBcZ7wjkClVYUGAhOO1ND96iIyEJod1gS5nEnxpqgG6Nb858tI
/3KcY39YGylJpFxan97t6x6fapOE9uBX/pcYtleHkD3Qfw5hyHmDEGOo73UmherC43Z/edmjPrd4
RheYENnxYNf6Q8+DnP8/AaA8novihx6A4F0fZLl1sq9nMZnnga/b7HTi+38wl/pxLwJimv57j2DN
7TBI3LaXqt9GWX0SFvbgUMboU4vDXQ40ujEw/MmPTHCEBtzOhAZaKU2oSnsRIG/EzS+XaU82smmR
FMnl4Er/Kj+BGM/XrT4Oq0Vn7xsAV2cwhrTRR6i9rP/UctWj/SuRnEiQCmcE8gVC83wP0nIB0Jkc
DdscMO4Hzeb8b9gT20kOGWY0NwSuWOBkHAxfeuqlkzq4dKEwN0ShsbaaL6f5tUyNlrCFLapRibME
Lk12/mgcH/q0zFFqK6gZ6aQLu+focDjDWjd8EStUh4qeoCwu+Ewg1KipOkwXgYsrDUtq0GDz/J1o
/lStyhQIemq3/DkWmQpnjTK4T7iIN1shv6Hm4ihdLGJVIRZAOpI+nnV+sASkx+kiDWnh7J4zuxkk
l3V7OCTwe8QdmW9S6NbQbTIP0TcZo2qOm2eLULRYMZ4xb/dmEfG0gASfYG2RoMR1fSaFvXRZ4SCD
h4YT+gHqEtAeCDBcuI5zsr4SPd4XXHp9netlNXLZTI69lD4tX1RYXH5Ry2xRqy+129SuYkrNC/Iv
0c3e9gzJWg6ItrEYUMyvfsLfWfCTFDdrBLVDqOEdX+M3jxYmClIU3sYaa3Ca41Ahgx9fJUL5ts+q
QHr9AiQjJNWrQN0uAChSIo6Zz5ezce9M9WOxG0YD+akzGitXWBRCFjyw9Km9l5qeUO71740bLrX8
NuH4wnzJ7uZ8QCbHSyJ4h+l7mseFLHMk26i+uK7IrLJuHnQVUMOtc8HN4BlxuA/nB5jbWkuAjLzK
OqrgeKDVxF89nE4YMuuBCP9vtO13CuUsKO3Vy6O7gFnfDjqbmMWFUQlXISv67prChmo1pYNfLJPD
Ql/ecosp+LD/+yrRmVsoWXCzldVWygsJ9yv/5hEYZn+ZlUEKxLpPEfAWtJRjmb14bJICqGj+y7BY
cpz+spoN3H++F3OZUDSwD4CpoMyWITgYOKgcSvNEmfx+dhlteiCW/mkIiRr78Q0LGgmNp8FrlO8x
vfJEtwj4ho12cxhpnnSL0Gv+BZvWBRdVVKyXrzRz9gHC5fmcWQi5UfQifuW0zZiNe1PLJzBebppZ
IgmcRG88HAKEMWzgPMsWcB0gwNNOVuhd5arj4522dQ7L71L4131exuhhcjJvBwRVBxhHeH+Zcabz
MiUJ31uNp+W2/dtQ4LQNxLqloiaQcxvkSw0dqPVeNd+NLllmPnilKv4RI0lgGCN2TnL2YpjiJQQB
z1LNYEluBvFnOijeXBt2b7XzXj9e1v3OVS1xW9MYsV43wuR9lZ4ENtDIbEmFP2yDDEe4gXgp0biA
khP+1/0gJoXXFdO8PMPeSQO8VDXa/ocbFe2pW0JLhCGxQvujEEDU7mCPtRrRcQ6TINTagmjn5i9B
VKE7t6gpvF2MIePMkIPCNjPOJi9RScoainiW4z6OUpzcLER0LvsrNQaGDk1/oMjpWCzzH/0ECc6a
xqu5GZ09taFTNeVE/R93IBggV8OveX2pGpFNTX4Ms/hDo6tt3698U7k1kkqqmjTZNyk8sZQMoLfC
BPJGnHEb5BoyFpFV+08WcqHzq1e/o1yLxSt43VGr5dwiRBTYWF/Taca8ucZh8cv/J8EyQdx/VuIi
nrV6gOJNnK4XmDrwDdnD0isdjxPVzfJ7Od+bx7n2uG39A3mQEmdxWcy0N118jZNzSAHlFy0mWv7E
dnogaGPvTULYFSP6hKta3+X23kOC6OX4iyVixZx6HSUd24zY/9pN1jgEPoepXBlm4OA/qzE4zSa2
WpsdJVa8E4MMzGyFp0bGRtUhg+FaXhrF6sXdBvsA1bYwn8qEhM1hcREhMguLXemun/nyuM6Xp8Qy
1zkEDycViGhMj2b8C4bU0AGudteI4EKdric+SWkuNRDCHJnvOJNXDBiYTqVMTF620AF82XgaWTWw
HCMvBGgtCEZrTxdx76ZY/dksvBgPn10JTydd85tjDVXTSglzMKYY7Qc/3iUeCR7k9g/oRYBoX+LX
KSMRxLCW5anlvBuZbdWV0EATFpTlDt7FWemIbwMv5p/6/Tc1DCqAVSZswfhfTqlLKrhV8aiYGYcF
NVzEZunB91gZWdsIrIW86f3Z/lLssvL9GKQnJFy19JzLHoYn3SFzhw6o93Yg94oWAijuRiUatg3Q
jMeAnUdAkmBm2ApjhMX03w3I3bqnkbpxlXHsjHh7Md/TtwsFTTm1S//pFyechCTngGAs6Yw53p+Z
F+noezdJzGquOvX7yY4KXPtTDQri4sfsj0Ji5Jz5tx7og6RjEPBWu22nIiu/EBhd2qUwAq7Sdbaw
vmn515HSTaJ9BH0oDwZV02oXz6Cap+t3Uum/pHC3Qnqr5IaHRiTZyXIVepuSQcMmFQ8OpASQwMqj
HSNoes/1S9NbAuw4emgnBi9tW+sFpmUuZ1LCX8fMbwoAV9slp6Oc/nJr4LfzcIC92VXFfqa3E86F
25SD9lVCMB52wdw2sv4i/9PpUHWxemfjUTgRDAh8PxIu6zEc1ZBsggVyuKo+vwR6IP/HdEa2KxYV
+iiz8DjbGnuONnZweD1MXdrWviWUjFF9+6Vxjw3s63V6YIWM9OfkSdegMCXCoBh2qX61uyXNp7xL
yNNcdp6oKfovAmKM109vSzrjbTtQFRpTWPhXAoEwJhf45x06/TJpkjLB15dmZVqR9uYmwuL5R0ZV
hB+jbTRA2lBdUUbcX26CGLXzlPGYWX1tKi3pkH3neKLXUMXBoPnlW17PfXRO8L/DQGmQTy99bxpw
NQTElhQjHcHhDAurRw41SL6lDzBbIHggezIt/4MFhSk+o1QeaGq+qYDDZQ+cYJipVGez/kXnWyDL
X0UN/p8AIllMtQ0Wg6Fphy/SQqRQIpMlLn2IUeyoEPydoqzkfqMACB+Ga+fNTg8khdBghbA1E0Vp
0DvqW/nK/uZ3S5SOVH1DStc+ZVhVFjGTgY0wtK19/6xLpxYV+pOn9dLD7W6f1U8GEK5RuvCrK1kF
xWBprkHNPFkEDWS0eFuJxGH6BIBl5ONzV+2Q+JMttKmuaC7Mqc+Yb8iPBt+vDxolVbpT10R8vKpE
Y/CZIAmNikkTjnxO8fPiPnSiP3y+RV3c5ilrr3IY3lwIl6BA4rJg4qFzKhHW9JLvefb1brJ0v87/
ZqmPypO+ayVm/lGE+ZImdfUenTM8TYn7hw9nijWdbi+K5Z5lwJpQguuKGWtcUJ7Mqs5jCKYbU0f+
kSXxeasNZNVdjqUHUn8g/sBLEQWcxlm9f6JrRzZM9/r72vNM7fpgpNf/vZqMDL8khYVD+dROWD2T
ij31cDI17rTE/+QAIV7HhpD/s/ujYD+UwN4e9sXRw6Fbd7s9qMw2pWcvq46NbMIaYDTtwCcW83Ib
KHQQiBoNuccviGfdiNc2Sk6mV9OqLnCTIHAa907YXoow83WDtTUtaZSPGbYNUakmp4cZ1JboqhUn
jDsLDwk+4lOhc3jLv989LhyaUv3LrWIX72UflN0e+8s2mWNFwDfNmlEV4cn6bL+wmw/QKI0upknZ
k/OwZxgQFkHCP4FBhQoGVh+11vpam1IcxjkfVbYmsE66x19AipgXFTk989yMr16Am9LV2y1s31A7
UJtRE9h9nX/2q/BN5Eb+zl7g1NP9HSgZ9eEPtXynwMDeft8UlLs4ufiJsIghqVXIO0zG3rm+uxz9
c1IhXwyfwOKRWr1j82nVPHtjJMKeXBAcLc73yj+9LcGLG+8YKqLeKZY1sUxqRpYo3sW0XY4DdDBd
Vu0JmgKdLRHUu0YiViSA0B/LwAohObfP2Dk6bdCeBfDfDo6T6DDgUM56Hu3V3uELsUyAv7pXrAfj
Ep7RhGkczF12RPdVx48Y3ojE6yxQv6krC/Dgb266CHqbFTTlcw3LKNUPbL0KZNPsFVVnnZzpOpWr
WT/EEJdkYDg1/EUlGEbsKtq0ROTt2atQgXRd8iHjrLzfIO3zJP48Yl4hLhm1TUyxlKe4ytq1qggT
fSWPkLzw5ZNy2yHnoDrCaw1IqzlviHTot+jPA2XyCmOS8CjRCbSCwxafRn0k9kZIKcZoSKOrAqyE
VYU6WlBd0VVbBoabU+kPrnHVJf808iaxLEKJEQEbNScz/NX5k+lLwe3jcPSs0/NDKnx8oHyaqhop
zfdm2w6xr3FVrU13HPl3WBd+jf3eCOIoBc7OYgORcrE9qZt7j+fQTMA64AOxQ6baG1JARCFWU4ET
VVocO352eK354Bgq3JqF2GHcwwvAxnSYb/46XzkZbq9sHhpdok/MkXOkn5QhvV+cy17PaMbzEtlW
3tuL1peMptV3Ci5gK9TT1djvXNMih0mjB+oIp1AvDX3jInjbfUmsifd/aCIPp2Gxnpb2K6zUD3zH
RWbadFvgprf9YzRb+mljpQsE3e5GgjrYQZhyibbBM+GNGvcftxFob3Y//1t0eDJx1RLCcpRBgtcW
7jZhxSG1omDVlH7BUe6ccEecyzO9lRd4+Mpt3cu1Xa/doJ46w/kB+XfIQBpi3tMFYxNF7EQMHuGU
YsQaN9nlYY04f3SY639Mj0NAz7MhRs+zCpiRR3KSqCJxMOmgju9DnhLff9subjZxCkyvIgKbvt+P
4dtzhXpbRqe4crkFptFpkzLKuhQs8GLzbwYgl6vZfoCC8n5xs18cc+rhUG//knlpe8/tKE04SfNI
Lo0tpoTeZm+YYSNNzXaTeY6rUZIBl7wm4y9yfzLqwmvywfKvFDdJ7WxRv81N2uICg5ulQqypMnFH
Q6l5hOl1Mf019NmYnRtPAi1ay4N0sMo+/NPfvYBmVeGvYTWc5mVfVIr08S8VlkIEWkWpyJqRid7x
c4XK88oE7Vt9DUqmCjuPUyJKy1UXu0SBw9by4KcniRiVIwa8XdXn5ZRETqXVMDW8Scme//sU62Zv
42B5/3OsvNa8XGvPM/qcZR8tJLiOqGUtwZHLVwy4m73Nj2LovUAqBdkxdH92rmTN9bxsWjLxYgTU
7+lShVp5Lut3qfjQVkV+Po2XxCt8CNKHsy6EzKq2LYT7fIgp4+KsUjaRXcMYjUjcQHfvlak2tqbT
e16OE2ZV3D9f448l3dFK9l4W/+TanaXblzju+kR3cgLadoN/Fzh2RPRbiqmc9c4/4zb6trwL/GNM
pQLWtj2hOUGSr+jwv4J7i+Y4t2iUJIkJ+p6NZffRu5b7xd5pzDupPey6f0RtxzRW4v5RZehRKLv5
TAiFEJnPBb03pEHRx3Gb3MCOAHtuJoXYRwkutg7bCb62kCL8ypIi4K50srRBvsV0fa2rTuoEa5ih
h1hhodSGhvh97FWs/BWnAEjzhDMvYNHJTyum3FqsjK5KYoPHqAC4AJxzVfgWQilaT1SMOLnDkZRx
Sqp/J6wyT5v4MD1tXfVcnNZLsRs8vQiEfcvAOXuXYTYHpLrE7qEUODNkHZqfJ8Bh7eEo15d7Accd
lRg5s18Dz2hsZRiDtYDn3p1zYroFTAomhUq+YPw8zCLzfGvUG5m24wJhIwNv78BAq4/WvyGyT3wQ
DiRdHM0e07pZJv/UwXa5n7ZiOHngBli6uGyW/WB3SZbGSK9TLSUx9wLO1M1av6LRPRSX4SJ0pf37
eim5WvZHrmdrLvHOVNqqxBL+L3RJn9dM7St3ePHxmRKaD6a1EiLVhbCgmX+k9ys+psZUqUp7WE4w
7g/hgwP+tK/QOCPv9SoylQ1TGwEE3P8Fy5AebkkbmPxPqtyriSkJSCxCyhJPRW0UnlGrpCIRgX9t
iPdJcy9qHqqdFr9e1UIReJJrFPhS/P8i/9LqOf5N2z8n1wgh8fVfiaHQmEbOTF9MD3CLgNkyJyaF
t6cQkIIqIyhiz1jx/OazS+Kp7wJEAZ1AB2qFVwPeawzygGYR652OjKfFwNJplPRuE8VnM9HnYuYf
+Ad1jcGTsL2L7CuxbYh3yeUFJ8IJZq2LOyJ+cAyjzkqrZrp8K8+8+htSOkRb12kbBBQ2A4CoC3u5
GLiAa/Y+4XNnGzEIHOfoRkpei63Wk2Tj0kpuU0rr/QD8EOGnqq3JYolsYimofzQ+8qKooHNyT5Id
insT5S64cnzcKMTG66KvrAEr8/Wta6nj9SQiv50k0GXlWCW+pFzPd992CDc79qEOp1zDRqXkHbza
ZpeWSHdanCz1EFtvwTw2Xpfg7PtBPWp5PJ2u8kRNHZIqmoJJXjOU81Qk1JtmztujR2LlNIcr8wCR
7qerJe1lsOkdUpWTZmDS8iiZtTWz8ptxcxhTV1avLO3412cU8PovsjWQfAkXQmXE5QB/P/Aq9bcm
r0fBOZ65702U6UX2cjlTpIhj13JPmAz9ka3Ip6ugxNSgcibKKaxtjNorEx/eI1gNH60sYMY0AN1t
xdtnDbYj3G6uuH50ejNjO1VUWzwP7WTrd/5FbI/8B12SkwczYqxwaYWPTgz6BpLTLJJ4inixy6Hg
Jhonj2gPWZHRz5pQj2w52fu1vNu1auKRerFtdPiX3Z7gnBFUA2KC7Mkhc1Ygd+U3RVnQOVwogxWG
VPTBtJefVrsDkiPcQBwAO4wRceq79ucma14Fo489lS+JwcvMULaIJbxNflM21g2bLL4Rcn0iMFEj
B4Mrok54N/qiVUZnbAuqtdc8wRmkM3F6iMmIsTFS3q1ixDDBjoAlrZWTYQjsjIqcPGcLF0VKNGQF
afnQtSv/Xe/jyd89eIUCJdFn/9j0kvVNFe5lAoJV3G8AkFpFx8bS/5PWZ98Kc1SxC68NzPEbovUm
KtFZVbXRPppFjW/I/vftiIy3ijLfoOQcPDWuoXcFxKI/fhw9yAqj74dzzR2CWhCn38+KZxtgDrSr
RReIoyqeF9B6d/n9JqW3BYZdXl47ZywPVWX4HvBx1u7MtuAHNFsQjCbMea3HY7MqczNy7NOS5SS4
1ygBN5UffmyHrqMiKZB1palDlx8ugIxbvS7RqZOAO/xawn4NoZlGaBLnNNYD4fqOatjHVMqKWApz
ZewFhnpxetKAjwHpAavEPiBNKjyow591SZIzwD6IFVd+lWaZA7fZfn+Uf76sUuN/KRNCM4T9rAxE
SHI0+6E6XBA26gQS67DA5XOKhzm+Wt0aLmnsZK8zZuqv9B5EaoWkxIgwyfdNBTmx/G5yFo8Jj313
VO82OXY8eCz4tQJKe0ldk9Y/h5OlguKUIdWLky/IIlr0zJRrjgwcYe0vU5tMt0a4mY5XgO6DJmDX
p3GKbnRqKl5SErDEB6BPFLyUqniJL7AL9UfuLRQpdzv1uBl3K2j2SMXAl8CNk2AXwh8d0rg1m8ro
95qB6784Lnd8vDzoaM3USISDrKOVlXEM9GRRU+DP1Fzn5CW1YhN1olj2RJEsk760O1oBxkxhPUFd
ozTbBMhv6zT0yZAD7aebrmgea2ipF7xT5rDmPBRo09yN22gq/vaKINrdWhKvGcpIC4WEOy6nRdAb
SmcZNP/4gPcjF6vIvT5geGQ0Ska4Yy6foiNBk6YhaMOtgq1Tk94ak/SiMHBTdc0lrrwdQeNrJ1tw
62UPNFc2WYtQAl/8I9kVLokUbNIxXEQ6hGmxO0D67glJNX9TIi76NK5oJgJnRzEfiVjVHpAoY78r
pVnzMBToQX/hMeDhKR0Gk3NeH96VamnQXSW2gjZM0jkbxxsWE6Bff54Dh0t6ozIrz314ZrOQUgGJ
6w23Aw7e8hC/WvPbTTEFrvkKRfG1n+L+IRPmaptCbSnfBHrmx4enjSDyj4z8jZ7zgDzp8aJX0NfW
1nOZkjl1fYp61Gl7ZiihEY5nsLHc8+yPSvVnxXFgFXvZCTzypaLiUCu/OV7G+js/sjazB7T09LgG
++JD2Xc3PmoFNpuwPiv9q0/lzapzKex6qremCYpMwY+vJlE6sKUdpoqwIFsjDMcDkELKnV/PLUkt
FfpW0cXd/5iH2V2mvyjH3Uv4ZgJY1UWd5D1sdH5csoVU6qttstU8IFbfTtsOTAtRcWwnqe9do0W8
D21ctHwhcK34dprp5UCM+W+0IVSxYF7SGQ+9S5lvNOnVaG2qrHQCJk4BmEcmX2geQe6siI1Zj9Ew
eiwzj9fBGcC6DShcXxBj70GouRflo0MBOBBRsXoJQ5Q6ge3BZ14MZCzT+TUqnqKeZYlqUW1YgDD4
kVZQAnkjat69D7qBkn6sWMZNEjCkza5HCMP56QiHNNiz8g0SzvVpd6Xh8OXef+xHuppAQqyLZhFb
f4RNkJuH4fpznwPLguB/dbo8kjd/dpgVlTwUJ71I6jGUoQEDreCB5EcIMmA4MUn1caloOnjHPmc4
OA59jX3tMeRrKjD0/M7ajldVRsomSqbk9VSkHGOrSSeSJpchp56Ap6pTexnk5BH/lQ4rUQ0gTEYU
XLPYCFfoBPjnVgnEvxEmw92fkN0OvD8ovb2O46BDVsefDo9k723RAFdaPLkC2d2WFhyc3ZbeN1mb
IgD8lOC28tR8D9Df08A2pBSOlU755ek3dw6gKLvLRLR2CPa0sO5pFE+P6uka0+/OQLZHAcUG+cs5
D9okii8QxOBwwcQ5gqzcNIz8qHttrPHO1kqFcHI+FwbdvI4x5haQu536LTcO4UE2P3H0vOL9d74J
Ioms0MyhuZq7PbaYvWnK7WEiHniQFXeFJ/3Fo3fIEAJ0QO648Q5IXuUlzgCajvhL8f5RbC33NbcL
reNbLsbkyWSMoIDtq5qPjv787kI3XW0YX67PSrl4YplAASIYjgGdFNwk7JuDSDYDW3BqRMdnPfkL
DOVc3pPyRbWCs2qedtzsBoejV8N9nQKSVvZlGcqK1RKpXdxpjV29lcd91bCfvhVUZkYldkHjGVSQ
DyyVAy/CaK+An0UkboMm1Fy6BBYe+4AIxmYNNJ41hHGbTL7Sbemy8eGg96b8f5RhRXNfqCXqGtbe
m8sz4jKrbZj4aGc8MAAlrbym8yR6AiuLGWrWEATdjO+MHat2xW69XYxRbUcNG3hEaBU7uBvpMTTk
168QNa6E0TOC/7zjVAuB51z6+/RIioyTf7XsjTUnToRr5Ubtc+9suLSKW85RegzSDYUVSf1T+w25
M3i8wBbb/VWPhzIvnk+QxmNiAWUaDxvwJOz4xVbPrueqlU1oF5gaCaTskbQWvM2FABnCW/JkgF42
+acrJzuN8utbLQMTyhS6V6v1PN9ghYkPMdzPI+qHbjNipDAvpNLmDMd44cE4k2VRbVbPkNEcNTwE
yczWZJl3W8Gii6ea25erRLfpgRZgVOu0N18Rtnno6lRcnZdKy5TUdNkpKOv7jV9spLnoOAMgEJG9
KQHt30UkuqcpYpP+zJE8hzOxxikXYkPCNP5Fa5FSmSe1w2HBZIdp9ajFxRrNU+PFnsqUHLpMGkRG
ROWGglox8HuRSmThCuL+7tUYX3ttBSKKtxMILhnJVILJtVREVErXMVs3GCUSKZv74MOGRuFYpz/o
2JarMf5BfuvKPaVOSLpISiw1QsbIuo2KxYHY6N/rLnaS/btQyV9HX20p3oIasHqMw0ZJOm2kBSCy
i1i0cFCJz1+Xz/3iv1rgZbA7NpNV8yomsJ1YrrEfb4V4W1+nhmg4BraK4G6sS83DyfZSUShbY16i
AD03EIa9bfLkajOXiR+9waI7ILzEU3V3+HvgVMfzkTeWFelUiq5oAW3FrxDR47bbb6jH6Hhfkvcm
CatjDGZn/AXpbjpZCwtAXRV4xAGKqN6wYzqGp3oFnMd3P4scqyqRGOODGxe+r8v4g7Vm2w2/us3A
rmh0uitGheFTVVRJ3RXzQo/lqIeqgIDcEieQmAHIQyd15hgJ31GwxcvRgYIRTdpOAkI0qFaypziD
eWtkriJORA2XE9jYNUVkIl0Lu7QkiE8VbxwB0R155gtFubu+0+kYmuiXq87qfnqk5PNf9YsFUfJ7
IavKtPinuQyuAD9YTnzNu4UqsTr92aq8czo5CmaRjBntCz1JTVksX5CjbRrENAKISAjHb0up3gq2
C+o3OSh/x8no0h+RndyqMLhT1s1tGMrg/U7SoqX56b4nw1/lcqRlzZ78gA1PKJu/aiVDTUahLF7c
YqAkVQN1g3Uu6OmsMfHwZKnodx7jh+Oba78ci3r5U3cqUDf0F3CVZR6tinsAYiZCPuIdBZ0Ps0P/
mvayS5cP5lDF8Lc6dT2/fVeVkIeAtm/rGoWbH6Elhc78Tpg7deWSAdwwVLdLiRZKp0t1k8LvaYPE
d3gNKZQ4cs4EGAENbCZ0iBWHvy+isHWVRbwMTpLeIc80VdKRZwMu/9mQWwCYakc5nC5PcJnhGvl9
KS+rmy3+iZyE25Gfuy2cDuH+7JbrQnNOKNM/CUG3PW81XvxoBMap9eVZPskAD6pd/7V85MH/HuZ1
BG+2mQDbCfbDk3/iNTUmRzapQTOk7n7QBTc+m94n0/Vgni7vrWhUEOK46zQX7E8kyodSkFl2T2J5
j9rU9u0iPzRes9+BX+79nJhxITmN6PJZ5/Iu1zb0MYwdjS6hIoeCpr9pORzuNkhF1TB1E2xuh6OR
KBeT7557DElXgpibChprl67CRizEtlpaF488K8hEsDTk2mWeqCiXGCGZBhhfGJwf5APQ+5TNWC0d
NDxcWLYNrNG3SWDEKdOqp6+OOUsRfGQxxRFDwmTGs++3Yo6b8gDfkMCE9GSnS0WUzn95iBQc8a9h
ihhJbDTpdT4OeA1cNXZoTLFtFJd8ZWTMkMBi8x67YZC09kmZrFStallz4bNlXoHzypUjcUaXr+lm
TCnArJdgdFwc3Bnz3+JYk+0qFgecTNFDuwAVT1UTlgSZ6X+cuKwzsjJfdikbE/CJFcv+aEXj3H2U
7batfscK0KXZqGY+aKKmPyaCLjvFcTNE9Nbl8BSt2qkvWj7SKZT2rdDxXZ+qgAh5fw93iwCOCftV
ZFPh1lLxuRjKGbGOwi9btSoHbvBUHDQK/BQjY/VsPPdE0MQLvLTO0F+0m2VHjeWonqcaEb8mN9Q0
n/a/GZgxzIxL3ZHq2Rp20YMArrONYRGkpeakVbH/YJ/iutZS+1Cs0DW6O6fDieedFcEEBytSGDm7
ivktz9+yTBlUz0MqFtxkzvQunj59EAXwOFAnpwcWAt/ljJqEpoxW3U5tDlsOQJeZEAA8K/HhJB4v
53jWm6mgqEgbGaFq2/pz/RL3Va5DAvQ8yeCIirg/vzaULH2m9lNdxORZe6bba54/19Xg3+iZXkiB
t0o3wD5UBSlYLoQlW2YJ2+uA7blnaAj3dkPFFWyDVf3b6p9L/eU6YFhzmsLxY7vibNIZcQfV/Nre
CtPYDy/nge0og/Mzbh5juYkwHuCd0CDnGDTJFuPgmqsxeHb6AibcJM/okzp8O3aG8xUVqJVAesVb
ZNDBrdvaFlntxMfxO6MLii7LsnBUqrZ14P8LhZ/ldY9uoA/hy9K/L8v+7Z+lsnDeRDcM/5a7wjzz
yzeTHPpTonV5QJmbBpy12wLfuVe9433ML0mL5gJJo9lymxUwekEeYyIe9DyvdVTfmWIeN3iEQKAn
BxiQ1ZSO2UjxewAX3M3cJvpdK1sLKcTmN3+FQhZuahCIbOTxZxREvmtCKeEtH+gi6MHbvJiRNB6n
Jx+NRRrKzeLQFVcmxhBGY2UbovHE+ZWyOef+azbpX9yf7Z9B/LznmUtfqqT9mJtJACuUeD2U5QrG
oOjpUjgl5I3jaz8c78DGTK5oOdFKXdg0lnE41lhhon2Oi62+IK+m352rdWNvH2wll0/OKwQy5Dy/
eVA4tmO8cPDVylvOkZqZX0dCG1hZgxEWPZi3BPY+OyPvrvpV9614qZOvXZPFqZLl0WJnfgza3a3U
Dua8MiwixJfOzjgD3NShi8jZtRRP5/+CIaYEmY5uj42LnliUMmOBo1oCN+kQxWUCX0vXo+vtK8Be
2ibYxj6+kcQr9ibxdlS/PBZD2mbk/oEjfQsLvbtEiQuDBE8WPiWwtSqyGQr/hb6/xfF3S8qaxvxR
R/TvZTc6RiS11aio9oCQnr5gAjbB1qRwh3vZtCT3DifwBXHRjYg6UdqG/4nxdI7SyItb5mlELKlg
rqPViDFTszWDQOt3g84MuPUigabRNtp5o9OjF95ojj8kvf5k/8Y+zkdH6vvrhKpLR9zECnnGcmba
i19ipdLqJ4l0Jf/iPyaFdyLg4zFcpMUJ8Snb9r8pRAMYvDfLLUacaydhaK/MYt8oqGrPMPVnXGHP
t6AVSX3K4iHpE4dTUwyPmzH2fNx+M3URt24adRfOLMELPt87asKYJH4+UlmqCNwqe8F4kpd53b56
iDUFf+N6qVtTURZBKhPXEAwyYQeiZPc/T1vI8HsQUZdbGglTOiiv0Eqxl0zf2AvJAkt4LEdBi8el
U6AYk6+NG9YlpdurOBkjCl7pshzBi35lNtDFcTi/19uP1d5f8TCd9cKPICLZnO1hBldy73V3OUIZ
dJUlA3g0cV4i6KtjguHKNRsowC3FKbY9UtbEveRzX14qKVx8wP4tycJ2Gj06bejf7+ebYVYj0gkv
9LXX9HyAapGwESQyvToTeFjbEAHfsR0coJFqwELqpozIpf+nWIirAxLYGgXuj0J32uMK0O3SoyKc
5/2qxunE0/c+1WgJTSTXZ+BcHk39vRJoWUgyQtTEa86UnUl/MbYl5SmVT5Qm4GZf5AJntoc87qTa
vKcDgaRUgftzZH0+gyNHTw6+n4wixaS1svYU41px1jPkzmWQDYOYd0mJyb067LcQ+mu+lVvh8cdE
T23DZo0rMY48CMzjtBHNr+Fh0TAEtuGMKiJHaNiCBEO6K/mupTdzSMydLm9rCrRejR5dbQCHESwu
CxG3SL/M7XqD9AewhkYDxIZpjA4CdhLfW1It41kvByIY0qAzbO0k59lSe9p0NCfZOa11keLqYaYg
pPb2vAeaObYF5RvyK8hDD0mupfoiGUY6fF8S/CbmcLX0T8I6kF8dvG107UEX4drHskdrp5dxcBSb
RpZrchUMCrzTyDcwKVqN0rmgvlZ1t8peV7erR1uM8TQ0jWkBkMK9vwXdjCpyuF80Hx/+eSQyu2kc
Kw3MbCuxi/YFdbheEJzzYzpIdV06zLXLh3qee7BsvVNIZU3me6mHa0qnKS4TiROJeDVspygJq/CE
GWG4UqTYMzh3jB6v5U/35h0fHJgQrbo/KhgLY1fD7Fu/ImlyuMT21P54er2nn7E1hrnnPLkWvb0i
wu7f9tSGQyYagGXej3AdknKClff9wPyJ8Ru2YilwpjLUjEeFScFW/WeKV7QExpReHaOUq/Ani62Z
07fznrTk346pSzYGWS4SStPTww5RHI7Rz7BzRGRVjC1b6EzhhGj0uX6DzfAtMqzsaQV8gmF1uyf5
RYApfM5IqBG869ctJih+HT9gDsL0Nt3WZQoev7ELeCU3WG3r6D3vwlkxA/b0g6u1PEQROQ3wA5jw
8jIa6zHi9Xqhudgrz1nZszrn9NphdMKFSQdfGKqofoxxR0+AcHsEZh7kd6zZUNO/M9/nLzFYUfkx
xrxBWHSaT7LT6Gyw61uhthOty1iR1D9Az4QKTI/NOdnW7UY+1rfWYVJa1A45zSur19JnwC4Yu5P6
qDJS5+f0hVdqtbsDc29nAmeR/VDY1lL0M2wxBCCxgdcWqQo1n6Qp1aFf6AyP6sLZn5RvDqv82+hx
bzt1G+3v7ILCz0ZSu0lY3WW7vU3okdaXekGeaWwbn3msoEpKn0C8Si5qMT73T97+Rm/gnU0F9tWn
JZ4Ee0LqUvOQcwH/mbDM+kW+OWKr7OVzNkIiyEuNSSq4WPIgflXF0tuxIiZRMP4lBDTdZ3l16tFT
5eM71zwZU0j2N8ae1GX2xaT33tXy1fkVmCamTBM+tqwcu6V2HzQldGcTatZnX4TZzGSNtWncqFPp
jPr3kfYsIFkN7KOFY7cbmfu4cJwd/Rlrh7FeJdPNRcSnaMqBWpwVVh5XLdaDFdURc2Fh16IeXVhc
UmIKZYaq9UeJU6FTzSdwgEJeYkFuRweInbglKAr3SCRuJPKpQItTefpMtLKO1xypHVXchaAnobZI
CRPZrtEr9YcmVPHsWRpPXxgSBa4HDSMqhg/2KSyF1ZUcdLIhWWJ7EcTQMBAemYl1eSORQGWdihkk
ZQLvyW/yFk4gi01wswZPJ+TVYifY14Aanbd8SOQcD2yIY7/2GycSxIPJDsVnxfeYe5plEW5aoEBj
botEjMBWHrQLHzEBY4UQB3ZB96W/bbxtZXPDqZmRuVfOpizEP0o3glaTSD9uxTNahK/IYcvszyq2
nEa6llVLEjoNJlRMUix9RP3XeY7f8gUDogz44Za3F4OpgdoKTfT17NEVW7BLY/vHZwgsFAbx/qSb
K5YItALqAMqFiTG4IHV8G+syJOlPC6pDnmJaXNd8xRIV/hqF+i3RyQusEr7HSHDRRRcm2vGMm0hE
VCVmdhfD2N9yocIcK+K9Je1BsVyTPZ5qrzIaLMSPbzZ4Z9QH2Pp1sXpKD2TnEqLOp+Mw5+BHjbkf
7a7j30CEvC0uk6r+OyF4du5drzcb7m1WYmIl35ZP5jNK9Q7kof6tT4t4oDCDgD8wM1bAmmAbD4d/
F87NzijIa3+CJ3eBjWIz8R9F+jBaqBBCUPpB6jFwjajlOwFNTGeIFhKsI2iwXx5c5mOCPqbYF7+/
Ut+X5NKUZUkohAXqT0zukTpzwEBiQHmUaQOBN1ABSYrElBwu7+UKkyOJLpKChEAaq3cn1Onv9FLE
KOE0vbUCPUObxkWklulV/1qeoDewH1Xl8vI4zQrY3BpA59VMziL3x/4sUF8nE1hvm2sQKAd6hVLo
LUXedJ+0x1DkYZm4OJFlgkKcWd9ayOhVwNYxnRqfSkImUGmyPR5oxdHW3BwkN5hpdDQGPdh8qiQP
RkWv9gTeFsGYoFLSfVkkIQki4FL1ikezu6fXN8g9t5wDZS9ES+hzjviPHEf59KD0AxHaMd5tv04j
ZcOLtiUEcpmyAWkc4MZb9Ft2wvIVsKaa6JHevylffXu0q0BMHJCReEVBRThcqjkPfdlnRJ//u4IJ
SK2m9awaWyMrOBy0AiY8BW5LTYSYRdmjhfaS9c0pJWs9IoHOnatmp40G5qixB+SvFQICD0eInJZv
JFbGpw5RoDIEkoFrHz+IEnkd6z34AoQnaMBPme8+Gz5pHgIh6bL9aVOkd9O1Tct6BjDlDrKbC+Sy
/qu0QZ9tuCT3RXZbCDxVu4HPTYgT6jHcnH2B1YW1mxEU92KluZ0CVf/+IoCs8YMg/vj03WSKxhK/
Nnl7wcCr0Evmz7VHdRo3SZpYh/n29XRcPQg56kWYZjauxYoOyXzfICgLnRo9E23ptVGT2Dgpeagd
TZgVwr9znIJA1Rv2y+bkFeEisRqyC2nfwZg9u6FplV2/ZuMG4bZaCcb5eNUoQw0KFy8sriUHdePo
ht7vy0UhK2qL7X55KswdHGvuyqrWPbG5rLX2y0l/EOAxZQOS/QOaaze1dmJy2IMGOJx40SXIIXQ7
dmUeiZ1SkFHuWwjOwvufzMNZQZPPjD98X7JkT279RqUh6VmIYeROxUP0bq8EY7z1iB4Z/Dc5fj8Z
MNLJNDPQfeBAMgD3dxndb3RiZRJekykwwiHFT6ao7XjM8afl2B1Vhi0QCBZOu+8DJAI4iZyN56zt
bgRYLWaAdNsrmBhGnyXmlvsFo1tcNvO6wEv6ilniTBR9GX7Oo/ph7wJ7yOlp5ltf9mXIGZASvKNW
tadmS6JQi1D9+yS7bvKPgdFJsTFEqcT92u3gnpZHphGIQcUNu373b8mZA7CGTV+UnKjFdKb/DO+K
WTudUEyYuQl1o5TxbJ3AJT5allt5jLp62WmK6GggaNdHgz/GnYIjF75LW2HGnSNJaYRi0fAP24nZ
Y0JMEI4kXbVmeIirFZMBYsd50JYgVhH3n2X3qJSXE6GQ5+08VextVNT661MV9mluko/rP0rslkKu
QYUh76m+qiYJXR0qNdRJ3CfxuUXvl7Fo0QkH6H6v7h41NgCo87cdgSU/fMUU82lIqyQcqMzNZGZd
WAflWYOVvi3jxq63cxjHObX2IPARq7/xvGVrPQgAtd6bHCDnXzJbtqnh8C8+aLkZerX3kxV6d10Z
KCa1Ce9Q+0/62ngdQaQgHID5AcGZEA9fpxA6NUwNNRSeZ4ysU4svmQ3m/LjEo+UC+twIaPPKgFHm
wxqB+F0jYwLAKeb/jOek1kPcqBF7SMEgzN5lufhWO0p3LE1BpXL1/JMxVY16qPPQDsOAhQU+n92V
H1ucabKSBaiDhQW8eWju5HBmS2Ve4FEGUiUrRlKOmavLTbSENOWi5d6qpFgsoglppZ4lPBfRgw53
2Mu6N3bsg7FwyVynrrV7UyH9MC6UuIas6rc9elF/GFs8eITVo7DLQE7onWqU84W5RzZqxV3mhFUg
7CnP7jZL1nvb3qnCCxalbDXIszOvP6fcts/3nHD6ujyxsU2nW649QF2auroOAJCg0OEg9E4s2ogL
UkI8LuBk/LqiwhmN0XTX3+DW3/ke3jB03vkwI89INIqdt4sQRlRrMALtY4UcvD3u70Pt7dw819Eo
hIVQHs7jbrIStmvGlctQ95OXoQLfP+4TRwuo0xySTXYJEzqLJKfLrZK51skXpMHrt/2VoKAHIW6U
UctU2OmDtVpLVB+f10hnaXz+EmtFQ6fjoTixSG2o4H5sLF5+AeX03H87Eu0UE4rqGp+CRVHddqOl
9ILSwag+UFDLEx+MQJeYykiBiaxeHGT75hKlvFpdHwS5HIxX9m0Ui3D5AI1b7+SPp2Gdv7ZJ1MUt
YmmcENLrGihW6QPXN8Je7TE8EpNuW05TpVvk9ZesbZKugJbUYKzksguiVyc8ebrzzTWHStjaFToH
ok2n5vv5B9GfWTNwol84NvvC7oZPyzx1xQQ1A+OoRSPXdei26fJWjUuIKQtqAkq2MDSP35rtOqO1
CuQ/bHiIFT2T4n58/IVA/pQ6U+TUySMC2qtfx6TnzOeIiw3P0/jCIK49az/6BbM9pUhpmRnOGY4i
fuc92cl9GRXWIEx0Np1YIiIFiint60OU8MtI4KpCwTktIbmhh9dur3WoXWM1jH5jY4gOSFGRM1Yf
ryU6PDiXG6pbbwt/fGHp/2YMxECOCl6YLCLdfS4liHP3Yd89t9EPrDQisOcqnfgAT+VrAz85Fqbe
ViqUIQ1+gAIbEUf3944jFwIi0k1ARo6cpe/BmAvON5abyH1s/xK1Oc37wS8SkpiXoHk94BQz04FJ
U82ef+VsCf6yyDpx2nrMaIMHWUy8FWqIpEyYMmNdGb1bV25JUS8UurBmaxABdeeG7U5g0ifUKUGk
JEcVrN2MjO+NlKtpmmWS8mEdXZkhSEre/beJ4ul/15JJzTFpw0flI2oumFokB5FkDzzvXRECNtm0
GBkrOJWSJtptUGRvQZiqAsybOCY6ZCh2HEgQ7ZkeoM1E/0o7oWNVEGIADPH8Vq4VgXNPL1tPterR
1Kep7g5JVrsyamZ6rag2SBrmK02GH9S/ZbrAX29GxwUUJWOOjd90JByYyQbkaEkNFRK5dihfSQL4
U1SBQc6JhZAyb1uAKyt6aZ8TF5r3Ye3BLR50Nt8ledDbrZULgFWPue9rZ2Tj370X0vKAdvlLdawd
uF8/FCrpkxKHNRNwbOtAngKdEW1j0NgKYb1ug6D+sC4RBiWu1Ccnd1aUkx4HKlGEcT1dxiyzhNgC
7Dc6elTaGpSss5FFVM9GwnY9dkCfdeWYhuJrP3JIX1EIAL5QBz7MtuKz/KRk4tSgbywAvocHnIPr
aGmNUSurr+R6tgfsAoaCwv5uKv4sYapZfbVTiONX9SNmiVagH3uMg+NXCO41xbSJaYO+Aj87LW3c
b17TTl/L192HeJPksnOIqAO6ayJ/hK++npHq55q5wKykE5omkQGZ2J0fTAuiIoDoFtO19jn0gWTL
ZeTtwQe1arbbNz/h6yClOwnW0h9kgBWkgWkRoGsclfcNvsQWds9xvGIc0hHMyXKAHKSx2GGiy5pA
1uSSGd5oW5EnPmBPSCmRPixJvNvGzqQjO+9fLTUutF+vXkIvS05DTpjUVKECXJUPfoMmj5ug7ygN
injTnydTHTuZvd027vPX+rzx3vVr+Ek1JCN6yXiN4mOnEgA3JnsWjArpuypLHFuBj5wvNroarrhw
1lP2mi2uXpoIVAwZi5WQn2MjOMpJU6Rp12DgRDaak5JtPu/qj5IT5LvDOVwPX8LOPeIIk02bUFO7
//ONH0Q6oy5lZjQQcLUDZ8jfruoTLOa/ZdsVqksjIt5z45MmZa/AcwS0ow8ROi31xJBe2v4YREcE
r6O2i0O6yM0J+clj8+ayzYJ4XwgyeSNkcdFvp617iyAwKjE2/xfHIZERrHY1VpYW7U8wx696veIO
IC4a1zJHL3yH0G5+1KG5zTHzMzoGTGOdZnBoO9dcGmIP6IJXBKfgsnKgQunWmnwGfdwR6PeBqW+I
0rWKscLdZnIna+8FV/U2vDIFUwYuTCJ8CZfvA7OxUY1myMCebVjNZpZXvkJ4r6C2KgfMHsxGKKAc
adc0TvR2OgGV5F7CEHZQLqWvL2Qsgu/FS1mJEnmtRlV1h7VvJGbF92Jal4vPDGxZwy+JcohsrR/d
RXF/6621dN66TZS0uBOBOSjeOyT8h5cAw4J2VsDlbFeoHpc31feFaOIzH+cLYR0uqcOOh6AmglUn
7QZkJthPx81lF4fovbn+ldRFRtksrbQCSY/DQCEleZOIelPzbWSIMwhzMBtEH3/0MqmTFFmrmBz0
yboN0GPDRgT6YebpuDpDnG85gCvtVM2id89Rp+Ifl2ec9XG9nm7OVfdpBfSbqaM4Xt4BVePwoEoX
t0s1DQYoljb6LgzYa1rKa8/F4vJKQ2qsEU7pVyBFViw0G/k5B2SKUjvr5m0DjQSpgIoF7bkQK/TG
xrdvvcgPX2JmXtMkHGdZ48hRQWvc15FqgLhSdXVyobHnOOpK7b/LV3TAQn8u7vrBG4VHF6x5EsKo
F5IBoK3IZtombhvWqLsfeeNZW97+oyMzljWjEdp+sPYg8tHr2FIoQPYSfchSmVrAe1x2EGtrV76r
8ea63tEdL2h/sqamp78BZp4KKAb4r3ez8Obb0as4oG1GAFpnhEKcdd1EqHHg+wEsrq7PqcaZPVxp
L7epQdXr0DMhG5x/Vk1tt8Bjz75a8oDMeSpX7jR2ssdlQZ3dNgCM+EgGDOIaV61I3Gxqq6KpwiSz
L1//N8T9eBoAIcOon+xzHBnYkPEHXfevEle4YBFNI7Ys8IcY9/i10nmr9ugNnpVy6kExLyKLCkNB
SVAKhErXGi+uZK9PMNpz1V79zaf59hI0nEI4f3/i5YUCYXMx7tWj0uJl3pu3xfS7YloWYMCF+7Ig
c1gCuwugqqSlAyg5JhhXkz2s5eaaKsU+PzzUP6DMG7JxgyTxgsRRbyhoZZkVFQRAZRySBvHWINzS
Msh4yyacgQRqfV6e2ot47MiQav4rf82nZEEP6wHWhwSyuyHl2wfUYXW+TXsYt2ZA28bpDUw6vU6z
bAd0XyfOlD/V49/TVvFaufw4Zf+99E1ic0M5FzciRF0HH/+iVnRbCRc44owOEUNYjbzivm4N476s
nnnW0M27q9hKY7flgPijsyWobKjhnKOqFK9FynNFv2I72SGdxfE3baeHfv1xYQpeSmmUOdJyn8zS
djoGna99UZWTtveezvnKdb9Dh/TSQOVwtFb0/ao6rodWRc7bChiP3+vyRoznK/JUtAmGoZCwhsW1
Q/tjzTThxPv3AIchTrhqW/GaSSjSMaiGXTsO+Fp9Hseun0rh60gz37bGpB2ud895HfUJ551XrLQY
uMgZQrd8LQ9YFedapZeNkyNc1YUNxTfEDbRFSeMepZnDoP7Gm3W6Xtsqt3yvNqzTzElsUsb5crwx
OkUYRwQfhvEk8Sdq28RAV6YHrRu4Wutu64A5VysY3zIgVu2pltYaIksOkfqJ7PDkxWXHqcG06PWT
NF2JwZG9QeA9V88BHzbJAhNYi33tngGYCdCDa21gx40mCKPR+ksAMO1YOAECgdYxZN8He6WcdEjM
K+Fq9Z/JbllYTZ6q/tQZ+EzOVcmfPfkrknMsGA/BmIJWoNJhElGe/SPKx+1QT63Uh7vE6bDETPV7
g0z4WKsiyHg7js1VGFeXJoY3qYECvrAyGj8L+lXjz6jQN3b0zR/8pRou3QG0I4Gd/1MYNnTfsKwF
6ZJ0mCOcr55CkqgDa3VZOAqumPcubUXMoyBs4ld6LVAChWExLIGAqkdIf2i69LKi1ONvTkNTbFqI
hwNPnQQF8asy7PsvqtAOOzx2DYTJmqqBgOijofS//BmmHB82s6Z9znqNuz4b06pc9OemoY1JXCpy
3gv6ZgPZME43knlWS2fhqVs/RrlcXxHPIPZmzpI+gBS2sw5ZSh09sUpVsuWg064dqG9ek5Cd9yda
my00ycMafRK9gbw3laRVpyE1TNVv73M4DWraRVHD+Fc1i4W5O0DeGKXc31ECwSRwzrE+MFfjMDjS
wkjf0h+it8uIqx5JPP20ue8/Ciu1N2Jvo5UJFyqQnaDPBbpp5Md+ClyGE5B5Gt2PgOcSBRjftSVN
XtNgTXiu6EOG+G28h5mj0qMpjin5XPcNJbyw6+EuGgyDenlfsl1rsqfh3W+dCCWU8wRZav17f9Io
WzQDKSNbPwic6pRbzh0izjdcXlclz8p7q0hY3ylmerFnQxuo4ZRge/urVVGF0A==
`protect end_protected

