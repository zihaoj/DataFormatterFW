

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lvSE1wnTbUzcyFaEkCK/oaIwLhSg0I6H5NtAJDSx1lTgwyyckziPTGY5rLYavTcVFBRHCSV5wXpw
oInm6nX4CQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
c46olHU3F8bCjhyybwcNX5+VAFexzs/MQFisGTAzMX/KyUASEQnIrxg8MhWz9kHjdnq6rKc37dVG
1ZjbIdn8SkMrZ6jO7IRmCdIwB2EJTzAsoK8YFSf+6vyLoMhBmoDwezZkm/1rHqzqGVbjJUUQF2G4
P62ohvDWyPWNNIgy8JA=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kk1hNe76KGY+Tdlckns92+3icZXVsH8SqvU4x4kYPRWgztibTY8vqSlNrsqzBHJdsETPt8u0QfLK
rDuQWNGJrxqMHSKFIsyfEfs0bmfsNV+V/rvrW3PMMpW1qQmLdTz2AR1aqM9ak/yz11TVvd+gg1S9
8e43wm8aETQxbosNdhrNLl9/0F06bpoxxaqy9pAztWtvjybX0PbWTo7mpZOZXhquCHhDCOgAUoVa
iqF4CjXc5CNxWspFmUpLkXJoG4RQW+ZSYUNweVqwAL+zY/NPkwMGzKXDJoB7oFe8gr5J6WuQwXzJ
K4AytURqWSKZO1uQyvsgQcXrmvaVAFUnfFq0/Q==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2meTUxRFJcrHQ0hBTBJTkVAXwoHUYJpgII5GQKJSLR9629yOWtHT1gVQQ+/1DiJqelxMhOcZUTQh
U57QePWpJ7XVAAehftRjhyRKZvvjOSXsylQSyb1EU5+M8QqtLhmpagSdkcuEV9aR6SlXtPWIwzSH
4izOxcUZHdfC9UgUzZY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lt1ufMLnNLe6MPpqKfqVCN/YfycsVOQhsMH0cw/qRDjacuyDA1nAr3hI5fo0QPXNktQ06ZB0rz0u
+2ScolNa5DnjA0UdgIGXLztxHTJ8oj+Me1AK1QclJZE9Fqj/ihlVWPX/SWC018RWnpzz+44QrVbR
6pYK2NFPTh+zRUOKCLlQSCa75ftb3OYecza1taUkBWsh2vJaK7Eo7Rco7jppMAvQKKHggXtDwbKk
/YzMfTJYfkOVud9zn1XPdRy+927MWTUJT4sKcU9WL+psbWvcWsIavw5oJ8LRjc2oHQ+z8fF8NEvV
PcXHGZfB8tkdxiwwYgEEQalcaKorac2nBssNUg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103072)
`protect data_block
1Vt4DVzWrS6ic3Zuc/inERarJW/5YcmImWa9Ikc6MqXQ0eVsJ4iK344P9bYwfABuQnOEiH7uHLGU
J+iVUljkmSew3DL2pIq6qq178/FngyKzPmOpq6E/GKoY9MRq4EhYSrQyNRGmJMALgfqu3zOXWlhe
WvZ2xZ9neBdR/46Lc4pegNnJiXC3f0aR/6OVdwuMPlDkHgofxi4X5By1/c1ws/e86Yd5+6rk5kNh
JaBfAfAw6LOBUQ8NYAG8IQwRnCtr0EZGx7S2hnvYY/CtFk/FlQpcVoPAUg22ai91u4hhCcTcDBVP
ogAPfvN+BkroQLW6MmvanEJZIcdM2rPy3B0HJy3jMYgnXWqfAp2oUF5d/mxLwdo94z6hD8YGNHGJ
z/oo+OnIEQdc9xb+eSr0FCWcMCUwR5r3XJ8hWLUxmFrRElFjzdURIXggitJyRJb9ZzgNJxKJtuG4
drlkjzKDrRx5lRfEGS4R8MvHP8+67DQUSYGUA0EjR7OASVRwDgBJNipZHQlgbSPGAghJJLi+Md2f
bONdo2z1c2W0vv6+VWQqyqfY+RfvhPfVbMZGvFioA2C0gGeSMHn7NgeL68jQtoS1PViOFl2SKvce
qv2mlIB5DF+m5O98bJhu9PXD0/qOL01n1XOlTN2qOc4oT9LU4yC7a+2eU3SX2yjJBWINDwY0Wd8/
e2Xg85B4nmvnvs34wb+Us9mwy4uk5lXA51iVK/tYaJkijGP2O56kBidfa6A/ny1eUqcJ8lXTgN38
IaTthmkA600VJ+NI2QJjJ1gqIBWURN1QSyr0abhKftn/fNiAeIUUqD6aiyfvGieoRRLzr/vmGird
Bu4+NCRzj7qUkj9Q8YxDkK+jEcGFZWG/6h4istRqOHCxooLIPCH5cA5azIoiHF12YBsIW1LBCCme
9mGcnKfEuD309ZwCj9m+Fqf1TNA+XOYLnUQDgexyBLsZC6DVgT/V7AvERDUzTCoE4Fw6n9PZa6wV
8ekmeYEyN2Xh3DlXQ/CWs64Ujgmmv205PHh5ai/YpbJu5JmOE7Fzbuf6PvW/dFfTI5tenDrd///X
CK4LzUVO8rwoWny10yQp9DPguTIk80BpjowFCrjueqMOwojFT7mxi6zuj30jdg3lKK3XvS/uhZ+U
m/ItPfw8jj0ZmVFAizf1xXyPv8Rb+g6PcsKKRkMCTafMPwvEHK0pfBxOuC1c3lDcL1trTcynOB3/
XLYRC5v41uBGlaLbUet/WK79+shEr+IdDXWHRxWBKxpf1sfaCV0IurD/HIrfWj1MEp8p6zxXbqhA
ZC1lil/k68KCCD+kGqm0ANcKfR2ef9AsvPoMjTR6S5SeYO36okfhnPWLLUCavnZ34G9W9oxRodTV
VigcGZJhl24Akuk4Vck40nP0mFHp6dGvFMF9f8O/MSMFE8snJCpeIHL4Gs0+Nj/nD1sHqY6H6sMO
vr8uAtRJAUHH+bXZnqz37kx1z2RgCL6ZO4MsrKtUUez6ZU6KUgLMfo3+Tz/x4CdbXv68TsQydg1c
JYPamQIyzaWY+f8D/Y5vMbK52GIi2Uai0M4YdKhmpz40RBFr65e6Q1MjREN5vrojWanbuszCsTLw
iuGaAWN3Vrv6lgsxxRNSXq8x2cjkR9G/QpGRdTENQXiCisgHC47SWURfphWDQiTuJL1v/0os/OTK
an+rgnDr2DcuF8F/Ux+RPDGq+w7MqxMUfht4w8vLLCsg/AEkwDF8Q14BdhDvNErQhHQJk+WmHRnL
AwXnNfM7E33J+u7gqdQZ25TWDIjxsA3i/PB4p3oFXCHaDxB9IHm4EdrK/uH8yERt0KKreiwIt8f7
MksU+Fvi1lilMIoDawizZ8JSQcxYbm2l1KdcF4lK7eFhPU94S7vZM2KW+KqPuHjNxi62gOU2+XY+
dy4VaCor7udQ2etqE6eorRe7hYVEIE2cJpQLGH1vc6AC9veavkZdrgiVktkCl5+KsFutTM1lS7Ma
hdxeMgt88rct10+vW7oDw+Rji7xdW2jIdveqPxBDseKOoUm/dpCuaikh9PcEHsljRIkIrxM2Npnh
1uSQHuLcCWQpa4FqoiVxOcdUyfAjOIwSC4aI1Z7myUDNcHt4GatV4cfUmSgaR3lwiDu1dYnNY3Rk
+FOmgMvU9fPe8Kzwdpb0ivekt4vIk8ui2NFXIdmngvorJS8F9n8K8dhEQRVzej3pSfpguaKFchcq
A8COW4ToQr83eCatmKcdBVf6XPZGBQrEL0MubWqdhdG7X3uKTDrb1uBcSbK9NWVkKADoo0YxCeBR
EkwxHcHjaMOM87Qw2BA1HOXT2Of3vt/bmV3Cru5c2eApWWHW61Z+CWpMItYL7RPLhB3dNz/P6MmE
wbMHKmu6LXCBO4NuLbyAhW/Wk1h2HFwrTzUS0fgyDoFsXxrsbVRZPYVcW6JEIe0CVE7f6tXy277H
+iss9n3m04tKFETnemThTwHl1EUEVvf4SC0jaZajdKugPT1IKjXsyXsq0BXcfcPXsp76w9/1bYjf
YVMkZPA4wPgXR3QcW840K2mFG95krJNRzmADDaHnRrjpbJ1Aoa+81mLzdF2rrE5kM004RLJcbMtQ
l2vxFmpBrJJGvsopgEMVpDSSYwEaGMbeDoc2T0fO+8R9PswYKuEtBtSjAxYaXr40aQWlmIR8WwLK
HfuJXxzDheb511Zj921+JSqWpC3bWs45RHQCCByWoQeSznFMO0hqxLoVw+RByi2aO6aLd4XLM3Gv
UwAxmqDNjwAfmRbwxuBvj959GQd3384LBc3UtvkDOLx3m5EtpkH/JucD0lk8ygUfJOIbL+LezGih
gUVUf7lOQzSsZMBw+d8RuJnVYKAzD2/xgA0P7tj+Q9NlkLA6PQYcjSd3ynl4ziTJDIqZ8aqCQNjo
QKBHn8rLGERT9i7JZbopeu6qthNVmQkFORj2G8NN4ryiNsAmIgYWIy23Vnk2ICCdJ4cOPXDZVCf2
oJbEQndUieh0XHwVOxan10d99pFFpolquHQGkPbhsfatgQR4IJvwgjD04JJWwyLWVMTycPnlKkwk
Zyf1MKanBMKUxzAbcjO3nw74kd4Y7TBwtwduDGA55GApmusnWYU4NqlC+NRbHPL7xPV/JoqjW6ok
xcr3mp1f5GgTOw8v/YhGLrCBfrkWOn04bPMoJpzVQJO1hjvOgpe+qhmCJKLgv2wbjNrrwohreLve
TiuRJOjZ2N7yhm8C0cOFr0aMp8FvSxc7PWVFh0qfxZ+N0/qOvK7g2FY857MNAOLWOknCQmxKhU7e
i56I4/mWmaN0yZk3z1xXNMK97wp0JkRfM/wDEOztuWTPDPYY8MMIW/uAMyJwX5FIxuM9Ue/9rHBZ
EVUdqD4ylNUnC+YVjpZcqUHFaJDR990nUIW3b6Gbf1wtkia5qf84MOSOr3det+Cr0A81T6lfGaWS
OA9c1ixy7ryjJe+JNrh1jt51COBxbZYUyrGFletAw+N4cjHd3fN8xlzVPTvH2ToMQDZSq6L8EIKT
V7ny+xDjmngemIYMFVAiPQKa31t0JK6DcmtJIiiM6DMnNkTWnosEnbAuXrkIhYO6opCur+Xk5qqE
6vljBXNU1GaftlCNLwJdEt4uFTn/ou+GI3z+1ofcM1xH9h8xUk7orSSL3RIsi7JdELoG9kq+DwSS
264g4Zr7ptjDlDlHGhvugrZlvxgnJREgSixwqaobQb6DT5YP98nNC9nWRsB7LJMEC7IUa7hHI1Bo
eCrC5C/VFdYotdxLY6Xk80uS4wv/kreisKX2uF1ksvuaW5Km+Ubyjg476Uq3gzJEwN6KRatgf/q2
/vLCp3uvU+DJJJVfGuUDOLO0lBlNh2PmecZfbgCvS3uR6vsFEWC9DFzXOYCzbIe9UPScPMEtKEpk
D3aBV28BcuLxh3ibkWt4FbK284bjLqafVWpT+jafGDY5q6FJC2EDMaRnj2QJ7wUF3cGe0vJLfKsR
L45pB4fySCmqdVOYQC0ObNyeROgUoeZNRASxPiKGZgUWjMmU/t2xE4UQUjd6BoC6A76RnGEpQIky
NS1zsD/3s6GNazaBWa9RsazIVWgasD9GPpXekrXPbR7UTC/8/cA7Tv5h5BhV90GmhZRm84S9VeO5
qShrmwgBKPDl565SW9VvLadWisjwZwlVs87wCriOYuSDbG5m4noKbCRh1g5Fr/dyeL1bWZFoWBnK
9Wcv48COoh3ERdS7oKhocW18KJsMxC73lBsj+1fyp3AOufFmEll0fQdNM+HmuGWme0UZVNs1Aw4c
tI5WWj9x9OOSgnLNisly2YmSlu5LthHpl+rPJUJ7Rwqy1Fkf9DAPtqiSgg1D+Nnqzv0yYun6Y4Rb
ei5tJyE7ZF4eph4YYUCbGy5aM3HOTJ3vzYMTjoHWaFkTHmeLv6Bt4l1jRGB0RJQewYt+xsuzVQT9
ClQLG7XdyAOnkqtqDjw8kSttTS9K2fw07JXKrNAT1fO06Ue68FXaXcO7K1kgt12X7C2Ph4oSO4bZ
CRGm6Gavu7K/XQYAdThaGdXXfV4CCuOHOx0PFiRLfxKabf38g+UMEPXQXkdlvBDQHGlXQuwOkcj7
6XGaWBkIy0f8cqhfznG5vfLgyvXzYLM7lnnc+rlynfTJICaeixVw2OMF5KU1lwsImQlb9Mex2oN3
40Puj2STAXE1Bc/Dlf03TjiCNzBRhgInNQC9JdExzaLkT5PHK7nmIQvK+X79FEr5EQfIioaAR/CD
SCNrq6MxlmbD6DeBfFo9PLueAljuquIr5hXvPDkZ4hEpNE5el7wEWgzcJqcVRh5nXpzRraQeCzBs
SAmi67UlNdEltfdy9Dsndd5r3vQFdyphbZW6lclDzphE+aJJu1NjqISCI0L/7Dd1bdkOpsp0cV5f
MXAxyVBtm4Cd/BprujNPsycvxAJxv/F8WrFmRxPoNdmqLJgyef25YrY9BkJpBmaqID2EEudg/H0o
3pPR7Fs/JQ9oaNCK00z0ZOYg9/K51xfYOJLttsGFtUNNxMugkbPzg6Hp1ZeTA5M728+NqeN2i2BN
wQMdUpeYP/5FmInIhZ0hC5dFN26j7uM804IBIwcIVq0lG3t4a3VouqwdoP89LEe5voUzTY1/KmEM
Z8yyimNoUd5M+cwQDagBwu5ny92ddSbZCsoCEvQRCIP8SMqwZ8efhpWJsLiK4G6dzWBScYinnV0F
I8qyAqZdgHb0AYiLxFLQ/tY0vdxTmu12Xq67RLKfl0IUsIDnK/oruI6il+qV+okKZxrAh1zwpT54
wdGf4B6rDhXz6pjuGg4zMK3ii9MU7TzYdfMrjiXY3KL4fhPgYZ+r9VanKN4uhrBz8iVyLTqx2iAe
SNLYo6qibC6HDVvIS4ZA0OEOciayAEpk2hw0otywlpSe5DCuwO6jmzcPZmpqyP703EhpsA8a1ONh
y5myew7BAmfdSscErs2mXYRC/Jeo0m3sz20UNOPLV1ojvTz0ZdvPtr2sheumSHmMfSOC3ly4eHZZ
917CZa/JOj1LnOIh5T5Pv5V86nCMenm71WVUHNSrQISgCpu3S0N2lyPnkzX+7rRrFEhYSH8fH3Zj
UyF2Dx2SYe0MeKabnyLNWacHgV+7DntX0jbPv6xO8e7tabcciNGx+PDcgdXCmA2pq7KtlqTkUAN4
I/OlLejFIxgA4xCqlmGQr/KtXt7XKWOWZauzjLO1udT8PZd7DzqY1LHgoxa3yFLv+jslRb7j+hfL
A0RHDAc2k85H7KbXNvjGvs6jWwqA37l5XPMmrZnFgSbhPVZ0HmtaXQm4EwEtX1uLn3QPMUhkWqMr
p9mHrnbOQWqwb7jnk6u4xyO8wis+2UVJ9xujgwyrvmRyYgWZzZ/YaQpZEI3qSpP6qBKMduzh+v/f
cf/Ub9iZ1ASJR1Q7/3IiPw6T7NgPQG5EmLJ9iMIptfhVzxKYbE2MNClK3gariClOFTV4awF7bi5c
DvQIxVoWHtAkKuGh//d5eMLKr7/mveJSRRY9ovEqkveQ86dpVdKbmG0F4wSmxs2KrtPfNmNdN52r
qobdLEVhlDjfS5hj6ZsigkWwy9qSz5PpHc4v8tNepFjhSR3nRG8t2AgPsE0XjtVO4M9i5yz+uty0
4MIPZVKKQfUlEpfU/Pp4DnAqqloJ/UIH732Y5XZqL4HXgu40jUb16nCPqRfxY5sNKJoUD10BcEvZ
qdtgw1GbGA0sLM7Chl5dcOohtcluX/sxuZXRjLrcV4P5usoKxkDe+KdKyhOiKHMPrFRHRfIf2KbX
kB18Sh9xJtr9rn0ImVszuESgKdsWRFFVLXJLHHmt8ayTZpJrZHU/fpwEPbWGj6QwP+UCDaVvOZr2
QqXYQoYzDw8YEHmMt1wa3gg94byzoeNhPLT9Txyk+UUfT8mXSYDmbvK9JqAf/OCaGz3BMgqZJYMg
ys3b82XIsxEIpk7eYkm48N1UJPrYW1OJ7jq1fbacEk9sSk93Vqx3/BSbmcpw897Log63Nqjvy0Ex
S/XqQkAzG7asnqs5UkOpN8DYqq4tzIGHvm+ARuJyG2dlhODGlV8x4KUL+aCsPbNAPBrCseFN/LpA
AivmeMXSS9th35VLBCydDII0dlS2ksjIAwgimLCWBRAZImTTwg1dLzH0/kNeF3osI/SjKkuCRgYE
ZOtullhXGOrrOkIThSpbLJu+QMwO23fJmIrRPiHI4AyFpa2iwP0EY3KKIGvh5eXON0LY/O2UDVyi
c0RYCFfEuj6wYGrgYfh2+tzygyijlW2WfA7X68flCQk2q3ERuMLO9xv2qPJvXhLulOv3vwjyEsWH
HTvE9MzxBMDNjeRUH2vM1uG6R1bQJNPztXgUcccx37DDhM2wjOG+cncLrQNmn7gx7XfrY9hspTy/
Zed2iYk6Crphp4Fxw8s6p7vu150PZk99zSLR1P1kPyvHt9c6LJIxLNxwh602og65BgjFntQK3GFe
gmPERz+TPjV5HEpV8zsgm/pqGpMWy0m054gnwbXJsUCA1ou786xrIoybn0rLoe+amrQHZwKajoVr
gZ4LnwJzvMthqcO8fgEVQOrKbDjlrZ3i8pHRjMEwDkjzu6jg4B/ymfsmVITrwCS9Hdd3+zVLiayQ
7OXX4idKEIrc6CEdcDhAHjRkhh/KNhXGy6YIXJxbD6rwugrjDXmcy28OZMTG37dDZSoOdkmrhHUH
rSkvOpG864xADMDk8S5jsB3pPpVdQWs16X4u7pRxSB46UNyDTOJf5/qOsF3FuMRVKvQKC3BBBWA0
Z4knG1rElLblZtotjwVLpt7g4uiERlu5zcdb9uqudzDpDkO0NtLP6v+WWWwdvMEC/WR4n18mIYwJ
/WZxys8oqQgzOlPgnG/huzF1z/L82NKaZVgoPf7okVVyCANg59OEaBQuTXzxA1HnbBlvHIZpg6I0
dpx3WT8vfQHNn8a97hk924EfyPXoN+88dml4WFh8EZdo7diTE1NJNY0B4mv1JUZVdEV2t9/o8Bf8
7FOOcjZwRxFWL6gOPD/8gD1brb9ApIRdb+G+J0rujlHZZ83W1YAVS2XUw6ovm/rNnaY4ZdNUPBSW
wH+2sBP9bsDGt1kpWHOADj95yDXdtCmWtcdRy9T5ZDHO8FTIszhfMePJKBi4FUKZbNyvygMifO4j
+PBHkLX9jtkQBO6lOwjYA32rknDHYn+MVAuoaTBHKRJO04+Z5ASPh7fFc2pqwb9X0Q5S/6ej+RYH
d9ciaKg8STJzEXI+cuNjbR8RIgRcam33twzPI+ww2sRiaW2d8m5N0Kmy5o/FLxH9NooQlklfDnrC
Jm78zdaeiiFZssthgAL2acZbacca89hxKU7wuSNqcLgjERXAzPH2glc24IxgRin4hncxY9p7WLUu
J8XL0JHeJ8LgQtDu1pWocfB3P+QCS9l8NUivTwsAitqRAD0g+n2Tzcs7ae3B25Zt+I0+nbf2Ksag
d8l/JFqqxudrw4NgUpzsFVc6VzQ8ndAjF2V5aee00ND4FAFWw8XjqICW6CfBBw7bX5bBW/6HY4sZ
7k+sNscwEw79UOEJNn8nqMW19A6eaEp4LP08O47w+Zh5VQQY9g/CPMYd9SrU/IyQEPNFyelDCM5B
WSLX6bPnhIoDzply0NXbfPrW5d7mR+CIp8pTUO9rBx7+ioaf4C5+RBRePfijouKmTA0LYK0oZOM2
CogzVmKQghiDXUk8/J5VPQIFRTforMKN1WYqr0JNV8MXJCyyWsFQyItnYw8vhinI7bbAMMKjS8r+
I+7MZCjZTHj6IDDRZ5QdFfu/jURW6wzdL0IJL44PH4IomW4orUX+iqC35SYAFDUMkagNeg+0ySjY
Gwqe6V6eYLcylg/Ayass+4GXOTtAMpcnRQ8KRSp554H+dcJWO3vVLso6uOcFdGNcrKBo4WEwWdxt
R+kwlncRseq02NzfnsyiDXm+ed7Q77MQwNLX23iYinlda6H+l6PWrTs5rvcFV0LsqBspG40T6ZxK
X7KM7RhzqZww4IXIZvyayhpnVuN/r5Wd9EtYAh3WVeO8UQ2MpgTzohn2UukX+weAcSegXjKLyw9m
JubFyatYMR5RG2DMZraUYxNOaqfTKbCBlOgIHa4Inp/3BQLhywoBg9Hh55ExWpiq7VJ04MKKqv9i
noXRZHKF3G7Li0Y+4RgDspvMFaWb/ytwlEcuAcXSksXq5yOEyTCAyadebWXDrjd0TEY/jhPi9j7o
J11vbuOyV/KteIQlyOFO5ihnT8Vs7I0RljcESXFqtQ40ssiBThGHbMEIFDK9fj1fJidA+735o3Q1
7h10RQCST/uAM77y9MxNoaux7axaqPxM4wdKsDfpN1yN29+28Trjslu7d8YuqzfgTEIPhbYW4ZaX
o7jB+fCYtmyBUFpGimVBMyX1uCEugTDHC7Hvde/F0rW6iIgbmju45R9u+N0mPrpkXweSgguGk/Zx
6mc7FEEGCVWtktMX1Vfa3B+nesN4iLIdfkkM0HCy1KPLEBLN/Y+iQy0qnKwX4lbeYZjhRSlt62zt
R3BaZU3kk68eJSc4yTNgVWgaEfAM39INOzPWXRTV59mBgs9oyMh0jF+bgoX0ZhdN0M9Tq/XRHT1A
yj7V1iC996B1KVhmKtrLKpGkJky+DXPZBJyiYDUFgdDofJrVOZduVwf3upSDc8if7Bfh4IM2AT4F
ibPeCVSAFUsjp3WaKgG8GI30HUlTCLP3u0YkI0Amum6uS1K+XiWreuzKds7LZPCD3nUZtMe6eU9O
NdJKX/G8asxwwzhSQvGEP+u+QMpWfEtFJOXGhm36XpMbMzQylnSxhi8KVkyt1kz/kKN0C9hIR4qd
+Mj8spADeLWFUN0AXBm91RpL9Sgub+aQWz18XAiHHlwdaIYJRNb6RDy8LXPEpCSrcTntbNFbsfWM
6hU69wHswZnyzBUy8rjta3/C18fV3SDUc8MqYJrOYY7FRUR4bJ9h4bc4FF5sPZiEsxAri6+tImGu
GKWwIy/Hu6tS85Ggl+8i2b1M2EySpwNcseoK1zCfwqMCmxS2UBHGH+CWsKtLbXtrPYNmjYRXbXVC
q3x3wK63Z/wxJCATaZFxjyUBDNfa8JP8p8lZe6o++EAspmqOKeJcHwBgEhdDPIpc0FAe/bc/+9K3
9tW6auswDP4QV2ZdWKqt3D9QAxct4FNw+jgqevzubVjhCXKffYSAIONJ7Mf0UQhD6EMKvF4I2+U3
Wrmqm+ACT5rZ5OnD8C/s1Z2BCUeqUEnhqc3uxF/3EZOc98SgL0PSnSasXES/JHNe+qSu+DS217T4
jHltNevIzKD3tPFFFlvM4111s5+oCXDaSRzDbcYk5QkaFr7Dc8SlDyADRGBGLM1XIFodB5ksBwR7
7mKf6KOKCXiebX5u28kznqY4PDpgUPh/7Vy7YhwLFSiAN4cokjEI8nV5AleLKqJvQ2KQ2QXzeckG
RSRp/Jwe4Pe5u0gJUUvBNaiO3VeiK5g8z6/CjIE0fs5GBexohAC1ktVTJ4evRSydm1GNnpFT7lwv
QWP69tGt5iY3MuhUCt8ZTTw9rHeecA7r5NI0Lj4o/0Jrm+jr3U54QHnypilfTRF/zr/WuKck3phE
W3arsMinW+Zxlydc0AljzKzIx/SaElOz6PklJ5bEovriWUlRbDjVdZYpNlgItul/fkzMvCZmiyI3
0CbTU9yyIj7S1N/Ny0w7d8BoVfh85rKReSanyCTX+hBLg5VUBKY09A+5mUIcgxb/3ViB3QLm2GVT
59bFl61hxMKpoPBXdBoy3ho96rKoulE8KwxEIW85ygGeOGjdkdToZRpK+lybi8uufaS3gaGx7K7A
hUPQ36uSj6VQ9ZY2voF+lgBGHuLTUhDVQpNwhCi2yWKESk8qWBHtl+nk7BfFY60kVBR6Lw8pwEmO
HHEqTIGJDwBnsHH6NyEEdUecfnKrnp5yORXjkPrKTNQF81Fs0vLBnGFRP3ONMDiwFxAwp5xgGEQf
HszRGV7Ez5K9dKPm1OPxhjP/TBmAt0NQhSWybW+hMydNjCZCPA7Y892CdTUMnyrEHPmwzGodWBDN
DkDXz8aVABA8iovU/H2tnf1RdvYs6A2Pfd9zM6fAbn8DNrqz5/ZB6zRJ0GqpLTb4MmyW7kkSxB4Q
ALFZh0vVF+5dah2yLD5BBF0pacq8hjHecSvX2wRW+cmKBBicEpR7uZOk6bBRzHmZDekpjh8yPvd0
cKN4YPoy312pznMntIUClZgWAq7otHDjYHLPtCvhOqjEmfg+w8h5cHoP71ja0AcrnEIyLqsnNUa5
CTLT98eWN/NsM4lBd4s302amroiOb8L4GEzhNUXTG705bUMn2OVAbQAnpreNiC0N3POtr8LD/KCH
B8zDbnVZtfYxPU0SusKkvD49Ht4oBHWuAiDm6zx+D8a8CtcHkIjYSbCC0r1oc+2hhXIq9k42Xhed
lZBTPaLVYE43CHhmO+CAysQg79vH4SBLlppbh8lOkmHv/AW2NRa67I5ppamQFCm4Dh4zhLT7QTym
bLeeIxKlCM02F4OOE5yW8EpWzbloUrlb9IkfReijXsRKtXlj1TM6V4UYuYBhSsG5u1tJoaDMfQkk
/LKfzAws9mrCJnNVMiJqlaMo1lgHKlJv9tRwm8NL3GpUxf3+FohooFDq+Bx840QiY+meKkAl6P2w
bff0G6sTftAsYwpwToVIKNyfNRHcUkvs+MXfyWbVJMV03qUkMZ4bPLW29vBqSvq+oFF/PvmftGzZ
BtkMMqdnBKM36+omk/FJP8cck4I+GF9/iELBfKwLKkJmyzJbxZLw3RWPB95lR8LmRUGcbYfyuF83
acNeq/QQcoKgc0eT7bdpzRRTIMFeJT/zK0jTCgdrPedZv3wOlljDWxQzJN63WAMEIp3IsJ5AJxYh
12tPUB8RIEokJNTeyoJsuXjJOqdaPTbvYmv40TFK24CAKQ8QruA/ZD5uRoVV27uw0iCALi9+gnlc
Xi3+rA+UHwyyCcNSx5pUDrUJWhbvQX5LxrYU/X1UiY/ALs7nVzNfXp0EaqcHgABKxnYdMuXW5F+u
lrOuHNogZhTBRUIBV1LAIVvb7AKlw6fKIUVdAlIP0Me672eNpkUK21CcrGMusCnRBnoX62ThiEGQ
mpXIStn+1mcUzFQXQafgtNbxfSE89bapX7SlIgvxf/rTc3EGwFw+cznwsUHWM667tP2ZkcFgnDZY
8i3LMmu2P4JEB7k7bhJlyHTjLWktsisIFDvhjaBRsMK+SLR84+hiouG86fnaS/SGiddHtRQFts1o
2cPFpZENwcD+fwJqSeH+OTNBTS9rd5lxSt6VyZbPlJxNifE9d0eORcz637S4yb1AiUqhDiiSQjNs
Oui2vUuzlKAmZjwT/Ks4S3fSaBo7v3LivWKn9MbGJq6exYuXUsFXMqlVk2y+JY42/J+zEbDipYRU
9agkweteOQ9qQnvy0Uavul1x0aZV9SCox5BWnCgjnz7fKRwFTTUhtnUBsECzD5Zl1EKL3bxFWOUT
xHydj1E+EAipE1QrXyEH374b9cmN9dEjYR3noumB9IheCeNO//AyGX3USYKToBTg+UN8Hrhrr+kp
613Gu9x4mB19bpgTFKfJYPTplwTUmM/Oh3SCI1P5DSDqmiLsknQqZ+YjwMRggBD53Q8Rf/CU/Fk/
lSc25PMm3DrppTff+QAs8o7BVxux0yiYecXUnd8oYZR0lT7NQ1AGxz8TJ5TaNXpQIZljn5DH4N0X
raMV7w9xsQXhGmWRS/DtQCP54Ck6uojeL3DWHUDQojmzfv/pIs/Ib0bDVt0w0GDHYx/okv5fD4DF
+2LhHMD3sQFNLWjuQ5LIB2AwkEQg3bHpRenfMf7qAOjKlVQ1dxO7i2Nir4LXwrC+Y6qeIChaWvOl
nOomQ14g1rhbyhnBOVU+GAd5BQKG4y4Y1ghx9mGeWTo8bH7LbvcZbdi1bFV8EQJ0+NpnE1n8R2HH
OpGhHCrdLn7e4d6rcCHE4jAVgPXKMr3sX/tmWnrpdutSQyoPyLoq9bYJpqFqTe9ZpvW3POjQq1bH
jsfZsreG/ms7uVwzUEIlhxfwdUj1yedvtucKdM+Rr8fZgvTzj7CEKkCiLG7UuwFbPzPkrYfPzEA0
t0JlwIVHkq1NS5BxWMCffnuYXKI3fM4ncjTxBcbTFhkw//0vggwyWJ61GlcDLJ/Cqj77p9prQAJH
r6ekSy9H6OilyARH8676uzUTD/vi2E9Zr8ivTl9qhpFxNhe4Dd3aaPMgKTrX5gF14u7Kt19cXdVB
EeujBBIXukbJ1rlCI6lkKL0GDjoFTZ6t1iEUAsiTvRqzF8c36psWn/jSgoLNoi7eQKgiOf5ykqHy
wookLt+B+f8sJu7KTifW/htXTmiLTDrXplRP0cSWG51yByHLe8dNGIPZasIrxXpvwy1VgQcjTUOI
eFd/2JJIr14xlpqUhThUolO407arIq3jEnMlYv8v4fhQSxkcjnk1JqbYJDGScpx9i6KV+QImCRog
ZwqINbGgYVaeeymnR5L2MTIFJsr4i+4jRiRWWZjoyGslVS6/XEoziTxiHSOWPvboaAZs1EKhH1x/
bjfSkWQ/YXkxb01t+KX7dwvTv93KL0THjrPsQrQs+LjcWsTzgSvJN7PT1SyQ7O8j2FeUGNXGbEVG
+qwSZ9/yAu9Th9Jy6t7S4SdraPt1dFtYLMDt3cB9jXFjbv3GHr6mLXLq7C1+lYCqWSXSE3VSGggK
uf2dZOP9Rwx/MzSJKLpnefBvfBPtg+iVKUpvg9xzGUmUgcJTj2vYcOKg2OoN3VKYmmFK/b1hS6NO
DQ+MGmgM5rFVo5LpN9JSVzbu/8LA9ab4nSpsvnVURP2VBppizMHfgRRKsWSUUnZd2qUjMaHkQLVp
6FdBCAl/+EFsHj8vmpPEK8X/h5q2+vfJ9BNJDVR8wjUxqS+hivZVe2S9VevpQoqcGfJWpWH7yveV
ldT1mNxirYh90zp2z1vbozDumrH+0zlYLG24PZ/P+Fdi32RCAyVPoTYmiM03ek6Ol6/qGSc+tRIO
xn4H3N/3dn9nMrUNJHgSZPEVS/v76sV7ehnlPGTW2Yte1+aOrsue0Xk2XG+wJLsXQb6jxmqN9gMK
6Coj4WcSuwXGYYm4HAh++4UpBJfejMttC6/ZochJgMhY/M2YQjLVLBGtIWYHWlx875r5w+Mp0QQY
pLuDYdg1hhvylRNTrDa7Nl297Hp/1PNQ3T+u73rxaK0EPq/a88bDTq3rHt8PPBN/gG/mjTYvk0T4
WnenFwxMI6dhtieabr2l2jOoAe1Qi3K6081LxoHGF6Vt9lOF1U3WacsIQ8RXbpC8lgEcBe8ywzab
mmbNaeAcfEutBzc2YSQsXuBD9iKppAymbj3PpODdO6NNIeF5M+YPKXP31kU/lFrgADY32LyDf5Xr
fJmf9e3NOp3STPrQYr9L78cwxmmsulnjAhYfyStybb6ky16MPSTvJ9MTGilVTzNFilnrgPPfDuje
ESHYxSoBTDnZHYmtaxDSl8DMGdi8ZYgB+KC72MG8wZkacf9xVIy7ARsi8pVQVwX+n98Wr2cHw4mN
j6fs65IMnsycZakNtUusgd+s7kezGhh2q9H+MKOSRs2m6QocTs1vzRXh8ooFda92SkeqdOo5YGuw
b+/H64skzbCoS1+dtExf05ZvS/4p4Gs4x8DX80QwGSz2KbQiPsWD1UhNIAkNh/B5nYXpmNi4tA7e
GVKNqgYFtTeO51/HVQo0ciWIgq9DRluoUJweUm8sg47K7CFL9+LfVDQ0M31fV749DN+MMJOPAH8i
ULCkVu4ngkfgcGvOHUxukN7dEYXvjbc8f/pBxmfjNrrTzvFCxL8Es3DxpJZRKWpxFVkVxP22xbsO
Y4XJrgCISz/VFYOnTp0vgpqphwpSBvOsrtjKz+lfWcdW9MUfMTRYBuAYOf1tzdDzH5P4IWLxR1EG
/I9+axuSf2NuOumOcaXKJ5vtBfzlk14zU3rhXLwutf9AwkdImjHI9dpu837mbR4nVcxoX9EP7TDS
GpAecm5XBFM55fDlCIqj1f9xsV/q5B+CJc+QUE4Zh3zkQ1NUHQgQAw4K87p7+BplJS2EdNMP1v2s
dKubSYEKIa05TG1gXjG88ZHoW5cd6mVJl80fb8avIwRt8Zy3Yhce3Hex7Gl03qYH1F/GrxrYtVNe
iyRRTpj4M9vnIExbU2amaSLVLJ2B8VCiT3gs1lW5vznTfpWbA/8Qfx4A3lw7+8O/sMAqx/KzT0Tn
3p2mioeDyaK9hHQo+V8J/CSkMWWWSFDR9fpQr9Tsordm8rSPqai704xkeqny8pqMqWAC2aJbyCmC
e52UIByJaOZRGC625zuhlPynkrZy74tmeSkiolmcMzSbE0/NpQ4+wFO3xQpNth9wDF2oAPjSCyaw
JTBLzFFtj87v1vtgOxh7Kgm3Z6++jlhXKV3qfHCjVMmHhvFn1eDPP4ZcpHrEl5zvF5kQCvIXFHAG
TlB9z7/6SuaP/ULWlfp5pfryRhnYVWgw8XcxxyoMF9OOVxe+Jdi/5KcT8W3ovvqUK/Gghhm5wgXB
MSy5NKT29FNkZEQKecRsgZFd9EMWYHnzgz3f80RefVnTL54kBoouVygHlX42S28Y7pvNkQQLCnjd
4qu+o0YwrEnUF1E8GNWfK1d2SNAWrU/SdxLf6a8MW6Xugpp3DUiD0Yz7kOS17nxDxyAgaUxVxsCK
lOzE4AL+rFgnsPmnhiwzEAupsAnJw6qx5UYOyTSxiPe1IOwSJcCcJth8k2GmKrngCv1FwukMy2Eu
KIFC7dAmAXOp23m8egtUZplttbIG/mRZi6MCBF6USo7XWHuV+gizygj8GMfN6EOCR2iWouoKP+GE
pbH/+QWtu5AzPbI8HbkJt1+HwZ93Kz81WUSIVQq79xDoPu/DcstYG2+PiRiF6Q3q02pa3zu0Ucea
sAfHigcEFkNcfCrQBUL4IamAwZwiTTbmMpPEPdl47WtPV0INXvh2KkuquIw8IrZfzLyozL1GfFMM
ecRKKTEih+QVXewBu6Goti2bvbXYFU9R5Z8xWMSDhX3/H3uEyJlLammtTiY5+9lfnP7NSHsU3Ya4
f98sZNlrgvakPuIJkrGD3hI0FWNzcBgIPfW1PjGcEZmKkIUuqjP4haIXziPz30rjnhHCmK3OtF9b
yDGpor9q4Pow+PQsX0VSNKWouNh0z5FCirT+AMKbfVA9s6EKhY5N42Gp3ENMR5rbPs1eci3+t7j8
y9Xh9gP866iwB4grIWuXbheD/Ul2E4Rd6+pKvVtDxOQmo0mOl0MwN5L/img0CyslfCQwZY2Yg6mO
lev/LtEEpUPDIWQyMa6BCJMe72bIuuHHb3spajNXA99mLn3CqELpFWd2t9d6qjR+ZSdSN1yreWEg
o63twZBfOIaiO94X/fZdx3iFTc5i7dbN7p7kRaesyDxUXdt7PwRQbNMbcjCGfJ2h23cYZhpOsY/Z
nMOROnpXlH3/vRQpFuBmQ64tBP0JEpxurvleoVTfEY26yxoxunITcyUGhLoLrmxJUiyDMLfRkuGu
Qpcwyky/DLh8+PQ6RjtHymJdLTO1SnQCCQvpvG0bL7RwLYDyCEwvSeLjzurbOT5+eyM8OvY25NCt
1axogRvHRXEHrms7bgOiNvamvdQEhIqm2k0GM2edwJSwao8jWkZffSkS6jFI7a/FGpLF//M4OaNd
hSh2748Qmn5k4XS6IUReaMi7o5/e4dVDCME9HzIHgcriAFSmo99U2FPoT3Ab7HUP9YYFyI9+QFN1
0qsKWZRQcPoNdouvv/0qMTqs4ykqhatMc/EW6rEHVWOXxjyEIiqcSbZSISWGOkB4xi4P5DbYzgRQ
Wq9m+B9yJDepQPo4fWeRaKsH1P7JcIhStOgaecF2ZQIzipVsM5hJ/Ydk4Z+tP1JM9iXJBIVfN4df
wwauF0v6mDlmiD9m4ySvooBaovnzZ+WnDs86iRzsxH/6vDGkBJWOgdr2/Pc+ukr3YXMH0FcCEi2v
XZYxUJuwWB/pTwM5gcMgXgywVHt4XEnJ4Fo3ho9VqLT9kLbDv/NYDq8CIhnhrubONi2op+uYwlpB
IZ4qY9M7DdQy5Kc6ueuvWEN9BO10ww3/0OO/9K+mzpaJ1u6BaXpVSm4VJ7BfKV7jc5XSmZGGCtCk
c1FTt1aGHLx8WoF5/quv9xy8FURvU6aVn8GGKCLaS3bASTSZdbe71gjQpsdhCoDP/D6BI5f0Sykz
YUXi0WX0L/hOG7K9WAQIYw/asvn5ioh3KHFqj+A1Qhk6K034NePXHBQiG+X+LfmW6IE1LpJqRhpf
4LUUAAMnxB8sCuXsOXNIsz7tUnnMJ81yPSoXArzRg8EQxfGBbQsV0wj6+/naxTNlXpGVmzhAu+0K
idr/VlRBpktk92VuPREQzwCwh3+XQ2iLkxNxL4vk+y+6Cp57lpZJ56UAz08ei+Vv2MoEcknps/NK
EssaPYGQ3ZUcFZD25waNMzphJVA5RiWm4Ex+La5bpsyhwSkWzyfHArN55doX5HIZLOQF0HQNCj7r
gbhhPpAK4K+UTv0A03LETSND8VvMFb0aBVyE+Cf+iZtgJMKVNZEywMwdUESuR6mmu5iSxBBsRHCj
PYuCO/yd6sO/gbkR5vzDOfMtzhE2capZUwytUyTIBfe+RmxMGQNglzLrj6mxaORu7na2MLVypCwG
3NrGSU+Z8smrn6q9fKYlUWX4jlt6coQUh5DU7oSQu/Kbq8maWW8b3YSSU8OHidpO8FI6E22EVviI
ZoxjdbdJHdcV/uYaOtagUdTQ8so4dE3HwVDXN9HF7DHU3tnkvouvC06EwRsc94IaLYvjQvaa1mCe
d90jrdVTbT+l4E8Z3zBXchdMteYOemrkzbtWwOSHOsNrTkaOmnlNQ39JdQt7T6g4vH4NxD/m/zlN
W69io0DW2zgM3YvYwLFa1O7y+im9qoHGw8aa9oanosnIXXeSK1qzdxvFwXnI/LiODv5RENnYHW2G
x24pPR8wqjZGTAyeCs91588GRe4IKgui7lnwj4VkEjWGwRc1YVHS3i52x+gSc2+ZJD/v7tai8v6P
OMs/ArPke/NqEON35XRmwnhlJ+ks/ZIgl3ATuRAu+YUAEQxf+MUwffU9iNgwD7bg2daSQTNXOrFv
oWDUot+wwyAtgiZ+PpbFSqB4Zd0T/WFj/Fy4/rQGGnSo/N/rnbN+woKR/C2qhsHI1caNbm+T4CPT
X5cRqrLmDtSAxdLD8um54Kbd8h2zFZZaUbAiLZMSRkWnMyck8ZeJSJvf0WhdUcqRu9i39T/nw2TY
Cbk6SgU0RAbaiLn2ZZt1WMYr4KB4ElUUvPfP8RdZoCdulaU/6HmW3V9iNhJwqufRVQqePMrV3A9q
Q98VSn3VMw//ZKdtA+looXf7gLXnRvd3GKe35WyEdC2KlHOkShB1Isu9tqzpUyRpuAXlTIbkLznm
WQdKq2DtIEkJqFuvu8yiUMbFDg5cMDN1iK16OxBNrfEhB8LEQsmYWuVuybz9IgWUGukoJgBgSMd6
cCjIWcs5oMkQ5VGlwuSU5zwHSNhB/3Gx+dTXT7CrrlCIBPJJHy1E8ZJeY4QJ9xNrTu0Ni+OtOcVv
BjiJWkolu1N+zQ8EZc9CIClFa5fxZw7J7xmsL6Cab6fEoA2d+ye0MqUzW3nk0LpYhkbNxdwoQoK0
3VV4HCdikCB5thSp8L59WRWgPJiyPZv/u8kG6+wIdVYd3w5L+LsXeiQk2BK6SgieDBSh4mzrKi0v
nK3OFmOiGGX0KwsTbYtuWKE0nYcY5u0c/u5e7/73u8hbO7cZ9AXdapu7vDMzpsIcvA2O38yO79xm
e33rHUXawgcBnvK8Ra5tk/jGsWwEPIJE5C88GSU2niLjTmcV0P416MoVZjbjg53KIdmjXkh2U5X1
JSREEv/N70sotkWVakZDd+zUsGA7/7NDIuW3HclgB+2ZGUKRgK0zfmI7tNuMhJU3C/efknotWDhP
sCXiGgfGigUY1cK9nOnlBVq+h5WYF7M/5HzZG9TQYVVPRaW02tAWAIjnjuKIM31lXNPvRF6YByzG
v3QilHsV7ebyChJToRSeU6XOaCaUMUaIXOrL9pZ9ZkaA9fLfwSgnZ3docjm5w/HtNOGS2JfiWuez
LIp6ITAvHk1tzottj5p7QmqqrJL2U/I9MzOrJxk2SzeqJkHkRtUdOkz6bmD/BVsG/mprrQ3Gk/TD
CC2YszIzqX7KMAqD2pI/XUgmwCEV+I08DeFDBbkgdkbw+fn3aE4DOogp7StrNz0S/qAf8/LIJoB/
bYDiJsMxiHPXXX914qfsu3jBs/XVSyHUf/iUQafp7ScqfJeZoWjYnvc+YPNZwOrhajPlV73XZewT
n4Ri3Ph1ltC4afymT2pY8+OkSrDqr0ZLYKgv2uv1d5K/vYlXoyCaT27soP6yHamG98qRm7szgeZb
7vKcd+xCwyHVDd1wCNmky1NHHk+pg14z84McTplc71znyjw2nzmD6pY9Jwcw1LlTLA6G7dBdOZhp
MMy4Oio2iBiN8bJmP8o8BefyVPfDRe0aNdAVCKZFfRleuvKxFqWKZiJ2Q1DuhPx4bIAQZeo3yixq
Krnh4EXEDKqjSbPw3THgmkjpE+Z6cdTyEy7S9OUCNNsqh8nLzHsay9PDvWfQnZVEJpqUnAehzSLE
6/Llcw6TEzO7S7OSD6j8TzXTYE7mktTcWoKzStOcsFINSqvW1scZdWSg86dIKAk4Z80+SM+iG6J4
2WL6ldN8DcoRcADJYPwCloWX1IFEmv0AVX4I1Iev0bIq4/nJUHQS0T1P71NNjaWqjLv0YbNyzShk
LjMHaegJrfLPHC99wpGfWOIsf47YFBF25os83zJK745YKkmeLyzhrRHC1XWFH8L6frQavbzLkpQs
dC1ovcZ1mADJUtPAtf63D6+wsW6jLc1Z3PntDMcn9HNoDjq0IgGDOKwTty7HndXSD9W7/0ZqM3se
i9nKYoslW7BOE3StYwWmdZJ9lXkLiQsmTQV+M9LiFlQACPnAA+wLlytF64FkTAdh2BptEolmpMUg
uBYiC9KWygtHpBz2UFWBZ3FvhxngWDgbm2VsQ1E42wWpHRJsPnRckfQUDGgSS6DffM4Ur0ALNnaw
dEOvmZiBP71b+M+DYu4A/B9jsEK6biT9Dj6bhg//pYPnYOuzRts3dlLSZjipElo6Ddxs6WUUY1TM
DqJLtfqzbXPdeigrkqY85OvBomloQUPuW5VhELFBLktMdPyDcv5GVkQAUkuJzqSO2JyXwMQ/hS6W
WA5nM6kVa3VR2gSW157faE85k4EuCon20Cvg2425Cx5F3etxXsNKDRO5eLVBUxu6WJt8bjxoOs4u
BqscjJaqlYbFlvP5U4TYevMaWOF0txlHLRbU90Z0AsNjAO5+c3asmG5jSECvv6NK0tXD92uHePJq
Vt6xGso3yolhzltCoFtNApTtdL3Q/mFKBwRXz3e5UlwviHRSnNIIOfhWbaK6kN+yC8SFvcqeB5XD
PWXhge0KmjCQCgK8Itg97gnKtcMfQEyAbMsl+I0erD2UeYD+tKgsIjTuA503MFUjlAk2JxI6sW78
DdJiLrp9Mmq5L4lUG5R/93mDfYCkQsHTqb3JfSBxvTQrX0/B6E3th/yHf7lDl7MyUx1pdBqQNznk
NWlQq6wBBQB3e/9aY6TcLEF45ygsubia/S2ARee0Q+dqD6NcqhOxzyGeSBIGSJgmIqQTFLt/PRwC
Xaq15UcnQlaCRZoeR0GM/hmFbWbvdfzoF0PMFNer7GQsOoGwK+CZd5MJp25LKsPfL8ZvEuQbe3Vg
dF2EoNq2lLmFsJo6kh9Jw2/OYFLxmlG6+MUKPmV9WANvVYaC4nrOOBcJTjsJMBOpLeTxELPT11nD
gqUjm5GSDyqBKYtG9WjhwQj1GWAsWM+KyURS9k7mHd8POy+erFv9U2VBJMFMwcKamEf4hA/EO95I
YKatbFonL4jq5Q2DjSdWzy2NFrT99fepTM8g/a6SgbR8lhqj2zBYPMfKtHJDMPxV8MnEUCsw8tdv
+oMn2xGW3UcJAmhvD/JUXHTz7aWMa1EfW64cHeJyq+NlKudPT/XdpLnUgjZeP2VSIMu43GgCd2gq
0XSo2tCnmB3y3Bl7+41/fUnP/JkDmWf2gDE4z+i22NR0BO6cwgtTrGqrQR+EjJdWVSi7u7UGnzw+
DlVIMmfG3gvRxqCdZCou0rkWk5lLFMys5pLs9OZ74l0yIqZ0Xn2bpdId4s141GTr9Sa2nN515Xvq
7YzwNJjfLAMAlIqus3KsUPi3P+HTa2XdO6vOFQV+8WZWUtZ60EhPowm4HcFVUiruFGzNu/0WVHDN
Bop8VztS0XcCkHfiMo+iqlSmf/OMWMVWO8fgeC8y8b6p4/9ExISBge1PPYlUpQ1mFwzp0/P/dJN9
1vGfllwZlqTSko0XheCHtYnnw4vb3v4T/XjY+0Nzic/saD309gwM48VkRnNm7QWRCrRIJwzrKRTi
tNJxlzQKDHv5GjByPD/rjIAEe+8MGALqiVXYyq1d7Wpskf7Z6nJC8YdkCUckFq5DrE4e7IuijUiT
xXcVUbCB+Y/cpAVXamAjhOzJa1UmZ1Gl+CQcgjavFAD1MudxFeWm4M3TZ/2xL/ErOtSI3tmav3sb
Y6sj2vP/XB0wsUbM/g2RRfrAFZWWX4gH/omX34SfuYROf4XZQ8FY35ERL7JrPPb8KzfprF9KNJW+
b+CKWE64UwV84TgsmQSv/8WUvwaClim4A34ygIisGg7nebGAWhvD6eyGLaLWDoSEfZaO6RWgpcoE
89sgQTeyWFWojaLhYphnK1H5XFq95tz7TrtZ1ylnbDdxe9YUzENWxAWAWdHS8JspC03lZWxnC1/M
5bkzCU2HVHO/MAov2bsGm2sUydegZjtsMsB64xOAnknTjCE8GXEoraxhfzjhyBoloWNGBz635Lxd
z49+WFgTXyqkhLtRBc6Xh9XrCpj9yDarKTAl8qaDlse5h3bruZ5Qn+cP97Xvj/Fl+FljTcJzltW1
5ajHVo/cngkaUuvQLx5AXSkTPlpfAe1/s/pizzV66R9p3+N6ybr18eS+VLf7Qy/BeEz0RGJZYAYo
EIw68moj9QnXH+xfcNKRO0ThP2t2eUAoIiTmhSAUhmBE+JfOpYNv3A2rYatQPUsLV97qBJplfcvH
LUjV84WaLKEEBDQ4NXoqiiANJFb1UEpsVeH8Vd6Lm/YV8v+7gXOSwbvGQ1kmrbppKvtMMSiBtbzd
TWxhM9n/V8Ysa7jMc329VX+3mfFuCpW7N0ovxYK84GQ19XtxkfMspIpljO2H6xrNWLL9g4+TMWsA
gqGjbSe9EdKs9V8SNkn7CmOADHRNm58Fqr84w8msJ/CnkZhoEF6MeMKCbRPufaop6K21YHAwVtcG
w0umXdQolLjRRWL2PrKCmtVvcrmXO7vsTIqtEzAN0Ktb3zMCwOmHeuFJRB60BdjVls+3N8nJ9ubr
v6Ogf49UbdUoa+QxiWOAXqmLuMoZmcH3EFf5IimqE8N72nIhKJqDDQYl9aCOU9nLBoqJnjOLYc9l
Y501yOe4Olu241uq6b1GGG7EDNAz3XYoAmiJTmcRO43UEViQ3RFBhryWESjEjWhIkp6H7lAfX3/Z
1Ykgw6baf/AZqHeyEsl6fTpOWyhMKFCmDkHBMKL/Q7jDnEP52Z09kxPupzXQRuDKMDm/1i5wyLNp
SpRxqM/GW8/OquYNAGVOEyQFDQDt2hNfeaM/382a3Ni2UZPiNhlgYYdIMCZurDWri8asaPWbcxDH
mWsfDp5065G/KxlUVd4/8ND2Fst9xUGz8WsL8SbtdyqoE7Ofi0qXyxSG6+Pz/OB9Z4RK6ZieHb/H
rfzfmhj536OUiKT1+xboBcbNHJ7bFyMKyACENna4dxx2GxPpMXn9KST/uC6L0NPEF8W3FKs1J9vS
pZNyB/JVD/xpWXFjd3eNd8EEa3LCRY0imB+RuEmJ928PrQNW0+HV9AIofx6ugjwjNO7OPbWmh9A6
Tz5y8+wbQmGM3rj172qw9WgYQsBSTk0qsxteAaHfqKUW+n4TBADA5sMl61z3+cINdJzHrvxwUj62
oktTPcpw3HS6FUSyv175i5wQ2y6ebnOjt1A0r6fB/Lg2KJoWyPXhqAYcfE4wdOvMqaMvwob6PwoZ
TlFdq3YL3mk9gRoEL1e9Ra7RTQAxNf8dMIafgyodmeXu0syEHLXOoQT+nIN9WN8BOhKw1VPQ873D
F+iaYfOq8yl0lFgkG7k5OWb35XrlSSI/2eooFhL1S6dRi09mltOxReJJHZ8O+IbGzQiyIjv0RTxn
GZE+V8HB/mBz29gDSPh9te5sa55+odXsPCaJjjly0sqbuAT9NY53FwP9TWq5A18RJmzzNs4fLKq7
0o4vCfiUbQrOLzxhZsZx30bkE6LDbd86zNHhXs5gZ+IZncrdHYKyx46W9hQewp1ZEz2rjzeQRSMr
b1GI3wqH9LOBPJ7ryRzHI8LIGebyb/sa9kD1X5zMvidaumXB2cqipt+UWMtFkjGKGq0ZqNeQ8Igd
TnFpAA6Hhy42VHLIa81rQfeVrD0cSmlHG1wbEDfMIY28kGK/vx+tQ/An5NPQP0q+zkbiQnguLCyf
Qtg3Zfd+n+jgZp8JV0O/3TFK5rAWpayieBEj4o/Akno7bdlxuhiz6YZfQwaI0fYcINJXXi4BoNkq
H631CEJGhwuB3Uu67cgfyCsUOwV1e4zqzVkVv3CL7m1mQjDLwqwWfexJMqQtwPxJAcbnePtXdfXe
bBEIisbbBad8juOfT3kgMUVE1ZDvgIzs12o3lD62y+jbDj2RwiMTdn7nGZhbykWo/QALWWyD900U
jy+fPSDPY9sTMZwJAp841D+qnPbDARmwaQrLtjY1IB4gk/c6ZR1OG5Z/OyGZFcBMyYmxHsFHbcrz
eFGmPF3JZ6a9fmIeN33LVA1NigBoZHfdoWIKiZ7OLBIImoaBBXd9OXt6TkuYMsNiW8q3VrkE2F5M
aIPqYt9864WYM/Yp5Oh9YTJ/gRfZF0DDXlok7ZJ6h6qu1BV3ofzjST/mnYaLThsC6SdQ258mOnZ9
DyWWuy+trGeaxy2eYqBrkAGnV+/zRFkYP1O5V89Xu4oGLUs5TuQs0DW1E47ggIrhGrG3gpbOyZUK
NYiJpcjsd3mndMFqjna03JQ+6CmMWTctpGQsruXepVvAN3ol3hmhOi3zfIcI/xAuUwsBLHFIl2Bi
d1n4JVxWsGU7mmGRvKSe7UmoSvXMUKQWYigEyCIB4S6OtQ9fvkzwhPh7sl1gp7ck+Rzahj91yAyz
W4wU6bXH1ftq4PlBZCGg+XvF7j2257m1Eo+jbFeMM2/dN2eUMUh8z7JI7iQogQwwKJaFFFPWdcGO
tUBN7YEdSUy/nEZMQ94CkRVbbk7Uhb/Ij0dKy7Ego4abdkBDLx2cwmuGO1CyKuDE6ybcZOvdFS7f
ccBK0vzYCBub6pQXoMKFahVgWpP9v5GSNzB9sFYKStj5jvQu6tvsPf7zSKXTOzdmdXn89c/bmnHs
o3ke+i9hpUZnkXuw/U6qxYG5qxKg/DJc8Mz6v5p4LMyl+oLNYG8Iy8xAt6GE4pJ2bm61AV8O6CKb
tiLI6ItPXl16XYHjhFvjrqtNHGNvZuOCaRjbQqm/hSb3aEuVrEJ2DYpyS3klBbKBlZjf5TwVEjGN
k3aJcrQFtmguLda6zq/jgO/B4AieV5gYfiFw/ogJgL8PllMB0Pjpga6gRQg2cMebRbPsW9kQa67d
pVvgsxgKy/5Y8g+GiQ8pUFktJUgovkmgmacl8KQxeYMcpBujs3xLLLYmCL/ljugGsikswxRlGjCr
qMx10ipkLAhXCt4+utc4qPrqnXeULEXs16K/oykZu0VXe1Tpytz1xFxPurZt7fe4J0Wd70y4dwHx
yYgqgfjY9w+Mssl3tj/iwySIiagzlpknYCHVD4NcK32LsVcDZOnGnubirtQBek/IvditwnzInX+P
mkzQVq2Q7ufFxZ3YFx6B6GYpvx5kmpAoZdiJ0CKr5DQEHkgzJ87O5MxHjXqFPAibCukjcq2l4dso
UEyCfmWLwgItXGX8dDCzpyFZLvuAu9DXvFKZJywsErlgp7Trv9CH6MaWCqOhkzYMkBU6s7lfeIEC
5HjGp9QsDDCaXqG0UTs9DSkcGQDEyHt3ciIzT42VKF2bUkYjybt7WWs8QBbRnhYEVKe4j39iRdRF
4W1GG2mMQB0qWB9mka5kLFPKTMyqxdY+lFxcWe0x7tMYc0mpu0bCk14l+YM0SUh4CAuf1pCiMAWA
y4UVBP/ZRjHJrvjmCBify/0JGkD3hGlGs1F6PdKs0oG8b5QNFifLXovg68r/wy4gsLumZKxxj3Qz
JeBTXhEE0qNUPH8h9fV1yp8UChmJgh620cuqK+4fLmHT2WpsImousCWXTviA0R7SSi1KM2MSKepw
UoiCjcxcfsGga40j2jpPInBjC/x3qKFo19jAxh7J2Y/7Kb8ENC0ILZ4Y4f3gMZI/RIrHthU7WdDm
tzNVlXKErNyOGmdDM29VIVmaek+tA4cu3JNgKobwlQwYva7agr1FQska4fHDTcsCLLql7/H/QnYZ
HoNOfE2sKA80/6jvFnULiPaUjs1LEF+0aUwdr+T9x/rmRPhUWxroxnE3IzfnmGBTDZkBeqn2MzAM
/KuDXhpHNBnX7Kh5WY9qXjpQwkU/VRHh3kJn/PtP1c4YcdQtkmhkrkFKC1IF++w+brjVaegLMbL1
J+tQ/Yij0j6wgdgIomoGvZMUcp954UHSMsWscKL0bwWoU5GrEl2kanvSQRTt+hOSaEvzt8eBHhKk
hVK/N5GB1CMxBc9yE7ejGvGOvvYNADJTPO0mv4eEO9s/ypX1+HPlYu7iugwbwgwNModdUGXElGnP
F6WSOcyxnUK2Q0kb/Ms6Xlq6C6Q6DDhFF1BkyrjmHiXbJq5ch+wXLUpBDa8BZEHkNWwM9Ta2JISJ
a3ouG4kNWlaNxBB/DSl3sKIHO0NjeQkkN1NDVrsSQNe1QGHSdLTS7Ug67qc2xADqR1V0274jbAzV
2kT1Kd8s49V0b6iVIcNKsGG9VZxfLAofZ00glRmgGDB0f79zG2fpSZQ3xP9vqP7y93XVoinymyc1
JpHAN1T6tycDjrFLOhOYsYPEP64Y03feGwbAo2cC2qz6ZM/O4JDXSQLS57/h09z3W2QCXY3rblax
ZgGFJxEiRyxXph2pJNz+63Q0uM6lsX9nN4YHNuwihR2rXNOz8MedRs4o4GmeZHxUgVjZnD9Z27+W
IaYBpNOwJzk/HfsSL6eIxhsAqTkoAbLZYQMgefkJMlbUE3YGFzJB2VqTpwC/knrvxbN6q+8bEIx1
xQgnKRqc9mFIaVNwbvrMgVHTyNOVLoRsYWWO54pVxLUiVMoyl+z2QAKwksg1dm9avrNG9EzEKqK0
tcnz8F8gT6l4luJ9h+EUJEeFr/T5vb6aeqElzLPtd9DhJ6ksaDg6eJS40g53uGR7RwbhvQGMeEyZ
Z+eKucGl+u0jxFdr9m80CTd5a1TBz8yubgQSX7NZ91TcQl/6jCfLUfcn0TtJrpBagTC0fBJZtYKH
YPCGgvPCFKjmKUYAii23knEn6piRExEKEF4rYZ7/FUJkZu+O4i8Lw3JruptBylLkO5s/g4r7TRpt
up0czo9a2aKOIzGVWVHZRjCOzNrMZXcGRhdKSi6ns9itMQtiVZSHZqKQV5HQ/++JpjE/pJA5CKSv
uJ5oKBJdzbL80V55lvaSblJyVIjawP0/3AdbWqh9fFh6X1mWEpFfV1cHZvwPnefgezsupiYNWQEi
4BiAeZS9n6qW40Gu1K6uvmK5HauULCvvQ//GqnRDN0zA8wG16mHomkRy4BpgYD436JwQavm1X1JK
lGFOgDanpQDW/JT1HBqDq00JKbm+FEv2K76ssdzEdAjBhMGRT3YeQZixQ0tXXZoR33hiZPwMmw1X
ovlU0BwDF2jG/Y33P0ov0OhUo5m8dXFEoTuN5uRHoMwjylbUbdZ5APzPg7AJ94EuGu+F2WP8RfVc
ErTjEhMMETHKP9R9i7P4jNhjVLGK98RVgd8NeMb1x8bjllJlfpK/pSuMmGWdqr1JSaqO4LjYZFLm
b4YacSM5S5o058dImQncUxxNVSWi+8ZYDmfXgPnwE8HwPc4h+dU7BzXXdshHMIbX1ySdDkhtRQJO
iaxF3XB/67ecK0/IHp019ij0OkDtULzMf5mmBu2DyURg8EfYol5481CBXQ97R4A87zH2d9I8gbPh
F8fBLHt1iDbLzf1H5sv4vrK9prz/8BRCw60dwrtjRnrk2fG1AzCkYbpANvch6SWrTDfWhR3fXHRX
5p4+00PUfTis+oN+3xL5tcFR8AAAtsKCHLfsuvMDM92Ua2BGw6baa6isMBkVcfQkyYj0lvz0h2SK
rH43aEPTyRSMpGOQQSTsS/OYCae7v1ethjhZHU/3kRfCIKVwYv7mxvcDdFlr2oG4JeAwQ2HsQ1Sx
geSyJU4+04t6k36gVdYfnZ8lq42NsZuYZYxzDI0fOlFqEKo9j10U69YMOiOe4QhAb8f/5reKLxMw
ciJYolLG3Y7MpLLdJOhqzdzj34EwGTdlxdqJirXAc3+6+4dHbusFc4y2o7xBlEui5B3RMUF4a+/P
UCtrA1xaXL4LRwxByiIdwxK4h/KS1LvJiyfEkDH6r3/Lmc6qhu0OsiGz00ci5CzS5Gtofce8Qoah
1Y+47yf8L4UwfFIPTllJYAkSl0jyn84MzjQabwbjb/vDmV8/j5jBk4DNRBaoeI0mpxwEuefKGAk4
0F7IiP1yf11dPS63uQoVEUJIUKbRpTBtRMH7yCYIgLwB366kUW7pf5gKR6rE9SEzJuKqKXyp8YZR
7yNR8B5K5Gx0XXYRPJBpDeYS4GkqjwK7+nO2e1L8WyGwkhNZ51FpJPBkfDklzD9LDFNjA4QWeh9Z
LFqwmjY1rUP4mSPT+SnV1S3QdcYl/USGUi8Sk+6v2r4kdS1sOE6MjUHJ8M5PhNOAomJaL6YexEMp
avcmsUDdUYtPy/EgfQSnZGOSRDJ8dPIL96UO1uS+5dQBTCo/9h5GNJG44eEbmFIjRKd9ntGEejkq
/noBZqrps9iylwVUPfMXCYFvJzVhFCYdZZf7YDWPYE5N8SdgdV/nYIzrGEdAgvglyOQNXK6F9cbG
vV4UFA5Nkg8H/IyxvcJzOlshTxnnABs3FONSZ4njeqgw5b2WE3uD9B9gcZuXBUdQIPGa/8V2kW0r
BRcaDhdz0FtWWgnW2hb5t9Kv+am0BUJIDLVtBFO3ALS7oTS1YHAycX7gYql7kBiuE6PSNvWI9qIX
N3xfRZIzs5abPDkP6YnUhUkm9narB21c+jQ6/jvrNjCbKr/CzZErhcF1SEjRWwsVdYzcfNgrhlxs
qlmNZ2Sc9SKysadVsyuEKH5DKHMksr9JK2ffwex0akLsLY+Aj4g9i6jW/4kGEK9gCsHJHggeGaz1
s21OGg3HsEfbejgAeFYq3JMfVAXUHW2Es4aloUZYCkocVXxsq/oMe+CrvtzNeY1Z2macJ28ljNPH
0gHI9vblqs7mv93N5bfDuok2pSQU5zWYR7V6wkOPtocFxbz33Bke8b2nkNi+rYukXwSaez+wAtr1
eGTLK6RXNqhVZlDM5Z8s9caDMOTQ2FFk3dzDfHHmKTzCD3gHZgIy+JxBgi/QzTwE0N2Sa8mln7kz
MYt6oH667PJVW7WyaiAQ5GLqHq57XONTgWpgtjh1tWsL+9BE07mA4ozIGxz/4I+azvhcxYDOcmfv
TwUz2ltFJq0/RGnadaS78iKS3BPNWrntcpEeZ1Y84V5HnoE9qQtT5MqHsi3ZVuxtIros/hx5Csh+
CGkKH/XQUPDur43JcMag/2euI5FuJsPDJUEmR3cfltYdWX+SVPRCV7M8cXRPiEwFFqOtcroChN0k
CzXA2968vG9diXwzfdSZtaJG4LgVJbneW9qno9og/1VptxMdPxDX4QN72XaZc3Uva/SKM4Cf9YdU
GxaIMQjklPzVcjZshIdT4mu8ZAxukuEq4wFIm0Iypsg3k0CbNBGUWaAZ5FHGcKq3gG3Dx0A+xc+S
YZquQkQ9kTDxUY0qg/Q86odp4asiIc+s+icW8hBeV9abTJCBIoJl0VCzODoworsNugHfrG1iCNEU
OVhiYQpwzXGG2tyiB09S8ZZJ+KA88iXPpmOnCEi7MnpJb+zQDMmxHQe812FhCdCeQTbL1QiOpOkP
a7p4W0gQFCQaDY1T1JgyFyYB6NBZVT5BECzvheERg0b3iqX3lxnuhQ4dlknAcAqD5kVfeVfKzU4T
GAU7LbSZAINEAOkO2dZGKrmPxix0i/KhQJxEQaiH2xZ3+ZSq0fbvcQo7tZHUtNRs++TjE2HxL+bo
W0P+5cOc2B51ruQYEOn2ObziLEmq6FT9qbKpg7p9bIX69Lo6mtCua1a9VOVD8PIQdK4nWB5P5LiZ
UOk4czOHpbpsk3EQl0bVAXHYJ09n2p7hhZFgnWGfRKHXRhCmCOH3WAJwWUlcAzH8qNDXu7o+n2po
LC3iKapB1/T/4McvYpT4cwcdLIrWvFciq7tCauNmm+GDEM35uC2up3lMY/1wej04V3ECsztrBQUa
GaakxB0M4HDXkN5Mue8jC/X+Vrs20ZUkqW8eIdEAXctGPATAEEjht35WngbSVbxWCOBbNvX+6GSw
DfSkBGJL4qrYSlxZfKoY/sSk1cyBlqe0RXJKhMd6uhjuTYiFZmcV6Lxk1o29Sj/n8Zx0pOnTr8Yt
g3+UIQjq9ffWM7/HFi9LkfeLXdlhT54mYqrkF4vTMs5Hl4E+DZrwYLhKwUMDMe+1BgAE7WEkXyZU
jdZ62EkveLw3QLpnvMM5C67KY9vvuOWA2fN+n8BTOaPPa3B2AYaJxbNFxQUFCbtp8pUabazeeUUR
SmdguIVt1hA/XS29UADi2ehl0RGXzrlHKOywlDIsjvB8eiRNf25FOfVC/TeR8yD0LRxbGFHJWO/L
bzc6exopCPMcQLaUunQ/auA65UL9F7tjoGGpy3XhXR2PfS++g+rywiFTQT26R2AnzLyvBU5wlnNN
bhSnOPDU8YRYmSHcnebFwByoCQg+K958G84L6jNGdNn4jkyXJBpyYTYLAphudh0AhkYmdhfo8v6f
Vugw5k7MxGdXsdxSzXTUv/fYCVLgphzIkOLv1VqnbN8RfpIYV4leGeZ+3reOCrAyVbxVWBxAbd8n
JvhSrkIL3eUp8cvtQSyHTORs/7OBXjzIhDciZNnjNBsBgEjR1m7NMLcl73Q3cX1R4Fq0f48n2/6g
uOsop9A27Y/4szqr2SxMj7OPDwVtsW6piXTAcC/+FIGuGAk/6kMX9KKtMHSprgptPAGQrHt9lW0w
m5Ju43lSK2MXnn5sXErui630eAkr9FXje1yCs9bh/E9Z6ukha+KDkq48OMkQibOLQPOH6JU65T5A
biLpofpOKm4xPINYhWJ6MysOUVxUxsQEKRPPlJ2LIh1QAqtAPMYAJP43ilujKG+W/T0ftcLmEUSW
f80QUruAiB/JrFGlr2Wt5U+ChTSNf4cqyQ0APyCw8CpiM8megQhXJXr4Ch5II+DZj9tQYB314DA8
UPAIU+EV7RjHu42Km2W7kAr1kq0w5L6d5aviKafyfLR6JMzfkHPL7LHiZ3JODiiYMsWEkJVbbfX1
LY+pxwxnQNQr2bNt90AzoP/oNUCaywhKyYlUfGLKYHXmOermYH7Z5bCWAkNT/eTG2rUI7ad/LXH+
p77yGp8s5bAMfs/ZhP+aSOogXsZAr4pXETkTB6vnqLHEOj5gCxFCY+kd/J/5cRlUnnNIeAcc7OXJ
gSxj4y3+zkhcLTJj/SC81qsKUiawenDSYdV5dGKzc0YIMDtgIeNJNOnqEZs7OJvOXbbYKE+VjbmI
sxaHYkO7cHCfCcP4h3p9Q19RbLfqQiX4x+oipDf0Xq+MV896I01qCQAbUc2N4fYnS9lTlYk07foU
x3XGYEIv/n92461R4Jkehqb01Ahut/Tz2GTyYWVLXByAOdP8aa/faTUzRhqSt5/71PtI1us0RX7F
obJsHz2EUKPjkAK3Rrp1SkSmtDa5SqXo4BezvWHED0wm+SxiU8wHvvOSgVsO+My5T/6UF+Oi8Pj7
diq6odgUsfqgzAuDE7clUynCxB0bzYj32vl5M+vwU+AmoYLryFX3u8LJENxq7zH6Wn0FEalqtQc2
i3d8wXCCwfXZkDoXArGYciZMCmd7nbPc5IK9LjiL2Fp5LvgPPbTpTIR+C287IzhWOIEcnSjZwSaq
ka2eKri/a9iLd7PMVw0YD4buxbrkOr3+NRkEkk8t2JINSUppLZabssyODJ4OU0Cho3higqWzQdBK
lPEo1QEuyNmZ50jM9z1fbldI1C9ffjzYkosta59S+8TsIzqmK6pA1A/PqKlH9xiUXVb9hU5j0EqC
iGKm9MzKrSQiG9J44ld3QCUkTQfdzSKzPCf3lue6x+952qezPiKYgp9xdMApl/mMUsMakJlBw3eZ
lwmr5MeLNQ0fGak/XYAkBiJy8hz5hq+s8dRrc/18nKwIkmkjH1KFsN1wvntHd0ExbmlpsYYSjb2v
XHrDsJeFq6yoxBomPi7GM8NY+UDIzWjCV5oVrPUl7Wfe84dEuCoCwgDAyAO5syhW5IERwwh9LFaP
RoG4B+bCYlgk7iN1OluVWehB5wisWJuUnnCfg4ZUYJ/5k56VHaSM37y+zlauYWyjjq1tC44AFCLf
3/81QwoiTmwHcVFoU6cYFVpNcBTBcIpFAvUiwPxe2d4Vc297qJ3C8k5sMLVkdIVDuJfKtZ1L5mGv
CWtqEYDIOLXPlEnsIp3pjYJ28A+tzuU1WY+mRw47IWmUTfSCYJuvLiqZazkF4mwubE6Dx646pYx+
UE1SjvRmp/jX4453PjafGfb0g4nuhWfnwb1xfiY1bXsCtRzPD7jrFPttNOuZohexvvhOO2zN6roF
i7pFrb3gTaVM9/2Sc3HKtjl1ZkqjDWmgtHAE0K8fONetl0yd3QOZOQOCtUJ/WRgp5rFFsudkJeLh
SsFta6ft+Z73olOFXR5c/lPZqF+di2JXGXf/+0Uyekjnx5Z05EE3Civ6Sq52Nv3ZqLt0Yu1Y9l3P
0MltBlIA8kp/UwDDp+IjetS+bt+zkUwiuAAx0f44z9yyV7Zjz8HbIbLE/1D9MGzz8nUiyMHBokYo
bI6Ww53YUYdoQjT6xA1iwHtz0ukhYSoR1XvnAcxEXXI+WEXvc/OxcE2WPPjcaCeoDsV7HR24JwoU
BzPeLsz6ybeQQ5L6ewxK6TEhusvCp0Jvnia3cQVrMdv1sFIglXb32x/Ttk4zYpdJw8GRqWxoHsuc
IH4F4uHdCuAcESuQcIJJ9I+6toS6ROM2XVQddgkH6D7mTUPdhbnHyNP5R7T8mU8OZMzg+3avsr9Z
XURHvfgrgwNS8ihRa6TEGX0VCpYXmgCpD52uLSXrbdbppfz+9wOvZV502pHyAJhuhnqelYKVZ3mX
elvfp6Kb9tDQouRFrNilBX4HLLfZbrRSdjrv2Ekb7QAulvRQfGWYMDszeopr2FPgkbTYiiCM0GjD
piHWW+/+NDNnoiv7K2DZZRc3EXIZmK5Ptray8ZKV8aoU2fmbqQ9Lp+xkUJlITY613uNlSUI50n9Q
H0wsGjWdDPxLV3XklEdiALCDdNY+5CZuOyMU2SD7MYpy+PBri0CIYUgGyt5cXMmv38bM1+5CQTDn
i2RoLhOakchG+Tb39VhWGPsKyh5CQtwbRCo8StZzgYe9owcnZOa3gpGIgokwdlSujk5fg7YbAduM
exA4zSVDLHG5Yeg0bHzuGzOulpZYmwRcqQbktVf/YmQjouQANHcV0VchIvLnRIQlRdbwWLh+e9m2
m9+gbMm6njYZf9fK362XDQsFi+AyzqWz2cVy3hfe1OmJXcsQJQMYs9a2rwPpD04my0lfq58CPI45
AOXnBWCwLc1V3cJGPSOps+iHAqYatSGUu9/gPJZ1AinuR9c0lY+J0zT2Ws/P/5n3IOiWTCS1PbON
sxER0Y5JMIUjAUoq99/WYQjZDOLmpZsWgU6NYZwpb4tVQjU1XS2sGhhop4lxL57pSbS9pHH1j13G
1ucu3a/bZLO0Sr8xSRHqBZ3dRNsfw/FGQ3YlDm8ppBq2EFyYoTAbh/FR79BJKA+hEVAQLbwRm62B
2qHeTAKDkwD70otJ7jtC2zl0cQvf1WLMhCp75toYG47Tu++cF9Cgb4Zrp5Qca7jvvqCGH0Aw+s7n
EFzr8tQ9gzQc4FJabU83vPW28YWSImdSMio1GX0rHsBcLjX2oVLzOoXgyAC9hvWKimmG36bJ+lVf
UEuL39XPGNfBtk8LMzp4+ajkZNt+vu0Th6ZvdASUgmqJ2cayckAM9tBg2u7+2QhR8T/z6SyMKxSY
bzmrSieX26AYGhX95DgYyZhhFYokRPBefBYx9amt7j54pnVaXVBsU/lkkMm9CSDeK9ik+YvRScLN
OqAJsolbwdW0NiBldQZn9q1kvVQ5Dmv3l5uI65DpYDf3djfe9ffOmyBWp6ZR3SymuJdnhaVMZbf2
ObW9ZeboSJjk/BLnp3fwZH0NmsLf7aPtgz+9z2p8zj88WScT+NVtb1x6GDdV8DMbanLB1E6MjQjq
RHf5OT0NM553uwD2uR6qJLzA8L02F0GkuzcYwD0qQ7hys9pLw74LBOrVNRpB8bwiELlCvGp1nUWx
38EJFbASbC692804egKgnMBJoSNOEIKU9R0z5Ms8cBo1NpahjEanFgnMZyLP2oqJjTEORkK5Jkhq
i0nadMEWIUDVB7rnbnHhpDbCorv59IP9iKQNoDukGaWYaKw+LYN4OConE7Ql8t8ybXXShdYJAZxV
puFx0BJ0Z1878QMCCKOtSHRqv1OUmFDGc9ryO5LuJuaYBsF+ZPXWVa0AOH5X5js8WwIBsBkOBRkO
Qw3R4qjZdpkKVXTy8DDjnWh5UvNMuMB7HkehdXcoWCTFlCRdwuluQDL4xga3XNYITFlLPWxVa8Zd
DcxtcXOKc2MjzUBE3250Z/A5dO4VjLsztJp3YGv1DZf5h8bqxqs6Zec4FHg/1YIo3jcc80IJ5LQW
V3tuM6b9CtLgziLS3FCHPvf1ppFN9Px3wMJLcnDGofx0CVXfd9Q9+sjRP3i9D5jOzIBdK3qbMgHn
gzud+JzzypbEJTSpIAZVDrmJgbiyYPeccDf2iWOwrx5GDYA1w0NhVUoOe6emPGBr9D90LA4xXJQ2
FNYyofaQlqzewMv48D57QjppQNjGrz3TijkC8DAmKdZxdFEvst5cvjEeF0RYT5idOD5nVmMKN1HH
bBRsBfjqmWM/HrAwh5NfzHGTQGFxg2E1izxQtFk/rNQ77mJporNSAU4S/31ipZyTSYy6ltgdXNTr
24yj80K0TKoMN51AaFuOFmqrHGxkZL82e8QO0Xwk6YkGDrEY12K4DtZxskd3ZkcIuM15bYdK4aqF
jtSztN/c8BoqU2y5ynA67vXvNWAOyUwaLp30JBPLr+u0ekL00WaYnQuQ2phS0RvesyXRpQQdgQtf
jHCSIh0zIoHytLHyvYCq0BwaTI1a2avPTr6bpAkTF9fZr5+mfXJzMgwdexV+iBx9YaKXh3LYr8Ts
v+MtnQgev4m2lidrYLqhgBx+pPoMBSGA1qUGaxSWiMzfIU9T0oFUYSuENi1se3dkpFBFz75ILZDG
jsah5WaOjv9sfHFILovf20TaMPuoh3srYKwg6AtAXnJ+HFsgjlMdC/CukRdkj+sMOTZiFgk1O7kA
9QRmTSOeVTSnBDW7CYi/eUVbE7OpyJVc11uoPd4t5LjtTGRNIAUvbYSqy1XPAUAYGsCmviwrdY5+
tLbKjKMmH15UcRThkXBZZP97akT1ovZpLYXSr7BO1ptRPNmWTcFR2rYzEyj26j7/uwD3SJ5vfKBa
1j5wf6wVDpBRlZrTz6P2zemYl7uuDhF+OoImYONy/e8ZIVw0oC7wRpKCbitm6fODZO7NIsul9Bsa
OCyjiwzgIkJWyFkraYPZ6LyH6IMVx8PKD64EfL701Ca7atIKGcRlUfZpwDVtO6QI1A8YplNk8lLc
H2titQBbVVJjFlweyv70eVuZLZr4LIcWrWLiPHrEVu79GNJJv4RC5QGNMQ8zq0C5SBA8S5oHSvkv
vBp8t7JYvRKXwI07UOV+Uul1GtpqvC0q8D7vqPOXAIZhdE9TAM3KMEm6T5Dt0vgrYuWVFfS3Zzwg
jR3eq7Knna4IB1cjlUkjY6Mlsc94J32zEI0DfGJFyNImQ2UFZ5TZWXrpRVhr0yOk/G2tQue1pvoA
ALOjRXDawBoiuOc6wgUQVwszN6KNHXA3qDLrV6xuS7f0/ncf2/M9mPhZH/2dVjP4NCFU0f5len86
tzBhL8rXxQ+QWJJTeYY+8K/zgO1j+O1A2kSACyz/Nxy1gy8X7lyUqzC8nBD6uzx2qqnLhv2hx0TI
a9Lr324/b0DeS/YcoaZcFda5SEDrNHzJxfYzmDKYCSqSD8BazkwX8L4j8bIgVxxaOrxYV8PvYn/V
ggGtGhSGiHK4Mm/5ALZA7JOi2LiCMQuBfH9rIR0skJXJ2vt98Rk0LM80JxZZo0yGlLbOx1S54AqQ
sRmVhGoF5zhKSo16LTYLeWmZKL5ItFrmdHyxmim94H0lFV7BZanenfe1/F9LFsoIqn7XOvwaUje2
B7i+l5jo06rN2IYQLDs3AhINpP/77OcLtmfx06WfST2MN+HztgQIZQcEAWw7krGKTP7v7gQr8adF
V7wKn9aN4wPxa6Ac+Nh6OjlAE2qXLRuA68JcWBdXJ3vQJqV3H/0gFpHq1zcfLsq+8AujkAH82wxH
F+E5/veAJTKNehk6V1Zi5R6KJgg6VaYwx8WIbJ5xxdul25r0MGYxy3kFKnD4QbUQtdXC6vwcWPOF
JrUph0ID4CU6yzhbhBoj+XgV7mJsRgY6NfbeNvFCGlePVgz2GzKDr+rVoyeIW8/+F84sTCW6juzC
BMcaGMCiUDQ6EkSDqiOX5MSg2H7gwCnu2wLLl5ajIJHpilM3fyflSMYHqeo2EJbQFV0Pvk8HaU/p
TPhgiEdbdrnru/D2ELo/oHbXL+O5yz4nx2evYfESjMXDK+YfuwNs9F+BNffJFiTsKMUR7+HAo9yA
bzNM2fEB5MXAdJkbxctO4Ed+7L88D3btl85gG62HKfq9WMxlf7yqtOpR6DQqvyoDqBydin7L4V4d
chCnc3b/WxYEInKkY+dRT9+4fZ3AQwU5A6C1orT2DIyOblFPa8NiMC9qSygex2EonBELRpdyCwel
O97QP3U0btxKquOpnrzqEf+hF1Aa7cwHzmEOG2anUEfPlQgbXoVpUkgLQHUwrGj6V6VVWtduyHGv
KLXvKm+Qa5VcJhuvtZ+KRbgxLXsVxv6H3bpzNvj/vS+4Q2rkzDcEDGc3DilYbxIRsWa+ABD5NCCd
3JJQENNkBemFDymYsLhVRoaOKn0m1PLd85TDzgM25B//OkodsbrpV5Y9UqyHxQ0R6EBI1x4CVQjT
C0HtxP7004OHGanjJD97BtW1Mt+sIDV+EusOok1MriXVBv7GAhTHP3BlIXLKeXsD/8Vupqr0ySTY
4UGV5Eo9/L05rlj1pCbIh2EhiohxZ8aQAca2hPneBSz/MsKy547k+ItvyXrJw4XnakL1qce3yman
53J7zJWzmFiMY43N9cUjKXLgMclwmHcIYOIA1Vxr8rPT+xsrUGs15A8w24Bq6Vdi+VPPibbcpYCj
pYrgPrv8r/jMwnMC1d1L0WSXeoc7PpsLmWJFh3/zb0SnGnI+fZOqe5LEyc3ZM0UZ9ZLbwPDlYEs4
m0TPNeC26chz+Icf/bwqWl8FbR8MgEpnNBughyr2ToEvhaUYmq+kAnqrtC8J2tEtnTNU5YW3nses
knnnfAYhBfy1RSNJ9pX3Rp1YJQyH2H2g7NrHdXBkZB2wJGsqR0ptUEbdabb4hfWqDJRS+CoBBtDC
+S2ruCXdYulOku5MLJyh8BTE4dmud3JeHoC0d58KEE7ff9dLcJ1OrcfIYDCJDpi6Tff6Is12OIJw
8fMriO6YKEYbrYHx4i4fYV3o9t+F40FpGbJAc465TmzgygP87Z78p4uIIQUb/PC2De40v+kXqHg/
Hy1TosN2i/u3d+CPn3I+snAGoa2IsDO6WBk80aHI1HCO0A6eOYhwz6QzylrsY5Bzf126QkT03xN3
lvWv2VJlFo55rc+6L6RgmbvBhiUQpPhqHhtkJb5NA1t97zPJFrmdGqoe8kAaw1B2jVRw81qDcQ4G
v/jPJsM0SquWqaUuPxHx3CbDCZOsXkUJs64YnmOEQLmxziq1B+da2aDixXDWizSNGTRKdJtPaeqN
WDCvfZzswbslOrgQIA+OJsrwrfJ+afPI2uFapRI1FNvMIaxDLrO0CvfCLwQWS8RSiZBk+5VSwPvy
OIdomGBsFQB/HhHJgZlcSxRsXoJt8CJ6Vlrww4pMHGo9DHTlOycrbC6TMYDcRiUeHkn5ioWWIlVV
7TT833YS40FW2vAVT4obMYHbAPgIT30QoXk8V9C579CbJEC9+oxGjXxkBly1aGBkZpPVGN6dSbgn
Ao2ifxM2G26pz+ny9EY7gKb+hLAeDfIriq6TStfRrXHUqQQarU/bzD3e4aB2HMY+1K3esum8h5Nt
+OyvmaAbGD8bXgOLtsO0xm3X5eJrBiUgBArcdrPESnnSrTwePZrjeNbuYcYU00w3oryB4iQY5d17
jyehyWIn+sk+kAjpGYMwskJn8fnmL2VwzB/d/XXPFDvigWXdT1EC/uIOa29rxE4ntNM5SP4/tmoj
SwL3zoLpa6ZDhZXbWVCbZ/X1KoSanwA5vtEZpj7ly8S3qOXkT80cjNgy6TaRUgzCbviG1s7ot0+Y
sbn8jsQzCToYMR4G1+oZuv62psGacPx+jNur0oo/vVLFi8cqQf/vuXUgTwxYQQRCO2VHvQt06un9
bpg5P5e6KlHVEKn87j70rIQFXxBecd2jug5k1ClxgvtmYZ/32A+5MQ8AsHCr/yy5JJQTXtFq4lC3
iG0RYIC5IwxVyy6ZtBSSUi8ivTb20wr2VKzHV75rfdxfcdI6IuZEMSTAulaZSQz/0OV1eCf9fho/
XBUz9APByspPCpnLa1NZhE2hr9ABdr3IGinVWQ3A4H9fGGgCT4pWeIwNg2VvL7cUc4XxHKwTM9ov
NieFBUiWeWfZuMojOSGVOXPp/bzW1p9AfyiriKB+6XnzDca0F5Eqbsq/nNkyEFT1LWsyfejr6aKy
Lx75seg2F0fg9A/kQpXhfoCrKFg7Qy+/fZ+HwhpGPPvC2S405Cqa1Zjsp/nw33/u1BfAJbcJuTUP
lJnR3jG8WrxPUp4Wp0jRfpXgXU+OslwsYsmFW/jv9kio1ZHMQ2VCuATJAgUtk88M4nU1ftsKhpOW
zNQIoyIwyK6nkv6iRljO6mUG+TGrPteDnkQHMEhjnPgeIQupoCeHe8vCuq65p5mIpVduI99yJcIU
iwp9yx9aAKX5yl+sObGFLzK1awfrNypDS6uEcZEuWSU22Rnydg5X2M5FCCOY6mT+42mBQ//roEIt
XOseByvYwAi62ah5sxz5mc1vw924/H0yx+vxFdJ5r329V+pXS/2Gu39s5YPeiQ8Cnu8yEJp6zTDV
WzQ5YSkTELIr8XkFquEI/NsQLxR+cFaNjl7HrTbk49/z1YDz1Hvj3M3EHQMLT+sfLPilB3U0bXp3
zh5PXp6u2vgdmZN/BsdEsK46bVTsqJmNfx5RsClDqWq2RI9o8Jrg6RHvQYUdtqa5EihGojquwEh+
hqTeXbOvn8gbq44Ko066tpCSpEHbirqfplXQwy0OCFKfYCT4KJwJ2fLLzQXLRAIKb+OTzzPVxtUa
pgHQJRez1q7UEkk0D4lYwUxvjpWEDZvxe0kd2U25w83LzB9xOgvCWCzfw5OuJvs8ITSHo1/Mnk0K
QgLXaotle/s6ZJmcd6cY9GNg/XYMLHAfVZm0y1ZM5kgcBZYXdxp99C6yWfchCO/3lfzSbEmALqry
tt7OlQvIX2bfnMDhI6xz7aGSbWQG+Q3u+Ok0O+BXyIkpeT105w2/hCqjrHaDytzneUm/x8mSgQbU
LCDXNLMNd36XUUKluhwS6Ml7UwxvuLYSm7C9SbCLFR29dVUM93V4e3xmIfA9kH1fvZNc1f4zPhlT
Tap70IL/NgHyKheMcPvUvIVQ7ttzfOk+931fesZMV4eBquCVsOFbv5WQIA4jRJrY4ZzJeuClpKnF
/h0zZVW+foeg0cB6HWrNM2ZSwmFLpN8yuZ/Kba3NyPGVJmz/angxocijgGlOqCR3RVtFh97Jt6NR
XfrwfJDfwtiAUxaYFwGZ4kW2oCOGv+fS1P8J6trLiZlzVpTNoUX6yXs7pssUKzLCLOypSaf09rl5
Oeyht8gkkRZE4RMtliBZ+CjYdphT0EobBcqg6F66X0wChpaMjfWTPTUZ6N6y/bVZAov0obgrbnyK
5pIkAP242b7oY7EfIbtdEMlMqZz+JkjBDoW6WJtGUmLSyJ9ob2C/VRX8/rN9M5cD7g+SSG64VxOC
bcl8akRBf0PiqA3unp9uZZwR2qB3uu+tA+MtDqWMIeED6pwsAizg/tpglw34rS2hAfUEBxIJKsKc
pboloGgqUhCEm7FA0NQALhG+d3TvqhYj5GTqXCYWeePBI5jEMExpih9JoOvEXIKMpGne19ynY31t
x6hJCIO3LDcIN0tdgLWyTrTtgo6GrnTTyRA/0ZyuqfHOAACoUAqeVmTOzQ1V+GAgY9tRPv9qC18m
C6XvdD1yV/YQmJqyz10+9U2eTXFt7mab5hIB9BMHdyRlq+G3Y6HDK3L+rJ3nVY2St0s4sbSfNKqB
CyPC+l1lAwC2kOzL0AgGAWMkHv+az4Yr70yOwJ5LzHNVEsG85Zjl7t1zJf7vhJ36WPUrpklDPM7D
sUJZb62+NpBbSEJJZSrMulsWjhl0I+gDSvRMmSvMp0bxRjCFYuWYxUgRAakayfiw2akNpJlHKwTk
zsbuWePgPiHX4W3brbJs6w875OT9VGjhcwg/nhNWBQ4dPkXvstg4SZncdI7pMWEMAbZjmLptHQvM
JfQ6NtZwPwah/oyxzWj7CH4r/Ii2UwljrG5/09t7kTBxIwRnxCXyGEcdd8NKMZ5chtwI4R3XshL6
tEU1jcNMI/gaR5cNp/DYJt+s7BJfhxBI4/M2Qq87AMYM07j0bj4GxJbybUE4nBo1o9rW/ZeBRpav
3NpSQhekwO40UTANETsPTV+huigltFWWbuzkVKqSjVgNx0alo+JQSmCMUqSmvzdQBFU5GzwHaTlT
aRfc9qE+QjJwdy3Ft2U5G3bKHCH+P4m1Cc9q3qtyoLHAyk+cjEnjGR56nwoC1MJ2BiyJJNPx/jab
z4JCbKNMDgHPOSub1DppIkq3Xw/I2Z1NFoodlGeJTFd4TQKuqlCYJ23AoOTJKEitotfKQt+C4wMu
ewFBcA16+KdDlD0xAKyuqd3bmo6r/Fjr90PwhS0Us0whulbjdqenCzaWXtyZ3dJYaWMtq2yz5yYV
s/wk4fbXNSZCZbJ6R/v17rAbsbDJa0DVR8o6k2c5vp97Kbxi9DlrwHLGhyBBBX3dxqmfXIklw7Hf
/QJRV+mtZa8SC4Dnid/FKXJvwzNx1HNME6wOkB/x7WoSWIqs3b4yzP3V/b50Y1xjA1MMp3kv5fPC
RE01H9p3v0BoMgkX4C3JylhJmFzj+rybaUiHW2kKRE3EL5r04kEvvfSL0a3oAh7r4tVD/wy2RX+S
oZ2DjWeXtG5sb6qaOZmBZuwd24NDcC7StR5kAl1ZzXGMO1feYMD4RkB9h8g7wZyicEaTUmjVGC0e
gFXm+3YziuZoxvqqPkcYXPeIMGu+BCITtKHwzDTu4eD4Tu2Kyx/+b++oeblZ2d7CDFx+z9E9cMlw
wFLxRnXzAVnA3c8Rc3ld9tf45bdC5lqYpH1zRJFvvCLtZqKv/ITwFc86wfYS2BhEIPkiM4xhNhRd
VuBTA1PMr3JW9u2vwlm8xlKM+sI+EXJu0M4kNfEcPs7V/TGJXIe71t7pvj37RQMMU8BrKZ86wLUV
bg6TWXFADXxYT7lIQmK7vGtZHQZa7r7ap1an4nQqGY449y04xE9sp5636hVTmuX+/HpSV6cSECSP
Yt4VV9/yuhQUS/Y7U28FGMfTpDTv2OZFZfJkG34YsU100nGwuDhrParUvJEyV6db7aIbcB6XmX/u
WxclbQmTDefqu5dgZcVkYOGaz2Zi2Gyi3fb4FCdsb4liwnAjkAq8NxtM9fFefeTNNvKKGKBpAjZ8
Kb23rNsiiXmvC5BaYu/rhWE7YzavcrpnjfSdpHGxa0nElpHxihNPR5EECJ5IIGMxKNtj5ibWoW7G
YRdxpsxvPbHO/Zf+T+WvDE5FICjjETM44WR9/gyTbvigIlH1rr5h7RBFjZ//PwvP/o6npxnP+Y0L
XQudbX/KzWYvL+cOuiNVSy3661Ntr9kyfdbHDH1bVzCulwQKLC7vzq51IgV+gOhs649+PjBlnb/s
V/qkpUKJOVJxwj+KaYmGuuaq48WDxHW4Tr+43QUjQATd6h+hH4DhptFHF5+rq60yZ5l0LsqwTy1H
vCuLldrvzsbIn75zw5c3tO7CsGnXFz5TGyj8aDyVZ2pbo2PN4l1ML9oURvCCWFyqcoWqN1dtvTcj
7GiTKDjXoy/pjmGkF82PMuU3Jo1SmHgZAQotnONtXJ7AB65A9JeXYSKTDI6ag/40IgaOkx0VEV5Z
ztLkqn65/5nxqWsWm6nSLi0CcmfUrUCUFQXTC5iYL/MWrstlx/YGnQKtPoMg6NBcM38FrANmXssC
w1pZXp91GW7NCjB0YH8MAsWoPWEoFIWJMfMyeJOl4nXztlOCog6oe1MhWte2uJrph1TUIf2NRFOb
9hDMuZEBWH5X/603w7ezgqldWcn7uJwTMPuo6fbu4FgdoZuvnpmNwzN3WZVgVIdWZ0ttjFg2hCGH
wjxWvqAvYsHPemZXQRs0XJEyWoV5BTEq/PenM+LrCCekfgMenfaCSLylR7xMIXlmRK8/BRZMZJfe
VjxcWP725qElLiHyo0RmUFzvArUzzdaqT+SezHSETJ0wP6Pjc7DkNKaDgEGvnXX2RlK5o4CKlRtH
PoxgQnQySonyyS0y8eI8sMKhmlW5/gvQJzlM3bZ9UcG6NWcJnT9UzVf1zbXHXTIbQpBBvT2Ho+iS
kdBS4kg1+6CWRCS2Ivuc9l0p+eXsxhZ/EPlIeM47h4pulaorH4uBO2i9B3y+IvT5IkMVWR5f3a9R
42nWbPbuIe8IrK3z+fIkHMsaUYD/98iyJOQtpldfCQBR129r+FnkjuSuHMmqGsKNsrneMGsHCDtk
vfHIqFtiOlAVqB4QYeKmZeK/rvbTE2/EHApMv29iXQk9GSstqaTxn9upG9cct3njgdu9u5q1byJZ
x+HTwP1JcNQzqCFetoZEQLlo8D83H0YtHGURZ+JwxhvrR1xd0h7pfG6YfXfAkn1zV4IL7iEJviZF
sQDAaWgGQ6URzdyNXAPHLGkfucowsq+g5UIw4e+yQcYIaPJJSpSwj1tLyuqf6C5Ybz8b4t+nsZR5
MgHsl2WaXMxTwvjKBX9TAz2GuGHmoGP1URs/5QII0TImvCO6zlKgiOfqXe0bM6///pFr70mgVEyJ
twUrtjGMebN+2AnEt5ubD1JCpnCNr4n5Inogh/pJxQZ8WfpG8PMw3EUvnAorrEfSJ91stucRSeEY
rw+R6tcO/GPVEMcDcP3F7EVh1bbqi15Col2BRFAqyjfJDJTLCF+Vb/73wBnNq6lUx+zFlSOvxqdb
W9YUAdO1LRKBQsfSWT0K5jCrqbPOM5Kv9WCpolS7gpZXnDoOH8Yo+tvq2U+3Tdq3ARnt6XAel9/4
YAx3+S2fl2CiSE7wj7docHKYfjn7kKS4kAjXBuxmzrUfZcsJIy1AK95mBoWs4YVjp6COfHPwL6KY
DpaZBosImkiXnXuLb1UpLjpMhtySR68rgFjsk7oQI8N/5z99LkAgn9MzWeHi77DyPbsUcOPcquPz
jbNI3UPpXzv/ZyrxkxNqFj+69ozvgCYKDDhOhV7MTSh+R/yndmys37D9zcGa7Z4kRR/LIjEPoacJ
jBc1INIiUoYL6xg808/s7IHd7ftrRoo/19Cg9qUiEuTXkTq8YVBg8u9NNmwh8g9bMVz1NNVcx0v6
hekOzxyYLb8/TBdg+PMhEEEIvIDK0FoWPMVveG6e4e8RG+bGCaAo3y7xsGRUyr7Bnloe1mtJdE1n
zrwihLIEQiuZkEGaKFrQlqzoMpziapF0vMKppyLHTRKkQdZaiOEPyds5plJXeuDBudIWdMt/AXeQ
B3pbrzDFt0NfpJAMTh2zGwRT6U7EpcsBTI+V+R8jWmJ/uiS4SU4lJhMEQo6UyXdKyZtYQgWyiGAw
mnfq0E8E0eeHunk1x4BmWZ/h8tAkPbFJRnCydA/5vu+PBgitDWMnSHbLaNUCu7RilXkiBZ3hmAbT
S6nxQj7hcsYgVcOCMTJRF3yA4S7OgosiPrU/70F4LD9BIoXnC1bT2cYl1hIswAsW+gzvNtsbjNPt
f0Ru9gAGsq+5ib3j9DTNrSZZWzgyRLbo0AcUZOJMmmB9xd0K46/uJbIig+IMvZtuDHqEeBEZE/r8
KUeHvdaIrcGi/6FEypTIK76ssWJS3/vbJnl+crY0w1jz9HSR53s6A1E+lsl1iYvHwMOO699kbB0h
4O1tpSSfQ8OHrqjInrjKgk8x2cr0Vgq/9JeUz+rdWqROpZ6UwYKBb5KCreKjgn51BXeHef2nq4AW
/DD7v1BCAoTDIvSFf6iiwHcvTlzOSIrWndFIozktGQLq8Ymb8f8kWbWTpUo6oxa6mQlO5HTGzooN
w3WiTby6JQKoJ4febt2BVFyAEjIKWjB5/l7v88thofyyGqngYbX9vO9ic1ZU61gcNwjG3Ml/pAgG
K7+Pz1hppmIsMizzDl3w3FOhK3fqhMUrvWg4puRAF9OeoSnWIBf4v5VSf50eYmvztHSp+wxLc0Xa
DanPDjmMl1r5Cljf3SyYPN0WxXBzRt1gTT88d2in21gTL4bDJhWqtTgtTqcHlxAzK/ELw0pnW36Y
OVUHaDT9PTT/SRNQjsknA+NBDDEiWguuLKztcixlWH/0RYxapCsH7WaHYSRCq0bfyirVjMXpKVwL
SglMFphm/zeDOfv2y3N6rF4HOfXLPB6wZ0SRRs0sTDb1q9ofOtJmX83Y+WfcAJkBHwHb68kyUNdH
q2Jxiq7nS67Px/2jtKPq3lB3mtJNf2ODuI3Zjyz/iDbqrJCsjo8zhH6XzGbfnlSxpd6uRAF+aaep
4U3CEG5HA5eCRPtlfEfO6pBftBKpfY0vLJ3ZgpF8K09kPQTxpYxvLKKrQZtZQaZt7JuuRJcidd1+
ZcPNYgwqM/v+/KY8P0dOIcKxraFKd20MiXnrph7TokboIg6o3DTo+a7zaKnpjremIBW/HsA5JyhF
9wPeBvD2UNqdj74O6KsW+Uib00OM5fjkAWZMLNOfU8m8jcvAN+bdsV8oaCx6Wi939Q9MNBc+dOts
vNMVETFvBH1cemzmOKVQPbjfiGtG45OGJ0B2KRjfK5fQfMdnIfxCcJ9bekr/LMWq/RD8qleA97um
ImiowsUVbwF3gS93PyRl3xg8220hIGKl3F1AqQkAsCdqfEAlVNcVUSzq0Qcd9qdVAT2IP/x786DF
2vy8W/bbrOnniUS3WhLFbo8+XIVZpnpFXh3Mz5RUDL0EpJGuBcUUpvoC/SaixWrm3k6Iq1V/yK9q
pvhN3z2BKi5y8eNlNabnIAUFGkWqYXzSJ7gcaI2GkMTk7LrY4D/Q6lC5cAg+bw9o+eu+sOa6PP/y
Zf6vX3t7GNHh4JWuj/Alt5h90+8dH86iMdEOf8z97wLnfI5QVOsIhvJUZuPNHurVs+fKCVeWzaO6
6Z0NoGBFh+kGrpAtAzELVEEge8/4rVGNbkVwWKSviHDBufltUB7tndp+82c882yOpaLzNvwothKP
8qfUEs3Dj5fRKu2j3aMioZlQHd4DVWuuaZAMO7sDOsgfngd7lexLXSHAWJzvnAfgWqhfwfF17QNu
w2FYHT22USitNcU11oiupmHnnLWUzFDSX5FTHkCqDjVmI0pHUk5tNG9vdmnCvsouGGjsMH64Ujov
E7XxAs9UtMmDWrhJYwtO1BFEOICnzIwdRizonYX4PTjXRavoxW6FUruAPSM0IouO1LYIzZ94NtN2
gMFNBX8bF+L57vusl8sR0jluR4+AW1/JZ7C8tGbR08xhmw6p0kjMBP/aEawGAYldk4CU2WhcbxHD
uk2yAwanqObCpnw5AWimnkgAmYyyDw2tUe0hZx7VgUdwyL70ppJt5TxCiQB7eRI1HYuRrY2Jc6XR
DdrprXIqY/n1WXwBaEZFAaPuMRSvTPZz0ewHL/lgpI3BeEDtJ9ksR/ct0SBcevIfUu34tZhjAPwD
xoktDYKpJrgIx98nbdHJIuqEyaHTRBqDmV3Sa/95nNgh8S4xM2uqv1CRgQyR5TKK31Vrf53AjyCz
nwCfQMsV8+Wy0yeHeAq55QJFFJ8QU/YbyKhFaYVzV7Z75E8Ayb4sdJ0es4uTzRrt6uk9xIdGfMtS
YdmWgnyN5TI1DmVdfZ+DeV9o7XpG+jFaygqNKvN18fafXf44LfaHMCtH54hWDSkUkTCNmyYHaHyw
NToAzjB8ylmDj5Bj3LcJ3NhqjWGizFsAcPKa/Fm8X12AM68os8OD1n+TQwq0wYaIEx2G7XbNMfZt
HEEJG8fE4YeEctfVR9/VN+7Kjls2LjkHEHOviBOkV9TrIhfEguvCPNVBRFFIYCx2ffy5L9gpxipy
SK3qIHyUaLCLc7+IgJAqFeRJU8e/5kdcbGtreWTBi3PTVZGuT+xgKcyv1jffAmoaJUiv8HvAM5JY
aGpQ3qd9NRaYKd1lkHquMOss4JdD1G4zoL7KTImnBcm6vM1h/HCn6h2vM6676s3539NklQMHC+9L
Zu4FiWlaXSD9fhfhMFfs4Xr2qTyLv8Q0voMw4RN72ov/w+YuLrtZmUPeNJzeHI4qI6c8myZcleWZ
lRTF/4yj8x4I3vtLXxaYcXtkXhPhR8AgxY/yKYEi4m8V7xuZMPr11wYgkX28UECoX3MCnGMjipcJ
3oy41OQgE/MpKWlZb1fflGE0ittLOz8gvKrcUp/j6wsKsobwR0BKIx25ZqPcNbovQKlsnKed8X9L
x2/SWEPWCNevLs6HvbhFl3qCUCFnD+6uhMorHD1oEj10pE24TmNxsQYdOWhtCv465vzayGk7JbLP
fL0usyNNwjP2xuwKmHwcvcFKc0F1duloWmjqi1im0c1iAC7gxvSobLYvBvRXCqdqa0gYdXH3yXHK
rIMv+q5V4cAcBVuDTNzWWkiNKEw195bBL5+fkl/16AVFbb8KRk6kuIP1n26kHFT3NrX7IHdF4494
WJffhXDBcv2kZdyBlUjRvhpqKKGfBMJqQ6Ovd5/AR5/6Zmql64dPcO82A4Ya47ywQTkvE5n3NN0T
SxmqF0z5OHART8yHjuipj2yd8kKSay6V2s9utRKv37LShHvw9B1fIRvceOxPeFLh3nBFoiU5LD2i
+enBDrz57q19rWmcTXjVqVbQEGVvfQJjfBs79Zo46oKg3BoGNQh+0Dbhvgnc+BfM8VbOYvevizla
n26hYAEDp2NRb23JjSe2T6U8wOyvltyfDXBcGpRzUDrnSSxnMnWpuJaIccXrg58AxRClsm32Qq9M
+JrTZotSnjxjbEztL+XeC2KZlgMzMwFOFyuQcBd+JYgCgNySBgzt8lFLrRclNl8a4gw1wFXOpQo3
8EiihfYrU+mmJ1nbVUrcv1kWXrco6o0C6HgZPwI5MmShZPdbMxKBmwswqisWklylOu6IvFwuf5S+
YdvW2V/w0RKeHs4hFM9fmUf/MsU5cn7zuze+6b+9uzDwNdXQ7b365pFwLbMTt0Ub36QhKB1vRTsq
yexc3kfmJCTMhQOPRjUBFQyQyxpXQluKa3VTGrg4jA8hSCqOeudnr06FX/JMpCldL3DL8bvHBweU
KGgdkYmygGfuU0gDOMDAPTiqCUjtU23TTXAoky63ScjXTPAipJ2AeHT8sPA9IT7pe0/QZYvjSVTU
K4XGItrCNYMSxG5FMMl9RvMxOC88m8i2wIp1zNbh88fHhjO9N3CXk8rNQ4TJWbiTSubUtDpIG7jd
uu0Of3or1JS06JBEFOPviBf/HIHhbthNidrCprQiq18kJjw/oO21+Yt9+/+Yjae7Ry79L7+Ns6pZ
HDzau5Q6//NNkCRgKDTA9dp3HtXlEwq9f/4scgTPfnWUTWTcoM1nUz9h1mmq9cP3CPLP/J104Y8E
qxwSU9BtV2i/vpOQpK3G2OugI43JKFqb0o83hJRCVfw+HakgsyeLGOdgG7yBjZ2kypPy+X1o58FA
kydYZ44Vx+3RL1m+BauESEMDL8foYLQJR/jwFyDWOkUjAYLB97BqyiduKyqTp9mC9LELdXiB3MRw
n1deMB5Hp0DAxs7wa6tEAT0HmRulixOujS1lBKkKvRjAqcPd9SLBVwSwBKCGrOZA8w3uDvHhGoqv
Uie9WRmcdT3uc9oh86zop/EbP2Xpf0gLnc3gc3aKgg1vUA2dYp0vrRW5ogBUi0EG+P51/zqtwbNq
HduakH92cZpNTFalnvipqM5dxNM8spiGhXoy8dtNZcVJggDQhdYUqN0OyJnZd1V+TESejIDLnyGr
Mt0YPCnu1drvrEa/aqWIQQSGMQ0jkt+jGlwAo8JR6egwG3SE+zryJP7r7u/vjrzvF8JNXXudZq8Y
tAbzqO6KdgDsjFSFTtZRbpbLEqcw/dv3tMPsKlNLgp6X7M4rjrWq0s+54t9XfxYHqRkGIrVwoAHZ
EDmpYcOAr028fYIBTk/H1hM9zQzIHDx8OCHg5ifCIRYjGoIwmvoRnt+ckRE8D1vbQaEuUQvBSgXZ
8nTVGZUJx6tGZzxluM3/M1fsHIy3yvRwaP4BNdF2PRTlBxGZIUkqPU+5CaHXe6VwSc/KhRQ89ih2
LRRPrN9AyuWx5RCe2Qlspw03h0J8EALlZwII6e5JNpzq11CDxR/Se+HN6tk7NL3Fto6aw13jfS9d
OGK5FZNVnlAgNCgPErOfi2Gc8X50uzZ3YDx/wGg0YJQVw8XF2RRGCAzXoQoTzL6pJABP/o/0xJ+x
NSiNkQX6NbBRLYSB3NjQvp5pRu1nGGKmzciCZoxde30XKKum1GXSfOVuVAzrMW2QeZoKdgdPpUpK
VnMHq9KiW/K04zDZ2EUVjRsofwguTcbjSJc2BdjqSBrstUMyKdGicjhyurngNKtIi61yiBpIg7rZ
/f6Fx7fIXHKlF56x0SGrtnKs+bcgFpuMPiSX4G5cwfQ1G8WbWdyuaUVctAofT6tZEp9nYbDU265M
psnKrainnV5Nmv51zavKJ8Fyc/YEVuqEdpIzIH3Vy0n9+6vbz9kObI0bsOM++SDZPlnI0n2dE5kQ
YsDi94dDHK3eKzFgXmIvMYMVBPBlpWC0jga6TuAPeGMzQg+Axb/WQrIvSN9ltRCB85lPDgKr0ywZ
fLEYzGaU/pdK7KYGC7E0oq07h1KO8wB5FNjiDNEti2I27I0D8oEOINAvIXjFmqXXGltu8EJHfxKW
VAgYcoVeCg6NcFGS8bfmiJ/gkYWBh74i3zrwVj6bKw52hyXHzVhs2V5+v+AUqIPzVArVT3t3AcmA
2K5tT/qM8zUwXIasGWY1ZEQMpa+PvGrDOmiukI4mEHiEIAS5ZbdBO7uOolRmDjSZugI4mHrIeiVZ
4d4b288HWSfXvNH597OI/NeUJ5b/udFRIyCASsSNgzaVoaxsQmEhcj6eMbomJ2vmYGhwgAvI/ypl
/7x7+FOWJHG+tRIAGTJ/EGRvfoi+Lh7+95pkOkoGsfsTIwPfE5CxhbK8hk6QT+mbjfZ7E5Bs/WUV
K+aVPo6MCC7fXzhr43tQ8ok18c9FvJ1FF/NXYxGIYPnZ8LzzHCMS9kH5mxbHet5j/VP0K3SYRyaJ
rmPlbzRZtC+sKepcrHtJEgPRjJDJTOv9Lo62c4gGfjY6fGTRCHv8r5VPvegBKInhaPppMD/uET75
RWNClzowY273tMPWFnHd7sckKKShyB/msijyGM+lAPDGKJXYyY1XYSthaNxruUZggKWEIpAAhOnL
58ijn7WkJxs7mIJqNlaC3iNiKA+ujTIrV3WwlOgX+DFw1RUA57DZ3GpALIPs9HM+pJedzgxxldGk
ysLlJ1r8vigJ2IvMHyUPooipzhgcQPwdVMzuWwNExuTI+pciifT1negfn2kqXNp7amimD1mkKZaI
jiD3tk/+kny6k/ECHUJR8PMU3L4tFfK5IHeqiHaGkfrxEo/naWisdhGfj9hHITIU7ojpu63nOY+p
SaTaWo6z4gjZfQWZZNaPFnAemLlLh9/JKMQsCgFmzY4MJw/dN05HGohKjQGZchw2Ma7jYLLcJvzr
uW7MkCZeTfIhyzaa97ddcuRGLbbdc4Z3w0quIYw/4WHF3iw2NgLDu4ZigEfs5Mk9RWSKjxKrFTg3
SGdnr6sl4QcEuuCrX2o+88DjwFAdZ3qzhynyX+iaF8LlX03G6ZLz1xAAY9I44tGfr+XjLs901aW2
3XMmBeUNflQgbNTe8i4dy12JpYaXge2vspn2WgQtT+Kwx4VeexsmZLkZqb3YCWTxYfea0oLomNrb
6Biurwa1AN5dTiPRB0ddMVJDyVaoN9H5Xt7uj0CLQCi7oRWiVJPC9ZZaA9hQP7wMH4HFXiPFCkrV
xgqPwgU1NeTvwUlWzmrMIt3piN7fwAFNG/0Thksa1s4yPFZuIWcQWtAHqHNQvKawgs3tk3qeqd2D
7LDo72WGFGsO+cl4cCZ/yYcUzZ/6L2Mz/VMLlW1W6dIln6p8CWpkY5FbW3R5x28FLdAc6TpWn2Yq
NYvOb82jrj4el32gcLv9RDx+ZwEmPt3vq7uQou/OFWz/ugNSNn2OHqtMcmj1rXUsK0Kh1cfLxbP5
jme5SfLK3PLs8tyKbRbS1hZ7V/v5mXWYnWttyZvkGiXrLL+fRICEuWUKD67hxbsOMfnXGQ2DHLTp
MVj5fG55o1eSfC3VPGmGzIaz/0lfIfn8CpBjgZit9SvVtn5UG0EhzcEBUEwKISw971srZ3sEluAL
nztGysZmr+QdmZDIUeh3uStUpH8B6lw0Z8CxAwhVtrehU3pQSKZTMZnp8YSPaOwdy9/svgEfZph2
pvzbp2u3NYimm8jRopEhMdEwaLCnnRAi9qNdCKyOux1BQUiKUdhdJ/k5LIyXW5zRPcW7FNqcH2dV
77TNFcbf+BEhAoCZKgRGCDwnZpQU6jbTaR76xNl2LE2rYSq7HBxIdZuZYlpMDPpLnrXtyw2GNg/Q
JElsyPhmy1kbSNumGbp3XRLGJPE6+w9Fuq95cGJ9Csh2+ktO3wwzzIzbyA+q/Re8Y4OT88tDu6fl
yqXWTQ7tqqnPrSH+bhEimhH2LkV/qbZ6Nxz7Boz0dLhgmGuRN7TJIpmQs5d3bc5eMKzcE4CMmKHA
Hd4gpXpDzl9KYpml2cwofB+86dxzFx+0TnKbTW7sYaW4jLz3Ld43mo3GGiLHiS8Of+JAJ+uMrd+e
iFRNg/JTkzSBugexfelfX4yuY7X3COSNp35ykIOSa10wYChw4M1kzDVf65PiLjvkNBWc6nlPE0CK
44rvNdWDcJNZdIhXs8svrG0UIrZxHlNug1qRUnu66xAiCisSSe8os3ilpMJ2NCqbMbT6MQA5gX6w
/RDCIqW4V5htizpEvfTaIAAipvpFR+El1RovvyObT3wZVFagbuRagLXA2DTC7FZz2Uvr0Vsaloiy
jP9xegNAudgZkzo5y4CN0h8SP5lVFQJSuBnHpCdZ8eHnKDiPgqMFlpX0l28G3chvdal6lyKD0/D+
KGaZG50zc9uD09dyIjVkWKKkkK6aINNqF+b0WyAaOMsePkpNKO+bYzXZzgF+3n16jbz/9D8xNTip
jj7XfMgqoNYuzvV59Z+V9ifVE0Johy3p6ch7fUnS4bhm21OKDVZIjS4F/W4iYYkHbTXno8CD9QZ7
73woic2JcYQ/R+y9hrQArUNnP43cBDZpHxXW4lX0HkW7VcAoEK2Cd8UPeih4wKFK0wQQrdcyIk18
m7ipOtW9UVTu4rkp+kqjbdwWMaCUWMWn+oGxkVqMyGJgFirrFeRzhizJU00la0t5wYLg39ESvbMZ
Zmfq+1iLuu3dBnXqJ+bg0Y17aLEt2I9DWp5TyZlIQ07bA9nlIOtCbbt5zdcapFp5uCLSbtAsAPKP
XECK0f0y3YzjkggtjlhXNrgChgmKDi2dhznK2kvSNVCnMXk+CwCET5wXlHWvzFIe3+NrcHXXLECi
MgKz5jnShQXGvnqoNnjdmykZikHPTRV+jkASxDgi52icVap0o3UdMyHqB9H4tOyoL9mjCqPj/I9X
GQZQqsV2M9mK7pkE+2Xahamm8J+EICKdJTMI+70Sym2pP1C1MF/Z7vkCoz3NQ2PoChJnALPpTXO7
+zYpzFiv816lggbEBTglBGA3LpgFFWFLVqxLuqsL1FkLy82L2hLFjCQN5mJU1zC0TVAjxf2roZSM
h7kkL8CLcbLkkI1OWr6WpE5ZlV9BrtJpn6AZBSt/u/htprp27sGGBrK7squ7So6TdlCkpTHZMVpW
R9kbVLbdVNTfIgysalZuq9Xh4vSc+AYBKx7o9hPd7Cm5rw8sVByq59Pim+PmuoI5dsJl55j54N/y
BwIwmxhdowyFVOAbM4sGTJJN+cEoduTJ4hX73PJTxeYPkYr+3oqal2bUQmVsTzQzdDwKYYCdO1Ky
W/A8gL7NobTXZLbVBULU0bm0b/lPrhDDEqsirUXY4QWLBiVYg4um6knK3hV33rFVR9FivilqBkSx
PtZ+EoHzInERnEz9HiPTMeZL9cB6riMwGkROQLBV05oJFP181bE9luC8WPPFb4DR6CMrMm+aFMIB
7Oq2cqSQnmzbuDrpSwfauQ+dfPU9MDreWdazpiYaiZ+PeWfXdkLa1XYX/qm1+xQkyIm5bPU8NyMk
bOE6eMnBSfnpig8yWw9IyNWKsAt/UggU5BRDz41MSOdEmMlbPWPnj8VUqYGVzwuk7NfFt9Rebo4i
D2HoWq9t0rk0QGhqdVTddi8TgbWFcBhkSJTHRF2k1YhIocGcbfrgoHSx74I9GQo+upinXoXpgSMr
sU8pNpSTkaOMZ+jdEGgUX8hkI0gXZZ/6A9kg6COHjlT7XQvTXnRXAlBjmJWnN/9hvw/wFeNe+VK0
F23mAwuDFebmI7H+m3eu4JlVebPeI60Urp8ljY8JaJm630eA2BiI1l63LKlWBvv9Ufq+PxtQUYux
KArx2/5woxgumkhNkPwDN7Sf+nwICy9QxqA+gF5o7zHI5kOS4WOwbVmCuzdmTt/vDheqoptHUvh0
5EVa3xh4CUN9a7PG4crPvu1wm/RBe6JSJeYCQM4NG0ys2U8DmGHNML1284A4S/JXQix8X32Ifcg9
XwXmaTkMCkyyKTcmeCesnrGVPvgLNBG8IQJcvL9AlvX9/zbq2MtYLEfq7wAA1ipLBpCRt+XNPfv/
b8L3DhpCBmuqJBKjEuGHYlpDZ3QZKjpDzk8tarGdyyiUoHI1pQFHsOlQx5/VRUq/bRFGR0z3HLo0
CsQYCsIYNEI9iaVQATFZLroV9+YSZajxBh2naRt+XCR0+Oq2/EGVD6g6wh/BcS14sJcCqNdXrBG+
oLrqtEozaaIfpVLY2c24msjpXIW+prOD/Tsdq+RVTu8rff9/EB+I2AWtjBHwXp5IapmnjYekE+xt
RZEdYrhSqSDEM82hD8wC5anq0SxVHqhHnKXBo/u5MyNSfFg621Ngp/1yiCB3eoynhvzmHSWDjKDn
q2U+Q/jr/xzRSGt66ehBhImy9HSiYHCLpjherOjqUStpUptcsOcS0RBiTM2Tl6qqCZi0ryR7XL7q
m9Uo/FfkOssxbiY7ZhQI+/Yftm/M0I766AshAOQNIIXKP7Td+qP6JSYAhLJ7pdRLiSXARGocIxp6
9mMrzXefF4d5CNjojXJ0u2Ub0TsBbOJE0MxeAwanESVgEbKxThZAOW+F3gO8RKv41yCowAfepqIV
RLut9sdRGGCmux1KWMHKDhQ/nU1tBmFTyKP8eLcdWOmXdIIydnYdwhjuN3gJHpPz3DnAYARBhpAu
Etk0tS4OoxP1pEaXJ/wJQ9D6+i8kPFeiG3Fsl+z7PediNWgBVKgyzC9oM7EaB9PWiih5ysgkCO8+
LulWRG3y7QaXNwcfp6n39iLiRRsgSVOac6ecUEQJWfF2kAWh1B8N1emJaByt5xrIc4SClzVmFpWS
+sQ1G3CeMGhN2Yn/57AbjmnchsAZThTx2qJv4n/e7T7SdRQsXghcUGO4iJShHj3nJ6pmzqc++mrx
XaRO24PHw5Vd34R7GcyGvOjT5el3BiHr1jOykgUOmm5gK2qd4WuvjnSiIUdYaZiz6I6LBwpjmUYy
H4Pk9YnOfeXMx29JU35mVEYdOdlxkr5dcL+Aa7zELcHjyaacraKvl9LAHyAZ0ZYYinuHjSkFTnxy
S/yscRGTG/uX3zOqOBoiV5JIKkogkmPA7cMrYgafmgYnQBNLEW5xZJw3o2iGgdmupY5PBH0CGZ+4
WI/Isv4eIjoaWdrjujbt1+4gbGOldvgjWydOxByZLsBE0liuMa8B4HWaqVCNaH5u4HO+aTGJf04X
gnDm7EHcRR8tju28MwuuiWdd6Pas3VqYyzZV057Gwqm3y04hyY6CcmrlRLP/UiPweITn2LZhGc5B
eCbcSvZn7R+s/+8cruQMTfhtOe22SCbcOgS4lEzxRGiv+RVE7BBY3URhd6nCAGY+T9sH51oTVtAW
CryaJCE8wNEauBFpiFsvds/3RYi5sJ5VE+mOn+N9qgfn/K2NKXCQmKUAd2S3HNKQEgF6s4QQuWaj
05tmWZzgwzZ0RBJNIaHUYvvtc77GOHRKLE3VAnTzbprRbcyZvvc8berVveUffpBLp8wUd8rVMn9F
pw2RJr+6NmOOiFciN1ssuLWlq6fw8x/aGRLJIS1rs6KxLXhIhFogV5ZSBOYLh4AjCzVwZ2EwdQsd
G6jjg60oUiLWkt3tLmidOGJ0Pzribf6KQvMxVH9YNJRGSY49YgJv1eqyduyvn17ZiKJGOJg4FvEn
q2Ryd3f6viFFmMDr8Qm73shrov8Rxx/trxlxWak/4BKCAZ7HFz+hxsv9bTykPJ8i1ZgjpOyM/rTl
4Jhj20cfgaNy5GzlqSVhkQTr4rvHZz5gtSOlgwd+oMXCOZscL7iUzMQ7mpQ33H8TgpswAK5uTZgF
Pvr7EhgpuJkt2mLqOYvCgi0GljXGngy9D2JSl2nLFPij9I64goNLEkp0KBnDIoexuxshP9x3P+1X
gZs1GVdWDEPkzmMHR5oG/kVnMi5eScE7BMJHu2sq125I/1Z5O51fo7X2Ur5Y58bsh3Fj8+V1VICM
sniysu7dwu8sU/guPH8WLQDPbDxemEmGWi/BMus8eY6ebHHv2VGLumWrb+ct7Cs7Bn1QFiq4lbTe
UXPvaiDs6RgTlntCuOKgSMEw/4IwGb/+zy+7VFAvfBp+6E0amfNOb3xVrD8cRjrLLEVbrwvEh6N4
38xl3bpOO3WmvzR8LRLqu7ET6hkYgHDK8fYQc/rZawtPF55PuFzyqMYmjvgFzZBsDTo6oQKAOCv5
KVw1TLT8SnDZGXANEUb/gGiz//1bobQ51qYpM7HKiZvO/W/Y+QPFqi1ltGrUBSGWOxWXJFRD3fyp
EY1qIIhyIiYdrpQ/0+2B7R9sO+qdMhUV99azZXxjAwVWiTJsBOovMasNwqus3A94bmlC7lPZBtPp
LR96pTiHTBUp2iAAL0ig7ne+oy9USpOwUfg+NDnBgKa9xpVmYczwCA/n/R2j2/2QhnYUs6x64bMK
nDxweveY95A+lrfClkAQ2cxCzemah8H5SU+b/8bLJ/bh7QByHzrnzgZUKXj6gp1vfEujNhithY3Y
C1pAIKk0EF7klUm2TnOTmKwgYJPeCJNNWkqF55e95Skx+YXW73f9gvSpQk5Z75M1prQnOliv1o2A
VLCyq3pTO3gcJmiR5zhj7z1xdkAb6NLDGQScD7KhdLGzYfg96GZG0V8V+jrAHgC3WagyL02TIYss
BogHrKIZ085HCtXTGoO+LagnGPc/cVVbh9T7EXNk62WN7A12IMAYgbSPPeoZzFeHg0NEKs3bra/m
fvyEVKSzZP+lKgP2gLnyKLlrwmg7S857hBjUJvvH/yxv1Qs+BErdr0hoExUiQETYdyd8Z8xWxE0e
aKUd6jOM4YLsiJgjTGbRLjC1o4KPxwuCrUYPacFEpEzQRBqBTTapdeZBSImePO4emGdl6o38aQQF
C4JFao2F2u7n+P96buVUqCNRC+iiOl3dt5K8aNdz0Z4wPrnY/b/RmznYaZ/4cPg2P0VkIfyA9C8x
LXbh0E/aC0V1N5wkKAc626neDPivv6sjCFGY3yQnRqZNJS5RJ5zKownqH1Vl55ji7J4gBxD9BLuI
OOGwq0SMfQkpeuHVGPnFvJwoC6xcJpwUn8m/pzbDdYgwgEo/reOLWcUj0bddX0YjwAtPSLyaPGZb
2Mn9t41qYXvzaktjI+jIRLNh7nfhO1emt8kxEgWqfkmW321d/LmtJKSpFGYCNbCAT/llpKsc1eIN
axq4mou3VxSAairS0z/UGretJbg+LorwtWiR6+mwgzAyDye9CNo9ueLEj8F2uLNfKAfrjOdiBA9A
wie3pWfiAKioeBqgPRSHCWo2uOEVV9/mCuBsrJ1jJkLUc0Txj/e71hn+pZ1asMpUP6jK6XyHOYsk
GuRFwgIrkad/Wa4Cxg5+UI3WhWOHSct6/moTWuCBsOZDxPTYpPKa/seKZ1Q/m2BIu/1thFA2RGOS
rmZE4ejbTZHffhTzb52kMDFu81T+NhK3liHom8dUFamQPaciz5ZJ6m85hmX0A28vPPqlr3SQtOEI
iN5k2/msHQauZvAfHFrkxXotl+bf8oogAaGDWzxks7s0JHDmq4REBaOod9LvorURVUEOLv5fpxJs
td9OeswNHOmDK5tPdPZNbOx9nbCkbdqM+v6JG4uqkjJd8Q7fqIsiXWehmCz3psNpi8VlDZHPrt4H
B5W03mfMTzQKgHOwlA9XVC+olHaazyELr1icDZkequ6xX4BsCRAmiDh+I8KaQv+HypirQsIntfrm
TDX4oh4N36DONCs1yNdpN9p1YST2iYe6g0prCiwWvVhTITS/9YqfCuehu2POtyiKCwFjK06B/KKV
qLiZ4uWtJNmwcT5lPLSMBZf3fdvTzYL2Jnkw5ctm0Nf7HzR5XdJ7X8wZfCbjp2e9KHpTnvbZLnO9
S/EjHvBAIA1qLiewO87KShnHBfmvd/tK9TRG8rqyMcd1pcbOeFNAxdVDOs5amvghEx4gfljMKLr5
itZ1+RYURz1V204vhmKQvrvaNOQ1A45slhcRfHy5FDymouUruSkHcD7pXciqCwTorOMC5FFXmFU7
ZJwx0E/uCcfyuYTWATA9HNaSD50lGu62Ap24opk6jZ5sREfVnmyVBwdzwcEv5dG4k+1mgy9AodWo
kY4ME9T0KEKyq3pUkIDi9RQfZAnofZ72Opdyn1x5K/H0T9Up6ojdwN8/B5IWqjEB3e/CP5lnQ4xL
KocdxQM+OSm8wGGhN5xPJAqGji7B4mPlfgatejRoxm8IUyoTISNy58IcXjdId435FSJXM6YHFWvj
Rpajq2ZljyzPr2Vapi+TGd7+pMhLANHdMUJ1RpmHA+bZmVvsgrjRka07cd6z0jCKkzHMVN+DrAl/
tHItf6oQQGj7kCHPip+UwQpGRG+Ms2QBNibrLhbYPl8x8GsWueflTT/AN+32DKF3lB4kPdGf9Fkq
nCBgyW0Ok1udyVDQCms0v/ZSJQu6kltu1ND/BvKk72nk7bvFuTK0C3kJRpwcYS/ci9nWcCXhdIho
weAuiNk0waxuqWE1qqArQnJfPeCpDSzde1Hlka02iiCjdT3I4zu98+rMv8Y1aHHx9PPaIhH00fBv
rv+MqrJKMvq2diPx2JDW88uIpVb09/P7y/twvqBQSUP4WmPpXd5imKZymLSeIgmM8NvAo1L/joWc
2h2cNq/4n81kwQgy2vXEDLTVEKdGH7mM41HeLgtmaIZVpxBNPKdbke0zZ1LzHDTbkjsmPGPdcS16
/2Ri0t4MdPr5GIqOy3+MxF1UkYKjrj4pVYGe8OseDlKOhbwdQitFakr8knHMGlmBIxMNVgx45NdV
CMW2L/CACA5ZG39uwnB9r2ehmtEmxqHlQkYRedPWr55g1iFId4TIEXoFtzscCUJHo4LtA7a8Zdtm
wNMz7xtgJd1HiEhtCrvndNVIt7fsjd8JPWb9t58pG6IzTPDnV04/Rwg2iJvL5cYhnCOjpzq3IbPo
Fk/V7WAHNh9H74ND6opdqOmQ5HPyrWMypdvW0OUuSH6TsRlx7tknI0PRpsS9S1A6xoK4xRgY7Xl8
67EkB+Mr/pgmCuxNOitV0yq/qr05NgvJPn0MITVSw+QK5Qxr5DlxFEx7sgoUneyZCuphGgB+k3Ny
5pUAY73+F7IfK+7o9aflB4TW2Hmn/uCuwaTjYGdlsCLsNEyIowUyPRePkvH9eYpZix64gSOb+OqM
4h6gy38IUYnGXJ+T5l8R5esdcki596X2eol/ymP4gJALOBp6IyyyrPjKyuUU6VrienMmZFqHZkH2
iYMIVguAepaTkjDLXNG0dqP/2KVNz5ZgQn4/0VxXr9mLm4MYFpbIfdNnbSJEoPg6q2aeEPeEMM++
slfGOpYlQEPbANyvcgoHMgTsgp3O3Z2Txq2uYYpixt7iMGz4qZ2dB+kW8E/S0tp9eJjuhl3iPZm/
/V1K754Fers1NztP0FQ1lRtNwM9dbaau0Hu9+cGBmWR+9QWfoT4KWP2Xxi2sy4TV0Teu34GBuyLM
tiJRMJskjfZMqcRwK7lgKk/3FVYvZrZnPDX/YVvZn/VNPozs/vjPRK91GAYCE3ARlCIUo4n318aG
O8R8cRuAIsiFbqCTxZCXBbeYbFOlPZF7uPH74ATpCm0+y88GfzB8xNq1yi483eiypTgWOwqts07k
EXgDzGSpEt6C+mDG/E3u9FDfS50isS3duqhk7+8tNh9Atu2uGu9CfJd9E9Y5U5l87K64kuQe543Y
N4O20qW9F7drbXMI5gBqUNencEwesoXVdsgCJmCz0uhcEb5T2rDvLXFLfKeMf8YEKSNwAnxk3aaP
Zn7VgT1gzlGRqaIdUqOpr3DOKfdHAlmWoJGL+VRq7j9tvWVewDdr4/pALql1ZNH84Iav5B1mKPhr
QZ95/A5c7TcuwEIXhtR6cSlkEiVYh2Xqw/+VNUdS6YH4BceUXvPJchf3ToRrtoutUReC4UqAubHM
0MX8kh1YO6O4Dq2QqniDC/UpEL3DfcbuwDQZRhXFL8kubxJPp+pxLfamGWpbvFjmA2qa6NWHbIRu
SS9OaBcj0+3gLxLnPzoBuDrauownmDtub+BX5okIHTnHhX7STM5GRoBBYZR5ZTJkG+JqkheOJ6no
aftx2KVXbRg5YS/PU4Dc0iWxK/rFHp6bGr1VwYg0r5PczoX2Gmpz5QZhuKvzNEBWsaQtsmTwPsw2
j83J+BL8l+Sd9xjFY3LaEM8EaFWMhJ5gOq+0B4F1fJ91tWV/blG5E8AmDmHZuGzdvMjJH9FORf6h
iDTFeGzDTqW4UBZAyKiPA/wo6ag+oaHEUdq2CDLfa6RSqD8TtkOs5yFYxmPSnYIVQn5tvfBspNlU
W7utPl9sUzx2qge6ESREsZmgdJSicvn5ULKkR3dREJxYSolGfBRRmscEJUybYVNX8qAuZpCpmK4B
fTWy/XN753WZxxO4paGoJnwYSlFdYgY48Hj0h5AhFujVmD5GfTKD5oJZdYZoCJ8OE2FPvzytxkca
3NqVoht0C3dIMaLWCI4yBGTn0yi63sCWrTCH3alj4nJPQb1UU2aHwfCwI8hcT/4T7ZXlXS9iB/t/
Er57yKFuOI2Eoe9bcHEYdibFlaDZ/JNWgBmkcoh38pdT/o60yAmD4FpptDd2isa2hON4GGvh2Ugy
gdgUDcK5x+3AIUHHVprqojp/HQsdlm/qtvumSzdPl+sXuNdcnFQ4sIKKqFZmCDclxW/DcxwuYbAV
RyJ5mTzNmmTgbna7gZfI3HxRfEhq3Rc0CtVY8QvsEEIflwZChU7mZfnNChQ5+SofkqIXZ3Vb+fM0
oMRT1OxqMLh8+GYRywGSDdr5TO8p1blo9MhXeCOmJuG2PsCUNLh/p//6SB+AJ3CVJiNrigR4gL0q
CyW9mlkA7ek3E5AsMuMH/tETrfkIMDuibHq+sN1xIqhOXViLZBvR0ayjd5Hhy2hK3Kvt6OdY9h6u
JUaM+LZPfHI4L/DbkuGdOpN0rFnmxnAK+w3CJwShtefc/BpNfYQidKfOez/VmtsDDSAsJjt7OsDR
bcOI5b7zh2oDMTRCdqbb4dLTIXakYFb3sD142iJ7J1XE08TiUpZXinyo+pYvs8cxHW06LXUnPTJF
w0nsurzhHOV/EB4Yzw8GwdYXobWHy4aw2kPGcq0XA1SOguiCrOIP5Xw8gcH8cCU7Uk0FMJQzeBFY
68qaVR0zDwuw/hnTVFge+oGSH4lBkGql24fgtEVHqtnlxJ7F8MYJBzU8bTgMl/JZmwAdeHrAWvll
eTUb9FaipEq5A4ToOT/fJ9gWPoBoEZWU9uXEAGfkgllB6wD0hAa+KW6Bs/8VZNyAGOkabAeaYBhV
ygeZtPiDPiAJJ7dHdKCAmPiCdWPIqeC1sFBKuXYPiX5bturDv8TYPmo94m8/RvKudqiXbya38Hni
g5VM62Jx9/JV09YMmsCq7g0q3irkFbD4IUfOJEBqWRk5f4zP1bl69J70+lFpJ6Dr17eaxbz41Ulj
tZDZi3f1dhtyTNTOlTXMSiSW9hWzsSUIwf94jOf0Q3/SgtSHy96Li+mM5IA6/htglmJz+K53suIO
qecIhxUu2WbHsd/D4cZm81c8jVtJFbBp6Kwhly0f2EMyRAYNffgxbwxG+qzSJXsQQPqIHsbJpgK6
OO5lYItGrszmRjl9pfhPP+IUAcI36vHrRmhOZJxwKW114SDeMlJCUQRK5djWXqQ4zCeA3AD5BOFI
mTn43oH+qRO+jmGWTF0P5+4fK/BfB89p9ssjynI4mzkope3wRCZwmfYqZhFz+i5HdaMJddg7n9a4
34vtJglJzF9sFK1aRNLKjszhZgcTSvWGDrtBPcJ7wW8KYrEtvktfHnGqpMizdxZpu3jXdMdIECht
GGcoKXppFD/xcDefZrM3KQU+BEOThd+JvlESsBhIf6hvRinB3Q3PMi0nFrYkcahYPEQTqrUcE7Oe
w0de2Jj1Qi4bnb+kKJpfspVhJYVSN3a9C/phB1qSWE5doOcqkE45/Pg+byvrsGvQbUzLBcTzzMDT
NScnpB1Wk7AigXsmxY0iuER0RKbuFl7VsXQXLvZLlWW1UIi+YkvPnjEuMTZMQ9P0MwptsmC2xyl4
WSrgSg9ktjSQm4NqQendvdXIxTOGprA+IcGf82cGiwmtVg8fTtxj3myv0eRG0JIDfkyVZV8473bH
MpiTKXQMFEpWFq8MCMLRFj0bkLhwffKo/0sxJap9T+KZbVBh22SachgsWyBCl3N49ux2pE89Oxzh
P66RTqjxtu7BJd5vH/IkKw2yb9Lvs091L++yovtWkmsHVLaqJz3ZyTkIkQTtNmGtLj+SMl1XB5lf
wwifZBdQK6LERObnJxAamRIz4aHcInkTse7ITAv/q1ePos5n7IBuevK504vxrcwwQeD2oPHZveDs
Hz10fhkSAzG+XHdQANDb4pgwL/XXLy8ZhYBOeop4vXAPr6VTiRhwg+koaSObCp+FdmgSsfDuEoai
t1rg7V3Ui8rHCHCbdPgEuRd6vEms+R4DwKoYrTEdm3FbdI3w7V8sx/hiQtT96UJSv06w0/qlNwPi
CoSAJN20dV/O2ztuJzUWmyGdBZprcK8w88eRiJIkl3O5LJJDSO1JIAzpW6/NbonbR9cDG9DyfWCu
oFYWag32Cr/g12L+89dwjNk4pCb2+jfF8l3Ff2DSCaqPQtmjgiFiLD68+B400oCov551UmUXAqRw
3dzn6gLzYT9+mdMR5j/5FZCKjEMzhlETkQIew11ADHpMspvnUw1eb2tJ1KLRZurFm8JPskUwrw7b
jY/dtRVLOwscsMbO6xks+p6zLqMrQ6ymwbTHz5hkZnADjWbZ4yaDFYcX9pxDYG9nF2pzGF5gOA4i
D0SrFMdB6FDwRYdQ82vdcFLAmjVc0Scsas2HenplNuD3yWYp2V8kAa/1qz+rJPJA8l+1kb9vHc0g
l+XWorCCsTllsrRpEhVLB3B8M0xI+RkawbEdVJNduqVYqoXz22/nYQrpvXHj22zoSrU0QOLvwydF
chHo7ohbQ33YhKUWPv9y1e+gAJ4yBKDZZni+3f26dEVaDBXmiWRKIdObNmBi04Q7pv+pSO7h2z+e
9PeqHyXs4q8ZSJLbyE1WOuK+DqpwJs5tPCTB8izD2wwvJBwZpyAH7q7E3MBLebQryCKTFKZ5TlgK
I7b1p0auiKb1pj6PIcsszrk52yxDYI9HitrIdGFBGyAp1D5hD8VRT0r0xzwx5r9vZ9lf1mZOumAr
xy7wCtGY3WbXTG85Uzi2/Xf5fA9ipDCHB8MfDhS3qddkQKy6CkWuK7gioAZb/XzyLtPR4FsqFm4R
J158RK16yhmrWa+YIUup/OdehNbcpl4bbYaGwzFzozEGzVc8ZUbYW9ms2jIZc47MPdL5wUDvfGTY
HfrGJtQoCwHxDnrYMz9FjWd4SKCorjXDajbetaFDf9y5l9f8UBcsKK8WF7D4GL5yPr3fWmQJpG5u
KJBnk9BNWTeqT3UTjsRqd2hNtHGlXcWbG7DrXQbowY5eJQ6/qsRzsFSI/Ck4ihXLNDkuFopB7oOj
miuEEnNCvGjG73w0xIBh5BP017/gnYMajnzGIYbgpjmtwIjzHdh9TM2ENTaVdiWCqV7qrcW4l1ej
gW+3MttEMa+WA11WumIMreItYWoU76DfJwMz8Kd0HkoXxBZzUlqEtjDMbVvxL7pd2YNapR/0Gnm3
9SFWOLF8IpIVPFH3a7zd0DonK/yUp2DS7Td3bfDIoY/Ek9fKlkiRK85R0GAUsDs9wOjljj/GGJnZ
OKLDKB0OYU9Cuoy/c5OioBXtd6Us/zPIVATddlBU/4MbiIUr6I3n6TEKf6YB+orZCAnYjKPns0R4
5OXzhsxERerGMzhd0nI7rB2cQHGAehhnm+yRnX4bhNs3SylNYTfZpv57pQBaglQtO0tmu49FMarE
NOaKrcJ04N589kmCR8CW6Pjzj/I+R3yVKN+6HkzlwipwBZBXwNDAZqh0PaQNCcpia0Y0J9Uxznx3
SfT5eh2zFhJk5c4OlHmwkj7w8elPmx3/AjhDtB2zzvk27ubwnTfKnEoPUvNRd/KEs805BjAMYxXZ
1XvoA4CJgeGagDqIsnm4GyK9S/MLIiy3rQ6813gs4ndaovcyADBQ0kMi6J/uZVRBfESZxksBSu7U
trOGR+5GKs0smS9qut9DmvicrW3l6qf1eRKOA5+3wRpxKu3/koz6Pxkht5+4+FfUHtqafWwNob4j
nf/1+LaaVlF8VFk6v9GlwCVtlDNLZA3XCUNPf4arnR/q6+PWFyrwWRMQaWda9uD08FYJ2aHAHsDZ
SnBBbLFDY4FyYs73XdAAtjftpBiTxY/tar9AbW5xXjzm8l6xX/IHjmqGIs6CUpGL1sF0wYcwr6Gv
Vp+uMZUSn1jXlAvRJ5/tIJf8m+rFnQrJn5vYew0HXTAC3TinOh2AeXX2ghZx7jmrHzXkMnv3L/aW
gxyFyP5SBcKT7nU06qpKAWNArszwbIMdMkJZurrwyQgGT2JGEidOhRLpwA/gECSi88rAJZzlKQAX
mocFFp18qlYEaZVyfva9SHkQZp9szbcemnyV3bJke6Eu2WvkqEnHDWVMhDodt92SagBVEaqjfp/l
/ekT00n0/hlKw7i4mgQGVU3Sw0sCqDdTWRV8KYX4SgwCtEO3NMb5OdbHnFgkOJSL6jopjbC347lo
o4gyVExVzemoJXdu5oxDrrjlYx65x0hH3gJ45wn4sLfoPjjkFxBX8i86lt2gc+P1xdhQqr4Vbj3M
NfDlZqBPyThrh1x4ew3g7BtfH6iXsPyyb3c0uVFSj3F/tyMLtshF3R9bd/4Fj2O1EoYgtqM33CKJ
PhEbnUTnvFOqiwMcXXR4x90zca1anxD4pjHnD+jfyYLBdi8zdyOZvPLfXjsGMBnx5lLJK8eHAnM0
KFr0YfEHXeyGYu7IrRvNSjWu4LSJoZ60wM3pzwWg/J+4R9rfUCe8TUm3cqv8hRT1CIaKcfz2JhL+
6K9BMl4D6u9xcsnkvvSrzU4eKTCVPv66v0YHdTMtF22xAXH6NiqQNqswsnh5rE0214G0LsYTAUJu
ozMb4M8oYJ/gPLjl1UewInRZqYdl7P8Bh9Qlw6cJNQ6HUBuGBhoPBiLQ1DdIgSmfd/AfSptnDMsb
aIiUM9C+nWmp2oSLHRr15O0ixJaLvqbqprIFUmrzoWF9jb06ZJTRltSM2ZmD7OLy/YWkvjnKrn/q
B78BoAHARtGiePaUKlrQsHQUndLtq4iz9RtjLrCjckgdIurWyKK7u6IvWClT75cZCMyKxjSPPU9x
bbome9sYQueyTrOan63k1wBXn9fK0jUEpKXPOUfIDQQmeXXh1nZYJAcmQaF1z/o7We2QKsy0xJnh
66wse3Et48YO7dE+XIvIZOCqfvMxbNKYxVF6lTwVrPmUhvALYqMZvXWAItoYTT0vNmNJ7RUrC40c
U0Bv0yPVTfJ2/91YEpMHkSat8A6TsACk24zRs3l8rvSI3wJHejtxCkXSmta6TF87OtXy1iKxHnqr
CbO+irEo69A0NGbgnT5bwsIzk8d7ARb8btUFEohbQ3Cmj4SNqGFFGPvLHv2lBtFPsE1fqDRMUMi6
qJXvdVCYipvKK43kVVpuC9+XxMpZLlMAyhYu/9g2xLVHPdRxNHQc710IggBZ4DXl7PmWdOUWW67C
a8I/GCpZX1S6eqYxZ9N0j1yPD8nAX6pAeoYDwYpLekajL1V7vC0MEFro+C680j4S1OruLctnWYYr
eJFtI/Q9f2mUHFiiVJAIRrTQm0D9mcehKW5PjmlO1Uu+x4GdgazN0a22RNiHiKlmDcmWEXCOSyn4
7N4nO2IbpzJNgYX245InT7yx99cHxl/Ya0tQwCG9+odPjTnbmbzvhMlbHRCO92xlGO4GF/Whlvec
IVSJlGx/nzCa9jmC057GgyfrDq+iKWwWaamFoYcf3ZCA0FC2RrfBgjiV7+yfS9ixB9LtNPqpl/zj
kqEGIOGezOY9yqMCJj3WhZpzSKE0PAjWCHR2oX1d7JZSZhaSKg6svYJZeAS3zVdIwdz1CwsaMPZ0
+Tv0FL6vp6g2/DxGjuFy8F5KXUCM+aEy/quGSEvz8AK5b6RUU2KG4N4qF9gfdUgh+dTQZcKt2N3R
pjJ1qQnXqi9VzvswTZcTvtKdjEKtJGqp4DdJ7KLiEO6jm9UeslwkEpPSXfjTNezViysq4TYQHONN
MJG3zyl7vRjy1wUGdWN4j6xyddYR0xhZmgXChry3MwEDIEz1GQsHdu3OroP3AqYbs7O6jFSEbyte
cuz+g/a8diInhOOmvzMdVolQ3Cd7JluX+sMkWOzx47d42KyDP/CDYt4R8e3aFkz8MNLS3HiOkeIS
HTR8ecD9jTybapm8rlKDpxcVGmkOXfai/Vaf158L5GxjfFP3xCgxSP3l+G8fwuqV2k6L3uiE019r
XwckUExln9saxASrU3QxhNrjDUXbDUkGtX2VXpr8RrpgB3lS0uuCNuOQb2kzkfVrIcjOva6WpR/x
x3wugxVhJQZ3iJfMf7oytgkmG58HpwWEbfeZQixpnk37Eb0w5sVbAggho35q7M5C2qDZPIsPLoRF
G5nOIDQ/JPxk5ZX3J+XhXtj6vFSNGAwjLx7ZT9IJCbXRVRlW9qYjqp6eFw9go9Ms6zCKUl+j7AiD
e6GqHcAMXm0ubBuDEzopNY0RvlX4TiAapXFPQhgnEdHRs6IniMFwuwukE5djCWFfzofnPPH6Obei
pPjkBlbQwQh0XDoP/PwbL90HjFoSIx4BFWe28AD34lhrzVP3RRZdz6q23OWAaGZc4HW/Z3ogpHoZ
UBc0SikYkQh1HqeXRiCv3hFd4LiiowGeWFwc7n8VTSRswB6gZUP4P6NZVzbFlupDLkbj8E3d1Nsa
UTnwm9Eo2VwEjhtECsPOUP+lH/9nQ0xzi/hVYB/k36PRkIfTnsvYhEDSy0oUcgU1ByI2iA8EeDfN
m+SYNAFMMRNnSMjQiGceviG7HTaEcYamEmi6S5krqa685ut/HKXrQ23jl3YjhiiniCIHure0W1vE
xCguCzZ0y/V/SJdylphCjWZYBEpiNOitNywC/fmcYlwlclJdvCCc0BtO0rC2+7MRvoY6JTEjndsS
vcZpZsnuhYV6X6XR27VxwjLxU+bpo5cRsFoMCgp0Oy+vI5lLBZkaZ4Vuma6aV2QL5EMtfStqYGg5
M/ScRHCIoD+LHvdd4Yd2wTRgcG93c66X9SX1dDhvuoCOKbp22qqTEKuG4dCVmOyiacJ38rKrcyEo
bp1GeX/+dhQ28BtxWUGSa6wokqWj1On/1DE1dJkGHMAn6RYi6BcJtdWaWh2099z+GmrvNfNBrqxe
8LLySZShxQ0KYAEpAVYOWIIC7qg4P2HjMRTKx27V/2a28sO6XesL8lubs+XeZ4U+qgO3BHO83Yth
s0zTPKO8v1j9a8eWO4N1KDbFyFTEiFh8Mv/c6VvwODrDFxild1iNcfpEbPc52do/hn9dfBUo0son
kiZ6VqnVDDtMst4EgMVYgj6eefRzetsX8S3HStBGD2GsH8gQogaNHBe7jlaIhrVXmV4C3xYGz3XR
VTxF0UeAygFDAzaviPIMphhCCPxyHGmfEPNm1DouwHzcPOkxnsyKNCZFsv2XkdsjDY6UqvOSkeq2
UfPng2+itPWvSeeNAE/z4Wtimtz74Ie07JVcaznenxD3vPGA1qpc/Q9rknoKh4Z94DhHnErQMvB7
QIxZVvRVglz/M1aBVNXMzxQ2Dr1skO64I/EzCqNwXLpFCrDxZCYkAy8O8dPKrqGv79EXdMWUkQtm
r8QsijBz0Ff+BZG27dg8vBqk5cK5qq+Yy0SlOkJOb20J5HVhIb05cr/mwGQfMRkk9gvdxm8aDR3k
2NeEuGwT4ZYNuno8IqQSgsA2Gy4NI/kFzXN6bATX12MDv3G6VF4l1RCjQpJ4cHVaZkLIjH/qAdRM
PHSwmcMq0cVgX/lX75vCrzLyymsqWdbhswP6Jgc6Nf6KsVlRzsoiSIsbsMcl/uabiL7YtPlj+lc4
pPfhr90ZDYtPIwoRRscBz/8cB9wKdaHqKl5HwhQfLXsHPV5EUcI5pXqFMR/N0oPc/fjVnJmsNe6B
JX2NBRLbysEoDdIRSSl3JteCoPMBLpvjykJ84wcZaaZzVT0fJ9A7hgQK3RxyQWgQ47sKtQuIS8wS
aAaLL1gDm7SVTMyPAZjcktL3aYrKiUVKBlURLXII6/ddovqvJ76nLX9HrnbF5Sw/DVQd1MDIYT5U
NVcC+Wm+Rzka3huvSJXWWYgz2S6tbGatjQy16gPsVG3yFWiJX5Gv7gAspZygo31h+7pb82uq4LjQ
/cMVksdJgCITlhslcIZrENny/z4B4ihIOq0t1183OsH/Jp1jYvxONq3YA2GMw75wAVTjE+SGr3tY
XhkYuI0kphdl454oOrBn9p9iPj9KHdCDuCKxthfbcSS37NEgbbe9Ezyy8jgjyD83ieo4Una7VGlV
rLTxGWAbsNuZCJ5kqpM8qA9eeZ9hBOuZsOx4+JvTa96PTNqP43UJ6og7EaSmTtHB0IXiMggUMVnY
AgPCbmp3tCrUaepX4yMhRL+18RQSKK8qYtb/+d/X2bOCDQNyh4/DK7vs0cY9RrN0VRAEPsTJ/MI+
5bQwBjbNbsEXBaR/i8/qoshMYtIbFfFCPbWtJNhr+S6j0avhlgSIN6ec0o+6Sb5WXMbxLx9K59XT
J/tOGYVgME+H2JuMbxAqessNC5tVVTqB4hWxkl0fi0UvvbXjwBZ6GL9vHF6s8G2A0G3sME2L0oqB
afBZlbDPrNwJf0WyOwT4TU5UQCBaCjQk9NsqjrnFkbwejrbcc7BhRYV6Wc2Y6FZoG5+/cTHJS1up
aES4Udm0ufek/h6TzrpYvQNlsUyziAYvjYojAvg+gBN0h/KPdpQr1jBru+7Xg436UhGwK1bxaevq
Fy2LcdL95zik6fcMd6mDjj7SojgySJiJKprB9Hb4f6JUXntrZnONR7/foO5Pdo7DXWGtnfg7Pdi2
LZVhnXxlPzfIrqAl627jfmx5L/m892oCJ3ywpS9BABHXUZs/4MPJJxEvICKoHFIMcsAURKW+l9eO
KKzg+8yto0xEGLmQBbFq7WkEN6BATbZ+EjgQon1vZ4d7MBlnsEbaFVeqI6WnScOcTc0+VITOAjGO
DASI71Y3sVBvaSQRcUU23L21imLC6tuYNOKF4+XkgcY4R7stjESwcnteXsSidfz1qkdNB5r8C2H7
PfiYSIeiwN4NJ04BE8Hhg47/ku3C1+vihzhiahFzYPu01+BUIrEDcC49M+tll1+jdHFdk7BhfZw3
kKebAkvkT+HCEV5/+Zyf+C4sH9F0iyIsq/L5zXzD3zAbCR4venP+uQeijRFHOLXKA63MC+Li3qxh
dcyBzs+2Qftdn339/PPUr2TcpBat7Ry2JNl56ULfDENGtjBUWmtOTLDCJmi0fPgjOrVoxiFc2hiQ
Z2eEIQV0Yl4Lmc0DW5/Ct8P5aPIWfA5ZzzpwmsuZlRbFakTgMgZHu2FZ6bbnvOK7HEQX/Ye6z7m5
sQU2fi+ixU+D/ipTebbTu9jNStgED6VzjSA0COtzGPiQpubcOyc+yVfDlGhNuK5P+I/8La5l1eNc
veVAdmfvmPT8Jh26IoMWCsBb2ZeFuRFvC85wMZ7yUmy7xG4lp40ik9mj7vMjPYoYoiXtKtG4NpmM
ip328GBFdPXCJ1upPEppRie1g34PKhxgdAo/Hxp6JSMKnb+ewEjpQAExMtH/RrwK/yyER+xZHzLB
3x6gxkdgFgVnzwHXQ1njWhTKH652dXcDW8Jvz1YkwUMMzzkw7L+nIdj00qG1pQ/jfrY40xfS9C7Q
FOrD6zcw3NWIUmwJVjwODoFGrXzsGa6Y711v1fElfSDn39YygY2DE9BTknaJwcvk55xMPlF0u97/
6GLxjJfIZVbfRjtUhNffMRPIrZ4c8gI3TDclziJaMe7FktIBarCS5KllndDwYTTewup3dced6+Q5
mY+hdamGaz9z/Q/J1MJO4G/Hf0pQUxbpoiSgoXo2Os9CHAcBjH7+vJm1jQyd8eefzvjwNkv6AbQu
enO4nN7Cy1J5yrkXX8lLAObfx7vX2faLKjsihq5yTFUvMPOvNq9QJEM9aoWPoGs9lPo9qkhijuUE
3NQUK4a1yWtEuZF+hxGerYorRTzvvrSTjNqTPJS3yozSl0auEumAUu0VbIQuncIb+5MrVPg76cIP
iC6Ex+95eAXdiW1kgZnJckz786ZChYKRGCMkLci+lumXlI7S5gdS4TakdhuLCzDFFa3Jps+z8+ht
uz2d6v4G+W8QKZRXmPH7bG2/QOPeGeSwpS+6KOBDUSUCys2VVLeRwpK//ohl6yJ2maC+JjSV2oF9
fRKjA/BtBwEQ/y6BtEzrKRGuRYMhPuV330TMJ8OA0sUg4Jlx33N7MfNMhOIrCab6u9kccUQFmsKh
Dt1928RcOba0GSYPvGtnoOS77v783I1fAPdBetM/fc/CorTZRlXbUbRqmwzUxNpTgODdztSuMJi1
3UGyRfBVsYtthJ5DbTgfBWPdu+1D+YRlzc3uzG8QogtMvCQJ8dPW9etC8AmJeX4cCq9ZAvNmv/vl
lu9gehiLNivbpbXec+c+dIGaKKfMgBCM24eKqxqNLzOnKS+eYAttC7kKq3a+1Q3oXkDSGXZpZpm0
IxD5zYJzQP5JMcma+OUBS3mnnb4kpFrQciGvJPSIGxr1brIXYZTvxCnC3mZ+t1R8BoitjqG3Js1C
S39H99EtcZD3QG2xy2vliExYl6is852bRz7aRFaY4m53B9UzrbybAYwSSZtd0azgblu6KcSJCxeL
wzDvMlFCAiyJJdx/oCtnCHBahfNQ/1oXnQsUsKKD19UsbRnd0hNhu6kt1m6GQjM1nhglDWR0MwBV
kDZ1USyEX8OS69/7uc0HF6oyqv9gDaGTxYfcewT5j1bRyZZ+bhlcoGQRuhfYAEAOrCPlhVaNWqG4
rh9tcpA6KfvWhowAWZmc7MoAuy9b1YGyxjR+uCKTqSBM9Sx81SC17W/6PqAjKhBac7tsMR9pc82u
fXyZAFb1csIDb2861MIrK1ULXoTEk/pUYJmdTjUh8c2lH80gYPUdglhMel2p7Z603C9/pjdhHr1N
uRKSSqjyPZMO/tNln4zpwRzoNv3HbtezNCjp8mFpFkkIx6IvOUmalMCoY2M+7xrRzlVfBCRNQ5eH
BrrsJW9HGNQztQtaKeNMBXqCF2rJCXeoVmf5jndARTYsa3fpLdg9jBWI84KFpurU4oM/bn+o2Rei
WshqC09YOuZ7yKYDIgRCfp19QffM1zFVmmdhuIOHi3pMFyegh8ARuJGUxOJUU8B5EI36jSCPW4RG
vteFVR5lr1M8bP/NktptjPn2eJEEXt+HvV06Jxiv9aw5kfIpFKtYmGGHAmBBRNbKp9ZE9vJRudh2
XUMfd+34/6/5gjqsohjseS26KjSrdgysJS9OQ1DHnRiZcb/8TLCimrrmaDrFJVRmgwV1Y/bnirdl
bfIeDD5PJOe8fFPUpr1tqd4tQS/SVqyX2LVM7J0KDKm78B9PiC0YEx6yI+dpYaSU4fJWnzobvpOC
D1jeuesNqZB3tIFfVAJJowVIq0QZ1VAagqFbF4AXSHLPM/bZlYMVekVNNi3TPu+N/JCDxLXteP7E
0jaPnpTfGdhEJhh9khEbTlD1BYLJ3Os6h7zTS1tNbuLrtB1eMTkQlMtACxgB+GW/uG4PKJ3FU/bX
2HBuutjwCQiLUzy6uxn/Oqb3m9MCAjHS2T2eRSYLh3FR1f9VS0ezl4MD7+qXJb3GGClWkz8Svc3t
uPg+ou1o2jg7XYg5DR8lTgBmyM2KXU7N671AFwuE4j/qirTNH1ppcbdOCDXw1Dtpn4YhkOzpWy7y
keFy62pBhgTZlkUn4fW/IPNiF/ryJNI2FeY6PUdZuGNXmlynxrwv22yvnPZKJmyddPEeMRO+88Hg
P95PBR5I66xFiJ02CnMo5bTOy0kRcxGD5BRHjeKxcqbf+NZ4BQybYUFjEJ2xn3opJU0Dv6rwB67O
oW621Pr8MXzQBFmVUJm/4Eflp1uhhqhwsnlXijCR5r1clnQU6ugwu/FELixzfX09N10gQKk0RBlw
wAGVFYTqR7ob8/IYSDQYC5OmEfjdgNmOM3VhvVVVTj73gBhpW5sbNQuz12OZg/yAYQ98MnPJmp1s
74A6JxegGhgP+XS3YUF2H0LsLqFq0pp3PiST4X+xmesTTlfNq9+BVfxVFHFo/MzNpDsEGdj39xAf
eYLO/KlXhDFKKc+NbwWAGAArn0c1jwj04ZaNCFPd3Hne4iUZV0q2gT+YI0a0Lq6e7RGxBOCv9DCg
KCpXrT6xvB2XarlQingnCIHaavDgq+J7wInNsTnuPOnFHooS0zj/MPqzuq4OeFwDNXhN5pqJ0yL6
yR6Q7GFIs0HKTqw3Ytc+OeMq5ih1dzPe8sJ0yyyPdA3xZUQH2ov0nKNnLRq1QhlM8jrTIMHeT8Xx
NgYzyomVrf4SchY2Nk1pz5i06wOS1eryCqZTSJEv2uBM7Vd7Ly81k8aA/qoh/dcdtzhWRNFapy1N
lN3NdYiSY0XrJqP0dOKheqnSMLR5AK9ztPGHJrEwqB55dtgiKOFDPTUUNeKiUDvjRSsRyUgDQ2xQ
lfBgji4kEDueYM7hY/fKGO/IRT/jP0zFVwqDxDQhZsKq0t0vl5ESjetG1zzgzo5/WBEjAJ9+dXiL
NC6UQosLWJO2D9UekZHE/mpRB1FNibWnFXbF36AXWRLGWmUwVcj2Wn9F+gm9sk/luAAdletmCxIp
mvAbm8X5VEezZ5TeJKCnn7Y8kb6Tnz5K5P1BnOFIbqTEI2RZ32OhX0IYCOlNNlYXOlXxrVe5D0LC
p0EN103idUvOhbM2CzyOtdGTQEjs6DOl1sEbkr6smie2sY787IqHNIMdYHAG9gjIJKwNqTZ7oxXK
HM/cA5F8BNUpw7z2T6fSlGDJS5uKc5SQ/UQSw0gLlaD+ucU+PWUFFES8mPT6b3o5N6qp19TTKDB6
K+8euy3Y/rtXZplJ17F7myi90ifhudAA2eKSGpO+vPb+lNbv1kM5kUn97puMkSAPcnWY3L7zvVlh
N88yia9euDfMJ6PckpnieLAlvx6Y7ABYUo7t7xo3wXKKtNMzKFXLPDLQvqa2y8VZf/c0IFxSmvu4
TDyYaTyf0YnEAVZH9IYwn0Ihuur4IQitSpAFdUuXjtMg5tQk27QuvjD7vpyNo7ac4/AA8Yt2gbdV
/P0XBo4vCm5xrt8R4uGAsB2N6dERtvz0+q/p4vE22954CD27JbW9gNCaDQvXNyX3rCdnvIZKgM1k
e/nMbPmEX8MlkdJHjpYL3KyM+sOEQ/2v2m6OlWQpF9XGpjohmdMOB/fOBZWJGrCWg/UmdH9rndKC
kRjxK9t2fps763wWRuqr+qeXLeatWAX+9ybmZ3RMVdLgIEjvYIT+inS51eBHR87vqBZ14RkU/83V
RzxD+jUGUxko9oOFDLYjQinbuS+bjI08GYSJ0kB3EwA+VFImunG2mrkZafdqIakN7RNsCHsRP2Vd
V5kD16yos/iaWPLX7rM4bnar07mXz9HzVRh5U8vj6d94pUJgemx0R6uUz/l2onItZxbCbm2eWh+M
e9Sjhh2TL4kA2/CJ7E8jWCmRbkMPiZr9q8RrfgyDyjNe/zDWBs+zShgz3YuXHufXIqNYMCWKrzvH
+hqKxUgytaECKhkHxGelNQhhGZEW+gqHWASGORodU0ea6e26ET1nB6U128D8fj6XIOhJyuTgJXjt
DgnIDKMGjhEiJjlQX1ihnQd94V+zij3jyMjNMaYhoAPQdmReB/SRA62BwKybLc1J6Xb+QGq/eXPv
ols0LTO+e1TswDNvCzSBGkW7dusif4QEaOlZ6h2DTspfDy2nr3VEj1Jok/YzipbNKojvCYQVwAc0
B8mcRQPi0JkaW1Y0yWqn1BEGcxLMTYAaGSs2kQplGl9mYE/znE4Ky+w0KjcqVS5upc7zf1mIddJM
kDmMxGAwaiG2f6uOOJBNEYBSDTCBS1hy8C3bWiX1dr3TOUeP/PlYIPdFlxFtqDUeIOB4vqJkh1Vn
VT4OInjDDhTeu9sN72jNMlDxoq62bpziZUUb8mA3UXvHFvoET1v0on0gpUUMzOPqG2d/9InaR0wU
VyjRTEQyOyVHceT4ufFQVWfGf09M5ZzrTBaTf4WxHXvuS58h86/alzWKq3AL6STGZTIG4pcYnzlb
JDWnA14Utp652raU/f+cHRx7/8FUlCtGKLqCrfIyfO/lAXRfsJ3e8tKj5bdYqX3FBI7TyqK0bqWH
srzYBcXTotPUDNGXbf8sc1DWsEghjtRblut6Zc1P1Wywfx2rq3B8Q8E6TsHwLmSi1sipbi7ND8JC
cecygBEqyBTC7881ERhImjTL1Np1FoR1dzERhVKyc251Jc8rnrjJ8sx4X16sNcIzf82W2FgpMw5Z
jtbgxMTHO/oXAc16SxupXYB9APTwYyPkfL/HEJB4KFourK6PKgi/AhfGHoqVJ4cjceb7UOgLsfgQ
uBFY+Wb+73LPVpJaUAHkJAQnazR9VrLKVja9kLrsETociL3OIcaENR+yhXOwkFQbvg0u7bJmomlb
jmhELWu1dwzvGEgpzC6+UO1jkhZaBTDkzrSbwVZaS8PdbaHffNfQ64bt45nk5UNpcZxwbma91m5p
5cqXduAqeTzmUceT54axhDKQ28PlRGJxnh31Adw9GyEz4DjfNXR5NEEFS+53E9/4faMm2h9kZRZx
TgNJXI97D399MFBGWogUYUmxk+HhJysvkK6PDFbIpxMN8W28y7hsSkYGZevifdwHEiEPf1mGzImF
FghIma3sSrQdrogIJlTNFyeMPRRO72s4rmoeTNYwKRh55k5KF+l6j/d/4Vrzgk1ljd0p9lQbSlZ+
UE4p1pJ6U7xr24WygMF9WJOmK1VY8asi6T2jj9qs2fPcfl4qoyuRnGWHG4LcTr06K3uR795S8bGI
a7PnfJOOBSq3W3Zs/TRdSnwULq11l4pLha3y/A0YVJtQ+HuAqDyy88ELcJvJV2ACVcPThlpi1CXU
2BiGR/lueV+i0GnZS6uuGypPBcs4o9GYvTsV7tg6J/xMVcHII/mPM6QErecIWrctyqbbt0dE/ob4
R6w411N0EQz39feD0AHCTr26QA2aurXfIRnT1oHjMlqPGcBlYzkUNebc1xZC0G461Rlo+m+SAk6i
xmiw0A70jOfhCSugR+dF7gELppo8mknNy/dD2W2MZ6SajmI5I5/OpsAFsLlYFW/4PLFWH3lseshP
JLER1xW/E1a5p8sEPZvCz7LLbYty3oPWcj257IgL5Nfr4Ot93qoeKOr8/4/YwpesO+UM2cBKMJKo
P11x5yUEM1DTmKaGsJOVL+a+Ff2H35gZ0qTQO04at5KU4AjvVzbA1cwWqWll6VBSy9v2sKZ8Q996
FoWhbyH7RyaZx77MEnstv5r82YRP948qpGVDXcU+gTpyjTxQocY0jnq0RKiq5T8T4DowidJGhHlB
Ilm1NvyB9NuFBlkfOn2DI1v+gjAr0Vi+ZwBIkug5oN0Wr9fWFthK0kcOd3naAMUM9Ku/Fa7r7ZvW
DPqpIRe9s7trZg3QqJlcumsZeK+yH5GQxBI5Q9lacgQsGdu2DDl1HhqdXiyHnjqBaL3i9LXRa1Xe
wIYMGDWRq0Rr9+cCU4B/vAlh44F7NeKo2ZwEonc8AS7x6lOVfr+H6iVAMxJZ+4mnhqmb5cE6Dzaa
gDCbnqanvtia1u8ShOtMXtnBydNe2feMBPBx9m42LZu6rNqnTDrOKriXbp/6eI3DTXuZ/DS5+Ezo
X0gtXcTTX6u3uil9O6Zn3JSHTa3U6OPWaVGN7JFvIur/Rta7folWrqV0xMUTsvweOb++JFkXWb44
XNX8DAUmSvqzEB2YlPcLGRXsSJnI3OT7O1SS0p72L6a+OIlhnXFJIJMs5KEq/zcfA5h2pr2susr6
b/POUfboQQwcc0+LvilkoAi47bYUPCw89W6tNr8vvr30fZuni2pccaUXZG11V7wKjBqcRT+eTT6Y
37cemvO/3oZ9VJl9kOfJuFA46/KA/zjt+6qlOtCNYZ8moHL1jX1JYzyq+KqBXSXQDpGeM+B1E824
HLes+uqsOpSp0Vsa0/kxTle13KLrHX7LT3yUhlYT4qTehO7o3CBBrtoE5EPO5KdZynfYqI6Gv6h6
l6A9fRAZbKuvyX0HW9y0wSle3zMqjYD1PrpJ3iVBAj8wKbZHlCA8GRjeQAiTuB7skjzIsllHwOAC
1MImE+H96P1azywCvGAsZMTkJq3rdHGg6xeq+FaF5zR2/Ra3ge91a0RwAa3cAqmxBgAblg8u5Uwu
zhNL/Rg+KmZGgdTFPXperL+NCdJeZxCEpOJnU3EIJTul/782JtLa/vn+nZLELjIYbb32ArB2lSSY
QpbLAXi9M00oTMjYIOSWNX+8sT2PzJm4EY4ltqFCOJvEBrVE9kKJZwDfsWixBcB+AmvZmtWEBwDY
mFabWOvaEXXRUkL9iiatDzVflDaz5fYymNBCPJicT+tSPwQAvN6L3Sw/7DlxEUPeW8Qfo6RnKwi8
b5Ywzf2dnr7KYtFqwwoNyCNbVzyK82ZFgmMQUwheEVCMPUn8VoiEV3pTzSbKUP4ZS4PQWNs3hil4
O7p/nSRujRjzmNJMu1wtFBg0OWUWVQ1JPeXjGuN5+Akb80zcdKIi67tpWXN5zBOfo9InOXrCsV0v
Hpam0BV7f5majtqfFP3t+9IFN6kQZSQohsf4zdujWB5oNs1+0UyGzhVq0OD07htZfbe4OmJFtjas
L6TyioI8Mz+SsqdFQTYp1GaQI1AFFtNIbkfNxKcJx6vAdDdbs++eE0GTjZLSzh91nXEzs+/2WEz9
HXurYPBme1GZckBAfXssVXpIIZUYNrXeNfMYQwVSUSNPubErU8Uo0FSfxo5jDhi1gBGjnpfNovSt
7Xrz1t7RBL1SqIEGGykNqxaWt5aTdljHViL6CLrc56M3JFe1tzb63CbEZM8MJMDgWhBlQNqT6dgF
sSNrPqw9ZS2NJ71G+Rn/6M62XLwNTHOlamHk4G3/7QIVR06ot7a5c42sYCgKYQP7N8wS45gpHsAH
5v5XxLeet3K7MQE4E4jCXroCH7MYoh1onbsWCef5S7B0ZgC/WoPBZWYQ2JxxhWRBgud++HcFAjqZ
vPJajiR/u/4jb47qo4LRbrBYUwSDeQgbFSIYo7QxXp0jNuXRTJgjI8EDtIIPQLnSYMuJIeFbjhAR
yq3Y/uycpMT41jv6LloYpnFdSwZRs+54LMho2PwT0VkS+91A0lY+TUMKnW/kMQ6CNXdINcgfrAEq
zvjYgLvjYDZzuexJMFoiTAOVPpyXKJyuGJfeKXFG3dIj8Aqy4HbV7tPvms0L1kuC6hxlLkxHM5ye
ggiPo8RJePDcEjfGeL2zzcBvRsyxcLO+sPxygG8EnloqyAOZ46tZGFT6mCdyIfl4WSZ3exynzWhn
kSfEjZv4IFDyJmc/CUobCm0UmHy2fF9AMOho48TV/5R8g0lJDxgulbT1yRVReIGYKK86ft9ZRlhL
daEV+QGCSRAuHiDrgmbCW046Yt5+L/RCuCjasdTSSbE1hgSTbiaKNUf8Ts8VZ/F0/RQB+FpA6Irr
ZiJNvE0QaEl7RNOyPoe3EBGqiTGr29uBaGOch/8GjMRf4WTJ/QNL11HyjhVE+g0Mj3b2N8x3RMtv
aG60bZx81b+g0EDFJ0mjMalv+mofQpX2TQyaz8xxW3xW/7H9jtJpOBzo0pOtAG9ss9ZPaAGY/gVH
bvpReSCrvunV2ZhMHBtyMvjcfnhKFrAaFZ8IdtwmtaMawxEuKd4HC8/AjXjBokyrwHlFh1qjDtyC
Mq7o64J33so9teQ1U8KZKY1q7XSY1jjuvkwi2ieijxSM/+ynCv8g3inb3+vX1y40kv0d0TTxB1kI
ppiNMzXLoJKmy7JufEFIGi5BLEngMZj/gG6+RRIFeR9c8MhL7miNrWGfz1IQ+ShbpkKRdp3t14hu
ijQtuppNuDfQHt4ikUz+lFr/Y07324fWo+zuuWjCUtaHL/yLopfAUh5QUrdR4d01M8J0Jj4bnAVx
qq2pMTvAY10JGVR2UUNKB6nCXKrVa1Jd9JWTHn7CUhsotkDuqBmleChGKXRa9jzE5/zCCFLKFG57
vnx7Oa1YELBGCR5gqrhNbi8l9s/dee/Cwnyzx+wIWN7pkFEbJBMQ/UmAqvntzxj9esafl9Z8blm+
DzDr2jOOnOd3iC8JDknYYPkO+C0kPSjO5KtrBqREwVynPy88clRXvcdK4rzUi2b7TZSnD1zDuLNu
z5gPEvdUP1+JUrDcrZnxKkJoc5xk+Sn1WMDeW/R+lD75aqwGcwGDkTx/WUE1hc/0SscjUFdb1fLX
V83jh1grnJYy8V1eBlrLxcmCdmSpnfh+sccWgrhfftww93VdrXdBpYhP7f5nXnH3nW3IrXNzgnfm
dKOq6BGr3LmVshKDE/Bsuy6m29jCXDWcDGoL3Ms7PJ6TYHo1IuaORoLrOU+CH3eKudG9MiYLtgZD
qKfSA2PpErUzBdwVSKNkOoVttm3CNsHmKfBC11aFllqamcLGMmqdinH4QXOBsWZH8MyOITr1XMUK
hOv9b1h537Ch5dHg7Us8WGKSiePTNpoJyH8fZH4C18osyai0gx8owx300eqLx65g66SV8hrpWAJy
DGc8/qPs6n5crqoPww1iGPFtNMbnPxxsBRL1rAp+SPFlA5jZE5D0Zvw2jmL1qFpgoPw/argF2S1D
Fn6XLcALHWsaF1Yij5GrctOshPqXgC1WSq1D2orLZv5v+RNGRBLgkuQDrYBcYIUsw5CQGvl9fqYo
egs2EBkXHgpV1lUA1UZHSuZeRntsYTHac5pQINCvlJXEOqzT6ZF1/X1REbltK6d4ON6IeKHR2Vqz
D4T71/TUXgt08l2k+5muzsVVzgA9Cu4bEuycJRULzYK6UjleJI1+3gF0eThUFRFklc3qcpMAqk+l
YNLiV9QFAcW6FzYIWB58bJl0hRdvHRSZWRVujZRVRe2/wVamafuFbEqIVccIyb6E7RmtN8la7z3M
bSYoEzpp13rpdyQjYVccD3MY4p0lN2L6vuTn2m5Pzl3VRhKgbCVEfBzJ/XcMejcgKWbVsUX1o4+q
bPiCI6WsXPezs+6WYtHd2UE/u5COcPupBO63tkVLLhfoYFsul21Q/pTCG5b2ydv1B/GXej7UfnZO
hH3ZZU3PraWWIylUUANHGgTNuPVsz2ugJ4u7Pek+hNpaTu0+f/LKC0Mve2ZhKrRt9b2zGxWav5pA
MtKGLCvm+hSES2LQqJizWVN+L2dkOSJEjoOegxHcGxy48+G/ET9Kqoe2CqRF2YeizUKwaoFesOBC
KnDilYaT2UGmVVRrnseJlh1OKCcmrby/6QW72Hz7vbOdLCMlipclwE3s75wva3+vVA5KzDB98n91
by731/sFeHP2kwJI8Jc2w/VDkfIakVGn0aFhEOTvm4Eyn453+4eKV0rVDze5VvzcpCXYNg0vraF9
XiSUGGvNKzScEOvnvJHXBlaoqWY9l1cev/t2lLhOgYDx7RcZ9iulxJklPhNdxFDvn/MCJReQlGAU
6YPd5UmInKeGj6pA7J0q8Eg4YHBftcvaxRmOAUTNLwpeBV+HZBYWGXunClT8s64wgiHFHaJgxMMG
4y6SxIwDhb3hbeqdBBp1CVxc57R8MrKudDJc0a7QZANIWCyURaL/gmGkT74A1LDeMZa14QeCD94F
Qp6nEucjxMkXmKZ16YqGUu6PKUAW1ZTfVVuPRmLOnBcvT9f75r9nxxVaema7fPlE1JYBp+O0BbDB
NOlwqaysQh0PTtKA7QvDXZL0t65cTQsiFZMvvDQyEscWbSrtU217Jao8ViBpAfNVO67hjFHNhcQY
389Pt/bKj17XuH9hodh8nFyYf4neOTWxeISYr3kQc3vg58bGG/SA65EWwBKeAYPPTlTD0b3EP+4Z
+7x8EYxJr0J/+Jb6OAmALTnzC/TJuXDEuCbjbC838d9SZopFZ9G3C21ZOkc5yFPLJRGgpTDP8UXs
4Oyut69XjSEV5ZXQG/km/yc9LQwLgWiKrzSCdH1UniE0+rlvXEN6cfviqyPGucY5ELDmDc6ip073
WurPJKjzr+tWRZGybLqwYdIw1/RtITrtOW6p+kn5Oglm5yL3SeLHx7i6XVnaTpHgGaBElGpCyhsW
l/Sa8CkVsK5vDpLI0MKIQlKsdfKu7bCDEXjmDGv5SuBO7qa9t0vXtg8+lpTFIjUW9vaCnTWtSJxl
ERgk7E2vNMjwRp1xb2jsyLn11ZuEZn2IhaoqyqbPgnkFXnu8p6whGQDjl/kvbgRHPCIvz4VS5Trf
ylKkv7+0c3F+0WbicY+lDo6P38J4tUma79wqP8hedSJaCw7c+KR7zTDhWHf150+L4RzBR5Cqmj9d
za485D2h968OtLac/P6IdCKF8XJpeP1E5xV7puFQz6tz7ZcctCUPLhhhKlCmQ7oUJbxxT7LPRy8U
v0np3DwM9AVZe1gVBY9mp9V2YWrf/8VJBa6+06MZuezdWzxYZoVhb5+jO1OQ2amD4BmoRosVGAoo
Cjf90XxArxz+elwl2c5KkyWJz7+aQg2k1jkbFkbDumeSwu3vGhfcxe7TjEiMl7yGE7UMMH8nXtBW
XFlOSMrJesZehHuCHkbkoOK0GSx98+go6nSyRdWux8qz8GLOC8lEhgrPfGFbesfKXkibXT0kGdNT
efZYcWpgsUbAJW0ebkjAmyRPcT7gTW4sMLH/5xVgsc7qlQ4wR/tR+5Skp/iEjRwZNpyVWTJZjOIo
HDdEsXCly7ctjnTJtjChr8qAyE8mka4t6zMbUsX/nc7b7vRzBGDcUB8A8xgILUPYlQnys7b5aJ67
lk1VW8i6eBG3TtDRfZjVLUXUPgpNM1HkuyuRovBCPe+eobWEh0BUbK19ccqdlQFfJAS/71SHBGXm
fVpRGimmrPlCa5NlARmUY8oeDrsVW5orFu2HdKkbygNi8F136RxViB9m3hD9tLc2QsSAomMSuzsM
jcJqUzdHeoUfY6pSbfnstzux9yOVDg6YA3fIwIfw/8lcPbf12Zs8nKsawl7wKk4nmXQqo14+wrG5
+nI+3GZhmPBUCaHYKXSbtmRqq8hsMQo2hfbayrtPe4K8jWzZkzoQyaxfeJPx35z9W+YA4hV4dVPt
guFmyqrUjKAT7/0gb2EccM5sYLSm7T2U2Cbcnu8ShRmWCzLLOdFhcfN7YRNpEFHUkBHkWaOKYBJp
1d64aaUcNIMRDF0k9avgPaPjk3YXcSt89qW0dIUktQzcyZbcsjJ0eIKGBtMRCCzjwA+9a3/noCY4
4TEydiA1NPm6aUtBns/J4RJS4c0qZ4J0jcWQeggpXuCkbuTX/DfezkBsoQDgtJxwSgAVmcOzjIeb
/LqyjvqHwriBNYkofBCG5awcWr21ytC6jpStjwMzMuxGaThduCH4hoxFSkJuiZhgjD9QEYSLmWjX
r0T1A9Sjy6UEBYwcpvsgXmU628T6UwexvCNg+wt21wEHqLWkyVAAlIXGEcC2e90xYnJo75qa315U
K9+AtkfFKHaiHrcWHono78b+aBiTsbEarSavMAFw5T5Bw4GFJDkWRB7F1+guMx8Wx2NfC7aN41uI
dSCnmS34b+dvSqZC3OJLmZz40AQtYrRSNci9Sc32D+SMvNPgLZ2V2WysHusJo3EwDnGxzclzOUEL
pdBZtRhb671IFixPyI5eiJEYKmi6hjVCeE+b7VpvCyMyqDikfvQ/T9YNifYaNM9M1QdbQALaDhvA
XhrzW2WBfsGUPYUjNf6eIiOa29RoFKyHE9LhIGXecmNXibezJkYEJhB0EeZWBWKirdQahgIseIGW
asjRjc8vamm0c9/Irgx89lT9FDR/krfIbKHFZpEc94pgCdZRHAAognS5RwLvSr8Vb2cCQBwh4JaQ
VmZQUKDir2Cxh+cYopPhZPka1KLn54+IV7j6jazY1JxObXt7PESO15ym3TBoLsP0OYp9FewvLSLA
Utao4vU5kThk5/XTglG5LRLLIM97fBNM2wF5Rke5VeT+aW+83xT1gXE0ZGqN1bdagJiSQ4Bp+1hr
8Exgglnzu7dXScWitEfDeIHRZ/pEIi7XL3YjVQx04rCXTM+JU49naM4v0t51eWRFSuJJATgQEhu5
eRVEbRRiSM00GobrnJruckMV6ssnGiByne7fM4emaPG9bjjEzQKno0PQQNPy6skC/E0ZN99TlAd2
zPy/PFlofctmdPN3t6fivQ467nsuWsmfYjgFeXQCGVcUSu61Vb++u5DpoAemWcAtocW6tQlW8mcR
xh8CnJp+DvGSBvhf5tLhslGWXmYcnGis+YPK9oF9xUEox1haKyMPWZUOqsISNeyZJQyRQWutm5yV
RfRFZsjkMTond+E+uJMgm/BwmjUjHFgNPshl31caijSU1w7o2zoxDDM9qYof0Psw31GHLEGLmFdg
AvRIcB1byt9zafcgXYCGSnH9PZLXRFocktNzjfEExmFvV1CU3MTA7gDgKLn/GnJ+Y+Fmf+W2bIkZ
8mvv/k+Y4aO7Tks2GWb3u5FTEXjB4otVWX80PYiPZtrgVBpuZQjpLy/bZey0jmow1I32vLUe33TQ
b9BRgY7WmodaykxbaZ5iegt8dZLCqEOezV1IF+153XVXHkw8VcouxJY5BuayzyfCjfTdHnIk72h2
3cNhPP0HaLYPD1Cq9hNTGU0VlvW6b5OBuTfT1uJJvBUdtblRaAFL/CL/DiUL54a5i4X8Y2nFmuWN
tGXx3ybiToIwvbckNtp+Lb24nGmJZMQpjjilfUMEugn+ryxaVUwsMkklsPz1Xu3eS58WwECIgkwn
xeJlS6xg1mT5O5APwqd+NvV+lkR/BklOKhhf8tGzZvNCU1WGB4XVpNKN7N8V2S1t8AKQ/NENsbfA
xBljuXe6hugzQOl0bM5nxyd/8KR1a/QUpDzVmu+FnjWvM5/VvQS/YKTPrw0tzmSKrU1IVwStMDIV
uOHB3O8nuG59jgLQFFBG2m5mxl1YKakWLhfgHmVaekRIPpafB/qgzkAzLngtKMvwaTJt/M1izo5V
8waMxH2X439Jx+Pw/nAdMntuGYF1yXlAHLtHLubEQQ4HVRw//U4ytYRB67PhqtDhGFYR/V2Vi2ep
sfO1nW7HnQw46yaMNTZdK1qltBUAjCfrohDJk4+HaqJRVX8LVIuebqMfPM/BOds8Zkl43ODnY5RM
yxW7ZNh2oMcScir2/Uz+w7jgwuPBB7QPXW9WCBxnZJYl98SlVd7KHcTDUrh93hOQf1uSsmk79nY3
ZS2ZnyvFmwg1YvRRCnYuALHtHdyUaN23FoZUomKFfaB7imVvORRXNoc02rm+QSaKTlm8YvFPW0Fm
kXagLwHj3XLSPoYFFWed2SZD6aKy3iwAphwZDSEAs6oJvFzqLick0u0EJpLF3GNtWAolNw19r9HL
RCDv+xKPI0e939x07ArMQFWasjCX2cehrm1XmgelP/QGSJk9nsdGCPZCVqsQoMOXaA/0lOfpgJpB
cu6+y8FgGkIBT+Eb00OSzMT6b3/HZSs80+0/D+Bqm+4pvSOxm991ssRSp/21HZJCK/e4bf0IfzNd
cI3HBGanuNK7fW9T7pSKtumh+Gi0OgHCXxyThzHXGXqQ1UE+iAHdtE35cyFkFU4Vc5GYwsiQ1EOL
U3ZyxBA8UXEyLcs3653aUnn5Y1Yr0ksdBqmhT4r6tWDKPeUE4UzYnZG5K3YY4I8duh9tU7zInwUl
gtSS5VG0dHQ3nJekxk4FpeT7yocYPcaIkfEjZ6CowfKq5xz8CINkwUsWOSK/ZAPmHK8XWYYlsC1X
cTr64mRAisI9w4TNslNv0OEcSnCIkVeQpCiTXWFriXvMdpBHJ68jPAezyCYHMOLWOslAA5TOmEgb
VV4M4hNDv0dILyfsUSMH+3kMb/i+qJCxnuP6lg1uNAe7dvBSR2RSjjXZAWAuuityl/cVNcjDCmBu
OC9c1IzkKp2eZEqu8GAiO2N3MDV4s/ibze3B5N+zS21RNbDoh1f4ih6rTArFgpdQuTHRSsprfQ5G
v+wbQXEjpJOLz18ew9oq/U5UWFb5vvvdtMUkF3T+vUb6TwllCpVrywDFOtBKVOCEC4HUQff9wFg9
Gf94denJjuhhY7Hj7MUusT9wp0BFPJsBhS2yspPtGJiU/2nwc5nE9brY1NAO+Ydvn2SFGGCysBIL
zZQwYfN3E+erRRsJaDRfP8mOnjkYUp3aGUT8pUyjMjBMTKm5Xu/N8ITnf7VhcdNGZe1gmJvCUrXp
Esf012fg8yI00ss9VDQus/etdvphjsjfgS28GPm8VOzotN4nzLjByc9WfANOIrzeZx4GkH0j8Mu4
5O0nwVow0fNyEVjWAXZ8zlzmcQbKl74aofPAnK4pxqSeiDKxB4eQnBHVbjuyl2eDbw6rgl4/4/8z
BnNAwQ3S08GnsI1W2BLXuALw+dDGTEN9yWL+RtxjQFENQDhyeOjgIDWlUUbzqe6kFq8UfcNSlvPC
k3PDXFwdX1lGAIXA90sfOUsujNHnLotrx7DdgSqeoh5yPqfLq6YuLFm+QIAsrNlWBAWjaHr18GUl
w5n2ker8mEKMVILx4Hy0Z0uG+eozo1OYsFZD+lWubHhxVs5yp5cTfebkA3ox1pmRxNPJ7uktKZyw
Pa2zyrKqVcqYrjIu8ad2YwNjuimaNKc8pZX3Fn8gWzoJE/j3qgX5KdKM9lI8CG0DzZnBNVgPysqC
A5iWc4hisI8W1FmLhepgeWMs43Q4CiG+Y+MXFnOkL5aMgwqOmPTpdhEnwNnpgGXtOmIBDhLGulGw
DCAHzz94ZIonHf1WEvGiDpN2r7fVM9u1yDo7SVz3qFj0pPAu3EKZ31IAoeUuzg6989PYVy6yqyZZ
iUdi3uWLbAzXR9Tw9KlYa0S6KU/zmZou6/1qLdwCYRz2LNUa7kwkfMNUSVN4iMPzUE+FBEYsLA+T
s/Yflc6OcJzvPv8krmfsIauyniu+r4OJmyJktQT6SH/fBbbki6eTpg9WTkM7ELyR9knmkiQirvL5
QjaTMOEkWfyJAuSRR8uvy79640qqTkh4jDNt/j+7FanNmTyCQ93DG9LPMCs9d04pstvYcf9lnYec
IG7fD6MdLbZ0vQzIA6M6kM0FTLp1EKp0VPTJ9eIgZ3hjak+/+hDt5UFLeeGw96HUEst7JZEU9SM3
BZgbwTKBBWYGksW1CzA8T/q3sHCHoLjFeJL23PcKW6CEYlVBltEptol6zEXFW5UpKMKPzX1xYvnh
lSt85WvfY6i9TqvbwdOaJO0djTg9KjKDRwvuwMP+9HaJLnmX9Dytg1NYLlR04etk36JPP2LdERU1
xHhn4vt2FwpFVsdyUxR87b7SvXGGimaH4bTYWpVWeMRQzy99TcMtGGioiVi1TreC++GTCpAH4FC8
3GVr5476qc3qSobWdQhHyHrCj1eTM32VG3KLaXzKPUSBSgwQKKVv20VSHKXJ1zq49yHB1IlMSwU6
SmtYaNpavQJTAHfWtSsLhn5tXwux02V+0xEEF+oDaZ0Xb4NzBdTx3H4EAZ4CASfZtONW41qd0B5J
7SKDHsKS0o5syJhctwndbG746Lm6VcWk7Lh/m+U1kuYYLcW3hTgfYg21uPp1y1c+cukRmk//oXVk
gB/G3t0mj2HPLN9ytst9ANQZfXbJsE54j/cvCLW50yt+T7dWpAK53VNgQKeh9fNFmowxVILUT6mm
z6+5rrKsDvpWPympOnuQ+bQrCgZhRImImjpXvgn/4D4WAiy5pPM8Fw7EzgwTdl+Ceif4CguDj6ui
W9GOF+Tx+YsVXA7g5iRC3ftG0l1W5nUYH0IbRULph6KCbndG+OFCPkdBozFYAySliwb6n3sKwXsx
T2IznJ24Si1CbKUUzIBF4npZr2gLZTebZztRfmmCK1rwNszieU96PPGZBzjKtBsv9fwOPpCARFKA
H6RzvYryTemOVXF/ngnD06ek9uYsSnSsBaV4e8bNUiFra4jMqQyq7zs85PTrbz/Pvp+B3QMgw4wW
elhm7FS9S2cO8jFFKaG7CgecOCTYxJp8eIKQ512h3RKdZLsCGf6aER68TVc21XWcYas/XgDBC8yp
9MUamOJJc+o1NMsk+3WzliZnS/MBcsXN8uz10/RoUvUIA8TYzYlNnjyrS7Oh/BZ/vZuGyhYq34+R
IqJonP6VCU0TIm/AbHEofmzwwf7WkaRRqFIr+AGzzWjsXjtL/J5omvX8TVpTk/T7iA7p0FZHZw+Y
QOvB4O+VACtHVNtco9XdMAz9UyfJTTBeS9NOeOnDBokL9NbYpqa+NRUUenpIXBzYaNF+DT4sohjH
em+qCACtwSQxkcXMRoTHEUyqp99RqwijXzjVgSKaQJTluch9GP4HNGM9TxWvK9SzcpaVXXni5UCm
XUWTgTuqt/jiUSOAf692SscTvm+b3KESsq9BFxSp1ySA4aaW97vQ4TWHKwMfUcPW7Db0MWoCPYRg
hib43q274UYmiNE5VQS+BcXLmWDS3uiSQDIifPxLGsw4NXI3Jmhmh46rtOGjAGnhX3bn2+zZZwyJ
qYSVt/jo8nYMrvF+l69MR+Ruddlpu3pfiEeLM49l6FhCpQgbNMeKUcj6zc3K4V9j0rWIZkzU9Zje
e9rFOgQAdrfnRZY/SjMrM73GIO88hFO05PaO+5bAEk3B5JTpSbYJh7sgXKx2qcUwS4leUDXgML55
c3jkVedyR6XKG4zE2Bhgsojdo76BQ05DX2tl2zC6cwufmw3ywFqVAs86rMuUc9WWdRmSQ5Vz6/ij
IkTJkntBb4ZoY+d5TjSpVW5ow6qLrvZUseDRyC0tQizR6aHtW268FLSoQeqqQ8vnYmgAMqXUlFKW
61bZ3JaeXWKTKCFRu2wTc13166AqUqvv82uOfLrRE8S/XLAJKLZLi2aGPhCeVQpBdfTgQAKKhage
aEceg+MwTSsE91Y/N9jSpkCSorqtzi8rjOslha5xfAKQRlM6O0gZ4fcbzGwA/O1Tx9DZHpKY9dFh
kExJDunis6arFRh/qL+ys2olcrh5Silxp9XhNNznVBiukDkaSnn2hp7SmaZAaD+liHrfr2TRr3qx
MPL6J3vC8lKkdB5xAxVb1fhSWQ/8AaDCpMrGUPP/Gi81cOcTUoLjiCRESd4y441g/ckmFFKwgLO1
uenAshH9/lvJChebmMcl+78UwPZQQFvtnIt/o2EQZQWyVZk/KMSpQDAn/hAk/S0j7t2IQIhZCLvk
jAqLWL9+jFaxrhEW87wOQv+s6dEWN8hHo1JJDhN2wTFA7S4dxX5lbyPyPCEuOSDJqRJCBdpsJBiO
8GHTXfnmbgU7bGuRJ8cfh8oeElkabL8NnHTgG2Q2CYoRmsRxBkPYuoHwi9MEeBIUZXmteke1hWPw
90ACNF3qKw4r8H6DMhv2hTHsZVkgeVw97kECiGTbClh3Z+PpPOwyykwBK3qq735k7H2Vj3DOObiT
FDY1j1oDmheocmRRYLdBjl97spa2XxDzu3v0zGvSVGAfifQf52PP1C4c+0GXlzwlWLb7smBn8As/
JEiItnFbAYcSaBFDx+mdNEa6Wr3hj71IgmmA2o0q+zQ9HqlF/Yra1BHlDMtpMiR6/oVjUoTpP2My
x51CA8EMxYJp9Ff0uSzlDv0VKuu8xrfH4lRojYTMlWxF44IjrI5S1f7IE19c0RBuAM/rQeJ3dH9W
zzIGwaSpXNbdQ4J05RDU5sbdpdw87b3tBZBOEpYT0nVWUaJErwo4YQmvLp+VjB7riFfiHDYLPTAv
6OhiuU962OHIlzJs2hJq2nhAd/ic0d2aZemRUmm6DDSAl34vRIukTs059uzwL3OijhYtKiNAADbc
JX6GcWFeE9J0HVsrVFzH2+CSnLv0lH+WqFgd1klzG6iLk9I32/fNHIqsR5PnBu+HmIRECvYNqiqt
YehHH+aa0Azl/KN/YrQ/w7xxp0xIL64TEqObOUi9ffeCxoJE6L6WAao7ooS9xWxUXvLoNotcSPT7
JfjBalxhCWNQV8mKI/6PMgN1mPxFhVDbkl8cfLSUGfDUmUEKqTcU3y2EWuza6NxQtqTJgll7jBrI
O9JT3+Yy3mfVOE98yOU7FSTkY5CiKzLhCNf1vIQEzOzavAQe5FtLxwmJxX995bAqpmyVydquQn3B
E4U913Y7RiPsh5JJpFihui0rvtjuCvqdA1ySQogeZ+VUVuwvhSNDhSckzv2R8Yu0CZMSF220xago
Uo6QtSkPv/4/HJVifIzOWGSoNuFer26XXblT4Gj3YE/OGlm+7qGcUgzBYWVDz1sqwh1fiCvOh+Mf
fG5fxnmpWPV2+pkFSFZmPuIr4GhhGHNIwRsUUNFYdufkZpU+a3nw/9Aqi6VYSnZXl+2YuYzv/6K9
c21mSecde0JPOApAVPj7X3M3QIBpu27+OujQ1i3LAI5hLOOB0Q+DL+KvdVZZbebeTqOYEnThDQmZ
9sjELfgNL16dshmKF0cxClqwthidttT5H8JeJ6D6JCRAIZRRoORBz4UYQcfiTAstGKmfFGXP7hh/
wc7sJlOzP5oR78sP6EQIZIythbCD540XRuyGXJ0hQOJUfu70CD164kp7l7r6L+GDrzhG1xM20IT5
1ayKgeAHlFSuEOyuL3CsmnOBtFEK6V10zcQilQHX0D4aqr15DRUZmy6YyVDmbbTKhLvmqmmxWimr
a78n+DN4Kr4ENhNKetRajq34XsLk+LnJ1+avxdaKnF5x3uSntYNzhxzAr3hRZpxJgzVtf4ysjoeW
wEeW1zSYIgbcWztnYde0ek7djxbLSyby3Xrnj9YVJmFURCPeZGbKl8NCKih0jU5akIJIV1eGWb7z
9YybFqf+/i0HRJ1yROZ74V0wiHLFfs705fUpki71KPnroJB+NPaQQ7g90GDENetlpwA2D6j5zTsC
oTqmsAs9pvOoEgkQqOXg2M/jnwU/GDe0/KZVn2eGUdUpfQAWgBspHj2V/48IcdojXuJFVpspfJTp
BMLijhfuv2A0DhReNNM53bIN20UmTq/yDlPAYGdHaPbrFhxOBfMWowTvcC3buBa576BUPGD2UQUe
LOg+iy4LCGFmTb3IgYX0kCKTigOA+WBI3JbD44C7dChr0QiDjvyev+jGdOPc8AA09BBmkW/KmmmV
6NYBkswhBoFBPDPGohsLKasU5pVQnpSpZczH0ejzpP8pEwuHRFVnocAmNJs8CuwycvjzuROzwA/z
1Yw37UJbLB1fcLNonfwZIEJyW8T2/XpuiiG3U22GmR8mX3XW2HDImq7at+ykglkPttlodCF1gpkE
hqCzMLNMpkNlYq7fX9hDLCoi1/P5esZ9qaylTxywmYYLAby9O0LFaOJ/vm0rKLeZx0hSUAElDeBL
cnQ2Jn/A1e/mir8hwjNZZBKR7zTSpgDHWz6X2ZucdDIkZEAdUdrsOYAZSIPz6sVkJKzuq92V5aQw
ukQBAfgmK3gnCStmiGocKNStqRCEiltNQpow2nawGdlJ7wsIiY5168cvRs+3ECnannPkqEGFQRcN
ePkH54FUJOTJ5DTiqwKa50ne8Qkz5jOKte/zxBy0aK19BJ9PBznbWE46PnmQtFcZR52KMukw4VbT
fExoPltTPAzWTe9g/HvpDrHLbRCj8OKi4qfOBllFhdQE6FLEVhu8sKHKuXVh0lX2ANYQyFerijXO
LWbeum2Bj0ie7lO1nn5RJzeXZcTRpQ5AlmUCOuhzruDh5hdYn0XRN7badnbDvC3gHnKOaFlJSikc
TWWli2qH06YDtu8rzP26/JJFjlbxXP7rC5FdchXPE+3USpqY9kd1MzUmOEomdcls3pDtEuwWA5HB
oHlkI8Ixm7hQkPaeE1BqCDJOtKY/zNauPsKD+F5vndlOPWnCtEXHDEr4f8yTZsrRwqSGjGL+YS+m
xisCqPiWOphHjvqdRCJm8a0Kg6Dlyu6cQQ05ZLDRc3E/sVavShq957T8sLbiUhlWCOapVRigyV8m
wEiuVheIrHFUkPH3B8Z9xyJ445m5DllnHbTGdk0vq+rPQkwtJMjFWQj2dVkzrYSlgphCfE6067fe
psLS2o8ggQbytrnyC9YFyw1u1bpMC41IFoKCzHPiNsjYYR6sB3+FntxIOJsCXiBuiHP/BKomb5A8
ro0CMdSMsrQFy6dWOXASlsKEqP6x0ILeMiKP5REell7CQKhS/OT9mtDhWnKfYOXlAlb6gpNtZcbU
QpNH/AGKw0EmJ74w89tMfb0Orh109zkoN8/9zCD05fT3KxtpFliMOixDXDbp6fp7q84qyzOhYNyg
0zMVYuEaUgxVuIt76o/lCBZc1BraAMK/18fsgJmBw0FkzyERfOvdRpJlsGFQyUmLL2ARoN3oN7Y/
NukWUjbnpG+m3OIM7fGxwBnKaXQG5bEioksnJ4BJm4bCTEmv3uG30pJROXuSx4l8yPuGNQH3Z1wj
dnOYBZ6oML9V3Qkc0Pr6e18c0lHHcEbeVV0ASsK1q/un1HXLuUjMXJT4sqGaRjt29XQJbn2We+b+
PgzOZRjGBd5wcXS4n+o+9DIPCJnU8uNJnbmaBFO9WIGiEATkmHKgpjtMkL2MMSMvnjaG5xj5kQSS
DiCsSqN9+p5mv/zQn0DrLkXzOjMYjDVltVyov0BudpMZdnnt8E8CkZjxDKlLaQ7FHJZWp0SvR15f
A+ZVD5p3xL5/NdYoUfmtuCNidYj0xWNAogCt2vz3UzIfpkWYctI0jpEx+OBvjr+8GyoAlYTtoHOL
DlGz1OE/WW8T26r8kx+JTlk9EQYf7suA59J4/PociS3gqDyR0ISOBl3V7H9EL3wymUSwMtUckz2K
3ZS+RBmKzd7plOToqRk8vKBEYry7T6o0aamawnr81H2uR2uCGGmccV4VKtriJiWF9U/hecwSKCX/
Ta0WqWc+lZwFp+mjQ1yJ71xq/17McuVI8r3LcqhDhQt35gXJal0CZa6bNr6QGTbRneezFwx02bPW
CP0snlXGpls8uYyzoXmHdEhm+EjhPgQU6JEKsCZu+QEXa8HbrYU+GZCDnKE6wVedw8MV9r6NLHt1
ip7+cJZQgOcppJcbx9wo5dNfLRU/92I+peCrkVKVn68uDOqsLf2zjqh8aeMrbFnA2hNxBlMnyELJ
JTWTDOnHPJ2Q2h87d9WqDmY8qneD5cy9OKNcuD005ZGHhcaRtmdEdBqAyARX7DuuhauT4o7zGxyl
h3wGVVc2se6zj0s8bTLRAT7MxBtHbaUPeaZ9n7QkqAGhnRGCgG3Mlea3eUHBF64E1/rGbkimgTVX
YT/zE+ZdhjroseCPX2t7wvHNBfLAe0r3+plI8zU5uRFfwpebypHKqMZ1pdkY+zS+xzpuiRCM625Q
3/WWIGTaT9ivZth+6EPt7eTIkJVCnA3psenw2IIbl2iD7ZiqUm4o0G3Ssxm9parvLmCowbx24zpl
oTHG/1M5LZkz47cGi0TPQHau9BN3yKbIR4gPDziKuJOLyyCUed+j/LfZNhHBUOmGpICLD1x9h9BB
zW+c7HRDeR+gQiliTE4M2ljw9Jyz2D8mKpkzhwyHVlNxWE0tFYQQNQgchU5wbXhyzwtlWMuXRiIW
xyvJjgzQ9Af1cOPIyF7QSGMforc8GAFqGs8a7yHTg/1P3wZO5LoGfZPeS5vUU1jB6c4T18STSUR1
NhuLtXzNcvyckA4/kFl4GQrm5p+uYZuTZbq94JPD/BCpaujKIXira+OKa/sKelr+gsA+11EUpzzx
ToxlRl8OY8ucwKa0/B9RhloKPzhJdG6cfTcx5kGE3tsER2vzkMa60I3QPxiZRg0ou1yXlLbexMC1
FWyUofh7ViX6aUrA+l6prm0hh9YzNMrHMWCQ1mfl0zQ1kZntjqaJC6ww3PcANCQvig/d7KH8EjDo
LZ8g914J6KUDxWpsFKNdgNA8HLeuZJFgtPCCaFOLmGba24Kl4TRQS+3vUvzdkHmHWLx358lJ+io3
GXeHsm9IFfF21QpXuneNQms419xCIIykzmWK2sTnRTBT2aV6Qio0Fn0yN286wJX24O3cNvfuJITr
XzqEf68jtBCOzBGEmEwKYFG/c80YNA8tjF1rcMVyEQ7YOSk8wwuqU9RDEQV8G3cFR0tbXgxeYVI6
i27w98ENXZ7kgt1Lgp5rzMOXoeYy/85B91nS03+hk9mPXypTbRK+80qTjcol75jn5amZpcWksYp0
HyWkdRDKnPbYlkcdAmxgwjcU5/s+zhBXCSAkAmhYnTWR/bRtfs8lAZUvWSz8xLUqgG45wxuyzHV3
Zn9+gBgX7fVbMJpo/5laxMyDXVdtIVc2v9BaYYfA6LxHypLkYs5VzRRfoccjREBa+l8XptOQRDQ4
mzl7U6VJV2GQ2Hz4J+p76KuAtcE5iicKTTbhVUmkzoBxhWCT9yVqMUVzpujApci94ffTQR2pXQUn
I7a1UnY9x9ETIAJM3tZDSt6OvPQWDyPs15XXQ/eo5Y6KWt+I8zlWLkr/3jVgMlYWS5xmkknUoG9W
YHe+i90Er84ye4TH5Ey+eV2yzerdRPPfq9VrSgW2gQrkxZ9nHaQe+PlErBYHxM7pfwKBuqxcpA6y
z5VQCdc4VBLaVZUiczuUanhxPBxeOxUnYUfjPvkC2iAAT7BNFBbzPv5mdpk8DPAdw4qXnGtTwz7S
b+uH3Pw7fuiNxCLwtypsg5daqjY640NglG3ubeF5+6KwX15S5shUSJaQ7PWOoFZgq29olM4nTDO2
zMG+tam60f88BhxBzc9f3fj8NRECDMog9R2kIJu/Tc1V7eWkcoMVF2TZ2A9RPmkoP+LAPp469hkb
JuBzyMeXrwLBJhPOo/xGt/5/GXqzKahJlYa35Vlk4r3V6Dr5Dg8hOme8mYRsBjQpXW/F7CBzzhiF
TG+8I59UIp6AB6+eslmZtZyFmU61EqRLIthMgyNZ7eRmliNWwQpcjKRPUTQlmsC3CiclhxmcEaYi
jfaw1l70pelV757Tb2qRPopVvAGhwJcZ5lH34E7VvqR6Gyqt1eRhat5GmccazlTbIjjSlgWEBpr1
aY+9QP4u6jDTG9s1DdXsfM0e3geSNdfEEpE9fUVuS4bCMX3IREkwt0IrY1hr0jWdJTsrGBxa/m68
LUEbyRgWd2bRRZ/gDUFucLNY4lzsjVWS0Olbh4hevh+xGnGTCVytbEX7KJK3oasCKk8YwUhODVN0
ZOBgYk7bFhsZnn/+hxugiQJR4xg0U05jexTtZeVyVBB+EdLsyLF0hvPfHKq3tkQ2vMuGNQjrZm1A
Ot/tcyVmk1iHf0Bwb3Qzf/PEvLvAQmAE42zbiTDCjPktiNQgXchNk6ul8Uf/auCSzq8MWfP5vrj+
nKThq9WhMGVu2vVetHaroE+Oq1GRIxnPn54r94zkgzmWnL9lJFFoycmax+K5LAGsSpj6PKpsngfB
XBCgH6cQd/h9AhTqgNygUVArwNEMD9ibL2HqCeuvMDz9QxrTU6/I0FDwuUyqwEULFy8gRBq8h0n0
E/u8jTlITohwpRX24FPaxuysaFMjBPiPDU6x6P9byljFJ1vCEUJWJEv1B0v9xo8IoIbKQoW2tjkN
XZ65A9a1EuAehnqsNaWFSbvDZRReJwGV5bjPdE1is9ff6aUtgatuslU9VXZoXmODWCaSuUItLZko
cPeNApdtlF3lPeQ5K1DtECUQwgUVE2svJeXiUiaV0EGjFQtW1qi4Fp6+kCLoSvh7rKDkHb6bojQ3
raTJv/vUaW9mreAGQzri1vfcdMvG749neplPpfg8N0PBRurtIgwSNEp5N/CuJssq9FqceLzcfEzI
4PxUYAn4JWgsUgEhpInJWCiIaFGFyUFEZqp5ghA3/nmObLpMMUlev/Utcqeh9xF36sxrHB9SBoEq
czlxED91YWkOiWnq2OjCHUo4zKLMOK9MzHCHDyD+X3uvyAbsjE0ZHKI8txZ3EnCcNdUmTY9VPOSx
fkhQUHC0AX2QzCIziVuNZ9bgy3An2iBOANdpk6f/hRr6a0uhkXhlXp3uVTdQEzRZqEd1SaFLDeiD
GMGPufI3e7pMUuTj7+9kV+6472pYg7xEq1/dw8jlZfpGv44QoPvZCsPNHeOWCtdSP/dgqoEpfFXd
n0NayCD+VJSxNiMnN8/K08GTiirnU9NNi1AI1AaOK64+7+zDh6B9JpptAOUoF4/cLot0ahItGETb
nBm2P5OsaccKq1fLvIsPrzEZK/5xPTnc1AX0Ze2vRoOvDtSf/zjHPr78WMRSORfWfw3nUJKY88dc
qRuRSZHu8cth0Hq8VOwVMD6xAsCHLChY2OTx+1tX3dAzHh+byRIwqe/JzGLa7wqbLk9002Zjzbor
DhnrbASJqI8m1o23uR/M+h+1E9+xSRBNSOdX6LuEA0CrsNlHswahpa6QbAkWRoa3NUOQOHh3PmWu
W1AtfXZEy91SQLNz/4RXwFSS+8UAThBhOVwW/iigD1RXMcLROc6ubRZdvoGjLpQovMfGK269L+b/
dT8YjE19SsNd9umSWUSlCV8AgTQnzujXTQe0k8WpYhhsuKKygx7yRoSFCh/n4v2P9f5tgaZZmHZt
Cx6gZRwtCrbTBXkIHuMwD5M2hPWmgAH2i3GYy3b2ZWtY0UW7NMEtnJmSxbbhdah5D7U3ruorThWm
hMBCRDVSMIwh7TYyb6Yebmqj1yRyfPjbj86pP60a+gRVuz9LU5jSx22d1fkiPNP3zyYufOTA6rsL
gFWrc7BcPha5ne81jFZbMYTx+GOAPrssAVzG9pTBN+AW9S3Fyjv6pj6kLutETyEsLJFqZcvgv9Ml
X2E/LFmaTmP7pXsRyIMimC9J2ANMr5ZMcW6YwgKGK25kD8i94cJcptgRGmtQe4nEVxESGwJ1nLp9
iPDVwHa/TM9ZGlX7Rg5QP3fWIXN5vUXfsuIONudOrTACUaCVP1RDndrjNtD3IHP1JGZkpfEDMP1i
DrLoHSgGrVHGYdCOWe+AUKsggU9I2I+DaHB4z+xmgJh0czVbW1atJFcHG496PyLScTdTMOMNOqfe
eEOrkF9AXduC6gHuDp84Jl6hGMLpjnffMm8C4t33L/QU98TKUihxvjXrX8uB/oiKtGcTZT34uy5m
56ed/hRMZJWg2rmnj478nCfRWJue1PaHM/iQHMA7/4jkA4xSBvr6iJzFNH5z6KpyFUCC8qxqFqp1
XIyA/E6Yk83V8ysBQFXoyVHY6Edvo7mg6ALociejmqBBPlhA7b4LwA11R7B1OsNudAsBSykhtZ2r
k4ONHEiqdE1aLdrwAgGZdmbWIpo4zYqGPWzW65wXXiCPml5zNDyklTmZH8B/U2BkjScpXx3dbZp4
dyykIjhHI4SWit1x4hkEU4Hptrqu0pehIvSA+RiAcUHIyAvRf5LjiCHeRbxMqNs0rJW2Ib+fJSAF
v83u4c1cqkpQJkwYteP5X0QaalcO81QYDQcWWIHDYVPN0BNeOfdfRNAenl1DrWwSWEYk4if2pvkd
aL0IvQTq91b1b//4bnYzLll0lVy6Ue9y+7V+CUs9QdFfKZsTJQrxSvOGJHhD01AKFiXMvsx8UV6O
aVug6u/Sf3GGy4XydLJZsPU9scQ4ibmcEdFl7ZbRtC/34+kBA/VyGHhaySeX2lqyF83ZGv/1/lW5
egsiieKN8RTe8Pz/kBAQY8gc6ZnLgZB1qwJFR7oOdyKEEkBLzUwmHLpHC6xMXzJKOicI5jl6wkV+
HX9W+rCj3VMLKIoV4llu1B2+SpwAC85arThDFN0FDMOx3MKKn30jc0B+glHpMSmudn5aXkE/0qOm
FGC3XIeLqpu7/AtSxPa8HxlYejNQW6X19RXo0UAEIi7H16J1O1CWVK5GfVrK9aG29WsSLa9JpRf4
M0Qoo4pFIZWfy0fB0n5Q1C3Lb6sH4EC2EGMQkYnBCT2Xjf4FocQYC+ucoyNMhH8gWoJ+rrtUOsq2
5KMUi0M+8rCEr81FBOO3+Nj8GVjtl/SdRQJJVc+NrNd9W+PlbiAn9Asj3oljejc9WH4QBye9jg0C
SFr70m4jtYXXuhk/66i+EZNYhDG0X/DQQMu2BAnwnfDgLAK0OEglyLoR7Rt3sH2kYKq7/J/lUOqJ
aX5NMCVxgYbDLP3SX8KKq3E4EhA8LmFaSycSYnMzXzVdOZXaJg6/mYMSGUyh7fr1kGMVG9+crRWw
WtmXtvGiup385Welpl1oVYpGU0diTvg32PiaY3XDZ1f/Ft8NIX5X3BORfAJnxaQnUwtf8f5dCUzH
VhCGZtvVCGUqB9dskHd0i+5NqYDZVPs3dufljVnSqUUcPjtQdteN1x18eq+//TWjfzjuXHrAAVm6
uJdSXhzvOyF0KDYDkosbhLk4aaKq77PNITN9bFjHM8+RmdYIYLJgrJaWsf/Pm1W3XqXpb8ZF2n7x
LjZFqURoW3/rMW7WQdfhgul/lbFhNwBAdn0NSmuw+UOQj5NLg4vxlnYzx2yuaJ+ugwkhiDa0sOtr
eicw4QAolMXBegSo45o3/5dgoEIz52/dtNNAitcAxbuBTtf/ihKuefk//niY0HQ7klBecWa1AMtS
8wnyM03P5L6uVzQLiaiml6AJRg6q4OvYAMnPgusPyPl1QaW+a7tMPYnDQtcX12fT/yFgMc6Mtz7L
vLSZq/QQUht85zmGU/TCftOlbwZA7/FOfVO/gGMF71Rkf2buUZ0ea2QVKCw1+kdRLpadaLt2IKC+
5i7dtfObu7S1/hk6oKgDT8Je6SobBNkqw8GtqUUWcoDxMesu7ocWThos3f10G1lmP+5tC1XKB859
5VilCedeACyDn2hIXg+Zk/7kpBpjxScBllMSyoslwIdwOiP4C3I5jegtKwgfSoNr9TP/OOnc610e
kRU33wVQi3Te0hB5SoLoeeNv+wINHZ/KaYjjJmLShYGg0GRnB0FDUH6vHzs+PClfxMbzr0vibcmo
/LTa0gZ+kAKpX/0AL6rMe7dOoAHx47gkuu3YXKy03JK+gEQV8JYkEx3ig90UXmiVFCDTbvS2+1rA
9Y09wktsEM2Sm2D9VpGqI3eYYTVpc4xzgEKVEJIR8sKllUUC55R5nAeL4P68PELbgzgb6pIFlklB
Gqg4qeZWlBM/6DVSL3/4tffOp0lhd04zRSUQN+0tOkV8juG7RdCvuxSOKg7Q/7DHTsDohHHw1ZyS
u2HNh3XHAA+wcNPgK1LImOitFXfU6tqfQKxaK6LL7q37b4oVyb/wsotgU/3j/TX6MzBIK0pEQXBe
KTTxfWUrVg09JAAcgi9tPiIBdoMa0G2Nuj45pWuC8Da1Ao8Vent4IosOIykqmMJIEbz2K152kYmT
j6Mdc3vOSw7zFkzJe1N5/OAZyWjb1NEJ8TySXQ5oxnbsj6+m6mcDcZVnfQTqpaQ5VyZLNTOAOmBo
/DWEbG9zg5irmTb/E81VPZTsPKIbAbsKWvMRlG8r3kFqU0ppq+2lhbjpxqPIuuSPuWPVSqPqShnS
sCjo+tdDBovVSWwZgGTMzbIwX3Mexlw5pQeYqGgaYEeanFtz7Rbvi7QgenJizWhdpucYsBG9qBc5
Vg4anpbKf8PEB6cqnlyIRhG+GMwCO011+UDeLKIrMfI2rqbNYXMXjibdHsl5U0z7mzzUNKtx6oH1
sv1ldWL2CAUEdV+e4j9yFwixcMNHFJ7zh3qxL/xOZ1ddpZcdOrI6OCdDfAQ6wgNZ0fHLuu2DdtUV
RinlY3lM8l7ysbLxY2wz15FMKXdr8+6o2a6LC/KimG0Lkn+SovHK3UOBsYe3g376ES2yU5Rh5OCb
Ov3WaYIJ+U5FKQD0b9MfcdxAenY2evYwtY6oM3p+XostPm/ei5DFdeNDmHDibh5qNvKY7jwiPsnS
BDQVoFpKrTTWK67MuwIcD+Af2XrOEGnJeoppIz221FIyCZdtq22qAvWDdB8UinTjJW5eiHspcJIK
CMzheooZO68PxWlz+DhazngB95MdBQ+na4OvbR5+9g87aQl1MPH9xluFl4wcsITkEfbqj05zgIQw
1WwtVi6kVOXWnh/2JQFuvZzyiG3uI5BIGZGAYMulabiBid87vO1ZlwY58nFfmQuAK/iSuaW5oAv0
Kr3++a/2Q88xatCy/iAQ8dsYPPwNyOeDpSKG9/eiAoYnWUh31Pa1T0ioECM2kUBZOonxNYSQSk3q
A7fwmH3CBRzrxBJ4a6nL5q9Wp434XdN9DIm/fEc8DchkJY798XVk+BNb0o3sf/41nnsSKwY6+knt
pHEV73KBXPwX6ai/Fo4lqZ++XbFtKfmP+/J8mA6gKmJF9cGnlpgfSZwKWGh0FFc70aQ9CEiZIaTn
BNoZRSLBNIRX3RY129Qy5ca0f+dedUBnDD2dAbYV8hThsXay7RfHGas1+lIpizcR3NCDqCjHfqyZ
XAUiwJGSX02LyDxt7bNhvKu0tQJRsI9C5VpiPmgEnFYr8iXnPy7T+uJfNgoqYw5RzpkNFrTgGAFY
tThW7txiuOKwwfrecifn7kBTodMG9EBgzohe3dICbzZ5e3UsufKYfBqq+EDEVQBSj1lE9YGKEo/q
PN1kTRIl0eJR1jXcRnf+2WwgaJ5IO4hyCNdKv9cwyfWc4dubt4c7kxxfPuzo0bJrDrvGUJIQjH+N
eOZymRO3CF/a9DAWiunmGVeZNRWq+D27gmgi8GGttrd4NZk5d+al1/WvqxEMWKv9ghU2smd6GvMM
R/OQ38tfiJrvCmWjph6t8hF56rFRsBMbFNFb0bKoxgyE6tQmBVIipQme9BcW2M/DO1z4xXVg7HOD
g4u9LF1x/lBRQ4vPjVaJTBO5e3J8v6KlcgIoUSTqijUkDggl5gdyPMiVZxxVUCCLLhhWpVsJ6fGg
qSxUkc74Hq7+5bboH21SzUvfXW40XDvlWwDAnFXAWQ/wEiIo/s2NhVBqCZRW9voGpt+M61AC3TvZ
pe0gv3zfs/LG9yExm5yAH7RyXJjkoeLMjPkn2a3tnEcMiwkIuPK7BRi9FE0AoPvMeuFMiT0zrSDw
8ieHw3b7vijOXeV27Lgdv6n2xGDR6/MoS+skLDijK1M7qkdhP+LxU6yF9OR1mAO2F3AXa1L2vZpC
de3jEFZoCEKo9ZWfvPg9JIFitxYoIjpY6Z4hC4ZoWYDlajfAvsfXnfV5zwUr+7FO3ZkTHeiba/2M
YAXbnnJbYsW1zJtPMZWPb4DFWuXKlZ2WPcLXj2Yo8LsCNXqlROA92o0gPDA5zPcKukEw+UfSgxDZ
FjqJZ3VonclEMZ10vTgDaIf+WqrePZhEuVnpib0V603qLwElCe/SFwqbMKUHCjiwLhIYhTv+uDH7
GmD31X3xaWyYPeWDxZE2rBPSQV+6u3pScYmLQNakFltmrRfaM4xZnN35rfT16vx079j5rZzH1VQX
odXfAjUbYvzwGeCo2jYxp4PbUrVNyIVZ1fp/Yvi7ieFIFTX9us6efODY8rBDZpzddt8IJrG9BIwC
yJRAi/Ir+zLdp0Z2OOg4p/21np7KnIN5o8FDitOj38bpg+sVRNK2gpU9BQmFtD+XI+JgvCt5k4gQ
uB4Q58aleyqqR3d+QVPrNCu7HZuWlgVVcBxl+88hBcIowNNO3su9FMw+1VtsgY3RfcDPwd/WKEaS
tVszzc8+TAvCXBp0A7w9buO2DCkjroWmthaB9yrgPWO0htx8Zv2TinWIVMBDOPX4GvtcMwsS0Sah
qe2r4fLDr+pfZlnoSNiZi1p7TDunPqO0/JTNJgAT8IYDU+AJWL6i/B7b163pjSDONLbWX5u6nEzr
BkDdmtUnO2RV6Od1eSgvR/B3N9xBfwlleDjeTd69BMXhtVjv1CZQbz1UsV4BzGgtasALuP3OtufZ
iQhC25bq1SF0QslRtI5g+B1Dc166ALcO+t8w1xW9M0DcxhyCku1ACXgCbVUBUGC39PuO0NZLIxyu
60xG4XvVaDkZ0NhGYoBsMhaqhfEYChXt33I5Qs3LbmsacZrs+iiekLsDqVTe873Ch/Jd7pIOWaRs
66/NE0LC2j+zase2mMA6qIyoNd0IV15+HYMC68wcLFaIRWaTmYvhghw4w0wqT1Mxk196cUCfqdvJ
EzqMRUHKp8na3T8J3+fR7/L20peHmtoKr/gAOuxUaS6n+mD+uu21lkIihv2mlzckD4wpwnPEtQLh
qt9ozTad3BBDdMaqrZIpdwkccCKwUmSolsv+lTFi0K1Ychcq6lIidBILdbleczVBDCeh0WlYz+uo
Z5MlnCpJ6dttXbOQpmfP/VzeXfNWsfOvw9VMNV5FJTGniqf9bt37W6xI9L/GqB49nqn89zd/dwR5
djmsEHkjW+eB5941hT29VP/nKQ1wsKT8NMcgzvJs01sdpi5iVJiX85Dz8HhmOA7Gu2UD7VR8RhPR
YE0gv2pghJ3Izl9PQg9qFnYtCrkaFMbHYY8SKwrEdBxazXBJ7yFQavF90as865cYVJVIwzBtLyI/
NMsRYsYSE9V/fIkbpVE+ZEHqxP6JTEYWtH3VGEFanojiK+sHWdoOt3hv0ymeGM8GZt79sqIgFZhX
fSEYafhoon0uAWGNCruFXekTlXWeEFQgor6eiyMebfTwsr3//Xd7YNO/gcRvPzyHQvgNsq9H6zEJ
xYO+NDR9UMPxEroMpdjmZ/laP5/we4PEeVOrnMejE3YvcpKG6Zpdcywm5itjCBKglJoRDRgKtQ0t
QJwfRftAeBhR7agz5XOR36uJVyLc11/em0FeXbOhp7xE/Kv/Ay5y2YSqNApsoNJ+u1HK9VC7yvtD
w0mkKhCBtG5GcdGwPN9rA5ZIQUa4BbcSV1leHGmdBngpaqCpLaVg2o4PZluHR97NRkno4u8mHMQP
wRc3+jOeboL1AipZEqs3lrNv2rT74F+/FzN6xLvwI4BkkGFLghyYYVUKcBPaPkMLW7phK2+14LgX
x5epNF2Z2g74Yj3ni7dujiJ14VX3SKP4V8M0QdkLfVCgvMXkLFwbMF9v5fQM4k7hcEKIBWLHJ6Nv
y2AUvWklki6dXhg8eI8m1DBN1Lq8gbrVk2X/UU7MH89PGwULfnrWh3qUA8rrS4okhL5m3M1jEfBv
N3lcAILnPwd9iIB9xOquf+PSv78YeTr3zZUKtKKzdU9phckJ8q1iqgk+xiMFiQxjv70jXZMc2RHm
jZ66fJzQku4FgncHp5ZnzX4WY5eF5pJjN1VszrL9R3wT853lYCEKj7nyGSjYJEgqztQeY70HCUbt
WAcS+br1VUi/ke+pSgBjGwPmY/854Odimn2M4ASpiE0YAGyeiUUSvYLP6sdJdUdHSYtY33117BxG
GDpnLgDmiaskGKS0iM9B9LOUl0WkY9CsBjYUq0uHdUadPvk6X+ard+rijjmkPzgRV8eAEsjOQapO
Y7AKTFTTTioopd9BvpSt4HAvLIvB83Mi4odUCv/AOTGY3M2nYz3H44BtHOMANTCdJzTEn+6EVacd
eNI2vb7Nmsnch0wn99KSiDjsriwCXCn+3km4uMZsb8QgU9p5/2BiJiMnwxvLR3jrAyjGugIz5t5U
5U6mR1GaK5t2LM6owe6Kqu05M60qzT5veVBDOJvepWtVs0hiRsnMKByHEN5EIS71IxieDw5kTxA4
MZZAFRAduSx0x5Wy66aYO4IvwXldlMEMzscDHPBuhukt58EcerN8GMOgE8+oud6olBd3HkX48f0f
KgAT1sOnm1iBMrOy5BZCHK2AAdEGFagcvfuOw4g6luNyeTjdS2DAj5dNFn+LYKZk/WO2nyvOCRsJ
XLInrjXtpDNmJ2PwfcT3oxfxcXT67NocuQ60SsX0xhkgUviQ6aLM4d/Nzgy2VrwQ78T2oxPh3WyI
xyF388CBWb1/7CAtUhR2KP5Y17w6XBY9D0OOT169ypYW9M97IjZwGzTNiRmTbLUrV396dctQeHY3
QHEnExqhL1gTMpDCSmRjyY6NnS3hljafYAxom4b2nNnm2328difZ4Rr+1jzys0Hy+RM8drO7hHoq
Ujrzb7FhddtPTSyaKk1YSLcgne72M29P0Q8Rn6JNUo3CgVoCkzQR4OOb3b+bYCG/N4nJrqzCZm/f
d6z4Ea1bbIA0LhKZzj1e8UDEYItewayXLM8aGG/wCjJ9LtUsJzh2c0WkXyF8eESlT1rQ0RadyMxZ
+bkWWWbkZgqnobg/sY3M/dx0qndc/vdWcK6pDe9YPyfGpn16tIitc7n1GukWmlzq09+MODrk1iUS
+TenKeKRYlxm6MMGit7T4/Mir7AeAsfN1BOg/wyFLQpDfe5Y8kTG9UCxqwnV3NlD9kGQ4WaxXTo+
8mA2EW9/Km73Y+w/WRdJFZxsfClVUOOWHER1nGJPC20hnxfS5Z5fZs287DijYT+VuLnW25m9dbIj
Ei0Iff1WWhw/UTeFGNFG01kqqjHkbzZAdSA8c8q7esq5pjLcKPH+xuJoC168awT/UIBdzNX9jdsw
d0FHiOCIhQgJUW9AwkqJlRi4uHOHHzwkIwDh1VB9UL1kMVmaeFcrCsoYTm8iRF+pWK2Oxg/F7UX9
H+nkH5JgtYkUjpvqn9kUCFm7yZ4J+dM1MedtGCwGHlob4JrnGhRbxqngzQg8jAXivTJBfSkz/+Uo
ZscNPiRN6+ESa29fsDGfyAvBxKQ9Fk7YG09Wh1eRQdx5gLrmxZUKxeH6kG8uEBCvKsx9Je5Tpi7Q
fe8BofQTB3ayuGJiFI36N6af4zQKT2p4gawSj6FakEUhnBr+98T2qay5ZK5nE5635uXHQN57quJU
RARey7DTJz6q3lMZJ5kTIwnfVi4lXfswUVUiBb7CeTjXnFknrrvZ39IJwIvLeaw+dNSM545QhOnW
1T0BwqWyddvFTsrDAXdkqb4Bozhfeq7bOm8kENF84y4ROvFmiAmQ+9VWdCvzmIb72s1f+e6e6uqn
1ows94UrgLnj7TAxO6jKLz+t2FPdYyDuA3QbfGh+MHB6kpp2AjAp4acmNpMKYqK+Jf7If5yYAIfx
58vxhDmpkZ57e1OsIQTxYTu26ZEqDnm0ADj3XFxpXSR9mN61MlhN4V9EFYiZGH+2sUcv/DAZly+y
no2b8heFD7PmJWAxotYv+6J6ix5FsDPfXnLZ2vPfqVyxBk2lPtOHRRMfriMQcb1U2AC6YRBsOAzP
2jcD9kYr/h/klNNb9xapXv9XcU1tb7Xs/KR6oSE508iTc+ov2BZ6hi4M/OdLqpUO6z9ghmvlqDQl
enEEj5yWZuJig0DV9eZRzWUkiwCtSnWx5wg0KCcqozwpCXPXXsrAwS2onkNQBJdleRvQ7HUABX59
xTGyoJlGHsEXel3a2x1H99aIoGZ8ymDkP+Hza6YbGG4dK2Q1NiEm95Cs8C2C0glenrgSSAepRGGB
rsGU5cineC0miM5+ECetTee2n4uJh8RH5gnB+0D6ug3zpDXUrtX2YvalX5FnBkw13bkyayO0/3Fu
rD1X95XrBwY4QIyF4FO9EZvl6Tjc+C0wq33J78pVduly++eXyc8Z7dIQdQYuIGP7etjg0PgrZ3GT
N8RWOgmWTdHserofZ8HSc/55x5v+NQ+2SQgJsQATXroCxMJavW+od74lbdTzOTZCqzFL6yKYEQED
4OjOZieSZ6SNk9mXiAXzJ6gZyIIGYbD0cejt4vmLylcIhMZN0cut4CL2zvFwfkFBg9nKjqe7tjNc
Oh7DB9UVxQPZfnLiPcSB3FoMy083o9hjBiqtKro1EwlV1VP83D59Oq/KNZuSCRTuD6x6DbuTMJQQ
Q2HEvyFZCYWSUWK46Y5j1w47ZOUnSbVP25HTd8tuAhiJKYFlNbLrKHw9aPOFEQsBy4Q4N6DSNKXn
HoVCwLyW1YEMKri+Lgr7oHp5t8C8kuN04uY82dMop9xAUijT4LQAMlrXpw8v0LUePB93DaSomARK
grOHWzbt9P0RXJGhqP8OA0gdHoLhHA2tIl4y/csqxBwRa5G2+TkGmQusgzKwtUeEeUkyNkgS0vL3
+iz6BXCLsgm0ptLgVuuHgEo7AczuvNgcHzyiIZ1pcEuyOqHAfY2qo8yNhrqRz+g54lCxNg2YJmWA
iLj1sX0gNTuXoE4rycK50q4OCK7N4IbG5sp7vvj+TnfREdLARX68oePIb9KZwsD/BSnqIir5Oomp
yYySR5WjvcRllrrHKvrwvYyLcqimlpxbmlfSKpKddoack4G6dMOg11zpSLlq5wKSiLvPdMcA8Aix
b3zI5lstZywLwlhro+k7IxvzB4JRj0vztLKPSMjlQJOaJAGXvoN5by8sJIB3jCP/Hq1nHc+A1YCw
VJ4z3e3r5qVcZzV5yeblRB4pR0vxOzJTrk1//Ra0qQ/GfxzQKesmsvpkoF9/LPuhlusI+sezr23I
6Z50rx9gdQY5KwFdGhhi3XnhQz5Uw1/oVy/QC8gPP4WkOPHpEAZdWvISB5LTahE2swKt/AGgKfQc
yfPwP8FF3Sn+rL1SLSjkwqyc5uy/zuzKgfQlFTSO3n3leYDTeg/0Tnw4tcpSpeuKaoE6c6Orlhpy
quUsEgwcWuGWfRYvc/doEQVGmzgMdhcnSaX3731WYCv7Uam1ZkTOv/nBbVlXMu1BUtzqI87IVwaA
DKNYsJIW8QukJ0Wf0u3Z/iGrusIwCVQE07dsskJOThD5AoPs41FScP3ddh08oer8veNaFz66VH34
+TmxIGtPeSkPMWVRRK8iyzsDTmX0toWLxzH7RMXktsPXSJwEZyf1up6uqVBJiiAzlcpw/B05j8mn
t5B24nYSkbhN+dVZn1AvTvyu/8oV/kKwVqaZJq5sPvYFQEDRvMKKCiACF8PGtVMVtoYZOIpWOtU0
MbnqeKPP/zuj5HdVCpleah9YIMDR56Zs4J1LWVug/4Au65r1vzBkH2hw1XktYkj8MOJnGKF1vnMJ
8ezNP8gQ5VatNbJDbXImLarr7OKfVK6fmiX3ycWWW02WjBt7nkFGfoxn+3qWDtsbLLiEzGm9/Gyh
ZwyKJAqKKAVd1osvELFAz/K/lYXv5i4BtF8XlNpcZWCDyXvKJG39M5bwIowHGN8u0o0e6V98/CKE
Y4mAAhcmq3F5ax58+ZvKkIzzGNkZ+Ccv2gHVU8CHtxna9kwUbFSxGE9q0eacKR/BmG7o3v3vCHqy
avo9aqiRa1TwCsA7aByVFN1uZuaZdqQFEME0tfV+eM21RfCbGZpiEs7H7fsXOEzEBZ3yX45WNniK
1uhwbud7F3HjlS1godGkJ9MKTB1TtAr4hMPgnyIU1Ntko+d2ZYrTjfpRmR2CytC4vZN7BlldMLzV
rLIHmhAzl+RJbWTqqjsUVhITBXFNCBZRD0F+TaeHzCarIwELYNIKX9rYI25VKzkd4HuBsKcM6FAs
Ocr1BnQsVSJ21+blHGKnsB0BCD/x/Eh3uATezFpwyvM3Cu99TswxLYImWWv4Z3vbiiInelqRl7ZY
uRkVtLoP2fEtL1kaoMGMNCwQ7iQv+J9Eo2psfEYMlxKQQQKO+WZLJHH+eIuqVzNep8QjAWgwM0gY
Q/9+GKm/+LOwz4zT75bToWvZ3NV8rl6Vd2c02pv0liARLKFmDBYIG4m1E+VDlbgFxompIW0I/ZCM
6f98oO4Hi/pBOknPmu8kdG6MxqyvuX9M3M4m09L8LzLflR/0VzEatqPadrIyfiM+qNrxsJZ9/A6Q
yfS61OWR0vDeLIwsNJl/xg7e+wRmuqpE0pblInqS55/2YvJ1WJCOjvuYvcizMbKNHo4fbcA7520w
07gB/fDpnKNsnAoXlcrHLj3dCywv7D1TYMDxnJ1uUHKPfPpgyBsj9v0harCbzrkbDhuHJskN3og7
dOdvKPrwG6o2wfdnDr0MpTTW82ctCjEMMW5sBjsoC4Zk8KvOiodwN8uK12nt5T4clySwo9F+hUCr
rGvbAer9rZ/R2A9TjQagIkjLlYouKE+uka2/bEj8OqWATwogfLv28Wo4BXgYEeRaYi6jm2ZbAStv
UELysO1Ft8QI8P7S7vvbyfs+Wv90RWzHcGM1Bq7dKucKnN22ULa7gA4z+Jh+sqjNdgYhYaNMhBQy
JgFsUWE+8iZ5+WP3z9VL+t9DS8Bl+OVqpVF6/SgH9WXzh5vwo2+nc8+vpUayYsqjqNGb+ihJd9Dm
/wpfawKlrQsqb/1jOlyQsSO07uKChixiOu4AhQeIQMrcopmlX/YczJKmhEM43K2pUoGw1X3x50xc
UdJcSIY+YUTDu2Y1swvUZbSbVroEsN4lIrHYU0FOyjbo4NcJkcAUEcpc1V+HtwcrN04lmOi9xRhs
ijQ6RO08u1eQEFfq18fo3JVv0rrnBDIyn+WILt5PR5hlMznQa96fYOsnBnv4CvL4LMwaa3BRaMnP
jnJzUgEFwiZtI/ihrqVeA6ene5/GIvrHGoSsVshRPGXryF1kIYt7QI3d3w0EscG7HbkK0Gumqeja
MZnhbv8IKjUfIDwyoGUdhexd/TMLLIDbzuXllwSh86HK+kGfNNaaNVgd/0Kyd8+Ix3y9uJURq24S
FBEzOEeEZovUGt0Xk0UJ1utWixjX/Xh0HeMVve4AS3JXn+TL/bhmbtJ7PDTEwHtrKyy+C7mX1mp0
kMi8+G9dH6YGSZcTai40Zi506NfC7gi9y8Y5UoI5cnhh8d9dmhv0L/CHp5sjK39dtMp7goo9iPyD
j7NNkda9v7vm1ZD7kl2zaLoOrmHXXoW14WCLKKPzVOhgMJvOAIWv+Rml4dz/ORDr3cXEmh5QR6j2
rWSn6fFlCzGtFHM3PMYUAktabWJhrQfB3pXic7hibdY4RdKiUV48RJBFe9w8ccqJAvKEwikKtLjY
HjmzesVvvcnwqd0mm8xlgqSl5lcX+YJ5sVUsH40eI/07Z8Da4BYNEYtg+kpLa52LJUIhkBb3Xp58
P1wUMR7lFB/sZ+HrLLvC3QG/jSGUoKBGltVpG9gYYMSUnYkhVtYvtWHZ4BDjFL4owqkgT1/yxjV4
/+vwcs8uBfNOx8b4BBy9Hqmhzw8IZuU0k622nVn+lSmsaq0MbWqxPU2r3kzjmSHZFWe5wAFmuuN2
GPArlnQCklgJN2QzDSlpuqUCQOXgx0d+7n7ExVeazhe44LmQiXHbxM7fcxq0rS+ZCA/urjhRaIaS
wgwvasyzWZxVuopFjfXYgmV1uOaSvNjrXN1P/g11O853/HnFuAnHJI53oMMUb2yCi60YYKAgzNyb
vPuptCKDtKq1Zicr5cEStw6fhkJl0UchUOFIsCohVCA0T1oqZ3HH805nyW5HbzZ8OT9RUzzmiUCd
aBCw18I8YIZ5y72bsA42Ie3rBG7sIBofXwQvjG8uJLMNnaQ2A/wO6yM8XY1Wmj5i06G8giNZBjzc
CsDVzFd+KcER1keCBqi0qFFitohrnEjIUJefFptt4T4hqC4lhfhmcFog531wp5mEu2V0aI2vf9xz
ZXNwWjrj1Vf52K/vx1mZ/92JtB/gbhmYcaxKvG6mNSVB2Pm3aTpZNUV7oS26dHqq54aPS4TqvfSg
xOh3KzyPygvbEWg7oYUjDJRws5JC+J+qEkWM0U3S2/ONfn/gwCeM2o7FnbXqSPkNrREnd3abQkM+
bKtlsScP8xzIdPEXDEYiwtTkwBtePZcOfBpORHRDdxuUonxjPgrwyDBJYjFQ8TCx3DcOIRc8njH4
4LedT2y1YKcFjOcJ91+HqUAnejQn+Qe7xck017hy4wnXpugHkD0BukQawH0t4sNGwActnSzxP/+P
OGgmwR9e5MjX8JiO3nlcyWLc/+t0X+K0mMocb7GMStTD//dig7xU/8exIzwIyN7rxbc7ZEck03D0
M20l7TRFVq4oMI1y3y48Cd8UWqdNE84SLY0PnCeCsQItfsJtC+04vuN4ZRyTEgcVd0zL9F5r59+4
m1W4hFFAKvw0591jWCLjEzwAmfkvoLg7oOpCIkpRshdWXF5BaPg0q04KeMNbWSfREC6OW+84rWDA
BjoEwlLQYaS8mqKpLnUnoWxK1YQf3Txpe1d1qoR5TGL0G35NUgOy9D8l1DnLF2sXvKJ9oUPg94cl
aZdCRgTsazWWCv4T0kQ8unoVFOSKNLCqksnXCTpLMTa1qX/WcO3yGfGzkPSvx3Ait9rflmS6JQ3Q
OOg3s2dl+39kGyD/0rGoaUSi8ovHkiZ5dORYTzrJ2lPfIq6PCrdyqxF/0r7EUcRht6fo7ZAi6rfo
Bcx5RU1Xo6wCnniI9OktiYhYyz7juU/ln4yZKZk8SSBxVCrYufa9CNlMU41vpZBV+ylKLZyzYgR/
PZL0SLK+HG+X95GPdQNS8O1jS8msaDGfV/UxNTDktIUPtV0Z471FhKBRapPrPdVcGLE2zWxi8DR7
22U+TlwNS7YYJ9yJ6hvdfne5OFiVqMF0nyeEVy/ULAzxSHriHg4bzfMz8/OWCBvQP1VNdDh7aiQB
/0BwkG0bTAMe07nu4HWLIK/HmjgA9VOd7wzOK0zZdO94BwJ4O2EPSMvS5Ja3VQO+7Pmc0dzyzIaC
xDCMQyQGT2ZgAoFKHAIb98d64m6Taw4fTNw2ay30wMl5OHAplQC3B8u9pnS08VyDUAIvP/LCBWAL
1EfaAf92rfRk1Bo+xqKRd7xes5JPD3a7nyOhDoA2c6oeQN/rxLBV9xzTWuE9zRWlOThyl0m7BRWm
Hhm/1+EBJpHCRGbUHqby5QpCcwzwnnlsH7c2C49hJor9bBHLMPSYTlgVUaWl9O0tlD91bQXLWY6x
eXiCefcTRWD7QBGksikiQF3W0ZlF01CBE/MO1SqrMNBqrWLZzmTEmQ6pjnXKwLZzbEyAypFtliMY
RlyVo3RgwzwUGzuPRmaZveUP2nFw0z1MJxCSOaQ5lerahp/IMej69nWARsLzvDWGQHb3saeUflHa
ancIc1Z8a9Gqh1TldCf0mGSLgo7yaABaq8NXm+nji98FmVEQW3le0pQxFNQnLwEL0mrQml++Y09v
2HXnjHQw2HYX63WPR7xGk58FAAjDZ352PxRse9ggQi2AT0gk7TZ9pR+esvwWukiiZR/CVoe2R25n
Oj98VMYco0BWegmZ+dXh3pXtdDHVaScmhF1CusmQARoeBr0uFh+eWFH2Ytb4Nz7Fc82Zp+d3eOG3
IGIf3J7zVgEu6Pw3r3P3KBUqH3TbvoQd1wX+fzaRzxtNmMQyS4W1ez42VR3ShQHEEq5eOWj7Vg9F
pCqWk9QpYNqLhP649I+dYI6sUO7DKDVyqIt1Lf8gSc6mdQTfQCyFRjaIpJ+NB4VXiymJv3l0ZpS6
XYSOGOAbLEdWMh4gnUiNCcAPeYDVt/p2aAE2EKwOTYFe/jRo/0YD0emDXZNoecnzyTtO3+1STrXD
aGG5bXmHdrHGejEbMfOrJetOsHiLuau9QzlpHn/BsaarMqLf5dnatU3CClS8xlQATI7dch/r+Pn9
7/V0+y2uDyAdtvNw77eCIy8o+sCBj7WJZUzlxKvvIDhCxU+M8Vxa3tQFZZaTfTjOFKvN9wclVuBn
ghXrxNhLZDLSH74D+YDL/YEG8Mvu/zJzVZLnmeIspmQbZiDuOErOtx42SHmns/OJE4hQ1FQSZORU
tTJghgkam0lSWVrzEXctu5AIV0nbxNxpoowfHhUvUBz4v2j0xIvBB9d2/VaBHss5w9+6rKUMS2EK
i8VxBtHgJ/v5m8EWctJZsUVNQU0eQUKUEWFkn6O6HVcTgGtzxhZKcdd4hzEzcRdTkn7v64pQ9w6O
E6o3q7558pV0jDj2EbAnOCX/jrLgpl6tKseIobHiiwqM2xxXrK4sdk80ggWQ3yqAQZmanWkeqsaI
ObvAvZBqbWXZrQYZf+xKugjO2HqwC01xJDDEBS4owMseiSG2WP27hnPUlUbg7gfCjrOJ5MWBw7ND
0l+LFKh6NH0BjImw3Zfop5T/A/y1J05RXOwYU0tomMSQE6XZGSfyuNqVAoIKxGVJ8NMqQjI7+V1S
4CRJ/TRFKOiMG4Ppod34YHhXxXQ4yE0ZkpmOquhoBucrgnyJyFSwlHDcDzrdRN/hO8YIgApqpfEM
8N0KbnqBeGO7vINhOT19rWLkPSf/sK81by7oo0gm7VSmEkJQ7g7oDLeUNTz1kd8xp5eKK8+r0yRv
7CPlomcA2t+wmh0ko4aU4GJfSOEAs+FELZPA+Rk4Nl1AWG0MzaPBCoHE+Td8vHvX/X5X+WQEl4Ec
+cDEf6sKVGruwC1GUrJv6w82iy2J0tVsB+pAnTxH5A11N8CrN+CcfpjsGnhsnEI51ejpQqj2x2Qf
T7h7wl/OY7WMpUz4jtP9UFvFXc8Nnioa+Cyry3h3GxsHlaawskcN4XRrhkRCtVQs5kxCFYvSx8GZ
a1ZrvMJyzqnLBOXuXI+w/rk7L2prddMRJw0GcYgK3YjbZGPp5S5MEIe3FxMFX9s94+IgTfYxsBbr
Fp70oa4j2bAyfRi1XyQ3FHEJri7+GWMnHAHE/XJCQc3ptVXbndj4v3YugJrDUicMISX770RPtfw9
yNoFz9WUTqPSOMH+dOentqxVPQwmerX/86FnpBHHdNgfDPPLsf9YhFbcorsI3PXo3KiWZMbPYaZL
t6j9KGXQb6Xz+qo4NuRfKkTqIKaMvuXKoS3cBta+RavfgfnqnAPm9VsntiHoYdw9NEIgj9MoSG0a
Ubw3MJKQvk4ThfTYA5xpcYpaU1T1y/JVxZDz0OwD1eeAtZHjFOVyzZsUwdWDWLInEIdMJfSDcm9x
jT9vaDOS84Z0HpBsrLhzOtuXX/UzMY8XwK812rLKlhR3KAY7OxF4LZcxiGDNAc45+FG/D4W05uuZ
48rpIthrZ2px4ADe5kvdvFwym0B361yuHcOjW24XmMVAEQtrHAVqKTaoWU5mGLxFN+7LTy1AYll8
hOV0rmO+foi34ZFnthppM66m9wF4EQA8uh9S5ahfs2qQnzANKOPbIjvT7aMePR3NRnnOwnYD8JPw
MxM3A6EKBwXmJ2JbXEDcD/AD2Zhij4TpqAUlJeyMe5JnT0fonnBIHPlEU0gw9qKY7j+JZvL7gICD
sM3l0wLw0HksG4aBlcLrEzRx91kn6GgiFMetOeO2yKTAm2Yna4PIIGAiwP45p0b/3J1AwiCUQMpn
DBtKejQPWTxWxzV4OfoGCE8OSWxdZg4Ujk97OVm6Q/G+v4Vf4uUiLSAFOiT+sG2P3ejCoIA6Qd6D
OJ2JXNyd3AljDp2xrDhapBzYuH7u0xvCvLBUQ7bebrNFMq9MswMmAC97eIQyG5oaGGZUmcWkct7O
ehBv4zegGRquAlfVJACJJu6GgFU4NQ/seo1kdAfNeF6KEtGO/eQyjKkdWPXVcKtukrTRf55JueWo
JSOjNOsgG8p2i+O2jeTWV5YVmSxqISdPW24DnIK/nUGPV/s+FoCmiMfyPZ/DlWpHB1SUCopqfdhK
Vv4stEH9e7e0x1UNyrFEDCzvX0qB4W/tJZJ+m0HnsxZpKIGPB+AJhqzXEnqR130tqPMjrdw0qkQj
kRaxxV+POvC4tqFSxcsXPXfBhrboD9xxe5Qla9O5iAue7RobXXL+ZgfbZ9n+lSBN3fe1HYBHBmct
JZO0Ww3gfTGI8R84xwt31NHL1WpQnqtjioaRkCCuzt2bcURpsOD2HmB9DuUSqIC6lF/Den5/uT7y
L7pOAQx1rNFTJfBaGiuhc6SEN6darIW3iRIy3OIa4qgUdI4Yll8mfswuJiL+NwNDw/+vZ1NC4tYL
NPiWQbjNOpQpiFFavMMBI5WYgyl6Rkfa+OtGvgx2RG0JvEpoy1KnAVtVbuuDDbj8w26BP6gphb5A
VhGWxAfwOtfQAb3DNPAr3IoV/AAzyP/HVWg4XHuGnSsh3sEsVfw5aEGYWe67ZVPoIG0MIteud13T
N1O2nWONhHa5u91C35egMbkc77qJqP3orK2DSpACqhXc5dk0DIDCA28862GFvpfwxQOEDfxtm60y
bYTeYAp/IKddbDyHVv3p8Yy8QqOcxxbb+H3LZQQOSoeUX0VpKFqNqcTRkwd9+qpofPTM6EtA8xW2
Cq7GTwIPS7B05tV9ZbiPlvcUasBTLasUHrzB1ik7jMA3Kjcz98UfKYbyS6OZFayF/HAjO/iVR9Tx
qAvpVEmOkGasn4OImmu41QNc28gL3WDcFB5WAXXOgX2us7189z6fUWxG8uQwoEwCF+yF5bfaMyih
UvG3Dm6O5sxjMjkEnyJbmPJWl3U/KTRwXh8vQLelnYLo+SMJ+UJf7zMNUs0tmfs1V75SYJzwLuWR
FT8/PooCSgYhD7yTAPFCHAzNctJlY6aSWRaGk7QdTPol4YuM3tN+z9DXSGO4OCRvrtrLAHiPAEy3
OtIaEYIddHjUvP54435WVvB3IXNFMiozVm0/DaIyTwIfz3VldAWbjVFBivH11LwaO3kC4+RewIX7
pJqQnOeVz7CgL5RvhzDFQ7lGuczaeAbs2EDrMxneV0+dbK/8T8XF6lrIUNkaiYpS4Cm1RZKjEFOT
V4b/o8Ar9UfK1E+jY3EynIVgmvBxoheK4fpgPaY13xo6QTrMm9kdWYNeqzK4J557PRUc20+XL30t
73XSQIFiPLxUHt5k7cwG/BSehWsEgJ3e85kDqXgsuw5gS4Zytw1DNhh4mbSooThIuwraVOxU0nwg
hErWiIOvzVrGtakVbtQMcM7I8059sygfICwxrma6hAZw5eCGcGJtBLcGvzqvWNjKc9sN9J/rFIaV
IU+3bpPJwyB3qs5koPs6ka+PQpQ+h2NyAqoVyNcdYAlgSwrKKX7OJ8Zg0UR34bfc2Sp3xhnziRrJ
vqKRTtWgsoodV/Y2pbBYimdNvEj5mg8abXPz+RRvtWzAbVLyOkZhKqPSU62v5LRCuiI3wpcRo5qM
Vg0g8RarLJ8YhdREJSy3b6z/aTcTc+67NWmScSmPspA2NecBtKbvWSesXKiQ3B+ID5tRJofdlMuB
zJrTIpcTctao+g4ra8c2ebraLBIvYmoDBqQ+5VnV+8Nq5T/HxSiDJgr1Zrl6U804HeAsgbSWGLoi
qs3RYDj+YxlVI7vQBjFIhO72sa0OG0uKdqnbW8fCklnE+dGRz9Yl2ogpdeG7JL+cbMhc2MRSyjMa
v6wFu94W5Qa3jJyLwUEcQFA9uPNXnPMQE128qwS5FsyMzeNEVX382JUb8H9uvwgasmSC03eMQcCq
wHOm8Uhqvuyud8Fp2kZgzebm9EsklGhmbIaU/q3CKCbViBOvDZXeSdfHx8tbGyHDZ9GLDtIuOfHJ
yykNMrFecin0aDBbfJw1ygiVj6NCguAFTfOUQucurlIZU3NY3b9NERnv1bJuX+g8C3nqlbbH8cKG
26wC5uZCQERXAXWaq7Uv0gwho6G4Zd0e7LioqWIWVHvH3hJiSPbNJJ4Spcofg3PLzgoSkIYXElvW
WjgOHDJEPLWSA5Bp1l6tHtKMEnXGe3ucypMF3W53G2GiEiQaIel6rkHAUcRu0VivReiWBWcNPL/a
OzUWqaXcZmBYwPSs0L4KPZ3k3nrCUidT7ikk3UAak9whI+RINLb0ioNV0/gYS4bP40+l1KPPz1Rv
k9OeEHETajB5fT7y29Hg9VGtQRMvLudCZ/BMaG/VGY3BX2n6jR7gb3fyqkAmCxN2uZj8o/XV6uP0
u1HLIQrwypr29pLA6imruRZdSY8KWno5KXnvLWhEfcEjk/jFvNKZCmy+oR+t7gJstApt8ijAEIfF
Z1WAisD/1+rwI71OMXW344hPtj7VWttV23vLKjzW2vibBJhLPziyvIbiCAEgw8E6N5z/4oZDm2IS
k3vNMDmETyjuZuwOuh1YDeaSyjVKBPKp7Mx+EVHpTDbjsFjVYmMTIv5GZOMH6PjzhseLtkBTPvmN
sY6q3MAAEsurcZxzHVIg/abDKjk1BbR6GsperUUKvHlJz7HhzNeoH3eFPlSgQPmQ6xt0+BjU1KXY
sQBb5fbgsW+YWGibkQsa9x6Ji+GbM1B2rk6W8kJEWVXvmagSQ2DVkaAEcSw0OPiVKLjdeh7xrzh6
tGkgOXB6ak51Ssm9EkHqqcA8m9/aRpKHZK65UJoUXAGyI2Flo/eniCC4GUO+uKP6Uk/qRTs4Ws71
L8cjF6/XhRwIO8TA1fZFBK0HOjaaw0G6rJ8t2+88zilKeyZR/NkDkpog+7soXoSBp7UGE0RMgBxf
fO+eCrkEUOV88/cpMJO4BP2pX/XT71nckQ2JUfkDPlUcF7edit/O6N2y0vNvz7S/A3AXmwEeE35C
KJMjm2QHlwqz0K1V6ME25ESMi/EauMiNQNSl8Vjv6JpZK/jFly7/6FTAc3lRr3VE3v4aKYwv/uxy
SpLIVYgtK/NLVxErPFe6K66mMT5JaoDBXaLvFODdFkdSNMgM4C2ssQutPxDBDOw6jZqp0z0exr59
e+QU3isD2pCChCRT+0A8Oi2w6xw7pEnXQ2Sf1xqaRtxTr8TBJiSpS+fqbaQD7tr06xS4BtlIuVhd
DPN6RnrR/dEIxtDAaks46/RnbAXsRLPQCs2nh/1NB+4gcOzyEubxj2/hqJ+IkJNz5z6PmSTfhn1S
JLvTEAuLerBUjQF+R1vOjAgw010mp4yqDkuyZ7naR2CbNkugOl21Q+f+um3J1Vqrze8UyyTFjuYH
9szrcaNVkrwUxpzpZHkFsz4s6asMSxqUyFa5aaj2pfLBppypd9kDeWxNRLPVKpGefB+C41jsPYxx
r9GHs9MuoWHw48Nd5rx/D9bK2yecgSoklGZnVwIzSJ9hTzLjZ7nSupDf1XmtBeuaW3uceZ4zF3bI
ZOtYTxXzjWIEghrrbgEtHFe8hi9UM+B5F6b4UBBM0T3ShtbUebhvn4yJoF4HouL932HwO9R074Et
3pAPrnkGHQ80RpbYWGzNRsEDMIojNzf1d+spYgTREPr+yLOXoAPV7OPYVMvDi1G0572K1VEDWHBX
f+j3VBVb5eOX1DFo1GcxBi988WS9q3C91fsIksFvI+zCL4Ohm45zq/XhvkU+IS8+7+ffXo47jL6n
KNDxpOFgrJD9OS2AvKODrmDBeYzTHhAyKxmg8dwQznaMYlwa6RGj+WxFt4EQ3pN8g62evXY6DjJh
v6kmiFRn/MMo7uyU4UcQi7wN6zILg1k3n19zGe3GekfnYzxZPnSA2RfxjMDYd8Hh1gOXnVGlGR9i
psv04hH5Izz7bUzBi7Hxsxth3zpPVXgS8TO//OfP0Vx2HUqPSnlC4I4RrVW01xpDmx8Fnrkq8FjZ
/GCyn6ngdLIjQwVe/S41XUqmWxukcnzIbHvQD21xlPvEVC74KLfg6BYgQhoKDocXyZVTkaQVdtMi
uWZSBcsLnJZo+OtbUs4nM4dkhvym5XU0U4+FQ7Dh5ptZdBLJ0na9NAswy/mfJKg10xQ93/+KwUzA
KSkqKPhXyKNgsHovAp0Xttxs1vuLN2vyTTTVQkk6SSYKCUaawBYcbHsNtg9R2Zmluz7eVLyY/QDD
17YuMZrw9SUBU+dpfWN1d0QKoUGtYyB6vhP3F8iIYm4xkBCAOng6c23HifY1dxGlVaITLj01mXJc
FGotzbNWB72N5Uz+DiaWbYO7jMYQf6z9Gfi+yPI6Cwy107x9nvEyENTH0Oi/nAy1+4a498IhQe86
0B1pCRVjwKwJP++NirW1nLics7sGCZmRN3TvGjDJmAqf8Z1E5/RywTGm01yhJ3IZsfBH8Li6cten
vukhBt4RVpMhNniEY62AOm7h750D3mO4Z3W4oWmfD/SHLVEeqnWzoNJdCi7NUTyg0Yd74KSCqG7Q
BIOloolukLhuvWwmUbzlSW1l2H+fJh1IArAwjbZ6PiZqyBK0R1Xvf0c4LWDyDJCwzqqKi6d1KNr/
zdhNnYLJaTSdQA2ppr5nDX6vJ7SYDpevAGi0nQd5CAfpEI4FKcDOI6rql0YS5TNxJM9LZTW9zYNo
8nZFcARg2wZ5b6vzTdKGUKo4xtPgOMNHF4TwSR7IVMZjAHozj/euARtatfRBHd0b/8x2BIMMJDQO
KZFAwx/ufQne801RfKLN8ihtTeTjzLPZE0Ns0icQaoPsywkWuOZRRwR4NFLkVFbuJqg8GbVVuh2t
GYPmrV1tBB1InAv+hkZ90jMmG432/W3wUDZXCThBiOxv0olV4ncxrepY4QZcrU0pLy52xM3ZimH1
ws0LgO6VNsGcLqpHrlOYzOxA1Sda1kWJqWK+Lo5g0QOiCrgsW/LcMB2PwEnwK0Aa5jRXvwLXp0YR
u+gbzWMM4vZE1YTUqb07EXn2H0aVS0sL/u4kOre2TiCBp5mf9cIeA8/GYLbnKD4H4rx4+IvDvnyf
MveHnbCZdZMRi1DELxC20iP0vdUA0H33s7+s/n4eqVUK7dOk3i1LdGDvra/1Pxla9maKAEI+X3v+
cPM0L4PA1M7k1yA3NJNe5WT74CUkYNzqf8/Fw0LWIqAeP7RE7+WYFFcg7kbkSIQhzPwcHhaBs5yx
5Ls2JOUiOtzrQxICn6b85SiyjzN4bDRRiT6ISBgyCBwkgT+019Pa5Pvnv6ZwGyCTnwz7n7GcaVV0
l8uabRwaMTmBltka6zJjg/pVRQt6je9wpSp69iT4gmSSFlB4PRoaExr+cjpPknwSRPeFlwBUoxk7
8QG0WLO7HYD914LuVPMl8UgmkK6vNM92bJfiMOB2P3Ibt86v8Im5WrD9fmfj+S35v4J50B0O7xhz
nhJ8L2b8sXaTDFPp05+OLio4HxcJRG5l7h+9nVcTC6I6r+2mKJmXC+hrpOqWQXncZTEh1O3fMSU+
0d6emEVP3MT/XCMHtgJcq7lCwRF/g/8BY1Ubt2JEphNRxEu6GNQAzD2POTwMaEJV6axkXSNoMIQ3
xSL584oHRMF8EtltZcMa41Di4V4iRI1PJTt8l8x0oaLIgKnDl9WK+bK4zi8gVVuYEU7auF6x7hrA
aFZvL1d7wvmMibQcoKhoD+2Xmi7G//INyepkP9761RmNQW63ZRTqFLfVRcj98Ik9Avdvld6fGLrK
oGLnz/psDGTTS6y4fb0Er35mfvJfKcNI+gKyyfZDGy1NXnVL5uCbZyb5ncrxvQ6T3zjp6TdHC7ZK
BSxV6pqE96v/ZrQ80OHLeg8l7OE5KkrmCut27qBXvY6wqj+xhhQAvESk/q29HAOdSlhp2C5bcHmz
gFz5w1pkS+wD901MMz5MfkS9ocPhpfxuWimoEcjQN5mqTQrgR+Ssf/FdZC7Ny+7ytLeZCX4MPvNq
aUz4S9iB1r0Hnki3JsOhbvA0sWdysYog7cXLmhpkDJAm9BkkjzjetlD/qcArB7PJ4JrKtfEGq3EQ
50gZsTRcAIoqW5fjz7r/vmLjwRnrIRLhMXMiIVSIfDNWnJlXwEA/7wpqVKLs2mua+s/awEd4PzEW
tpUQ0KxuToL5GrTqeRyqiGq+U5s2LqphJ42xsmNopINBrBpOKm3w+XgtNHWWDagWWFfQQ7uP9bRK
zti/fb4Kr4BmA2Er40xFlHAIssXF2z/1RTdSCKk9oFt4AhQcET9rsdmYdxSTmqYWe6RAOApfFQYd
/bvT9aOWJvW+1lZVmaw6jX+kXHJm0SD7WJ8pEsRDiB6vQwR7JjQXPJeBlRoaTy8MmzwGib3dV+uV
kEiZ75UVcW38IOh3Agq/muhjspKvHABJ4E81IvSppVyeXjkPp/84br/VHBa3O+4mMfCtBiWpJU9N
yRBDmBGq2VD79v5LMqwIwDVfB/UFuTdSPWpQFj9scM2xaSVh3TTTR+xPUfVTOEJlGHnc1Bh+AZL5
hXVbeiBDjNB/PLyePBPrvDGM0GeYJM9wUgvhDTcOleaL81Xj1iuSNAtTzmpZWy156q2bzjdNeFgV
thOL5Bmstjcf+tf8mQq3brQTQVcdFnxGhHSD5p/OOXypyaoVE/mtAsjg1rUCn8JJXbaLVtjkCbL7
2418hY7K1+UTgF3l4v4K990/7NF+xfWJ3N7SeTp5vULiTHEEC3QVbyywovIpWyTs+SSnyOUmVGks
hH4xU8dyW1woJHe53HH50F6VIxS/YNR4VJ9FKog5ZpzHYCBVIsTFCnfcl18aD7CNqOTJQ8cnpw1R
k15jM/eQxyzCGHN2aJOcsOp3qAMNqvSSFC2TrEQ8uEHqXfiE96XgL1K3n6q3z04mB7zlfYR0eSdV
VfwumJywe3ahmCqKOqJY8YyDL9UtxFkuHhM5+aUztSC1OtU2qOK2MoRB84mP/un61eAJ5WPIbhyj
Ys8795PSqPEKniYV63+BzfO2BeNi8X5F/PZ2Q4mMWkEeGRlVw192CfuCT9/akw+g2zl8+dbmt/lg
47ZfL+ysIBF9Tqh+yy3dNbHditMN6sVUQRncYSkWdDoCAkxKg9gUt4iiw7/bKTBWU6f3dFaSuOwk
MZW8oR+7j4V9vkN1JQJtoZqJJVTFFL1Iv3SsSeRntZAdKEqFUQbGpI22/s4uF7GUWFqWLkWmpByW
fYYeJKpnrpMrIfFITaBy35Cb6t1Z8y1Ct7lKuERCfgrrU91jGwfc0oHV9NzRRl5PB3IiGq3gOW6i
y5Y+F4KpgzULpdWgJ/4/gTbpsDlupsY/r5bUtLrKbXjfxf6FaonNxsP2mJP4FUtZNkxFVDYxnyTe
khEMIaOVYZMcOTbUvIgBWNzGLj1+vglWrYjhjBthDU98Yacw12xE+yt2CUHsq6IyU3RecZV15r4T
DVkWguZOofuxlpD90r2NHh0eT+aRGpuuaS9Xw9Py8pGzlmYPqhOgSXCNqfzlrU/OyIZ9eomX7EPG
U9uWMYZyMadhxX1mfl4+yA9mrV7LnRs9AibbR1J3DZVFTrX90ET8nTQZ70HNwNxiqA5Tnastx5hb
ggCI5wdkE+6+kgd0qat10ncC394/LcF2tXivxD/R1xVcyGK+aDC9N94kcdF0k15q3zWUSm9TTHvs
kh43uNKaaE+gR0sVD5i7Z4RIvjQ+1JFmS04oc1rhyluYjdm1/QfdJFmR41pTCnEcbHsCj4pah2wf
ZSPJ0KEhcrD5KH4O/JnBTtzTuVOqKgt/Vc7OIptohEHrwXLVJ7KpHWYWmBHjgJAFVQRpOu0AnQJv
aLkCx5bbYQdY2EfS5TbOW3+v+nTlqhWPgjTyALiz3lz28H/CoJW5U/iSQDDVzjqHugzenRckBzGQ
bhtjGKFsBoxPwXRSS3pNY9EWsFAtJJ25OtrHw1Qput4G/at9AWnm5ENNTIronyOH1+xyKCnTB0HT
szrdJi82RshBMeiy6g3za/p8Ns0dmkVk2nEphOmngXBuUbJ8YTY+JX1ynkpTBPBlcOlSQ2PM3WVe
kSu3gPKth1jC5DXHCYYoP22RL6QpFMD6jHj2y0HYobSgZaY/Z2KoTrnkayTF0bpxvMy2+mj8sAYc
ZoLI1WhrCaSMy8Li7hLElNds138oSepTEVUviPJcqEz6CY2i25toJvBQgpeCmdfYHdNCV7ztdK7Z
9pK9qm48zStkQq0wEUv8ngyBNK7aRPknZcRXp9Rosjgk7RNLQPSGwzX3HsEThkhggkjyVRo23arX
m+FAQ/teXmQVH+n6UaSZbCxGR0rqEurYKbUDBG4UJRhACcFGx+l2ySnzdELbgxNphihlaBZRI7Yz
08VylnV9b0zPlqU03drZ+4XNlhdp4/p47qCJfuSMI1/ME4ocdG3He4ylKSlKKaDJfW9qQcvW8VkK
PDOciO2ufV7SIysNlUcd9WQU48GpOsQKmfAOA0dCSCmIbBhcKZhJu0o0PsUqnZWHga3Mm7kezAjN
8kwRoVoRxY6SWo7xzm5kodLqKx5DiBPN95c//wCpZ7ZBtGEMgpHwCnhq46EZh7N+1K7FMQ1JnbzS
kQVhE/UIiI/W59MgU/wookLCmxnogDAn3b8NgsnpRkjS/6b3Qr3BMeIc1WPt+4QO0rmb4xr3fzXh
xoZ0EbYFJnFvyyFGPWiVe22NzqV4eUr2xx2AdSHkDUqE5fVmLCrvnJ7WYH5ZOfOm+obJxOmiUM09
jkzGNOUsnb/SVz0dRSxbUmGRvwNDFEWiKVmlhMPzFN0fuA4T9/zrpeF3bqFM4e0rhTiKch5rBNNj
ngvucHJuRyt1QUocfGlRpGr5DHLqQ2WplUMytH3oU+xbHWg57FnMZD6wFND0WKkEVsOQOCCDLAS/
3/iFHam9HP1G4e7rNqLLwRscFgDNRmrDcBTnoX6kN8nu/Pl+TgfnpAUIz/V5qK2CtydX6n/HE0hw
lPfA8xyXUzFElS6ZH/Wk5zzDnmPvae8byU9A1HTbUURJhEP3qbQ9LM/4vT4pO3Scfm5F5MLZgyZO
YI80KTp/drNAsc88bcMQup9uw44WQzlZ0icVsZ7cLk7lflRdZIRISGxtI3DLhzUiYck4fiihtQ/y
xH9HeHocsxFzZNKRyaCLUB4tpiaAHcv1yCjPog3PmvkPP6FPg9AaYfXqWsi6+JRlJ7IxkFftnipR
Mmcs/+hsB3P3OhuK41oc88NJNvJ25r3QsLeUigPJLOjGTVdBN+tg0Dyju2WF9DWK8q8RzQKq4yJI
z36AQrhN1yEerT1z7HJOOBTULTZ3RF9jiOXGlp7e/UblprOUZaga7JCEnK51ECsE52gupaW8GoAq
3bzAHn3WuhwZbDZroqdG52gdn3cPkSyawSX5oy/AqZdSyqe3AlmaO9EwFUthsKtklRKXru8FMLKC
mORzvGxh+aD8YIWmRqVnYFimwdynNFXIZKTvpyX7s/bQe1SiFJ/92K8K3paZCuFmOqx+zWVmbp6r
JSVut3IETIaBnJHvGV8tTNxHJdEETXZju8FX1Uh6SfN95bq24rAdWXXhfs8tqB3Olv3KAtJlVKUe
7CBAoSsGQHfvEyyLKBhomnS33xxYAHha/oQuUqIoROxs54xpVR64gocMW5OYVAlF45aYBraaq/kO
P0DB8zALBsamMahvBskA7KR+jdyHpvcGj3VjyBBZoNS8kTFYr46gjeWoXUEAehaNTLdrXLn4KbPk
UkWsFFuMXtMRjYUgPDxOG2QForXOfNG80RsdaLTfbL4iWqozlSvzEscHuoryT4NZf4groG+FwpmE
PdQQLjME4KsT69x10WDTYWiOPFek/SPu6WgSZpz/AAs+W1usgAm/baKw+mkk9MLI2VPDvfnfNpLD
M8Fb2won6w/xdhyC0RvfsAwoH5Vh4fEB0U0SiIVb3Xqirhb9ZkJjwC2H36yKmricHHbUrse2L9X+
KNygt3kTh7okeTOUwluGzhzn/M14a/CP35NtC1mKayvb7FgpDc2QLBQRIv9bddSYSRD6CzqYBk1C
e3JFuM/CuLbrTYPGj4DPtiPG4l5Alf2IjQJXqUukWWVESo49Fk8Nw1XMEdePF9HmmSQFphOP5g6v
MFUDfo/xcGDHuw0QlELH4Y7LORzmfKPAYLGDdcAuHbA8abzDJiwqfRpwBLKc9u+tyO8Nde+j7cwW
MMZZdkB7PsbIwpD+KjxSn3ctdQkvJSciU790NpzYaikvTF0RRwVBC3sYZfrAMX89FGNq6aNH9SHl
XbuwEQAptfGBLf2p5pOO084UgI2d+OAZhsMLJ5kLxAXYQptrB9aTv+PhVaQpHX0OaYkrl9qIh7Ry
2fAbLBbY+fX0p1hy+nP0ZiEJAJMuuRQVAN5ED1lVt4mBkVyakGpxbmItNzuJOtE09PBFUImyjSCc
gwU3IiLc5xXpmTVi1oZ66w93tq/gQTuHqSg+HKBwvfwWXKf1ryxIw70M+SfdfdiEzo8MOVhBWiAb
ecgf0gq6FZ0rpYffYJVHLpyA+gwIUspk9D7+PR5zIc5AecuUQn+RvwpCpnKJbv2oDlDH2ZLc+UZj
i8RSz8iWQHSjmYavKALHr77wskhMauGyouURZt8L4JZnp57Q6hwleCPj/ab5b+WiKTKfvNQSItRl
CBkJeGTlbmlc+vR/sh83/yEz0G0xUIhwiTjdKD14co5ME2NbBkeSxsLKXg15zvaNtq4xbnLM4Zdo
60d1fVd1zev63t8vez/HzxlWJb5HKIJFMbnZVMqZ+Z9lfwJw3Uf3uqwYkZmOBVc9Ux0ufQ3HwbC8
TJTLH6QK5P99rwjg8BfT9eldK3z8hbilnkpHrQMy97FE811sfK+oltKCUgLKttT6YmQPqD2k8Rew
4EhjhPhEHrY27oYKV17BvKu8zH5k62jbBnVNV66ouTRLRZFlOuTaK6T8kkQIgGk1+Rs7KJJNcLGd
nxSu0/JhvY9ZTudeKR3l2UErnmyT6/7jCq2Ia+yDcLvITLNOOyiPJitzDKGP39WW5CAhoqTJK5VV
ksEehSIb7O3CUWik7DgqE0FcgOKhihHeVY7Ux/y6Pnhb3Bzb+swuTR8NEZdCcfxg1p1OOApcRq3a
knqeCwm1IO2W8XjECXod5R+5Z5BbdFu03Cr2xE+V/Zsz4GAFJ77WXWFhvw7Rl6rgoKdRFPsgoxm7
iW230qLMVoIISW7ERCLTK6O0ZvCFB6lRkkB9Et3bqXEsiW/oAcke4gHzny6MZoVW9jnzU73AIMw7
2o4k1G++97ekAutefAdXPUeXBm9cHYxaFLLpiX2qW9lThIaDmHlfx4dw9Bgo+PnfQJ8Ui2T/BRGs
XP6w4ajE3bVrfM+2LpeDggv1d1Gpw/5FxxE04xzlQnaUevT7gvndokaYesjnEWXD2+881VfN2yFy
cr3SxvQUPmxa4uJ2m6MAvxdjfJv6anMesHKFYRmG0w7Ev1BUWb3XgpMCdelj8l/QWvIJxmNkQGK+
sA5WEU4nXQlpEB1/cUtUYU6y8oy9bldjVOsQBMX2XoahyZOKAF8F4zvj/CCNwHhFAjb6tP+7A65y
5Yz6tY2PjdEgCURQ7q4bdiqWAv6/CMEAFCTiNCZOMgFm5J9na5kTRMCZZRcMOkQI3jJCKBdKq44x
r/7ChmG99mQICwtPjiYqcc647ZxOkRcbkWMJT4iZjAMY8NmMtZC4FAhn0R5r8z9qlpSzOIosTxCs
v73V1/XgUyP47yXSZTsVRsAHAfdPyGs0gm4iCn6CH07tTvj8DgCFV0Ms/km/9edIY/qxXWQamQ+1
moanpsdaNP7+qB3+ssqOth26vXNCOAet2pip5l4A1EZQg1M4GS3zHk3qsiD3OU7978pxB546mLjb
/y8Tw777g50fg7zW8Hq1qU5xvHvjTD8fK3zHkNbFjHJ6Rcec301XnWJt+FQHBB1YNXdVZIvt/I/l
4NtNfssgvg3pTettUgyrPCZNSFYlz+Ru5J+t+g3gIDkmuBORovti3mtG6T9WLhL1hdqm0YL57MS+
kFFjooMyueovLJEQFs7lZqhApanXN/L4B8XOs5o272mEIVJqfpzxHzliD3vLvUMUDiVqeqLB6KYV
/fL6xLu9U8FwJWCS+EciAcgsH5vntOLCUkAvf10XTt9u5dkvS0FOJkty5nxDpqY7/ApIeYPZRtb/
1y/SBG+8FtJ7k6Emd6UKJYso8QQ9vltQAsV0l7Nt57n5dK1ChtSpOH2Wzff77Lmep467M78WhZfw
oQ6IsgImjci8loeUH3ldRprcSXYNmYMj8P0ZenAbat9slT5okfec9MXSWrUN4PMCB4csafQJIHBQ
HFjgNK+rxXz+75EflX3CquJxh+3ULZPYKG6rAA/VjpJAJqzaSsr+VErM2CQp35vNsUJWurToZ5gz
z1LKGYuaKiZkGnpVrkL633O1fqW5lmoRK5k+UTfN9rSw7uCD45ldHSKtiR2fGJHPm9XhDhUEbFxt
+gEYXv3/xIGGUpNsyFxJOPntjc8rWDYrvcqF2kk+nMP/LYIuGpyc7Kr+15fF8+0z5eEXy4vJxIaE
ZJ2EMmZoVo09qtPoHoViZot3iAMqkVzlCh+RJdtwBjKL9Q+Mk24ZXS7wA+wIo4rAjjWE0EMDSX3S
cynf+irMXYqDuKDc91zHNLgUAivPnweUt/zwQ3rTps7QsQXa/3M+oRnHBdRLuGO7aWNIVqYSgRog
oJl0Zdh73tWMfPZ2jO/k934m62x08Jv0WIZrXOkwhIPH3hn/QN96PIMleom0+GLpqK+sr5kQx+VG
Jq+WzwcL02x7C2GBoPQV0V0f6rHZnJK1f90WIz0lYaj+aHH22xyGVPqiZMEeo7smwBhZ8oLN/hps
cOtlyOuQSGOBX5JsECjtpEOT3lqznezIH21toNrTBkGI82wExPMLrcRsnPuqqFTDlljuIV2uhGeO
2X1FOL6oD6NM+bW7Rk1rAePwUGuhrsnzfUazL6YiFDPgUYdU7Vu62VKMontwmBGkf3ALkXDnWnr/
WIqwifahBn4iBguP+lrYYqo5wSBz7scUi5ZnFECwteTk6biQayQa5HYwO2NvfnHHGFo497JYh4Gz
2sOWdG3VqIWfU9ryk05OWudQtdlUWjH3RkOm4nyv+Oq+uAkD8p+w4FD6kdLsfx9/9C0u1p+2KMEd
h8L0vrMQJYU9PCvobb5oU+ZwWvN1PVK+ewiO/2WW8thrATxoRqwCbX4eIXu9Kl/z8N+JNQbi3dIc
tPfTgBkx9ofhCdLo+7OXKWEobKKcmNrn+RAr6wQZUQTBzER5SrZ+EKuO8sQXAWvr+x8ysOf0RW0d
UMwp4uebT6F/i2wTH4bq69Wit/roz0dTkAOIfS89Y8TnodZM8RY189KuSckdRJgj/6J75fl/x3/N
m+GRTOOafDsj9g56FUyRF+rthSgWgOSCTV2h/VnheHU3lYryG+cX62S/vOX6ulWU5cN+f7IRSrZR
DvQ6j6DejCk0/uKA8o5LBY5ljMMF1Bi7OhThinP6VJI5vPoxaUHzdX5jz5J+v6h9BMt5nZzLdADi
4skriNPAv70GMGwqu2WRX7CZ9pSPn+4PzVGcCs0vwOIMTxNCUHUJsuuEJ+xoGtsgylCUyBLaz1O+
F25YKqpePTh2n3zFHp9Aql7B61MO6SR3XaWUQmnMK+TFMeBoiDZNFgxLXyPLNTPJAgupMjhsjtd/
PEUPr+JvkvGQgBbTeR68V+OFZuvIwCzJ1JQEiTOxZ+3vDrEyNPNbYj8tN4y0FfSOrr036upghOAr
/tN6litUYv6BUt/pwrzJ3cdr3axgGHxsTAQmzgHkODgVXha4sSTz2C9SRFmwKURYKgHalgXA7aZ6
smu6oiabB2g7z0K5jrn/sBApWxQPResKvpj+rM0oIv+Puk3HuSbw6ziwfF0U8mY2JRNAbd2TB+aL
Su254gJ1yC9hfBjRARbFm5vIK0xTMXO9vsf+JHToGYA4RAHjSQkCWt1NhK2TFW97oqYiUtKtfQ2L
bEket9pkpvT0JA3IR03wJKgxxIrdVkkFLq7nza7qWmtJrsBoWeUhKO1H+c3To+LFyIXyR+nV5IZv
Yvt84NWcJEnjcTeRQ4IMP6tABYqbtP9TidLfQU4kRHPqmvvwrAhoCq2Zvh7F0Cx6EdN+fjwnI2wF
UT6+qGukIRGLQsfzeLueWowGKFfyeMZ6LkZr40jgBF3Zp+xSJfvokXW+5kmnVgMJ2UsQpSzAtLC3
fBwGnLRpYRwNHuFk0M45aejDuzvCBNreZchNxguOu05q7A2sOEHBDsT5DoQ9ahs9Lt5vvZQqeFOI
xuoMqv1WSPIHPTBGHXPjVlwWxTKprYqNcChNPfRfsQWB7xq2SSVR2PlKK5RIYxqL4F5CcMtCP+Zs
tOhGO8xpp4Q8ntvnKJaBn+T2r5hLV6KYxG0cRBpVou8B9DY+sh4PSrJkYFquETIcSTlbqE/jihBB
oCdg1KmVTRbF8jDz5RKB5cI42u5R18AbtJzqm6MAhMIFldOo5ChFn6mfZZk1rokSZJd/IJaAFl2l
lYxXc2EkziBVU8PaDsYZAtg/7VI4PjwdYLrYM+NQ8dm8NMoX+nQzPTOtDNW5FKwVZUaLLn4uzsFc
tBRabcFmdIt7PwtQekitHWsO32stcK67GeSK7FR8jVwJcfauADr3E1fp13Y28ZTyEQjhQLud6a8i
gxODoXmOiifqZWgHklbTjqovf9TMiuZ2q8DCiwxHQi3fO/7mfy0QO2Zwn3Wvueoi1l6J9te+dWhK
vSl48IiacnNasJTLUi1XG2oEfAMKvP69z7/jFfOd/EN2s8EJa9xn6kbH2PJ2yedyJ6bcn6ZbjsYd
jdVe89lLCOjBCxf/qNcUTQchS6wKZD355uSHPYEEpK113SmTZdxfYnbIopDjGDmHUmmcJG47fblp
RCOUataajAr7bVQDbtxlv3Ax6yxTtbUZJK4+8pcwO0hYksvJtlI1KeabRs9gYd5b3Oh5cu84IhqG
4Skuav46Yjl7CHw76rmoahcJAV9xelvjoT1y6qDQM2kI7RizZqtH2Tga9SyAzBJO4eToF8AGmxpk
v93HMXTwnjoX7X/qA3MzzHa9H/YHFVGZWLk8IXiP0thbWxMraaSDfWe8nhTKjqOIclpTLeIdtpyU
8QqYBr3Il3HrE//Us6jXsWrTFZo/PoEYycSQ1sl0pWeuvvNESBm2abQuZJPTJbgT4bpDg7JmhbeT
AumQvpyfAZElOKRMRjrg+FuDmqVn+AyRAwaXmbexPidAv962Q0XoZWC5po40G3X7oeVP/bpdw7Qk
bojz9S6J51AOOWqnov1jeX2lvwsHkGKoYhqBkMyK7a+xLMK2cnoKDo/9fuB02zPiNtLe/Qp7gcVj
3VRxvb53clivq+Ej+0uIp+M4CAgL+yFkahPc+/NtE7+p4tpkl6jWGG2dEkdBWxcFFs2U003LhEm/
N/HHwNP+2lljT5x8ZCN9gjSysg+LcKStv2Nv0y6yaqbfH3TB8oaGkpl1OjjBw/0H9AylKn1VXTEy
TybQb/9+MPLASbUx/uccf13lMH/6O5X9Q28WlZktzSXx9mU62d4iiRMY8pVCxE46ZvW7nZOk5sIr
sgfSPNa4EygXVZi0cyFPV8prB4wSIg/idqPrU9g7fmsvGbyhBZk4JLg5x8Iko7ptGgxZkQacpBFf
KXvppG4gpsCBGpJdtOwHa/IpEOlALVelDfplAM+fuAcngBmIh9kOj5x027hnpmXnxhkyrmF9FOaT
BO8KaQYFHjcUXyTIJKhCnmN0J+Pqy75/RzCc5PZBMIVhw+DDD1eYLYujEbUjMKq1TtoQ24U9BFuC
dI5QNbaRodyMFrEO4P05CuXzlWPf2hkuqHZoWN2GZKjIT1B9uRg1PHl0b33rN1aP3gKI0JzPVabQ
VRV+vlYP6f2qVWY3dQCDxnr7wqzwctRTgEj2FhCoJ9OtnT7CrrRARwkOmr4JxD79L8hyPf5wxfi8
GIl/fmyMNcIrk4r9qfkGnAnrlRSyRBzhfDJMh7ELtoC5eMFWQviV9JiNDL7209jJgbNCc0a5/hu+
p0xq32ULB202+U7X4VlAK1WHLvynJ7TkMp+8L4EGAca7hXp7iDRO3Qs1TeyrLAxpYbhh/3no2c7B
KpgpER2a/IVCndcbqrjyEkONPcopDGqLihbFOxdDWvgHSdtQsFEdvbIpvaDaAU+lcEF/HkddfPaO
On1yUG47y2L3mSNKFAaCUnQF/BHmcxFh99oMiU1t89beJi9bMrqbb442t59QqjVsCby9SWVRz7P1
YZb76rny2o1ELDUVjYd8k3ORQXiTGGgPUrLBXF6nNGqf/3YE1z1kNyZVllP3iObnqCHKwfZ5+AyX
nnkGIuydanCm16BUwcSQNJ23MQFr8f7ZaF27DspeHvtNkalsMJfXOahobkKb3c5FzsJHcCF8NOWx
yzEWe5+XLf/oU/t/chb7MRXa/lOZXdi2Sv599RGy7L6SNCp6E4O3BIILV4T7GSxFabMe33/3ICgJ
+afRqCEJMIa8ier9DjdvV54212sZuQEucYE5ZI/fz+K0Zpcgcn1GXyvGuUt21LB71XaAyAelQ/Hx
nu+rcjKr4wtEFGrQKH99mLJAjcc+2xwh8/HHgMvuX0z9xO1dsqfZ/l//3C5yX9EFStHLVLO7zfBU
txxrI0NajSZ8KILSKQXC9c7AoK64gRNX4MuW+vL9uiVAgiEIEyWFEez4qDtFmI7MtnwPEPYz/PYO
Fff7q44bd+jHfvnNEAT76Dzg4fcKosCwrl0V0MqnkRljGE9jEw2C1kteNC7N3ZmGK3D9AOwe8UpR
OisBZEldHxPpQ5Bgf2W06qfERW+SOEq4pO0mDpJ/4/YJ6siTKpmyWdnwtHImKICy/0JMs+JYFwyz
8xnC+Z5nCCk5rrAFaalWrdIqw47ia+n8ItvJ9GJEGpNVqjYJCz/o2eMnUnOF22Vx6VQZsuiTp49r
kXLPm14jvr1vMlKKvvbdF0FjP2J/N3jVYGUn6dNvph4Iv4bmz+gGSr6YRx0BEoU8AlHLk0rtb+aU
uu5UWFuS+ILWPH3FeMHDxdoqCufYWBzTPdC0chwfLZEkGVexK5X+nqvNmfCS2qGccEmnipoNhAVk
avGtfP6mMBZIpqK0ZjNQITeTbv+5UCZHDnXY3nYca1MG9/jRzUY099JedkCnlb5zM1AuPsMgNbm8
qzn767snWRHxQO7Ij9PF08urJ+2gzGfQ2vUvVyYQq9Z9ivss3P93Cc6Bef1fay/BcEb4siEjwK3T
FSdOg10ovisWEK/pFQv9mpgN8f6YeNa9R7NGawxnfe5tI7olUllaJgR0kZc8/SvVqosYRPN1svcp
97elKlLvdmrc7P/iX3c/Ut6kkQPzzLptxyzz9600F+vkk2U+9vrQrt7kD+7cVfX8J0hH3blYthLK
/qSpXGju9uRkVADW4CZdLWFGr2jZGxP/0/B+p9j3I2RKKlcgtnuZcDdQ7uJHRXVUlLn02lhV+cPN
0ANz3fpTdBL7T8vZz7WobQv3Ir9ZB98OkWvfJpDOl1t2Ha9cgt9VmK1+sz7qB5PCOaunb01xHA/T
JGWtKFqe7U4cf6r/kbusKOhGkiuf60P1yE4MjDqnL1EIb2UZ21u7yy3stemB49gSmN/IItb7/RRV
CH1nfuxL6sbmbJTlX7XeKBQf13JCCGJcuPdWV54o+uWk8qC43Pucd1pWJTH7xD4jUZPeRNgdTxER
43s0UCmlx/alb1IS8WaRfAvlzLgp/g7MvZO9aO2wGdT3b+uao7rCDO8ODqDkBAxp6F69BfsAVFAx
b79KupgPIyfiFtbUMZCPoObxm8y+VgVxT48gugX2MnpG+mBP2EBB+nc2t3BghExPohJuQz1Fci1v
3aw9xAkur8qHbu2MClLCghDYsN906WLL1uVM+GPHrqEf9nQICkzgomgVvRr0iyljzprLLawLkUbX
q3DkPVFxAebd7boCvGL3FngcmavnWou/utBshjdJNvFDaeMc5t1XSagYsvfLxJ0B6mce4Kn7NsAQ
A284YWSlS5Jf1HhUoB3OVIxw2m4ff2BrI5bRQGJ8/Mu1YwMzLpfVw5SVhB2sbFOOWA+GKhQN6oTx
uGHmIJZyMSOPuf1br+B92v/UL5UfxJjIF8C0fQgUG9K+KLiDNvQRN3c6qa0gFdfC+lXr4ReeQ4pR
Tj5FgAgGCDu+JLvHlo9CLEOCsvs+ReeYCPeEkEL2rlCa0HSlHkOrhyj6QAlrn9YB4/Vwy9seJpba
I0afpoMCe+vmm+9jcuRcx0/ngMxpVENzSYJjBI2exwuobtPk7sxKwNfpCuxyqpzz4x1rwz1tiBY6
l1QRQgZwzPtbstZRRth2vzZln+pFQvr1+9Gm64sIJTMGwbRoAasGTD6zu1/r9fDrQmyAgI959eNN
s7mSEixitVR94HJght767j1El4soVzNh9WK/0qsrLz0gCNujwYFsfAA0tZRWCzy1rZDW77lIrBst
Z4TnZuHjigEQZ53hSg/5O+Hqd7zj2/FQYFwh+nlgfxlEzQH75AHoRF2UXZoKWIRfZbZp0ukknltA
VWEX04CIX3n+M+pGMI3jMlGGXKjg3/Bxs5TgMr4w5CKu+3zaXlIxgKXtDO2QaE9L0LBwJQhbs5eH
wN2cpKN8rBAhbiseWFqDpekUxTe0J1aRdGu+34rdxBOBQnrre66QKrGFpGnwPopOpHj1J3nQ75jU
6Wz22O9XI0V+D4iqgXlydEDDJjuyPrFspbRQ2Xo1XhevmwsPz6PikPcABRb7vehoee6aE/fVoZR2
55gXA5XDXkZP6QW79IRvIBYY7K/6GIoReMkRg/IN2BAkZFAugbWnXNMSd6GwCXtXTOMQiAoQMoWm
jSZVZftafRlNE/0bn3WbXr7kNsa+GjbrUzier/BE+MVczFoeaRiucHvfEbUyPvBqf1WCbxzJrUrw
VUpkPghHaxtVvNQBBpvV39PLVi5KncR66HRofageD6Q1fXpo1RVmyxHAQI9qIkJtROdfL7qAHtZ1
ocFCQo8qltwK86tRduo+Cq6FRTH2mQTmDdE22yy2qSf05SlUrPgPlNPnGMWTY0sbxY9OWruedqer
uI3jVR81SNLZlPJYZm6viJgJ5KhWGTTwrCAtmWDwQYis8v1J0RilobcGEOakXRCI9GnfFRcMpN8u
71eKst+o2RU8MrDatT4d+RIEDZiVlDy9JK6OvW8MQmsJtr6CZpSRL0CNeWFCH77E7SrnDyzrC/Mo
aSHY1Q6ESfM4rig+nr9ZNoFJof3cgxAkuy0uWI35sj7ivGKNAiM9iVEN723ii/RILK2tYobBBz0n
AxhCuWEoMJXNplNzbrGuoqBq5GNI2arRPUIwvvGBM41Blax91FvFTDTXt3yARndPPiow3hLqmqBS
twBI3QYotPqIHZ88MF63Rg81iDovGO6s3Z1cbT5b1YM9m6zxYjLkVKCuq+XnNR9BHgH2E6f949Uk
55wum0ugr5bm2mmPsiteFHNuB2tLwwhd2oXh/2YFIX5blniqJPh5wR2FzbQdQLH0JR9miOWUamvp
+lD0nfzknlb3T4pSQfQwmyPmM4LdUS66BCnDqvsywiKDI8Q1863Y4UAMXxjaUFoCC7hXv/wZEroo
ViJyP4GVT7gmdkBCTCSGUmI2KJfkL/Bu0V9ZQLem9n1AJjWoeWXaqAdqai5I/ARRrwkmV/9TCj9+
DpgsLq9CoiF1DlefZnpU9AZlpZlABrJ+pJiA91LxCggJCz8XbAA15YSrn4Tr2yEv6QalP+pUxG2Y
nxkRAX7NgkUdo2M8w46oYq9+A4aPmQJ7VQemNyQig1dP8oXpDXE6rfGYtbQSSjLa9BFZl6aDI/2L
RmeuG5aQLIw/InhplG2vZkcxZw+r+nW9VoVb+0wgMfm1qNz+ww8637t7z/cQ3kKpb20IB5syyEBl
8QaIrVaGzmC+N23D4M3qykMRYm5tNWASuvWLyEd/dTPSuduCK3Fw1RCbF0gEa+7+wq/fkg8iVIDY
uZf4elip3IYdaVC3B/4rui3cLctebN4hGGypNr/3LDtwOFxruu3TxdYqaYnV4FOpz95gKjxZoOnZ
Q/Qvd7P09nFS6Mg62Bu17cAo+fGBbWzi9LiHjpZDYInHZ7zq8eWa9KeyAgUezJUR54pIbMjm5cYe
yCst6QMBzdfYgISnO79BFSoya4w2diJJWzs9P0kKFAEiVukpKen7tXod7uxU73bvIkYXsYuNyKXe
phOgm9WKiInldWD7f68CQ1Uj6wrktRxXyKsko46dvYasO7mY39FnVAT/RDZzQxziYcgXFhCUWUwY
A9sdeBUCBlnTkS8znUa0JBql6ZfMkj3MpmcNu8D/Q57PpvISyUDroYlmPSv9XmxXtTfxJlhN25Th
355EOXPefNWTTGz6Cc1EkhOAcfONAZVS1JmF6hZvYIKKQGfc5FlYcFw1D9Z+8hIMWkYTKYWI3T77
mSFBcTA83Rbj4uRc6Z/w5sV4ariHwdDLPd3bz8BvN/uyTMGbaShucFsz1+KybiWtEy7+DNY1e36D
BzzxLwlf8944U0KB/N81prwSGn93GBC+g4oN5ONENvWVwDzcaVooOkLEFxgalFthV5dL79qsdQyh
WSlvXUendCEz7z3Wy/HgMZhkZEcWU4RYZfZotoUdQPwAVMOSM/MkyUk6lF3/8Xk+34t86X5npQzl
TUn9IfJDxWRPEMks5ONQyglzX374uGa2AepQ/rTVU6Z9bgWgIs9MFNqrgUxkZmIJQNcfSHjiIWPw
alrQ0qkZWp3yEStL4SUxe3hWTaYqnn8LAnKdfC/24dExRD7JgSmIduo3tmETinnx4A4tY/3uCsv0
SOITu5E8YtuLLqh4cQ4u8iKkKdTY6BHsS4+5wBKfNlYZecrc9WMc1BkwbCQIZjAFRLJEg1XKS6OZ
td1CG/W9bseyXfl1B0JeByUMIiNCqoQGvaNE4zy+OHNh5wJC4XtevrFjn0z6kh/H92rckh0lQWQr
hBYKsmURUEt1s7dvTUqzpAjL4rTlFQ6DjUf7YeHk6Gt/uj5zLYi5t2cr6o9QP52BvF6CEthW7S1l
lrVCRMZ1lY3Tsy2yL39VhrjzQVRfCzFlmBiMSWOtJhkGonURfdRuAzluUlFid+c620eiXAcW5vcL
a1h1cMQ2tNclyQNTXTwglbb1xFl3YQmbJlScYh4EGOMTSjvWR5ftuUaGcrbEX0/O2E9MTJeMoLUf
rEYR40DcWgZ1vlCDGaq1WGCDRWpDN6Lfc5nvgN+3XK+wbBFvPR+0/Lr9JN3064za/seqEEyIwMU9
TACarnlFwXnim/BHQ5bV28vya2/3ykgqeLngu6qJ3bkXGVsx70TSvV7LgSRYzaiPgxfbs96Gp/No
H4FY9HQ0RG4DTSc1RFomD5Y7F93xZvx9k0HH4u2sdpV4FyAapIxD2nFx7cDf4I8x0NGglUdypm8f
CNakmLaPjAseuYQyuQ7V74hCjl8ykHUQDJo9D3A9OMISJygAEJvjaLkK8bFEA6STEi0WLl3LcJPD
B1nLPcqg+TTlp90FX5jVW9ZtjWeEyeGXUp6PNMLDPqt6D9GrRE0C8vCde7Qx2JMcRZ6GgIzSkrdn
lEwqCFC/rYPvxPYtr/WYpFLg4W01puvSYPebN5CZ5it35effjwgWZ/R+Phm3yOVPQ5kZZPqLPplN
M+7dGzK7oL+bsK0iFgnjw4EJDAW6/4zEAqfGikeM2YHbkllZ5736QGhM3OCy7/jP04kcOWoVs+gE
k3LcNDS1XQjVCs3xPwnwvTmNWtviQX9tWnENeaE8XH4OdrvHUt/eWq7p6L/3YkcpWucMl5CMv8VS
yOIqyFyBoxxMvpiEPfASt+s7hOTgTj8vq5cb/AzJ+CwdlTrErjqyamMRYsXr0W7/MMlVeWLDZygI
ZHaNdjjduEaWgEHeli3VmtUilztaZuWFtIVoe30Ok4lrmwljLSOvmo0mzFMNbYKQn181oAciT3hv
cYKNSNvtmtn0+EP+3TE2WQMyJD0F6ayCORkE9AZ1fqWGq1T63x5T5RskzVGYin5QvA6Po/215Wri
D6+mKCWYGU7gHcFOevZDYmkxCiMBVcToGL1PK5c2pD+tMVRFCkrl8hycv871j4cO2vb0nzpvL9vl
VPbACyxN7TniZAFyQS27WLV+UrMc/klPAak/XTx5f2RC7HDC5P4E1sGl+5FEJfoMtsYnXe2nFLtS
cInEqQWutxZ3wa6p33BaSKslnaynybDxucpy9/CvpHb+TLRdU8j02OTNw6aicFya3hgifZhPK1u9
kRrYP7XJJu9OqT3xzsH2MuiugSeidYT2649zmGoTX63lKPWAoRkHj83Akk5kuUkIT0XXG0caHT7h
2T7DGZSm7cE9AopVJQ1b0cpkDOD4uh8L8uhK5ZLJWn69HGHzQV2r6JJMuSOX16ntXIGsmEL3YGct
i4xHYIJppMNq9SkgIO9PZGW9GTs6P7elhl1bUi12y58vGWKp/IALkiudPStdGH0RiCbN2C2GZV/n
qFUu1wFRPxvcDvLOk3b17+2mPdtHfGUz1ULpT9CNxfQXurZmf5oI9Aob+ySjoaDCX35nZiOSLGw9
LGnYkA8mFggdDmck3fZepGLFbiLKHzkQanohQjLDopVqFF3J4SfmxCnWc7jZi/Nu3wFNv9LlM/Si
jUEc7gIGGyYJu6EHn5OPVyrctFJX12MnC24dRxbMfStKoHrNdDnMVHzp4CO6R8hXYUZjVss1Wfeb
vpxYgZNSaDfS/ZvDBA5VZq+QATPDW3WF18TOxc4HC8k3+1aHE/6YoFlOfMIiQUfSsOmGt4k4duZs
h7zolS2gGfWWMdytedo5r6AdxHIcI6rVK9poJV+6Pyoa66inbmQgphYSu09Ia5hxocNmFgOxo5kO
80XKzKTOHEAKz3mWyiWet66kgp9pcNICs1TnuEkn6lUrKumJoxGZO3iuzAg4Bly2KaBxqgHvebsy
Dw9X+Bdse+ycnyIIPuLuqalI7XiV4EHAGYvkPnqzciJFI1P2douDsPEo84J8JCwlPvrRCFv2WQcs
8+Sc5qINmo9LreChQobpWOZJofqQzu/fGxhujbAc+AEU4qmfkzhVSqCmyxZEVxnRTKFAWxaG/Zi/
DWENKb1eKU8Ecg5DtwWtubT9bKXMt/gygf+pMRYQ5YYgNUTLMECslLzedrw7iF4crokOaNdfTgnw
s3YlqC8rcCijlNd6rH/4yW9ZYs5vXJwonA6bf9Y+uNDy6g+0W+KfasA/23hjdx3dhseUq/NXLR4J
2dp+jbqHe0bfe95EEHIXr+t/3LbNg/DFSi8sH9JSay1+n4DA18RT99gWOeIC7bzP55Ad9bn5L8Ts
aRkdJT5LzoxtGsvJ873wGdwIFGa8b0TlsyAf9brvrUp8vkp+33udHjVMzQ6pXHmohYzA+1U7Dp7R
Df9qqaATcmqreK5RwPqFbaxSC8bKf4UKFx7BQ2qMh9SSi6bgifESX8WqS2NbyXCQx23ae5HIOsxM
lm+CT10cWLWCyLYMmPkI+ASHq+2s2DsXFh655Qv3xE1f4sgxVyhevHcGOnr69i+iTk+TPCJMcYG5
ZEz87m+8dYcIxnUR8Sv3jElgMoZpxQ7SiLvBVDTmTpM/FKACehZvAn1Vbnx2Tkn4v+AUSHr8O7Tu
mZq/0mYQDAcx+6vqJLw7moqyrOz279Tj+TXQXlb3DOHmf2UJt3T5qLPoZyHzvEJmVBOnthR9zO6R
ciIuXcILT4KKsFc6S3smbwVQIV7/BqejOYKUiDve6nOlW4KP1QhPz2IPX82DIZcWIh//dsJqGeCc
bB6DM9EvLa95LS2GO5oZt69xvChIuTyU9IIFa3FkhORH/2Hpg/LwG+HBEntHDc2MrM1UHs1GPK/t
ed5LLlVkGK3FjnPwiDYfbdFjQJ/A8bkoO9t52zzzRC06LJzXimLGO9keKiMAoT9K/mVdzc9H1rwF
dk/64FT3zWf2lwMl34JzBFX1sbm+kevqWCwQxzb9cxT8LS5kI0KKwGTGsIzqZeofwZ/hPrjWlsCJ
guYDDdy38KUG9DwMyk4FuORYI1btyb+cURSmG/F2RyMmGTdgpeWI8L7GHC3UEJ+Xa3I2dnqlowFi
xG5ekmAFp9BiIWhRna5DMuBoXmTmmKtz5NR7o0Gakqwct2FNJjBSn5B2HRtr8hcmtWawM0M3Q+YQ
MrXchASWWFXvtR3EFMZNmbFLugDG38x86+OGjSeGSweywYHVh7Oh44s1/p81Hl79U8hAPEg6o1p3
qFvC2l9++EPaMedc/v4XXH4GWFD1xqgRbbvCd25UIqpz5HSj9t60mxh+XFcCdwfSxQQ4JKzg5BX3
ErZENNRmRzm80VL0KfT6BetnqbXxoWeprXlTNuNz6O8mNpEuvf1D10FzOsRWKN0U2E2Hd8rAcsYi
wfJnjw+EjYluCRzbj+0FTyJD7+ie4rELfQZZUOIB/dQxJJo+DXk2areMTpIPFwEGUju8J9O9lo1z
HyKSSK3Tg32ZGjcrHjPEsS7n+iSVc1qNIO5oUOoWOrYZNhNA7cWLEuiBzA2r0CVP1Dr+ktQo9Ssq
lp1RRIqLLtS/OOmqdTzTjrxRcN3Q2i3zp/Eyb6sZhsblrI0vYa8iyDmA2u291l6okDro5WxJ4DlE
Pv5wcMIEV4MDWHejQ0HV8SKHblQ+YnNKCdzfo6RZ1LNDkxoF77bP569qNUDUnztGafJrBtCiOVOB
NC1EVvhMGtn6Vfvq0MYWMPjgCDP2iQ7r2XFY0Izc8aXKhjGd/Ca9UBn/DNiL6Cd7pOi4iLttv2ft
bmO8Sdhmn2OB5Jkrlet/3xgf015K55F8ZCq481LJb4R/CFk1+T4ns8zXtiDnR13DM6VDj7o9NGUj
2Qmb9fZMe9BQZ7AILQ1FA9BOws6u4CIxHge1+tByIZVxCZxx91zPdqXYKvMy5BjdspKbnEve34Sr
jEHSinbDVO+lpOWPppWePM2zGNx145iG19LnrQITQvj3CNiHbuoeaC31lgG3paYx4HUd5yLR5QWp
HtSz1vjO6fPKGfU4rljmbCPTCkUfmGkSdRo97UOz0ZflLZcvXPMNYYGEoL/AnG9PYTeKuG6cLD4a
UbioH2+soNAM65DkNosv+TldFkSif9fsVhkFi3zdvNfJZCL2C+KMVHPgqKz4giCAXjMy2wNgDfJh
FtP5igIhTby9s5je4CH8IxRiwfzQrgdL7r02Kh/kWRYXychh9PZ2GUQ1QqstCn6QqMFnRJzRcaJ1
X23HcudvSoZ6Z8Fc2q4VACBQClNSL20CKhUojSUP1eN98Six89+tK1syM6PUrf0+JyaI+YUnAEcc
x8sNGvn2gjn1Y8rEJNItiGdPIZcA8jr/Q88NwJSfopSuu8WHRHKmcnKk9NwVClrIeCBrDVSlrlT+
gXp1DUuoYoe2whODt/URNRvBtmFqJamfJ4RJ7msnYREJ0y/uQ2R5LT0uxlYol08mH+hvxp6kvv4z
e8yVjRSgHW+5YFASdvy9K3KhOXZumhl1LOxX9Vq3kF9JFRwyreuBqHZLTd6UjZKB4LTWfsg1Dp+E
ZXKZ/9OIDi8wx3s9hL8ot42a325oZRMOqe4cbpDt6gsn+HOKf01jRfijqiYyngD9c/crpdaIyG4Y
2F5poigV/I+VPbmSjJBpBpTHMGMagCd4NGGR8G5v+vT9g8hEehVFEK/v8Nf10agvdf3f83f1MzPJ
Bz1S76FupcXTjj8cfju+8eGbRkZWo4MJasLnYOqV2qnLJrCr836ONjD0eZwUvKX1NT5EPaZ9ltvp
HlNDMi6iAs2KtBXddn4RwPCX8GC9IPGEPDz1WwWQIlhIoByNliPrFtpvNvQClRT6eW7QCP8zdi4C
HP1dfCfMBBsC+AEOd8lJrwTiZzgaq/aPPGTTbKSfJrdiTJ8J7ga8Vl3I1QjEHCNNN1RfFK07vTeH
Xcx0RKMAaITjp5XuRU/HQxJ+3o6gEyHyt3reP2haKpg+NmGZltC4wZuwFGq0kmTHklfQ9KwnaXJg
hO1ouB+vIETNcbqd4YfyNE24nWjKWM48Bwm+OOGEdj5RRhpagjTytmmPjTYy+bA3ShiU6ZNUtzYb
3EtgjeXYzd2WJGrmoqVwzSfPfdIv2lFgRYZvKm6ctyTKUHlHr6+c29nPxJbjD6qZAp3pRt0j5I+1
y3HqShl2R0EsibNioRQbrdxkpva1Sf5Crayz8diTs1W1bMX3JDu6hkigqNh35BJIeJld+DQRdkH2
y5Dohu2/uFNHLkj+K9QlpPgPMCey/7iyhaO6YoQDjrcOa9wzdvrKuElnyWjtqq1A6HmwwEJicLp/
3oM+p+tVrEAnB9dOiqf0M5+LOtTLBZ9qVjw5Zxjmi8/OjgkPVlWDHOYvoovr3/yifav6ah4O2zPC
EeWnxBS3hKHudwTjoBvr3KYVeB4liLeAdsjhBopYq0Bht6SMS/mTeSb9g71jIeVvZCvm6Bpur5cU
SlB9DuZv8aR35mc4sGtW+Il7Z+VFlXdsxj06ERcVXnXoTWfvRMIR/mTenI7iOluJ5+0RnUlrhqAO
QBekrX7R8NTfR3Yykg6CvOsC9YyQN1P1UpPNDlG0g10S6+7RKX9yvj79Tl+1o2gBFyJLWjN17ISS
Hd/QZVoEGbNoaAw0lfjbFYxtZQjILLDnKgiqrFvu0F55VKDF19eDGxbi/oMRXZdaclZtCCrAvgF8
LIkOyfFds/ncfVMjM3zq+Dmg1Ra0L2vzfD6kTJI8VNItyQ/1qWqGsdfSdiKiPlX9KWmKsia23uJK
HTs8EeQCn7/AoY2BfiAYYlUSB+V1wHHF4HaE6HrowVCdbpN97kUsfa2ONSKHhuVI1rxJ39lGPkrk
8peh0yc2ThP5ZlJDK+MzJN2+btKdo+GLVMgL9rQCNx7CrY0U3XVSsNll5KPMuLxdM6+wI9Mfzmyz
7QYEoy4Yi4hec2liE9GbtHUVL7M/UUNedOXxG7ohK3gp+gf4QwR9ckwOlT/QIlUtiROxcrI6Y/KN
pgu1HJil8xMWd3eXDqZak6XRUbZc4c10iih3lqMUT1w7hA7nWL+O7qeP6dN+lWNw/ltuiMa5QUN8
hNNpzoVIsKQQyDqDY8PSntmyPMicKNtXh/jidEwj7zirQgybur+WhJAOGUvFFo3ApnpUX5IRg1w5
CEO6UcyNaioDpdc7PXvhSy5h1/olG1hp6KQg1jeGE08ZXQ1Db50FWt65GBLEJnv6HifxM3lia4t1
fKcHIyYOUQepq4punHBHnsN2dfBQ2E+MSaX5JlXyJOEyKkiOSOk1bs+/Rqgk0ZY7nU1STDM0zUhk
YcaqiZGYEoL00aU1yHqdmANPUHQTbh9WxzKUpgzXn4ZiZnOmQyjZ58x966QE8rOCpN5h56HjmnNG
4MM24JYEYEBNYOjoTYfUnhNnxv4TIEhuBM22i0Ytfy/ORsdxEZm88grePOLQQnqFNYq04sIgNbnk
GBhZ3HIs8lybmsukN7S9JImDThMOK4rFv/ZT2edWw4mcaPERijdrfEsJZNh13e67mMXq+ecvs2S9
v8l69c6V7iAZfCRgYTvDAEVzzXghjGYqi11UM5gVtvMhopVA+1nPLxq0NNk/C8avbkQOMkRRRHZt
FObUxxQEIIhdfGNqxbs/59e3ELGst2gBKc+bzbbZWd693j0JBPqQnI4QZrseLb3xQX1/8xkd75tR
1yznHK4SAkcdGps6ZRNEYlMCB95XSZLjMpMfaRL60NdeohHFGE1q7X8eO/NT4sC0zalG9neTuRN6
oGdMOUIWSk9wcbLZsH49dWo3xULhmomIljQtkwPcol/SHcWL5T0mxPmBe2+pT9CW51UXlRxnxzSv
g0MV4OzWwzi/KK/DaCW9TQndQEGbxFnRBzdsMZjsE9auZmj4q3lxmEAlgREjL2j+2XIXkexX8Uyy
OcNiRUQylNFN0Lqp0747xT8xZsmK0u+p15XCqCzhSJy/SZtA1GQeIBjmmFNPt/niI5W+G1dmNN/q
dPIHcsTQY0NSDDdiN9rFchCRITpiRD8jXiJOMUcrJ1Sh67h/kX3dtGYgY6Bm8oWUYGhlwgpYSQvG
6d6AxN9BjypF8DJv0DaFjqG7MZgqGNhplOtOsTqI4H6zFuST5rfYUdsJCnjYyqhe2x+mVYmLDX4U
pIR2PV/9rwTn3yu3lQ3f73AUOv0JbNEaY7SZvcjLdrjGA7ySCZx9KpxA0hK+bRGnlbo3RTGjshHI
ZLoLMFVVIN9LEMcrObMGM4Q+ROi62E504VIQojedbWy1Z58FXJgmTFoTUYT2bM3kEx+DGLfVBQNI
03UcSAAVIeF6oUqmJMb1R5576VsL0j7ygCKQIoytgofHZnQTn7arvhThFDgRc9G6k7MI1QSFV+Y5
8R6rWLwKDujuF1X0O+s4ng==
`protect end_protected

