

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gxJVQBcSQzsbwH1GLrg1ZESzDvrkikrA6vdLpp95ue41M0lmLElFgzzCnPkJPvxfP02JEfCkzu1s
pXyOx1+/ZQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
as6UL1EJsW9MY/SAJjdc4y/0ZbchfPWRZ1fO8sgcSvmzT8PhDxHiE2Qv094M2Mf5UxTO1pmguf74
HRrcuhkl5xTcz3SUgEh1WqTgvNR8v3I22HLFetAdFeAfwtFZ8WvCSLor3Yg5WhjacxKzsx/R+B3A
Ic1e9ERorPLK+2OWDXk=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VKtFT/ad0mndSTNYku9P/p8pTsvri9shyNk13WEjbKiIq+gQoaEMBYqKlUj1txesDW5BSN/vb2L8
WcR0ho1RI1AGo8y9tYmqORrdmk40Vs1+gqMQCfIiZwlKBZmVSoyHFg/uvBbeY40omXist3OrVmLk
ek7TtttpRm83fmMK7OGVEehvqtEULYY3DOqBcu2re7sG7LxKpszndoH7kfBnWA+R4Uc33vWeadnd
g6Oz3503o4HZjTYzqaI83vGJuKxDWF5lpNA6grtaK6MLeulhLJkFI34NJnCbFwlIH0j/a6X/NOK9
kE/9xzaRMrt2DXPz06r1p9zWXUaXULkLZNJGCQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fSxesrZXgYAQp6z3s+Mn8TPb3bLkqza8nC5XgxzWq/mXl1dMa5Ml2g5M80mUOlkXRmUOZymc+Bc4
WM2y1HxgX5+JsAIjs1wpPrFSHzjHRcHcvowsTXhTMQ12m5t3+UzDaDcRPweSUjf18fqi6cqE3nVU
Sfah17SHXQ+D8FjN0Ig=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Pw16GfE5lmct+1yHq5aabqWplAJ9NyQFSmc7ZK86jiJfkiQiewcVOFWOaoYaAbWH8NvRlUTWxPDY
IJZow2AxlsHQYg/BVCCfi6Nou6nItiOvPTdaycyuC2yVki71gI8y/Hb3VqhrwCJyz+gO8RezkRKT
K7icG5iNkHF95Ybco1baJF1EsxTsjmFbbCqBjLdWPS+4hZQmoZ3Ifbb7SnBR+mh541FCQTCGTC2j
d/LaIIFECqkijQ+ZFSd6r4keOeZDRlAd90xaWc9YbUz8EcXsrFGvk0cfiELaenio+xWCzcCA4xZj
1RA4VErN6S6k0GdYguQHKTjRx2AHdBSjKkPAZg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8720)
`protect data_block
vB6MA/ATm8/E+Sp3xOHp091V1w00VGLw9MJG5AQBxw66ogRajUy6/R3IAOgIPLnA2+Ueb+//G8dZ
7dZgZpGXLWzhsuivn/52dr1KqHHZyH9Z2UrvKpPbeGNxTx8aQ1T8/UvmhoLWtaGJddslWZzUBo1M
pPRy9UwoWrmPlTz88eWyZbN0zmpefxg6OydL7A8NV4u6D8VP/n/GgJWuZmC2FYd95GxXx4+NpEbg
Mez1UvsYO5LVqMUwe2QhZ0i3fe+Yh1lh0qfrMi6qcL7OA4aazg1ynBZhNrUYDzt+q99Sc/RvthSQ
gS6F4dnX3ncI1vilFILat6DudHJw2uhos0/Lie4gTEhdhb/zbDusT3kbWVrRl7oYAehuk+0iT5/F
OHFfReNi5u4q4n7+6L9NQFtqfkbeTXura2dA99FMv+ACE7z7KGSZn1lfD/DEPsitiI8lpZeKCH4q
qEZu1eUDPt9okQe3kSJcATTNzpWlYTqODBvuHnL8LpFQtv/xZDx+CyFmS8KkwJBrQ7m+S4qJuvho
gPHVuVzEt+mqfxRcHFTR63ad4TSGJ0M9nOo54VvvRA4QdHguunQzxaJgwnkbsuMkoKQ7/5tHVh4v
Iz6Q0+Z/hdYx1TOOKa0DtA/BZiXpFQDGO/kdXxDF2gJsjBmFnd39fUrdywjftDhlxKaGGwt3AMyy
UWOg4Qs4qfOGrxZQH2NG2w1cplNcLi9bO6C1tUJTVJrkdcpEq3nmHNucJ+tYt8MrL1n9aegsjCWJ
lVMr2MFW+XpBFXL9OGJrjNCP3rX8zWPko6FFaWYMhWwMYBddit618X6RtkvrkCqb+ET/AQaGuK0H
V2xEdtPeMAL+4kvv+mWmM9+/XVYeM2T4BzF+uDkevP9PQRdCSCm2+sI9LwW4UqZjfdBnEUoJkQoG
H0ZDxTpEwyAEo/MIi5KLEyb1gT8ghb/Jig1wkJGItF53o9VinXCOSelAugiukzkdw1qfVWvn9N7o
YSrKqZXRFAzqUVT1BE7Lc+44yojXz90Qv8PJWvHBm6FQDLYFXKPf0BG6yA4Z05Fhlp3w7JkjKVVK
c2Z7oKwgfAf5BzjmiHLUXbLI6n1/bMFNStKVcKXU7UEVuc8153uCYUubXbl1T16XJ5Wc6XIvBFaB
FbfX0Os1NUJv3siWy7NjhKVEcYqo22x0oc/AvaPFvcwNyVr9okyaC32/8jtLDy/ObcGeN+K41+i8
w7ZSpoMomBT08Hb8TGOL0ZQjqNvWSa//hfNR4JzRZ4VAqRH1h/XT7PJMHu1TSLxK77NY4IyJYX97
8+gEUniSv6oPF8sb/BGo8LI3ZAYj55gyGPCM42PCw+8b4qYlW94WdLQpug0Zd1zGi2aeH7seF4US
eKfoHt5DmyOIOrl78UJwxQEABUhz2ViELhoU5c1pyGhflKt3Jq8jm78b/XckOFM4/KlNIrShqjEB
b+rwJyV23S4eMqw/LG9OmejyeySlGQlcTRgni7o4JjbX5y0B5mZor0UWyceA4kgaxHgA5dR+NIAj
HJxf2Zy8aERdeJDaqbtzuU9hC8oqwDz5mTe5jX18tylffVmAeA8Ky0yKFnNUumk4fjxYOLWEvnjo
1xf/k6cescGy45Ji96qsx+fZps66+Top0kQjVZmu1UbDzFPyNusAyHz/bklaoiKA5XibUjPT2ULj
7hm58GBoFpUU5eo5bNVvhJ8LyfUj+o+nGGFYGwp5SBgjsLKnAki2vwZ8XLtzKaGZqNMoApxALRqT
F9J9WjDKYx+zborYRZtGgll8HxqpEYJ/QBSoLZUAeEj8slzhkYUcMaDdYvzNrJVtGS1X7KQ4dr99
4kQgsaQ4dWbEcZa2o+Ik7oxJnQvixDI3f0XLiPpyr5NXCdm4UPZqDaAfywuDG0ch9F4eMKPSLepi
vfk+rkSJcDJL48cF0DjUouccDBuMZ01gttDtWgv4L8gKpDBJo1ZKXkjnFMOV+qiBP7U8ROtXqAuq
YNT6wwr6PjAfj1Lju2V8FXYNGfjKcT1swiETCmj2QxIhvkCk223hf14KMKC+hx2O+BDtsu9LRdmB
cqK7irff0shpul1JlWbY4B1g3CSYkF1b8sCwDV4Fa4g5oj5BO6OdRcCrCZ0Pl/dl0Njvdz87aSne
cstUZriAHhbfAMLjYyeyw3e2oMAIGNX1T4MWUEGasnvVhk7xn50d8IEOpEfimu5nK6vyIvE5s+1S
0JmW5jIo/P5AX/2+6bynRsDqMXs7jPlzxGKjTmKxEg8ZntbICXjJW+F6bXpruLo3EjsBRpyJWh+U
pNYHiNHLG2WteDfXKP2j+GZVzLJI9wUMAD5i5jueuuS7+PrPV9Iq/kFsJ5XenSU3nHPnRnuQN8kR
ijoS2IsB9+34Ys6bhXzatsSKzn8jz1vpGlFN/M1jHiLycoiTH1QVic0gWmK1/hvB/5hKFmfeDBUO
ytxtkd9A+2tICpeUO3ILPTOONLazXyWpP6ifFOuAFb/cnZZf8vKkSTBCUdUUAbKtIcD+7blAu6JV
L2BzxOL6ge5cxaihWILKrAA/9Lt6/q0W1PtFaV2BzCysyrhTSbSfMYjJi1eBmaahfHnFIXeSy6Y8
3x4TxQm6AKrey+llfwlRTjc4dc1SuWNkZxZbUzmT3E0s/a52QLctWY6uL+/Ifhaj4orRc+UnEzjr
cf8VoftcNQW036dGzAo3Qiw0izvwxNm7oS9X/lsEYyYyqZ4kMmDv6Q6Lf5AK+xKSR+rcNxX6a1oI
+Am0rrW0tq2iWLswyRF+JKw5xNxA2FvfY03JF6MKabXvBkRempV78Jx9ZSR28dgH+brCGs4/ZEAz
uyj+qBd+fnMfoCcNNNutlWCxwZtTYU3KuhIhid592eXnQvm3BRGMGmwqBiViRomGahUy4m7MxnqZ
urQBYgb+4Pb9lb8fX7RemSCgy7HMrNzVH1z8D2qVm1ESQX37i7dQx8BttiyPSMjfpz858sNDCJEL
1NHkB6nubKs/XC4UmSd8ZqmmEboSr4uPLjixyPtacy0B8F9cOxqKjmb1qKAp0N9SAwrJL/kMjUHc
amxnQ7FeOX/VZhmzuHAtf2M4filzNAaoaKtXLsGP8HgY7Ga9LfWQiFi+QGgvv/C12MSi8NNjbpSp
6mmpXtUz14c7gpmkUX+BGn2Gok/lNMhvW5IMlvAtSu2ZwzzmlL4qvn8aLjxml9MKwIq69BoxCtGD
bdQaar7XRXELLSqh8dyTu7dY/5FyNjMKeT8/UmOhrwZhVDrrW1ysvt0rftqbzb9ad6ZC1/noRABm
gzQU/7FfOjKyUSpEXncpDjypW1gKiYOuk7SlntRbgnNGVAczkKaU31QVOA9wRgIUAMthlmCLZB00
stV7WbPR0Uewmq/wBxEBsNQrZklX1PpBLYhczh3Jgu6I0UG+RUCkrbUYf97EgBQHp9ejuhb+6HZe
aJPl7xUaf8SgO3V9TM9fqSYDI88ETFgDs2tF1ZRszuHKEO0lm6khBrkpO9yF3Lw8AkHWOR+i0UTk
hSGAz1ukuz4IW0USXU1wOy8rH5vZXOhY3PhEQSwStXSpq+JjyDVQACe2kkkkmbtbwbFUzPqlc7L0
Ht9zKRplDcXRYx8QNmYQMiA0saWNC+Gsr/7pPfu/xcWz3w1DlBjFdEVeH08ETk+Fc4+cqCNL6gT/
FP/D7j0BeZsPLdWk3GnPYSjEVjFsP16aKcJWaWO+xPG2I/qBnE4lz8daQ+PXU2aQwBu9s7VKfYVq
tZYdiKRZLq/6PzOvG+CZxHEfOYaOtLXw5xSsjL0aOB113N31xKxkkVgU3kVvEmWV/+Weve5gTRwQ
L2qHm+EHOX7DccUji6LO1pWLpHlogZK781czmBVS6AiwbRIT1ehTs3nZYidwUUcKK/1ayul/yfIo
scKGMbK9hLOqWjNJrVdfiGrv2jzA+tkE30s+SXdHHl4n4InAg0RGaSA7GvHJoaVAbJPcpGKFA82u
fzOTcShejVf/IJHiEbFzQNn4VJXkNdRITaPE4wIR3FNHyldLakAaeQd8JhiHmO2WbdFpAxv6D+z8
OP8xROKUfMA9Ol6Ck8tb3zLK3aJzNPNNuybpFrQX6+/Nq3QRNXMM2g6dgyaK0WfdrtuNfO8XFPqS
LjTFwrUGY/fHtPzyq0CDlQkEBI9J0jJBxerfjlNwMAVDvdYgLneXAh1Nm5CgO8hoyLBYQv/cAhpD
SeclGNuDG06+FChTtTqtg05dKFUYB5nN56nAA2ibwUgB+8bbF7Dpr/C+3wlH29iX6q8nlQjFoUAw
EEY9zrABlC/1kLieYj7cQYvThPdLMJgxqv3L/LJMbECHTXcX/7WyKESzgK1XUzNbgyPfJx+7Y7YN
rH3KVXuBW7Aifkv7eKNOba1Zg0gRixEvJvjdrE4gDNBGStp/iCH7i/Gd8rHx1thmB8aJqyTpAreD
aK6Sho70V7eutpZTebiI7L7jZeafDdhOLILF3yY0YYnROYOooO9zjwvTNQjZpHooZUhVRnQmevZw
weRS1YoNnSww4pnBnN5NKGmIf1VfSQ/qjCZzfK3aKgqSDPox8i1PlXjEJm8Vhf1jLXX2z9Le84au
PsSj+wI/mxOSqeuKtfGu9xvNxGN8RKaInQyf3tDHGQMYEBz+cMC2LSnPnCVi1MlqEV9/vjoggPxt
uhZfp+N5C2ACsTjH6083xiQclLWtXXto3b8G5+7WgDNWFlVJBWB2FXDa7sfGxXySKBBDSi4hFlPm
vVQHLF+398ucTo0hjwMcRtKZlLne5rrSrJopNBzkAe7VtaO1wPlf0w1IP8nWRiBrDesKEa8uhThO
Fxieo9x3VcsWjKoR6E5x5WLdblyPWt5mHiJK6KTarFZMtLySGT3Bg9CoS+sZHnCgmYXTVcZonVRs
HY5ZqCVPhdO/M2EEo6HHLMuB6Y23LJArMLnYI0gHS9MPrc4t9BRQBXxuDlpBrAi4/PTGNr7wE58M
ssCv4UdJpi7UR3PGY0wZfa7c+qKiWUM+Bw29DVR26OvCqFpDg812EQHNjbpXDZd9JfO3Wqd649bc
r5Tr/v1mixQtOK36vD/sr+aWVWsx81CHU0QvRvJ/daVyFE1eNbV575b8sviA1D7dzOywSzRAmDrW
sRPxZjZCQl6Lg8aR5gj5TpNyzwGAr95kRKv9icdfC33RScGVqvQ4dhimzk5nYo+boipkPqQUBBvA
odcjhTeHRMABJT7yF/QKORBCRUt/LEfpQqFMCAv3k6plGNU+a39QG5F8rgklbRg5VxlZfJdM8aZy
PE5y3uVo0ltFz6dpTv2d4RVwtzZB1/Bd2enijeGNhCJHpUZKRhUhKWVIKc1U14V9fvQGmC9TaRpR
z2FjeNE8GIJjt80HFFgYHwJx5c7a+1IUQjlv0kxmOaFLqn0ZzZxKD9RXi9CSoLlceSbIYll/2MZ9
qwWYZQI6sHuCit+fbOOY+G4bedXgUEJXESIrIr5XKVDtApkGHpMS12s5PQa0GzU6RCyiyoFZiMqk
oRf0uT0wY2TSxyW0zb5ZHbnZMk4FGSohTFUWNqbaW1iVp1jK+C7KCSNMXjTG6zHWweK6W29/RPty
Jw8KE96caOASnVxQeYqb++zPIEz+mouUJwW9H5squxwgHfCS6pzY1COQJwv/H6pk/OKFXOU13NyK
7AQDXLyJxO5gQM3hbyJV6L4REXwIh8gRgm9PYQBZHhiftVo65aihbB86yHV9AOyEKWjgPzUWP6ys
TAWz1Rk1trX+6Ps5sVRVEPPHdTsO0Y8/pKjlhiOCE35drFi3Z72P2p0G0teu5QoWJd04MFT/oqI3
hpvX6lXjuNej6864MEGwEBInkA8BOAGFpa1AsoDXVycErUsdJToWKmK7kGi3YjCWLvLxBcmGmGv7
cNJqtn+Mqwo0vzLpAcBxYF9CevXb/BA3Sn6HNNYolWuKf9/G5BVWBtNyuajHoFEYfvdCmf+3DRYC
JSyQb+cV20VB7kiteGBkMv5LfVH4V5SZssLSdjdp00IMxKiWqpEPTRJOGdbTLGky/h0EXIJwI73X
7kzeJyQZe0XNDxbAGhVToipJCAPJeC9+e8htF7YK+oOSJYOKD2+I0tNnUHwoaeC2pQ9cITXxYT+4
bDEEmfLdcAeZqwJtGc4AzuqHoxtnO15FrV53OIhUJ45+dx4HNTMvsWHv3ot+Hd8HujUiEbyCF+/N
yrpQ4oeJG9oUJzfE5mRk1ZLSXe94j61joI04LCGB8VQecr5sgUdYTjF71fprkpBYQTMqF8PIs2Fo
fC1PXSxDL76hoIFIJU2Ea3ruxSYr2gJmRqpLQ8Ud7wA8o0hev8Ln4/1ACqq+iygCmE+gHYdEqkRH
gH/IF0Um1SS5KNrNUKhwC3oISC81GLG8CFb3g/lF2ZERQRzjA/w9GT4CPsuf8F6OqM2LuGWpB5mQ
zNjxLdl/VuNCSfAQbOVUtlpszORPRXEXwRC5lxUz9VCfqOHlqhfMUp4nJvV6o3LzX2lZ+QXPBsDa
WI0B7o4rIJeGnV86qSFQ3Lh2/LWDIekJn5YmudcxwT+txLpxOKr2kZUOFfWYM6Ssa4eOaxFOHwic
7cXmG6IKMk8uwjXYNsc9VOLNFXlJu+TdhbO4GavHKyGjBAcNpghw+Rp0ojFoLHfv+GKgm8Jjhahg
bzeenahlFgfVKc1E4J4pH/Xg3HL2ZhKnvKti17dBNibNyaxAjrBT4qG15lBT+vf3xhqp1XZXVxmV
0/SEJOt9AkGadNa6jIJJtBsxFn0+6bpMVyzKTZJwNEBAnhOBd3Cja6ArW122VbjeQbkQ34AcAQCQ
IIUBkXfd3RmV2DLEarhjNkeaA/5JDqxS7dt2G8fbsMISdpCr9F2ccK79KNMxxem79ibtztsNca5f
FoK9n4YwzxszzQdjtNjYG4Y021sq4TRXxZ4yzxWr9E8abmD8HqGU0E9ZuXveRaSdsJIwbsvEnmcY
YLt4wqg8YhwbXnvTxQQBbZNzzpaHFWNc4BXNj23NZbhTNw0VrwHwL7hpMT7cQzoSQvcINuLrePYQ
lhUxaLz5sKPFD/RJO5g54T/up30m7ofwmhsUCrH6E5e9uk1bCmtsnXc7BG1FBAGlTcF9LaSuyxwU
tmj99LTT8rS629ptcLAbYOHGn623NYJTAnb0fG/PpUEaU2MciGVeYB/G8AQV5MNcyfz0oJk3ukJT
uQRUHALHzdl5Z7YBLnzKkGBDMa8bJs4kKNdNy27Tw6tqy7zUS2XJvDng6ka62Xhp7NZagS/yhTUP
8YLlOaA03BVgWXx7Qig5SSuxliQlhuKSYnNvqYQ6AQnsVYwOEkWXHMdhatw3fU8DhnSQapnj+Fes
kvHt5na9iYk42MQ1P3/JGtTnRVAbIwX6zJrFz+pjwz+mqZrRD8OgvGmksM5TZ+XLGIkntu+eGGEH
js34h9LQB5DK0o858i5W0ovyfzovBBCmwwIy5h/uqhJllzZqGqwYqnOdMaud0/8jYTQ5gfE5t/oZ
k6MvIsOHDCdH4t7IUWtsMs4Z1KXBluvLbOqITDamezX4iAB0sImWf62reTZ5iayfd41XLihtrxGL
dH210lKrFRX4KMLtpzyc2ot/GBQM4rHFDAbYsVOW59WENRQUy+T3FMyXEBHZG8hXf+gY0y1AwNdU
Mgx6zgTl+5nOvdxES2JzqZGPQD0ouTzwFj5PXOufPTTgnHv+sWs2mFcrB7MpX6pJvW1YrTgcegwx
zgIFzlnDZom9q+3CoNgsLz8V93UgrGjKsWJctGpUcdu7CyulgBwLkJ+C3YArVgegLWfOEyoIhsXx
2aTPntOAd2xdvR9fYLjeyJN0wnOQDsKwJf26kVGr8jk3dC1/uoJDzEP9/6L4rxpzWFrHK/6Fm4AD
EPGnXnRNwsswFT+XZv0jkf1641qpHWHwKXHcwI5yPO37Qmvqe2Xk4H9s1ueaUkcxwVUYox/A9ien
p5U1KM1d6h5rW1a29qu37twL39jF96UuJjufw4erz7Fq8aOwqnq1fQJ21h/MeHb9c0ZXEvMiVjY/
L+PD7yvs1+mWXNnXr+CI/KlGcToCfPVEP5pg06YjQTGiKRAHarqw6/AFDxOk6h1aMnBFL8UGyDra
PYQs1KsjnS9k+bhLdSZhwMBvPoFExE9KqFZpUuczX+2+3/PWGNtpUU0dGgn35GpzPNcr25PKuxWY
KTwXpW8QUo7MDG7KNfH0EVTYYkNJLPsaia17Bl5SByXcAX8ugpFnVp7RrdhHIotrbQDDy1vTkd8A
f/OyFSCHpnxkrdkQF6rnhBDcmqjwQTQFqznCQyunXFacyKV2d4c52LYxxM50GmFIJ66zQdRA7Wog
Af/KszwZXDJ9xQFmH3bz8hNnc1y5rztQhhpTg+6XYg1XTZhsBCtTV8eft/NgAag1aOE7nuM4Kd/3
U9ptct2Pul0E59/TNQc2XIkT6ITDDbiF3M4jRi1z75rCnBKUhrsWnVyktz5haWl40r7oXFoJcw4R
v6w6KMly9iFRqIW4kVdrntQSHkz9sKf7yqx8tYR9pGnbIunyT1V/C1y74zkA/Rrgw98L2jiXaUYQ
XGPhvlvSjXCZ7m+z2Q6Sho/f2A0+jFmKVXQMNpYTslObzh0UUV6HejY3E5PUMBGc5g1HSL4GExQC
x7DanB0JqKctBFYprhUCsIk7sH3SXVpfeMVDcrjRQJWwYugwr3ed3ceuBweU7NJk01AGS2dnYWAe
tNOk4RNOtzVtKEMngoKyU+gK8y/1wYBZPb/t/Te0LGlRGhsa8dDxPpz3pRFn8q9xWU9NbT69gVqY
DrEV0iLfmwN7LxKRhRDhu+D0utk5ZAPe0Ho1KhAOJzNhr15laAQBdfmw0KUSquVU1OYYc2CrQXue
1QP/yPfaTsRwZtSxkfA550TPPrJrukxZuRBs+dZrnA8L73RnyE7eDvDafGe7a44RfxW82SLVtdVW
YY+hw/Lk/B+6zsknRlmPBL6tevuG7QRsRpwQ+wAbOCV8HpMbo/Oky6mcIBapjo5L2PXzMZV2FMZ5
mSP1WvzNxREtRXgNS/NYeMQ0xlB/m27hCFyD3S+69FZPYC1zwZ9+Cv3W/2m5+26IxaZYmSnm6Rk7
SIjkuiFwJ7r51ULSYe+h6z1cW+ewUxOI4bONRL5i7o4+Ps8HDYuSWEjDIi+LkrAni0vhM6u2pZkI
pu3sgrEjN/8Anlj0jyChzJqAbuCRH7cJ5vFHBIXvqI55s4KI68jQCxb5G4IGzll0MTdjnN5GE8BQ
y6B944P0NYavRtmOMyTlDuVGICrxHbwizKiSVXgwUrZ/0QpR06Moz49Tv/zYETH/XI5pUz5xucO8
rDsln+CANUH9pTAkLF4zm03dx2ePRb67HhMM4XqpYciOf8QQwfrTP4wuz/7RAJ98F/b1tVe7ZKeH
o8hqh4P5/izxuidodkJHQeboIFhdSBTCJsc9NYdyyjEdl88yqUwWxvvmcWsFi9ljRDRmW/RbcoEo
aABVMpJlcwZQ0x4eiLz8Emz82rQrfa7BrhTHE3xQy05OSMwEI+r9aojWKKYZ7cH3IY5isZYMIJ6l
yk6EyFjEMk6AR6O1HulpiWB8GsIyZmaVL+Do4FDaV7oFStWWDUF8gLhjlmkzjf0zChvxHe1PqlQM
c6Swa+0nIx2wKVeUDzqmS0OqeiQE3dXZNJ3pwBbYrydQmuZq//S+KjdGi3sQ3gRfZ2AgrEPvsMyP
w6LwjE9eccAkuhCxDr6vJMlEHHC5wdtlbUH+jmhw8ZHrwhOR43jn0JgSRbjKYdd0ys23Kekjl1wR
90C7DEYsoW/8bKLwmg7Lb8GUl44f/v2gxWotRSsAlkKkJVmV1uGhHrrzK8/tqt1OUPyDKDZ9gM3U
/rX2zLkFfbhKOnWxEvPrCI0iM5iUva4Kdpt859YB2wudV76CFYqlrXYaPRHuRkscbKxTl72J8zL9
r9FxFHwi/G5pjxpaNeLXcsN/O/UVm5CK5ITjyuQMP5PZ2ZCA+fuVLKuVFZZGZz/2Ix5xa54UVAs/
KlwZLGadqEeMEcCAMoz8V1FyedywoIS4+/IqxLGNcyNCnfx8xSZZWYUOddpzxc7GiR0lLxqFAHzI
wYYdv1xMoR66mcrUcuOaq38jqxX7kqr9+yTErFCfY066rEVvCkdeeFaHjTUwsZaiJlr70Ys5wDsr
SoCjvRyC4+nGWRboazFcg/BzSrVzHmOMMUBhAVd/Wrbz0s+42K8M0lQ3T6V3vjvJCABZK0z1kbQ2
v+XYqNrY/O71LIxckl3yWqcGuaDm7kfmiyqV5mZmZp3WduKAqGf85BLwPRKfjrZt7JYOM1tIWAZ2
lzDTyMCMFFXeiD/+ApDAXAn6nqa5MWya4lnQxcbz43oQjvDzIL1QjvojjloVozRdHYX1r5aCyQJk
EITmSvvBfZQv+gnROYco/aW9x6BxuW6V7tozyuJM40Rq5Vp/e+1jquXy94WJbLV2GFBg1gKue4wj
QtiyJqntzxKKmWH1mHpZfQTvyfCj06RA2Xd0d02zylL7FOGr+byJF7No/Ts4aXOSTcwOfeSwMs9g
VYW6zf4qdMRhNWWLR4UOMotIF0DPX+5xRO+TizriW3X93I306YGWBSSs14iLpCmPosGaFHC1aCqR
3Noaa7QYQ3va6JbA3CPKHubrkVr38bezmkZeT3OhHWjW0OrzryUcoNCtYccv7Yd/1Y3jOCjEcxuU
vGlFplPQy9WInym1epgyfyDpcAhEqLVnJxN8ECoo9ad2wnl8F4jA+iJ6v0VArLTF+JtDSQCSmbBM
ex3N+8GWgobX7B/CWX45o8e2ap4o4WOw3Lj2Wx83ZWzXc2QSx1hfEJ8nrI5RaYVyhlgrCRqDg2Wr
SX3weac/nZvL63qFrAdqkDReueXDTuSP424UI0f/gzBUI4KAgtQU8gkQ7SXzKGaiRkn4qZ2ECx+W
q3mnriF0VqUVu1nQ3XjzYlT19jJ3GLf2id7YSbUz3wqDzL1uMnXEz8esV/+42ELzuZaCFskWAO4n
mgWzc0eVu7cQwG1PvY+zbJaKEg3R5om5QG50DsgqQx6b4AGeWJBsXnrmkdlMHMRz3C9CvJJgIRWt
CGXC84GN3mpbU/U2VSM8itd99E4w9bM2SA9cG6dNKVjiMG7MiNqLzrexL094Tr/mPOnIm8hdPAyM
tGXeoXT32BgFJ7BOk+BFv6KcADL+sluLm+sxaUvO8keMnKiUQOcyXONC9nMrpQqBGQRq1jG6mAJf
PqwUaSC/B1s0iKl+PH0xhs356DC1aXKd8syhSk6/QQsEBK6Ij9cOFVGwdsHAL27SykdZs1tT2ksf
VyMEsXLdGtkd73G5yJTcKktUkEgFWyv3HjUx1yymr+VxyUxesZoycgoeB9Wn3/izJHg3KcJaDEZp
f+caALq82YTIMQJjYKVs8HB28C6/0iVz1s1AzYofsBM7ZXcwb/DUw8VPinVXp+nywKH/yiGPdrjw
xUQKU7vzDjiTzoD/SrHhFcImcIxMMUCuWkg4hiarA3FHVpdVB9fMDYDGfMjjeOyzAyi3emNTYzHF
FmhJ52kQMrqm/NddxOv4d7rgD/K7OR4MySPl0ri/tB+5QXyQ/zlQjzfJ4DX2S1sgF4lLg7hqvKoe
HSgZ2S0bo9JfkasE+htZdxk8FDNsRwV4X9Q7c480KoUk0tRkBR5mZMlzO3XM9Tq6YsCKzjOgNNQ=
`protect end_protected

