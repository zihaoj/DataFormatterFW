------------------------------------------------------------------------------
-- PulsarII
------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

package FmcConstants is
  
  --################################################################################################################
  --########################## PARAMETER TO BE GENERATED by ../src/ software FROM here #############################
  --################################################################################################################
  -- number of lvds pairs between main FPGA and Mezzanine Cards
  constant lvds_pairs_for_rx_in_each_fpga : integer := 12;
  constant lvds_pairs_for_rx_in_each_mezzanine : integer :=24;
  constant total_low_pin_count_fmc : integer := 34;
  constant num_fpga_per_fmc  : integer := 2;
  constant num_fmc_per_board : integer := 4;
  constant num_fpga_on_board : integer := num_fpga_per_fmc*num_fmc_per_board;
  constant num_fmc_per_mainfpga : integer := 2;
  constant num_fpga_for_each_mainfpga : integer := num_fpga_per_fmc*num_fmc_per_mainfpga;
  constant width_of_decoded_word : integer := 32; -- DATA FORMAT DETERMINATION

  constant lvds_pairs_for_tx_in_each_fpga : integer := 3; 
  constant lvds_pairs_for_tx_in_each_mezzanine : integer :=lvds_pairs_for_tx_in_each_fpga*num_fpga_per_fmc;

  -- per clock means,
  -- sent data during one clock cycle
  constant data_width_in_each_clockcycle : integer :=8;
  constant ctrl_width_in_each_clockcycle : integer :=3; -- to be 2
  constant word_width_in_each_clockcycle : integer := data_width_in_each_clockcycle + ctrl_width_in_each_clockcycle;
  constant bitpos_in_txline_spy_freeze   : integer := 0;
  constant bitpos_in_txline_sct_hold     : integer := 1;
  constant bitpos_in_txline_pix_hold     : integer := 2;

  type lvds_pairs_for_each_fpga_t is array (0 to num_fpga_for_each_mainfpga-1)
    of std_logic_vector(lvds_pairs_for_rx_in_each_fpga-1 downto 0);
  type lvds_pairs_for_each_fmc_t is array (0 to num_fmc_per_mainfpga-1)
    of std_logic_vector(lvds_pairs_for_rx_in_each_mezzanine-1 downto 0);
  type rx_fmc_to_fpga_bit_mapping_array_t is array (0 to lvds_pairs_for_rx_in_each_fpga-1)
    of integer range 0 to total_low_pin_count_fmc-1;
  type data_type_for_imfpga_output_lanes_t is array (0 to num_fpga_for_each_mainfpga-1)
    of std_logic_vector(width_of_decoded_word-1 downto 0);
  type data_type_for_imfpga_input_lanes_t  is array (0 to num_fpga_for_each_mainfpga-1)
    of std_logic_vector(lvds_pairs_for_rx_in_each_fpga-1 downto 0);
  type data_type_for_imfpga_output_lanes_tx_t  is array (0 to num_fpga_for_each_mainfpga-1)
    of std_logic_vector(lvds_pairs_for_tx_in_each_fpga-1 downto 0);

  type data_type_for_fullwidth_data_from_imfpga_t  is array (0 to num_fpga_for_each_mainfpga-1)
    of std_logic_vector(2*lvds_pairs_for_rx_in_each_fpga-1 downto 0);

  type tx_fmc_to_fpga_bit_mapping_array_t is array (0 to lvds_pairs_for_tx_in_each_fpga-1)
    of integer range 0 to total_low_pin_count_fmc-1;

  -- ########################################################
  -- <config> From this line :: FROM FTK IM Schematics in LA pin count (0 - 33)
  -- ########################################################
  constant rx_fmc_to_fpga0_bit_mapping_in_all_FMC_LA_pin_count : rx_fmc_to_fpga_bit_mapping_array_t
    := (7, 8, 9, 11, 12, 13, 14, 15, 2, 3, 6, 10);
  constant rx_fmc_to_fpga1_bit_mapping_in_all_FMC_LA_pin_count : rx_fmc_to_fpga_bit_mapping_array_t
    := (29, 25, 22, 33, 26, 24, 28, 31, 19, 21, 27, 30);
  constant tx_fmc_to_fpga0_bit_mapping_in_all_FMC_LA_pin_count : tx_fmc_to_fpga_bit_mapping_array_t
    := (5, 0, 16);
  constant tx_fmc_to_fpga1_bit_mapping_in_all_FMC_LA_pin_count : tx_fmc_to_fpga_bit_mapping_array_t
    := (20, 18, 32);
  constant tx_clock_forward_bit_position_in_all_FMC_LA_pin_count : integer := 1;
  -- ########################################################
  -- <config> Until this line :: FROM FTK IM Schematics in LA pin count (0 - 33)
  -- ########################################################

  -- ########################################################
  -- <config> From this line :: FROM FTK IM Schematics
  -- NEEDED to encode the data to match the interface format (to divide the
  -- data into FPGA units)
  -- ########################################################
  constant rx_fmc_to_fpga0_bit_mapping : rx_fmc_to_fpga_bit_mapping_array_t
    := (0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11);
  constant rx_fmc_to_fpga1_bit_mapping : rx_fmc_to_fpga_bit_mapping_array_t
    := (12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23);
  constant tx_fmc_to_fpga0_bit_mapping : tx_fmc_to_fpga_bit_mapping_array_t
    := (0, 1, 2);
  constant tx_fmc_to_fpga1_bit_mapping : tx_fmc_to_fpga_bit_mapping_array_t
    := (3, 4, 5);
  -- ########################################################
  -- <config> Until this line :: FROM FTK IM Schematics
  -- ########################################################




  type fpga_to_data_bit_mapping_array_t is array (0 to data_width_in_each_clockcycle-1) of integer range 0 to 2*lvds_pairs_for_rx_in_each_fpga-1;
  type fpga_to_ctrl_bit_mapping_array_t is array (0 to ctrl_width_in_each_clockcycle-1) of integer range 0 to 2*lvds_pairs_for_rx_in_each_fpga-1;

  -- ########################################################
  -- <config> From this line :: FROM Bit assignment in FPGA logic NOTE
  -- total number of bit should be equarl to or less than 2*lvds_pairs_for_rx_in_each_fpga
  -- ########################################################
  constant detword_to_data_bit_mapping : fpga_to_data_bit_mapping_array_t := (0, 1, 2, 3, 4, 5, 6, 7);
  constant detword_to_ctrl_bit_mapping : fpga_to_ctrl_bit_mapping_array_t := (8, 9, 10);
  -- ########################################################
  -- <config> Until this line :: FROM Bit assignment in FPGA logic
  -- ########################################################


  -- ###############################################################################################
  type fpga_to_det_mapping_array_t is array (0 to word_width_in_each_clockcycle-1) of integer range 0 to 2*lvds_pairs_for_rx_in_each_fpga-1;

  -- ########################################################
  -- <config> From this line :: FTKIM-DF pin assignment
  -- ########################################################
  constant fpga_to_sctword_bit_mapping : fpga_to_det_mapping_array_t := (0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10);
  constant fpga_to_pixword_bit_mapping : fpga_to_det_mapping_array_t := (12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22);
  constant fpga_to_parity_sct_bit_mapping : integer :=11;
  constant fpga_to_parity_pix_bit_mapping : integer :=23;
  constant fpga_to_soft_reset0_bit_mapping : integer :=4;
  constant fpga_to_soft_reset1_bit_mapping : integer :=23;
  -- ########################################################
  -- <config> From this line :: FTKIM-DF pin assignment
  -- ########################################################

  -- ########################################################
  -- <config> From this line :: FROM IM - DF bit assignment
  -- ########################################################
  constant ctrl_invalid_word         : std_logic_vector(ctrl_width_in_each_clockcycle-1 downto 0) := "000";
  constant ctrl_first_byte_of_data   : std_logic_vector(ctrl_width_in_each_clockcycle-1 downto 0) := "110";
  constant ctrl_another_byte_of_data : std_logic_vector(ctrl_width_in_each_clockcycle-1 downto 0) := "010";
  constant ctrl_first_byte_of_ctrl   : std_logic_vector(ctrl_width_in_each_clockcycle-1 downto 0) := "111";
  constant ctrl_another_byte_of_ctrl : std_logic_vector(ctrl_width_in_each_clockcycle-1 downto 0) := "011";
  constant ctrl_idleword             : std_logic_vector(ctrl_width_in_each_clockcycle-1 downto 0) := "101";
  constant data_idleword             : std_logic_vector(data_width_in_each_clockcycle-1 downto 0) := "01010101";
  -- ########################################################
  -- <config> Until this line :: FROM IM - DF bit assignment
  -- ########################################################


  -- ########################################################
  -- <config> From this line :: FROM Pulsar IIb Schematics
  -- ########################################################
  constant swap_mask_fmc1 : std_logic_vector(total_low_pin_count_fmc-1 downto 0) :="0111111110101110101011010000000001";

  constant swap_mask_fmc2 : std_logic_vector(total_low_pin_count_fmc-1 downto 0) :="0000101000100000000100001000001010";
  constant swap_mask_fmc1_soft_reset0 : std_logic :='0';
  constant swap_mask_fmc2_soft_reset0 : std_logic :='0';
  constant swap_mask_fmc1_soft_reset1 : std_logic :='1';
  constant swap_mask_fmc2_soft_reset1 : std_logic :='1';

  -- ###############################################################################################
  constant number_of_banks_for_each_fpga : integer := 3;
  type bank_position_map_from_fmc_t is array(total_low_pin_count_fmc-1 downto 0) of integer;
  constant bank_position_fmc1 : bank_position_map_from_fmc_t := (2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 2, 0, 1, 1, 1, 1, 2, 0, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, 0, 0, 0);
  -- 0 for Bank17 / 1 for Bank19
  constant bank_position_fmc2 : bank_position_map_from_fmc_t := (2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 0, 0);
  -- ########################################################
  -- <config> Until this line :: FROM Pulsar IIb Schematics
  -- ########################################################


  constant swap_mask_tx_clk_forward : std_logic_vector(0 to num_fmc_per_mainfpga-1) :=
    (swap_mask_fmc1(tx_clock_forward_bit_position_in_all_FMC_LA_pin_count),
     swap_mask_fmc2(tx_clock_forward_bit_position_in_all_FMC_LA_pin_count)
     );



  -- ###############################################################################################
  constant swap_mask_fmc2_clk0 : std_logic := '0';
  constant swap_mask_fmc2_clk1 : std_logic := '0';

  constant swap_mask_fmc1_clk0 : std_logic := '0';
  constant swap_mask_fmc1_clk1 : std_logic := '0';
  --################################################################################################################
  --########################## PARAMETER TO BE GENERATED by ../src/ software UNTIL here ############################
  --################################################################################################################

  
  -- ###############################################################################################
  -- FPGA-by-FPGA (RX)
  -- ###############################################################################################
  impure function ExtractFMCRXVectorComponent_FMCToFPGA
    (info               : in std_logic_vector;
     bit_mapping_on_fmc : in rx_fmc_to_fpga_bit_mapping_array_t) return std_logic_vector;
  
  constant rx_swap_mask_fmc1_fpga0 : std_logic_vector(lvds_pairs_for_rx_in_each_fpga-1 downto 0)
    := ExtractFMCRXVectorComponent_FMCToFPGA(swap_mask_fmc1, rx_fmc_to_fpga0_bit_mapping_in_all_FMC_LA_pin_count);
  constant rx_swap_mask_fmc1_fpga1 : std_logic_vector(lvds_pairs_for_rx_in_each_fpga-1 downto 0)
    := ExtractFMCRXVectorComponent_FMCToFPGA(swap_mask_fmc1, rx_fmc_to_fpga1_bit_mapping_in_all_FMC_LA_pin_count);
  constant rx_swap_mask_fmc2_fpga0 : std_logic_vector(lvds_pairs_for_rx_in_each_fpga-1 downto 0)
    := ExtractFMCRXVectorComponent_FMCToFPGA(swap_mask_fmc2, rx_fmc_to_fpga0_bit_mapping_in_all_FMC_LA_pin_count);
  constant rx_swap_mask_fmc2_fpga1 : std_logic_vector(lvds_pairs_for_rx_in_each_fpga-1 downto 0)
    := ExtractFMCRXVectorComponent_FMCToFPGA(swap_mask_fmc2, rx_fmc_to_fpga1_bit_mapping_in_all_FMC_LA_pin_count);
  
  -- ###############################################################################################
  -- FPGA-by-FPGA (TX)
  -- ###############################################################################################
  impure function ExtractFMCTXVectorComponent_FMCToFPGA
    (info               : in std_logic_vector;
     bit_mapping_on_fmc : in tx_fmc_to_fpga_bit_mapping_array_t) return std_logic_vector;
  
  constant tx_swap_mask_fmc1_fpga0 : std_logic_vector(lvds_pairs_for_tx_in_each_fpga-1 downto 0)
    := ExtractFMCTXVectorComponent_FMCToFPGA(swap_mask_fmc1, tx_fmc_to_fpga0_bit_mapping_in_all_FMC_LA_pin_count);
  constant tx_swap_mask_fmc1_fpga1 : std_logic_vector(lvds_pairs_for_tx_in_each_fpga-1 downto 0)
    := ExtractFMCTXVectorComponent_FMCToFPGA(swap_mask_fmc1, tx_fmc_to_fpga1_bit_mapping_in_all_FMC_LA_pin_count);
  constant tx_swap_mask_fmc2_fpga0 : std_logic_vector(lvds_pairs_for_tx_in_each_fpga-1 downto 0)
    := ExtractFMCTXVectorComponent_FMCToFPGA(swap_mask_fmc2, tx_fmc_to_fpga0_bit_mapping_in_all_FMC_LA_pin_count);
  constant tx_swap_mask_fmc2_fpga1 : std_logic_vector(lvds_pairs_for_tx_in_each_fpga-1 downto 0)
    := ExtractFMCTXVectorComponent_FMCToFPGA(swap_mask_fmc2, tx_fmc_to_fpga1_bit_mapping_in_all_FMC_LA_pin_count);
  
  type bank_position_map_from_fpga_t is array (lvds_pairs_for_rx_in_each_fpga-1 downto 0) of integer;
  impure function ExtractFMCRXBankPosition_FMCToFPGA (info               : in bank_position_map_from_fmc_t;
                                                 bit_mapping_on_fmc : in rx_fmc_to_fpga_bit_mapping_array_t) return bank_position_map_from_fpga_t;
  constant bank_position_fmc1_fpga0 : bank_position_map_from_fpga_t
    := ExtractFMCRXBankPosition_FMCToFPGA(bank_position_fmc1, rx_fmc_to_fpga0_bit_mapping_in_all_FMC_LA_pin_count);
  constant bank_position_fmc1_fpga1 : bank_position_map_from_fpga_t
    := ExtractFMCRXBankPosition_FMCToFPGA(bank_position_fmc1, rx_fmc_to_fpga1_bit_mapping_in_all_FMC_LA_pin_count);
  constant bank_position_fmc2_fpga0 : bank_position_map_from_fpga_t
    := ExtractFMCRXBankPosition_FMCToFPGA(bank_position_fmc2, rx_fmc_to_fpga0_bit_mapping_in_all_FMC_LA_pin_count);
  constant bank_position_fmc2_fpga1 : bank_position_map_from_fpga_t
    := ExtractFMCRXBankPosition_FMCToFPGA(bank_position_fmc2, rx_fmc_to_fpga1_bit_mapping_in_all_FMC_LA_pin_count);
  
  constant swap_mask_clk : std_logic_vector(0 to num_fpga_for_each_mainfpga-1) :=
    (swap_mask_fmc1_clk0, swap_mask_fmc1_clk1, swap_mask_fmc2_clk0, swap_mask_fmc2_clk1);
  
  type map_fpga_to_rx_swap_mask_t is array (0 to num_fpga_for_each_mainfpga-1) of std_logic_vector(lvds_pairs_for_rx_in_each_fpga-1 downto 0);
  constant rx_swap_mask_channel_in_fpga : map_fpga_to_rx_swap_mask_t :=
    (rx_swap_mask_fmc1_fpga0, rx_swap_mask_fmc1_fpga1, rx_swap_mask_fmc2_fpga0, rx_swap_mask_fmc2_fpga1);
  
  type map_fpga_to_tx_swap_mask_t is array (0 to num_fpga_for_each_mainfpga-1) of std_logic_vector(lvds_pairs_for_tx_in_each_fpga-1 downto 0);
  constant tx_swap_mask_channel_in_fpga : map_fpga_to_tx_swap_mask_t :=
    (tx_swap_mask_fmc1_fpga0, tx_swap_mask_fmc1_fpga1, tx_swap_mask_fmc2_fpga0, tx_swap_mask_fmc2_fpga1);  

  type map_fpga_to_bank_position_t is array (0 to num_fpga_for_each_mainfpga-1) of bank_position_map_from_fpga_t;
  constant bank_position_in_fpga : map_fpga_to_bank_position_t := 
    (bank_position_fmc1_fpga0, bank_position_fmc1_fpga1, bank_position_fmc2_fpga0, bank_position_fmc2_fpga1);
  
  constant IsSctFIFO : integer := 1;
  constant IsPixFIFO : integer := 0;
  
  type rx_fmc_to_fpga_bit_channel_mapping is array(0 to num_fpga_per_fmc-1) of rx_fmc_to_fpga_bit_mapping_array_t;
  constant rx_fmc_to_fpgas_bit_mapping_in_all_FMC_LA_pin_count : rx_fmc_to_fpga_bit_channel_mapping
    := (rx_fmc_to_fpga0_bit_mapping_in_all_FMC_LA_pin_count,
        rx_fmc_to_fpga1_bit_mapping_in_all_FMC_LA_pin_count);
  type tx_fmc_to_fpga_bit_channel_mapping is array(0 to num_fpga_per_fmc-1) of tx_fmc_to_fpga_bit_mapping_array_t;  
  constant tx_fmc_to_fpgas_bit_mapping_in_all_FMC_LA_pin_count : tx_fmc_to_fpga_bit_channel_mapping
    := (tx_fmc_to_fpga0_bit_mapping_in_all_FMC_LA_pin_count,
        tx_fmc_to_fpga1_bit_mapping_in_all_FMC_LA_pin_count);

  constant swap_mask_test_mezzanine_la : std_logic_vector(total_low_pin_count_fmc-1 downto 0) :=
    "0100"&       -- LA33 - LA30 @ mezzanine
    "1000010001"& -- LA29 - LA20 @ mezzanine
    "0101011011"& -- LA19 - LA10 @ mezzanine
    "1101101010"; -- LA09 - LA00 @ mezzanine
  
  constant swap_mask_test_mezzanine_clk : std_logic_vector(num_fpga_per_fmc-1 downto 0) := "00";

  type swap_mask_for_total_low_pin_count is array(0 to num_fmc_per_mainfpga-1) of std_logic_vector(total_low_pin_count_fmc-1 downto 0);
  constant swap_mask_fmcs : swap_mask_for_total_low_pin_count := (swap_mask_fmc1, swap_mask_fmc2);
  
  constant fmc_phase_scan_pattern_id_for_normal_data    : integer := 0;
  constant fmc_phase_scan_pattern_id_for_test_pattern_1 : integer := 1;
  constant fmc_phase_scan_pattern_id_for_test_pattern_2 : integer := 2;

  constant FMC_BANK_IOSTANDARD : string := "LVDS";
  
end FmcConstants;


package body FmcConstants is
  -- ########################################################
  impure function ExtractFMCTXVectorComponent_FMCToFPGA (info               : in std_logic_vector;
                                                         bit_mapping_on_fmc : in tx_fmc_to_fpga_bit_mapping_array_t)
    return std_logic_vector is
    variable output_vector : std_logic_vector(lvds_pairs_for_tx_in_each_fpga-1 downto 0);
  begin
    for i in output_vector'range loop
      output_vector(i) := info(bit_mapping_on_fmc(i));
    end loop;
    return output_vector;
  end function;

-- ########################################################
  impure function ExtractFMCRXVectorComponent_FMCToFPGA (info               : in std_logic_vector;
                                                         bit_mapping_on_fmc : in rx_fmc_to_fpga_bit_mapping_array_t)
    return std_logic_vector is
    variable output_vector : std_logic_vector(lvds_pairs_for_rx_in_each_fpga-1 downto 0);
  begin
    for i in output_vector'range loop
      output_vector(i) := info(bit_mapping_on_fmc(i));
    end loop;
    return output_vector;
  end function;
  
  -- ########################################################  
  impure function ExtractFMCRXBankPosition_FMCToFPGA (info               : in bank_position_map_from_fmc_t;
                                                      bit_mapping_on_fmc : in rx_fmc_to_fpga_bit_mapping_array_t)
    return bank_position_map_from_fpga_t is
    variable output_vector : bank_position_map_from_fpga_t;
  begin
    for i in output_vector'range loop
      output_vector(i) := info(bit_mapping_on_fmc(i));
    end loop;
    return output_vector;
  end function;
    
end package body;
